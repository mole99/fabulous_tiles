magic
tech ihp-sg13g2
magscale 1 2
timestamp 1743695088
<< metal1 >>
rect 1152 10604 38112 10628
rect 1152 10564 4928 10604
rect 4968 10564 5010 10604
rect 5050 10564 5092 10604
rect 5132 10564 5174 10604
rect 5214 10564 5256 10604
rect 5296 10564 20048 10604
rect 20088 10564 20130 10604
rect 20170 10564 20212 10604
rect 20252 10564 20294 10604
rect 20334 10564 20376 10604
rect 20416 10564 35168 10604
rect 35208 10564 35250 10604
rect 35290 10564 35332 10604
rect 35372 10564 35414 10604
rect 35454 10564 35496 10604
rect 35536 10564 38112 10604
rect 1152 10540 38112 10564
rect 2235 10436 2277 10445
rect 2235 10396 2236 10436
rect 2276 10396 2277 10436
rect 2235 10387 2277 10396
rect 3963 10436 4005 10445
rect 3963 10396 3964 10436
rect 4004 10396 4005 10436
rect 3963 10387 4005 10396
rect 5691 10436 5733 10445
rect 5691 10396 5692 10436
rect 5732 10396 5733 10436
rect 5691 10387 5733 10396
rect 7419 10436 7461 10445
rect 7419 10396 7420 10436
rect 7460 10396 7461 10436
rect 7419 10387 7461 10396
rect 9147 10436 9189 10445
rect 9147 10396 9148 10436
rect 9188 10396 9189 10436
rect 9147 10387 9189 10396
rect 10875 10436 10917 10445
rect 10875 10396 10876 10436
rect 10916 10396 10917 10436
rect 10875 10387 10917 10396
rect 12603 10436 12645 10445
rect 12603 10396 12604 10436
rect 12644 10396 12645 10436
rect 12603 10387 12645 10396
rect 14331 10436 14373 10445
rect 14331 10396 14332 10436
rect 14372 10396 14373 10436
rect 14331 10387 14373 10396
rect 16059 10436 16101 10445
rect 16059 10396 16060 10436
rect 16100 10396 16101 10436
rect 16059 10387 16101 10396
rect 17787 10436 17829 10445
rect 17787 10396 17788 10436
rect 17828 10396 17829 10436
rect 17787 10387 17829 10396
rect 19515 10436 19557 10445
rect 19515 10396 19516 10436
rect 19556 10396 19557 10436
rect 19515 10387 19557 10396
rect 21243 10436 21285 10445
rect 21243 10396 21244 10436
rect 21284 10396 21285 10436
rect 21243 10387 21285 10396
rect 22971 10436 23013 10445
rect 22971 10396 22972 10436
rect 23012 10396 23013 10436
rect 22971 10387 23013 10396
rect 24699 10436 24741 10445
rect 24699 10396 24700 10436
rect 24740 10396 24741 10436
rect 24699 10387 24741 10396
rect 26427 10436 26469 10445
rect 26427 10396 26428 10436
rect 26468 10396 26469 10436
rect 26427 10387 26469 10396
rect 28155 10436 28197 10445
rect 28155 10396 28156 10436
rect 28196 10396 28197 10436
rect 28155 10387 28197 10396
rect 29883 10436 29925 10445
rect 29883 10396 29884 10436
rect 29924 10396 29925 10436
rect 29883 10387 29925 10396
rect 31611 10436 31653 10445
rect 31611 10396 31612 10436
rect 31652 10396 31653 10436
rect 31611 10387 31653 10396
rect 33339 10436 33381 10445
rect 33339 10396 33340 10436
rect 33380 10396 33381 10436
rect 33339 10387 33381 10396
rect 35067 10436 35109 10445
rect 35067 10396 35068 10436
rect 35108 10396 35109 10436
rect 35067 10387 35109 10396
rect 36315 10436 36357 10445
rect 36315 10396 36316 10436
rect 36356 10396 36357 10436
rect 36315 10387 36357 10396
rect 36795 10436 36837 10445
rect 36795 10396 36796 10436
rect 36836 10396 36837 10436
rect 36795 10387 36837 10396
rect 2475 10184 2517 10193
rect 2475 10144 2476 10184
rect 2516 10144 2517 10184
rect 2475 10135 2517 10144
rect 4203 10184 4245 10193
rect 4203 10144 4204 10184
rect 4244 10144 4245 10184
rect 4203 10135 4245 10144
rect 5931 10184 5973 10193
rect 5931 10144 5932 10184
rect 5972 10144 5973 10184
rect 5931 10135 5973 10144
rect 7659 10184 7701 10193
rect 7659 10144 7660 10184
rect 7700 10144 7701 10184
rect 7659 10135 7701 10144
rect 9387 10184 9429 10193
rect 9387 10144 9388 10184
rect 9428 10144 9429 10184
rect 9387 10135 9429 10144
rect 11115 10184 11157 10193
rect 11115 10144 11116 10184
rect 11156 10144 11157 10184
rect 11115 10135 11157 10144
rect 12843 10184 12885 10193
rect 12843 10144 12844 10184
rect 12884 10144 12885 10184
rect 12843 10135 12885 10144
rect 14571 10184 14613 10193
rect 14571 10144 14572 10184
rect 14612 10144 14613 10184
rect 14571 10135 14613 10144
rect 16299 10184 16341 10193
rect 16299 10144 16300 10184
rect 16340 10144 16341 10184
rect 16299 10135 16341 10144
rect 18027 10184 18069 10193
rect 18027 10144 18028 10184
rect 18068 10144 18069 10184
rect 18027 10135 18069 10144
rect 19803 10184 19845 10193
rect 19803 10144 19804 10184
rect 19844 10144 19845 10184
rect 19803 10135 19845 10144
rect 21483 10184 21525 10193
rect 21483 10144 21484 10184
rect 21524 10144 21525 10184
rect 21483 10135 21525 10144
rect 23211 10184 23253 10193
rect 23211 10144 23212 10184
rect 23252 10144 23253 10184
rect 23211 10135 23253 10144
rect 24939 10184 24981 10193
rect 24939 10144 24940 10184
rect 24980 10144 24981 10184
rect 24939 10135 24981 10144
rect 26667 10184 26709 10193
rect 26667 10144 26668 10184
rect 26708 10144 26709 10184
rect 26667 10135 26709 10144
rect 28395 10184 28437 10193
rect 28395 10144 28396 10184
rect 28436 10144 28437 10184
rect 28395 10135 28437 10144
rect 30123 10184 30165 10193
rect 30123 10144 30124 10184
rect 30164 10144 30165 10184
rect 30123 10135 30165 10144
rect 31851 10184 31893 10193
rect 31851 10144 31852 10184
rect 31892 10144 31893 10184
rect 31851 10135 31893 10144
rect 33579 10184 33621 10193
rect 33579 10144 33580 10184
rect 33620 10144 33621 10184
rect 33579 10135 33621 10144
rect 35307 10184 35349 10193
rect 35307 10144 35308 10184
rect 35348 10144 35349 10184
rect 35307 10135 35349 10144
rect 36075 10184 36117 10193
rect 36075 10144 36076 10184
rect 36116 10144 36117 10184
rect 36075 10135 36117 10144
rect 36459 10184 36501 10193
rect 36459 10144 36460 10184
rect 36500 10144 36501 10184
rect 36459 10135 36501 10144
rect 37035 10184 37077 10193
rect 37035 10144 37036 10184
rect 37076 10144 37077 10184
rect 37035 10135 37077 10144
rect 37419 10184 37461 10193
rect 37419 10144 37420 10184
rect 37460 10144 37461 10184
rect 37419 10135 37461 10144
rect 37803 10184 37845 10193
rect 37803 10144 37804 10184
rect 37844 10144 37845 10184
rect 37803 10135 37845 10144
rect 36699 10100 36741 10109
rect 36699 10060 36700 10100
rect 36740 10060 36741 10100
rect 36699 10051 36741 10060
rect 37659 10016 37701 10025
rect 37659 9976 37660 10016
rect 37700 9976 37701 10016
rect 37659 9967 37701 9976
rect 38043 10016 38085 10025
rect 38043 9976 38044 10016
rect 38084 9976 38085 10016
rect 38043 9967 38085 9976
rect 1152 9848 38112 9872
rect 1152 9808 3688 9848
rect 3728 9808 3770 9848
rect 3810 9808 3852 9848
rect 3892 9808 3934 9848
rect 3974 9808 4016 9848
rect 4056 9808 18808 9848
rect 18848 9808 18890 9848
rect 18930 9808 18972 9848
rect 19012 9808 19054 9848
rect 19094 9808 19136 9848
rect 19176 9808 33928 9848
rect 33968 9808 34010 9848
rect 34050 9808 34092 9848
rect 34132 9808 34174 9848
rect 34214 9808 34256 9848
rect 34296 9808 38112 9848
rect 1152 9784 38112 9808
rect 36891 9680 36933 9689
rect 36891 9640 36892 9680
rect 36932 9640 36933 9680
rect 36891 9631 36933 9640
rect 37275 9680 37317 9689
rect 37275 9640 37276 9680
rect 37316 9640 37317 9680
rect 37275 9631 37317 9640
rect 36651 9512 36693 9521
rect 36651 9472 36652 9512
rect 36692 9472 36693 9512
rect 36651 9463 36693 9472
rect 37035 9512 37077 9521
rect 37035 9472 37036 9512
rect 37076 9472 37077 9512
rect 37035 9463 37077 9472
rect 37419 9512 37461 9521
rect 37419 9472 37420 9512
rect 37460 9472 37461 9512
rect 37419 9463 37461 9472
rect 37803 9512 37845 9521
rect 37803 9472 37804 9512
rect 37844 9472 37845 9512
rect 37803 9463 37845 9472
rect 37659 9260 37701 9269
rect 37659 9220 37660 9260
rect 37700 9220 37701 9260
rect 37659 9211 37701 9220
rect 38043 9260 38085 9269
rect 38043 9220 38044 9260
rect 38084 9220 38085 9260
rect 38043 9211 38085 9220
rect 1152 9092 38112 9116
rect 1152 9052 4928 9092
rect 4968 9052 5010 9092
rect 5050 9052 5092 9092
rect 5132 9052 5174 9092
rect 5214 9052 5256 9092
rect 5296 9052 20048 9092
rect 20088 9052 20130 9092
rect 20170 9052 20212 9092
rect 20252 9052 20294 9092
rect 20334 9052 20376 9092
rect 20416 9052 35168 9092
rect 35208 9052 35250 9092
rect 35290 9052 35332 9092
rect 35372 9052 35414 9092
rect 35454 9052 35496 9092
rect 35536 9052 38112 9092
rect 1152 9028 38112 9052
rect 5499 8924 5541 8933
rect 5499 8884 5500 8924
rect 5540 8884 5541 8924
rect 5499 8875 5541 8884
rect 6651 8924 6693 8933
rect 6651 8884 6652 8924
rect 6692 8884 6693 8924
rect 6651 8875 6693 8884
rect 8187 8924 8229 8933
rect 8187 8884 8188 8924
rect 8228 8884 8229 8924
rect 8187 8875 8229 8884
rect 16923 8924 16965 8933
rect 16923 8884 16924 8924
rect 16964 8884 16965 8924
rect 16923 8875 16965 8884
rect 17883 8924 17925 8933
rect 17883 8884 17884 8924
rect 17924 8884 17925 8924
rect 17883 8875 17925 8884
rect 18747 8924 18789 8933
rect 18747 8884 18748 8924
rect 18788 8884 18789 8924
rect 18747 8875 18789 8884
rect 20091 8924 20133 8933
rect 20091 8884 20092 8924
rect 20132 8884 20133 8924
rect 20091 8875 20133 8884
rect 28251 8924 28293 8933
rect 28251 8884 28252 8924
rect 28292 8884 28293 8924
rect 28251 8875 28293 8884
rect 13083 8840 13125 8849
rect 13083 8800 13084 8840
rect 13124 8800 13125 8840
rect 13083 8791 13125 8800
rect 14907 8840 14949 8849
rect 14907 8800 14908 8840
rect 14948 8800 14949 8840
rect 14907 8791 14949 8800
rect 15291 8840 15333 8849
rect 15291 8800 15292 8840
rect 15332 8800 15333 8840
rect 15291 8791 15333 8800
rect 16827 8840 16869 8849
rect 16827 8800 16828 8840
rect 16868 8800 16869 8840
rect 16827 8791 16869 8800
rect 18363 8840 18405 8849
rect 18363 8800 18364 8840
rect 18404 8800 18405 8840
rect 18363 8791 18405 8800
rect 22683 8840 22725 8849
rect 22683 8800 22684 8840
rect 22724 8800 22725 8840
rect 22683 8791 22725 8800
rect 5259 8672 5301 8681
rect 5259 8632 5260 8672
rect 5300 8632 5301 8672
rect 5259 8623 5301 8632
rect 6411 8672 6453 8681
rect 6411 8632 6412 8672
rect 6452 8632 6453 8672
rect 6411 8623 6453 8632
rect 7947 8672 7989 8681
rect 7947 8632 7948 8672
rect 7988 8632 7989 8672
rect 7947 8623 7989 8632
rect 12843 8672 12885 8681
rect 12843 8632 12844 8672
rect 12884 8632 12885 8672
rect 12843 8623 12885 8632
rect 13227 8672 13269 8681
rect 13227 8632 13228 8672
rect 13268 8632 13269 8672
rect 13227 8623 13269 8632
rect 13899 8672 13941 8681
rect 13899 8632 13900 8672
rect 13940 8632 13941 8672
rect 13899 8623 13941 8632
rect 14139 8672 14181 8681
rect 14139 8632 14140 8672
rect 14180 8632 14181 8672
rect 14139 8623 14181 8632
rect 14667 8672 14709 8681
rect 14667 8632 14668 8672
rect 14708 8632 14709 8672
rect 14667 8623 14709 8632
rect 15051 8672 15093 8681
rect 15051 8632 15052 8672
rect 15092 8632 15093 8672
rect 15051 8623 15093 8632
rect 15531 8672 15573 8681
rect 15531 8632 15532 8672
rect 15572 8632 15573 8672
rect 15531 8623 15573 8632
rect 15771 8672 15813 8681
rect 15771 8632 15772 8672
rect 15812 8632 15813 8672
rect 15771 8623 15813 8632
rect 16587 8672 16629 8681
rect 16587 8632 16588 8672
rect 16628 8632 16629 8672
rect 16587 8623 16629 8632
rect 17163 8672 17205 8681
rect 17163 8632 17164 8672
rect 17204 8632 17205 8672
rect 17163 8623 17205 8632
rect 17643 8672 17685 8681
rect 17643 8632 17644 8672
rect 17684 8632 17685 8672
rect 17643 8623 17685 8632
rect 18123 8672 18165 8681
rect 18123 8632 18124 8672
rect 18164 8632 18165 8672
rect 18123 8623 18165 8632
rect 18507 8672 18549 8681
rect 18507 8632 18508 8672
rect 18548 8632 18549 8672
rect 18507 8623 18549 8632
rect 18987 8672 19029 8681
rect 18987 8632 18988 8672
rect 19028 8632 19029 8672
rect 18987 8623 19029 8632
rect 19227 8672 19269 8681
rect 19227 8632 19228 8672
rect 19268 8632 19269 8672
rect 19227 8623 19269 8632
rect 19498 8672 19556 8673
rect 19498 8632 19507 8672
rect 19547 8632 19556 8672
rect 19498 8631 19556 8632
rect 19882 8672 19940 8673
rect 19882 8632 19891 8672
rect 19931 8632 19940 8672
rect 19882 8631 19940 8632
rect 20523 8672 20565 8681
rect 20523 8632 20524 8672
rect 20564 8632 20565 8672
rect 20523 8623 20565 8632
rect 20907 8672 20949 8681
rect 20907 8632 20908 8672
rect 20948 8632 20949 8672
rect 20907 8623 20949 8632
rect 21147 8672 21189 8681
rect 21147 8632 21148 8672
rect 21188 8632 21189 8672
rect 21147 8623 21189 8632
rect 21771 8672 21813 8681
rect 21771 8632 21772 8672
rect 21812 8632 21813 8672
rect 21771 8623 21813 8632
rect 22923 8672 22965 8681
rect 22923 8632 22924 8672
rect 22964 8632 22965 8672
rect 22923 8623 22965 8632
rect 24315 8672 24357 8681
rect 24315 8632 24316 8672
rect 24356 8632 24357 8672
rect 24315 8623 24357 8632
rect 24555 8672 24597 8681
rect 24555 8632 24556 8672
rect 24596 8632 24597 8672
rect 24555 8623 24597 8632
rect 25131 8672 25173 8681
rect 25131 8632 25132 8672
rect 25172 8632 25173 8672
rect 25131 8623 25173 8632
rect 25371 8672 25413 8681
rect 25371 8632 25372 8672
rect 25412 8632 25413 8672
rect 25371 8623 25413 8632
rect 25803 8672 25845 8681
rect 25803 8632 25804 8672
rect 25844 8632 25845 8672
rect 25803 8623 25845 8632
rect 27435 8672 27477 8681
rect 27435 8632 27436 8672
rect 27476 8632 27477 8672
rect 27435 8623 27477 8632
rect 27819 8672 27861 8681
rect 27819 8632 27820 8672
rect 27860 8632 27861 8672
rect 27819 8623 27861 8632
rect 28042 8672 28100 8673
rect 28042 8632 28051 8672
rect 28091 8632 28100 8672
rect 28042 8631 28100 8632
rect 29067 8672 29109 8681
rect 29067 8632 29068 8672
rect 29108 8632 29109 8672
rect 29067 8623 29109 8632
rect 29307 8672 29349 8681
rect 29307 8632 29308 8672
rect 29348 8632 29349 8672
rect 29307 8623 29349 8632
rect 37419 8672 37461 8681
rect 37419 8632 37420 8672
rect 37460 8632 37461 8672
rect 37419 8623 37461 8632
rect 37803 8672 37845 8681
rect 37803 8632 37804 8672
rect 37844 8632 37845 8672
rect 37803 8623 37845 8632
rect 38043 8672 38085 8681
rect 38043 8632 38044 8672
rect 38084 8632 38085 8672
rect 38043 8623 38085 8632
rect 20763 8588 20805 8597
rect 20763 8548 20764 8588
rect 20804 8548 20805 8588
rect 20763 8539 20805 8548
rect 25563 8588 25605 8597
rect 25563 8548 25564 8588
rect 25604 8548 25605 8588
rect 25563 8539 25605 8548
rect 27195 8588 27237 8597
rect 27195 8548 27196 8588
rect 27236 8548 27237 8588
rect 27195 8539 27237 8548
rect 27579 8588 27621 8597
rect 27579 8548 27580 8588
rect 27620 8548 27621 8588
rect 27579 8539 27621 8548
rect 37659 8588 37701 8597
rect 37659 8548 37660 8588
rect 37700 8548 37701 8588
rect 37659 8539 37701 8548
rect 13467 8504 13509 8513
rect 13467 8464 13468 8504
rect 13508 8464 13509 8504
rect 13467 8455 13509 8464
rect 19707 8504 19749 8513
rect 19707 8464 19708 8504
rect 19748 8464 19749 8504
rect 19707 8455 19749 8464
rect 22011 8504 22053 8513
rect 22011 8464 22012 8504
rect 22052 8464 22053 8504
rect 22011 8455 22053 8464
rect 1152 8336 38112 8360
rect 1152 8296 3688 8336
rect 3728 8296 3770 8336
rect 3810 8296 3852 8336
rect 3892 8296 3934 8336
rect 3974 8296 4016 8336
rect 4056 8296 18808 8336
rect 18848 8296 18890 8336
rect 18930 8296 18972 8336
rect 19012 8296 19054 8336
rect 19094 8296 19136 8336
rect 19176 8296 33928 8336
rect 33968 8296 34010 8336
rect 34050 8296 34092 8336
rect 34132 8296 34174 8336
rect 34214 8296 34256 8336
rect 34296 8296 38112 8336
rect 1152 8272 38112 8296
rect 29211 8168 29253 8177
rect 29211 8128 29212 8168
rect 29252 8128 29253 8168
rect 29211 8119 29253 8128
rect 10683 8084 10725 8093
rect 10683 8044 10684 8084
rect 10724 8044 10725 8084
rect 10683 8035 10725 8044
rect 11355 8084 11397 8093
rect 11355 8044 11356 8084
rect 11396 8044 11397 8084
rect 11355 8035 11397 8044
rect 10443 8000 10485 8009
rect 10443 7960 10444 8000
rect 10484 7960 10485 8000
rect 10443 7951 10485 7960
rect 11115 8000 11157 8009
rect 11115 7960 11116 8000
rect 11156 7960 11157 8000
rect 11115 7951 11157 7960
rect 11499 8000 11541 8009
rect 11499 7960 11500 8000
rect 11540 7960 11541 8000
rect 11499 7951 11541 7960
rect 29451 8000 29493 8009
rect 29451 7960 29452 8000
rect 29492 7960 29493 8000
rect 29451 7951 29493 7960
rect 37419 8000 37461 8009
rect 37419 7960 37420 8000
rect 37460 7960 37461 8000
rect 37419 7951 37461 7960
rect 37803 8000 37845 8009
rect 37803 7960 37804 8000
rect 37844 7960 37845 8000
rect 37803 7951 37845 7960
rect 37659 7832 37701 7841
rect 37659 7792 37660 7832
rect 37700 7792 37701 7832
rect 37659 7783 37701 7792
rect 11739 7748 11781 7757
rect 11739 7708 11740 7748
rect 11780 7708 11781 7748
rect 11739 7699 11781 7708
rect 38043 7748 38085 7757
rect 38043 7708 38044 7748
rect 38084 7708 38085 7748
rect 38043 7699 38085 7708
rect 1152 7580 38112 7604
rect 1152 7540 4928 7580
rect 4968 7540 5010 7580
rect 5050 7540 5092 7580
rect 5132 7540 5174 7580
rect 5214 7540 5256 7580
rect 5296 7540 20048 7580
rect 20088 7540 20130 7580
rect 20170 7540 20212 7580
rect 20252 7540 20294 7580
rect 20334 7540 20376 7580
rect 20416 7540 35168 7580
rect 35208 7540 35250 7580
rect 35290 7540 35332 7580
rect 35372 7540 35414 7580
rect 35454 7540 35496 7580
rect 35536 7540 38112 7580
rect 1152 7516 38112 7540
rect 6027 7160 6069 7169
rect 6027 7120 6028 7160
rect 6068 7120 6069 7160
rect 6027 7111 6069 7120
rect 37419 7160 37461 7169
rect 37419 7120 37420 7160
rect 37460 7120 37461 7160
rect 37419 7111 37461 7120
rect 37803 7160 37845 7169
rect 37803 7120 37804 7160
rect 37844 7120 37845 7160
rect 37803 7111 37845 7120
rect 38043 7160 38085 7169
rect 38043 7120 38044 7160
rect 38084 7120 38085 7160
rect 38043 7111 38085 7120
rect 5787 7076 5829 7085
rect 5787 7036 5788 7076
rect 5828 7036 5829 7076
rect 5787 7027 5829 7036
rect 37659 6992 37701 7001
rect 37659 6952 37660 6992
rect 37700 6952 37701 6992
rect 37659 6943 37701 6952
rect 1152 6824 38112 6848
rect 1152 6784 3688 6824
rect 3728 6784 3770 6824
rect 3810 6784 3852 6824
rect 3892 6784 3934 6824
rect 3974 6784 4016 6824
rect 4056 6784 18808 6824
rect 18848 6784 18890 6824
rect 18930 6784 18972 6824
rect 19012 6784 19054 6824
rect 19094 6784 19136 6824
rect 19176 6784 33928 6824
rect 33968 6784 34010 6824
rect 34050 6784 34092 6824
rect 34132 6784 34174 6824
rect 34214 6784 34256 6824
rect 34296 6784 38112 6824
rect 1152 6760 38112 6784
rect 2619 6656 2661 6665
rect 2619 6616 2620 6656
rect 2660 6616 2661 6656
rect 2619 6607 2661 6616
rect 27483 6656 27525 6665
rect 27483 6616 27484 6656
rect 27524 6616 27525 6656
rect 27483 6607 27525 6616
rect 2859 6488 2901 6497
rect 2859 6448 2860 6488
rect 2900 6448 2901 6488
rect 2859 6439 2901 6448
rect 27723 6488 27765 6497
rect 27723 6448 27724 6488
rect 27764 6448 27765 6488
rect 27723 6439 27765 6448
rect 31467 6488 31509 6497
rect 31467 6448 31468 6488
rect 31508 6448 31509 6488
rect 31467 6439 31509 6448
rect 37419 6488 37461 6497
rect 37419 6448 37420 6488
rect 37460 6448 37461 6488
rect 37419 6439 37461 6448
rect 37803 6488 37845 6497
rect 37803 6448 37804 6488
rect 37844 6448 37845 6488
rect 37803 6439 37845 6448
rect 38043 6488 38085 6497
rect 38043 6448 38044 6488
rect 38084 6448 38085 6488
rect 38043 6439 38085 6448
rect 31707 6236 31749 6245
rect 31707 6196 31708 6236
rect 31748 6196 31749 6236
rect 31707 6187 31749 6196
rect 37659 6236 37701 6245
rect 37659 6196 37660 6236
rect 37700 6196 37701 6236
rect 37659 6187 37701 6196
rect 1152 6068 38112 6092
rect 1152 6028 4928 6068
rect 4968 6028 5010 6068
rect 5050 6028 5092 6068
rect 5132 6028 5174 6068
rect 5214 6028 5256 6068
rect 5296 6028 20048 6068
rect 20088 6028 20130 6068
rect 20170 6028 20212 6068
rect 20252 6028 20294 6068
rect 20334 6028 20376 6068
rect 20416 6028 35168 6068
rect 35208 6028 35250 6068
rect 35290 6028 35332 6068
rect 35372 6028 35414 6068
rect 35454 6028 35496 6068
rect 35536 6028 38112 6068
rect 1152 6004 38112 6028
rect 38043 5816 38085 5825
rect 38043 5776 38044 5816
rect 38084 5776 38085 5816
rect 38043 5767 38085 5776
rect 2667 5648 2709 5657
rect 2667 5608 2668 5648
rect 2708 5608 2709 5648
rect 2667 5599 2709 5608
rect 2907 5648 2949 5657
rect 2907 5608 2908 5648
rect 2948 5608 2949 5648
rect 2907 5599 2949 5608
rect 37419 5648 37461 5657
rect 37419 5608 37420 5648
rect 37460 5608 37461 5648
rect 37419 5599 37461 5608
rect 37803 5648 37845 5657
rect 37803 5608 37804 5648
rect 37844 5608 37845 5648
rect 37803 5599 37845 5608
rect 37659 5564 37701 5573
rect 37659 5524 37660 5564
rect 37700 5524 37701 5564
rect 37659 5515 37701 5524
rect 1152 5312 38112 5336
rect 1152 5272 3688 5312
rect 3728 5272 3770 5312
rect 3810 5272 3852 5312
rect 3892 5272 3934 5312
rect 3974 5272 4016 5312
rect 4056 5272 18808 5312
rect 18848 5272 18890 5312
rect 18930 5272 18972 5312
rect 19012 5272 19054 5312
rect 19094 5272 19136 5312
rect 19176 5272 33928 5312
rect 33968 5272 34010 5312
rect 34050 5272 34092 5312
rect 34132 5272 34174 5312
rect 34214 5272 34256 5312
rect 34296 5272 38112 5312
rect 1152 5248 38112 5272
rect 7899 5144 7941 5153
rect 7899 5104 7900 5144
rect 7940 5104 7941 5144
rect 7899 5095 7941 5104
rect 8379 5144 8421 5153
rect 8379 5104 8380 5144
rect 8420 5104 8421 5144
rect 8379 5095 8421 5104
rect 10395 5144 10437 5153
rect 10395 5104 10396 5144
rect 10436 5104 10437 5144
rect 10395 5095 10437 5104
rect 27867 5144 27909 5153
rect 27867 5104 27868 5144
rect 27908 5104 27909 5144
rect 27867 5095 27909 5104
rect 33627 5144 33669 5153
rect 33627 5104 33628 5144
rect 33668 5104 33669 5144
rect 33627 5095 33669 5104
rect 38043 5144 38085 5153
rect 38043 5104 38044 5144
rect 38084 5104 38085 5144
rect 38043 5095 38085 5104
rect 16251 5060 16293 5069
rect 16251 5020 16252 5060
rect 16292 5020 16293 5060
rect 16251 5011 16293 5020
rect 7275 4976 7317 4985
rect 7275 4936 7276 4976
rect 7316 4936 7317 4976
rect 7275 4927 7317 4936
rect 7659 4976 7701 4985
rect 7659 4936 7660 4976
rect 7700 4936 7701 4976
rect 7659 4927 7701 4936
rect 8139 4976 8181 4985
rect 8139 4936 8140 4976
rect 8180 4936 8181 4976
rect 8139 4927 8181 4936
rect 8523 4976 8565 4985
rect 8523 4936 8524 4976
rect 8564 4936 8565 4976
rect 8523 4927 8565 4936
rect 8907 4976 8949 4985
rect 8907 4936 8908 4976
rect 8948 4936 8949 4976
rect 8907 4927 8949 4936
rect 9291 4976 9333 4985
rect 9291 4936 9292 4976
rect 9332 4936 9333 4976
rect 9291 4927 9333 4936
rect 9771 4976 9813 4985
rect 9771 4936 9772 4976
rect 9812 4936 9813 4976
rect 9771 4927 9813 4936
rect 10155 4976 10197 4985
rect 10155 4936 10156 4976
rect 10196 4936 10197 4976
rect 10155 4927 10197 4936
rect 13131 4976 13173 4985
rect 13131 4936 13132 4976
rect 13172 4936 13173 4976
rect 13131 4927 13173 4936
rect 13371 4976 13413 4985
rect 13371 4936 13372 4976
rect 13412 4936 13413 4976
rect 13371 4927 13413 4936
rect 16011 4976 16053 4985
rect 16011 4936 16012 4976
rect 16052 4936 16053 4976
rect 16011 4927 16053 4936
rect 17067 4976 17109 4985
rect 17067 4936 17068 4976
rect 17108 4936 17109 4976
rect 17067 4927 17109 4936
rect 17643 4976 17685 4985
rect 17643 4936 17644 4976
rect 17684 4936 17685 4976
rect 17643 4927 17685 4936
rect 18027 4976 18069 4985
rect 18027 4936 18028 4976
rect 18068 4936 18069 4976
rect 18027 4927 18069 4936
rect 21963 4976 22005 4985
rect 21963 4936 21964 4976
rect 22004 4936 22005 4976
rect 21963 4927 22005 4936
rect 22347 4976 22389 4985
rect 22347 4936 22348 4976
rect 22388 4936 22389 4976
rect 22347 4927 22389 4936
rect 25707 4976 25749 4985
rect 25707 4936 25708 4976
rect 25748 4936 25749 4976
rect 25707 4927 25749 4936
rect 26187 4976 26229 4985
rect 26187 4936 26188 4976
rect 26228 4936 26229 4976
rect 26187 4927 26229 4936
rect 28107 4976 28149 4985
rect 28107 4936 28108 4976
rect 28148 4936 28149 4976
rect 28107 4927 28149 4936
rect 31275 4976 31317 4985
rect 31275 4936 31276 4976
rect 31316 4936 31317 4976
rect 31275 4927 31317 4936
rect 33387 4976 33429 4985
rect 33387 4936 33388 4976
rect 33428 4936 33429 4976
rect 33387 4927 33429 4936
rect 37419 4976 37461 4985
rect 37419 4936 37420 4976
rect 37460 4936 37461 4976
rect 37419 4927 37461 4936
rect 37803 4976 37845 4985
rect 37803 4936 37804 4976
rect 37844 4936 37845 4976
rect 37803 4927 37845 4936
rect 10011 4808 10053 4817
rect 10011 4768 10012 4808
rect 10052 4768 10053 4808
rect 10011 4759 10053 4768
rect 37659 4808 37701 4817
rect 37659 4768 37660 4808
rect 37700 4768 37701 4808
rect 37659 4759 37701 4768
rect 7515 4724 7557 4733
rect 7515 4684 7516 4724
rect 7556 4684 7557 4724
rect 7515 4675 7557 4684
rect 8763 4724 8805 4733
rect 8763 4684 8764 4724
rect 8804 4684 8805 4724
rect 8763 4675 8805 4684
rect 9147 4724 9189 4733
rect 9147 4684 9148 4724
rect 9188 4684 9189 4724
rect 9147 4675 9189 4684
rect 9531 4724 9573 4733
rect 9531 4684 9532 4724
rect 9572 4684 9573 4724
rect 9531 4675 9573 4684
rect 17307 4724 17349 4733
rect 17307 4684 17308 4724
rect 17348 4684 17349 4724
rect 17307 4675 17349 4684
rect 17883 4724 17925 4733
rect 17883 4684 17884 4724
rect 17924 4684 17925 4724
rect 17883 4675 17925 4684
rect 18267 4724 18309 4733
rect 18267 4684 18268 4724
rect 18308 4684 18309 4724
rect 18267 4675 18309 4684
rect 22203 4724 22245 4733
rect 22203 4684 22204 4724
rect 22244 4684 22245 4724
rect 22203 4675 22245 4684
rect 22587 4724 22629 4733
rect 22587 4684 22588 4724
rect 22628 4684 22629 4724
rect 22587 4675 22629 4684
rect 25947 4724 25989 4733
rect 25947 4684 25948 4724
rect 25988 4684 25989 4724
rect 25947 4675 25989 4684
rect 26427 4724 26469 4733
rect 26427 4684 26428 4724
rect 26468 4684 26469 4724
rect 26427 4675 26469 4684
rect 31515 4724 31557 4733
rect 31515 4684 31516 4724
rect 31556 4684 31557 4724
rect 31515 4675 31557 4684
rect 1152 4556 38112 4580
rect 1152 4516 4928 4556
rect 4968 4516 5010 4556
rect 5050 4516 5092 4556
rect 5132 4516 5174 4556
rect 5214 4516 5256 4556
rect 5296 4516 20048 4556
rect 20088 4516 20130 4556
rect 20170 4516 20212 4556
rect 20252 4516 20294 4556
rect 20334 4516 20376 4556
rect 20416 4516 35168 4556
rect 35208 4516 35250 4556
rect 35290 4516 35332 4556
rect 35372 4516 35414 4556
rect 35454 4516 35496 4556
rect 35536 4516 38112 4556
rect 1152 4492 38112 4516
rect 26139 4388 26181 4397
rect 26139 4348 26140 4388
rect 26180 4348 26181 4388
rect 26139 4339 26181 4348
rect 13275 4304 13317 4313
rect 13275 4264 13276 4304
rect 13316 4264 13317 4304
rect 13275 4255 13317 4264
rect 18651 4304 18693 4313
rect 18651 4264 18652 4304
rect 18692 4264 18693 4304
rect 18651 4255 18693 4264
rect 22491 4304 22533 4313
rect 22491 4264 22492 4304
rect 22532 4264 22533 4304
rect 22491 4255 22533 4264
rect 23643 4304 23685 4313
rect 23643 4264 23644 4304
rect 23684 4264 23685 4304
rect 23643 4255 23685 4264
rect 32475 4304 32517 4313
rect 32475 4264 32476 4304
rect 32516 4264 32517 4304
rect 32475 4255 32517 4264
rect 32859 4304 32901 4313
rect 32859 4264 32860 4304
rect 32900 4264 32901 4304
rect 32859 4255 32901 4264
rect 38043 4304 38085 4313
rect 38043 4264 38044 4304
rect 38084 4264 38085 4304
rect 38043 4255 38085 4264
rect 8235 4136 8277 4145
rect 8235 4096 8236 4136
rect 8276 4096 8277 4136
rect 8235 4087 8277 4096
rect 8619 4136 8661 4145
rect 8619 4096 8620 4136
rect 8660 4096 8661 4136
rect 8619 4087 8661 4096
rect 9963 4136 10005 4145
rect 9963 4096 9964 4136
rect 10004 4096 10005 4136
rect 9963 4087 10005 4096
rect 10347 4136 10389 4145
rect 10347 4096 10348 4136
rect 10388 4096 10389 4136
rect 10347 4087 10389 4096
rect 11883 4136 11925 4145
rect 11883 4096 11884 4136
rect 11924 4096 11925 4136
rect 11883 4087 11925 4096
rect 12267 4136 12309 4145
rect 12267 4096 12268 4136
rect 12308 4096 12309 4136
rect 12267 4087 12309 4096
rect 12651 4136 12693 4145
rect 12651 4096 12652 4136
rect 12692 4096 12693 4136
rect 12651 4087 12693 4096
rect 13035 4136 13077 4145
rect 13035 4096 13036 4136
rect 13076 4096 13077 4136
rect 13035 4087 13077 4096
rect 13419 4136 13461 4145
rect 13419 4096 13420 4136
rect 13460 4096 13461 4136
rect 13419 4087 13461 4096
rect 13803 4136 13845 4145
rect 13803 4096 13804 4136
rect 13844 4096 13845 4136
rect 13803 4087 13845 4096
rect 14379 4136 14421 4145
rect 14379 4096 14380 4136
rect 14420 4096 14421 4136
rect 14379 4087 14421 4096
rect 16107 4136 16149 4145
rect 16107 4096 16108 4136
rect 16148 4096 16149 4136
rect 16107 4087 16149 4096
rect 16491 4136 16533 4145
rect 16491 4096 16492 4136
rect 16532 4096 16533 4136
rect 16491 4087 16533 4096
rect 16875 4136 16917 4145
rect 16875 4096 16876 4136
rect 16916 4096 16917 4136
rect 16875 4087 16917 4096
rect 17259 4136 17301 4145
rect 17259 4096 17260 4136
rect 17300 4096 17301 4136
rect 17259 4087 17301 4096
rect 17643 4136 17685 4145
rect 17643 4096 17644 4136
rect 17684 4096 17685 4136
rect 17643 4087 17685 4096
rect 18027 4136 18069 4145
rect 18027 4096 18028 4136
rect 18068 4096 18069 4136
rect 18027 4087 18069 4096
rect 18411 4136 18453 4145
rect 18411 4096 18412 4136
rect 18452 4096 18453 4136
rect 18411 4087 18453 4096
rect 18795 4136 18837 4145
rect 18795 4096 18796 4136
rect 18836 4096 18837 4136
rect 18795 4087 18837 4096
rect 19179 4136 19221 4145
rect 19179 4096 19180 4136
rect 19220 4096 19221 4136
rect 19179 4087 19221 4096
rect 19419 4136 19461 4145
rect 19419 4096 19420 4136
rect 19460 4096 19461 4136
rect 19419 4087 19461 4096
rect 19755 4136 19797 4145
rect 19755 4096 19756 4136
rect 19796 4096 19797 4136
rect 19755 4087 19797 4096
rect 21099 4136 21141 4145
rect 21099 4096 21100 4136
rect 21140 4096 21141 4136
rect 21099 4087 21141 4096
rect 21483 4136 21525 4145
rect 21483 4096 21484 4136
rect 21524 4096 21525 4136
rect 21483 4087 21525 4096
rect 21867 4136 21909 4145
rect 21867 4096 21868 4136
rect 21908 4096 21909 4136
rect 21867 4087 21909 4096
rect 22251 4136 22293 4145
rect 22251 4096 22252 4136
rect 22292 4096 22293 4136
rect 22251 4087 22293 4096
rect 22635 4136 22677 4145
rect 22635 4096 22636 4136
rect 22676 4096 22677 4136
rect 22635 4087 22677 4096
rect 23019 4136 23061 4145
rect 23019 4096 23020 4136
rect 23060 4096 23061 4136
rect 23019 4087 23061 4096
rect 23403 4136 23445 4145
rect 23403 4096 23404 4136
rect 23444 4096 23445 4136
rect 23403 4087 23445 4096
rect 23787 4136 23829 4145
rect 23787 4096 23788 4136
rect 23828 4096 23829 4136
rect 23787 4087 23829 4096
rect 24171 4136 24213 4145
rect 24171 4096 24172 4136
rect 24212 4096 24213 4136
rect 24171 4087 24213 4096
rect 25899 4136 25941 4145
rect 25899 4096 25900 4136
rect 25940 4096 25941 4136
rect 25899 4087 25941 4096
rect 27243 4136 27285 4145
rect 27243 4096 27244 4136
rect 27284 4096 27285 4136
rect 27243 4087 27285 4096
rect 28587 4136 28629 4145
rect 28587 4096 28588 4136
rect 28628 4096 28629 4136
rect 28587 4087 28629 4096
rect 29643 4136 29685 4145
rect 29643 4096 29644 4136
rect 29684 4096 29685 4136
rect 29643 4087 29685 4096
rect 31563 4136 31605 4145
rect 31563 4096 31564 4136
rect 31604 4096 31605 4136
rect 31563 4087 31605 4096
rect 32235 4136 32277 4145
rect 32235 4096 32236 4136
rect 32276 4096 32277 4136
rect 32235 4087 32277 4096
rect 32619 4136 32661 4145
rect 32619 4096 32620 4136
rect 32660 4096 32661 4136
rect 32619 4087 32661 4096
rect 33003 4136 33045 4145
rect 33003 4096 33004 4136
rect 33044 4096 33045 4136
rect 33003 4087 33045 4096
rect 37035 4136 37077 4145
rect 37035 4096 37036 4136
rect 37076 4096 37077 4136
rect 37035 4087 37077 4096
rect 37419 4136 37461 4145
rect 37419 4096 37420 4136
rect 37460 4096 37461 4136
rect 37419 4087 37461 4096
rect 37803 4136 37845 4145
rect 37803 4096 37804 4136
rect 37844 4096 37845 4136
rect 37803 4087 37845 4096
rect 12123 4052 12165 4061
rect 12123 4012 12124 4052
rect 12164 4012 12165 4052
rect 12123 4003 12165 4012
rect 14043 4052 14085 4061
rect 14043 4012 14044 4052
rect 14084 4012 14085 4052
rect 14043 4003 14085 4012
rect 14619 4052 14661 4061
rect 14619 4012 14620 4052
rect 14660 4012 14661 4052
rect 14619 4003 14661 4012
rect 24411 4052 24453 4061
rect 24411 4012 24412 4052
rect 24452 4012 24453 4052
rect 24411 4003 24453 4012
rect 31803 4052 31845 4061
rect 31803 4012 31804 4052
rect 31844 4012 31845 4052
rect 31803 4003 31845 4012
rect 33243 4052 33285 4061
rect 33243 4012 33244 4052
rect 33284 4012 33285 4052
rect 33243 4003 33285 4012
rect 37659 4052 37701 4061
rect 37659 4012 37660 4052
rect 37700 4012 37701 4052
rect 37659 4003 37701 4012
rect 8475 3968 8517 3977
rect 8475 3928 8476 3968
rect 8516 3928 8517 3968
rect 8475 3919 8517 3928
rect 8859 3968 8901 3977
rect 8859 3928 8860 3968
rect 8900 3928 8901 3968
rect 8859 3919 8901 3928
rect 10203 3968 10245 3977
rect 10203 3928 10204 3968
rect 10244 3928 10245 3968
rect 10203 3919 10245 3928
rect 10587 3968 10629 3977
rect 10587 3928 10588 3968
rect 10628 3928 10629 3968
rect 10587 3919 10629 3928
rect 12507 3968 12549 3977
rect 12507 3928 12508 3968
rect 12548 3928 12549 3968
rect 12507 3919 12549 3928
rect 12891 3968 12933 3977
rect 12891 3928 12892 3968
rect 12932 3928 12933 3968
rect 12891 3919 12933 3928
rect 13659 3968 13701 3977
rect 13659 3928 13660 3968
rect 13700 3928 13701 3968
rect 13659 3919 13701 3928
rect 16347 3968 16389 3977
rect 16347 3928 16348 3968
rect 16388 3928 16389 3968
rect 16347 3919 16389 3928
rect 16731 3968 16773 3977
rect 16731 3928 16732 3968
rect 16772 3928 16773 3968
rect 16731 3919 16773 3928
rect 17115 3968 17157 3977
rect 17115 3928 17116 3968
rect 17156 3928 17157 3968
rect 17115 3919 17157 3928
rect 17499 3968 17541 3977
rect 17499 3928 17500 3968
rect 17540 3928 17541 3968
rect 17499 3919 17541 3928
rect 17883 3968 17925 3977
rect 17883 3928 17884 3968
rect 17924 3928 17925 3968
rect 17883 3919 17925 3928
rect 18267 3968 18309 3977
rect 18267 3928 18268 3968
rect 18308 3928 18309 3968
rect 18267 3919 18309 3928
rect 19035 3968 19077 3977
rect 19035 3928 19036 3968
rect 19076 3928 19077 3968
rect 19035 3919 19077 3928
rect 19995 3968 20037 3977
rect 19995 3928 19996 3968
rect 20036 3928 20037 3968
rect 19995 3919 20037 3928
rect 21339 3968 21381 3977
rect 21339 3928 21340 3968
rect 21380 3928 21381 3968
rect 21339 3919 21381 3928
rect 21723 3968 21765 3977
rect 21723 3928 21724 3968
rect 21764 3928 21765 3968
rect 21723 3919 21765 3928
rect 22107 3968 22149 3977
rect 22107 3928 22108 3968
rect 22148 3928 22149 3968
rect 22107 3919 22149 3928
rect 22875 3968 22917 3977
rect 22875 3928 22876 3968
rect 22916 3928 22917 3968
rect 22875 3919 22917 3928
rect 23259 3968 23301 3977
rect 23259 3928 23260 3968
rect 23300 3928 23301 3968
rect 23259 3919 23301 3928
rect 24027 3968 24069 3977
rect 24027 3928 24028 3968
rect 24068 3928 24069 3968
rect 24027 3919 24069 3928
rect 27483 3968 27525 3977
rect 27483 3928 27484 3968
rect 27524 3928 27525 3968
rect 27483 3919 27525 3928
rect 28347 3968 28389 3977
rect 28347 3928 28348 3968
rect 28388 3928 28389 3968
rect 28347 3919 28389 3928
rect 29403 3968 29445 3977
rect 29403 3928 29404 3968
rect 29444 3928 29445 3968
rect 29403 3919 29445 3928
rect 37275 3968 37317 3977
rect 37275 3928 37276 3968
rect 37316 3928 37317 3968
rect 37275 3919 37317 3928
rect 1152 3800 38112 3824
rect 1152 3760 3688 3800
rect 3728 3760 3770 3800
rect 3810 3760 3852 3800
rect 3892 3760 3934 3800
rect 3974 3760 4016 3800
rect 4056 3760 18808 3800
rect 18848 3760 18890 3800
rect 18930 3760 18972 3800
rect 19012 3760 19054 3800
rect 19094 3760 19136 3800
rect 19176 3760 33928 3800
rect 33968 3760 34010 3800
rect 34050 3760 34092 3800
rect 34132 3760 34174 3800
rect 34214 3760 34256 3800
rect 34296 3760 38112 3800
rect 1152 3736 38112 3760
rect 27579 3632 27621 3641
rect 27579 3592 27580 3632
rect 27620 3592 27621 3632
rect 27579 3583 27621 3592
rect 28923 3632 28965 3641
rect 28923 3592 28924 3632
rect 28964 3592 28965 3632
rect 28923 3583 28965 3592
rect 30843 3632 30885 3641
rect 30843 3592 30844 3632
rect 30884 3592 30885 3632
rect 30843 3583 30885 3592
rect 31995 3632 32037 3641
rect 31995 3592 31996 3632
rect 32036 3592 32037 3632
rect 31995 3583 32037 3592
rect 38043 3632 38085 3641
rect 38043 3592 38044 3632
rect 38084 3592 38085 3632
rect 38043 3583 38085 3592
rect 13035 3464 13077 3473
rect 13035 3424 13036 3464
rect 13076 3424 13077 3464
rect 13035 3415 13077 3424
rect 13419 3464 13461 3473
rect 13419 3424 13420 3464
rect 13460 3424 13461 3464
rect 13419 3415 13461 3424
rect 13659 3464 13701 3473
rect 13659 3424 13660 3464
rect 13700 3424 13701 3464
rect 13659 3415 13701 3424
rect 17739 3464 17781 3473
rect 17739 3424 17740 3464
rect 17780 3424 17781 3464
rect 17739 3415 17781 3424
rect 18123 3464 18165 3473
rect 18123 3424 18124 3464
rect 18164 3424 18165 3464
rect 18123 3415 18165 3424
rect 21867 3464 21909 3473
rect 21867 3424 21868 3464
rect 21908 3424 21909 3464
rect 21867 3415 21909 3424
rect 22251 3464 22293 3473
rect 22251 3424 22252 3464
rect 22292 3424 22293 3464
rect 22251 3415 22293 3424
rect 27819 3464 27861 3473
rect 27819 3424 27820 3464
rect 27860 3424 27861 3464
rect 27819 3415 27861 3424
rect 29163 3464 29205 3473
rect 29163 3424 29164 3464
rect 29204 3424 29205 3464
rect 29163 3415 29205 3424
rect 31083 3464 31125 3473
rect 31083 3424 31084 3464
rect 31124 3424 31125 3464
rect 31083 3415 31125 3424
rect 31755 3464 31797 3473
rect 31755 3424 31756 3464
rect 31796 3424 31797 3464
rect 31755 3415 31797 3424
rect 37419 3464 37461 3473
rect 37419 3424 37420 3464
rect 37460 3424 37461 3464
rect 37419 3415 37461 3424
rect 37803 3464 37845 3473
rect 37803 3424 37804 3464
rect 37844 3424 37845 3464
rect 37803 3415 37845 3424
rect 13275 3296 13317 3305
rect 13275 3256 13276 3296
rect 13316 3256 13317 3296
rect 13275 3247 13317 3256
rect 17979 3296 18021 3305
rect 17979 3256 17980 3296
rect 18020 3256 18021 3296
rect 17979 3247 18021 3256
rect 18363 3296 18405 3305
rect 18363 3256 18364 3296
rect 18404 3256 18405 3296
rect 18363 3247 18405 3256
rect 22107 3212 22149 3221
rect 22107 3172 22108 3212
rect 22148 3172 22149 3212
rect 22107 3163 22149 3172
rect 22491 3212 22533 3221
rect 22491 3172 22492 3212
rect 22532 3172 22533 3212
rect 22491 3163 22533 3172
rect 37659 3212 37701 3221
rect 37659 3172 37660 3212
rect 37700 3172 37701 3212
rect 37659 3163 37701 3172
rect 1152 3044 38112 3068
rect 1152 3004 4928 3044
rect 4968 3004 5010 3044
rect 5050 3004 5092 3044
rect 5132 3004 5174 3044
rect 5214 3004 5256 3044
rect 5296 3004 20048 3044
rect 20088 3004 20130 3044
rect 20170 3004 20212 3044
rect 20252 3004 20294 3044
rect 20334 3004 20376 3044
rect 20416 3004 35168 3044
rect 35208 3004 35250 3044
rect 35290 3004 35332 3044
rect 35372 3004 35414 3044
rect 35454 3004 35496 3044
rect 35536 3004 38112 3044
rect 1152 2980 38112 3004
rect 38043 2792 38085 2801
rect 38043 2752 38044 2792
rect 38084 2752 38085 2792
rect 38043 2743 38085 2752
rect 18027 2624 18069 2633
rect 18027 2584 18028 2624
rect 18068 2584 18069 2624
rect 18027 2575 18069 2584
rect 18411 2624 18453 2633
rect 18411 2584 18412 2624
rect 18452 2584 18453 2624
rect 18411 2575 18453 2584
rect 18795 2624 18837 2633
rect 18795 2584 18796 2624
rect 18836 2584 18837 2624
rect 18795 2575 18837 2584
rect 19179 2624 19221 2633
rect 19179 2584 19180 2624
rect 19220 2584 19221 2624
rect 19179 2575 19221 2584
rect 19563 2624 19605 2633
rect 19563 2584 19564 2624
rect 19604 2584 19605 2624
rect 19563 2575 19605 2584
rect 19947 2624 19989 2633
rect 19947 2584 19948 2624
rect 19988 2584 19989 2624
rect 19947 2575 19989 2584
rect 21675 2624 21717 2633
rect 21675 2584 21676 2624
rect 21716 2584 21717 2624
rect 21675 2575 21717 2584
rect 22059 2624 22101 2633
rect 22059 2584 22060 2624
rect 22100 2584 22101 2624
rect 22059 2575 22101 2584
rect 22443 2624 22485 2633
rect 22443 2584 22444 2624
rect 22484 2584 22485 2624
rect 22443 2575 22485 2584
rect 22762 2624 22820 2625
rect 22762 2584 22771 2624
rect 22811 2584 22820 2624
rect 22762 2583 22820 2584
rect 23211 2624 23253 2633
rect 23211 2584 23212 2624
rect 23252 2584 23253 2624
rect 23211 2575 23253 2584
rect 23595 2624 23637 2633
rect 23595 2584 23596 2624
rect 23636 2584 23637 2624
rect 23595 2575 23637 2584
rect 23979 2624 24021 2633
rect 23979 2584 23980 2624
rect 24020 2584 24021 2624
rect 23979 2575 24021 2584
rect 24363 2624 24405 2633
rect 24363 2584 24364 2624
rect 24404 2584 24405 2624
rect 24363 2575 24405 2584
rect 24747 2624 24789 2633
rect 24747 2584 24748 2624
rect 24788 2584 24789 2624
rect 24747 2575 24789 2584
rect 25131 2624 25173 2633
rect 25131 2584 25132 2624
rect 25172 2584 25173 2624
rect 25131 2575 25173 2584
rect 25515 2624 25557 2633
rect 25515 2584 25516 2624
rect 25556 2584 25557 2624
rect 25515 2575 25557 2584
rect 25899 2624 25941 2633
rect 25899 2584 25900 2624
rect 25940 2584 25941 2624
rect 25899 2575 25941 2584
rect 26283 2624 26325 2633
rect 26283 2584 26284 2624
rect 26324 2584 26325 2624
rect 26283 2575 26325 2584
rect 26667 2624 26709 2633
rect 26667 2584 26668 2624
rect 26708 2584 26709 2624
rect 26667 2575 26709 2584
rect 27051 2624 27093 2633
rect 27051 2584 27052 2624
rect 27092 2584 27093 2624
rect 27051 2575 27093 2584
rect 27435 2624 27477 2633
rect 27435 2584 27436 2624
rect 27476 2584 27477 2624
rect 27435 2575 27477 2584
rect 37035 2624 37077 2633
rect 37035 2584 37036 2624
rect 37076 2584 37077 2624
rect 37035 2575 37077 2584
rect 37419 2624 37461 2633
rect 37419 2584 37420 2624
rect 37460 2584 37461 2624
rect 37419 2575 37461 2584
rect 37803 2624 37845 2633
rect 37803 2584 37804 2624
rect 37844 2584 37845 2624
rect 37803 2575 37845 2584
rect 37659 2540 37701 2549
rect 37659 2500 37660 2540
rect 37700 2500 37701 2540
rect 37659 2491 37701 2500
rect 17787 2456 17829 2465
rect 17787 2416 17788 2456
rect 17828 2416 17829 2456
rect 17787 2407 17829 2416
rect 18171 2456 18213 2465
rect 18171 2416 18172 2456
rect 18212 2416 18213 2456
rect 18171 2407 18213 2416
rect 18555 2456 18597 2465
rect 18555 2416 18556 2456
rect 18596 2416 18597 2456
rect 18555 2407 18597 2416
rect 18939 2456 18981 2465
rect 18939 2416 18940 2456
rect 18980 2416 18981 2456
rect 18939 2407 18981 2416
rect 19323 2456 19365 2465
rect 19323 2416 19324 2456
rect 19364 2416 19365 2456
rect 19323 2407 19365 2416
rect 19707 2456 19749 2465
rect 19707 2416 19708 2456
rect 19748 2416 19749 2456
rect 19707 2407 19749 2416
rect 21435 2456 21477 2465
rect 21435 2416 21436 2456
rect 21476 2416 21477 2456
rect 21435 2407 21477 2416
rect 21819 2456 21861 2465
rect 21819 2416 21820 2456
rect 21860 2416 21861 2456
rect 21819 2407 21861 2416
rect 22203 2456 22245 2465
rect 22203 2416 22204 2456
rect 22244 2416 22245 2456
rect 22203 2407 22245 2416
rect 22587 2456 22629 2465
rect 22587 2416 22588 2456
rect 22628 2416 22629 2456
rect 22587 2407 22629 2416
rect 22971 2456 23013 2465
rect 22971 2416 22972 2456
rect 23012 2416 23013 2456
rect 22971 2407 23013 2416
rect 23355 2456 23397 2465
rect 23355 2416 23356 2456
rect 23396 2416 23397 2456
rect 23355 2407 23397 2416
rect 23739 2456 23781 2465
rect 23739 2416 23740 2456
rect 23780 2416 23781 2456
rect 23739 2407 23781 2416
rect 24123 2456 24165 2465
rect 24123 2416 24124 2456
rect 24164 2416 24165 2456
rect 24123 2407 24165 2416
rect 24507 2456 24549 2465
rect 24507 2416 24508 2456
rect 24548 2416 24549 2456
rect 24507 2407 24549 2416
rect 24891 2456 24933 2465
rect 24891 2416 24892 2456
rect 24932 2416 24933 2456
rect 24891 2407 24933 2416
rect 25275 2456 25317 2465
rect 25275 2416 25276 2456
rect 25316 2416 25317 2456
rect 25275 2407 25317 2416
rect 25659 2456 25701 2465
rect 25659 2416 25660 2456
rect 25700 2416 25701 2456
rect 25659 2407 25701 2416
rect 26043 2456 26085 2465
rect 26043 2416 26044 2456
rect 26084 2416 26085 2456
rect 26043 2407 26085 2416
rect 26427 2456 26469 2465
rect 26427 2416 26428 2456
rect 26468 2416 26469 2456
rect 26427 2407 26469 2416
rect 26811 2456 26853 2465
rect 26811 2416 26812 2456
rect 26852 2416 26853 2456
rect 26811 2407 26853 2416
rect 27195 2456 27237 2465
rect 27195 2416 27196 2456
rect 27236 2416 27237 2456
rect 27195 2407 27237 2416
rect 37275 2456 37317 2465
rect 37275 2416 37276 2456
rect 37316 2416 37317 2456
rect 37275 2407 37317 2416
rect 1152 2288 38112 2312
rect 1152 2248 3688 2288
rect 3728 2248 3770 2288
rect 3810 2248 3852 2288
rect 3892 2248 3934 2288
rect 3974 2248 4016 2288
rect 4056 2248 18808 2288
rect 18848 2248 18890 2288
rect 18930 2248 18972 2288
rect 19012 2248 19054 2288
rect 19094 2248 19136 2288
rect 19176 2248 33928 2288
rect 33968 2248 34010 2288
rect 34050 2248 34092 2288
rect 34132 2248 34174 2288
rect 34214 2248 34256 2288
rect 34296 2248 38112 2288
rect 1152 2224 38112 2248
rect 38043 2120 38085 2129
rect 38043 2080 38044 2120
rect 38084 2080 38085 2120
rect 38043 2071 38085 2080
rect 22011 2036 22053 2045
rect 22011 1996 22012 2036
rect 22052 1996 22053 2036
rect 22011 1987 22053 1996
rect 23163 2036 23205 2045
rect 23163 1996 23164 2036
rect 23204 1996 23205 2036
rect 23163 1987 23205 1996
rect 27003 2036 27045 2045
rect 27003 1996 27004 2036
rect 27044 1996 27045 2036
rect 27003 1987 27045 1996
rect 17067 1952 17109 1961
rect 17067 1912 17068 1952
rect 17108 1912 17109 1952
rect 17067 1903 17109 1912
rect 17451 1952 17493 1961
rect 17451 1912 17452 1952
rect 17492 1912 17493 1952
rect 17451 1903 17493 1912
rect 17866 1952 17924 1953
rect 17866 1912 17875 1952
rect 17915 1912 17924 1952
rect 17866 1911 17924 1912
rect 18219 1952 18261 1961
rect 18219 1912 18220 1952
rect 18260 1912 18261 1952
rect 18219 1903 18261 1912
rect 18603 1952 18645 1961
rect 18603 1912 18604 1952
rect 18644 1912 18645 1952
rect 18603 1903 18645 1912
rect 18987 1952 19029 1961
rect 18987 1912 18988 1952
rect 19028 1912 19029 1952
rect 18987 1903 19029 1912
rect 19371 1952 19413 1961
rect 19371 1912 19372 1952
rect 19412 1912 19413 1952
rect 19371 1903 19413 1912
rect 19755 1952 19797 1961
rect 19755 1912 19756 1952
rect 19796 1912 19797 1952
rect 19755 1903 19797 1912
rect 20139 1952 20181 1961
rect 20139 1912 20140 1952
rect 20180 1912 20181 1952
rect 20139 1903 20181 1912
rect 20715 1952 20757 1961
rect 20715 1912 20716 1952
rect 20756 1912 20757 1952
rect 20715 1903 20757 1912
rect 21099 1952 21141 1961
rect 21099 1912 21100 1952
rect 21140 1912 21141 1952
rect 21099 1903 21141 1912
rect 21483 1952 21525 1961
rect 21483 1912 21484 1952
rect 21524 1912 21525 1952
rect 21483 1903 21525 1912
rect 21867 1952 21909 1961
rect 21867 1912 21868 1952
rect 21908 1912 21909 1952
rect 21867 1903 21909 1912
rect 22251 1952 22293 1961
rect 22251 1912 22252 1952
rect 22292 1912 22293 1952
rect 22251 1903 22293 1912
rect 22635 1952 22677 1961
rect 22635 1912 22636 1952
rect 22676 1912 22677 1952
rect 22635 1903 22677 1912
rect 23019 1952 23061 1961
rect 23019 1912 23020 1952
rect 23060 1912 23061 1952
rect 23019 1903 23061 1912
rect 23403 1952 23445 1961
rect 23403 1912 23404 1952
rect 23444 1912 23445 1952
rect 23403 1903 23445 1912
rect 23787 1952 23829 1961
rect 23787 1912 23788 1952
rect 23828 1912 23829 1952
rect 23787 1903 23829 1912
rect 24171 1952 24213 1961
rect 24171 1912 24172 1952
rect 24212 1912 24213 1952
rect 24171 1903 24213 1912
rect 24555 1952 24597 1961
rect 24555 1912 24556 1952
rect 24596 1912 24597 1952
rect 24555 1903 24597 1912
rect 24939 1952 24981 1961
rect 24939 1912 24940 1952
rect 24980 1912 24981 1952
rect 24939 1903 24981 1912
rect 25323 1952 25365 1961
rect 25323 1912 25324 1952
rect 25364 1912 25365 1952
rect 25323 1903 25365 1912
rect 25707 1952 25749 1961
rect 25707 1912 25708 1952
rect 25748 1912 25749 1952
rect 25707 1903 25749 1912
rect 26091 1952 26133 1961
rect 26091 1912 26092 1952
rect 26132 1912 26133 1952
rect 26091 1903 26133 1912
rect 26475 1952 26517 1961
rect 26475 1912 26476 1952
rect 26516 1912 26517 1952
rect 26475 1903 26517 1912
rect 26859 1952 26901 1961
rect 26859 1912 26860 1952
rect 26900 1912 26901 1952
rect 26859 1903 26901 1912
rect 27243 1952 27285 1961
rect 27243 1912 27244 1952
rect 27284 1912 27285 1952
rect 27243 1903 27285 1912
rect 27627 1952 27669 1961
rect 27627 1912 27628 1952
rect 27668 1912 27669 1952
rect 27627 1903 27669 1912
rect 28011 1952 28053 1961
rect 28011 1912 28012 1952
rect 28052 1912 28053 1952
rect 28011 1903 28053 1912
rect 28395 1952 28437 1961
rect 28395 1912 28396 1952
rect 28436 1912 28437 1952
rect 28395 1903 28437 1912
rect 36651 1952 36693 1961
rect 36651 1912 36652 1952
rect 36692 1912 36693 1952
rect 36651 1903 36693 1912
rect 37035 1952 37077 1961
rect 37035 1912 37036 1952
rect 37076 1912 37077 1952
rect 37035 1903 37077 1912
rect 37419 1952 37461 1961
rect 37419 1912 37420 1952
rect 37460 1912 37461 1952
rect 37419 1903 37461 1912
rect 37803 1952 37845 1961
rect 37803 1912 37804 1952
rect 37844 1912 37845 1952
rect 37803 1903 37845 1912
rect 19611 1784 19653 1793
rect 19611 1744 19612 1784
rect 19652 1744 19653 1784
rect 19611 1735 19653 1744
rect 20379 1784 20421 1793
rect 20379 1744 20380 1784
rect 20420 1744 20421 1784
rect 20379 1735 20421 1744
rect 21243 1784 21285 1793
rect 21243 1744 21244 1784
rect 21284 1744 21285 1784
rect 21243 1735 21285 1744
rect 22395 1784 22437 1793
rect 22395 1744 22396 1784
rect 22436 1744 22437 1784
rect 22395 1735 22437 1744
rect 23547 1784 23589 1793
rect 23547 1744 23548 1784
rect 23588 1744 23589 1784
rect 23547 1735 23589 1744
rect 24699 1784 24741 1793
rect 24699 1744 24700 1784
rect 24740 1744 24741 1784
rect 24699 1735 24741 1744
rect 25851 1784 25893 1793
rect 25851 1744 25852 1784
rect 25892 1744 25893 1784
rect 25851 1735 25893 1744
rect 27387 1784 27429 1793
rect 27387 1744 27388 1784
rect 27428 1744 27429 1784
rect 27387 1735 27429 1744
rect 36891 1784 36933 1793
rect 36891 1744 36892 1784
rect 36932 1744 36933 1784
rect 36891 1735 36933 1744
rect 37659 1784 37701 1793
rect 37659 1744 37660 1784
rect 37700 1744 37701 1784
rect 37659 1735 37701 1744
rect 17307 1700 17349 1709
rect 17307 1660 17308 1700
rect 17348 1660 17349 1700
rect 17307 1651 17349 1660
rect 17691 1700 17733 1709
rect 17691 1660 17692 1700
rect 17732 1660 17733 1700
rect 17691 1651 17733 1660
rect 18075 1700 18117 1709
rect 18075 1660 18076 1700
rect 18116 1660 18117 1700
rect 18075 1651 18117 1660
rect 18459 1700 18501 1709
rect 18459 1660 18460 1700
rect 18500 1660 18501 1700
rect 18459 1651 18501 1660
rect 18843 1700 18885 1709
rect 18843 1660 18844 1700
rect 18884 1660 18885 1700
rect 18843 1651 18885 1660
rect 19227 1700 19269 1709
rect 19227 1660 19228 1700
rect 19268 1660 19269 1700
rect 19227 1651 19269 1660
rect 19995 1700 20037 1709
rect 19995 1660 19996 1700
rect 20036 1660 20037 1700
rect 19995 1651 20037 1660
rect 20475 1700 20517 1709
rect 20475 1660 20476 1700
rect 20516 1660 20517 1700
rect 20475 1651 20517 1660
rect 20859 1700 20901 1709
rect 20859 1660 20860 1700
rect 20900 1660 20901 1700
rect 20859 1651 20901 1660
rect 21627 1700 21669 1709
rect 21627 1660 21628 1700
rect 21668 1660 21669 1700
rect 21627 1651 21669 1660
rect 22779 1700 22821 1709
rect 22779 1660 22780 1700
rect 22820 1660 22821 1700
rect 22779 1651 22821 1660
rect 23931 1700 23973 1709
rect 23931 1660 23932 1700
rect 23972 1660 23973 1700
rect 23931 1651 23973 1660
rect 24315 1700 24357 1709
rect 24315 1660 24316 1700
rect 24356 1660 24357 1700
rect 24315 1651 24357 1660
rect 25083 1700 25125 1709
rect 25083 1660 25084 1700
rect 25124 1660 25125 1700
rect 25083 1651 25125 1660
rect 25467 1700 25509 1709
rect 25467 1660 25468 1700
rect 25508 1660 25509 1700
rect 25467 1651 25509 1660
rect 26235 1700 26277 1709
rect 26235 1660 26236 1700
rect 26276 1660 26277 1700
rect 26235 1651 26277 1660
rect 26619 1700 26661 1709
rect 26619 1660 26620 1700
rect 26660 1660 26661 1700
rect 26619 1651 26661 1660
rect 27771 1700 27813 1709
rect 27771 1660 27772 1700
rect 27812 1660 27813 1700
rect 27771 1651 27813 1660
rect 28155 1700 28197 1709
rect 28155 1660 28156 1700
rect 28196 1660 28197 1700
rect 28155 1651 28197 1660
rect 37275 1700 37317 1709
rect 37275 1660 37276 1700
rect 37316 1660 37317 1700
rect 37275 1651 37317 1660
rect 1152 1532 38112 1556
rect 1152 1492 4928 1532
rect 4968 1492 5010 1532
rect 5050 1492 5092 1532
rect 5132 1492 5174 1532
rect 5214 1492 5256 1532
rect 5296 1492 20048 1532
rect 20088 1492 20130 1532
rect 20170 1492 20212 1532
rect 20252 1492 20294 1532
rect 20334 1492 20376 1532
rect 20416 1492 35168 1532
rect 35208 1492 35250 1532
rect 35290 1492 35332 1532
rect 35372 1492 35414 1532
rect 35454 1492 35496 1532
rect 35536 1492 38112 1532
rect 1152 1468 38112 1492
<< via1 >>
rect 4928 10564 4968 10604
rect 5010 10564 5050 10604
rect 5092 10564 5132 10604
rect 5174 10564 5214 10604
rect 5256 10564 5296 10604
rect 20048 10564 20088 10604
rect 20130 10564 20170 10604
rect 20212 10564 20252 10604
rect 20294 10564 20334 10604
rect 20376 10564 20416 10604
rect 35168 10564 35208 10604
rect 35250 10564 35290 10604
rect 35332 10564 35372 10604
rect 35414 10564 35454 10604
rect 35496 10564 35536 10604
rect 2236 10396 2276 10436
rect 3964 10396 4004 10436
rect 5692 10396 5732 10436
rect 7420 10396 7460 10436
rect 9148 10396 9188 10436
rect 10876 10396 10916 10436
rect 12604 10396 12644 10436
rect 14332 10396 14372 10436
rect 16060 10396 16100 10436
rect 17788 10396 17828 10436
rect 19516 10396 19556 10436
rect 21244 10396 21284 10436
rect 22972 10396 23012 10436
rect 24700 10396 24740 10436
rect 26428 10396 26468 10436
rect 28156 10396 28196 10436
rect 29884 10396 29924 10436
rect 31612 10396 31652 10436
rect 33340 10396 33380 10436
rect 35068 10396 35108 10436
rect 36316 10396 36356 10436
rect 36796 10396 36836 10436
rect 2476 10144 2516 10184
rect 4204 10144 4244 10184
rect 5932 10144 5972 10184
rect 7660 10144 7700 10184
rect 9388 10144 9428 10184
rect 11116 10144 11156 10184
rect 12844 10144 12884 10184
rect 14572 10144 14612 10184
rect 16300 10144 16340 10184
rect 18028 10144 18068 10184
rect 19804 10144 19844 10184
rect 21484 10144 21524 10184
rect 23212 10144 23252 10184
rect 24940 10144 24980 10184
rect 26668 10144 26708 10184
rect 28396 10144 28436 10184
rect 30124 10144 30164 10184
rect 31852 10144 31892 10184
rect 33580 10144 33620 10184
rect 35308 10144 35348 10184
rect 36076 10144 36116 10184
rect 36460 10144 36500 10184
rect 37036 10144 37076 10184
rect 37420 10144 37460 10184
rect 37804 10144 37844 10184
rect 36700 10060 36740 10100
rect 37660 9976 37700 10016
rect 38044 9976 38084 10016
rect 3688 9808 3728 9848
rect 3770 9808 3810 9848
rect 3852 9808 3892 9848
rect 3934 9808 3974 9848
rect 4016 9808 4056 9848
rect 18808 9808 18848 9848
rect 18890 9808 18930 9848
rect 18972 9808 19012 9848
rect 19054 9808 19094 9848
rect 19136 9808 19176 9848
rect 33928 9808 33968 9848
rect 34010 9808 34050 9848
rect 34092 9808 34132 9848
rect 34174 9808 34214 9848
rect 34256 9808 34296 9848
rect 36892 9640 36932 9680
rect 37276 9640 37316 9680
rect 36652 9472 36692 9512
rect 37036 9472 37076 9512
rect 37420 9472 37460 9512
rect 37804 9472 37844 9512
rect 37660 9220 37700 9260
rect 38044 9220 38084 9260
rect 4928 9052 4968 9092
rect 5010 9052 5050 9092
rect 5092 9052 5132 9092
rect 5174 9052 5214 9092
rect 5256 9052 5296 9092
rect 20048 9052 20088 9092
rect 20130 9052 20170 9092
rect 20212 9052 20252 9092
rect 20294 9052 20334 9092
rect 20376 9052 20416 9092
rect 35168 9052 35208 9092
rect 35250 9052 35290 9092
rect 35332 9052 35372 9092
rect 35414 9052 35454 9092
rect 35496 9052 35536 9092
rect 5500 8884 5540 8924
rect 6652 8884 6692 8924
rect 8188 8884 8228 8924
rect 16924 8884 16964 8924
rect 17884 8884 17924 8924
rect 18748 8884 18788 8924
rect 20092 8884 20132 8924
rect 28252 8884 28292 8924
rect 13084 8800 13124 8840
rect 14908 8800 14948 8840
rect 15292 8800 15332 8840
rect 16828 8800 16868 8840
rect 18364 8800 18404 8840
rect 22684 8800 22724 8840
rect 5260 8632 5300 8672
rect 6412 8632 6452 8672
rect 7948 8632 7988 8672
rect 12844 8632 12884 8672
rect 13228 8632 13268 8672
rect 13900 8632 13940 8672
rect 14140 8632 14180 8672
rect 14668 8632 14708 8672
rect 15052 8632 15092 8672
rect 15532 8632 15572 8672
rect 15772 8632 15812 8672
rect 16588 8632 16628 8672
rect 17164 8632 17204 8672
rect 17644 8632 17684 8672
rect 18124 8632 18164 8672
rect 18508 8632 18548 8672
rect 18988 8632 19028 8672
rect 19228 8632 19268 8672
rect 19507 8632 19547 8672
rect 19891 8632 19931 8672
rect 20524 8632 20564 8672
rect 20908 8632 20948 8672
rect 21148 8632 21188 8672
rect 21772 8632 21812 8672
rect 22924 8632 22964 8672
rect 24316 8632 24356 8672
rect 24556 8632 24596 8672
rect 25132 8632 25172 8672
rect 25372 8632 25412 8672
rect 25804 8632 25844 8672
rect 27436 8632 27476 8672
rect 27820 8632 27860 8672
rect 28051 8632 28091 8672
rect 29068 8632 29108 8672
rect 29308 8632 29348 8672
rect 37420 8632 37460 8672
rect 37804 8632 37844 8672
rect 38044 8632 38084 8672
rect 20764 8548 20804 8588
rect 25564 8548 25604 8588
rect 27196 8548 27236 8588
rect 27580 8548 27620 8588
rect 37660 8548 37700 8588
rect 13468 8464 13508 8504
rect 19708 8464 19748 8504
rect 22012 8464 22052 8504
rect 3688 8296 3728 8336
rect 3770 8296 3810 8336
rect 3852 8296 3892 8336
rect 3934 8296 3974 8336
rect 4016 8296 4056 8336
rect 18808 8296 18848 8336
rect 18890 8296 18930 8336
rect 18972 8296 19012 8336
rect 19054 8296 19094 8336
rect 19136 8296 19176 8336
rect 33928 8296 33968 8336
rect 34010 8296 34050 8336
rect 34092 8296 34132 8336
rect 34174 8296 34214 8336
rect 34256 8296 34296 8336
rect 29212 8128 29252 8168
rect 10684 8044 10724 8084
rect 11356 8044 11396 8084
rect 10444 7960 10484 8000
rect 11116 7960 11156 8000
rect 11500 7960 11540 8000
rect 29452 7960 29492 8000
rect 37420 7960 37460 8000
rect 37804 7960 37844 8000
rect 37660 7792 37700 7832
rect 11740 7708 11780 7748
rect 38044 7708 38084 7748
rect 4928 7540 4968 7580
rect 5010 7540 5050 7580
rect 5092 7540 5132 7580
rect 5174 7540 5214 7580
rect 5256 7540 5296 7580
rect 20048 7540 20088 7580
rect 20130 7540 20170 7580
rect 20212 7540 20252 7580
rect 20294 7540 20334 7580
rect 20376 7540 20416 7580
rect 35168 7540 35208 7580
rect 35250 7540 35290 7580
rect 35332 7540 35372 7580
rect 35414 7540 35454 7580
rect 35496 7540 35536 7580
rect 6028 7120 6068 7160
rect 37420 7120 37460 7160
rect 37804 7120 37844 7160
rect 38044 7120 38084 7160
rect 5788 7036 5828 7076
rect 37660 6952 37700 6992
rect 3688 6784 3728 6824
rect 3770 6784 3810 6824
rect 3852 6784 3892 6824
rect 3934 6784 3974 6824
rect 4016 6784 4056 6824
rect 18808 6784 18848 6824
rect 18890 6784 18930 6824
rect 18972 6784 19012 6824
rect 19054 6784 19094 6824
rect 19136 6784 19176 6824
rect 33928 6784 33968 6824
rect 34010 6784 34050 6824
rect 34092 6784 34132 6824
rect 34174 6784 34214 6824
rect 34256 6784 34296 6824
rect 2620 6616 2660 6656
rect 27484 6616 27524 6656
rect 2860 6448 2900 6488
rect 27724 6448 27764 6488
rect 31468 6448 31508 6488
rect 37420 6448 37460 6488
rect 37804 6448 37844 6488
rect 38044 6448 38084 6488
rect 31708 6196 31748 6236
rect 37660 6196 37700 6236
rect 4928 6028 4968 6068
rect 5010 6028 5050 6068
rect 5092 6028 5132 6068
rect 5174 6028 5214 6068
rect 5256 6028 5296 6068
rect 20048 6028 20088 6068
rect 20130 6028 20170 6068
rect 20212 6028 20252 6068
rect 20294 6028 20334 6068
rect 20376 6028 20416 6068
rect 35168 6028 35208 6068
rect 35250 6028 35290 6068
rect 35332 6028 35372 6068
rect 35414 6028 35454 6068
rect 35496 6028 35536 6068
rect 38044 5776 38084 5816
rect 2668 5608 2708 5648
rect 2908 5608 2948 5648
rect 37420 5608 37460 5648
rect 37804 5608 37844 5648
rect 37660 5524 37700 5564
rect 3688 5272 3728 5312
rect 3770 5272 3810 5312
rect 3852 5272 3892 5312
rect 3934 5272 3974 5312
rect 4016 5272 4056 5312
rect 18808 5272 18848 5312
rect 18890 5272 18930 5312
rect 18972 5272 19012 5312
rect 19054 5272 19094 5312
rect 19136 5272 19176 5312
rect 33928 5272 33968 5312
rect 34010 5272 34050 5312
rect 34092 5272 34132 5312
rect 34174 5272 34214 5312
rect 34256 5272 34296 5312
rect 7900 5104 7940 5144
rect 8380 5104 8420 5144
rect 10396 5104 10436 5144
rect 27868 5104 27908 5144
rect 33628 5104 33668 5144
rect 38044 5104 38084 5144
rect 16252 5020 16292 5060
rect 7276 4936 7316 4976
rect 7660 4936 7700 4976
rect 8140 4936 8180 4976
rect 8524 4936 8564 4976
rect 8908 4936 8948 4976
rect 9292 4936 9332 4976
rect 9772 4936 9812 4976
rect 10156 4936 10196 4976
rect 13132 4936 13172 4976
rect 13372 4936 13412 4976
rect 16012 4936 16052 4976
rect 17068 4936 17108 4976
rect 17644 4936 17684 4976
rect 18028 4936 18068 4976
rect 21964 4936 22004 4976
rect 22348 4936 22388 4976
rect 25708 4936 25748 4976
rect 26188 4936 26228 4976
rect 28108 4936 28148 4976
rect 31276 4936 31316 4976
rect 33388 4936 33428 4976
rect 37420 4936 37460 4976
rect 37804 4936 37844 4976
rect 10012 4768 10052 4808
rect 37660 4768 37700 4808
rect 7516 4684 7556 4724
rect 8764 4684 8804 4724
rect 9148 4684 9188 4724
rect 9532 4684 9572 4724
rect 17308 4684 17348 4724
rect 17884 4684 17924 4724
rect 18268 4684 18308 4724
rect 22204 4684 22244 4724
rect 22588 4684 22628 4724
rect 25948 4684 25988 4724
rect 26428 4684 26468 4724
rect 31516 4684 31556 4724
rect 4928 4516 4968 4556
rect 5010 4516 5050 4556
rect 5092 4516 5132 4556
rect 5174 4516 5214 4556
rect 5256 4516 5296 4556
rect 20048 4516 20088 4556
rect 20130 4516 20170 4556
rect 20212 4516 20252 4556
rect 20294 4516 20334 4556
rect 20376 4516 20416 4556
rect 35168 4516 35208 4556
rect 35250 4516 35290 4556
rect 35332 4516 35372 4556
rect 35414 4516 35454 4556
rect 35496 4516 35536 4556
rect 26140 4348 26180 4388
rect 13276 4264 13316 4304
rect 18652 4264 18692 4304
rect 22492 4264 22532 4304
rect 23644 4264 23684 4304
rect 32476 4264 32516 4304
rect 32860 4264 32900 4304
rect 38044 4264 38084 4304
rect 8236 4096 8276 4136
rect 8620 4096 8660 4136
rect 9964 4096 10004 4136
rect 10348 4096 10388 4136
rect 11884 4096 11924 4136
rect 12268 4096 12308 4136
rect 12652 4096 12692 4136
rect 13036 4096 13076 4136
rect 13420 4096 13460 4136
rect 13804 4096 13844 4136
rect 14380 4096 14420 4136
rect 16108 4096 16148 4136
rect 16492 4096 16532 4136
rect 16876 4096 16916 4136
rect 17260 4096 17300 4136
rect 17644 4096 17684 4136
rect 18028 4096 18068 4136
rect 18412 4096 18452 4136
rect 18796 4096 18836 4136
rect 19180 4096 19220 4136
rect 19420 4096 19460 4136
rect 19756 4096 19796 4136
rect 21100 4096 21140 4136
rect 21484 4096 21524 4136
rect 21868 4096 21908 4136
rect 22252 4096 22292 4136
rect 22636 4096 22676 4136
rect 23020 4096 23060 4136
rect 23404 4096 23444 4136
rect 23788 4096 23828 4136
rect 24172 4096 24212 4136
rect 25900 4096 25940 4136
rect 27244 4096 27284 4136
rect 28588 4096 28628 4136
rect 29644 4096 29684 4136
rect 31564 4096 31604 4136
rect 32236 4096 32276 4136
rect 32620 4096 32660 4136
rect 33004 4096 33044 4136
rect 37036 4096 37076 4136
rect 37420 4096 37460 4136
rect 37804 4096 37844 4136
rect 12124 4012 12164 4052
rect 14044 4012 14084 4052
rect 14620 4012 14660 4052
rect 24412 4012 24452 4052
rect 31804 4012 31844 4052
rect 33244 4012 33284 4052
rect 37660 4012 37700 4052
rect 8476 3928 8516 3968
rect 8860 3928 8900 3968
rect 10204 3928 10244 3968
rect 10588 3928 10628 3968
rect 12508 3928 12548 3968
rect 12892 3928 12932 3968
rect 13660 3928 13700 3968
rect 16348 3928 16388 3968
rect 16732 3928 16772 3968
rect 17116 3928 17156 3968
rect 17500 3928 17540 3968
rect 17884 3928 17924 3968
rect 18268 3928 18308 3968
rect 19036 3928 19076 3968
rect 19996 3928 20036 3968
rect 21340 3928 21380 3968
rect 21724 3928 21764 3968
rect 22108 3928 22148 3968
rect 22876 3928 22916 3968
rect 23260 3928 23300 3968
rect 24028 3928 24068 3968
rect 27484 3928 27524 3968
rect 28348 3928 28388 3968
rect 29404 3928 29444 3968
rect 37276 3928 37316 3968
rect 3688 3760 3728 3800
rect 3770 3760 3810 3800
rect 3852 3760 3892 3800
rect 3934 3760 3974 3800
rect 4016 3760 4056 3800
rect 18808 3760 18848 3800
rect 18890 3760 18930 3800
rect 18972 3760 19012 3800
rect 19054 3760 19094 3800
rect 19136 3760 19176 3800
rect 33928 3760 33968 3800
rect 34010 3760 34050 3800
rect 34092 3760 34132 3800
rect 34174 3760 34214 3800
rect 34256 3760 34296 3800
rect 27580 3592 27620 3632
rect 28924 3592 28964 3632
rect 30844 3592 30884 3632
rect 31996 3592 32036 3632
rect 38044 3592 38084 3632
rect 13036 3424 13076 3464
rect 13420 3424 13460 3464
rect 13660 3424 13700 3464
rect 17740 3424 17780 3464
rect 18124 3424 18164 3464
rect 21868 3424 21908 3464
rect 22252 3424 22292 3464
rect 27820 3424 27860 3464
rect 29164 3424 29204 3464
rect 31084 3424 31124 3464
rect 31756 3424 31796 3464
rect 37420 3424 37460 3464
rect 37804 3424 37844 3464
rect 13276 3256 13316 3296
rect 17980 3256 18020 3296
rect 18364 3256 18404 3296
rect 22108 3172 22148 3212
rect 22492 3172 22532 3212
rect 37660 3172 37700 3212
rect 4928 3004 4968 3044
rect 5010 3004 5050 3044
rect 5092 3004 5132 3044
rect 5174 3004 5214 3044
rect 5256 3004 5296 3044
rect 20048 3004 20088 3044
rect 20130 3004 20170 3044
rect 20212 3004 20252 3044
rect 20294 3004 20334 3044
rect 20376 3004 20416 3044
rect 35168 3004 35208 3044
rect 35250 3004 35290 3044
rect 35332 3004 35372 3044
rect 35414 3004 35454 3044
rect 35496 3004 35536 3044
rect 38044 2752 38084 2792
rect 18028 2584 18068 2624
rect 18412 2584 18452 2624
rect 18796 2584 18836 2624
rect 19180 2584 19220 2624
rect 19564 2584 19604 2624
rect 19948 2584 19988 2624
rect 21676 2584 21716 2624
rect 22060 2584 22100 2624
rect 22444 2584 22484 2624
rect 22771 2584 22811 2624
rect 23212 2584 23252 2624
rect 23596 2584 23636 2624
rect 23980 2584 24020 2624
rect 24364 2584 24404 2624
rect 24748 2584 24788 2624
rect 25132 2584 25172 2624
rect 25516 2584 25556 2624
rect 25900 2584 25940 2624
rect 26284 2584 26324 2624
rect 26668 2584 26708 2624
rect 27052 2584 27092 2624
rect 27436 2584 27476 2624
rect 37036 2584 37076 2624
rect 37420 2584 37460 2624
rect 37804 2584 37844 2624
rect 37660 2500 37700 2540
rect 17788 2416 17828 2456
rect 18172 2416 18212 2456
rect 18556 2416 18596 2456
rect 18940 2416 18980 2456
rect 19324 2416 19364 2456
rect 19708 2416 19748 2456
rect 21436 2416 21476 2456
rect 21820 2416 21860 2456
rect 22204 2416 22244 2456
rect 22588 2416 22628 2456
rect 22972 2416 23012 2456
rect 23356 2416 23396 2456
rect 23740 2416 23780 2456
rect 24124 2416 24164 2456
rect 24508 2416 24548 2456
rect 24892 2416 24932 2456
rect 25276 2416 25316 2456
rect 25660 2416 25700 2456
rect 26044 2416 26084 2456
rect 26428 2416 26468 2456
rect 26812 2416 26852 2456
rect 27196 2416 27236 2456
rect 37276 2416 37316 2456
rect 3688 2248 3728 2288
rect 3770 2248 3810 2288
rect 3852 2248 3892 2288
rect 3934 2248 3974 2288
rect 4016 2248 4056 2288
rect 18808 2248 18848 2288
rect 18890 2248 18930 2288
rect 18972 2248 19012 2288
rect 19054 2248 19094 2288
rect 19136 2248 19176 2288
rect 33928 2248 33968 2288
rect 34010 2248 34050 2288
rect 34092 2248 34132 2288
rect 34174 2248 34214 2288
rect 34256 2248 34296 2288
rect 38044 2080 38084 2120
rect 22012 1996 22052 2036
rect 23164 1996 23204 2036
rect 27004 1996 27044 2036
rect 17068 1912 17108 1952
rect 17452 1912 17492 1952
rect 17875 1912 17915 1952
rect 18220 1912 18260 1952
rect 18604 1912 18644 1952
rect 18988 1912 19028 1952
rect 19372 1912 19412 1952
rect 19756 1912 19796 1952
rect 20140 1912 20180 1952
rect 20716 1912 20756 1952
rect 21100 1912 21140 1952
rect 21484 1912 21524 1952
rect 21868 1912 21908 1952
rect 22252 1912 22292 1952
rect 22636 1912 22676 1952
rect 23020 1912 23060 1952
rect 23404 1912 23444 1952
rect 23788 1912 23828 1952
rect 24172 1912 24212 1952
rect 24556 1912 24596 1952
rect 24940 1912 24980 1952
rect 25324 1912 25364 1952
rect 25708 1912 25748 1952
rect 26092 1912 26132 1952
rect 26476 1912 26516 1952
rect 26860 1912 26900 1952
rect 27244 1912 27284 1952
rect 27628 1912 27668 1952
rect 28012 1912 28052 1952
rect 28396 1912 28436 1952
rect 36652 1912 36692 1952
rect 37036 1912 37076 1952
rect 37420 1912 37460 1952
rect 37804 1912 37844 1952
rect 19612 1744 19652 1784
rect 20380 1744 20420 1784
rect 21244 1744 21284 1784
rect 22396 1744 22436 1784
rect 23548 1744 23588 1784
rect 24700 1744 24740 1784
rect 25852 1744 25892 1784
rect 27388 1744 27428 1784
rect 36892 1744 36932 1784
rect 37660 1744 37700 1784
rect 17308 1660 17348 1700
rect 17692 1660 17732 1700
rect 18076 1660 18116 1700
rect 18460 1660 18500 1700
rect 18844 1660 18884 1700
rect 19228 1660 19268 1700
rect 19996 1660 20036 1700
rect 20476 1660 20516 1700
rect 20860 1660 20900 1700
rect 21628 1660 21668 1700
rect 22780 1660 22820 1700
rect 23932 1660 23972 1700
rect 24316 1660 24356 1700
rect 25084 1660 25124 1700
rect 25468 1660 25508 1700
rect 26236 1660 26276 1700
rect 26620 1660 26660 1700
rect 27772 1660 27812 1700
rect 28156 1660 28196 1700
rect 37276 1660 37316 1700
rect 4928 1492 4968 1532
rect 5010 1492 5050 1532
rect 5092 1492 5132 1532
rect 5174 1492 5214 1532
rect 5256 1492 5296 1532
rect 20048 1492 20088 1532
rect 20130 1492 20170 1532
rect 20212 1492 20252 1532
rect 20294 1492 20334 1532
rect 20376 1492 20416 1532
rect 35168 1492 35208 1532
rect 35250 1492 35290 1532
rect 35332 1492 35372 1532
rect 35414 1492 35454 1532
rect 35496 1492 35536 1532
<< metal2 >>
rect 0 11192 90 11212
rect 39174 11192 39264 11212
rect 0 11152 20524 11192
rect 20564 11152 20573 11192
rect 36931 11152 36940 11192
rect 36980 11152 39264 11192
rect 0 11132 90 11152
rect 39174 11132 39264 11152
rect 0 10856 90 10876
rect 39174 10856 39264 10876
rect 0 10816 8620 10856
rect 8660 10816 8669 10856
rect 11395 10816 11404 10856
rect 11444 10816 28012 10856
rect 28052 10816 28061 10856
rect 36355 10816 36364 10856
rect 36404 10816 39264 10856
rect 0 10796 90 10816
rect 39174 10796 39264 10816
rect 14563 10732 14572 10772
rect 14612 10732 27148 10772
rect 27188 10732 27197 10772
rect 31651 10732 31660 10772
rect 31700 10732 37804 10772
rect 37844 10732 37853 10772
rect 15331 10648 15340 10688
rect 15380 10648 36500 10688
rect 4919 10564 4928 10604
rect 4968 10564 5010 10604
rect 5050 10564 5092 10604
rect 5132 10564 5174 10604
rect 5214 10564 5256 10604
rect 5296 10564 5305 10604
rect 20039 10564 20048 10604
rect 20088 10564 20130 10604
rect 20170 10564 20212 10604
rect 20252 10564 20294 10604
rect 20334 10564 20376 10604
rect 20416 10564 20425 10604
rect 20524 10564 28684 10604
rect 28724 10564 28733 10604
rect 35159 10564 35168 10604
rect 35208 10564 35250 10604
rect 35290 10564 35332 10604
rect 35372 10564 35414 10604
rect 35454 10564 35496 10604
rect 35536 10564 35545 10604
rect 0 10520 90 10540
rect 0 10480 652 10520
rect 692 10480 701 10520
rect 2860 10480 14668 10520
rect 14708 10480 14717 10520
rect 0 10460 90 10480
rect 2179 10396 2188 10436
rect 2228 10396 2236 10436
rect 2276 10396 2359 10436
rect 2860 10352 2900 10480
rect 3907 10396 3916 10436
rect 3956 10396 3964 10436
rect 4004 10396 4087 10436
rect 5635 10396 5644 10436
rect 5684 10396 5692 10436
rect 5732 10396 5815 10436
rect 7363 10396 7372 10436
rect 7412 10396 7420 10436
rect 7460 10396 7543 10436
rect 9091 10396 9100 10436
rect 9140 10396 9148 10436
rect 9188 10396 9271 10436
rect 10819 10396 10828 10436
rect 10868 10396 10876 10436
rect 10916 10396 10999 10436
rect 12547 10396 12556 10436
rect 12596 10396 12604 10436
rect 12644 10396 12727 10436
rect 14275 10396 14284 10436
rect 14324 10396 14332 10436
rect 14372 10396 14455 10436
rect 16003 10396 16012 10436
rect 16052 10396 16060 10436
rect 16100 10396 16183 10436
rect 17731 10396 17740 10436
rect 17780 10396 17788 10436
rect 17828 10396 17911 10436
rect 19459 10396 19468 10436
rect 19508 10396 19516 10436
rect 19556 10396 19639 10436
rect 20524 10352 20564 10564
rect 36460 10520 36500 10648
rect 39174 10520 39264 10540
rect 21955 10480 21964 10520
rect 22004 10480 33140 10520
rect 36460 10480 37172 10520
rect 37315 10480 37324 10520
rect 37364 10480 39264 10520
rect 21187 10396 21196 10436
rect 21236 10396 21244 10436
rect 21284 10396 21367 10436
rect 22841 10396 22924 10436
rect 22964 10396 22972 10436
rect 23012 10396 23021 10436
rect 24643 10396 24652 10436
rect 24692 10396 24700 10436
rect 24740 10396 24823 10436
rect 26371 10396 26380 10436
rect 26420 10396 26428 10436
rect 26468 10396 26551 10436
rect 28099 10396 28108 10436
rect 28148 10396 28156 10436
rect 28196 10396 28279 10436
rect 29827 10396 29836 10436
rect 29876 10396 29884 10436
rect 29924 10396 30007 10436
rect 31555 10396 31564 10436
rect 31604 10396 31612 10436
rect 31652 10396 31735 10436
rect 33100 10352 33140 10480
rect 33283 10396 33292 10436
rect 33332 10396 33340 10436
rect 33380 10396 33463 10436
rect 35011 10396 35020 10436
rect 35060 10396 35068 10436
rect 35108 10396 35191 10436
rect 36233 10396 36316 10436
rect 36356 10396 36364 10436
rect 36404 10396 36413 10436
rect 36739 10396 36748 10436
rect 36788 10396 36796 10436
rect 36836 10396 36919 10436
rect 172 10312 2900 10352
rect 12940 10312 20564 10352
rect 21388 10312 22636 10352
rect 22676 10312 22685 10352
rect 33100 10312 36500 10352
rect 0 10184 90 10204
rect 172 10184 212 10312
rect 12940 10184 12980 10312
rect 16300 10228 20140 10268
rect 20180 10228 20189 10268
rect 16300 10184 16340 10228
rect 21388 10184 21428 10312
rect 21484 10228 25900 10268
rect 25940 10228 25949 10268
rect 28003 10228 28012 10268
rect 28052 10228 36116 10268
rect 21484 10184 21524 10228
rect 36076 10184 36116 10228
rect 36460 10184 36500 10312
rect 37132 10184 37172 10480
rect 39174 10460 39264 10480
rect 39174 10184 39264 10204
rect 0 10144 212 10184
rect 2467 10144 2476 10184
rect 2516 10144 2668 10184
rect 2708 10144 2717 10184
rect 4073 10144 4204 10184
rect 4244 10144 4253 10184
rect 5801 10144 5932 10184
rect 5972 10144 5981 10184
rect 7529 10144 7660 10184
rect 7700 10144 7709 10184
rect 9379 10144 9388 10184
rect 9428 10144 9437 10184
rect 11107 10144 11116 10184
rect 11156 10144 11165 10184
rect 12835 10144 12844 10184
rect 12884 10144 12980 10184
rect 14441 10144 14572 10184
rect 14612 10144 14621 10184
rect 16291 10144 16300 10184
rect 16340 10144 16349 10184
rect 18019 10144 18028 10184
rect 18068 10144 19660 10184
rect 19700 10144 19709 10184
rect 19795 10144 19804 10184
rect 19844 10144 19892 10184
rect 19939 10144 19948 10184
rect 19988 10144 21428 10184
rect 21475 10144 21484 10184
rect 21524 10144 21533 10184
rect 23081 10144 23212 10184
rect 23252 10144 23261 10184
rect 24931 10144 24940 10184
rect 24980 10144 26380 10184
rect 26420 10144 26429 10184
rect 26537 10144 26668 10184
rect 26708 10144 26717 10184
rect 28265 10144 28396 10184
rect 28436 10144 28445 10184
rect 29993 10144 30124 10184
rect 30164 10144 30173 10184
rect 31721 10144 31852 10184
rect 31892 10144 31901 10184
rect 32899 10144 32908 10184
rect 32948 10144 33580 10184
rect 33620 10144 33629 10184
rect 35299 10144 35308 10184
rect 35348 10144 35357 10184
rect 36067 10144 36076 10184
rect 36116 10144 36125 10184
rect 36451 10144 36460 10184
rect 36500 10144 36509 10184
rect 36556 10144 37036 10184
rect 37076 10144 37085 10184
rect 37132 10144 37420 10184
rect 37460 10144 37469 10184
rect 37673 10144 37804 10184
rect 37844 10144 37853 10184
rect 38284 10144 39264 10184
rect 0 10124 90 10144
rect 9388 10100 9428 10144
rect 5731 10060 5740 10100
rect 5780 10060 9428 10100
rect 11116 10100 11156 10144
rect 19852 10100 19892 10144
rect 35308 10100 35348 10144
rect 36556 10100 36596 10144
rect 38284 10100 38324 10144
rect 39174 10124 39264 10144
rect 11116 10060 15820 10100
rect 15860 10060 15869 10100
rect 19852 10060 24268 10100
rect 24308 10060 24317 10100
rect 27916 10060 28100 10100
rect 32515 10060 32524 10100
rect 32564 10060 35348 10100
rect 35587 10060 35596 10100
rect 35636 10060 36596 10100
rect 36691 10060 36700 10100
rect 36740 10060 38324 10100
rect 14947 9976 14956 10016
rect 14996 9976 21964 10016
rect 22004 9976 22013 10016
rect 27916 9932 27956 10060
rect 28060 10016 28100 10060
rect 28060 9976 37228 10016
rect 37268 9976 37277 10016
rect 37420 9976 37556 10016
rect 37651 9976 37660 10016
rect 37700 9976 37709 10016
rect 38035 9976 38044 10016
rect 38084 9976 38764 10016
rect 38804 9976 38813 10016
rect 37420 9932 37460 9976
rect 16867 9892 16876 9932
rect 16916 9892 27956 9932
rect 28195 9892 28204 9932
rect 28244 9892 37460 9932
rect 0 9848 90 9868
rect 0 9808 2900 9848
rect 3679 9808 3688 9848
rect 3728 9808 3770 9848
rect 3810 9808 3852 9848
rect 3892 9808 3934 9848
rect 3974 9808 4016 9848
rect 4056 9808 4065 9848
rect 18799 9808 18808 9848
rect 18848 9808 18890 9848
rect 18930 9808 18972 9848
rect 19012 9808 19054 9848
rect 19094 9808 19136 9848
rect 19176 9808 19185 9848
rect 24067 9808 24076 9848
rect 24116 9808 29260 9848
rect 29300 9808 29309 9848
rect 33919 9808 33928 9848
rect 33968 9808 34010 9848
rect 34050 9808 34092 9848
rect 34132 9808 34174 9848
rect 34214 9808 34256 9848
rect 34296 9808 34305 9848
rect 0 9788 90 9808
rect 2860 9764 2900 9808
rect 37516 9764 37556 9976
rect 37660 9848 37700 9976
rect 39174 9848 39264 9868
rect 37660 9808 39264 9848
rect 39174 9788 39264 9808
rect 2860 9724 15052 9764
rect 15092 9724 15101 9764
rect 17155 9724 17164 9764
rect 17204 9724 24364 9764
rect 24404 9724 24413 9764
rect 24547 9724 24556 9764
rect 24596 9724 29452 9764
rect 29492 9724 29501 9764
rect 37516 9724 37804 9764
rect 37844 9724 37853 9764
rect 10723 9640 10732 9680
rect 10772 9640 36652 9680
rect 36692 9640 36701 9680
rect 36809 9640 36892 9680
rect 36932 9640 36940 9680
rect 36980 9640 36989 9680
rect 37193 9640 37276 9680
rect 37316 9640 37324 9680
rect 37364 9640 37373 9680
rect 8227 9556 8236 9596
rect 8276 9556 37076 9596
rect 0 9512 90 9532
rect 37036 9512 37076 9556
rect 39174 9512 39264 9532
rect 0 9472 18988 9512
rect 19028 9472 19037 9512
rect 19084 9472 21004 9512
rect 21044 9472 21053 9512
rect 21187 9472 21196 9512
rect 21236 9472 24308 9512
rect 24355 9472 24364 9512
rect 24404 9472 27724 9512
rect 27764 9472 27773 9512
rect 27820 9472 36652 9512
rect 36692 9472 36701 9512
rect 37027 9472 37036 9512
rect 37076 9472 37085 9512
rect 37219 9472 37228 9512
rect 37268 9472 37420 9512
rect 37460 9472 37469 9512
rect 37603 9472 37612 9512
rect 37652 9472 37804 9512
rect 37844 9472 37853 9512
rect 38755 9472 38764 9512
rect 38804 9472 39264 9512
rect 0 9452 90 9472
rect 19084 9428 19124 9472
rect 835 9388 844 9428
rect 884 9388 19124 9428
rect 20131 9388 20140 9428
rect 20180 9388 23020 9428
rect 23060 9388 23069 9428
rect 24268 9344 24308 9472
rect 27820 9428 27860 9472
rect 39174 9452 39264 9472
rect 24451 9388 24460 9428
rect 24500 9388 27860 9428
rect 30211 9388 30220 9428
rect 30260 9388 31660 9428
rect 31700 9388 31709 9428
rect 36652 9388 37708 9428
rect 37748 9388 37757 9428
rect 36652 9344 36692 9388
rect 931 9304 940 9344
rect 980 9304 19468 9344
rect 19508 9304 19517 9344
rect 19564 9304 22924 9344
rect 22964 9304 22973 9344
rect 24268 9304 36692 9344
rect 36748 9304 37900 9344
rect 37940 9304 37949 9344
rect 19564 9260 19604 9304
rect 36748 9260 36788 9304
rect 19171 9220 19180 9260
rect 19220 9220 19604 9260
rect 30787 9220 30796 9260
rect 30836 9220 36788 9260
rect 37651 9220 37660 9260
rect 37700 9220 37709 9260
rect 38035 9220 38044 9260
rect 38084 9220 38668 9260
rect 38708 9220 38717 9260
rect 0 9176 90 9196
rect 37660 9176 37700 9220
rect 39174 9176 39264 9196
rect 0 9136 16588 9176
rect 16628 9136 16637 9176
rect 18787 9136 18796 9176
rect 18836 9136 22924 9176
rect 22964 9136 22973 9176
rect 37660 9136 39264 9176
rect 0 9116 90 9136
rect 39174 9116 39264 9136
rect 4919 9052 4928 9092
rect 4968 9052 5010 9092
rect 5050 9052 5092 9092
rect 5132 9052 5174 9092
rect 5214 9052 5256 9092
rect 5296 9052 5305 9092
rect 15715 9052 15724 9092
rect 15764 9052 19660 9092
rect 19700 9052 19709 9092
rect 19756 9052 19988 9092
rect 20039 9052 20048 9092
rect 20088 9052 20130 9092
rect 20170 9052 20212 9092
rect 20252 9052 20294 9092
rect 20334 9052 20376 9092
rect 20416 9052 20425 9092
rect 25795 9052 25804 9092
rect 25844 9052 28972 9092
rect 29012 9052 29021 9092
rect 35159 9052 35168 9092
rect 35208 9052 35250 9092
rect 35290 9052 35332 9092
rect 35372 9052 35414 9092
rect 35454 9052 35496 9092
rect 35536 9052 35545 9092
rect 19756 9008 19796 9052
rect 172 8968 17300 9008
rect 0 8840 90 8860
rect 172 8840 212 8968
rect 5491 8884 5500 8924
rect 5540 8884 5740 8924
rect 5780 8884 5789 8924
rect 6643 8884 6652 8924
rect 6692 8884 7660 8924
rect 7700 8884 7709 8924
rect 8105 8884 8188 8924
rect 8228 8884 8236 8924
rect 8276 8884 8285 8924
rect 15811 8884 15820 8924
rect 15860 8884 16924 8924
rect 16964 8884 16973 8924
rect 0 8800 212 8840
rect 1411 8800 1420 8840
rect 1460 8800 12940 8840
rect 12980 8800 12989 8840
rect 13075 8800 13084 8840
rect 13124 8800 14380 8840
rect 14420 8800 14429 8840
rect 14825 8800 14908 8840
rect 14948 8800 14956 8840
rect 14996 8800 15005 8840
rect 15283 8800 15292 8840
rect 15332 8800 15340 8840
rect 15380 8800 15463 8840
rect 16745 8800 16828 8840
rect 16868 8800 16876 8840
rect 16916 8800 16925 8840
rect 0 8780 90 8800
rect 643 8716 652 8756
rect 692 8716 7988 8756
rect 10051 8716 10060 8756
rect 10100 8716 13940 8756
rect 7948 8672 7988 8716
rect 13900 8672 13940 8716
rect 17260 8672 17300 8968
rect 18604 8968 19796 9008
rect 19948 9008 19988 9052
rect 19948 8968 25228 9008
rect 25268 8968 25277 9008
rect 27811 8968 27820 9008
rect 27860 8968 29644 9008
rect 29684 8968 29693 9008
rect 30211 8968 30220 9008
rect 30260 8968 37844 9008
rect 18604 8924 18644 8968
rect 17875 8884 17884 8924
rect 17924 8884 18644 8924
rect 18739 8884 18748 8924
rect 18788 8884 18796 8924
rect 18836 8884 18919 8924
rect 20083 8884 20092 8924
rect 20132 8884 20620 8924
rect 20660 8884 20669 8924
rect 28243 8884 28252 8924
rect 28292 8884 30796 8924
rect 30836 8884 30845 8924
rect 33100 8884 37612 8924
rect 37652 8884 37661 8924
rect 33100 8840 33140 8884
rect 18355 8800 18364 8840
rect 18404 8800 21580 8840
rect 21620 8800 21629 8840
rect 22627 8800 22636 8840
rect 22676 8800 22684 8840
rect 22724 8800 22807 8840
rect 25219 8800 25228 8840
rect 25268 8800 33140 8840
rect 37420 8800 37516 8840
rect 37556 8800 37565 8840
rect 37420 8756 37460 8800
rect 17731 8716 17740 8756
rect 17780 8716 20948 8756
rect 20995 8716 21004 8756
rect 21044 8716 21812 8756
rect 23107 8716 23116 8756
rect 23156 8716 25268 8756
rect 20908 8672 20948 8716
rect 21772 8672 21812 8716
rect 5251 8632 5260 8672
rect 5300 8632 5740 8672
rect 5780 8632 5789 8672
rect 6281 8632 6412 8672
rect 6452 8632 6461 8672
rect 7939 8632 7948 8672
rect 7988 8632 7997 8672
rect 8131 8632 8140 8672
rect 8180 8632 12844 8672
rect 12884 8632 12893 8672
rect 13097 8632 13228 8672
rect 13268 8632 13277 8672
rect 13891 8632 13900 8672
rect 13940 8632 13949 8672
rect 14131 8632 14140 8672
rect 14180 8632 14284 8672
rect 14324 8632 14333 8672
rect 14537 8632 14668 8672
rect 14708 8632 14717 8672
rect 14921 8632 15052 8672
rect 15092 8632 15101 8672
rect 15401 8632 15532 8672
rect 15572 8632 15581 8672
rect 15763 8632 15772 8672
rect 15812 8632 15820 8672
rect 15860 8632 15943 8672
rect 16579 8632 16588 8672
rect 16628 8632 16759 8672
rect 17033 8632 17164 8672
rect 17204 8632 17213 8672
rect 17260 8632 17644 8672
rect 17684 8632 17693 8672
rect 17740 8632 18124 8672
rect 18164 8632 18173 8672
rect 18220 8632 18508 8672
rect 18548 8632 18557 8672
rect 18857 8632 18988 8672
rect 19028 8632 19037 8672
rect 19171 8632 19180 8672
rect 19220 8632 19228 8672
rect 19268 8632 19351 8672
rect 19498 8632 19507 8672
rect 19547 8632 19564 8672
rect 19604 8632 19687 8672
rect 19756 8632 19891 8672
rect 19931 8632 19940 8672
rect 20393 8632 20524 8672
rect 20564 8632 20573 8672
rect 20899 8632 20908 8672
rect 20948 8632 20957 8672
rect 21065 8632 21148 8672
rect 21188 8632 21196 8672
rect 21236 8632 21245 8672
rect 21763 8632 21772 8672
rect 21812 8632 21821 8672
rect 22915 8632 22924 8672
rect 22964 8632 24076 8672
rect 24116 8632 24125 8672
rect 24259 8632 24268 8672
rect 24308 8632 24316 8672
rect 24356 8632 24439 8672
rect 24547 8632 24556 8672
rect 24596 8632 24727 8672
rect 25001 8632 25132 8672
rect 25172 8632 25181 8672
rect 17740 8588 17780 8632
rect 17251 8548 17260 8588
rect 17300 8548 17780 8588
rect 0 8504 90 8524
rect 18220 8504 18260 8632
rect 19756 8588 19796 8632
rect 25228 8588 25268 8716
rect 25708 8716 37460 8756
rect 25708 8672 25748 8716
rect 37804 8672 37844 8968
rect 39174 8840 39264 8860
rect 38659 8800 38668 8840
rect 38708 8800 39264 8840
rect 39174 8780 39264 8800
rect 25363 8632 25372 8672
rect 25412 8632 25748 8672
rect 25795 8632 25804 8672
rect 25844 8632 25975 8672
rect 26083 8632 26092 8672
rect 26132 8632 27380 8672
rect 27427 8632 27436 8672
rect 27476 8632 27764 8672
rect 27811 8632 27820 8672
rect 27860 8632 27991 8672
rect 28042 8632 28051 8672
rect 28091 8632 28108 8672
rect 28148 8632 28231 8672
rect 28300 8632 28780 8672
rect 28820 8632 28829 8672
rect 28937 8632 29068 8672
rect 29108 8632 29117 8672
rect 29299 8632 29308 8672
rect 29348 8632 33484 8672
rect 33524 8632 33533 8672
rect 36643 8632 36652 8672
rect 36692 8632 37420 8672
rect 37460 8632 37469 8672
rect 37795 8632 37804 8672
rect 37844 8632 37853 8672
rect 38035 8632 38044 8672
rect 38084 8632 39148 8672
rect 39188 8632 39197 8672
rect 27340 8588 27380 8632
rect 27724 8588 27764 8632
rect 28300 8588 28340 8632
rect 19651 8548 19660 8588
rect 19700 8548 19796 8588
rect 20755 8548 20764 8588
rect 20804 8548 24460 8588
rect 24500 8548 24509 8588
rect 25228 8548 25564 8588
rect 25604 8548 25613 8588
rect 27065 8548 27148 8588
rect 27188 8548 27196 8588
rect 27236 8548 27245 8588
rect 27340 8548 27580 8588
rect 27620 8548 27629 8588
rect 27724 8548 28340 8588
rect 37651 8548 37660 8588
rect 37700 8548 38516 8588
rect 38476 8504 38516 8548
rect 39174 8504 39264 8524
rect 0 8464 2420 8504
rect 13459 8464 13468 8504
rect 13508 8464 13996 8504
rect 14036 8464 14045 8504
rect 17155 8464 17164 8504
rect 17204 8464 18260 8504
rect 19699 8464 19708 8504
rect 19748 8464 19756 8504
rect 19796 8464 19879 8504
rect 22003 8464 22012 8504
rect 22052 8464 28204 8504
rect 28244 8464 28253 8504
rect 38476 8464 39264 8504
rect 0 8444 90 8464
rect 2380 8420 2420 8464
rect 39174 8444 39264 8464
rect 2380 8380 2860 8420
rect 2900 8380 2909 8420
rect 12940 8380 15724 8420
rect 15764 8380 15773 8420
rect 3679 8296 3688 8336
rect 3728 8296 3770 8336
rect 3810 8296 3852 8336
rect 3892 8296 3934 8336
rect 3974 8296 4016 8336
rect 4056 8296 4065 8336
rect 0 8168 90 8188
rect 12940 8168 12980 8380
rect 18799 8296 18808 8336
rect 18848 8296 18890 8336
rect 18930 8296 18972 8336
rect 19012 8296 19054 8336
rect 19094 8296 19136 8336
rect 19176 8296 19185 8336
rect 33919 8296 33928 8336
rect 33968 8296 34010 8336
rect 34050 8296 34092 8336
rect 34132 8296 34174 8336
rect 34214 8296 34256 8336
rect 34296 8296 34305 8336
rect 39174 8168 39264 8188
rect 0 8128 12980 8168
rect 28675 8128 28684 8168
rect 28724 8128 29212 8168
rect 29252 8128 29261 8168
rect 39139 8128 39148 8168
rect 39188 8128 39264 8168
rect 0 8108 90 8128
rect 39174 8108 39264 8128
rect 10601 8044 10684 8084
rect 10724 8044 10732 8084
rect 10772 8044 10781 8084
rect 11273 8044 11356 8084
rect 11396 8044 11404 8084
rect 11444 8044 11453 8084
rect 13987 8044 13996 8084
rect 14036 8044 37844 8084
rect 37804 8000 37844 8044
rect 2947 7960 2956 8000
rect 2996 7960 10444 8000
rect 10484 7960 10493 8000
rect 11107 7960 11116 8000
rect 11156 7960 11165 8000
rect 11491 7960 11500 8000
rect 11540 7960 11549 8000
rect 28675 7960 28684 8000
rect 28724 7960 29452 8000
rect 29492 7960 29501 8000
rect 37411 7960 37420 8000
rect 37460 7960 37469 8000
rect 37795 7960 37804 8000
rect 37844 7960 37853 8000
rect 11116 7916 11156 7960
rect 8611 7876 8620 7916
rect 8660 7876 11156 7916
rect 0 7832 90 7852
rect 11500 7832 11540 7960
rect 0 7792 11540 7832
rect 0 7772 90 7792
rect 11731 7708 11740 7748
rect 11780 7708 12980 7748
rect 12940 7664 12980 7708
rect 37420 7664 37460 7960
rect 39174 7832 39264 7852
rect 37651 7792 37660 7832
rect 37700 7792 39264 7832
rect 39174 7772 39264 7792
rect 38035 7708 38044 7748
rect 38084 7708 38093 7748
rect 12940 7624 37460 7664
rect 4919 7540 4928 7580
rect 4968 7540 5010 7580
rect 5050 7540 5092 7580
rect 5132 7540 5174 7580
rect 5214 7540 5256 7580
rect 5296 7540 5305 7580
rect 20039 7540 20048 7580
rect 20088 7540 20130 7580
rect 20170 7540 20212 7580
rect 20252 7540 20294 7580
rect 20334 7540 20376 7580
rect 20416 7540 20425 7580
rect 35159 7540 35168 7580
rect 35208 7540 35250 7580
rect 35290 7540 35332 7580
rect 35372 7540 35414 7580
rect 35454 7540 35496 7580
rect 35536 7540 35545 7580
rect 0 7496 90 7516
rect 38044 7496 38084 7708
rect 39174 7496 39264 7516
rect 0 7456 13228 7496
rect 13268 7456 13277 7496
rect 38044 7456 39264 7496
rect 0 7436 90 7456
rect 39174 7436 39264 7456
rect 0 7160 90 7180
rect 39174 7160 39264 7180
rect 0 7120 2900 7160
rect 5897 7120 6028 7160
rect 6068 7120 6077 7160
rect 14371 7120 14380 7160
rect 14420 7120 37420 7160
rect 37460 7120 37469 7160
rect 37795 7120 37804 7160
rect 37844 7120 37853 7160
rect 38035 7120 38044 7160
rect 38084 7120 39264 7160
rect 0 7100 90 7120
rect 2860 6992 2900 7120
rect 37804 7076 37844 7120
rect 39174 7100 39264 7120
rect 5779 7036 5788 7076
rect 5828 7036 5932 7076
rect 5972 7036 5981 7076
rect 12940 7036 17260 7076
rect 17300 7036 17309 7076
rect 21571 7036 21580 7076
rect 21620 7036 37844 7076
rect 12940 6992 12980 7036
rect 2860 6952 12980 6992
rect 37651 6952 37660 6992
rect 37700 6952 38612 6992
rect 2860 6868 8140 6908
rect 8180 6868 8189 6908
rect 0 6824 90 6844
rect 2860 6824 2900 6868
rect 38572 6824 38612 6952
rect 39174 6824 39264 6844
rect 0 6784 2900 6824
rect 3679 6784 3688 6824
rect 3728 6784 3770 6824
rect 3810 6784 3852 6824
rect 3892 6784 3934 6824
rect 3974 6784 4016 6824
rect 4056 6784 4065 6824
rect 18799 6784 18808 6824
rect 18848 6784 18890 6824
rect 18930 6784 18972 6824
rect 19012 6784 19054 6824
rect 19094 6784 19136 6824
rect 19176 6784 19185 6824
rect 33919 6784 33928 6824
rect 33968 6784 34010 6824
rect 34050 6784 34092 6824
rect 34132 6784 34174 6824
rect 34214 6784 34256 6824
rect 34296 6784 34305 6824
rect 38572 6784 39264 6824
rect 0 6764 90 6784
rect 39174 6764 39264 6784
rect 2537 6616 2620 6656
rect 2660 6616 2668 6656
rect 2708 6616 2717 6656
rect 23203 6616 23212 6656
rect 23252 6616 27484 6656
rect 27524 6616 27533 6656
rect 22915 6532 22924 6572
rect 22964 6532 37460 6572
rect 0 6488 90 6508
rect 37420 6488 37460 6532
rect 39174 6488 39264 6508
rect 0 6448 844 6488
rect 884 6448 893 6488
rect 2851 6448 2860 6488
rect 2900 6448 2956 6488
rect 2996 6448 3031 6488
rect 27715 6448 27724 6488
rect 27764 6448 29836 6488
rect 29876 6448 29885 6488
rect 31459 6448 31468 6488
rect 31508 6448 31517 6488
rect 37411 6448 37420 6488
rect 37460 6448 37469 6488
rect 37673 6448 37804 6488
rect 37844 6448 37853 6488
rect 38035 6448 38044 6488
rect 38084 6448 39264 6488
rect 0 6428 90 6448
rect 31468 6404 31508 6448
rect 39174 6428 39264 6448
rect 547 6364 556 6404
rect 596 6364 31508 6404
rect 31699 6196 31708 6236
rect 31748 6196 35980 6236
rect 36020 6196 36029 6236
rect 37651 6196 37660 6236
rect 37700 6196 38900 6236
rect 0 6152 90 6172
rect 38860 6152 38900 6196
rect 39174 6152 39264 6172
rect 0 6112 17164 6152
rect 17204 6112 17213 6152
rect 38860 6112 39264 6152
rect 0 6092 90 6112
rect 39174 6092 39264 6112
rect 4919 6028 4928 6068
rect 4968 6028 5010 6068
rect 5050 6028 5092 6068
rect 5132 6028 5174 6068
rect 5214 6028 5256 6068
rect 5296 6028 5305 6068
rect 20039 6028 20048 6068
rect 20088 6028 20130 6068
rect 20170 6028 20212 6068
rect 20252 6028 20294 6068
rect 20334 6028 20376 6068
rect 20416 6028 20425 6068
rect 35159 6028 35168 6068
rect 35208 6028 35250 6068
rect 35290 6028 35332 6068
rect 35372 6028 35414 6068
rect 35454 6028 35496 6068
rect 35536 6028 35545 6068
rect 0 5816 90 5836
rect 39174 5816 39264 5836
rect 0 5776 15532 5816
rect 15572 5776 15581 5816
rect 38035 5776 38044 5816
rect 38084 5776 39264 5816
rect 0 5756 90 5776
rect 39174 5756 39264 5776
rect 7660 5692 8812 5732
rect 8852 5692 8861 5732
rect 15811 5692 15820 5732
rect 15860 5692 37844 5732
rect 2537 5608 2668 5648
rect 2708 5608 2717 5648
rect 2899 5608 2908 5648
rect 2948 5608 4204 5648
rect 4244 5608 4253 5648
rect 7660 5564 7700 5692
rect 37804 5648 37844 5692
rect 1219 5524 1228 5564
rect 1268 5524 7700 5564
rect 7756 5608 10060 5648
rect 10100 5608 10109 5648
rect 14275 5608 14284 5648
rect 14324 5608 37420 5648
rect 37460 5608 37469 5648
rect 37795 5608 37804 5648
rect 37844 5608 37853 5648
rect 0 5480 90 5500
rect 7756 5480 7796 5608
rect 9187 5524 9196 5564
rect 9236 5524 16972 5564
rect 17012 5524 17021 5564
rect 37651 5524 37660 5564
rect 37700 5524 38708 5564
rect 38668 5480 38708 5524
rect 39174 5480 39264 5500
rect 0 5440 7796 5480
rect 8236 5440 9868 5480
rect 9908 5440 9917 5480
rect 12940 5440 16340 5480
rect 16867 5440 16876 5480
rect 16916 5440 22348 5480
rect 22388 5440 22397 5480
rect 38668 5440 39264 5480
rect 0 5420 90 5440
rect 3679 5272 3688 5312
rect 3728 5272 3770 5312
rect 3810 5272 3852 5312
rect 3892 5272 3934 5312
rect 3974 5272 4016 5312
rect 4056 5272 4065 5312
rect 0 5144 90 5164
rect 8236 5144 8276 5440
rect 12940 5396 12980 5440
rect 8620 5356 12980 5396
rect 8620 5144 8660 5356
rect 16300 5312 16340 5440
rect 39174 5420 39264 5440
rect 20131 5356 20140 5396
rect 20180 5356 24172 5396
rect 24212 5356 24221 5396
rect 8899 5272 8908 5312
rect 8948 5272 9964 5312
rect 10004 5272 10013 5312
rect 10147 5272 10156 5312
rect 10196 5272 16204 5312
rect 16244 5272 16253 5312
rect 16300 5272 17836 5312
rect 17876 5272 17885 5312
rect 18799 5272 18808 5312
rect 18848 5272 18890 5312
rect 18930 5272 18972 5312
rect 19012 5272 19054 5312
rect 19094 5272 19136 5312
rect 19176 5272 19185 5312
rect 19276 5272 31316 5312
rect 33919 5272 33928 5312
rect 33968 5272 34010 5312
rect 34050 5272 34092 5312
rect 34132 5272 34174 5312
rect 34214 5272 34256 5312
rect 34296 5272 34305 5312
rect 8803 5188 8812 5228
rect 8852 5188 13268 5228
rect 16483 5188 16492 5228
rect 16532 5188 18220 5228
rect 18260 5188 18269 5228
rect 13228 5144 13268 5188
rect 19276 5144 19316 5272
rect 0 5104 1420 5144
rect 1460 5104 1469 5144
rect 7891 5104 7900 5144
rect 7940 5104 8276 5144
rect 8371 5104 8380 5144
rect 8420 5104 8660 5144
rect 8707 5104 8716 5144
rect 8756 5104 9812 5144
rect 10387 5104 10396 5144
rect 10436 5104 13036 5144
rect 13076 5104 13085 5144
rect 13228 5104 19316 5144
rect 22156 5188 24940 5228
rect 24980 5188 24989 5228
rect 0 5084 90 5104
rect 8524 5020 9484 5060
rect 9524 5020 9533 5060
rect 8524 4976 8564 5020
rect 9772 4976 9812 5104
rect 22156 5060 22196 5188
rect 26371 5104 26380 5144
rect 26420 5104 27868 5144
rect 27908 5104 27917 5144
rect 11875 5020 11884 5060
rect 11924 5020 16052 5060
rect 16243 5020 16252 5060
rect 16292 5020 22196 5060
rect 23020 5020 26228 5060
rect 16012 4976 16052 5020
rect 7267 4936 7276 4976
rect 7316 4936 7325 4976
rect 7651 4936 7660 4976
rect 7700 4936 7948 4976
rect 7988 4936 7997 4976
rect 8131 4936 8140 4976
rect 8180 4936 8468 4976
rect 8515 4936 8524 4976
rect 8564 4936 8573 4976
rect 8899 4936 8908 4976
rect 8948 4936 8957 4976
rect 9091 4936 9100 4976
rect 9140 4936 9292 4976
rect 9332 4936 9341 4976
rect 9763 4936 9772 4976
rect 9812 4936 9821 4976
rect 9955 4936 9964 4976
rect 10004 4936 10156 4976
rect 10196 4936 10205 4976
rect 11395 4936 11404 4976
rect 11444 4936 13132 4976
rect 13172 4936 13181 4976
rect 13289 4936 13372 4976
rect 13412 4936 13420 4976
rect 13460 4936 13469 4976
rect 16003 4936 16012 4976
rect 16052 4936 16061 4976
rect 16937 4936 17068 4976
rect 17108 4936 17117 4976
rect 17251 4936 17260 4976
rect 17300 4936 17644 4976
rect 17684 4936 17693 4976
rect 17897 4936 17932 4976
rect 17972 4936 18028 4976
rect 18068 4936 18077 4976
rect 18211 4936 18220 4976
rect 18260 4936 21964 4976
rect 22004 4936 22013 4976
rect 22217 4936 22348 4976
rect 22388 4936 22397 4976
rect 7276 4892 7316 4936
rect 8428 4892 8468 4936
rect 8908 4892 8948 4936
rect 23020 4892 23060 5020
rect 26188 4976 26228 5020
rect 31276 4976 31316 5272
rect 39174 5144 39264 5164
rect 33619 5104 33628 5144
rect 33668 5104 35596 5144
rect 35636 5104 35645 5144
rect 38035 5104 38044 5144
rect 38084 5104 39264 5144
rect 39174 5084 39264 5104
rect 7276 4852 8140 4892
rect 8180 4852 8189 4892
rect 8428 4852 8812 4892
rect 8852 4852 8861 4892
rect 8908 4852 9292 4892
rect 9332 4852 9341 4892
rect 9388 4852 11636 4892
rect 11683 4852 11692 4892
rect 11732 4852 23060 4892
rect 24364 4936 25708 4976
rect 25748 4936 25757 4976
rect 26179 4936 26188 4976
rect 26228 4936 26237 4976
rect 28099 4936 28108 4976
rect 28148 4936 30028 4976
rect 30068 4936 30077 4976
rect 31267 4936 31276 4976
rect 31316 4936 31325 4976
rect 31372 4936 33388 4976
rect 33428 4936 33437 4976
rect 37356 4936 37420 4976
rect 37460 4936 37516 4976
rect 37556 4936 37591 4976
rect 37673 4936 37708 4976
rect 37748 4936 37804 4976
rect 37844 4936 37853 4976
rect 0 4808 90 4828
rect 9388 4808 9428 4852
rect 11596 4808 11636 4852
rect 24364 4808 24404 4936
rect 31372 4892 31412 4936
rect 31363 4852 31372 4892
rect 31412 4852 31421 4892
rect 39174 4808 39264 4828
rect 0 4768 364 4808
rect 404 4768 413 4808
rect 2860 4768 9428 4808
rect 10003 4768 10012 4808
rect 10052 4768 11540 4808
rect 11596 4768 24404 4808
rect 37651 4768 37660 4808
rect 37700 4768 39264 4808
rect 0 4748 90 4768
rect 2860 4640 2900 4768
rect 11500 4724 11540 4768
rect 39174 4748 39264 4768
rect 7507 4684 7516 4724
rect 7556 4684 8660 4724
rect 8755 4684 8764 4724
rect 8804 4684 9004 4724
rect 9044 4684 9053 4724
rect 9139 4684 9148 4724
rect 9188 4684 9196 4724
rect 9236 4684 9319 4724
rect 9523 4684 9532 4724
rect 9572 4684 10292 4724
rect 11500 4684 13132 4724
rect 13172 4684 13181 4724
rect 13315 4684 13324 4724
rect 13364 4684 17164 4724
rect 17204 4684 17213 4724
rect 17299 4684 17308 4724
rect 17348 4684 17780 4724
rect 17875 4684 17884 4724
rect 17924 4684 18164 4724
rect 18259 4684 18268 4724
rect 18308 4684 20660 4724
rect 22195 4684 22204 4724
rect 22244 4684 22484 4724
rect 22579 4684 22588 4724
rect 22628 4684 25132 4724
rect 25172 4684 25181 4724
rect 25939 4684 25948 4724
rect 25988 4684 26324 4724
rect 26419 4684 26428 4724
rect 26468 4684 27764 4724
rect 31507 4684 31516 4724
rect 31556 4684 32332 4724
rect 32372 4684 32381 4724
rect 1411 4600 1420 4640
rect 1460 4600 2900 4640
rect 8620 4556 8660 4684
rect 10252 4640 10292 4684
rect 8803 4600 8812 4640
rect 8852 4600 9676 4640
rect 9716 4600 9725 4640
rect 10252 4600 12844 4640
rect 12884 4600 12893 4640
rect 4919 4516 4928 4556
rect 4968 4516 5010 4556
rect 5050 4516 5092 4556
rect 5132 4516 5174 4556
rect 5214 4516 5256 4556
rect 5296 4516 5305 4556
rect 8620 4516 12748 4556
rect 12788 4516 12797 4556
rect 0 4472 90 4492
rect 0 4432 268 4472
rect 308 4432 317 4472
rect 2860 4432 11692 4472
rect 11732 4432 11741 4472
rect 13411 4432 13420 4472
rect 13460 4432 16012 4472
rect 16052 4432 16061 4472
rect 16108 4432 16588 4472
rect 16628 4432 16637 4472
rect 0 4412 90 4432
rect 2860 4388 2900 4432
rect 16108 4388 16148 4432
rect 1315 4348 1324 4388
rect 1364 4348 2900 4388
rect 8995 4348 9004 4388
rect 9044 4348 13036 4388
rect 13076 4348 13085 4388
rect 14467 4348 14476 4388
rect 14516 4348 16148 4388
rect 17740 4388 17780 4684
rect 18124 4472 18164 4684
rect 20620 4556 20660 4684
rect 22444 4640 22484 4684
rect 22444 4600 25516 4640
rect 25556 4600 25565 4640
rect 20039 4516 20048 4556
rect 20088 4516 20130 4556
rect 20170 4516 20212 4556
rect 20252 4516 20294 4556
rect 20334 4516 20376 4556
rect 20416 4516 20425 4556
rect 20620 4516 24556 4556
rect 24596 4516 24605 4556
rect 26284 4472 26324 4684
rect 27724 4640 27764 4684
rect 27724 4600 33196 4640
rect 33236 4600 33245 4640
rect 35159 4516 35168 4556
rect 35208 4516 35250 4556
rect 35290 4516 35332 4556
rect 35372 4516 35414 4556
rect 35454 4516 35496 4556
rect 35536 4516 35545 4556
rect 39174 4472 39264 4492
rect 18124 4432 21292 4472
rect 21332 4432 21341 4472
rect 26284 4432 37612 4472
rect 37652 4432 37661 4472
rect 38668 4432 39264 4472
rect 17740 4348 21100 4388
rect 21140 4348 21149 4388
rect 21676 4348 23212 4388
rect 23252 4348 23261 4388
rect 26131 4348 26140 4388
rect 26180 4348 26708 4388
rect 21676 4304 21716 4348
rect 26668 4304 26708 4348
rect 38668 4304 38708 4432
rect 39174 4412 39264 4432
rect 10051 4264 10060 4304
rect 10100 4264 12980 4304
rect 13267 4264 13276 4304
rect 13316 4264 14284 4304
rect 14324 4264 14333 4304
rect 18643 4264 18652 4304
rect 18692 4264 21716 4304
rect 22483 4264 22492 4304
rect 22532 4264 23500 4304
rect 23540 4264 23549 4304
rect 23635 4264 23644 4304
rect 23684 4264 26572 4304
rect 26612 4264 26621 4304
rect 26668 4264 27052 4304
rect 27092 4264 27101 4304
rect 32393 4264 32476 4304
rect 32516 4264 32524 4304
rect 32564 4264 32573 4304
rect 32777 4264 32860 4304
rect 32900 4264 32908 4304
rect 32948 4264 32957 4304
rect 38035 4264 38044 4304
rect 38084 4264 38708 4304
rect 8515 4180 8524 4220
rect 8564 4180 10004 4220
rect 10819 4180 10828 4220
rect 10868 4180 12692 4220
rect 0 4136 90 4156
rect 9964 4136 10004 4180
rect 12652 4136 12692 4180
rect 12940 4136 12980 4264
rect 13123 4180 13132 4220
rect 13172 4180 13844 4220
rect 14083 4180 14092 4220
rect 14132 4180 16916 4220
rect 13804 4136 13844 4180
rect 16876 4136 16916 4180
rect 19468 4180 22444 4220
rect 22484 4180 22493 4220
rect 22627 4180 22636 4220
rect 22676 4180 27284 4220
rect 30979 4180 30988 4220
rect 31028 4180 32660 4220
rect 33475 4180 33484 4220
rect 33524 4180 37460 4220
rect 19468 4136 19508 4180
rect 27244 4136 27284 4180
rect 32620 4136 32660 4180
rect 37420 4136 37460 4180
rect 39174 4136 39264 4156
rect 0 4096 172 4136
rect 212 4096 221 4136
rect 7555 4096 7564 4136
rect 7604 4096 8236 4136
rect 8276 4096 8285 4136
rect 8611 4096 8620 4136
rect 8660 4096 8669 4136
rect 9955 4096 9964 4136
rect 10004 4096 10013 4136
rect 10339 4096 10348 4136
rect 10388 4096 10397 4136
rect 11203 4096 11212 4136
rect 11252 4096 11884 4136
rect 11924 4096 11933 4136
rect 11980 4096 12268 4136
rect 12308 4096 12317 4136
rect 12643 4096 12652 4136
rect 12692 4096 12701 4136
rect 12940 4096 13036 4136
rect 13076 4096 13085 4136
rect 13289 4096 13420 4136
rect 13460 4096 13469 4136
rect 13795 4096 13804 4136
rect 13844 4096 13853 4136
rect 14249 4096 14380 4136
rect 14420 4096 14429 4136
rect 15977 4096 16108 4136
rect 16148 4096 16157 4136
rect 16483 4096 16492 4136
rect 16532 4096 16684 4136
rect 16724 4096 16733 4136
rect 16867 4096 16876 4136
rect 16916 4096 16925 4136
rect 17251 4096 17260 4136
rect 17300 4096 17356 4136
rect 17396 4096 17431 4136
rect 17513 4096 17644 4136
rect 17684 4096 17693 4136
rect 17897 4096 18028 4136
rect 18068 4096 18077 4136
rect 18211 4096 18220 4136
rect 18260 4096 18412 4136
rect 18452 4096 18461 4136
rect 18665 4096 18700 4136
rect 18740 4096 18796 4136
rect 18836 4096 18845 4136
rect 19171 4096 19180 4136
rect 19220 4096 19229 4136
rect 19411 4096 19420 4136
rect 19460 4096 19508 4136
rect 19555 4096 19564 4136
rect 19604 4096 19756 4136
rect 19796 4096 19805 4136
rect 20803 4096 20812 4136
rect 20852 4096 21100 4136
rect 21140 4096 21149 4136
rect 21475 4096 21484 4136
rect 21524 4096 21533 4136
rect 21737 4096 21868 4136
rect 21908 4096 21917 4136
rect 22243 4096 22252 4136
rect 22292 4096 22348 4136
rect 22388 4096 22423 4136
rect 22540 4096 22636 4136
rect 22676 4096 22685 4136
rect 22889 4096 22924 4136
rect 22964 4096 23020 4136
rect 23060 4096 23124 4136
rect 23395 4096 23404 4136
rect 23444 4096 23453 4136
rect 23657 4096 23788 4136
rect 23828 4096 23837 4136
rect 24163 4096 24172 4136
rect 24212 4096 24268 4136
rect 24308 4096 24343 4136
rect 25891 4096 25900 4136
rect 25940 4096 26188 4136
rect 26228 4096 26237 4136
rect 27235 4096 27244 4136
rect 27284 4096 27293 4136
rect 28457 4096 28588 4136
rect 28628 4096 28637 4136
rect 29635 4096 29644 4136
rect 29684 4096 29693 4136
rect 29923 4096 29932 4136
rect 29972 4096 31564 4136
rect 31604 4096 31613 4136
rect 31660 4096 32236 4136
rect 32276 4096 32285 4136
rect 32611 4096 32620 4136
rect 32660 4096 32669 4136
rect 32873 4096 33004 4136
rect 33044 4096 33053 4136
rect 35971 4096 35980 4136
rect 36020 4096 37036 4136
rect 37076 4096 37085 4136
rect 37411 4096 37420 4136
rect 37460 4096 37469 4136
rect 37795 4096 37804 4136
rect 37844 4096 37900 4136
rect 37940 4096 37975 4136
rect 38764 4096 39264 4136
rect 0 4076 90 4096
rect 8620 4052 8660 4096
rect 10348 4052 10388 4096
rect 11980 4052 12020 4096
rect 19180 4052 19220 4096
rect 21484 4052 21524 4096
rect 22540 4052 22580 4096
rect 23404 4052 23444 4096
rect 29644 4052 29684 4096
rect 31660 4052 31700 4096
rect 38764 4052 38804 4096
rect 39174 4076 39264 4096
rect 7747 4012 7756 4052
rect 7796 4012 8660 4052
rect 8716 4012 10388 4052
rect 11011 4012 11020 4052
rect 11060 4012 12020 4052
rect 12115 4012 12124 4052
rect 12164 4012 12940 4052
rect 12980 4012 12989 4052
rect 14035 4012 14044 4052
rect 14084 4012 14516 4052
rect 14611 4012 14620 4052
rect 14660 4012 18604 4052
rect 18644 4012 18653 4052
rect 19180 4012 19852 4052
rect 19892 4012 19901 4052
rect 20611 4012 20620 4052
rect 20660 4012 21524 4052
rect 21763 4012 21772 4052
rect 21812 4012 22580 4052
rect 22627 4012 22636 4052
rect 22676 4012 23444 4052
rect 24403 4012 24412 4052
rect 24452 4012 27244 4052
rect 27284 4012 27293 4052
rect 27340 4012 29684 4052
rect 31171 4012 31180 4052
rect 31220 4012 31700 4052
rect 31795 4012 31804 4052
rect 31844 4012 33140 4052
rect 33235 4012 33244 4052
rect 33284 4012 37420 4052
rect 37460 4012 37469 4052
rect 37651 4012 37660 4052
rect 37700 4012 38804 4052
rect 8467 3928 8476 3968
rect 8516 3928 8620 3968
rect 8660 3928 8669 3968
rect 8716 3884 8756 4012
rect 14476 3968 14516 4012
rect 27340 3968 27380 4012
rect 33100 3968 33140 4012
rect 8851 3928 8860 3968
rect 8900 3928 10100 3968
rect 10195 3928 10204 3968
rect 10244 3928 10484 3968
rect 10579 3928 10588 3968
rect 10628 3928 11788 3968
rect 11828 3928 11837 3968
rect 12499 3928 12508 3968
rect 12548 3928 12748 3968
rect 12788 3928 12797 3968
rect 12883 3928 12892 3968
rect 12932 3928 12941 3968
rect 13651 3928 13660 3968
rect 13700 3928 14420 3968
rect 14476 3928 15916 3968
rect 15956 3928 15965 3968
rect 16217 3928 16300 3968
rect 16340 3928 16348 3968
rect 16388 3928 16397 3968
rect 16723 3928 16732 3968
rect 16772 3928 17012 3968
rect 17107 3928 17116 3968
rect 17156 3928 17396 3968
rect 17491 3928 17500 3968
rect 17540 3928 17780 3968
rect 17875 3928 17884 3968
rect 17924 3928 18164 3968
rect 18259 3928 18268 3968
rect 18308 3928 18508 3968
rect 18548 3928 18557 3968
rect 19027 3928 19036 3968
rect 19076 3928 19660 3968
rect 19700 3928 19709 3968
rect 19865 3928 19948 3968
rect 19988 3928 19996 3968
rect 20036 3928 20045 3968
rect 20131 3928 20140 3968
rect 20180 3928 21004 3968
rect 21044 3928 21053 3968
rect 21331 3928 21340 3968
rect 21380 3928 21388 3968
rect 21428 3928 21511 3968
rect 21715 3928 21724 3968
rect 21764 3928 22004 3968
rect 22099 3928 22108 3968
rect 22148 3928 22540 3968
rect 22580 3928 22589 3968
rect 22867 3928 22876 3968
rect 22916 3928 23060 3968
rect 23251 3928 23260 3968
rect 23300 3928 23540 3968
rect 24019 3928 24028 3968
rect 24068 3928 26228 3968
rect 27331 3928 27340 3968
rect 27380 3928 27389 3968
rect 27475 3928 27484 3968
rect 27524 3928 28012 3968
rect 28052 3928 28061 3968
rect 28195 3928 28204 3968
rect 28244 3928 28348 3968
rect 28388 3928 28397 3968
rect 28771 3928 28780 3968
rect 28820 3928 29404 3968
rect 29444 3928 29453 3968
rect 33100 3928 34540 3968
rect 34580 3928 34589 3968
rect 37267 3928 37276 3968
rect 37316 3928 37940 3968
rect 8323 3844 8332 3884
rect 8372 3844 8756 3884
rect 0 3800 90 3820
rect 0 3760 940 3800
rect 980 3760 989 3800
rect 3679 3760 3688 3800
rect 3728 3760 3770 3800
rect 3810 3760 3852 3800
rect 3892 3760 3934 3800
rect 3974 3760 4016 3800
rect 4056 3760 4065 3800
rect 0 3740 90 3760
rect 10060 3548 10100 3928
rect 10444 3632 10484 3928
rect 12892 3884 12932 3928
rect 14380 3884 14420 3928
rect 16972 3884 17012 3928
rect 12892 3844 13804 3884
rect 13844 3844 13853 3884
rect 14380 3844 16780 3884
rect 16820 3844 16829 3884
rect 16972 3844 17164 3884
rect 17204 3844 17213 3884
rect 11587 3676 11596 3716
rect 11636 3676 14380 3716
rect 14420 3676 14429 3716
rect 14851 3676 14860 3716
rect 14900 3676 15820 3716
rect 15860 3676 15869 3716
rect 10444 3592 13516 3632
rect 13556 3592 13565 3632
rect 13699 3592 13708 3632
rect 13748 3592 16684 3632
rect 16724 3592 16733 3632
rect 17356 3548 17396 3928
rect 17740 3632 17780 3928
rect 18124 3716 18164 3928
rect 21964 3884 22004 3928
rect 20035 3844 20044 3884
rect 20084 3844 20908 3884
rect 20948 3844 20957 3884
rect 21964 3844 22732 3884
rect 22772 3844 22781 3884
rect 23020 3800 23060 3928
rect 23500 3884 23540 3928
rect 26188 3884 26228 3928
rect 23500 3844 26092 3884
rect 26132 3844 26141 3884
rect 26188 3844 31564 3884
rect 31604 3844 31613 3884
rect 18799 3760 18808 3800
rect 18848 3760 18890 3800
rect 18930 3760 18972 3800
rect 19012 3760 19054 3800
rect 19094 3760 19136 3800
rect 19176 3760 19185 3800
rect 19651 3760 19660 3800
rect 19700 3760 22828 3800
rect 22868 3760 22877 3800
rect 23020 3760 26476 3800
rect 26516 3760 26525 3800
rect 33919 3760 33928 3800
rect 33968 3760 34010 3800
rect 34050 3760 34092 3800
rect 34132 3760 34174 3800
rect 34214 3760 34256 3800
rect 34296 3760 34305 3800
rect 18124 3676 21484 3716
rect 21524 3676 21533 3716
rect 23491 3676 23500 3716
rect 23540 3676 26284 3716
rect 26324 3676 26333 3716
rect 33100 3676 37844 3716
rect 17740 3592 21196 3632
rect 21236 3592 21245 3632
rect 21379 3592 21388 3632
rect 21428 3592 23884 3632
rect 23924 3592 23933 3632
rect 26659 3592 26668 3632
rect 26708 3592 27580 3632
rect 27620 3592 27629 3632
rect 28387 3592 28396 3632
rect 28436 3592 28924 3632
rect 28964 3592 28973 3632
rect 30115 3592 30124 3632
rect 30164 3592 30844 3632
rect 30884 3592 30893 3632
rect 31843 3592 31852 3632
rect 31892 3592 31996 3632
rect 32036 3592 32045 3632
rect 33100 3548 33140 3676
rect 10060 3508 17260 3548
rect 17300 3508 17309 3548
rect 17356 3508 20140 3548
rect 20180 3508 20189 3548
rect 23020 3508 33140 3548
rect 0 3464 90 3484
rect 23020 3464 23060 3508
rect 37804 3464 37844 3676
rect 37900 3464 37940 3928
rect 39174 3800 39264 3820
rect 38668 3760 39264 3800
rect 38668 3632 38708 3760
rect 39174 3740 39264 3760
rect 38035 3592 38044 3632
rect 38084 3592 38708 3632
rect 39174 3464 39264 3484
rect 0 3424 556 3464
rect 596 3424 605 3464
rect 9859 3424 9868 3464
rect 9908 3424 13036 3464
rect 13076 3424 13085 3464
rect 13411 3424 13420 3464
rect 13460 3424 13469 3464
rect 13651 3424 13660 3464
rect 13700 3424 13996 3464
rect 14036 3424 14045 3464
rect 14179 3424 14188 3464
rect 14228 3424 17740 3464
rect 17780 3424 17789 3464
rect 18115 3424 18124 3464
rect 18164 3424 18173 3464
rect 18307 3424 18316 3464
rect 18356 3424 20524 3464
rect 20564 3424 20573 3464
rect 21379 3424 21388 3464
rect 21428 3424 21868 3464
rect 21908 3424 21917 3464
rect 22121 3424 22252 3464
rect 22292 3424 22301 3464
rect 22348 3424 23060 3464
rect 27811 3424 27820 3464
rect 27860 3424 27869 3464
rect 29155 3424 29164 3464
rect 29204 3424 30412 3464
rect 30452 3424 30461 3464
rect 30595 3424 30604 3464
rect 30644 3424 31084 3464
rect 31124 3424 31133 3464
rect 31747 3424 31756 3464
rect 31796 3424 31805 3464
rect 32323 3424 32332 3464
rect 32372 3424 37420 3464
rect 37460 3424 37469 3464
rect 37795 3424 37804 3464
rect 37844 3424 37853 3464
rect 37900 3424 39264 3464
rect 0 3404 90 3424
rect 13420 3380 13460 3424
rect 18124 3380 18164 3424
rect 10627 3340 10636 3380
rect 10676 3340 13460 3380
rect 13891 3340 13900 3380
rect 13940 3340 18164 3380
rect 18220 3340 19700 3380
rect 19747 3340 19756 3380
rect 19796 3340 21908 3380
rect 18220 3296 18260 3340
rect 19660 3296 19700 3340
rect 21868 3296 21908 3340
rect 22348 3296 22388 3424
rect 27820 3380 27860 3424
rect 31756 3380 31796 3424
rect 39174 3404 39264 3424
rect 22723 3340 22732 3380
rect 22772 3340 26860 3380
rect 26900 3340 26909 3380
rect 27820 3340 30316 3380
rect 30356 3340 30365 3380
rect 30787 3340 30796 3380
rect 30836 3340 31796 3380
rect 10243 3256 10252 3296
rect 10292 3256 13132 3296
rect 13172 3256 13181 3296
rect 13267 3256 13276 3296
rect 13316 3256 14380 3296
rect 14420 3256 14429 3296
rect 14563 3256 14572 3296
rect 14612 3256 17740 3296
rect 17780 3256 17789 3296
rect 17971 3256 17980 3296
rect 18020 3256 18260 3296
rect 18355 3256 18364 3296
rect 18404 3256 19604 3296
rect 19660 3256 21676 3296
rect 21716 3256 21725 3296
rect 21868 3256 22388 3296
rect 22531 3256 22540 3296
rect 22580 3256 25900 3296
rect 25940 3256 25949 3296
rect 19564 3212 19604 3256
rect 12739 3172 12748 3212
rect 12788 3172 14612 3212
rect 19564 3172 21964 3212
rect 22004 3172 22013 3212
rect 22099 3172 22108 3212
rect 22148 3172 22388 3212
rect 22483 3172 22492 3212
rect 22532 3172 25708 3212
rect 25748 3172 25757 3212
rect 37651 3172 37660 3212
rect 37700 3172 37940 3212
rect 0 3128 90 3148
rect 14572 3128 14612 3172
rect 22348 3128 22388 3172
rect 37900 3128 37940 3172
rect 39174 3128 39264 3148
rect 0 3088 1228 3128
rect 1268 3088 1277 3128
rect 8611 3088 8620 3128
rect 8660 3088 14476 3128
rect 14516 3088 14525 3128
rect 14572 3088 19756 3128
rect 19796 3088 19805 3128
rect 19948 3088 21580 3128
rect 21620 3088 21629 3128
rect 22348 3088 24748 3128
rect 24788 3088 24797 3128
rect 37900 3088 39264 3128
rect 0 3068 90 3088
rect 19948 3044 19988 3088
rect 39174 3068 39264 3088
rect 4919 3004 4928 3044
rect 4968 3004 5010 3044
rect 5050 3004 5092 3044
rect 5132 3004 5174 3044
rect 5214 3004 5256 3044
rect 5296 3004 5305 3044
rect 11779 3004 11788 3044
rect 11828 3004 18508 3044
rect 18548 3004 18557 3044
rect 18787 3004 18796 3044
rect 18836 3004 19988 3044
rect 20039 3004 20048 3044
rect 20088 3004 20130 3044
rect 20170 3004 20212 3044
rect 20252 3004 20294 3044
rect 20334 3004 20376 3044
rect 20416 3004 20425 3044
rect 22732 3004 29932 3044
rect 29972 3004 29981 3044
rect 35159 3004 35168 3044
rect 35208 3004 35250 3044
rect 35290 3004 35332 3044
rect 35372 3004 35414 3044
rect 35454 3004 35496 3044
rect 35536 3004 35545 3044
rect 13507 2920 13516 2960
rect 13556 2920 17164 2960
rect 17204 2920 17213 2960
rect 17731 2920 17740 2960
rect 17780 2920 20716 2960
rect 20756 2920 20765 2960
rect 16195 2836 16204 2876
rect 16244 2836 19660 2876
rect 19700 2836 19709 2876
rect 19939 2836 19948 2876
rect 19988 2836 22156 2876
rect 22196 2836 22205 2876
rect 22339 2836 22348 2876
rect 22388 2836 22540 2876
rect 22580 2836 22589 2876
rect 0 2792 90 2812
rect 22732 2792 22772 3004
rect 39174 2792 39264 2812
rect 0 2752 22772 2792
rect 38035 2752 38044 2792
rect 38084 2752 39264 2792
rect 0 2732 90 2752
rect 39174 2732 39264 2752
rect 14467 2668 14476 2708
rect 14516 2668 18452 2708
rect 18499 2668 18508 2708
rect 18548 2668 19988 2708
rect 21283 2668 21292 2708
rect 21332 2668 22820 2708
rect 23011 2668 23020 2708
rect 23060 2668 24308 2708
rect 34531 2668 34540 2708
rect 34580 2668 37844 2708
rect 18412 2624 18452 2668
rect 19948 2624 19988 2668
rect 22780 2624 22820 2668
rect 18019 2584 18028 2624
rect 18068 2584 18124 2624
rect 18164 2584 18199 2624
rect 18403 2584 18412 2624
rect 18452 2584 18461 2624
rect 18787 2584 18796 2624
rect 18836 2584 18845 2624
rect 19171 2584 19180 2624
rect 19220 2584 19229 2624
rect 19555 2584 19564 2624
rect 19604 2584 19660 2624
rect 19700 2584 19735 2624
rect 19939 2584 19948 2624
rect 19988 2584 19997 2624
rect 20131 2584 20140 2624
rect 20180 2584 21388 2624
rect 21428 2584 21437 2624
rect 21545 2584 21676 2624
rect 21716 2584 21725 2624
rect 21929 2584 21964 2624
rect 22004 2584 22060 2624
rect 22100 2584 22109 2624
rect 22313 2584 22444 2624
rect 22484 2584 22493 2624
rect 22762 2584 22771 2624
rect 22811 2584 22820 2624
rect 23203 2584 23212 2624
rect 23252 2584 23383 2624
rect 23587 2584 23596 2624
rect 23636 2584 23645 2624
rect 23971 2584 23980 2624
rect 24020 2584 24029 2624
rect 18796 2540 18836 2584
rect 19180 2540 19220 2584
rect 23596 2540 23636 2584
rect 23980 2540 24020 2584
rect 13027 2500 13036 2540
rect 13076 2500 18836 2540
rect 19084 2500 19220 2540
rect 23500 2500 23636 2540
rect 23884 2500 24020 2540
rect 24268 2540 24308 2668
rect 37804 2624 37844 2668
rect 24355 2584 24364 2624
rect 24404 2584 24535 2624
rect 24617 2584 24748 2624
rect 24788 2584 24797 2624
rect 25001 2584 25132 2624
rect 25172 2584 25181 2624
rect 25385 2584 25516 2624
rect 25556 2584 25565 2624
rect 25769 2584 25900 2624
rect 25940 2584 25949 2624
rect 26153 2584 26284 2624
rect 26324 2584 26333 2624
rect 26537 2584 26668 2624
rect 26708 2584 26717 2624
rect 26921 2584 27052 2624
rect 27092 2584 27101 2624
rect 27427 2584 27436 2624
rect 27476 2584 28204 2624
rect 28244 2584 28253 2624
rect 33187 2584 33196 2624
rect 33236 2584 37036 2624
rect 37076 2584 37085 2624
rect 37289 2584 37420 2624
rect 37460 2584 37469 2624
rect 37795 2584 37804 2624
rect 37844 2584 37853 2624
rect 24268 2500 33140 2540
rect 37651 2500 37660 2540
rect 37700 2500 38708 2540
rect 0 2456 90 2476
rect 0 2416 3532 2456
rect 3572 2416 3581 2456
rect 17657 2416 17740 2456
rect 17780 2416 17788 2456
rect 17828 2416 17837 2456
rect 18041 2416 18124 2456
rect 18164 2416 18172 2456
rect 18212 2416 18221 2456
rect 18425 2416 18508 2456
rect 18548 2416 18556 2456
rect 18596 2416 18605 2456
rect 18691 2416 18700 2456
rect 18740 2416 18940 2456
rect 18980 2416 18989 2456
rect 0 2396 90 2416
rect 19084 2372 19124 2500
rect 19193 2416 19276 2456
rect 19316 2416 19324 2456
rect 19364 2416 19373 2456
rect 19577 2416 19660 2456
rect 19700 2416 19708 2456
rect 19748 2416 19757 2456
rect 21305 2416 21388 2456
rect 21428 2416 21436 2456
rect 21476 2416 21485 2456
rect 21689 2416 21772 2456
rect 21812 2416 21820 2456
rect 21860 2416 21869 2456
rect 22073 2416 22156 2456
rect 22196 2416 22204 2456
rect 22244 2416 22253 2456
rect 22457 2416 22540 2456
rect 22580 2416 22588 2456
rect 22628 2416 22637 2456
rect 22841 2416 22924 2456
rect 22964 2416 22972 2456
rect 23012 2416 23021 2456
rect 23225 2416 23308 2456
rect 23348 2416 23356 2456
rect 23396 2416 23405 2456
rect 23500 2372 23540 2500
rect 23609 2416 23692 2456
rect 23732 2416 23740 2456
rect 23780 2416 23789 2456
rect 16003 2332 16012 2372
rect 16052 2332 19124 2372
rect 23011 2332 23020 2372
rect 23060 2332 23540 2372
rect 3679 2248 3688 2288
rect 3728 2248 3770 2288
rect 3810 2248 3852 2288
rect 3892 2248 3934 2288
rect 3974 2248 4016 2288
rect 4056 2248 4065 2288
rect 17443 2248 17452 2288
rect 17492 2248 18412 2288
rect 18452 2248 18461 2288
rect 18799 2248 18808 2288
rect 18848 2248 18890 2288
rect 18930 2248 18972 2288
rect 19012 2248 19054 2288
rect 19094 2248 19136 2288
rect 19176 2248 19185 2288
rect 19276 2248 20140 2288
rect 20180 2248 20189 2288
rect 19276 2204 19316 2248
rect 23884 2204 23924 2500
rect 23993 2416 24076 2456
rect 24116 2416 24124 2456
rect 24164 2416 24173 2456
rect 24377 2416 24460 2456
rect 24500 2416 24508 2456
rect 24548 2416 24557 2456
rect 24761 2416 24844 2456
rect 24884 2416 24892 2456
rect 24932 2416 24941 2456
rect 25145 2416 25228 2456
rect 25268 2416 25276 2456
rect 25316 2416 25325 2456
rect 25529 2416 25612 2456
rect 25652 2416 25660 2456
rect 25700 2416 25709 2456
rect 25913 2416 25996 2456
rect 26036 2416 26044 2456
rect 26084 2416 26093 2456
rect 26297 2416 26380 2456
rect 26420 2416 26428 2456
rect 26468 2416 26477 2456
rect 26681 2416 26764 2456
rect 26804 2416 26812 2456
rect 26852 2416 26861 2456
rect 27065 2416 27148 2456
rect 27188 2416 27196 2456
rect 27236 2416 27245 2456
rect 33100 2372 33140 2500
rect 38668 2456 38708 2500
rect 39174 2456 39264 2476
rect 37267 2416 37276 2456
rect 37316 2416 38380 2456
rect 38420 2416 38429 2456
rect 38668 2416 39264 2456
rect 39174 2396 39264 2416
rect 33100 2332 37460 2372
rect 33919 2248 33928 2288
rect 33968 2248 34010 2288
rect 34050 2248 34092 2288
rect 34132 2248 34174 2288
rect 34214 2248 34256 2288
rect 34296 2248 34305 2288
rect 14275 2164 14284 2204
rect 14324 2164 18356 2204
rect 18595 2164 18604 2204
rect 18644 2164 19316 2204
rect 21091 2164 21100 2204
rect 21140 2164 23924 2204
rect 23971 2164 23980 2204
rect 24020 2164 33140 2204
rect 0 2120 90 2140
rect 18316 2120 18356 2164
rect 0 2080 12980 2120
rect 17347 2080 17356 2120
rect 17396 2080 18260 2120
rect 18316 2080 21716 2120
rect 22051 2080 22060 2120
rect 22100 2080 22676 2120
rect 23107 2080 23116 2120
rect 23156 2080 23828 2120
rect 24163 2080 24172 2120
rect 24212 2080 25364 2120
rect 0 2060 90 2080
rect 0 1784 90 1804
rect 12940 1784 12980 2080
rect 18220 2036 18260 2080
rect 17827 1996 17836 2036
rect 17876 1996 17972 2036
rect 18220 1996 19028 2036
rect 20707 1996 20716 2036
rect 20756 1996 20803 2036
rect 17932 1952 17972 1996
rect 18988 1952 19028 1996
rect 20716 1952 20756 1996
rect 21676 1952 21716 2080
rect 21955 1996 21964 2036
rect 22004 1996 22012 2036
rect 22052 1996 22135 2036
rect 22636 1952 22676 2080
rect 22723 1996 22732 2036
rect 22772 1996 22781 2036
rect 23011 1996 23020 2036
rect 23060 1996 23164 2036
rect 23204 1996 23213 2036
rect 22732 1952 22772 1996
rect 23788 1952 23828 2080
rect 25324 1952 25364 2080
rect 33100 2036 33140 2164
rect 37420 2120 37460 2332
rect 39174 2120 39264 2140
rect 37420 2080 37844 2120
rect 38035 2080 38044 2120
rect 38084 2080 39264 2120
rect 26179 1996 26188 2036
rect 26228 1996 27004 2036
rect 27044 1996 27053 2036
rect 27235 1996 27244 2036
rect 27284 1996 27668 2036
rect 33100 1996 37076 2036
rect 27628 1952 27668 1996
rect 37036 1952 37076 1996
rect 37804 1952 37844 2080
rect 39174 2060 39264 2080
rect 16579 1912 16588 1952
rect 16628 1912 17068 1952
rect 17108 1912 17117 1952
rect 17443 1912 17452 1952
rect 17492 1912 17548 1952
rect 17588 1912 17623 1952
rect 17866 1912 17875 1952
rect 17915 1912 17972 1952
rect 18211 1912 18220 1952
rect 18260 1912 18316 1952
rect 18356 1912 18391 1952
rect 18508 1912 18604 1952
rect 18644 1912 18653 1952
rect 18979 1912 18988 1952
rect 19028 1912 19037 1952
rect 19241 1912 19372 1952
rect 19412 1912 19421 1952
rect 19625 1912 19756 1952
rect 19796 1912 19805 1952
rect 20009 1912 20044 1952
rect 20084 1912 20140 1952
rect 20180 1912 20189 1952
rect 20707 1912 20716 1952
rect 20756 1912 20765 1952
rect 20969 1912 21004 1952
rect 21044 1912 21100 1952
rect 21140 1912 21149 1952
rect 21475 1912 21484 1952
rect 21524 1912 21533 1952
rect 21676 1912 21868 1952
rect 21908 1912 21917 1952
rect 22243 1912 22252 1952
rect 22292 1912 22301 1952
rect 22627 1912 22636 1952
rect 22676 1912 22685 1952
rect 22732 1912 23020 1952
rect 23060 1912 23069 1952
rect 23395 1912 23404 1952
rect 23444 1912 23453 1952
rect 23779 1912 23788 1952
rect 23828 1912 23837 1952
rect 24041 1912 24172 1952
rect 24212 1912 24221 1952
rect 24425 1912 24556 1952
rect 24596 1912 24605 1952
rect 24809 1912 24940 1952
rect 24980 1912 24989 1952
rect 25315 1912 25324 1952
rect 25364 1912 25373 1952
rect 25577 1912 25708 1952
rect 25748 1912 25757 1952
rect 25961 1912 26092 1952
rect 26132 1912 26141 1952
rect 26345 1912 26476 1952
rect 26516 1912 26525 1952
rect 26729 1912 26860 1952
rect 26900 1912 26909 1952
rect 27235 1912 27244 1952
rect 27284 1912 27293 1952
rect 27619 1912 27628 1952
rect 27668 1912 27677 1952
rect 27881 1912 28012 1952
rect 28052 1912 28061 1952
rect 28387 1912 28396 1952
rect 28436 1912 28780 1952
rect 28820 1912 28829 1952
rect 31555 1912 31564 1952
rect 31604 1912 36652 1952
rect 36692 1912 36701 1952
rect 37027 1912 37036 1952
rect 37076 1912 37085 1952
rect 37411 1912 37420 1952
rect 37460 1912 37612 1952
rect 37652 1912 37661 1952
rect 37795 1912 37804 1952
rect 37844 1912 37853 1952
rect 18508 1868 18548 1912
rect 21484 1868 21524 1912
rect 22252 1868 22292 1912
rect 23404 1868 23444 1912
rect 27244 1868 27284 1912
rect 13219 1828 13228 1868
rect 13268 1828 18548 1868
rect 18700 1828 19564 1868
rect 19604 1828 19613 1868
rect 20515 1828 20524 1868
rect 20564 1828 21524 1868
rect 21667 1828 21676 1868
rect 21716 1828 22292 1868
rect 22819 1828 22828 1868
rect 22868 1828 23444 1868
rect 23971 1828 23980 1868
rect 24020 1828 27284 1868
rect 18700 1784 18740 1828
rect 39174 1784 39264 1804
rect 0 1744 1420 1784
rect 1460 1744 1469 1784
rect 12940 1744 18740 1784
rect 19603 1744 19612 1784
rect 19652 1744 19852 1784
rect 19892 1744 19901 1784
rect 20371 1744 20380 1784
rect 20420 1744 20428 1784
rect 20468 1744 20551 1784
rect 20611 1744 20620 1784
rect 20660 1744 21244 1784
rect 21284 1744 21293 1784
rect 21571 1744 21580 1784
rect 21620 1744 22396 1784
rect 22436 1744 22445 1784
rect 22723 1744 22732 1784
rect 22772 1744 23548 1784
rect 23588 1744 23597 1784
rect 23875 1744 23884 1784
rect 23924 1744 24700 1784
rect 24740 1744 24749 1784
rect 25027 1744 25036 1784
rect 25076 1744 25852 1784
rect 25892 1744 25901 1784
rect 26563 1744 26572 1784
rect 26612 1744 27388 1784
rect 27428 1744 27437 1784
rect 36883 1744 36892 1784
rect 36932 1744 37516 1784
rect 37556 1744 37565 1784
rect 37651 1744 37660 1784
rect 37700 1744 39264 1784
rect 0 1724 90 1744
rect 39174 1724 39264 1744
rect 17299 1660 17308 1700
rect 17348 1660 17548 1700
rect 17588 1660 17597 1700
rect 17683 1660 17692 1700
rect 17732 1660 17932 1700
rect 17972 1660 17981 1700
rect 18067 1660 18076 1700
rect 18116 1660 18316 1700
rect 18356 1660 18365 1700
rect 18451 1660 18460 1700
rect 18500 1660 18604 1700
rect 18644 1660 18653 1700
rect 18835 1660 18844 1700
rect 18884 1660 19084 1700
rect 19124 1660 19133 1700
rect 19219 1660 19228 1700
rect 19268 1660 19468 1700
rect 19508 1660 19517 1700
rect 19865 1660 19948 1700
rect 19988 1660 19996 1700
rect 20036 1660 20045 1700
rect 20467 1660 20476 1700
rect 20516 1660 20524 1700
rect 20564 1660 20647 1700
rect 20803 1660 20812 1700
rect 20852 1660 20860 1700
rect 20900 1660 20983 1700
rect 21091 1660 21100 1700
rect 21140 1660 21628 1700
rect 21668 1660 21677 1700
rect 21955 1660 21964 1700
rect 22004 1660 22780 1700
rect 22820 1660 22829 1700
rect 23107 1660 23116 1700
rect 23156 1660 23932 1700
rect 23972 1660 23981 1700
rect 24076 1660 24316 1700
rect 24356 1660 24365 1700
rect 24460 1660 25084 1700
rect 25124 1660 25133 1700
rect 25228 1660 25468 1700
rect 25508 1660 25517 1700
rect 25612 1660 26236 1700
rect 26276 1660 26285 1700
rect 26380 1660 26620 1700
rect 26660 1660 26669 1700
rect 27148 1660 27772 1700
rect 27812 1660 27821 1700
rect 27916 1660 28156 1700
rect 28196 1660 28205 1700
rect 37267 1660 37276 1700
rect 37316 1660 38284 1700
rect 38324 1660 38333 1700
rect 24076 1616 24116 1660
rect 24460 1616 24500 1660
rect 25228 1616 25268 1660
rect 25612 1616 25652 1660
rect 26380 1616 26420 1660
rect 27148 1616 27188 1660
rect 27916 1616 27956 1660
rect 3523 1576 3532 1616
rect 3572 1576 23444 1616
rect 23491 1576 23500 1616
rect 23540 1576 24116 1616
rect 24259 1576 24268 1616
rect 24308 1576 24500 1616
rect 24643 1576 24652 1616
rect 24692 1576 25268 1616
rect 25411 1576 25420 1616
rect 25460 1576 25652 1616
rect 25795 1576 25804 1616
rect 25844 1576 26420 1616
rect 26947 1576 26956 1616
rect 26996 1576 27188 1616
rect 27331 1576 27340 1616
rect 27380 1576 27956 1616
rect 4919 1492 4928 1532
rect 4968 1492 5010 1532
rect 5050 1492 5092 1532
rect 5132 1492 5174 1532
rect 5214 1492 5256 1532
rect 5296 1492 5305 1532
rect 14371 1492 14380 1532
rect 14420 1492 19988 1532
rect 20039 1492 20048 1532
rect 20088 1492 20130 1532
rect 20170 1492 20212 1532
rect 20252 1492 20294 1532
rect 20334 1492 20376 1532
rect 20416 1492 20425 1532
rect 0 1448 90 1468
rect 19948 1448 19988 1492
rect 23404 1448 23444 1576
rect 24268 1492 33004 1532
rect 33044 1492 33053 1532
rect 35159 1492 35168 1532
rect 35208 1492 35250 1532
rect 35290 1492 35332 1532
rect 35372 1492 35414 1532
rect 35454 1492 35496 1532
rect 35536 1492 35545 1532
rect 24268 1448 24308 1492
rect 39174 1448 39264 1468
rect 0 1408 1324 1448
rect 1364 1408 1373 1448
rect 12355 1408 12364 1448
rect 12404 1408 17644 1448
rect 17684 1408 17693 1448
rect 19948 1408 21676 1448
rect 21716 1408 21725 1448
rect 23404 1408 24308 1448
rect 38371 1408 38380 1448
rect 38420 1408 39264 1448
rect 0 1388 90 1408
rect 39174 1388 39264 1408
rect 12547 1324 12556 1364
rect 12596 1324 18028 1364
rect 18068 1324 18077 1364
rect 15619 1156 15628 1196
rect 15668 1156 20716 1196
rect 20756 1156 20765 1196
rect 0 1112 90 1132
rect 39174 1112 39264 1132
rect 0 1072 1420 1112
rect 1460 1072 1469 1112
rect 16387 1072 16396 1112
rect 16436 1072 21868 1112
rect 21908 1072 21917 1112
rect 37507 1072 37516 1112
rect 37556 1072 39264 1112
rect 0 1052 90 1072
rect 39174 1052 39264 1072
rect 12739 988 12748 1028
rect 12788 988 18220 1028
rect 18260 988 18269 1028
rect 15235 904 15244 944
rect 15284 904 21484 944
rect 21524 904 21533 944
rect 12163 820 12172 860
rect 12212 820 17836 860
rect 17876 820 17885 860
rect 0 776 90 796
rect 39174 776 39264 796
rect 0 736 16108 776
rect 16148 736 16157 776
rect 16771 736 16780 776
rect 16820 736 22828 776
rect 22868 736 22877 776
rect 38275 736 38284 776
rect 38324 736 39264 776
rect 0 716 90 736
rect 39174 716 39264 736
rect 16195 652 16204 692
rect 16244 652 22444 692
rect 22484 652 22493 692
rect 17155 568 17164 608
rect 17204 568 22252 608
rect 22292 568 22301 608
rect 15811 484 15820 524
rect 15860 484 22636 524
rect 22676 484 22685 524
rect 13507 400 13516 440
rect 13556 400 19756 440
rect 19796 400 19805 440
rect 15427 316 15436 356
rect 15476 316 21292 356
rect 21332 316 21341 356
rect 23020 148 26284 188
rect 26324 148 26333 188
rect 23020 104 23060 148
rect 15043 64 15052 104
rect 15092 64 23060 104
<< via2 >>
rect 20524 11152 20564 11192
rect 36940 11152 36980 11192
rect 8620 10816 8660 10856
rect 11404 10816 11444 10856
rect 28012 10816 28052 10856
rect 36364 10816 36404 10856
rect 14572 10732 14612 10772
rect 27148 10732 27188 10772
rect 31660 10732 31700 10772
rect 37804 10732 37844 10772
rect 15340 10648 15380 10688
rect 4928 10564 4968 10604
rect 5010 10564 5050 10604
rect 5092 10564 5132 10604
rect 5174 10564 5214 10604
rect 5256 10564 5296 10604
rect 20048 10564 20088 10604
rect 20130 10564 20170 10604
rect 20212 10564 20252 10604
rect 20294 10564 20334 10604
rect 20376 10564 20416 10604
rect 28684 10564 28724 10604
rect 35168 10564 35208 10604
rect 35250 10564 35290 10604
rect 35332 10564 35372 10604
rect 35414 10564 35454 10604
rect 35496 10564 35536 10604
rect 652 10480 692 10520
rect 14668 10480 14708 10520
rect 2188 10396 2228 10436
rect 3916 10396 3956 10436
rect 5644 10396 5684 10436
rect 7372 10396 7412 10436
rect 9100 10396 9140 10436
rect 10828 10396 10868 10436
rect 12556 10396 12596 10436
rect 14284 10396 14324 10436
rect 16012 10396 16052 10436
rect 17740 10396 17780 10436
rect 19468 10396 19508 10436
rect 21964 10480 22004 10520
rect 37324 10480 37364 10520
rect 21196 10396 21236 10436
rect 22924 10396 22964 10436
rect 24652 10396 24692 10436
rect 26380 10396 26420 10436
rect 28108 10396 28148 10436
rect 29836 10396 29876 10436
rect 31564 10396 31604 10436
rect 33292 10396 33332 10436
rect 35020 10396 35060 10436
rect 36364 10396 36404 10436
rect 36748 10396 36788 10436
rect 22636 10312 22676 10352
rect 20140 10228 20180 10268
rect 25900 10228 25940 10268
rect 28012 10228 28052 10268
rect 2668 10144 2708 10184
rect 4204 10144 4244 10184
rect 5932 10144 5972 10184
rect 7660 10144 7700 10184
rect 14572 10144 14612 10184
rect 19660 10144 19700 10184
rect 19948 10144 19988 10184
rect 23212 10144 23252 10184
rect 26380 10144 26420 10184
rect 26668 10144 26708 10184
rect 28396 10144 28436 10184
rect 30124 10144 30164 10184
rect 31852 10144 31892 10184
rect 32908 10144 32948 10184
rect 37804 10144 37844 10184
rect 5740 10060 5780 10100
rect 15820 10060 15860 10100
rect 24268 10060 24308 10100
rect 32524 10060 32564 10100
rect 35596 10060 35636 10100
rect 14956 9976 14996 10016
rect 21964 9976 22004 10016
rect 37228 9976 37268 10016
rect 38764 9976 38804 10016
rect 16876 9892 16916 9932
rect 28204 9892 28244 9932
rect 3688 9808 3728 9848
rect 3770 9808 3810 9848
rect 3852 9808 3892 9848
rect 3934 9808 3974 9848
rect 4016 9808 4056 9848
rect 18808 9808 18848 9848
rect 18890 9808 18930 9848
rect 18972 9808 19012 9848
rect 19054 9808 19094 9848
rect 19136 9808 19176 9848
rect 24076 9808 24116 9848
rect 29260 9808 29300 9848
rect 33928 9808 33968 9848
rect 34010 9808 34050 9848
rect 34092 9808 34132 9848
rect 34174 9808 34214 9848
rect 34256 9808 34296 9848
rect 15052 9724 15092 9764
rect 17164 9724 17204 9764
rect 24364 9724 24404 9764
rect 24556 9724 24596 9764
rect 29452 9724 29492 9764
rect 37804 9724 37844 9764
rect 10732 9640 10772 9680
rect 36652 9640 36692 9680
rect 36940 9640 36980 9680
rect 37324 9640 37364 9680
rect 8236 9556 8276 9596
rect 18988 9472 19028 9512
rect 21004 9472 21044 9512
rect 21196 9472 21236 9512
rect 24364 9472 24404 9512
rect 27724 9472 27764 9512
rect 37228 9472 37268 9512
rect 37612 9472 37652 9512
rect 38764 9472 38804 9512
rect 844 9388 884 9428
rect 20140 9388 20180 9428
rect 23020 9388 23060 9428
rect 24460 9388 24500 9428
rect 30220 9388 30260 9428
rect 31660 9388 31700 9428
rect 37708 9388 37748 9428
rect 940 9304 980 9344
rect 19468 9304 19508 9344
rect 22924 9304 22964 9344
rect 37900 9304 37940 9344
rect 19180 9220 19220 9260
rect 30796 9220 30836 9260
rect 38668 9220 38708 9260
rect 16588 9136 16628 9176
rect 18796 9136 18836 9176
rect 22924 9136 22964 9176
rect 4928 9052 4968 9092
rect 5010 9052 5050 9092
rect 5092 9052 5132 9092
rect 5174 9052 5214 9092
rect 5256 9052 5296 9092
rect 15724 9052 15764 9092
rect 19660 9052 19700 9092
rect 20048 9052 20088 9092
rect 20130 9052 20170 9092
rect 20212 9052 20252 9092
rect 20294 9052 20334 9092
rect 20376 9052 20416 9092
rect 25804 9052 25844 9092
rect 28972 9052 29012 9092
rect 35168 9052 35208 9092
rect 35250 9052 35290 9092
rect 35332 9052 35372 9092
rect 35414 9052 35454 9092
rect 35496 9052 35536 9092
rect 5740 8884 5780 8924
rect 7660 8884 7700 8924
rect 8236 8884 8276 8924
rect 15820 8884 15860 8924
rect 1420 8800 1460 8840
rect 12940 8800 12980 8840
rect 14380 8800 14420 8840
rect 14956 8800 14996 8840
rect 15340 8800 15380 8840
rect 16876 8800 16916 8840
rect 652 8716 692 8756
rect 10060 8716 10100 8756
rect 25228 8968 25268 9008
rect 27820 8968 27860 9008
rect 29644 8968 29684 9008
rect 30220 8968 30260 9008
rect 18796 8884 18836 8924
rect 20620 8884 20660 8924
rect 30796 8884 30836 8924
rect 37612 8884 37652 8924
rect 21580 8800 21620 8840
rect 22636 8800 22676 8840
rect 25228 8800 25268 8840
rect 37516 8800 37556 8840
rect 17740 8716 17780 8756
rect 21004 8716 21044 8756
rect 23116 8716 23156 8756
rect 5740 8632 5780 8672
rect 6412 8632 6452 8672
rect 8140 8632 8180 8672
rect 13228 8632 13268 8672
rect 14284 8632 14324 8672
rect 14668 8632 14708 8672
rect 15052 8632 15092 8672
rect 15532 8632 15572 8672
rect 15820 8632 15860 8672
rect 16588 8632 16628 8672
rect 17164 8632 17204 8672
rect 18988 8632 19028 8672
rect 19180 8632 19220 8672
rect 19564 8632 19604 8672
rect 20524 8632 20564 8672
rect 21196 8632 21236 8672
rect 24076 8632 24116 8672
rect 24268 8632 24308 8672
rect 24556 8632 24596 8672
rect 25132 8632 25172 8672
rect 17260 8548 17300 8588
rect 38668 8800 38708 8840
rect 25804 8632 25844 8672
rect 26092 8632 26132 8672
rect 27820 8632 27860 8672
rect 28108 8632 28148 8672
rect 28780 8632 28820 8672
rect 29068 8632 29108 8672
rect 33484 8632 33524 8672
rect 36652 8632 36692 8672
rect 39148 8632 39188 8672
rect 19660 8548 19700 8588
rect 24460 8548 24500 8588
rect 27148 8548 27188 8588
rect 13996 8464 14036 8504
rect 17164 8464 17204 8504
rect 19756 8464 19796 8504
rect 28204 8464 28244 8504
rect 2860 8380 2900 8420
rect 15724 8380 15764 8420
rect 3688 8296 3728 8336
rect 3770 8296 3810 8336
rect 3852 8296 3892 8336
rect 3934 8296 3974 8336
rect 4016 8296 4056 8336
rect 18808 8296 18848 8336
rect 18890 8296 18930 8336
rect 18972 8296 19012 8336
rect 19054 8296 19094 8336
rect 19136 8296 19176 8336
rect 33928 8296 33968 8336
rect 34010 8296 34050 8336
rect 34092 8296 34132 8336
rect 34174 8296 34214 8336
rect 34256 8296 34296 8336
rect 28684 8128 28724 8168
rect 39148 8128 39188 8168
rect 10732 8044 10772 8084
rect 11404 8044 11444 8084
rect 13996 8044 14036 8084
rect 2956 7960 2996 8000
rect 28684 7960 28724 8000
rect 8620 7876 8660 7916
rect 4928 7540 4968 7580
rect 5010 7540 5050 7580
rect 5092 7540 5132 7580
rect 5174 7540 5214 7580
rect 5256 7540 5296 7580
rect 20048 7540 20088 7580
rect 20130 7540 20170 7580
rect 20212 7540 20252 7580
rect 20294 7540 20334 7580
rect 20376 7540 20416 7580
rect 35168 7540 35208 7580
rect 35250 7540 35290 7580
rect 35332 7540 35372 7580
rect 35414 7540 35454 7580
rect 35496 7540 35536 7580
rect 13228 7456 13268 7496
rect 6028 7120 6068 7160
rect 14380 7120 14420 7160
rect 5932 7036 5972 7076
rect 17260 7036 17300 7076
rect 21580 7036 21620 7076
rect 8140 6868 8180 6908
rect 3688 6784 3728 6824
rect 3770 6784 3810 6824
rect 3852 6784 3892 6824
rect 3934 6784 3974 6824
rect 4016 6784 4056 6824
rect 18808 6784 18848 6824
rect 18890 6784 18930 6824
rect 18972 6784 19012 6824
rect 19054 6784 19094 6824
rect 19136 6784 19176 6824
rect 33928 6784 33968 6824
rect 34010 6784 34050 6824
rect 34092 6784 34132 6824
rect 34174 6784 34214 6824
rect 34256 6784 34296 6824
rect 2668 6616 2708 6656
rect 23212 6616 23252 6656
rect 22924 6532 22964 6572
rect 844 6448 884 6488
rect 2956 6448 2996 6488
rect 29836 6448 29876 6488
rect 37804 6448 37844 6488
rect 556 6364 596 6404
rect 35980 6196 36020 6236
rect 17164 6112 17204 6152
rect 4928 6028 4968 6068
rect 5010 6028 5050 6068
rect 5092 6028 5132 6068
rect 5174 6028 5214 6068
rect 5256 6028 5296 6068
rect 20048 6028 20088 6068
rect 20130 6028 20170 6068
rect 20212 6028 20252 6068
rect 20294 6028 20334 6068
rect 20376 6028 20416 6068
rect 35168 6028 35208 6068
rect 35250 6028 35290 6068
rect 35332 6028 35372 6068
rect 35414 6028 35454 6068
rect 35496 6028 35536 6068
rect 15532 5776 15572 5816
rect 8812 5692 8852 5732
rect 15820 5692 15860 5732
rect 2668 5608 2708 5648
rect 4204 5608 4244 5648
rect 1228 5524 1268 5564
rect 10060 5608 10100 5648
rect 14284 5608 14324 5648
rect 9196 5524 9236 5564
rect 16972 5524 17012 5564
rect 9868 5440 9908 5480
rect 16876 5440 16916 5480
rect 22348 5440 22388 5480
rect 3688 5272 3728 5312
rect 3770 5272 3810 5312
rect 3852 5272 3892 5312
rect 3934 5272 3974 5312
rect 4016 5272 4056 5312
rect 20140 5356 20180 5396
rect 24172 5356 24212 5396
rect 8908 5272 8948 5312
rect 9964 5272 10004 5312
rect 10156 5272 10196 5312
rect 16204 5272 16244 5312
rect 17836 5272 17876 5312
rect 18808 5272 18848 5312
rect 18890 5272 18930 5312
rect 18972 5272 19012 5312
rect 19054 5272 19094 5312
rect 19136 5272 19176 5312
rect 33928 5272 33968 5312
rect 34010 5272 34050 5312
rect 34092 5272 34132 5312
rect 34174 5272 34214 5312
rect 34256 5272 34296 5312
rect 8812 5188 8852 5228
rect 16492 5188 16532 5228
rect 18220 5188 18260 5228
rect 1420 5104 1460 5144
rect 8716 5104 8756 5144
rect 13036 5104 13076 5144
rect 24940 5188 24980 5228
rect 9484 5020 9524 5060
rect 26380 5104 26420 5144
rect 11884 5020 11924 5060
rect 7948 4936 7988 4976
rect 9100 4936 9140 4976
rect 9964 4936 10004 4976
rect 11404 4936 11444 4976
rect 13420 4936 13460 4976
rect 17068 4936 17108 4976
rect 17260 4936 17300 4976
rect 17932 4936 17972 4976
rect 18220 4936 18260 4976
rect 22348 4936 22388 4976
rect 35596 5104 35636 5144
rect 8140 4852 8180 4892
rect 8812 4852 8852 4892
rect 9292 4852 9332 4892
rect 11692 4852 11732 4892
rect 30028 4936 30068 4976
rect 37516 4936 37556 4976
rect 37708 4936 37748 4976
rect 31372 4852 31412 4892
rect 364 4768 404 4808
rect 9004 4684 9044 4724
rect 9196 4684 9236 4724
rect 13132 4684 13172 4724
rect 13324 4684 13364 4724
rect 17164 4684 17204 4724
rect 25132 4684 25172 4724
rect 32332 4684 32372 4724
rect 1420 4600 1460 4640
rect 8812 4600 8852 4640
rect 9676 4600 9716 4640
rect 12844 4600 12884 4640
rect 4928 4516 4968 4556
rect 5010 4516 5050 4556
rect 5092 4516 5132 4556
rect 5174 4516 5214 4556
rect 5256 4516 5296 4556
rect 12748 4516 12788 4556
rect 268 4432 308 4472
rect 11692 4432 11732 4472
rect 13420 4432 13460 4472
rect 16012 4432 16052 4472
rect 16588 4432 16628 4472
rect 1324 4348 1364 4388
rect 9004 4348 9044 4388
rect 13036 4348 13076 4388
rect 14476 4348 14516 4388
rect 25516 4600 25556 4640
rect 20048 4516 20088 4556
rect 20130 4516 20170 4556
rect 20212 4516 20252 4556
rect 20294 4516 20334 4556
rect 20376 4516 20416 4556
rect 24556 4516 24596 4556
rect 33196 4600 33236 4640
rect 35168 4516 35208 4556
rect 35250 4516 35290 4556
rect 35332 4516 35372 4556
rect 35414 4516 35454 4556
rect 35496 4516 35536 4556
rect 21292 4432 21332 4472
rect 37612 4432 37652 4472
rect 21100 4348 21140 4388
rect 23212 4348 23252 4388
rect 10060 4264 10100 4304
rect 14284 4264 14324 4304
rect 23500 4264 23540 4304
rect 26572 4264 26612 4304
rect 27052 4264 27092 4304
rect 32524 4264 32564 4304
rect 32908 4264 32948 4304
rect 8524 4180 8564 4220
rect 10828 4180 10868 4220
rect 13132 4180 13172 4220
rect 14092 4180 14132 4220
rect 22444 4180 22484 4220
rect 22636 4180 22676 4220
rect 30988 4180 31028 4220
rect 33484 4180 33524 4220
rect 172 4096 212 4136
rect 7564 4096 7604 4136
rect 11212 4096 11252 4136
rect 13420 4096 13460 4136
rect 14380 4096 14420 4136
rect 16108 4096 16148 4136
rect 16684 4096 16724 4136
rect 17356 4096 17396 4136
rect 17644 4096 17684 4136
rect 18028 4096 18068 4136
rect 18220 4096 18260 4136
rect 18700 4096 18740 4136
rect 19564 4096 19604 4136
rect 20812 4096 20852 4136
rect 21868 4096 21908 4136
rect 22348 4096 22388 4136
rect 22924 4096 22964 4136
rect 23788 4096 23828 4136
rect 24268 4096 24308 4136
rect 26188 4096 26228 4136
rect 28588 4096 28628 4136
rect 29932 4096 29972 4136
rect 33004 4096 33044 4136
rect 35980 4096 36020 4136
rect 37900 4096 37940 4136
rect 7756 4012 7796 4052
rect 11020 4012 11060 4052
rect 12940 4012 12980 4052
rect 18604 4012 18644 4052
rect 19852 4012 19892 4052
rect 20620 4012 20660 4052
rect 21772 4012 21812 4052
rect 22636 4012 22676 4052
rect 27244 4012 27284 4052
rect 31180 4012 31220 4052
rect 37420 4012 37460 4052
rect 8620 3928 8660 3968
rect 11788 3928 11828 3968
rect 12748 3928 12788 3968
rect 15916 3928 15956 3968
rect 16300 3928 16340 3968
rect 18508 3928 18548 3968
rect 19660 3928 19700 3968
rect 19948 3928 19988 3968
rect 20140 3928 20180 3968
rect 21004 3928 21044 3968
rect 21388 3928 21428 3968
rect 22540 3928 22580 3968
rect 27340 3928 27380 3968
rect 28012 3928 28052 3968
rect 28204 3928 28244 3968
rect 28780 3928 28820 3968
rect 34540 3928 34580 3968
rect 8332 3844 8372 3884
rect 940 3760 980 3800
rect 3688 3760 3728 3800
rect 3770 3760 3810 3800
rect 3852 3760 3892 3800
rect 3934 3760 3974 3800
rect 4016 3760 4056 3800
rect 13804 3844 13844 3884
rect 16780 3844 16820 3884
rect 17164 3844 17204 3884
rect 11596 3676 11636 3716
rect 14380 3676 14420 3716
rect 14860 3676 14900 3716
rect 15820 3676 15860 3716
rect 13516 3592 13556 3632
rect 13708 3592 13748 3632
rect 16684 3592 16724 3632
rect 20044 3844 20084 3884
rect 20908 3844 20948 3884
rect 22732 3844 22772 3884
rect 26092 3844 26132 3884
rect 31564 3844 31604 3884
rect 18808 3760 18848 3800
rect 18890 3760 18930 3800
rect 18972 3760 19012 3800
rect 19054 3760 19094 3800
rect 19136 3760 19176 3800
rect 19660 3760 19700 3800
rect 22828 3760 22868 3800
rect 26476 3760 26516 3800
rect 33928 3760 33968 3800
rect 34010 3760 34050 3800
rect 34092 3760 34132 3800
rect 34174 3760 34214 3800
rect 34256 3760 34296 3800
rect 21484 3676 21524 3716
rect 23500 3676 23540 3716
rect 26284 3676 26324 3716
rect 21196 3592 21236 3632
rect 21388 3592 21428 3632
rect 23884 3592 23924 3632
rect 26668 3592 26708 3632
rect 28396 3592 28436 3632
rect 30124 3592 30164 3632
rect 31852 3592 31892 3632
rect 17260 3508 17300 3548
rect 20140 3508 20180 3548
rect 556 3424 596 3464
rect 9868 3424 9908 3464
rect 13996 3424 14036 3464
rect 14188 3424 14228 3464
rect 18316 3424 18356 3464
rect 20524 3424 20564 3464
rect 21388 3424 21428 3464
rect 22252 3424 22292 3464
rect 30412 3424 30452 3464
rect 30604 3424 30644 3464
rect 32332 3424 32372 3464
rect 10636 3340 10676 3380
rect 13900 3340 13940 3380
rect 19756 3340 19796 3380
rect 22732 3340 22772 3380
rect 26860 3340 26900 3380
rect 30316 3340 30356 3380
rect 30796 3340 30836 3380
rect 10252 3256 10292 3296
rect 13132 3256 13172 3296
rect 14380 3256 14420 3296
rect 14572 3256 14612 3296
rect 17740 3256 17780 3296
rect 21676 3256 21716 3296
rect 22540 3256 22580 3296
rect 25900 3256 25940 3296
rect 12748 3172 12788 3212
rect 21964 3172 22004 3212
rect 25708 3172 25748 3212
rect 1228 3088 1268 3128
rect 8620 3088 8660 3128
rect 14476 3088 14516 3128
rect 19756 3088 19796 3128
rect 21580 3088 21620 3128
rect 24748 3088 24788 3128
rect 4928 3004 4968 3044
rect 5010 3004 5050 3044
rect 5092 3004 5132 3044
rect 5174 3004 5214 3044
rect 5256 3004 5296 3044
rect 11788 3004 11828 3044
rect 18508 3004 18548 3044
rect 18796 3004 18836 3044
rect 20048 3004 20088 3044
rect 20130 3004 20170 3044
rect 20212 3004 20252 3044
rect 20294 3004 20334 3044
rect 20376 3004 20416 3044
rect 29932 3004 29972 3044
rect 35168 3004 35208 3044
rect 35250 3004 35290 3044
rect 35332 3004 35372 3044
rect 35414 3004 35454 3044
rect 35496 3004 35536 3044
rect 13516 2920 13556 2960
rect 17164 2920 17204 2960
rect 17740 2920 17780 2960
rect 20716 2920 20756 2960
rect 16204 2836 16244 2876
rect 19660 2836 19700 2876
rect 19948 2836 19988 2876
rect 22156 2836 22196 2876
rect 22348 2836 22388 2876
rect 22540 2836 22580 2876
rect 14476 2668 14516 2708
rect 18508 2668 18548 2708
rect 21292 2668 21332 2708
rect 23020 2668 23060 2708
rect 34540 2668 34580 2708
rect 18124 2584 18164 2624
rect 19660 2584 19700 2624
rect 20140 2584 20180 2624
rect 21388 2584 21428 2624
rect 21676 2584 21716 2624
rect 21964 2584 22004 2624
rect 22444 2584 22484 2624
rect 23212 2584 23252 2624
rect 13036 2500 13076 2540
rect 24364 2584 24404 2624
rect 24748 2584 24788 2624
rect 25132 2584 25172 2624
rect 25516 2584 25556 2624
rect 25900 2584 25940 2624
rect 26284 2584 26324 2624
rect 26668 2584 26708 2624
rect 27052 2584 27092 2624
rect 28204 2584 28244 2624
rect 33196 2584 33236 2624
rect 37420 2584 37460 2624
rect 3532 2416 3572 2456
rect 17740 2416 17780 2456
rect 18124 2416 18164 2456
rect 18508 2416 18548 2456
rect 18700 2416 18740 2456
rect 19276 2416 19316 2456
rect 19660 2416 19700 2456
rect 21388 2416 21428 2456
rect 21772 2416 21812 2456
rect 22156 2416 22196 2456
rect 22540 2416 22580 2456
rect 22924 2416 22964 2456
rect 23308 2416 23348 2456
rect 23692 2416 23732 2456
rect 16012 2332 16052 2372
rect 23020 2332 23060 2372
rect 3688 2248 3728 2288
rect 3770 2248 3810 2288
rect 3852 2248 3892 2288
rect 3934 2248 3974 2288
rect 4016 2248 4056 2288
rect 17452 2248 17492 2288
rect 18412 2248 18452 2288
rect 18808 2248 18848 2288
rect 18890 2248 18930 2288
rect 18972 2248 19012 2288
rect 19054 2248 19094 2288
rect 19136 2248 19176 2288
rect 20140 2248 20180 2288
rect 24076 2416 24116 2456
rect 24460 2416 24500 2456
rect 24844 2416 24884 2456
rect 25228 2416 25268 2456
rect 25612 2416 25652 2456
rect 25996 2416 26036 2456
rect 26380 2416 26420 2456
rect 26764 2416 26804 2456
rect 27148 2416 27188 2456
rect 38380 2416 38420 2456
rect 33928 2248 33968 2288
rect 34010 2248 34050 2288
rect 34092 2248 34132 2288
rect 34174 2248 34214 2288
rect 34256 2248 34296 2288
rect 14284 2164 14324 2204
rect 18604 2164 18644 2204
rect 21100 2164 21140 2204
rect 23980 2164 24020 2204
rect 17356 2080 17396 2120
rect 22060 2080 22100 2120
rect 23116 2080 23156 2120
rect 24172 2080 24212 2120
rect 17836 1996 17876 2036
rect 20716 1996 20756 2036
rect 21964 1996 22004 2036
rect 22732 1996 22772 2036
rect 23020 1996 23060 2036
rect 26188 1996 26228 2036
rect 27244 1996 27284 2036
rect 16588 1912 16628 1952
rect 17548 1912 17588 1952
rect 18316 1912 18356 1952
rect 19372 1912 19412 1952
rect 19756 1912 19796 1952
rect 20044 1912 20084 1952
rect 21004 1912 21044 1952
rect 24172 1912 24212 1952
rect 24556 1912 24596 1952
rect 24940 1912 24980 1952
rect 25708 1912 25748 1952
rect 26092 1912 26132 1952
rect 26476 1912 26516 1952
rect 26860 1912 26900 1952
rect 28012 1912 28052 1952
rect 28780 1912 28820 1952
rect 31564 1912 31604 1952
rect 37612 1912 37652 1952
rect 13228 1828 13268 1868
rect 19564 1828 19604 1868
rect 20524 1828 20564 1868
rect 21676 1828 21716 1868
rect 22828 1828 22868 1868
rect 23980 1828 24020 1868
rect 1420 1744 1460 1784
rect 19852 1744 19892 1784
rect 20428 1744 20468 1784
rect 20620 1744 20660 1784
rect 21580 1744 21620 1784
rect 22732 1744 22772 1784
rect 23884 1744 23924 1784
rect 25036 1744 25076 1784
rect 26572 1744 26612 1784
rect 37516 1744 37556 1784
rect 17548 1660 17588 1700
rect 17932 1660 17972 1700
rect 18316 1660 18356 1700
rect 18604 1660 18644 1700
rect 19084 1660 19124 1700
rect 19468 1660 19508 1700
rect 19948 1660 19988 1700
rect 20524 1660 20564 1700
rect 20812 1660 20852 1700
rect 21100 1660 21140 1700
rect 21964 1660 22004 1700
rect 23116 1660 23156 1700
rect 38284 1660 38324 1700
rect 3532 1576 3572 1616
rect 23500 1576 23540 1616
rect 24268 1576 24308 1616
rect 24652 1576 24692 1616
rect 25420 1576 25460 1616
rect 25804 1576 25844 1616
rect 26956 1576 26996 1616
rect 27340 1576 27380 1616
rect 4928 1492 4968 1532
rect 5010 1492 5050 1532
rect 5092 1492 5132 1532
rect 5174 1492 5214 1532
rect 5256 1492 5296 1532
rect 14380 1492 14420 1532
rect 20048 1492 20088 1532
rect 20130 1492 20170 1532
rect 20212 1492 20252 1532
rect 20294 1492 20334 1532
rect 20376 1492 20416 1532
rect 33004 1492 33044 1532
rect 35168 1492 35208 1532
rect 35250 1492 35290 1532
rect 35332 1492 35372 1532
rect 35414 1492 35454 1532
rect 35496 1492 35536 1532
rect 1324 1408 1364 1448
rect 12364 1408 12404 1448
rect 17644 1408 17684 1448
rect 21676 1408 21716 1448
rect 38380 1408 38420 1448
rect 12556 1324 12596 1364
rect 18028 1324 18068 1364
rect 15628 1156 15668 1196
rect 20716 1156 20756 1196
rect 1420 1072 1460 1112
rect 16396 1072 16436 1112
rect 21868 1072 21908 1112
rect 37516 1072 37556 1112
rect 12748 988 12788 1028
rect 18220 988 18260 1028
rect 15244 904 15284 944
rect 21484 904 21524 944
rect 12172 820 12212 860
rect 17836 820 17876 860
rect 16108 736 16148 776
rect 16780 736 16820 776
rect 22828 736 22868 776
rect 38284 736 38324 776
rect 16204 652 16244 692
rect 22444 652 22484 692
rect 17164 568 17204 608
rect 22252 568 22292 608
rect 15820 484 15860 524
rect 22636 484 22676 524
rect 13516 400 13556 440
rect 19756 400 19796 440
rect 15436 316 15476 356
rect 21292 316 21332 356
rect 26284 148 26324 188
rect 15052 64 15092 104
<< metal3 >>
rect 2168 12100 2248 12180
rect 3896 12100 3976 12180
rect 5624 12100 5704 12180
rect 7352 12100 7432 12180
rect 9080 12100 9160 12180
rect 10808 12100 10888 12180
rect 12536 12100 12616 12180
rect 14264 12100 14344 12180
rect 15992 12100 16072 12180
rect 17720 12100 17800 12180
rect 19448 12100 19528 12180
rect 21176 12100 21256 12180
rect 22904 12100 22984 12180
rect 24632 12100 24712 12180
rect 26360 12100 26440 12180
rect 28088 12100 28168 12180
rect 29816 12100 29896 12180
rect 31544 12100 31624 12180
rect 33272 12100 33352 12180
rect 35000 12100 35080 12180
rect 36728 12100 36808 12180
rect 652 10520 692 10529
rect 364 8840 404 8849
rect 268 8756 308 8765
rect 172 8672 212 8681
rect 172 4136 212 8632
rect 268 4472 308 8716
rect 364 4808 404 8800
rect 652 8756 692 10480
rect 2188 10436 2228 12100
rect 2188 10387 2228 10396
rect 3916 10436 3956 12100
rect 4928 10604 5296 10613
rect 4968 10564 5010 10604
rect 5050 10564 5092 10604
rect 5132 10564 5174 10604
rect 5214 10564 5256 10604
rect 4928 10555 5296 10564
rect 3916 10387 3956 10396
rect 5644 10436 5684 12100
rect 5644 10387 5684 10396
rect 7372 10436 7412 12100
rect 7372 10387 7412 10396
rect 8620 10856 8660 10865
rect 2668 10184 2708 10193
rect 652 8707 692 8716
rect 844 9428 884 9437
rect 844 6488 884 9388
rect 844 6439 884 6448
rect 940 9344 980 9353
rect 364 4759 404 4768
rect 556 6404 596 6413
rect 268 4423 308 4432
rect 172 4087 212 4096
rect 556 3464 596 6364
rect 940 3800 980 9304
rect 1420 8840 1460 8849
rect 940 3751 980 3760
rect 1228 5564 1268 5573
rect 556 3415 596 3424
rect 1228 3128 1268 5524
rect 1420 5144 1460 8800
rect 2668 6656 2708 10144
rect 4204 10184 4244 10193
rect 3688 9848 4056 9857
rect 3728 9808 3770 9848
rect 3810 9808 3852 9848
rect 3892 9808 3934 9848
rect 3974 9808 4016 9848
rect 3688 9799 4056 9808
rect 2860 8420 2900 8429
rect 2900 8380 2996 8420
rect 2860 8371 2900 8380
rect 2956 8000 2996 8380
rect 3688 8336 4056 8345
rect 3728 8296 3770 8336
rect 3810 8296 3852 8336
rect 3892 8296 3934 8336
rect 3974 8296 4016 8336
rect 3688 8287 4056 8296
rect 2956 7951 2996 7960
rect 3688 6824 4056 6833
rect 3728 6784 3770 6824
rect 3810 6784 3852 6824
rect 3892 6784 3934 6824
rect 3974 6784 4016 6824
rect 3688 6775 4056 6784
rect 2668 6607 2708 6616
rect 2956 6488 2996 6497
rect 1420 5095 1460 5104
rect 2668 5648 2708 5657
rect 1420 4640 1460 4649
rect 1228 3079 1268 3088
rect 1324 4388 1364 4397
rect 1324 1448 1364 4348
rect 1420 1784 1460 4600
rect 1420 1735 1460 1744
rect 1324 1399 1364 1408
rect 1420 1112 1460 1121
rect 1420 977 1460 1072
rect 2668 188 2708 5608
rect 2956 2900 2996 6448
rect 4204 5648 4244 10144
rect 5932 10184 5972 10193
rect 5740 10100 5780 10109
rect 4928 9092 5296 9101
rect 4968 9052 5010 9092
rect 5050 9052 5092 9092
rect 5132 9052 5174 9092
rect 5214 9052 5256 9092
rect 4928 9043 5296 9052
rect 5740 8924 5780 10060
rect 5740 8875 5780 8884
rect 5740 8672 5780 8681
rect 4928 7580 5296 7589
rect 4968 7540 5010 7580
rect 5050 7540 5092 7580
rect 5132 7540 5174 7580
rect 5214 7540 5256 7580
rect 4928 7531 5296 7540
rect 4928 6068 5296 6077
rect 4968 6028 5010 6068
rect 5050 6028 5092 6068
rect 5132 6028 5174 6068
rect 5214 6028 5256 6068
rect 4928 6019 5296 6028
rect 4204 5599 4244 5608
rect 3688 5312 4056 5321
rect 3728 5272 3770 5312
rect 3810 5272 3852 5312
rect 3892 5272 3934 5312
rect 3974 5272 4016 5312
rect 3688 5263 4056 5272
rect 4928 4556 5296 4565
rect 4968 4516 5010 4556
rect 5050 4516 5092 4556
rect 5132 4516 5174 4556
rect 5214 4516 5256 4556
rect 4928 4507 5296 4516
rect 3688 3800 4056 3809
rect 3728 3760 3770 3800
rect 3810 3760 3852 3800
rect 3892 3760 3934 3800
rect 3974 3760 4016 3800
rect 3688 3751 4056 3760
rect 4928 3044 5296 3053
rect 4968 3004 5010 3044
rect 5050 3004 5092 3044
rect 5132 3004 5174 3044
rect 5214 3004 5256 3044
rect 4928 2995 5296 3004
rect 2668 139 2708 148
rect 2860 2860 2996 2900
rect 2860 104 2900 2860
rect 3532 2456 3572 2465
rect 3532 1616 3572 2416
rect 3688 2288 4056 2297
rect 3728 2248 3770 2288
rect 3810 2248 3852 2288
rect 3892 2248 3934 2288
rect 3974 2248 4016 2288
rect 3688 2239 4056 2248
rect 3532 1567 3572 1576
rect 4928 1532 5296 1541
rect 4968 1492 5010 1532
rect 5050 1492 5092 1532
rect 5132 1492 5174 1532
rect 5214 1492 5256 1532
rect 4928 1483 5296 1492
rect 5740 272 5780 8632
rect 5932 7076 5972 10144
rect 7660 10184 7700 10193
rect 7660 8924 7700 10144
rect 7660 8875 7700 8884
rect 8236 9596 8276 9605
rect 8236 8924 8276 9556
rect 8236 8875 8276 8884
rect 6412 8672 6452 8681
rect 5932 7027 5972 7036
rect 6028 7160 6068 7169
rect 6028 356 6068 7120
rect 6412 440 6452 8632
rect 8140 8672 8180 8681
rect 8140 6908 8180 8632
rect 8620 7916 8660 10816
rect 9100 10436 9140 12100
rect 9100 10387 9140 10396
rect 10828 10436 10868 12100
rect 10828 10387 10868 10396
rect 11404 10856 11444 10865
rect 10732 9680 10772 9689
rect 8620 7867 8660 7876
rect 10060 8756 10100 8765
rect 8140 6859 8180 6868
rect 8812 5732 8852 5741
rect 8812 5228 8852 5692
rect 10060 5648 10100 8716
rect 10732 8084 10772 9640
rect 10732 8035 10772 8044
rect 11404 8084 11444 10816
rect 12556 10436 12596 12100
rect 12556 10387 12596 10396
rect 14284 10436 14324 12100
rect 14284 10387 14324 10396
rect 14572 10772 14612 10781
rect 14572 10184 14612 10732
rect 15340 10688 15380 10697
rect 14572 10135 14612 10144
rect 14668 10520 14708 10529
rect 12940 8924 12980 8933
rect 12940 8840 12980 8884
rect 12940 8789 12980 8800
rect 14380 8840 14420 8849
rect 11404 8035 11444 8044
rect 13228 8672 13268 8681
rect 13228 7496 13268 8632
rect 14284 8672 14324 8681
rect 13996 8504 14036 8513
rect 13996 8084 14036 8464
rect 13996 8035 14036 8044
rect 13228 7447 13268 7456
rect 10060 5599 10100 5608
rect 14284 5648 14324 8632
rect 14380 7160 14420 8800
rect 14668 8672 14708 10480
rect 14956 10016 14996 10025
rect 14956 8840 14996 9976
rect 14956 8791 14996 8800
rect 15052 9764 15092 9773
rect 14668 8623 14708 8632
rect 15052 8672 15092 9724
rect 15340 8840 15380 10648
rect 16012 10436 16052 12100
rect 16012 10387 16052 10396
rect 17740 10436 17780 12100
rect 17740 10387 17780 10396
rect 19468 10436 19508 12100
rect 20524 11192 20564 11201
rect 20048 10604 20416 10613
rect 20088 10564 20130 10604
rect 20170 10564 20212 10604
rect 20252 10564 20294 10604
rect 20334 10564 20376 10604
rect 20048 10555 20416 10564
rect 19468 10387 19508 10396
rect 20140 10268 20180 10277
rect 19660 10184 19700 10193
rect 19948 10184 19988 10193
rect 19700 10144 19948 10184
rect 19660 10135 19700 10144
rect 19948 10135 19988 10144
rect 15820 10100 15860 10109
rect 15340 8791 15380 8800
rect 15724 9092 15764 9101
rect 15052 8623 15092 8632
rect 15532 8672 15572 8681
rect 14380 7111 14420 7120
rect 15532 5816 15572 8632
rect 15724 8420 15764 9052
rect 15820 8924 15860 10060
rect 16876 9932 16916 9941
rect 15820 8875 15860 8884
rect 16588 9176 16628 9185
rect 15724 8371 15764 8380
rect 15820 8672 15860 8681
rect 15532 5767 15572 5776
rect 15820 5732 15860 8632
rect 16588 8672 16628 9136
rect 16876 8840 16916 9892
rect 18808 9848 19176 9857
rect 18848 9808 18890 9848
rect 18930 9808 18972 9848
rect 19012 9808 19054 9848
rect 19094 9808 19136 9848
rect 18808 9799 19176 9808
rect 16876 8791 16916 8800
rect 17164 9764 17204 9773
rect 16588 8623 16628 8632
rect 17164 8672 17204 9724
rect 18988 9512 19028 9521
rect 18796 9176 18836 9185
rect 17740 8924 17780 8933
rect 17740 8756 17780 8884
rect 18796 8924 18836 9136
rect 18796 8875 18836 8884
rect 17740 8707 17780 8716
rect 17164 8623 17204 8632
rect 18988 8672 19028 9472
rect 20140 9428 20180 10228
rect 20140 9379 20180 9388
rect 19468 9344 19508 9353
rect 19508 9304 19604 9344
rect 19468 9295 19508 9304
rect 18988 8623 19028 8632
rect 19180 9260 19220 9269
rect 19180 8672 19220 9220
rect 19180 8623 19220 8632
rect 19564 8672 19604 9304
rect 19564 8623 19604 8632
rect 19660 9092 19700 9101
rect 17260 8588 17300 8597
rect 17164 8504 17204 8513
rect 17164 6152 17204 8464
rect 17260 7076 17300 8548
rect 19660 8588 19700 9052
rect 20048 9092 20416 9101
rect 20088 9052 20130 9092
rect 20170 9052 20212 9092
rect 20252 9052 20294 9092
rect 20334 9052 20376 9092
rect 20048 9043 20416 9052
rect 20524 8672 20564 11152
rect 21196 10436 21236 12100
rect 21196 10387 21236 10396
rect 21964 10520 22004 10529
rect 21964 10016 22004 10480
rect 22924 10436 22964 12100
rect 22924 10387 22964 10396
rect 24652 10436 24692 12100
rect 24652 10387 24692 10396
rect 26380 10436 26420 12100
rect 28012 10856 28052 10865
rect 26380 10387 26420 10396
rect 27148 10772 27188 10781
rect 21964 9967 22004 9976
rect 22636 10352 22676 10361
rect 21004 9512 21044 9521
rect 20620 9008 20660 9017
rect 20620 8924 20660 8968
rect 20620 8873 20660 8884
rect 21004 8756 21044 9472
rect 21004 8707 21044 8716
rect 21196 9512 21236 9521
rect 20524 8623 20564 8632
rect 21196 8672 21236 9472
rect 21196 8623 21236 8632
rect 21580 8840 21620 8849
rect 19660 8539 19700 8548
rect 19756 8504 19796 8513
rect 18808 8336 19176 8345
rect 18848 8296 18890 8336
rect 18930 8296 18972 8336
rect 19012 8296 19054 8336
rect 19094 8296 19136 8336
rect 18808 8287 19176 8296
rect 17260 7027 17300 7036
rect 18808 6824 19176 6833
rect 18848 6784 18890 6824
rect 18930 6784 18972 6824
rect 19012 6784 19054 6824
rect 19094 6784 19136 6824
rect 18808 6775 19176 6784
rect 17164 6103 17204 6112
rect 15820 5683 15860 5692
rect 14284 5599 14324 5608
rect 9196 5564 9236 5573
rect 8812 5179 8852 5188
rect 8908 5312 8948 5321
rect 8716 5144 8756 5153
rect 7948 4976 7988 4985
rect 6412 391 6452 400
rect 7564 4136 7604 4145
rect 6028 307 6068 316
rect 5740 223 5780 232
rect 7564 80 7604 4096
rect 7756 4052 7796 4061
rect 7756 80 7796 4012
rect 7948 80 7988 4936
rect 8140 4892 8180 4901
rect 8140 80 8180 4852
rect 8524 4220 8564 4229
rect 8332 3884 8372 3893
rect 8332 80 8372 3844
rect 8524 80 8564 4180
rect 8620 3968 8660 3977
rect 8620 3128 8660 3928
rect 8620 3079 8660 3088
rect 8716 80 8756 5104
rect 8812 4892 8852 4901
rect 8812 4640 8852 4852
rect 8812 4591 8852 4600
rect 8908 80 8948 5272
rect 9100 4976 9140 4985
rect 9004 4724 9044 4733
rect 9004 4388 9044 4684
rect 9004 4339 9044 4348
rect 9100 80 9140 4936
rect 9196 4724 9236 5524
rect 16972 5564 17012 5573
rect 9868 5480 9908 5489
rect 16876 5480 16916 5489
rect 9908 5440 10196 5480
rect 9868 5431 9908 5440
rect 9964 5312 10004 5321
rect 9484 5060 9524 5069
rect 9196 4675 9236 4684
rect 9292 4892 9332 4901
rect 9292 80 9332 4852
rect 9484 80 9524 5020
rect 9964 4976 10004 5272
rect 10156 5312 10196 5440
rect 10156 5263 10196 5272
rect 13036 5440 13268 5480
rect 13036 5144 13076 5440
rect 13036 5095 13076 5104
rect 11884 5060 11924 5069
rect 9964 4927 10004 4936
rect 11404 4976 11444 4985
rect 9676 4640 9716 4649
rect 9676 80 9716 4600
rect 10060 4304 10100 4313
rect 9868 3464 9908 3473
rect 9868 80 9908 3424
rect 10060 80 10100 4264
rect 10828 4220 10868 4229
rect 10444 4136 10484 4145
rect 10252 3296 10292 3305
rect 10252 80 10292 3256
rect 10444 80 10484 4096
rect 10636 3380 10676 3389
rect 10636 80 10676 3340
rect 10828 80 10868 4180
rect 11212 4136 11252 4145
rect 11020 4052 11060 4061
rect 11020 80 11060 4012
rect 11212 80 11252 4096
rect 11404 80 11444 4936
rect 11692 4892 11732 4901
rect 11692 4472 11732 4852
rect 11692 4423 11732 4432
rect 11788 3968 11828 3977
rect 11596 3716 11636 3725
rect 11596 80 11636 3676
rect 11788 3044 11828 3928
rect 11788 2995 11828 3004
rect 11884 1448 11924 5020
rect 11788 1408 11924 1448
rect 11980 4976 12020 4985
rect 11788 80 11828 1408
rect 11980 80 12020 4936
rect 13132 4724 13172 4733
rect 12748 4640 12788 4651
rect 12748 4556 12788 4600
rect 12748 4507 12788 4516
rect 12844 4640 12884 4649
rect 12844 4472 12884 4600
rect 13132 4589 13172 4684
rect 12844 4423 12884 4432
rect 13036 4388 13076 4397
rect 12940 4052 12980 4061
rect 12748 3968 12788 3977
rect 12748 3212 12788 3928
rect 12940 3917 12980 4012
rect 12748 3163 12788 3172
rect 12940 3212 12980 3221
rect 12364 1448 12404 1457
rect 12172 860 12212 869
rect 12172 80 12212 820
rect 12364 80 12404 1408
rect 12556 1364 12596 1373
rect 12556 80 12596 1324
rect 12748 1028 12788 1037
rect 12748 80 12788 988
rect 12940 80 12980 3172
rect 13036 2540 13076 4348
rect 13132 4220 13172 4229
rect 13132 3296 13172 4180
rect 13132 3247 13172 3256
rect 13036 2491 13076 2500
rect 13228 1868 13268 5440
rect 13420 5396 13460 5405
rect 13420 4976 13460 5356
rect 16204 5312 16244 5321
rect 16204 5177 16244 5272
rect 16492 5228 16532 5237
rect 13420 4927 13460 4936
rect 13228 1819 13268 1828
rect 13324 4724 13364 4733
rect 13324 1532 13364 4684
rect 16204 4724 16244 4733
rect 14476 4640 14516 4649
rect 13420 4472 13460 4481
rect 13420 4337 13460 4432
rect 14476 4388 14516 4600
rect 14476 4339 14516 4348
rect 16012 4472 16052 4481
rect 14284 4304 14324 4313
rect 14092 4220 14132 4229
rect 13420 4136 13460 4145
rect 13420 4001 13460 4096
rect 13804 3884 13844 3893
rect 13516 3632 13556 3641
rect 13516 2960 13556 3592
rect 13516 2911 13556 2920
rect 13708 3632 13748 3641
rect 13132 1492 13364 1532
rect 13420 2708 13460 2717
rect 13132 80 13172 1492
rect 13420 1448 13460 2668
rect 13324 1408 13460 1448
rect 13324 80 13364 1408
rect 13516 440 13556 449
rect 13516 80 13556 400
rect 13708 80 13748 3592
rect 13804 2036 13844 3844
rect 13996 3464 14036 3473
rect 13804 1987 13844 1996
rect 13900 3380 13940 3389
rect 13900 80 13940 3340
rect 13996 3329 14036 3424
rect 14092 80 14132 4180
rect 14188 3464 14228 3473
rect 14188 440 14228 3424
rect 14284 2204 14324 4264
rect 15820 4220 15860 4229
rect 14380 4136 14420 4145
rect 14380 3716 14420 4096
rect 14380 3667 14420 3676
rect 14860 3716 14900 3725
rect 14572 3464 14612 3473
rect 14284 2155 14324 2164
rect 14380 3296 14420 3305
rect 14380 1532 14420 3256
rect 14572 3296 14612 3424
rect 14572 3247 14612 3256
rect 14476 3128 14516 3137
rect 14476 2708 14516 3088
rect 14476 2659 14516 2668
rect 14572 2960 14612 2969
rect 14380 1483 14420 1492
rect 14572 440 14612 2920
rect 14188 400 14324 440
rect 14284 80 14324 400
rect 14476 400 14612 440
rect 14668 524 14708 533
rect 14476 80 14516 400
rect 14668 80 14708 484
rect 14860 80 14900 3676
rect 15820 3716 15860 4180
rect 15916 3968 15956 3977
rect 15916 3833 15956 3928
rect 15820 3667 15860 3676
rect 16012 2372 16052 4432
rect 16012 2323 16052 2332
rect 16108 4136 16148 4145
rect 16012 1448 16052 1457
rect 15628 1196 15668 1205
rect 15244 944 15284 953
rect 15052 104 15092 113
rect 2860 55 2900 64
rect 7544 0 7624 80
rect 7736 0 7816 80
rect 7928 0 8008 80
rect 8120 0 8200 80
rect 8312 0 8392 80
rect 8504 0 8584 80
rect 8696 0 8776 80
rect 8888 0 8968 80
rect 9080 0 9160 80
rect 9272 0 9352 80
rect 9464 0 9544 80
rect 9656 0 9736 80
rect 9848 0 9928 80
rect 10040 0 10120 80
rect 10232 0 10312 80
rect 10424 0 10504 80
rect 10616 0 10696 80
rect 10808 0 10888 80
rect 11000 0 11080 80
rect 11192 0 11272 80
rect 11384 0 11464 80
rect 11576 0 11656 80
rect 11768 0 11848 80
rect 11960 0 12040 80
rect 12152 0 12232 80
rect 12344 0 12424 80
rect 12536 0 12616 80
rect 12728 0 12808 80
rect 12920 0 13000 80
rect 13112 0 13192 80
rect 13304 0 13384 80
rect 13496 0 13576 80
rect 13688 0 13768 80
rect 13880 0 13960 80
rect 14072 0 14152 80
rect 14264 0 14344 80
rect 14456 0 14536 80
rect 14648 0 14728 80
rect 14840 0 14920 80
rect 15032 64 15052 80
rect 15244 80 15284 904
rect 15436 356 15476 365
rect 15436 80 15476 316
rect 15628 80 15668 1156
rect 15820 524 15860 533
rect 15820 80 15860 484
rect 16012 80 16052 1408
rect 16108 776 16148 4096
rect 16204 2876 16244 4684
rect 16204 2827 16244 2836
rect 16300 3968 16340 3977
rect 16300 2456 16340 3928
rect 16300 2407 16340 2416
rect 16108 727 16148 736
rect 16396 1112 16436 1121
rect 16204 692 16244 701
rect 16204 80 16244 652
rect 16396 80 16436 1072
rect 16492 440 16532 5188
rect 16588 4472 16628 4481
rect 16588 1952 16628 4432
rect 16684 4136 16724 4145
rect 16684 3632 16724 4096
rect 16780 3884 16820 3893
rect 16780 3749 16820 3844
rect 16684 3583 16724 3592
rect 16876 2900 16916 5440
rect 16972 4388 17012 5524
rect 17836 5312 17876 5321
rect 17068 4976 17108 4985
rect 17260 4976 17300 4985
rect 17068 4841 17108 4936
rect 17164 4936 17260 4976
rect 17164 4724 17204 4936
rect 17260 4927 17300 4936
rect 17164 4675 17204 4684
rect 16972 4348 17108 4388
rect 16876 2860 17012 2900
rect 16588 1903 16628 1912
rect 16780 776 16820 785
rect 16492 400 16628 440
rect 16588 80 16628 400
rect 16780 80 16820 736
rect 16972 80 17012 2860
rect 17068 1952 17108 4348
rect 17356 4136 17396 4145
rect 17164 3884 17204 3893
rect 17164 3632 17204 3844
rect 17164 3583 17204 3592
rect 17260 3548 17300 3557
rect 17260 3044 17300 3508
rect 17356 3212 17396 4096
rect 17356 3163 17396 3172
rect 17644 4136 17684 4145
rect 17260 3004 17492 3044
rect 17164 2960 17204 2969
rect 17204 2920 17396 2960
rect 17164 2911 17204 2920
rect 17356 2120 17396 2920
rect 17452 2900 17492 3004
rect 17452 2860 17588 2900
rect 17356 2071 17396 2080
rect 17452 2288 17492 2297
rect 17068 1903 17108 1912
rect 17452 1448 17492 2248
rect 17548 1952 17588 2860
rect 17548 1903 17588 1912
rect 17356 1408 17492 1448
rect 17548 1700 17588 1709
rect 17164 608 17204 617
rect 17164 80 17204 568
rect 17356 80 17396 1408
rect 17548 80 17588 1660
rect 17644 1448 17684 4096
rect 17740 3296 17780 3305
rect 17740 2960 17780 3256
rect 17740 2911 17780 2920
rect 17644 1399 17684 1408
rect 17740 2456 17780 2465
rect 17740 80 17780 2416
rect 17836 2036 17876 5272
rect 18124 5312 18164 5321
rect 17836 1987 17876 1996
rect 17932 4976 17972 4985
rect 17932 1868 17972 4936
rect 17836 1828 17972 1868
rect 18028 4136 18068 4145
rect 17836 860 17876 1828
rect 17836 811 17876 820
rect 17932 1700 17972 1709
rect 17932 80 17972 1660
rect 18028 1364 18068 4096
rect 18124 2624 18164 5272
rect 18808 5312 19176 5321
rect 18848 5272 18890 5312
rect 18930 5272 18972 5312
rect 19012 5272 19054 5312
rect 19094 5272 19136 5312
rect 18808 5263 19176 5272
rect 18220 5228 18260 5237
rect 18220 4976 18260 5188
rect 18220 4927 18260 4936
rect 18124 2575 18164 2584
rect 18220 4136 18260 4145
rect 18028 1315 18068 1324
rect 18124 2456 18164 2465
rect 18124 80 18164 2416
rect 18220 1028 18260 4096
rect 18700 4136 18740 4145
rect 18604 4052 18644 4061
rect 18508 3968 18548 3977
rect 18316 3884 18356 3893
rect 18316 3464 18356 3844
rect 18508 3884 18548 3928
rect 18508 3833 18548 3844
rect 18316 3415 18356 3424
rect 18508 3044 18548 3053
rect 18508 2708 18548 3004
rect 18508 2659 18548 2668
rect 18412 2624 18452 2633
rect 18412 2288 18452 2584
rect 18412 2239 18452 2248
rect 18508 2456 18548 2465
rect 18316 1952 18356 2047
rect 18316 1903 18356 1912
rect 18220 979 18260 988
rect 18316 1700 18356 1709
rect 18316 80 18356 1660
rect 18508 80 18548 2416
rect 18604 2204 18644 4012
rect 18700 2708 18740 4096
rect 19564 4136 19604 4145
rect 19372 4052 19412 4061
rect 18808 3800 19176 3809
rect 18848 3760 18890 3800
rect 18930 3760 18972 3800
rect 19012 3760 19054 3800
rect 19094 3760 19136 3800
rect 18808 3751 19176 3760
rect 18796 3632 18836 3641
rect 18796 3044 18836 3592
rect 18796 2995 18836 3004
rect 18700 2659 18740 2668
rect 18604 2155 18644 2164
rect 18700 2456 18740 2465
rect 18604 1700 18644 1709
rect 18604 1196 18644 1660
rect 18700 1280 18740 2416
rect 19276 2456 19316 2465
rect 18808 2288 19176 2297
rect 18848 2248 18890 2288
rect 18930 2248 18972 2288
rect 19012 2248 19054 2288
rect 19094 2248 19136 2288
rect 18808 2239 19176 2248
rect 19084 1700 19124 1709
rect 18700 1240 18932 1280
rect 18604 1156 18740 1196
rect 18700 80 18740 1156
rect 18892 80 18932 1240
rect 19084 80 19124 1660
rect 19276 80 19316 2416
rect 19372 1952 19412 4012
rect 19372 1903 19412 1912
rect 19564 1868 19604 4096
rect 19660 3968 19700 3977
rect 19660 3800 19700 3928
rect 19660 3751 19700 3760
rect 19756 3380 19796 8464
rect 20048 7580 20416 7589
rect 20088 7540 20130 7580
rect 20170 7540 20212 7580
rect 20252 7540 20294 7580
rect 20334 7540 20376 7580
rect 20048 7531 20416 7540
rect 21580 7076 21620 8800
rect 22636 8840 22676 10312
rect 25900 10268 25940 10277
rect 23212 10184 23252 10193
rect 22924 9428 22964 9439
rect 22924 9344 22964 9388
rect 22924 9295 22964 9304
rect 23020 9428 23060 9437
rect 22636 8791 22676 8800
rect 22924 9176 22964 9185
rect 23020 9176 23060 9388
rect 23020 9136 23156 9176
rect 21580 7027 21620 7036
rect 22924 6572 22964 9136
rect 23116 8756 23156 9136
rect 23116 8707 23156 8716
rect 23212 6656 23252 10144
rect 24268 10100 24308 10109
rect 24076 9848 24116 9857
rect 24076 8672 24116 9808
rect 24076 8623 24116 8632
rect 24268 8672 24308 10060
rect 24364 9764 24404 9773
rect 24364 9512 24404 9724
rect 24364 9463 24404 9472
rect 24556 9764 24596 9773
rect 24268 8623 24308 8632
rect 24460 9428 24500 9437
rect 24460 8588 24500 9388
rect 24556 8672 24596 9724
rect 25804 9092 25844 9101
rect 25228 9008 25268 9017
rect 24556 8623 24596 8632
rect 25132 8840 25172 8849
rect 25132 8672 25172 8800
rect 25228 8840 25268 8968
rect 25228 8791 25268 8800
rect 25132 8623 25172 8632
rect 25804 8672 25844 9052
rect 25900 8672 25940 10228
rect 26380 10184 26420 10193
rect 26092 8672 26132 8681
rect 25900 8632 26092 8672
rect 25804 8623 25844 8632
rect 26092 8623 26132 8632
rect 24460 8539 24500 8548
rect 23212 6607 23252 6616
rect 22924 6523 22964 6532
rect 20048 6068 20416 6077
rect 20088 6028 20130 6068
rect 20170 6028 20212 6068
rect 20252 6028 20294 6068
rect 20334 6028 20376 6068
rect 20048 6019 20416 6028
rect 22348 5480 22388 5489
rect 20140 5396 20180 5405
rect 20140 5261 20180 5356
rect 22348 4976 22388 5440
rect 22348 4927 22388 4936
rect 24172 5396 24212 5405
rect 20048 4556 20416 4565
rect 20088 4516 20130 4556
rect 20170 4516 20212 4556
rect 20252 4516 20294 4556
rect 20334 4516 20376 4556
rect 20048 4507 20416 4516
rect 21292 4472 21332 4481
rect 21100 4388 21140 4397
rect 20812 4136 20852 4145
rect 19756 3331 19796 3340
rect 19852 4052 19892 4061
rect 19756 3128 19796 3137
rect 19660 2876 19700 2885
rect 19660 2624 19700 2836
rect 19660 2575 19700 2584
rect 19564 1819 19604 1828
rect 19660 2456 19700 2465
rect 19468 1700 19508 1709
rect 19468 80 19508 1660
rect 19660 80 19700 2416
rect 19756 1952 19796 3088
rect 19756 1903 19796 1912
rect 19852 1952 19892 4012
rect 20620 4052 20660 4061
rect 19948 3968 19988 3977
rect 19948 2876 19988 3928
rect 20140 3968 20180 3977
rect 20044 3884 20084 3893
rect 20044 3749 20084 3844
rect 20140 3833 20180 3928
rect 20140 3548 20180 3557
rect 20140 3212 20180 3508
rect 20140 3163 20180 3172
rect 20524 3464 20564 3473
rect 20048 3044 20416 3053
rect 20088 3004 20130 3044
rect 20170 3004 20212 3044
rect 20252 3004 20294 3044
rect 20334 3004 20376 3044
rect 20048 2995 20416 3004
rect 19948 2827 19988 2836
rect 20140 2624 20180 2633
rect 20140 2489 20180 2584
rect 20140 2288 20180 2297
rect 20140 2153 20180 2248
rect 19852 1903 19892 1912
rect 20044 2036 20084 2045
rect 20044 1952 20084 1996
rect 20044 1901 20084 1912
rect 19756 1784 19796 1793
rect 19756 440 19796 1744
rect 19756 391 19796 400
rect 19852 1784 19892 1793
rect 19852 80 19892 1744
rect 20428 1784 20468 1879
rect 20524 1868 20564 3424
rect 20620 1952 20660 4012
rect 20716 2960 20756 2969
rect 20716 2036 20756 2920
rect 20716 1987 20756 1996
rect 20620 1903 20660 1912
rect 20812 1868 20852 4096
rect 21004 3968 21044 3977
rect 20524 1819 20564 1828
rect 20716 1828 20852 1868
rect 20908 3884 20948 3893
rect 20908 1868 20948 3844
rect 21004 1952 21044 3928
rect 21100 2204 21140 4348
rect 21100 2155 21140 2164
rect 21196 3632 21236 3641
rect 21196 2204 21236 3592
rect 21292 2708 21332 4432
rect 23212 4388 23252 4397
rect 22444 4220 22484 4229
rect 21868 4136 21908 4145
rect 21772 4052 21812 4061
rect 21388 3968 21428 3977
rect 21388 3632 21428 3928
rect 21388 3583 21428 3592
rect 21484 3716 21524 3725
rect 21292 2659 21332 2668
rect 21388 3464 21428 3473
rect 21388 2624 21428 3424
rect 21388 2575 21428 2584
rect 21196 2155 21236 2164
rect 21292 2540 21332 2549
rect 21004 1903 21044 1912
rect 21196 2036 21236 2045
rect 20428 1735 20468 1744
rect 20620 1784 20660 1793
rect 19948 1700 19988 1709
rect 19948 860 19988 1660
rect 20524 1700 20564 1709
rect 20048 1532 20416 1541
rect 20088 1492 20130 1532
rect 20170 1492 20212 1532
rect 20252 1492 20294 1532
rect 20334 1492 20376 1532
rect 20048 1483 20416 1492
rect 20236 860 20276 869
rect 20524 860 20564 1660
rect 19948 820 20084 860
rect 20044 80 20084 820
rect 20236 80 20276 820
rect 20428 820 20564 860
rect 20428 80 20468 820
rect 20620 80 20660 1744
rect 20716 1196 20756 1828
rect 20908 1819 20948 1828
rect 20716 1147 20756 1156
rect 20812 1700 20852 1709
rect 21100 1700 21140 1709
rect 20812 80 20852 1660
rect 21004 1660 21100 1700
rect 21004 80 21044 1660
rect 21100 1651 21140 1660
rect 21196 80 21236 1996
rect 21292 356 21332 2500
rect 21292 307 21332 316
rect 21388 2456 21428 2465
rect 21388 80 21428 2416
rect 21484 2372 21524 3676
rect 21676 3296 21716 3305
rect 21580 3128 21620 3137
rect 21580 2993 21620 3088
rect 21676 2624 21716 3256
rect 21772 2624 21812 4012
rect 21868 2792 21908 4096
rect 22348 4136 22388 4145
rect 22252 3464 22292 3473
rect 21868 2743 21908 2752
rect 21964 3212 22004 3221
rect 21964 2624 22004 3172
rect 21772 2584 21908 2624
rect 21676 2575 21716 2584
rect 21484 2323 21524 2332
rect 21772 2456 21812 2465
rect 21484 1952 21524 1961
rect 21484 944 21524 1912
rect 21676 1868 21716 1877
rect 21484 895 21524 904
rect 21580 1784 21620 1793
rect 21580 80 21620 1744
rect 21676 1448 21716 1828
rect 21676 1399 21716 1408
rect 21772 80 21812 2416
rect 21868 1112 21908 2584
rect 21964 2575 22004 2584
rect 22060 3212 22100 3221
rect 22060 2120 22100 3172
rect 22156 2876 22196 2885
rect 22156 2741 22196 2836
rect 22060 2071 22100 2080
rect 22156 2456 22196 2465
rect 21964 2036 22004 2045
rect 21964 1901 22004 1996
rect 21868 1063 21908 1072
rect 21964 1700 22004 1709
rect 21964 80 22004 1660
rect 22156 80 22196 2416
rect 22252 608 22292 3424
rect 22348 2876 22388 4096
rect 22348 2827 22388 2836
rect 22348 2708 22388 2717
rect 22348 2204 22388 2668
rect 22444 2624 22484 4180
rect 22636 4220 22676 4315
rect 22636 4171 22676 4180
rect 22924 4136 22964 4145
rect 22636 4052 22676 4061
rect 22540 3968 22580 3977
rect 22540 3296 22580 3928
rect 22540 3247 22580 3256
rect 22540 2876 22580 2885
rect 22540 2624 22580 2836
rect 22636 2792 22676 4012
rect 22732 3884 22772 3893
rect 22732 3380 22772 3844
rect 22732 3331 22772 3340
rect 22828 3800 22868 3809
rect 22636 2743 22676 2752
rect 22732 3128 22772 3137
rect 22540 2584 22676 2624
rect 22444 2575 22484 2584
rect 22540 2456 22580 2465
rect 22348 2164 22484 2204
rect 22252 559 22292 568
rect 22348 2036 22388 2045
rect 22348 80 22388 1996
rect 22444 692 22484 2164
rect 22444 643 22484 652
rect 22540 80 22580 2416
rect 22636 524 22676 2584
rect 22732 2036 22772 3088
rect 22732 1987 22772 1996
rect 22828 1868 22868 3760
rect 22924 2792 22964 4096
rect 22924 2743 22964 2752
rect 23020 2708 23060 2717
rect 23020 2573 23060 2668
rect 23212 2624 23252 4348
rect 23500 4304 23540 4313
rect 23500 3716 23540 4264
rect 23500 3667 23540 3676
rect 23788 4136 23828 4145
rect 23212 2575 23252 2584
rect 22828 1819 22868 1828
rect 22924 2456 22964 2465
rect 22636 475 22676 484
rect 22732 1784 22772 1793
rect 22732 80 22772 1744
rect 22828 1700 22868 1709
rect 22828 776 22868 1660
rect 22828 727 22868 736
rect 22924 80 22964 2416
rect 23308 2456 23348 2465
rect 23020 2372 23060 2381
rect 23020 2237 23060 2332
rect 23116 2204 23156 2215
rect 23116 2120 23156 2164
rect 23116 2071 23156 2080
rect 23020 2036 23060 2045
rect 23020 1901 23060 1996
rect 23116 1700 23156 1709
rect 23116 80 23156 1660
rect 23308 80 23348 2416
rect 23692 2456 23732 2465
rect 23500 1616 23540 1625
rect 23500 80 23540 1576
rect 23692 80 23732 2416
rect 23788 1112 23828 4096
rect 23884 3632 23924 3641
rect 23884 2036 23924 3592
rect 23980 2456 24020 2465
rect 23980 2204 24020 2416
rect 23980 2155 24020 2164
rect 24076 2456 24116 2465
rect 23884 1996 24020 2036
rect 23980 1868 24020 1996
rect 23980 1819 24020 1828
rect 23788 1063 23828 1072
rect 23884 1784 23924 1793
rect 23884 80 23924 1744
rect 24076 80 24116 2416
rect 24172 2120 24212 5356
rect 24940 5228 24980 5237
rect 24556 4556 24596 4565
rect 24172 2071 24212 2080
rect 24268 4136 24308 4145
rect 24172 1952 24212 1961
rect 24172 1868 24212 1912
rect 24268 1952 24308 4096
rect 24364 2624 24404 2633
rect 24364 2288 24404 2584
rect 24364 2239 24404 2248
rect 24460 2456 24500 2465
rect 24268 1903 24308 1912
rect 24172 1817 24212 1828
rect 24268 1616 24308 1625
rect 24268 80 24308 1576
rect 24460 80 24500 2416
rect 24556 1952 24596 4516
rect 24748 3128 24788 3137
rect 24748 2624 24788 3088
rect 24748 2575 24788 2584
rect 24556 1903 24596 1912
rect 24844 2456 24884 2465
rect 24652 1616 24692 1625
rect 24652 80 24692 1576
rect 24844 80 24884 2416
rect 24940 1952 24980 5188
rect 26380 5144 26420 10144
rect 26380 5095 26420 5104
rect 26668 10184 26708 10193
rect 25132 4724 25172 4733
rect 25132 2624 25172 4684
rect 25132 2575 25172 2584
rect 25516 4640 25556 4649
rect 25516 2624 25556 4600
rect 26572 4304 26612 4313
rect 26188 4136 26228 4145
rect 26092 3884 26132 3893
rect 25900 3296 25940 3305
rect 25516 2575 25556 2584
rect 25708 3212 25748 3221
rect 24940 1903 24980 1912
rect 25228 2456 25268 2465
rect 25036 1784 25076 1793
rect 25036 80 25076 1744
rect 25228 80 25268 2416
rect 25612 2456 25652 2465
rect 25420 1616 25460 1625
rect 25420 80 25460 1576
rect 25612 80 25652 2416
rect 25708 1952 25748 3172
rect 25900 2624 25940 3256
rect 25900 2575 25940 2584
rect 25708 1903 25748 1912
rect 25996 2456 26036 2465
rect 25804 1616 25844 1625
rect 25804 80 25844 1576
rect 25996 80 26036 2416
rect 26092 1952 26132 3844
rect 26188 2204 26228 4096
rect 26476 3800 26516 3809
rect 26284 3716 26324 3725
rect 26284 2624 26324 3676
rect 26284 2575 26324 2584
rect 26380 2456 26420 2465
rect 26188 2164 26324 2204
rect 26092 1903 26132 1912
rect 26188 2036 26228 2045
rect 26188 80 26228 1996
rect 26284 188 26324 2164
rect 26284 139 26324 148
rect 26380 80 26420 2416
rect 26476 1952 26516 3760
rect 26572 2900 26612 4264
rect 26668 3632 26708 10144
rect 27148 8588 27188 10732
rect 28012 10268 28052 10816
rect 28108 10436 28148 12100
rect 28108 10387 28148 10396
rect 28684 10604 28724 10613
rect 28012 10219 28052 10228
rect 28396 10184 28436 10193
rect 28204 9932 28244 9941
rect 27148 8539 27188 8548
rect 27724 9512 27764 9521
rect 27724 6320 27764 9472
rect 27820 9008 27860 9017
rect 27820 8672 27860 8968
rect 27820 8623 27860 8632
rect 28108 8756 28148 8767
rect 28108 8672 28148 8716
rect 28108 8623 28148 8632
rect 28204 8504 28244 9892
rect 28204 8455 28244 8464
rect 27724 6280 28340 6320
rect 26668 3583 26708 3592
rect 27052 4304 27092 4313
rect 26860 3380 26900 3389
rect 26572 2860 26708 2900
rect 26668 2624 26708 2860
rect 26668 2575 26708 2584
rect 26476 1903 26516 1912
rect 26764 2456 26804 2465
rect 26572 1784 26612 1793
rect 26572 80 26612 1744
rect 26764 80 26804 2416
rect 26860 1952 26900 3340
rect 27052 2624 27092 4264
rect 27052 2575 27092 2584
rect 27244 4052 27284 4061
rect 26860 1903 26900 1912
rect 27148 2456 27188 2465
rect 26956 1616 26996 1625
rect 26956 80 26996 1576
rect 27148 80 27188 2416
rect 27244 2036 27284 4012
rect 27340 3968 27380 3977
rect 27340 2960 27380 3928
rect 27340 2911 27380 2920
rect 28012 3968 28052 3977
rect 27244 1987 27284 1996
rect 28012 1952 28052 3928
rect 28204 3968 28244 3977
rect 28204 2624 28244 3928
rect 28300 2900 28340 6280
rect 28396 3632 28436 10144
rect 28684 8168 28724 10564
rect 29836 10436 29876 12100
rect 29836 10387 29876 10396
rect 31564 10436 31604 12100
rect 31564 10387 31604 10396
rect 31660 10772 31700 10781
rect 30124 10184 30164 10193
rect 29260 9848 29300 9857
rect 28972 9092 29012 9101
rect 28780 8672 28820 8681
rect 28820 8632 28916 8672
rect 28780 8623 28820 8632
rect 28684 8119 28724 8128
rect 28684 8000 28724 8009
rect 28396 3583 28436 3592
rect 28588 4136 28628 4145
rect 28300 2860 28532 2900
rect 28204 2575 28244 2584
rect 28012 1903 28052 1912
rect 27340 1616 27380 1625
rect 27340 80 27380 1576
rect 28108 440 28148 449
rect 27916 356 27956 365
rect 27724 188 27764 197
rect 27532 104 27572 113
rect 15092 64 15112 80
rect 15032 0 15112 64
rect 15224 0 15304 80
rect 15416 0 15496 80
rect 15608 0 15688 80
rect 15800 0 15880 80
rect 15992 0 16072 80
rect 16184 0 16264 80
rect 16376 0 16456 80
rect 16568 0 16648 80
rect 16760 0 16840 80
rect 16952 0 17032 80
rect 17144 0 17224 80
rect 17336 0 17416 80
rect 17528 0 17608 80
rect 17720 0 17800 80
rect 17912 0 17992 80
rect 18104 0 18184 80
rect 18296 0 18376 80
rect 18488 0 18568 80
rect 18680 0 18760 80
rect 18872 0 18952 80
rect 19064 0 19144 80
rect 19256 0 19336 80
rect 19448 0 19528 80
rect 19640 0 19720 80
rect 19832 0 19912 80
rect 20024 0 20104 80
rect 20216 0 20296 80
rect 20408 0 20488 80
rect 20600 0 20680 80
rect 20792 0 20872 80
rect 20984 0 21064 80
rect 21176 0 21256 80
rect 21368 0 21448 80
rect 21560 0 21640 80
rect 21752 0 21832 80
rect 21944 0 22024 80
rect 22136 0 22216 80
rect 22328 0 22408 80
rect 22520 0 22600 80
rect 22712 0 22792 80
rect 22904 0 22984 80
rect 23096 0 23176 80
rect 23288 0 23368 80
rect 23480 0 23560 80
rect 23672 0 23752 80
rect 23864 0 23944 80
rect 24056 0 24136 80
rect 24248 0 24328 80
rect 24440 0 24520 80
rect 24632 0 24712 80
rect 24824 0 24904 80
rect 25016 0 25096 80
rect 25208 0 25288 80
rect 25400 0 25480 80
rect 25592 0 25672 80
rect 25784 0 25864 80
rect 25976 0 26056 80
rect 26168 0 26248 80
rect 26360 0 26440 80
rect 26552 0 26632 80
rect 26744 0 26824 80
rect 26936 0 27016 80
rect 27128 0 27208 80
rect 27320 0 27400 80
rect 27512 64 27532 80
rect 27724 80 27764 148
rect 27916 80 27956 316
rect 28108 80 28148 400
rect 28300 272 28340 281
rect 28300 80 28340 232
rect 28492 80 28532 2860
rect 28588 524 28628 4096
rect 28588 475 28628 484
rect 28684 80 28724 7960
rect 28780 3968 28820 3977
rect 28780 1952 28820 3928
rect 28780 1903 28820 1912
rect 28876 80 28916 8632
rect 28972 2900 29012 9052
rect 29068 8672 29108 8681
rect 29068 8537 29108 8632
rect 28972 2860 29108 2900
rect 29068 80 29108 2860
rect 29260 80 29300 9808
rect 29452 9764 29492 9773
rect 29452 80 29492 9724
rect 29644 9008 29684 9017
rect 29644 80 29684 8968
rect 29836 6488 29876 6497
rect 29836 80 29876 6448
rect 30028 4976 30068 4985
rect 29932 4136 29972 4145
rect 29932 3044 29972 4096
rect 29932 2995 29972 3004
rect 30028 80 30068 4936
rect 30124 3632 30164 10144
rect 30220 9428 30260 9437
rect 30220 9293 30260 9388
rect 31660 9428 31700 10732
rect 33292 10436 33332 12100
rect 33292 10387 33332 10396
rect 35020 10436 35060 12100
rect 36364 10856 36404 10865
rect 35168 10604 35536 10613
rect 35208 10564 35250 10604
rect 35290 10564 35332 10604
rect 35372 10564 35414 10604
rect 35454 10564 35496 10604
rect 35168 10555 35536 10564
rect 35020 10387 35060 10396
rect 36364 10436 36404 10816
rect 36364 10387 36404 10396
rect 36748 10436 36788 12100
rect 36748 10387 36788 10396
rect 36940 11192 36980 11201
rect 31660 9379 31700 9388
rect 31852 10184 31892 10193
rect 30796 9260 30836 9269
rect 30220 9008 30260 9017
rect 30220 8873 30260 8968
rect 30796 8924 30836 9220
rect 30796 8875 30836 8884
rect 31372 4892 31412 4901
rect 30124 3583 30164 3592
rect 30988 4220 31028 4229
rect 30412 3464 30452 3473
rect 30316 3380 30356 3389
rect 30316 440 30356 3340
rect 30220 400 30356 440
rect 30220 80 30260 400
rect 30412 80 30452 3424
rect 30604 3464 30644 3473
rect 30604 80 30644 3424
rect 30796 3380 30836 3389
rect 30796 80 30836 3340
rect 30988 80 31028 4180
rect 31180 4052 31220 4061
rect 31180 80 31220 4012
rect 31372 80 31412 4852
rect 31564 3884 31604 3893
rect 31564 1952 31604 3844
rect 31852 3632 31892 10144
rect 32908 10184 32948 10193
rect 32524 10100 32564 10109
rect 31852 3583 31892 3592
rect 32332 4724 32372 4733
rect 32332 3464 32372 4684
rect 32524 4304 32564 10060
rect 32524 4255 32564 4264
rect 32908 4304 32948 10144
rect 35596 10100 35636 10109
rect 33928 9848 34296 9857
rect 33968 9808 34010 9848
rect 34050 9808 34092 9848
rect 34132 9808 34174 9848
rect 34214 9808 34256 9848
rect 33928 9799 34296 9808
rect 35168 9092 35536 9101
rect 35208 9052 35250 9092
rect 35290 9052 35332 9092
rect 35372 9052 35414 9092
rect 35454 9052 35496 9092
rect 35168 9043 35536 9052
rect 33484 8672 33524 8681
rect 32908 4255 32948 4264
rect 33196 4640 33236 4649
rect 32332 3415 32372 3424
rect 33004 4136 33044 4145
rect 31564 1903 31604 1912
rect 33004 1532 33044 4096
rect 33196 2624 33236 4600
rect 33484 4220 33524 8632
rect 33928 8336 34296 8345
rect 33968 8296 34010 8336
rect 34050 8296 34092 8336
rect 34132 8296 34174 8336
rect 34214 8296 34256 8336
rect 33928 8287 34296 8296
rect 35168 7580 35536 7589
rect 35208 7540 35250 7580
rect 35290 7540 35332 7580
rect 35372 7540 35414 7580
rect 35454 7540 35496 7580
rect 35168 7531 35536 7540
rect 33928 6824 34296 6833
rect 33968 6784 34010 6824
rect 34050 6784 34092 6824
rect 34132 6784 34174 6824
rect 34214 6784 34256 6824
rect 33928 6775 34296 6784
rect 35168 6068 35536 6077
rect 35208 6028 35250 6068
rect 35290 6028 35332 6068
rect 35372 6028 35414 6068
rect 35454 6028 35496 6068
rect 35168 6019 35536 6028
rect 33928 5312 34296 5321
rect 33968 5272 34010 5312
rect 34050 5272 34092 5312
rect 34132 5272 34174 5312
rect 34214 5272 34256 5312
rect 33928 5263 34296 5272
rect 35596 5144 35636 10060
rect 36652 9680 36692 9689
rect 36652 8672 36692 9640
rect 36940 9680 36980 11152
rect 37804 10772 37844 10781
rect 37324 10520 37364 10529
rect 36940 9631 36980 9640
rect 37228 10016 37268 10025
rect 37228 9512 37268 9976
rect 37324 9680 37364 10480
rect 37804 10184 37844 10732
rect 37804 10135 37844 10144
rect 38764 10016 38804 10025
rect 37324 9631 37364 9640
rect 37804 9764 37844 9773
rect 37228 9463 37268 9472
rect 37612 9512 37652 9521
rect 37612 8924 37652 9472
rect 37612 8875 37652 8884
rect 37708 9428 37748 9437
rect 36652 8623 36692 8632
rect 37516 8840 37556 8849
rect 35596 5095 35636 5104
rect 35980 6236 36020 6245
rect 35168 4556 35536 4565
rect 35208 4516 35250 4556
rect 35290 4516 35332 4556
rect 35372 4516 35414 4556
rect 35454 4516 35496 4556
rect 35168 4507 35536 4516
rect 33484 4171 33524 4180
rect 35980 4136 36020 6196
rect 37516 4976 37556 8800
rect 37516 4927 37556 4936
rect 37708 4976 37748 9388
rect 37804 6488 37844 9724
rect 38764 9512 38804 9976
rect 38764 9463 38804 9472
rect 37804 6439 37844 6448
rect 37900 9344 37940 9353
rect 37708 4927 37748 4936
rect 35980 4087 36020 4096
rect 37612 4472 37652 4481
rect 37420 4052 37460 4061
rect 37460 4012 37556 4052
rect 37420 3984 37460 4012
rect 34540 3968 34580 3977
rect 33928 3800 34296 3809
rect 33968 3760 34010 3800
rect 34050 3760 34092 3800
rect 34132 3760 34174 3800
rect 34214 3760 34256 3800
rect 33928 3751 34296 3760
rect 34540 2708 34580 3928
rect 35168 3044 35536 3053
rect 35208 3004 35250 3044
rect 35290 3004 35332 3044
rect 35372 3004 35414 3044
rect 35454 3004 35496 3044
rect 35168 2995 35536 3004
rect 34540 2659 34580 2668
rect 33196 2575 33236 2584
rect 37420 2624 37460 2633
rect 37516 2624 37556 4012
rect 37460 2584 37556 2624
rect 37420 2556 37460 2584
rect 33928 2288 34296 2297
rect 33968 2248 34010 2288
rect 34050 2248 34092 2288
rect 34132 2248 34174 2288
rect 34214 2248 34256 2288
rect 33928 2239 34296 2248
rect 37612 1952 37652 4432
rect 37900 4136 37940 9304
rect 38668 9260 38708 9269
rect 38668 8840 38708 9220
rect 38668 8791 38708 8800
rect 39148 8672 39188 8681
rect 39148 8168 39188 8632
rect 39148 8119 39188 8128
rect 37900 4087 37940 4096
rect 37612 1903 37652 1912
rect 38380 2456 38420 2465
rect 37516 1784 37556 1793
rect 33004 1483 33044 1492
rect 35168 1532 35536 1541
rect 35208 1492 35250 1532
rect 35290 1492 35332 1532
rect 35372 1492 35414 1532
rect 35454 1492 35496 1532
rect 35168 1483 35536 1492
rect 37516 1112 37556 1744
rect 37516 1063 37556 1072
rect 38284 1700 38324 1709
rect 38284 776 38324 1660
rect 38380 1448 38420 2416
rect 38380 1399 38420 1408
rect 38284 727 38324 736
rect 27572 64 27592 80
rect 27512 0 27592 64
rect 27704 0 27784 80
rect 27896 0 27976 80
rect 28088 0 28168 80
rect 28280 0 28360 80
rect 28472 0 28552 80
rect 28664 0 28744 80
rect 28856 0 28936 80
rect 29048 0 29128 80
rect 29240 0 29320 80
rect 29432 0 29512 80
rect 29624 0 29704 80
rect 29816 0 29896 80
rect 30008 0 30088 80
rect 30200 0 30280 80
rect 30392 0 30472 80
rect 30584 0 30664 80
rect 30776 0 30856 80
rect 30968 0 31048 80
rect 31160 0 31240 80
rect 31352 0 31432 80
<< via3 >>
rect 364 8800 404 8840
rect 268 8716 308 8756
rect 172 8632 212 8672
rect 4928 10564 4968 10604
rect 5010 10564 5050 10604
rect 5092 10564 5132 10604
rect 5174 10564 5214 10604
rect 5256 10564 5296 10604
rect 3688 9808 3728 9848
rect 3770 9808 3810 9848
rect 3852 9808 3892 9848
rect 3934 9808 3974 9848
rect 4016 9808 4056 9848
rect 3688 8296 3728 8336
rect 3770 8296 3810 8336
rect 3852 8296 3892 8336
rect 3934 8296 3974 8336
rect 4016 8296 4056 8336
rect 3688 6784 3728 6824
rect 3770 6784 3810 6824
rect 3852 6784 3892 6824
rect 3934 6784 3974 6824
rect 4016 6784 4056 6824
rect 1420 1072 1460 1112
rect 4928 9052 4968 9092
rect 5010 9052 5050 9092
rect 5092 9052 5132 9092
rect 5174 9052 5214 9092
rect 5256 9052 5296 9092
rect 4928 7540 4968 7580
rect 5010 7540 5050 7580
rect 5092 7540 5132 7580
rect 5174 7540 5214 7580
rect 5256 7540 5296 7580
rect 4928 6028 4968 6068
rect 5010 6028 5050 6068
rect 5092 6028 5132 6068
rect 5174 6028 5214 6068
rect 5256 6028 5296 6068
rect 3688 5272 3728 5312
rect 3770 5272 3810 5312
rect 3852 5272 3892 5312
rect 3934 5272 3974 5312
rect 4016 5272 4056 5312
rect 4928 4516 4968 4556
rect 5010 4516 5050 4556
rect 5092 4516 5132 4556
rect 5174 4516 5214 4556
rect 5256 4516 5296 4556
rect 3688 3760 3728 3800
rect 3770 3760 3810 3800
rect 3852 3760 3892 3800
rect 3934 3760 3974 3800
rect 4016 3760 4056 3800
rect 4928 3004 4968 3044
rect 5010 3004 5050 3044
rect 5092 3004 5132 3044
rect 5174 3004 5214 3044
rect 5256 3004 5296 3044
rect 2668 148 2708 188
rect 3688 2248 3728 2288
rect 3770 2248 3810 2288
rect 3852 2248 3892 2288
rect 3934 2248 3974 2288
rect 4016 2248 4056 2288
rect 4928 1492 4968 1532
rect 5010 1492 5050 1532
rect 5092 1492 5132 1532
rect 5174 1492 5214 1532
rect 5256 1492 5296 1532
rect 12940 8884 12980 8924
rect 20048 10564 20088 10604
rect 20130 10564 20170 10604
rect 20212 10564 20252 10604
rect 20294 10564 20334 10604
rect 20376 10564 20416 10604
rect 18808 9808 18848 9848
rect 18890 9808 18930 9848
rect 18972 9808 19012 9848
rect 19054 9808 19094 9848
rect 19136 9808 19176 9848
rect 17740 8884 17780 8924
rect 20048 9052 20088 9092
rect 20130 9052 20170 9092
rect 20212 9052 20252 9092
rect 20294 9052 20334 9092
rect 20376 9052 20416 9092
rect 20620 8968 20660 9008
rect 18808 8296 18848 8336
rect 18890 8296 18930 8336
rect 18972 8296 19012 8336
rect 19054 8296 19094 8336
rect 19136 8296 19176 8336
rect 18808 6784 18848 6824
rect 18890 6784 18930 6824
rect 18972 6784 19012 6824
rect 19054 6784 19094 6824
rect 19136 6784 19176 6824
rect 6412 400 6452 440
rect 6028 316 6068 356
rect 5740 232 5780 272
rect 2860 64 2900 104
rect 10444 4096 10484 4136
rect 11980 4936 12020 4976
rect 13132 4684 13172 4724
rect 12748 4600 12788 4640
rect 12844 4432 12884 4472
rect 12940 4012 12980 4052
rect 12940 3172 12980 3212
rect 13420 5356 13460 5396
rect 16204 5272 16244 5312
rect 16204 4684 16244 4724
rect 14476 4600 14516 4640
rect 13420 4432 13460 4472
rect 13420 4096 13460 4136
rect 13420 2668 13460 2708
rect 13996 3424 14036 3464
rect 13804 1996 13844 2036
rect 15820 4180 15860 4220
rect 14572 3424 14612 3464
rect 14572 2920 14612 2960
rect 14668 484 14708 524
rect 15916 3928 15956 3968
rect 16012 1408 16052 1448
rect 16300 2416 16340 2456
rect 16780 3844 16820 3884
rect 17068 4936 17108 4976
rect 17164 3592 17204 3632
rect 17356 3172 17396 3212
rect 17068 1912 17108 1952
rect 18124 5272 18164 5312
rect 18808 5272 18848 5312
rect 18890 5272 18930 5312
rect 18972 5272 19012 5312
rect 19054 5272 19094 5312
rect 19136 5272 19176 5312
rect 18316 3844 18356 3884
rect 18508 3844 18548 3884
rect 18412 2584 18452 2624
rect 18316 1912 18356 1952
rect 19372 4012 19412 4052
rect 18808 3760 18848 3800
rect 18890 3760 18930 3800
rect 18972 3760 19012 3800
rect 19054 3760 19094 3800
rect 19136 3760 19176 3800
rect 18796 3592 18836 3632
rect 18700 2668 18740 2708
rect 18808 2248 18848 2288
rect 18890 2248 18930 2288
rect 18972 2248 19012 2288
rect 19054 2248 19094 2288
rect 19136 2248 19176 2288
rect 20048 7540 20088 7580
rect 20130 7540 20170 7580
rect 20212 7540 20252 7580
rect 20294 7540 20334 7580
rect 20376 7540 20416 7580
rect 22924 9388 22964 9428
rect 25132 8800 25172 8840
rect 20048 6028 20088 6068
rect 20130 6028 20170 6068
rect 20212 6028 20252 6068
rect 20294 6028 20334 6068
rect 20376 6028 20416 6068
rect 20140 5356 20180 5396
rect 20048 4516 20088 4556
rect 20130 4516 20170 4556
rect 20212 4516 20252 4556
rect 20294 4516 20334 4556
rect 20376 4516 20416 4556
rect 20140 3928 20180 3968
rect 20044 3844 20084 3884
rect 20140 3172 20180 3212
rect 20048 3004 20088 3044
rect 20130 3004 20170 3044
rect 20212 3004 20252 3044
rect 20294 3004 20334 3044
rect 20376 3004 20416 3044
rect 20140 2584 20180 2624
rect 20140 2248 20180 2288
rect 19852 1912 19892 1952
rect 20044 1996 20084 2036
rect 19756 1744 19796 1784
rect 20620 1912 20660 1952
rect 21196 2164 21236 2204
rect 21292 2500 21332 2540
rect 21196 1996 21236 2036
rect 20908 1828 20948 1868
rect 20428 1744 20468 1784
rect 20048 1492 20088 1532
rect 20130 1492 20170 1532
rect 20212 1492 20252 1532
rect 20294 1492 20334 1532
rect 20376 1492 20416 1532
rect 20236 820 20276 860
rect 21580 3088 21620 3128
rect 21868 2752 21908 2792
rect 21484 2332 21524 2372
rect 21484 1912 21524 1952
rect 22060 3172 22100 3212
rect 22156 2836 22196 2876
rect 21964 1996 22004 2036
rect 22348 2668 22388 2708
rect 22636 4180 22676 4220
rect 22636 2752 22676 2792
rect 22732 3088 22772 3128
rect 22348 1996 22388 2036
rect 22924 2752 22964 2792
rect 23020 2668 23060 2708
rect 22828 1660 22868 1700
rect 23020 2332 23060 2372
rect 23116 2164 23156 2204
rect 23020 1996 23060 2036
rect 23980 2416 24020 2456
rect 23788 1072 23828 1112
rect 24364 2248 24404 2288
rect 24268 1912 24308 1952
rect 24172 1828 24212 1868
rect 28108 8716 28148 8756
rect 27340 2920 27380 2960
rect 28108 400 28148 440
rect 27916 316 27956 356
rect 27724 148 27764 188
rect 27532 64 27572 104
rect 28300 232 28340 272
rect 28588 484 28628 524
rect 29068 8632 29108 8672
rect 30220 9388 30260 9428
rect 35168 10564 35208 10604
rect 35250 10564 35290 10604
rect 35332 10564 35372 10604
rect 35414 10564 35454 10604
rect 35496 10564 35536 10604
rect 30220 8968 30260 9008
rect 33928 9808 33968 9848
rect 34010 9808 34050 9848
rect 34092 9808 34132 9848
rect 34174 9808 34214 9848
rect 34256 9808 34296 9848
rect 35168 9052 35208 9092
rect 35250 9052 35290 9092
rect 35332 9052 35372 9092
rect 35414 9052 35454 9092
rect 35496 9052 35536 9092
rect 33928 8296 33968 8336
rect 34010 8296 34050 8336
rect 34092 8296 34132 8336
rect 34174 8296 34214 8336
rect 34256 8296 34296 8336
rect 35168 7540 35208 7580
rect 35250 7540 35290 7580
rect 35332 7540 35372 7580
rect 35414 7540 35454 7580
rect 35496 7540 35536 7580
rect 33928 6784 33968 6824
rect 34010 6784 34050 6824
rect 34092 6784 34132 6824
rect 34174 6784 34214 6824
rect 34256 6784 34296 6824
rect 35168 6028 35208 6068
rect 35250 6028 35290 6068
rect 35332 6028 35372 6068
rect 35414 6028 35454 6068
rect 35496 6028 35536 6068
rect 33928 5272 33968 5312
rect 34010 5272 34050 5312
rect 34092 5272 34132 5312
rect 34174 5272 34214 5312
rect 34256 5272 34296 5312
rect 35168 4516 35208 4556
rect 35250 4516 35290 4556
rect 35332 4516 35372 4556
rect 35414 4516 35454 4556
rect 35496 4516 35536 4556
rect 33928 3760 33968 3800
rect 34010 3760 34050 3800
rect 34092 3760 34132 3800
rect 34174 3760 34214 3800
rect 34256 3760 34296 3800
rect 35168 3004 35208 3044
rect 35250 3004 35290 3044
rect 35332 3004 35372 3044
rect 35414 3004 35454 3044
rect 35496 3004 35536 3044
rect 33928 2248 33968 2288
rect 34010 2248 34050 2288
rect 34092 2248 34132 2288
rect 34174 2248 34214 2288
rect 34256 2248 34296 2288
rect 35168 1492 35208 1532
rect 35250 1492 35290 1532
rect 35332 1492 35372 1532
rect 35414 1492 35454 1532
rect 35496 1492 35536 1532
<< metal4 >>
rect 4919 10564 4928 10604
rect 4968 10564 5010 10604
rect 5050 10564 5092 10604
rect 5132 10564 5174 10604
rect 5214 10564 5256 10604
rect 5296 10564 5305 10604
rect 20039 10564 20048 10604
rect 20088 10564 20130 10604
rect 20170 10564 20212 10604
rect 20252 10564 20294 10604
rect 20334 10564 20376 10604
rect 20416 10564 20425 10604
rect 35159 10564 35168 10604
rect 35208 10564 35250 10604
rect 35290 10564 35332 10604
rect 35372 10564 35414 10604
rect 35454 10564 35496 10604
rect 35536 10564 35545 10604
rect 3679 9808 3688 9848
rect 3728 9808 3770 9848
rect 3810 9808 3852 9848
rect 3892 9808 3934 9848
rect 3974 9808 4016 9848
rect 4056 9808 4065 9848
rect 18799 9808 18808 9848
rect 18848 9808 18890 9848
rect 18930 9808 18972 9848
rect 19012 9808 19054 9848
rect 19094 9808 19136 9848
rect 19176 9808 19185 9848
rect 33919 9808 33928 9848
rect 33968 9808 34010 9848
rect 34050 9808 34092 9848
rect 34132 9808 34174 9848
rect 34214 9808 34256 9848
rect 34296 9808 34305 9848
rect 22915 9388 22924 9428
rect 22964 9388 30220 9428
rect 30260 9388 30269 9428
rect 4919 9052 4928 9092
rect 4968 9052 5010 9092
rect 5050 9052 5092 9092
rect 5132 9052 5174 9092
rect 5214 9052 5256 9092
rect 5296 9052 5305 9092
rect 20039 9052 20048 9092
rect 20088 9052 20130 9092
rect 20170 9052 20212 9092
rect 20252 9052 20294 9092
rect 20334 9052 20376 9092
rect 20416 9052 20425 9092
rect 35159 9052 35168 9092
rect 35208 9052 35250 9092
rect 35290 9052 35332 9092
rect 35372 9052 35414 9092
rect 35454 9052 35496 9092
rect 35536 9052 35545 9092
rect 20611 8968 20620 9008
rect 20660 8968 30220 9008
rect 30260 8968 30269 9008
rect 12931 8884 12940 8924
rect 12980 8884 17740 8924
rect 17780 8884 17789 8924
rect 355 8800 364 8840
rect 404 8800 25132 8840
rect 25172 8800 25181 8840
rect 259 8716 268 8756
rect 308 8716 28108 8756
rect 28148 8716 28157 8756
rect 163 8632 172 8672
rect 212 8632 29068 8672
rect 29108 8632 29117 8672
rect 3679 8296 3688 8336
rect 3728 8296 3770 8336
rect 3810 8296 3852 8336
rect 3892 8296 3934 8336
rect 3974 8296 4016 8336
rect 4056 8296 4065 8336
rect 18799 8296 18808 8336
rect 18848 8296 18890 8336
rect 18930 8296 18972 8336
rect 19012 8296 19054 8336
rect 19094 8296 19136 8336
rect 19176 8296 19185 8336
rect 33919 8296 33928 8336
rect 33968 8296 34010 8336
rect 34050 8296 34092 8336
rect 34132 8296 34174 8336
rect 34214 8296 34256 8336
rect 34296 8296 34305 8336
rect 4919 7540 4928 7580
rect 4968 7540 5010 7580
rect 5050 7540 5092 7580
rect 5132 7540 5174 7580
rect 5214 7540 5256 7580
rect 5296 7540 5305 7580
rect 20039 7540 20048 7580
rect 20088 7540 20130 7580
rect 20170 7540 20212 7580
rect 20252 7540 20294 7580
rect 20334 7540 20376 7580
rect 20416 7540 20425 7580
rect 35159 7540 35168 7580
rect 35208 7540 35250 7580
rect 35290 7540 35332 7580
rect 35372 7540 35414 7580
rect 35454 7540 35496 7580
rect 35536 7540 35545 7580
rect 3679 6784 3688 6824
rect 3728 6784 3770 6824
rect 3810 6784 3852 6824
rect 3892 6784 3934 6824
rect 3974 6784 4016 6824
rect 4056 6784 4065 6824
rect 18799 6784 18808 6824
rect 18848 6784 18890 6824
rect 18930 6784 18972 6824
rect 19012 6784 19054 6824
rect 19094 6784 19136 6824
rect 19176 6784 19185 6824
rect 33919 6784 33928 6824
rect 33968 6784 34010 6824
rect 34050 6784 34092 6824
rect 34132 6784 34174 6824
rect 34214 6784 34256 6824
rect 34296 6784 34305 6824
rect 4919 6028 4928 6068
rect 4968 6028 5010 6068
rect 5050 6028 5092 6068
rect 5132 6028 5174 6068
rect 5214 6028 5256 6068
rect 5296 6028 5305 6068
rect 20039 6028 20048 6068
rect 20088 6028 20130 6068
rect 20170 6028 20212 6068
rect 20252 6028 20294 6068
rect 20334 6028 20376 6068
rect 20416 6028 20425 6068
rect 35159 6028 35168 6068
rect 35208 6028 35250 6068
rect 35290 6028 35332 6068
rect 35372 6028 35414 6068
rect 35454 6028 35496 6068
rect 35536 6028 35545 6068
rect 13411 5356 13420 5396
rect 13460 5356 20140 5396
rect 20180 5356 20189 5396
rect 3679 5272 3688 5312
rect 3728 5272 3770 5312
rect 3810 5272 3852 5312
rect 3892 5272 3934 5312
rect 3974 5272 4016 5312
rect 4056 5272 4065 5312
rect 16195 5272 16204 5312
rect 16244 5272 18124 5312
rect 18164 5272 18173 5312
rect 18799 5272 18808 5312
rect 18848 5272 18890 5312
rect 18930 5272 18972 5312
rect 19012 5272 19054 5312
rect 19094 5272 19136 5312
rect 19176 5272 19185 5312
rect 33919 5272 33928 5312
rect 33968 5272 34010 5312
rect 34050 5272 34092 5312
rect 34132 5272 34174 5312
rect 34214 5272 34256 5312
rect 34296 5272 34305 5312
rect 11971 4936 11980 4976
rect 12020 4936 17068 4976
rect 17108 4936 17117 4976
rect 13123 4684 13132 4724
rect 13172 4684 16204 4724
rect 16244 4684 16253 4724
rect 12739 4600 12748 4640
rect 12788 4600 14476 4640
rect 14516 4600 14525 4640
rect 4919 4516 4928 4556
rect 4968 4516 5010 4556
rect 5050 4516 5092 4556
rect 5132 4516 5174 4556
rect 5214 4516 5256 4556
rect 5296 4516 5305 4556
rect 20039 4516 20048 4556
rect 20088 4516 20130 4556
rect 20170 4516 20212 4556
rect 20252 4516 20294 4556
rect 20334 4516 20376 4556
rect 20416 4516 20425 4556
rect 35159 4516 35168 4556
rect 35208 4516 35250 4556
rect 35290 4516 35332 4556
rect 35372 4516 35414 4556
rect 35454 4516 35496 4556
rect 35536 4516 35545 4556
rect 12835 4432 12844 4472
rect 12884 4432 13420 4472
rect 13460 4432 13469 4472
rect 15811 4180 15820 4220
rect 15860 4180 22636 4220
rect 22676 4180 22685 4220
rect 10435 4096 10444 4136
rect 10484 4096 13420 4136
rect 13460 4096 13469 4136
rect 12931 4012 12940 4052
rect 12980 4012 19372 4052
rect 19412 4012 19421 4052
rect 15907 3928 15916 3968
rect 15956 3928 20140 3968
rect 20180 3928 20189 3968
rect 16771 3844 16780 3884
rect 16820 3844 18316 3884
rect 18356 3844 18365 3884
rect 18499 3844 18508 3884
rect 18548 3844 20044 3884
rect 20084 3844 20093 3884
rect 3679 3760 3688 3800
rect 3728 3760 3770 3800
rect 3810 3760 3852 3800
rect 3892 3760 3934 3800
rect 3974 3760 4016 3800
rect 4056 3760 4065 3800
rect 18799 3760 18808 3800
rect 18848 3760 18890 3800
rect 18930 3760 18972 3800
rect 19012 3760 19054 3800
rect 19094 3760 19136 3800
rect 19176 3760 19185 3800
rect 33919 3760 33928 3800
rect 33968 3760 34010 3800
rect 34050 3760 34092 3800
rect 34132 3760 34174 3800
rect 34214 3760 34256 3800
rect 34296 3760 34305 3800
rect 17155 3592 17164 3632
rect 17204 3592 18796 3632
rect 18836 3592 18845 3632
rect 13987 3424 13996 3464
rect 14036 3424 14572 3464
rect 14612 3424 14621 3464
rect 12931 3172 12940 3212
rect 12980 3172 17356 3212
rect 17396 3172 17405 3212
rect 20131 3172 20140 3212
rect 20180 3172 22060 3212
rect 22100 3172 22109 3212
rect 21571 3088 21580 3128
rect 21620 3088 22732 3128
rect 22772 3088 22781 3128
rect 4919 3004 4928 3044
rect 4968 3004 5010 3044
rect 5050 3004 5092 3044
rect 5132 3004 5174 3044
rect 5214 3004 5256 3044
rect 5296 3004 5305 3044
rect 20039 3004 20048 3044
rect 20088 3004 20130 3044
rect 20170 3004 20212 3044
rect 20252 3004 20294 3044
rect 20334 3004 20376 3044
rect 20416 3004 20425 3044
rect 35159 3004 35168 3044
rect 35208 3004 35250 3044
rect 35290 3004 35332 3044
rect 35372 3004 35414 3044
rect 35454 3004 35496 3044
rect 35536 3004 35545 3044
rect 14563 2920 14572 2960
rect 14612 2920 27340 2960
rect 27380 2920 27389 2960
rect 22147 2836 22156 2876
rect 22196 2836 22772 2876
rect 21859 2752 21868 2792
rect 21908 2752 21917 2792
rect 22627 2752 22636 2792
rect 22676 2752 22685 2792
rect 21868 2708 21908 2752
rect 13411 2668 13420 2708
rect 13460 2668 18700 2708
rect 18740 2668 18749 2708
rect 21868 2668 22348 2708
rect 22388 2668 22397 2708
rect 18403 2584 18412 2624
rect 18452 2584 20140 2624
rect 20180 2584 20189 2624
rect 22636 2540 22676 2752
rect 22732 2708 22772 2836
rect 22829 2752 22924 2792
rect 22964 2752 22973 2792
rect 22732 2668 23020 2708
rect 23060 2668 23069 2708
rect 21283 2500 21292 2540
rect 21332 2500 22676 2540
rect 16291 2416 16300 2456
rect 16340 2416 23980 2456
rect 24020 2416 24029 2456
rect 21475 2332 21484 2372
rect 21524 2332 23020 2372
rect 23060 2332 23069 2372
rect 3679 2248 3688 2288
rect 3728 2248 3770 2288
rect 3810 2248 3852 2288
rect 3892 2248 3934 2288
rect 3974 2248 4016 2288
rect 4056 2248 4065 2288
rect 18799 2248 18808 2288
rect 18848 2248 18890 2288
rect 18930 2248 18972 2288
rect 19012 2248 19054 2288
rect 19094 2248 19136 2288
rect 19176 2248 19185 2288
rect 20131 2248 20140 2288
rect 20180 2248 24364 2288
rect 24404 2248 24413 2288
rect 33919 2248 33928 2288
rect 33968 2248 34010 2288
rect 34050 2248 34092 2288
rect 34132 2248 34174 2288
rect 34214 2248 34256 2288
rect 34296 2248 34305 2288
rect 21187 2164 21196 2204
rect 21236 2164 23116 2204
rect 23156 2164 23165 2204
rect 13795 1996 13804 2036
rect 13844 1996 20044 2036
rect 20084 1996 20093 2036
rect 21187 1996 21196 2036
rect 21236 1996 21964 2036
rect 22004 1996 22013 2036
rect 22339 1996 22348 2036
rect 22388 1996 23020 2036
rect 23060 1996 23069 2036
rect 17059 1912 17068 1952
rect 17108 1912 18316 1952
rect 18356 1912 18365 1952
rect 19843 1912 19852 1952
rect 19892 1912 19901 1952
rect 20611 1912 20620 1952
rect 20660 1912 20669 1952
rect 21475 1912 21484 1952
rect 21524 1912 24268 1952
rect 24308 1912 24317 1952
rect 19852 1784 19892 1912
rect 19747 1744 19756 1784
rect 19796 1744 19892 1784
rect 20419 1744 20428 1784
rect 20468 1744 20524 1784
rect 20564 1744 20573 1784
rect 4919 1492 4928 1532
rect 4968 1492 5010 1532
rect 5050 1492 5092 1532
rect 5132 1492 5174 1532
rect 5214 1492 5256 1532
rect 5296 1492 5305 1532
rect 20039 1492 20048 1532
rect 20088 1492 20130 1532
rect 20170 1492 20212 1532
rect 20252 1492 20294 1532
rect 20334 1492 20376 1532
rect 20416 1492 20425 1532
rect 20620 1448 20660 1912
rect 20899 1828 20908 1868
rect 20948 1828 24172 1868
rect 24212 1828 24221 1868
rect 22819 1660 22828 1700
rect 22868 1660 22924 1700
rect 22964 1660 22973 1700
rect 35159 1492 35168 1532
rect 35208 1492 35250 1532
rect 35290 1492 35332 1532
rect 35372 1492 35414 1532
rect 35454 1492 35496 1532
rect 35536 1492 35545 1532
rect 16003 1408 16012 1448
rect 16052 1408 20660 1448
rect 1411 1072 1420 1112
rect 1460 1072 23788 1112
rect 23828 1072 23837 1112
rect 20227 820 20236 860
rect 20276 820 20524 860
rect 20564 820 20573 860
rect 14659 484 14668 524
rect 14708 484 28588 524
rect 28628 484 28637 524
rect 6403 400 6412 440
rect 6452 400 28108 440
rect 28148 400 28157 440
rect 6019 316 6028 356
rect 6068 316 27916 356
rect 27956 316 27965 356
rect 5731 232 5740 272
rect 5780 232 28300 272
rect 28340 232 28349 272
rect 2659 148 2668 188
rect 2708 148 27724 188
rect 27764 148 27773 188
rect 2851 64 2860 104
rect 2900 64 27532 104
rect 27572 64 27581 104
<< via4 >>
rect 4928 10564 4968 10604
rect 5010 10564 5050 10604
rect 5092 10564 5132 10604
rect 5174 10564 5214 10604
rect 5256 10564 5296 10604
rect 20048 10564 20088 10604
rect 20130 10564 20170 10604
rect 20212 10564 20252 10604
rect 20294 10564 20334 10604
rect 20376 10564 20416 10604
rect 35168 10564 35208 10604
rect 35250 10564 35290 10604
rect 35332 10564 35372 10604
rect 35414 10564 35454 10604
rect 35496 10564 35536 10604
rect 3688 9808 3728 9848
rect 3770 9808 3810 9848
rect 3852 9808 3892 9848
rect 3934 9808 3974 9848
rect 4016 9808 4056 9848
rect 18808 9808 18848 9848
rect 18890 9808 18930 9848
rect 18972 9808 19012 9848
rect 19054 9808 19094 9848
rect 19136 9808 19176 9848
rect 33928 9808 33968 9848
rect 34010 9808 34050 9848
rect 34092 9808 34132 9848
rect 34174 9808 34214 9848
rect 34256 9808 34296 9848
rect 4928 9052 4968 9092
rect 5010 9052 5050 9092
rect 5092 9052 5132 9092
rect 5174 9052 5214 9092
rect 5256 9052 5296 9092
rect 20048 9052 20088 9092
rect 20130 9052 20170 9092
rect 20212 9052 20252 9092
rect 20294 9052 20334 9092
rect 20376 9052 20416 9092
rect 35168 9052 35208 9092
rect 35250 9052 35290 9092
rect 35332 9052 35372 9092
rect 35414 9052 35454 9092
rect 35496 9052 35536 9092
rect 3688 8296 3728 8336
rect 3770 8296 3810 8336
rect 3852 8296 3892 8336
rect 3934 8296 3974 8336
rect 4016 8296 4056 8336
rect 18808 8296 18848 8336
rect 18890 8296 18930 8336
rect 18972 8296 19012 8336
rect 19054 8296 19094 8336
rect 19136 8296 19176 8336
rect 33928 8296 33968 8336
rect 34010 8296 34050 8336
rect 34092 8296 34132 8336
rect 34174 8296 34214 8336
rect 34256 8296 34296 8336
rect 4928 7540 4968 7580
rect 5010 7540 5050 7580
rect 5092 7540 5132 7580
rect 5174 7540 5214 7580
rect 5256 7540 5296 7580
rect 20048 7540 20088 7580
rect 20130 7540 20170 7580
rect 20212 7540 20252 7580
rect 20294 7540 20334 7580
rect 20376 7540 20416 7580
rect 35168 7540 35208 7580
rect 35250 7540 35290 7580
rect 35332 7540 35372 7580
rect 35414 7540 35454 7580
rect 35496 7540 35536 7580
rect 3688 6784 3728 6824
rect 3770 6784 3810 6824
rect 3852 6784 3892 6824
rect 3934 6784 3974 6824
rect 4016 6784 4056 6824
rect 18808 6784 18848 6824
rect 18890 6784 18930 6824
rect 18972 6784 19012 6824
rect 19054 6784 19094 6824
rect 19136 6784 19176 6824
rect 33928 6784 33968 6824
rect 34010 6784 34050 6824
rect 34092 6784 34132 6824
rect 34174 6784 34214 6824
rect 34256 6784 34296 6824
rect 4928 6028 4968 6068
rect 5010 6028 5050 6068
rect 5092 6028 5132 6068
rect 5174 6028 5214 6068
rect 5256 6028 5296 6068
rect 20048 6028 20088 6068
rect 20130 6028 20170 6068
rect 20212 6028 20252 6068
rect 20294 6028 20334 6068
rect 20376 6028 20416 6068
rect 35168 6028 35208 6068
rect 35250 6028 35290 6068
rect 35332 6028 35372 6068
rect 35414 6028 35454 6068
rect 35496 6028 35536 6068
rect 3688 5272 3728 5312
rect 3770 5272 3810 5312
rect 3852 5272 3892 5312
rect 3934 5272 3974 5312
rect 4016 5272 4056 5312
rect 18808 5272 18848 5312
rect 18890 5272 18930 5312
rect 18972 5272 19012 5312
rect 19054 5272 19094 5312
rect 19136 5272 19176 5312
rect 33928 5272 33968 5312
rect 34010 5272 34050 5312
rect 34092 5272 34132 5312
rect 34174 5272 34214 5312
rect 34256 5272 34296 5312
rect 4928 4516 4968 4556
rect 5010 4516 5050 4556
rect 5092 4516 5132 4556
rect 5174 4516 5214 4556
rect 5256 4516 5296 4556
rect 20048 4516 20088 4556
rect 20130 4516 20170 4556
rect 20212 4516 20252 4556
rect 20294 4516 20334 4556
rect 20376 4516 20416 4556
rect 35168 4516 35208 4556
rect 35250 4516 35290 4556
rect 35332 4516 35372 4556
rect 35414 4516 35454 4556
rect 35496 4516 35536 4556
rect 3688 3760 3728 3800
rect 3770 3760 3810 3800
rect 3852 3760 3892 3800
rect 3934 3760 3974 3800
rect 4016 3760 4056 3800
rect 18808 3760 18848 3800
rect 18890 3760 18930 3800
rect 18972 3760 19012 3800
rect 19054 3760 19094 3800
rect 19136 3760 19176 3800
rect 33928 3760 33968 3800
rect 34010 3760 34050 3800
rect 34092 3760 34132 3800
rect 34174 3760 34214 3800
rect 34256 3760 34296 3800
rect 4928 3004 4968 3044
rect 5010 3004 5050 3044
rect 5092 3004 5132 3044
rect 5174 3004 5214 3044
rect 5256 3004 5296 3044
rect 20048 3004 20088 3044
rect 20130 3004 20170 3044
rect 20212 3004 20252 3044
rect 20294 3004 20334 3044
rect 20376 3004 20416 3044
rect 35168 3004 35208 3044
rect 35250 3004 35290 3044
rect 35332 3004 35372 3044
rect 35414 3004 35454 3044
rect 35496 3004 35536 3044
rect 22924 2752 22964 2792
rect 3688 2248 3728 2288
rect 3770 2248 3810 2288
rect 3852 2248 3892 2288
rect 3934 2248 3974 2288
rect 4016 2248 4056 2288
rect 18808 2248 18848 2288
rect 18890 2248 18930 2288
rect 18972 2248 19012 2288
rect 19054 2248 19094 2288
rect 19136 2248 19176 2288
rect 33928 2248 33968 2288
rect 34010 2248 34050 2288
rect 34092 2248 34132 2288
rect 34174 2248 34214 2288
rect 34256 2248 34296 2288
rect 20524 1744 20564 1784
rect 4928 1492 4968 1532
rect 5010 1492 5050 1532
rect 5092 1492 5132 1532
rect 5174 1492 5214 1532
rect 5256 1492 5296 1532
rect 20048 1492 20088 1532
rect 20130 1492 20170 1532
rect 20212 1492 20252 1532
rect 20294 1492 20334 1532
rect 20376 1492 20416 1532
rect 22924 1660 22964 1700
rect 35168 1492 35208 1532
rect 35250 1492 35290 1532
rect 35332 1492 35372 1532
rect 35414 1492 35454 1532
rect 35496 1492 35536 1532
rect 20524 820 20564 860
<< metal5 >>
rect 3652 9848 4092 12180
rect 3652 9808 3688 9848
rect 3728 9808 3770 9848
rect 3810 9808 3852 9848
rect 3892 9808 3934 9848
rect 3974 9808 4016 9848
rect 4056 9808 4092 9848
rect 3652 8336 4092 9808
rect 3652 8296 3688 8336
rect 3728 8296 3770 8336
rect 3810 8296 3852 8336
rect 3892 8296 3934 8336
rect 3974 8296 4016 8336
rect 4056 8296 4092 8336
rect 3652 6824 4092 8296
rect 3652 6784 3688 6824
rect 3728 6784 3770 6824
rect 3810 6784 3852 6824
rect 3892 6784 3934 6824
rect 3974 6784 4016 6824
rect 4056 6784 4092 6824
rect 3652 5312 4092 6784
rect 3652 5272 3688 5312
rect 3728 5272 3770 5312
rect 3810 5272 3852 5312
rect 3892 5272 3934 5312
rect 3974 5272 4016 5312
rect 4056 5272 4092 5312
rect 3652 3800 4092 5272
rect 3652 3760 3688 3800
rect 3728 3760 3770 3800
rect 3810 3760 3852 3800
rect 3892 3760 3934 3800
rect 3974 3760 4016 3800
rect 4056 3760 4092 3800
rect 3652 2288 4092 3760
rect 3652 2248 3688 2288
rect 3728 2248 3770 2288
rect 3810 2248 3852 2288
rect 3892 2248 3934 2288
rect 3974 2248 4016 2288
rect 4056 2248 4092 2288
rect 3652 0 4092 2248
rect 4892 10604 5332 12180
rect 4892 10564 4928 10604
rect 4968 10564 5010 10604
rect 5050 10564 5092 10604
rect 5132 10564 5174 10604
rect 5214 10564 5256 10604
rect 5296 10564 5332 10604
rect 4892 9092 5332 10564
rect 4892 9052 4928 9092
rect 4968 9052 5010 9092
rect 5050 9052 5092 9092
rect 5132 9052 5174 9092
rect 5214 9052 5256 9092
rect 5296 9052 5332 9092
rect 4892 7580 5332 9052
rect 4892 7540 4928 7580
rect 4968 7540 5010 7580
rect 5050 7540 5092 7580
rect 5132 7540 5174 7580
rect 5214 7540 5256 7580
rect 5296 7540 5332 7580
rect 4892 6068 5332 7540
rect 4892 6028 4928 6068
rect 4968 6028 5010 6068
rect 5050 6028 5092 6068
rect 5132 6028 5174 6068
rect 5214 6028 5256 6068
rect 5296 6028 5332 6068
rect 4892 4556 5332 6028
rect 4892 4516 4928 4556
rect 4968 4516 5010 4556
rect 5050 4516 5092 4556
rect 5132 4516 5174 4556
rect 5214 4516 5256 4556
rect 5296 4516 5332 4556
rect 4892 3044 5332 4516
rect 4892 3004 4928 3044
rect 4968 3004 5010 3044
rect 5050 3004 5092 3044
rect 5132 3004 5174 3044
rect 5214 3004 5256 3044
rect 5296 3004 5332 3044
rect 4892 1532 5332 3004
rect 4892 1492 4928 1532
rect 4968 1492 5010 1532
rect 5050 1492 5092 1532
rect 5132 1492 5174 1532
rect 5214 1492 5256 1532
rect 5296 1492 5332 1532
rect 4892 0 5332 1492
rect 18772 9848 19212 12180
rect 18772 9808 18808 9848
rect 18848 9808 18890 9848
rect 18930 9808 18972 9848
rect 19012 9808 19054 9848
rect 19094 9808 19136 9848
rect 19176 9808 19212 9848
rect 18772 8336 19212 9808
rect 18772 8296 18808 8336
rect 18848 8296 18890 8336
rect 18930 8296 18972 8336
rect 19012 8296 19054 8336
rect 19094 8296 19136 8336
rect 19176 8296 19212 8336
rect 18772 6824 19212 8296
rect 18772 6784 18808 6824
rect 18848 6784 18890 6824
rect 18930 6784 18972 6824
rect 19012 6784 19054 6824
rect 19094 6784 19136 6824
rect 19176 6784 19212 6824
rect 18772 5312 19212 6784
rect 18772 5272 18808 5312
rect 18848 5272 18890 5312
rect 18930 5272 18972 5312
rect 19012 5272 19054 5312
rect 19094 5272 19136 5312
rect 19176 5272 19212 5312
rect 18772 3800 19212 5272
rect 18772 3760 18808 3800
rect 18848 3760 18890 3800
rect 18930 3760 18972 3800
rect 19012 3760 19054 3800
rect 19094 3760 19136 3800
rect 19176 3760 19212 3800
rect 18772 2288 19212 3760
rect 18772 2248 18808 2288
rect 18848 2248 18890 2288
rect 18930 2248 18972 2288
rect 19012 2248 19054 2288
rect 19094 2248 19136 2288
rect 19176 2248 19212 2288
rect 18772 0 19212 2248
rect 20012 10604 20452 12180
rect 20012 10564 20048 10604
rect 20088 10564 20130 10604
rect 20170 10564 20212 10604
rect 20252 10564 20294 10604
rect 20334 10564 20376 10604
rect 20416 10564 20452 10604
rect 20012 9092 20452 10564
rect 20012 9052 20048 9092
rect 20088 9052 20130 9092
rect 20170 9052 20212 9092
rect 20252 9052 20294 9092
rect 20334 9052 20376 9092
rect 20416 9052 20452 9092
rect 20012 7580 20452 9052
rect 20012 7540 20048 7580
rect 20088 7540 20130 7580
rect 20170 7540 20212 7580
rect 20252 7540 20294 7580
rect 20334 7540 20376 7580
rect 20416 7540 20452 7580
rect 20012 6068 20452 7540
rect 20012 6028 20048 6068
rect 20088 6028 20130 6068
rect 20170 6028 20212 6068
rect 20252 6028 20294 6068
rect 20334 6028 20376 6068
rect 20416 6028 20452 6068
rect 20012 4556 20452 6028
rect 20012 4516 20048 4556
rect 20088 4516 20130 4556
rect 20170 4516 20212 4556
rect 20252 4516 20294 4556
rect 20334 4516 20376 4556
rect 20416 4516 20452 4556
rect 20012 3044 20452 4516
rect 20012 3004 20048 3044
rect 20088 3004 20130 3044
rect 20170 3004 20212 3044
rect 20252 3004 20294 3044
rect 20334 3004 20376 3044
rect 20416 3004 20452 3044
rect 20012 1532 20452 3004
rect 33892 9848 34332 12180
rect 33892 9808 33928 9848
rect 33968 9808 34010 9848
rect 34050 9808 34092 9848
rect 34132 9808 34174 9848
rect 34214 9808 34256 9848
rect 34296 9808 34332 9848
rect 33892 8336 34332 9808
rect 33892 8296 33928 8336
rect 33968 8296 34010 8336
rect 34050 8296 34092 8336
rect 34132 8296 34174 8336
rect 34214 8296 34256 8336
rect 34296 8296 34332 8336
rect 33892 6824 34332 8296
rect 33892 6784 33928 6824
rect 33968 6784 34010 6824
rect 34050 6784 34092 6824
rect 34132 6784 34174 6824
rect 34214 6784 34256 6824
rect 34296 6784 34332 6824
rect 33892 5312 34332 6784
rect 33892 5272 33928 5312
rect 33968 5272 34010 5312
rect 34050 5272 34092 5312
rect 34132 5272 34174 5312
rect 34214 5272 34256 5312
rect 34296 5272 34332 5312
rect 33892 3800 34332 5272
rect 33892 3760 33928 3800
rect 33968 3760 34010 3800
rect 34050 3760 34092 3800
rect 34132 3760 34174 3800
rect 34214 3760 34256 3800
rect 34296 3760 34332 3800
rect 22924 2792 22964 2801
rect 20012 1492 20048 1532
rect 20088 1492 20130 1532
rect 20170 1492 20212 1532
rect 20252 1492 20294 1532
rect 20334 1492 20376 1532
rect 20416 1492 20452 1532
rect 20012 0 20452 1492
rect 20524 1784 20564 1793
rect 20524 860 20564 1744
rect 22924 1700 22964 2752
rect 22924 1651 22964 1660
rect 33892 2288 34332 3760
rect 33892 2248 33928 2288
rect 33968 2248 34010 2288
rect 34050 2248 34092 2288
rect 34132 2248 34174 2288
rect 34214 2248 34256 2288
rect 34296 2248 34332 2288
rect 20524 811 20564 820
rect 33892 0 34332 2248
rect 35132 10604 35572 12180
rect 35132 10564 35168 10604
rect 35208 10564 35250 10604
rect 35290 10564 35332 10604
rect 35372 10564 35414 10604
rect 35454 10564 35496 10604
rect 35536 10564 35572 10604
rect 35132 9092 35572 10564
rect 35132 9052 35168 9092
rect 35208 9052 35250 9092
rect 35290 9052 35332 9092
rect 35372 9052 35414 9092
rect 35454 9052 35496 9092
rect 35536 9052 35572 9092
rect 35132 7580 35572 9052
rect 35132 7540 35168 7580
rect 35208 7540 35250 7580
rect 35290 7540 35332 7580
rect 35372 7540 35414 7580
rect 35454 7540 35496 7580
rect 35536 7540 35572 7580
rect 35132 6068 35572 7540
rect 35132 6028 35168 6068
rect 35208 6028 35250 6068
rect 35290 6028 35332 6068
rect 35372 6028 35414 6068
rect 35454 6028 35496 6068
rect 35536 6028 35572 6068
rect 35132 4556 35572 6028
rect 35132 4516 35168 4556
rect 35208 4516 35250 4556
rect 35290 4516 35332 4556
rect 35372 4516 35414 4556
rect 35454 4516 35496 4556
rect 35536 4516 35572 4556
rect 35132 3044 35572 4516
rect 35132 3004 35168 3044
rect 35208 3004 35250 3044
rect 35290 3004 35332 3044
rect 35372 3004 35414 3044
rect 35454 3004 35496 3044
rect 35536 3004 35572 3044
rect 35132 1532 35572 3004
rect 35132 1492 35168 1532
rect 35208 1492 35250 1532
rect 35290 1492 35332 1532
rect 35372 1492 35414 1532
rect 35454 1492 35496 1532
rect 35536 1492 35572 1532
rect 35132 0 35572 1492
use sg13g2_buf_1  _000_
timestamp 1676381911
transform 1 0 16032 0 -1 4536
box -48 -56 432 834
use sg13g2_buf_1  _001_
timestamp 1676381911
transform 1 0 23712 0 -1 4536
box -48 -56 432 834
use sg13g2_buf_1  _002_
timestamp 1676381911
transform 1 0 26112 0 1 4536
box -48 -56 432 834
use sg13g2_buf_1  _003_
timestamp 1676381911
transform 1 0 25632 0 1 4536
box -48 -56 432 834
use sg13g2_buf_1  _004_
timestamp 1676381911
transform 1 0 19680 0 -1 4536
box -48 -56 432 834
use sg13g2_buf_1  _005_
timestamp 1676381911
transform 1 0 32928 0 -1 4536
box -48 -56 432 834
use sg13g2_buf_1  _006_
timestamp 1676381911
transform 1 0 31488 0 -1 4536
box -48 -56 432 834
use sg13g2_buf_1  _007_
timestamp 1676381911
transform 1 0 31200 0 1 4536
box -48 -56 432 834
use sg13g2_buf_1  _008_
timestamp 1676381911
transform 1 0 31392 0 1 6048
box -48 -56 432 834
use sg13g2_buf_1  _009_
timestamp 1676381911
transform 1 0 19392 0 -1 9072
box -48 -56 432 834
use sg13g2_buf_1  _010_
timestamp 1676381911
transform 1 0 28992 0 -1 9072
box -48 -56 432 834
use sg13g2_buf_1  _011_
timestamp 1676381911
transform 1 0 27936 0 -1 9072
box -48 -56 432 834
use sg13g2_buf_1  _012_
timestamp 1676381911
transform 1 0 25056 0 -1 9072
box -48 -56 432 834
use sg13g2_buf_1  _013_
timestamp 1676381911
transform 1 0 20832 0 -1 9072
box -48 -56 432 834
use sg13g2_buf_1  _014_
timestamp 1676381911
transform 1 0 13824 0 -1 9072
box -48 -56 432 834
use sg13g2_buf_1  _015_
timestamp 1676381911
transform 1 0 15456 0 -1 9072
box -48 -56 432 834
use sg13g2_buf_1  _016_
timestamp 1676381911
transform 1 0 18432 0 -1 9072
box -48 -56 432 834
use sg13g2_buf_1  _017_
timestamp 1676381911
transform 1 0 21696 0 -1 9072
box -48 -56 432 834
use sg13g2_buf_1  _018_
timestamp 1676381911
transform 1 0 12768 0 -1 9072
box -48 -56 432 834
use sg13g2_buf_1  _019_
timestamp 1676381911
transform 1 0 18048 0 -1 9072
box -48 -56 432 834
use sg13g2_buf_1  _020_
timestamp 1676381911
transform 1 0 13152 0 -1 9072
box -48 -56 432 834
use sg13g2_buf_1  _021_
timestamp 1676381911
transform 1 0 11424 0 1 7560
box -48 -56 432 834
use sg13g2_buf_1  _022_
timestamp 1676381911
transform 1 0 19776 0 -1 9072
box -48 -56 432 834
use sg13g2_buf_1  _023_
timestamp 1676381911
transform 1 0 10368 0 1 7560
box -48 -56 432 834
use sg13g2_buf_1  _024_
timestamp 1676381911
transform 1 0 17568 0 -1 9072
box -48 -56 432 834
use sg13g2_buf_1  _025_
timestamp 1676381911
transform 1 0 16512 0 -1 9072
box -48 -56 432 834
use sg13g2_buf_1  _026_
timestamp 1676381911
transform 1 0 18912 0 -1 9072
box -48 -56 432 834
use sg13g2_buf_1  _027_
timestamp 1676381911
transform 1 0 14976 0 -1 9072
box -48 -56 432 834
use sg13g2_buf_1  _028_
timestamp 1676381911
transform 1 0 14592 0 -1 9072
box -48 -56 432 834
use sg13g2_buf_1  _029_
timestamp 1676381911
transform 1 0 7872 0 -1 9072
box -48 -56 432 834
use sg13g2_buf_1  _030_
timestamp 1676381911
transform 1 0 11040 0 1 7560
box -48 -56 432 834
use sg13g2_buf_1  _031_
timestamp 1676381911
transform 1 0 20448 0 -1 9072
box -48 -56 432 834
use sg13g2_buf_1  _032_
timestamp 1676381911
transform 1 0 2592 0 -1 6048
box -48 -56 432 834
use sg13g2_buf_1  _033_
timestamp 1676381911
transform -1 0 6144 0 -1 7560
box -48 -56 432 834
use sg13g2_buf_1  _034_
timestamp 1676381911
transform 1 0 6336 0 -1 9072
box -48 -56 432 834
use sg13g2_buf_1  _035_
timestamp 1676381911
transform 1 0 5184 0 -1 9072
box -48 -56 432 834
use sg13g2_buf_1  _036_
timestamp 1676381911
transform -1 0 17280 0 -1 9072
box -48 -56 432 834
use sg13g2_buf_1  _037_
timestamp 1676381911
transform -1 0 29568 0 1 7560
box -48 -56 432 834
use sg13g2_buf_1  _038_
timestamp 1676381911
transform -1 0 27552 0 -1 9072
box -48 -56 432 834
use sg13g2_buf_1  _039_
timestamp 1676381911
transform -1 0 25920 0 -1 9072
box -48 -56 432 834
use sg13g2_buf_1  _040_
timestamp 1676381911
transform -1 0 23040 0 -1 9072
box -48 -56 432 834
use sg13g2_buf_1  _041_
timestamp 1676381911
transform -1 0 24672 0 -1 9072
box -48 -56 432 834
use sg13g2_buf_1  _042_
timestamp 1676381911
transform -1 0 27936 0 -1 9072
box -48 -56 432 834
use sg13g2_buf_1  _043_
timestamp 1676381911
transform -1 0 27840 0 1 6048
box -48 -56 432 834
use sg13g2_buf_1  _044_
timestamp 1676381911
transform -1 0 28224 0 1 4536
box -48 -56 432 834
use sg13g2_buf_1  _045_
timestamp 1676381911
transform -1 0 27936 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  _046_
timestamp 1676381911
transform -1 0 29280 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  _047_
timestamp 1676381911
transform -1 0 31200 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  _048_
timestamp 1676381911
transform 1 0 31680 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  _049_
timestamp 1676381911
transform 1 0 32544 0 -1 4536
box -48 -56 432 834
use sg13g2_buf_1  _050_
timestamp 1676381911
transform 1 0 32160 0 -1 4536
box -48 -56 432 834
use sg13g2_buf_1  _051_
timestamp 1676381911
transform 1 0 33312 0 1 4536
box -48 -56 432 834
use sg13g2_buf_1  _052_
timestamp 1676381911
transform 1 0 7200 0 1 4536
box -48 -56 432 834
use sg13g2_buf_1  _053_
timestamp 1676381911
transform 1 0 7584 0 1 4536
box -48 -56 432 834
use sg13g2_buf_1  _054_
timestamp 1676381911
transform 1 0 8544 0 -1 4536
box -48 -56 432 834
use sg13g2_buf_1  _055_
timestamp 1676381911
transform 1 0 8160 0 -1 4536
box -48 -56 432 834
use sg13g2_buf_1  _056_
timestamp 1676381911
transform 1 0 8064 0 1 4536
box -48 -56 432 834
use sg13g2_buf_1  _057_
timestamp 1676381911
transform 1 0 8448 0 1 4536
box -48 -56 432 834
use sg13g2_buf_1  _058_
timestamp 1676381911
transform 1 0 8832 0 1 4536
box -48 -56 432 834
use sg13g2_buf_1  _059_
timestamp 1676381911
transform 1 0 9216 0 1 4536
box -48 -56 432 834
use sg13g2_buf_1  _060_
timestamp 1676381911
transform 1 0 10080 0 1 4536
box -48 -56 432 834
use sg13g2_buf_1  _061_
timestamp 1676381911
transform 1 0 9696 0 1 4536
box -48 -56 432 834
use sg13g2_buf_1  _062_
timestamp 1676381911
transform 1 0 9888 0 -1 4536
box -48 -56 432 834
use sg13g2_buf_1  _063_
timestamp 1676381911
transform 1 0 10272 0 -1 4536
box -48 -56 432 834
use sg13g2_buf_1  _064_
timestamp 1676381911
transform 1 0 11808 0 -1 4536
box -48 -56 432 834
use sg13g2_buf_1  _065_
timestamp 1676381911
transform 1 0 12192 0 -1 4536
box -48 -56 432 834
use sg13g2_buf_1  _066_
timestamp 1676381911
transform 1 0 12576 0 -1 4536
box -48 -56 432 834
use sg13g2_buf_1  _067_
timestamp 1676381911
transform 1 0 13344 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  _068_
timestamp 1676381911
transform 1 0 13344 0 -1 4536
box -48 -56 432 834
use sg13g2_buf_1  _069_
timestamp 1676381911
transform 1 0 13728 0 -1 4536
box -48 -56 432 834
use sg13g2_buf_1  _070_
timestamp 1676381911
transform 1 0 12960 0 -1 4536
box -48 -56 432 834
use sg13g2_buf_1  _071_
timestamp 1676381911
transform 1 0 12960 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  _072_
timestamp 1676381911
transform 1 0 17664 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  _073_
timestamp 1676381911
transform 1 0 16800 0 -1 4536
box -48 -56 432 834
use sg13g2_buf_1  _074_
timestamp 1676381911
transform 1 0 18048 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  _075_
timestamp 1676381911
transform 1 0 16416 0 -1 4536
box -48 -56 432 834
use sg13g2_buf_1  _076_
timestamp 1676381911
transform 1 0 19104 0 -1 4536
box -48 -56 432 834
use sg13g2_buf_1  _077_
timestamp 1676381911
transform 1 0 18720 0 -1 4536
box -48 -56 432 834
use sg13g2_buf_1  _078_
timestamp 1676381911
transform 1 0 17568 0 1 4536
box -48 -56 432 834
use sg13g2_buf_1  _079_
timestamp 1676381911
transform 1 0 17184 0 -1 4536
box -48 -56 432 834
use sg13g2_buf_1  _080_
timestamp 1676381911
transform 1 0 18336 0 -1 4536
box -48 -56 432 834
use sg13g2_buf_1  _081_
timestamp 1676381911
transform 1 0 17952 0 -1 4536
box -48 -56 432 834
use sg13g2_buf_1  _082_
timestamp 1676381911
transform 1 0 17568 0 -1 4536
box -48 -56 432 834
use sg13g2_buf_1  _083_
timestamp 1676381911
transform 1 0 17952 0 1 4536
box -48 -56 432 834
use sg13g2_buf_1  _084_
timestamp 1676381911
transform 1 0 16992 0 1 4536
box -48 -56 432 834
use sg13g2_buf_1  _085_
timestamp 1676381911
transform 1 0 15936 0 1 4536
box -48 -56 432 834
use sg13g2_buf_1  _086_
timestamp 1676381911
transform 1 0 14304 0 -1 4536
box -48 -56 432 834
use sg13g2_buf_1  _087_
timestamp 1676381911
transform 1 0 13056 0 1 4536
box -48 -56 432 834
use sg13g2_buf_1  _088_
timestamp 1676381911
transform 1 0 21792 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  _089_
timestamp 1676381911
transform 1 0 22176 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  _090_
timestamp 1676381911
transform 1 0 22272 0 1 4536
box -48 -56 432 834
use sg13g2_buf_1  _091_
timestamp 1676381911
transform 1 0 22944 0 -1 4536
box -48 -56 432 834
use sg13g2_buf_1  _092_
timestamp 1676381911
transform 1 0 21888 0 1 4536
box -48 -56 432 834
use sg13g2_buf_1  _093_
timestamp 1676381911
transform 1 0 22560 0 -1 4536
box -48 -56 432 834
use sg13g2_buf_1  _094_
timestamp 1676381911
transform 1 0 21792 0 -1 4536
box -48 -56 432 834
use sg13g2_buf_1  _095_
timestamp 1676381911
transform 1 0 21408 0 -1 4536
box -48 -56 432 834
use sg13g2_buf_1  _096_
timestamp 1676381911
transform 1 0 22176 0 -1 4536
box -48 -56 432 834
use sg13g2_buf_1  _097_
timestamp 1676381911
transform 1 0 21024 0 -1 4536
box -48 -56 432 834
use sg13g2_buf_1  _098_
timestamp 1676381911
transform 1 0 23328 0 -1 4536
box -48 -56 432 834
use sg13g2_buf_1  _099_
timestamp 1676381911
transform 1 0 24096 0 -1 4536
box -48 -56 432 834
use sg13g2_buf_1  _100_
timestamp 1676381911
transform 1 0 25824 0 -1 4536
box -48 -56 432 834
use sg13g2_buf_1  _101_
timestamp 1676381911
transform 1 0 27168 0 -1 4536
box -48 -56 432 834
use sg13g2_buf_1  _102_
timestamp 1676381911
transform -1 0 28704 0 -1 4536
box -48 -56 432 834
use sg13g2_buf_1  _103_
timestamp 1676381911
transform -1 0 29760 0 -1 4536
box -48 -56 432 834
use sg13g2_buf_1  _104_
timestamp 1676381911
transform -1 0 2976 0 1 6048
box -48 -56 432 834
use sg13g2_decap_8  FILLER_0_0
timestamp 1679581782
transform 1 0 1152 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_7
timestamp 1679581782
transform 1 0 1824 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_14
timestamp 1679581782
transform 1 0 2496 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_21
timestamp 1679581782
transform 1 0 3168 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_28
timestamp 1679581782
transform 1 0 3840 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_35
timestamp 1679581782
transform 1 0 4512 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_42
timestamp 1679581782
transform 1 0 5184 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_49
timestamp 1679581782
transform 1 0 5856 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_56
timestamp 1679581782
transform 1 0 6528 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_63
timestamp 1679581782
transform 1 0 7200 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_70
timestamp 1679581782
transform 1 0 7872 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_77
timestamp 1679581782
transform 1 0 8544 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_84
timestamp 1679581782
transform 1 0 9216 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_91
timestamp 1679581782
transform 1 0 9888 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_98
timestamp 1679581782
transform 1 0 10560 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_105
timestamp 1679581782
transform 1 0 11232 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_112
timestamp 1679581782
transform 1 0 11904 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_119
timestamp 1679581782
transform 1 0 12576 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_126
timestamp 1679581782
transform 1 0 13248 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_133
timestamp 1679581782
transform 1 0 13920 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_140
timestamp 1679581782
transform 1 0 14592 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_147
timestamp 1679581782
transform 1 0 15264 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_154
timestamp 1679581782
transform 1 0 15936 0 1 1512
box -48 -56 720 834
use sg13g2_decap_4  FILLER_0_161
timestamp 1679577901
transform 1 0 16608 0 1 1512
box -48 -56 432 834
use sg13g2_decap_8  FILLER_0_285
timestamp 1679581782
transform 1 0 28512 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_292
timestamp 1679581782
transform 1 0 29184 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_299
timestamp 1679581782
transform 1 0 29856 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_306
timestamp 1679581782
transform 1 0 30528 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_313
timestamp 1679581782
transform 1 0 31200 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_320
timestamp 1679581782
transform 1 0 31872 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_327
timestamp 1679581782
transform 1 0 32544 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_334
timestamp 1679581782
transform 1 0 33216 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_341
timestamp 1679581782
transform 1 0 33888 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_348
timestamp 1679581782
transform 1 0 34560 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_355
timestamp 1679581782
transform 1 0 35232 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_362
timestamp 1679581782
transform 1 0 35904 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_0
timestamp 1679581782
transform 1 0 1152 0 -1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_7
timestamp 1679581782
transform 1 0 1824 0 -1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_14
timestamp 1679581782
transform 1 0 2496 0 -1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_21
timestamp 1679581782
transform 1 0 3168 0 -1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_28
timestamp 1679581782
transform 1 0 3840 0 -1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_35
timestamp 1679581782
transform 1 0 4512 0 -1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_42
timestamp 1679581782
transform 1 0 5184 0 -1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_49
timestamp 1679581782
transform 1 0 5856 0 -1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_56
timestamp 1679581782
transform 1 0 6528 0 -1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_63
timestamp 1679581782
transform 1 0 7200 0 -1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_70
timestamp 1679581782
transform 1 0 7872 0 -1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_77
timestamp 1679581782
transform 1 0 8544 0 -1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_84
timestamp 1679581782
transform 1 0 9216 0 -1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_91
timestamp 1679581782
transform 1 0 9888 0 -1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_98
timestamp 1679581782
transform 1 0 10560 0 -1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_105
timestamp 1679581782
transform 1 0 11232 0 -1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_112
timestamp 1679581782
transform 1 0 11904 0 -1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_119
timestamp 1679581782
transform 1 0 12576 0 -1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_126
timestamp 1679581782
transform 1 0 13248 0 -1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_133
timestamp 1679581782
transform 1 0 13920 0 -1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_140
timestamp 1679581782
transform 1 0 14592 0 -1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_147
timestamp 1679581782
transform 1 0 15264 0 -1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_154
timestamp 1679581782
transform 1 0 15936 0 -1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_161
timestamp 1679581782
transform 1 0 16608 0 -1 3024
box -48 -56 720 834
use sg13g2_decap_4  FILLER_1_168
timestamp 1679577901
transform 1 0 17280 0 -1 3024
box -48 -56 432 834
use sg13g2_fill_1  FILLER_1_172
timestamp 1677579658
transform 1 0 17664 0 -1 3024
box -48 -56 144 834
use sg13g2_decap_8  FILLER_1_197
timestamp 1679581782
transform 1 0 20064 0 -1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_204
timestamp 1679581782
transform 1 0 20736 0 -1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_275
timestamp 1679581782
transform 1 0 27552 0 -1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_282
timestamp 1679581782
transform 1 0 28224 0 -1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_289
timestamp 1679581782
transform 1 0 28896 0 -1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_296
timestamp 1679581782
transform 1 0 29568 0 -1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_303
timestamp 1679581782
transform 1 0 30240 0 -1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_310
timestamp 1679581782
transform 1 0 30912 0 -1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_317
timestamp 1679581782
transform 1 0 31584 0 -1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_324
timestamp 1679581782
transform 1 0 32256 0 -1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_331
timestamp 1679581782
transform 1 0 32928 0 -1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_338
timestamp 1679581782
transform 1 0 33600 0 -1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_345
timestamp 1679581782
transform 1 0 34272 0 -1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_352
timestamp 1679581782
transform 1 0 34944 0 -1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_359
timestamp 1679581782
transform 1 0 35616 0 -1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_366
timestamp 1679581782
transform 1 0 36288 0 -1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_0
timestamp 1679581782
transform 1 0 1152 0 1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_7
timestamp 1679581782
transform 1 0 1824 0 1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_14
timestamp 1679581782
transform 1 0 2496 0 1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_21
timestamp 1679581782
transform 1 0 3168 0 1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_28
timestamp 1679581782
transform 1 0 3840 0 1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_35
timestamp 1679581782
transform 1 0 4512 0 1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_42
timestamp 1679581782
transform 1 0 5184 0 1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_49
timestamp 1679581782
transform 1 0 5856 0 1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_56
timestamp 1679581782
transform 1 0 6528 0 1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_63
timestamp 1679581782
transform 1 0 7200 0 1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_70
timestamp 1679581782
transform 1 0 7872 0 1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_77
timestamp 1679581782
transform 1 0 8544 0 1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_84
timestamp 1679581782
transform 1 0 9216 0 1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_91
timestamp 1679581782
transform 1 0 9888 0 1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_98
timestamp 1679581782
transform 1 0 10560 0 1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_105
timestamp 1679581782
transform 1 0 11232 0 1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_112
timestamp 1679581782
transform 1 0 11904 0 1 3024
box -48 -56 720 834
use sg13g2_decap_4  FILLER_2_119
timestamp 1679577901
transform 1 0 12576 0 1 3024
box -48 -56 432 834
use sg13g2_decap_8  FILLER_2_131
timestamp 1679581782
transform 1 0 13728 0 1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_138
timestamp 1679581782
transform 1 0 14400 0 1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_145
timestamp 1679581782
transform 1 0 15072 0 1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_152
timestamp 1679581782
transform 1 0 15744 0 1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_159
timestamp 1679581782
transform 1 0 16416 0 1 3024
box -48 -56 720 834
use sg13g2_decap_4  FILLER_2_166
timestamp 1679577901
transform 1 0 17088 0 1 3024
box -48 -56 432 834
use sg13g2_fill_2  FILLER_2_170
timestamp 1677580104
transform 1 0 17472 0 1 3024
box -48 -56 240 834
use sg13g2_decap_8  FILLER_2_180
timestamp 1679581782
transform 1 0 18432 0 1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_187
timestamp 1679581782
transform 1 0 19104 0 1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_194
timestamp 1679581782
transform 1 0 19776 0 1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_201
timestamp 1679581782
transform 1 0 20448 0 1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_208
timestamp 1679581782
transform 1 0 21120 0 1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_223
timestamp 1679581782
transform 1 0 22560 0 1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_230
timestamp 1679581782
transform 1 0 23232 0 1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_237
timestamp 1679581782
transform 1 0 23904 0 1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_244
timestamp 1679581782
transform 1 0 24576 0 1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_251
timestamp 1679581782
transform 1 0 25248 0 1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_258
timestamp 1679581782
transform 1 0 25920 0 1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_265
timestamp 1679581782
transform 1 0 26592 0 1 3024
box -48 -56 720 834
use sg13g2_fill_2  FILLER_2_272
timestamp 1677580104
transform 1 0 27264 0 1 3024
box -48 -56 240 834
use sg13g2_fill_1  FILLER_2_274
timestamp 1677579658
transform 1 0 27456 0 1 3024
box -48 -56 144 834
use sg13g2_decap_8  FILLER_2_279
timestamp 1679581782
transform 1 0 27936 0 1 3024
box -48 -56 720 834
use sg13g2_fill_2  FILLER_2_286
timestamp 1677580104
transform 1 0 28608 0 1 3024
box -48 -56 240 834
use sg13g2_fill_1  FILLER_2_288
timestamp 1677579658
transform 1 0 28800 0 1 3024
box -48 -56 144 834
use sg13g2_decap_8  FILLER_2_293
timestamp 1679581782
transform 1 0 29280 0 1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_300
timestamp 1679581782
transform 1 0 29952 0 1 3024
box -48 -56 720 834
use sg13g2_fill_2  FILLER_2_307
timestamp 1677580104
transform 1 0 30624 0 1 3024
box -48 -56 240 834
use sg13g2_decap_4  FILLER_2_313
timestamp 1679577901
transform 1 0 31200 0 1 3024
box -48 -56 432 834
use sg13g2_fill_1  FILLER_2_317
timestamp 1677579658
transform 1 0 31584 0 1 3024
box -48 -56 144 834
use sg13g2_decap_8  FILLER_2_322
timestamp 1679581782
transform 1 0 32064 0 1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_329
timestamp 1679581782
transform 1 0 32736 0 1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_336
timestamp 1679581782
transform 1 0 33408 0 1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_343
timestamp 1679581782
transform 1 0 34080 0 1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_350
timestamp 1679581782
transform 1 0 34752 0 1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_357
timestamp 1679581782
transform 1 0 35424 0 1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_364
timestamp 1679581782
transform 1 0 36096 0 1 3024
box -48 -56 720 834
use sg13g2_decap_4  FILLER_2_371
timestamp 1679577901
transform 1 0 36768 0 1 3024
box -48 -56 432 834
use sg13g2_fill_2  FILLER_2_375
timestamp 1677580104
transform 1 0 37152 0 1 3024
box -48 -56 240 834
use sg13g2_decap_8  FILLER_3_0
timestamp 1679581782
transform 1 0 1152 0 -1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_7
timestamp 1679581782
transform 1 0 1824 0 -1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_14
timestamp 1679581782
transform 1 0 2496 0 -1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_21
timestamp 1679581782
transform 1 0 3168 0 -1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_28
timestamp 1679581782
transform 1 0 3840 0 -1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_35
timestamp 1679581782
transform 1 0 4512 0 -1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_42
timestamp 1679581782
transform 1 0 5184 0 -1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_49
timestamp 1679581782
transform 1 0 5856 0 -1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_56
timestamp 1679581782
transform 1 0 6528 0 -1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_63
timestamp 1679581782
transform 1 0 7200 0 -1 4536
box -48 -56 720 834
use sg13g2_fill_2  FILLER_3_70
timestamp 1677580104
transform 1 0 7872 0 -1 4536
box -48 -56 240 834
use sg13g2_fill_1  FILLER_3_72
timestamp 1677579658
transform 1 0 8064 0 -1 4536
box -48 -56 144 834
use sg13g2_decap_8  FILLER_3_81
timestamp 1679581782
transform 1 0 8928 0 -1 4536
box -48 -56 720 834
use sg13g2_fill_2  FILLER_3_88
timestamp 1677580104
transform 1 0 9600 0 -1 4536
box -48 -56 240 834
use sg13g2_fill_1  FILLER_3_90
timestamp 1677579658
transform 1 0 9792 0 -1 4536
box -48 -56 144 834
use sg13g2_decap_8  FILLER_3_99
timestamp 1679581782
transform 1 0 10656 0 -1 4536
box -48 -56 720 834
use sg13g2_decap_4  FILLER_3_106
timestamp 1679577901
transform 1 0 11328 0 -1 4536
box -48 -56 432 834
use sg13g2_fill_1  FILLER_3_110
timestamp 1677579658
transform 1 0 11712 0 -1 4536
box -48 -56 144 834
use sg13g2_fill_2  FILLER_3_135
timestamp 1677580104
transform 1 0 14112 0 -1 4536
box -48 -56 240 834
use sg13g2_decap_8  FILLER_3_141
timestamp 1679581782
transform 1 0 14688 0 -1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_148
timestamp 1679581782
transform 1 0 15360 0 -1 4536
box -48 -56 720 834
use sg13g2_fill_2  FILLER_3_191
timestamp 1677580104
transform 1 0 19488 0 -1 4536
box -48 -56 240 834
use sg13g2_decap_8  FILLER_3_197
timestamp 1679581782
transform 1 0 20064 0 -1 4536
box -48 -56 720 834
use sg13g2_fill_2  FILLER_3_204
timestamp 1677580104
transform 1 0 20736 0 -1 4536
box -48 -56 240 834
use sg13g2_fill_1  FILLER_3_206
timestamp 1677579658
transform 1 0 20928 0 -1 4536
box -48 -56 144 834
use sg13g2_decap_8  FILLER_3_243
timestamp 1679581782
transform 1 0 24480 0 -1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_250
timestamp 1679581782
transform 1 0 25152 0 -1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_261
timestamp 1679581782
transform 1 0 26208 0 -1 4536
box -48 -56 720 834
use sg13g2_fill_2  FILLER_3_268
timestamp 1677580104
transform 1 0 26880 0 -1 4536
box -48 -56 240 834
use sg13g2_fill_1  FILLER_3_270
timestamp 1677579658
transform 1 0 27072 0 -1 4536
box -48 -56 144 834
use sg13g2_decap_8  FILLER_3_275
timestamp 1679581782
transform 1 0 27552 0 -1 4536
box -48 -56 720 834
use sg13g2_fill_1  FILLER_3_282
timestamp 1677579658
transform 1 0 28224 0 -1 4536
box -48 -56 144 834
use sg13g2_decap_8  FILLER_3_287
timestamp 1679581782
transform 1 0 28704 0 -1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_298
timestamp 1679581782
transform 1 0 29760 0 -1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_305
timestamp 1679581782
transform 1 0 30432 0 -1 4536
box -48 -56 720 834
use sg13g2_decap_4  FILLER_3_312
timestamp 1679577901
transform 1 0 31104 0 -1 4536
box -48 -56 432 834
use sg13g2_fill_2  FILLER_3_320
timestamp 1677580104
transform 1 0 31872 0 -1 4536
box -48 -56 240 834
use sg13g2_fill_1  FILLER_3_322
timestamp 1677579658
transform 1 0 32064 0 -1 4536
box -48 -56 144 834
use sg13g2_decap_8  FILLER_3_335
timestamp 1679581782
transform 1 0 33312 0 -1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_342
timestamp 1679581782
transform 1 0 33984 0 -1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_349
timestamp 1679581782
transform 1 0 34656 0 -1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_356
timestamp 1679581782
transform 1 0 35328 0 -1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_363
timestamp 1679581782
transform 1 0 36000 0 -1 4536
box -48 -56 720 834
use sg13g2_fill_2  FILLER_3_370
timestamp 1677580104
transform 1 0 36672 0 -1 4536
box -48 -56 240 834
use sg13g2_fill_1  FILLER_3_372
timestamp 1677579658
transform 1 0 36864 0 -1 4536
box -48 -56 144 834
use sg13g2_decap_8  FILLER_4_0
timestamp 1679581782
transform 1 0 1152 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_7
timestamp 1679581782
transform 1 0 1824 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_14
timestamp 1679581782
transform 1 0 2496 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_21
timestamp 1679581782
transform 1 0 3168 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_28
timestamp 1679581782
transform 1 0 3840 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_35
timestamp 1679581782
transform 1 0 4512 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_42
timestamp 1679581782
transform 1 0 5184 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_49
timestamp 1679581782
transform 1 0 5856 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_56
timestamp 1679581782
transform 1 0 6528 0 1 4536
box -48 -56 720 834
use sg13g2_fill_1  FILLER_4_71
timestamp 1677579658
transform 1 0 7968 0 1 4536
box -48 -56 144 834
use sg13g2_fill_1  FILLER_4_88
timestamp 1677579658
transform 1 0 9600 0 1 4536
box -48 -56 144 834
use sg13g2_decap_8  FILLER_4_97
timestamp 1679581782
transform 1 0 10464 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_104
timestamp 1679581782
transform 1 0 11136 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_111
timestamp 1679581782
transform 1 0 11808 0 1 4536
box -48 -56 720 834
use sg13g2_decap_4  FILLER_4_118
timestamp 1679577901
transform 1 0 12480 0 1 4536
box -48 -56 432 834
use sg13g2_fill_2  FILLER_4_122
timestamp 1677580104
transform 1 0 12864 0 1 4536
box -48 -56 240 834
use sg13g2_decap_8  FILLER_4_128
timestamp 1679581782
transform 1 0 13440 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_135
timestamp 1679581782
transform 1 0 14112 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_142
timestamp 1679581782
transform 1 0 14784 0 1 4536
box -48 -56 720 834
use sg13g2_decap_4  FILLER_4_149
timestamp 1679577901
transform 1 0 15456 0 1 4536
box -48 -56 432 834
use sg13g2_fill_1  FILLER_4_153
timestamp 1677579658
transform 1 0 15840 0 1 4536
box -48 -56 144 834
use sg13g2_decap_8  FILLER_4_158
timestamp 1679581782
transform 1 0 16320 0 1 4536
box -48 -56 720 834
use sg13g2_fill_2  FILLER_4_169
timestamp 1677580104
transform 1 0 17376 0 1 4536
box -48 -56 240 834
use sg13g2_decap_8  FILLER_4_179
timestamp 1679581782
transform 1 0 18336 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_186
timestamp 1679581782
transform 1 0 19008 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_193
timestamp 1679581782
transform 1 0 19680 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_200
timestamp 1679581782
transform 1 0 20352 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_207
timestamp 1679581782
transform 1 0 21024 0 1 4536
box -48 -56 720 834
use sg13g2_fill_2  FILLER_4_214
timestamp 1677580104
transform 1 0 21696 0 1 4536
box -48 -56 240 834
use sg13g2_decap_8  FILLER_4_224
timestamp 1679581782
transform 1 0 22656 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_231
timestamp 1679581782
transform 1 0 23328 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_238
timestamp 1679581782
transform 1 0 24000 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_245
timestamp 1679581782
transform 1 0 24672 0 1 4536
box -48 -56 720 834
use sg13g2_fill_2  FILLER_4_252
timestamp 1677580104
transform 1 0 25344 0 1 4536
box -48 -56 240 834
use sg13g2_fill_1  FILLER_4_254
timestamp 1677579658
transform 1 0 25536 0 1 4536
box -48 -56 144 834
use sg13g2_fill_1  FILLER_4_259
timestamp 1677579658
transform 1 0 26016 0 1 4536
box -48 -56 144 834
use sg13g2_decap_8  FILLER_4_264
timestamp 1679581782
transform 1 0 26496 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_271
timestamp 1679581782
transform 1 0 27168 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_282
timestamp 1679581782
transform 1 0 28224 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_289
timestamp 1679581782
transform 1 0 28896 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_296
timestamp 1679581782
transform 1 0 29568 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_303
timestamp 1679581782
transform 1 0 30240 0 1 4536
box -48 -56 720 834
use sg13g2_fill_2  FILLER_4_310
timestamp 1677580104
transform 1 0 30912 0 1 4536
box -48 -56 240 834
use sg13g2_fill_1  FILLER_4_312
timestamp 1677579658
transform 1 0 31104 0 1 4536
box -48 -56 144 834
use sg13g2_decap_8  FILLER_4_317
timestamp 1679581782
transform 1 0 31584 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_324
timestamp 1679581782
transform 1 0 32256 0 1 4536
box -48 -56 720 834
use sg13g2_decap_4  FILLER_4_331
timestamp 1679577901
transform 1 0 32928 0 1 4536
box -48 -56 432 834
use sg13g2_decap_8  FILLER_4_339
timestamp 1679581782
transform 1 0 33696 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_346
timestamp 1679581782
transform 1 0 34368 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_353
timestamp 1679581782
transform 1 0 35040 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_360
timestamp 1679581782
transform 1 0 35712 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_367
timestamp 1679581782
transform 1 0 36384 0 1 4536
box -48 -56 720 834
use sg13g2_fill_2  FILLER_4_374
timestamp 1677580104
transform 1 0 37056 0 1 4536
box -48 -56 240 834
use sg13g2_fill_1  FILLER_4_376
timestamp 1677579658
transform 1 0 37248 0 1 4536
box -48 -56 144 834
use sg13g2_decap_8  FILLER_5_0
timestamp 1679581782
transform 1 0 1152 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_7
timestamp 1679581782
transform 1 0 1824 0 -1 6048
box -48 -56 720 834
use sg13g2_fill_1  FILLER_5_14
timestamp 1677579658
transform 1 0 2496 0 -1 6048
box -48 -56 144 834
use sg13g2_decap_8  FILLER_5_19
timestamp 1679581782
transform 1 0 2976 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_26
timestamp 1679581782
transform 1 0 3648 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_33
timestamp 1679581782
transform 1 0 4320 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_40
timestamp 1679581782
transform 1 0 4992 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_47
timestamp 1679581782
transform 1 0 5664 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_54
timestamp 1679581782
transform 1 0 6336 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_61
timestamp 1679581782
transform 1 0 7008 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_68
timestamp 1679581782
transform 1 0 7680 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_75
timestamp 1679581782
transform 1 0 8352 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_82
timestamp 1679581782
transform 1 0 9024 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_89
timestamp 1679581782
transform 1 0 9696 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_96
timestamp 1679581782
transform 1 0 10368 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_103
timestamp 1679581782
transform 1 0 11040 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_110
timestamp 1679581782
transform 1 0 11712 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_117
timestamp 1679581782
transform 1 0 12384 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_124
timestamp 1679581782
transform 1 0 13056 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_131
timestamp 1679581782
transform 1 0 13728 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_138
timestamp 1679581782
transform 1 0 14400 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_145
timestamp 1679581782
transform 1 0 15072 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_152
timestamp 1679581782
transform 1 0 15744 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_159
timestamp 1679581782
transform 1 0 16416 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_166
timestamp 1679581782
transform 1 0 17088 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_173
timestamp 1679581782
transform 1 0 17760 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_180
timestamp 1679581782
transform 1 0 18432 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_187
timestamp 1679581782
transform 1 0 19104 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_194
timestamp 1679581782
transform 1 0 19776 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_201
timestamp 1679581782
transform 1 0 20448 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_208
timestamp 1679581782
transform 1 0 21120 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_215
timestamp 1679581782
transform 1 0 21792 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_222
timestamp 1679581782
transform 1 0 22464 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_229
timestamp 1679581782
transform 1 0 23136 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_236
timestamp 1679581782
transform 1 0 23808 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_243
timestamp 1679581782
transform 1 0 24480 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_250
timestamp 1679581782
transform 1 0 25152 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_257
timestamp 1679581782
transform 1 0 25824 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_264
timestamp 1679581782
transform 1 0 26496 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_271
timestamp 1679581782
transform 1 0 27168 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_278
timestamp 1679581782
transform 1 0 27840 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_285
timestamp 1679581782
transform 1 0 28512 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_292
timestamp 1679581782
transform 1 0 29184 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_299
timestamp 1679581782
transform 1 0 29856 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_306
timestamp 1679581782
transform 1 0 30528 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_313
timestamp 1679581782
transform 1 0 31200 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_320
timestamp 1679581782
transform 1 0 31872 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_327
timestamp 1679581782
transform 1 0 32544 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_334
timestamp 1679581782
transform 1 0 33216 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_341
timestamp 1679581782
transform 1 0 33888 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_348
timestamp 1679581782
transform 1 0 34560 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_355
timestamp 1679581782
transform 1 0 35232 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_362
timestamp 1679581782
transform 1 0 35904 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_369
timestamp 1679581782
transform 1 0 36576 0 -1 6048
box -48 -56 720 834
use sg13g2_fill_1  FILLER_5_376
timestamp 1677579658
transform 1 0 37248 0 -1 6048
box -48 -56 144 834
use sg13g2_decap_8  FILLER_6_0
timestamp 1679581782
transform 1 0 1152 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_7
timestamp 1679581782
transform 1 0 1824 0 1 6048
box -48 -56 720 834
use sg13g2_fill_1  FILLER_6_14
timestamp 1677579658
transform 1 0 2496 0 1 6048
box -48 -56 144 834
use sg13g2_decap_8  FILLER_6_19
timestamp 1679581782
transform 1 0 2976 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_26
timestamp 1679581782
transform 1 0 3648 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_33
timestamp 1679581782
transform 1 0 4320 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_40
timestamp 1679581782
transform 1 0 4992 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_47
timestamp 1679581782
transform 1 0 5664 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_54
timestamp 1679581782
transform 1 0 6336 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_61
timestamp 1679581782
transform 1 0 7008 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_68
timestamp 1679581782
transform 1 0 7680 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_75
timestamp 1679581782
transform 1 0 8352 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_82
timestamp 1679581782
transform 1 0 9024 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_89
timestamp 1679581782
transform 1 0 9696 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_96
timestamp 1679581782
transform 1 0 10368 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_103
timestamp 1679581782
transform 1 0 11040 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_110
timestamp 1679581782
transform 1 0 11712 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_117
timestamp 1679581782
transform 1 0 12384 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_124
timestamp 1679581782
transform 1 0 13056 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_131
timestamp 1679581782
transform 1 0 13728 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_138
timestamp 1679581782
transform 1 0 14400 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_145
timestamp 1679581782
transform 1 0 15072 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_152
timestamp 1679581782
transform 1 0 15744 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_159
timestamp 1679581782
transform 1 0 16416 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_166
timestamp 1679581782
transform 1 0 17088 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_173
timestamp 1679581782
transform 1 0 17760 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_180
timestamp 1679581782
transform 1 0 18432 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_187
timestamp 1679581782
transform 1 0 19104 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_194
timestamp 1679581782
transform 1 0 19776 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_201
timestamp 1679581782
transform 1 0 20448 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_208
timestamp 1679581782
transform 1 0 21120 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_215
timestamp 1679581782
transform 1 0 21792 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_222
timestamp 1679581782
transform 1 0 22464 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_229
timestamp 1679581782
transform 1 0 23136 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_236
timestamp 1679581782
transform 1 0 23808 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_243
timestamp 1679581782
transform 1 0 24480 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_250
timestamp 1679581782
transform 1 0 25152 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_257
timestamp 1679581782
transform 1 0 25824 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_264
timestamp 1679581782
transform 1 0 26496 0 1 6048
box -48 -56 720 834
use sg13g2_fill_2  FILLER_6_271
timestamp 1677580104
transform 1 0 27168 0 1 6048
box -48 -56 240 834
use sg13g2_fill_1  FILLER_6_273
timestamp 1677579658
transform 1 0 27360 0 1 6048
box -48 -56 144 834
use sg13g2_decap_8  FILLER_6_278
timestamp 1679581782
transform 1 0 27840 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_285
timestamp 1679581782
transform 1 0 28512 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_292
timestamp 1679581782
transform 1 0 29184 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_299
timestamp 1679581782
transform 1 0 29856 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_306
timestamp 1679581782
transform 1 0 30528 0 1 6048
box -48 -56 720 834
use sg13g2_fill_2  FILLER_6_313
timestamp 1677580104
transform 1 0 31200 0 1 6048
box -48 -56 240 834
use sg13g2_decap_8  FILLER_6_319
timestamp 1679581782
transform 1 0 31776 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_326
timestamp 1679581782
transform 1 0 32448 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_333
timestamp 1679581782
transform 1 0 33120 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_340
timestamp 1679581782
transform 1 0 33792 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_347
timestamp 1679581782
transform 1 0 34464 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_354
timestamp 1679581782
transform 1 0 35136 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_361
timestamp 1679581782
transform 1 0 35808 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_368
timestamp 1679581782
transform 1 0 36480 0 1 6048
box -48 -56 720 834
use sg13g2_fill_2  FILLER_6_375
timestamp 1677580104
transform 1 0 37152 0 1 6048
box -48 -56 240 834
use sg13g2_decap_8  FILLER_7_0
timestamp 1679581782
transform 1 0 1152 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_7
timestamp 1679581782
transform 1 0 1824 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_14
timestamp 1679581782
transform 1 0 2496 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_21
timestamp 1679581782
transform 1 0 3168 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_28
timestamp 1679581782
transform 1 0 3840 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_35
timestamp 1679581782
transform 1 0 4512 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_4  FILLER_7_42
timestamp 1679577901
transform 1 0 5184 0 -1 7560
box -48 -56 432 834
use sg13g2_fill_2  FILLER_7_46
timestamp 1677580104
transform 1 0 5568 0 -1 7560
box -48 -56 240 834
use sg13g2_decap_8  FILLER_7_52
timestamp 1679581782
transform 1 0 6144 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_59
timestamp 1679581782
transform 1 0 6816 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_66
timestamp 1679581782
transform 1 0 7488 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_73
timestamp 1679581782
transform 1 0 8160 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_80
timestamp 1679581782
transform 1 0 8832 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_87
timestamp 1679581782
transform 1 0 9504 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_94
timestamp 1679581782
transform 1 0 10176 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_101
timestamp 1679581782
transform 1 0 10848 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_108
timestamp 1679581782
transform 1 0 11520 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_115
timestamp 1679581782
transform 1 0 12192 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_122
timestamp 1679581782
transform 1 0 12864 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_129
timestamp 1679581782
transform 1 0 13536 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_136
timestamp 1679581782
transform 1 0 14208 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_143
timestamp 1679581782
transform 1 0 14880 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_150
timestamp 1679581782
transform 1 0 15552 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_157
timestamp 1679581782
transform 1 0 16224 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_164
timestamp 1679581782
transform 1 0 16896 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_171
timestamp 1679581782
transform 1 0 17568 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_178
timestamp 1679581782
transform 1 0 18240 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_185
timestamp 1679581782
transform 1 0 18912 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_192
timestamp 1679581782
transform 1 0 19584 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_199
timestamp 1679581782
transform 1 0 20256 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_206
timestamp 1679581782
transform 1 0 20928 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_213
timestamp 1679581782
transform 1 0 21600 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_220
timestamp 1679581782
transform 1 0 22272 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_227
timestamp 1679581782
transform 1 0 22944 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_234
timestamp 1679581782
transform 1 0 23616 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_241
timestamp 1679581782
transform 1 0 24288 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_248
timestamp 1679581782
transform 1 0 24960 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_255
timestamp 1679581782
transform 1 0 25632 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_262
timestamp 1679581782
transform 1 0 26304 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_269
timestamp 1679581782
transform 1 0 26976 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_276
timestamp 1679581782
transform 1 0 27648 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_283
timestamp 1679581782
transform 1 0 28320 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_290
timestamp 1679581782
transform 1 0 28992 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_297
timestamp 1679581782
transform 1 0 29664 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_304
timestamp 1679581782
transform 1 0 30336 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_311
timestamp 1679581782
transform 1 0 31008 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_318
timestamp 1679581782
transform 1 0 31680 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_325
timestamp 1679581782
transform 1 0 32352 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_332
timestamp 1679581782
transform 1 0 33024 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_339
timestamp 1679581782
transform 1 0 33696 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_346
timestamp 1679581782
transform 1 0 34368 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_353
timestamp 1679581782
transform 1 0 35040 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_360
timestamp 1679581782
transform 1 0 35712 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_367
timestamp 1679581782
transform 1 0 36384 0 -1 7560
box -48 -56 720 834
use sg13g2_fill_2  FILLER_7_374
timestamp 1677580104
transform 1 0 37056 0 -1 7560
box -48 -56 240 834
use sg13g2_fill_1  FILLER_7_376
timestamp 1677579658
transform 1 0 37248 0 -1 7560
box -48 -56 144 834
use sg13g2_decap_8  FILLER_8_0
timestamp 1679581782
transform 1 0 1152 0 1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_7
timestamp 1679581782
transform 1 0 1824 0 1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_14
timestamp 1679581782
transform 1 0 2496 0 1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_21
timestamp 1679581782
transform 1 0 3168 0 1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_28
timestamp 1679581782
transform 1 0 3840 0 1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_35
timestamp 1679581782
transform 1 0 4512 0 1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_42
timestamp 1679581782
transform 1 0 5184 0 1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_49
timestamp 1679581782
transform 1 0 5856 0 1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_56
timestamp 1679581782
transform 1 0 6528 0 1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_63
timestamp 1679581782
transform 1 0 7200 0 1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_70
timestamp 1679581782
transform 1 0 7872 0 1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_77
timestamp 1679581782
transform 1 0 8544 0 1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_84
timestamp 1679581782
transform 1 0 9216 0 1 7560
box -48 -56 720 834
use sg13g2_decap_4  FILLER_8_91
timestamp 1679577901
transform 1 0 9888 0 1 7560
box -48 -56 432 834
use sg13g2_fill_1  FILLER_8_95
timestamp 1677579658
transform 1 0 10272 0 1 7560
box -48 -56 144 834
use sg13g2_fill_2  FILLER_8_100
timestamp 1677580104
transform 1 0 10752 0 1 7560
box -48 -56 240 834
use sg13g2_fill_1  FILLER_8_102
timestamp 1677579658
transform 1 0 10944 0 1 7560
box -48 -56 144 834
use sg13g2_decap_8  FILLER_8_111
timestamp 1679581782
transform 1 0 11808 0 1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_118
timestamp 1679581782
transform 1 0 12480 0 1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_125
timestamp 1679581782
transform 1 0 13152 0 1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_132
timestamp 1679581782
transform 1 0 13824 0 1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_139
timestamp 1679581782
transform 1 0 14496 0 1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_146
timestamp 1679581782
transform 1 0 15168 0 1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_153
timestamp 1679581782
transform 1 0 15840 0 1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_160
timestamp 1679581782
transform 1 0 16512 0 1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_167
timestamp 1679581782
transform 1 0 17184 0 1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_174
timestamp 1679581782
transform 1 0 17856 0 1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_181
timestamp 1679581782
transform 1 0 18528 0 1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_188
timestamp 1679581782
transform 1 0 19200 0 1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_195
timestamp 1679581782
transform 1 0 19872 0 1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_202
timestamp 1679581782
transform 1 0 20544 0 1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_209
timestamp 1679581782
transform 1 0 21216 0 1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_216
timestamp 1679581782
transform 1 0 21888 0 1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_223
timestamp 1679581782
transform 1 0 22560 0 1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_230
timestamp 1679581782
transform 1 0 23232 0 1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_237
timestamp 1679581782
transform 1 0 23904 0 1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_244
timestamp 1679581782
transform 1 0 24576 0 1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_251
timestamp 1679581782
transform 1 0 25248 0 1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_258
timestamp 1679581782
transform 1 0 25920 0 1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_265
timestamp 1679581782
transform 1 0 26592 0 1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_272
timestamp 1679581782
transform 1 0 27264 0 1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_279
timestamp 1679581782
transform 1 0 27936 0 1 7560
box -48 -56 720 834
use sg13g2_decap_4  FILLER_8_286
timestamp 1679577901
transform 1 0 28608 0 1 7560
box -48 -56 432 834
use sg13g2_fill_2  FILLER_8_290
timestamp 1677580104
transform 1 0 28992 0 1 7560
box -48 -56 240 834
use sg13g2_decap_8  FILLER_8_296
timestamp 1679581782
transform 1 0 29568 0 1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_303
timestamp 1679581782
transform 1 0 30240 0 1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_310
timestamp 1679581782
transform 1 0 30912 0 1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_317
timestamp 1679581782
transform 1 0 31584 0 1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_324
timestamp 1679581782
transform 1 0 32256 0 1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_331
timestamp 1679581782
transform 1 0 32928 0 1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_338
timestamp 1679581782
transform 1 0 33600 0 1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_345
timestamp 1679581782
transform 1 0 34272 0 1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_352
timestamp 1679581782
transform 1 0 34944 0 1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_359
timestamp 1679581782
transform 1 0 35616 0 1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_366
timestamp 1679581782
transform 1 0 36288 0 1 7560
box -48 -56 720 834
use sg13g2_decap_4  FILLER_8_373
timestamp 1679577901
transform 1 0 36960 0 1 7560
box -48 -56 432 834
use sg13g2_decap_8  FILLER_9_0
timestamp 1679581782
transform 1 0 1152 0 -1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_7
timestamp 1679581782
transform 1 0 1824 0 -1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_14
timestamp 1679581782
transform 1 0 2496 0 -1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_21
timestamp 1679581782
transform 1 0 3168 0 -1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_28
timestamp 1679581782
transform 1 0 3840 0 -1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_35
timestamp 1679581782
transform 1 0 4512 0 -1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_46
timestamp 1679581782
transform 1 0 5568 0 -1 9072
box -48 -56 720 834
use sg13g2_fill_1  FILLER_9_53
timestamp 1677579658
transform 1 0 6240 0 -1 9072
box -48 -56 144 834
use sg13g2_decap_8  FILLER_9_58
timestamp 1679581782
transform 1 0 6720 0 -1 9072
box -48 -56 720 834
use sg13g2_decap_4  FILLER_9_65
timestamp 1679577901
transform 1 0 7392 0 -1 9072
box -48 -56 432 834
use sg13g2_fill_1  FILLER_9_69
timestamp 1677579658
transform 1 0 7776 0 -1 9072
box -48 -56 144 834
use sg13g2_decap_8  FILLER_9_74
timestamp 1679581782
transform 1 0 8256 0 -1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_81
timestamp 1679581782
transform 1 0 8928 0 -1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_88
timestamp 1679581782
transform 1 0 9600 0 -1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_95
timestamp 1679581782
transform 1 0 10272 0 -1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_102
timestamp 1679581782
transform 1 0 10944 0 -1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_109
timestamp 1679581782
transform 1 0 11616 0 -1 9072
box -48 -56 720 834
use sg13g2_decap_4  FILLER_9_116
timestamp 1679577901
transform 1 0 12288 0 -1 9072
box -48 -56 432 834
use sg13g2_fill_1  FILLER_9_120
timestamp 1677579658
transform 1 0 12672 0 -1 9072
box -48 -56 144 834
use sg13g2_fill_2  FILLER_9_129
timestamp 1677580104
transform 1 0 13536 0 -1 9072
box -48 -56 240 834
use sg13g2_fill_1  FILLER_9_131
timestamp 1677579658
transform 1 0 13728 0 -1 9072
box -48 -56 144 834
use sg13g2_decap_4  FILLER_9_136
timestamp 1679577901
transform 1 0 14208 0 -1 9072
box -48 -56 432 834
use sg13g2_fill_1  FILLER_9_148
timestamp 1677579658
transform 1 0 15360 0 -1 9072
box -48 -56 144 834
use sg13g2_decap_8  FILLER_9_153
timestamp 1679581782
transform 1 0 15840 0 -1 9072
box -48 -56 720 834
use sg13g2_fill_2  FILLER_9_168
timestamp 1677580104
transform 1 0 17280 0 -1 9072
box -48 -56 240 834
use sg13g2_fill_1  FILLER_9_170
timestamp 1677579658
transform 1 0 17472 0 -1 9072
box -48 -56 144 834
use sg13g2_fill_1  FILLER_9_175
timestamp 1677579658
transform 1 0 17952 0 -1 9072
box -48 -56 144 834
use sg13g2_fill_1  FILLER_9_184
timestamp 1677579658
transform 1 0 18816 0 -1 9072
box -48 -56 144 834
use sg13g2_fill_1  FILLER_9_189
timestamp 1677579658
transform 1 0 19296 0 -1 9072
box -48 -56 144 834
use sg13g2_fill_2  FILLER_9_198
timestamp 1677580104
transform 1 0 20160 0 -1 9072
box -48 -56 240 834
use sg13g2_fill_1  FILLER_9_200
timestamp 1677579658
transform 1 0 20352 0 -1 9072
box -48 -56 144 834
use sg13g2_decap_4  FILLER_9_209
timestamp 1679577901
transform 1 0 21216 0 -1 9072
box -48 -56 432 834
use sg13g2_fill_1  FILLER_9_213
timestamp 1677579658
transform 1 0 21600 0 -1 9072
box -48 -56 144 834
use sg13g2_decap_4  FILLER_9_218
timestamp 1679577901
transform 1 0 22080 0 -1 9072
box -48 -56 432 834
use sg13g2_fill_2  FILLER_9_222
timestamp 1677580104
transform 1 0 22464 0 -1 9072
box -48 -56 240 834
use sg13g2_decap_8  FILLER_9_228
timestamp 1679581782
transform 1 0 23040 0 -1 9072
box -48 -56 720 834
use sg13g2_decap_4  FILLER_9_235
timestamp 1679577901
transform 1 0 23712 0 -1 9072
box -48 -56 432 834
use sg13g2_fill_2  FILLER_9_239
timestamp 1677580104
transform 1 0 24096 0 -1 9072
box -48 -56 240 834
use sg13g2_decap_4  FILLER_9_245
timestamp 1679577901
transform 1 0 24672 0 -1 9072
box -48 -56 432 834
use sg13g2_fill_1  FILLER_9_253
timestamp 1677579658
transform 1 0 25440 0 -1 9072
box -48 -56 144 834
use sg13g2_decap_8  FILLER_9_258
timestamp 1679581782
transform 1 0 25920 0 -1 9072
box -48 -56 720 834
use sg13g2_decap_4  FILLER_9_265
timestamp 1679577901
transform 1 0 26592 0 -1 9072
box -48 -56 432 834
use sg13g2_fill_2  FILLER_9_269
timestamp 1677580104
transform 1 0 26976 0 -1 9072
box -48 -56 240 834
use sg13g2_decap_8  FILLER_9_283
timestamp 1679581782
transform 1 0 28320 0 -1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_294
timestamp 1679581782
transform 1 0 29376 0 -1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_301
timestamp 1679581782
transform 1 0 30048 0 -1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_308
timestamp 1679581782
transform 1 0 30720 0 -1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_315
timestamp 1679581782
transform 1 0 31392 0 -1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_322
timestamp 1679581782
transform 1 0 32064 0 -1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_329
timestamp 1679581782
transform 1 0 32736 0 -1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_336
timestamp 1679581782
transform 1 0 33408 0 -1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_343
timestamp 1679581782
transform 1 0 34080 0 -1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_350
timestamp 1679581782
transform 1 0 34752 0 -1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_357
timestamp 1679581782
transform 1 0 35424 0 -1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_364
timestamp 1679581782
transform 1 0 36096 0 -1 9072
box -48 -56 720 834
use sg13g2_decap_4  FILLER_9_371
timestamp 1679577901
transform 1 0 36768 0 -1 9072
box -48 -56 432 834
use sg13g2_fill_2  FILLER_9_375
timestamp 1677580104
transform 1 0 37152 0 -1 9072
box -48 -56 240 834
use sg13g2_decap_8  FILLER_10_0
timestamp 1679581782
transform 1 0 1152 0 1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_7
timestamp 1679581782
transform 1 0 1824 0 1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_14
timestamp 1679581782
transform 1 0 2496 0 1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_21
timestamp 1679581782
transform 1 0 3168 0 1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_28
timestamp 1679581782
transform 1 0 3840 0 1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_35
timestamp 1679581782
transform 1 0 4512 0 1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_42
timestamp 1679581782
transform 1 0 5184 0 1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_49
timestamp 1679581782
transform 1 0 5856 0 1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_56
timestamp 1679581782
transform 1 0 6528 0 1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_63
timestamp 1679581782
transform 1 0 7200 0 1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_70
timestamp 1679581782
transform 1 0 7872 0 1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_77
timestamp 1679581782
transform 1 0 8544 0 1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_84
timestamp 1679581782
transform 1 0 9216 0 1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_91
timestamp 1679581782
transform 1 0 9888 0 1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_98
timestamp 1679581782
transform 1 0 10560 0 1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_105
timestamp 1679581782
transform 1 0 11232 0 1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_112
timestamp 1679581782
transform 1 0 11904 0 1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_119
timestamp 1679581782
transform 1 0 12576 0 1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_126
timestamp 1679581782
transform 1 0 13248 0 1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_133
timestamp 1679581782
transform 1 0 13920 0 1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_140
timestamp 1679581782
transform 1 0 14592 0 1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_147
timestamp 1679581782
transform 1 0 15264 0 1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_154
timestamp 1679581782
transform 1 0 15936 0 1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_161
timestamp 1679581782
transform 1 0 16608 0 1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_168
timestamp 1679581782
transform 1 0 17280 0 1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_175
timestamp 1679581782
transform 1 0 17952 0 1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_182
timestamp 1679581782
transform 1 0 18624 0 1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_189
timestamp 1679581782
transform 1 0 19296 0 1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_196
timestamp 1679581782
transform 1 0 19968 0 1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_203
timestamp 1679581782
transform 1 0 20640 0 1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_210
timestamp 1679581782
transform 1 0 21312 0 1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_217
timestamp 1679581782
transform 1 0 21984 0 1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_224
timestamp 1679581782
transform 1 0 22656 0 1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_231
timestamp 1679581782
transform 1 0 23328 0 1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_238
timestamp 1679581782
transform 1 0 24000 0 1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_245
timestamp 1679581782
transform 1 0 24672 0 1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_252
timestamp 1679581782
transform 1 0 25344 0 1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_259
timestamp 1679581782
transform 1 0 26016 0 1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_266
timestamp 1679581782
transform 1 0 26688 0 1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_273
timestamp 1679581782
transform 1 0 27360 0 1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_280
timestamp 1679581782
transform 1 0 28032 0 1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_287
timestamp 1679581782
transform 1 0 28704 0 1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_294
timestamp 1679581782
transform 1 0 29376 0 1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_301
timestamp 1679581782
transform 1 0 30048 0 1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_308
timestamp 1679581782
transform 1 0 30720 0 1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_315
timestamp 1679581782
transform 1 0 31392 0 1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_322
timestamp 1679581782
transform 1 0 32064 0 1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_329
timestamp 1679581782
transform 1 0 32736 0 1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_336
timestamp 1679581782
transform 1 0 33408 0 1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_343
timestamp 1679581782
transform 1 0 34080 0 1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_350
timestamp 1679581782
transform 1 0 34752 0 1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_357
timestamp 1679581782
transform 1 0 35424 0 1 9072
box -48 -56 720 834
use sg13g2_decap_4  FILLER_10_364
timestamp 1679577901
transform 1 0 36096 0 1 9072
box -48 -56 432 834
use sg13g2_fill_1  FILLER_10_368
timestamp 1677579658
transform 1 0 36480 0 1 9072
box -48 -56 144 834
use sg13g2_decap_8  FILLER_11_0
timestamp 1679581782
transform 1 0 1152 0 -1 10584
box -48 -56 720 834
use sg13g2_decap_4  FILLER_11_7
timestamp 1679577901
transform 1 0 1824 0 -1 10584
box -48 -56 432 834
use sg13g2_decap_8  FILLER_11_15
timestamp 1679581782
transform 1 0 2592 0 -1 10584
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_22
timestamp 1679581782
transform 1 0 3264 0 -1 10584
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_33
timestamp 1679581782
transform 1 0 4320 0 -1 10584
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_40
timestamp 1679581782
transform 1 0 4992 0 -1 10584
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_51
timestamp 1679581782
transform 1 0 6048 0 -1 10584
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_58
timestamp 1679581782
transform 1 0 6720 0 -1 10584
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_69
timestamp 1679581782
transform 1 0 7776 0 -1 10584
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_76
timestamp 1679581782
transform 1 0 8448 0 -1 10584
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_87
timestamp 1679581782
transform 1 0 9504 0 -1 10584
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_94
timestamp 1679581782
transform 1 0 10176 0 -1 10584
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_105
timestamp 1679581782
transform 1 0 11232 0 -1 10584
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_112
timestamp 1679581782
transform 1 0 11904 0 -1 10584
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_123
timestamp 1679581782
transform 1 0 12960 0 -1 10584
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_130
timestamp 1679581782
transform 1 0 13632 0 -1 10584
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_141
timestamp 1679581782
transform 1 0 14688 0 -1 10584
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_148
timestamp 1679581782
transform 1 0 15360 0 -1 10584
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_159
timestamp 1679581782
transform 1 0 16416 0 -1 10584
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_166
timestamp 1679581782
transform 1 0 17088 0 -1 10584
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_177
timestamp 1679581782
transform 1 0 18144 0 -1 10584
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_184
timestamp 1679581782
transform 1 0 18816 0 -1 10584
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_195
timestamp 1679581782
transform 1 0 19872 0 -1 10584
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_202
timestamp 1679581782
transform 1 0 20544 0 -1 10584
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_213
timestamp 1679581782
transform 1 0 21600 0 -1 10584
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_220
timestamp 1679581782
transform 1 0 22272 0 -1 10584
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_231
timestamp 1679581782
transform 1 0 23328 0 -1 10584
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_238
timestamp 1679581782
transform 1 0 24000 0 -1 10584
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_249
timestamp 1679581782
transform 1 0 25056 0 -1 10584
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_256
timestamp 1679581782
transform 1 0 25728 0 -1 10584
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_267
timestamp 1679581782
transform 1 0 26784 0 -1 10584
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_274
timestamp 1679581782
transform 1 0 27456 0 -1 10584
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_285
timestamp 1679581782
transform 1 0 28512 0 -1 10584
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_292
timestamp 1679581782
transform 1 0 29184 0 -1 10584
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_303
timestamp 1679581782
transform 1 0 30240 0 -1 10584
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_310
timestamp 1679581782
transform 1 0 30912 0 -1 10584
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_321
timestamp 1679581782
transform 1 0 31968 0 -1 10584
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_328
timestamp 1679581782
transform 1 0 32640 0 -1 10584
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_339
timestamp 1679581782
transform 1 0 33696 0 -1 10584
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_346
timestamp 1679581782
transform 1 0 34368 0 -1 10584
box -48 -56 720 834
use sg13g2_decap_4  FILLER_11_357
timestamp 1679577901
transform 1 0 35424 0 -1 10584
box -48 -56 432 834
use sg13g2_fill_2  FILLER_11_361
timestamp 1677580104
transform 1 0 35808 0 -1 10584
box -48 -56 240 834
use sg13g2_fill_2  FILLER_11_375
timestamp 1677580104
transform 1 0 37152 0 -1 10584
box -48 -56 240 834
use sg13g2_buf_1  output1
timestamp 1676381911
transform 1 0 36960 0 1 1512
box -48 -56 432 834
use sg13g2_buf_1  output2
timestamp 1676381911
transform 1 0 37344 0 -1 4536
box -48 -56 432 834
use sg13g2_buf_1  output3
timestamp 1676381911
transform 1 0 37728 0 -1 4536
box -48 -56 432 834
use sg13g2_buf_1  output4
timestamp 1676381911
transform 1 0 37344 0 1 4536
box -48 -56 432 834
use sg13g2_buf_1  output5
timestamp 1676381911
transform 1 0 37728 0 1 4536
box -48 -56 432 834
use sg13g2_buf_1  output6
timestamp 1676381911
transform 1 0 37344 0 -1 6048
box -48 -56 432 834
use sg13g2_buf_1  output7
timestamp 1676381911
transform 1 0 37728 0 -1 6048
box -48 -56 432 834
use sg13g2_buf_1  output8
timestamp 1676381911
transform 1 0 37344 0 1 6048
box -48 -56 432 834
use sg13g2_buf_1  output9
timestamp 1676381911
transform 1 0 37728 0 1 6048
box -48 -56 432 834
use sg13g2_buf_1  output10
timestamp 1676381911
transform 1 0 37344 0 -1 7560
box -48 -56 432 834
use sg13g2_buf_1  output11
timestamp 1676381911
transform 1 0 37728 0 -1 7560
box -48 -56 432 834
use sg13g2_buf_1  output12
timestamp 1676381911
transform 1 0 36576 0 1 1512
box -48 -56 432 834
use sg13g2_buf_1  output13
timestamp 1676381911
transform 1 0 37728 0 1 7560
box -48 -56 432 834
use sg13g2_buf_1  output14
timestamp 1676381911
transform 1 0 37344 0 1 7560
box -48 -56 432 834
use sg13g2_buf_1  output15
timestamp 1676381911
transform 1 0 37728 0 -1 9072
box -48 -56 432 834
use sg13g2_buf_1  output16
timestamp 1676381911
transform 1 0 37344 0 -1 9072
box -48 -56 432 834
use sg13g2_buf_1  output17
timestamp 1676381911
transform 1 0 37728 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  output18
timestamp 1676381911
transform 1 0 37344 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  output19
timestamp 1676381911
transform 1 0 37728 0 -1 10584
box -48 -56 432 834
use sg13g2_buf_1  output20
timestamp 1676381911
transform 1 0 37344 0 -1 10584
box -48 -56 432 834
use sg13g2_buf_1  output21
timestamp 1676381911
transform 1 0 36384 0 -1 10584
box -48 -56 432 834
use sg13g2_buf_1  output22
timestamp 1676381911
transform 1 0 36960 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  output23
timestamp 1676381911
transform 1 0 36960 0 -1 3024
box -48 -56 432 834
use sg13g2_buf_1  output24
timestamp 1676381911
transform 1 0 36000 0 -1 10584
box -48 -56 432 834
use sg13g2_buf_1  output25
timestamp 1676381911
transform 1 0 36576 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  output26
timestamp 1676381911
transform 1 0 37344 0 1 1512
box -48 -56 432 834
use sg13g2_buf_1  output27
timestamp 1676381911
transform 1 0 37728 0 1 1512
box -48 -56 432 834
use sg13g2_buf_1  output28
timestamp 1676381911
transform 1 0 37344 0 -1 3024
box -48 -56 432 834
use sg13g2_buf_1  output29
timestamp 1676381911
transform 1 0 37728 0 -1 3024
box -48 -56 432 834
use sg13g2_buf_1  output30
timestamp 1676381911
transform 1 0 37344 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  output31
timestamp 1676381911
transform 1 0 36960 0 -1 4536
box -48 -56 432 834
use sg13g2_buf_1  output32
timestamp 1676381911
transform 1 0 37728 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  output33
timestamp 1676381911
transform -1 0 4320 0 -1 10584
box -48 -56 432 834
use sg13g2_buf_1  output34
timestamp 1676381911
transform -1 0 21600 0 -1 10584
box -48 -56 432 834
use sg13g2_buf_1  output35
timestamp 1676381911
transform -1 0 23328 0 -1 10584
box -48 -56 432 834
use sg13g2_buf_1  output36
timestamp 1676381911
transform -1 0 25056 0 -1 10584
box -48 -56 432 834
use sg13g2_buf_1  output37
timestamp 1676381911
transform -1 0 26784 0 -1 10584
box -48 -56 432 834
use sg13g2_buf_1  output38
timestamp 1676381911
transform -1 0 28512 0 -1 10584
box -48 -56 432 834
use sg13g2_buf_1  output39
timestamp 1676381911
transform -1 0 30240 0 -1 10584
box -48 -56 432 834
use sg13g2_buf_1  output40
timestamp 1676381911
transform -1 0 31968 0 -1 10584
box -48 -56 432 834
use sg13g2_buf_1  output41
timestamp 1676381911
transform -1 0 33696 0 -1 10584
box -48 -56 432 834
use sg13g2_buf_1  output42
timestamp 1676381911
transform -1 0 35424 0 -1 10584
box -48 -56 432 834
use sg13g2_buf_1  output43
timestamp 1676381911
transform -1 0 37152 0 -1 10584
box -48 -56 432 834
use sg13g2_buf_1  output44
timestamp 1676381911
transform -1 0 6048 0 -1 10584
box -48 -56 432 834
use sg13g2_buf_1  output45
timestamp 1676381911
transform -1 0 7776 0 -1 10584
box -48 -56 432 834
use sg13g2_buf_1  output46
timestamp 1676381911
transform -1 0 9504 0 -1 10584
box -48 -56 432 834
use sg13g2_buf_1  output47
timestamp 1676381911
transform -1 0 11232 0 -1 10584
box -48 -56 432 834
use sg13g2_buf_1  output48
timestamp 1676381911
transform -1 0 12960 0 -1 10584
box -48 -56 432 834
use sg13g2_buf_1  output49
timestamp 1676381911
transform -1 0 14688 0 -1 10584
box -48 -56 432 834
use sg13g2_buf_1  output50
timestamp 1676381911
transform -1 0 16416 0 -1 10584
box -48 -56 432 834
use sg13g2_buf_1  output51
timestamp 1676381911
transform -1 0 18144 0 -1 10584
box -48 -56 432 834
use sg13g2_buf_1  output52
timestamp 1676381911
transform -1 0 19872 0 -1 10584
box -48 -56 432 834
use sg13g2_buf_1  output53
timestamp 1676381911
transform 1 0 16992 0 1 1512
box -48 -56 432 834
use sg13g2_buf_1  output54
timestamp 1676381911
transform -1 0 18144 0 -1 3024
box -48 -56 432 834
use sg13g2_buf_1  output55
timestamp 1676381911
transform 1 0 17376 0 1 1512
box -48 -56 432 834
use sg13g2_buf_1  output56
timestamp 1676381911
transform -1 0 18528 0 -1 3024
box -48 -56 432 834
use sg13g2_buf_1  output57
timestamp 1676381911
transform 1 0 17760 0 1 1512
box -48 -56 432 834
use sg13g2_buf_1  output58
timestamp 1676381911
transform -1 0 18912 0 -1 3024
box -48 -56 432 834
use sg13g2_buf_1  output59
timestamp 1676381911
transform 1 0 18144 0 1 1512
box -48 -56 432 834
use sg13g2_buf_1  output60
timestamp 1676381911
transform -1 0 19296 0 -1 3024
box -48 -56 432 834
use sg13g2_buf_1  output61
timestamp 1676381911
transform 1 0 18528 0 1 1512
box -48 -56 432 834
use sg13g2_buf_1  output62
timestamp 1676381911
transform -1 0 19680 0 -1 3024
box -48 -56 432 834
use sg13g2_buf_1  output63
timestamp 1676381911
transform 1 0 18912 0 1 1512
box -48 -56 432 834
use sg13g2_buf_1  output64
timestamp 1676381911
transform -1 0 20064 0 -1 3024
box -48 -56 432 834
use sg13g2_buf_1  output65
timestamp 1676381911
transform 1 0 19296 0 1 1512
box -48 -56 432 834
use sg13g2_buf_1  output66
timestamp 1676381911
transform 1 0 19680 0 1 1512
box -48 -56 432 834
use sg13g2_buf_1  output67
timestamp 1676381911
transform 1 0 20064 0 1 1512
box -48 -56 432 834
use sg13g2_buf_1  output68
timestamp 1676381911
transform -1 0 20832 0 1 1512
box -48 -56 432 834
use sg13g2_buf_1  output69
timestamp 1676381911
transform -1 0 21600 0 1 1512
box -48 -56 432 834
use sg13g2_buf_1  output70
timestamp 1676381911
transform -1 0 21216 0 1 1512
box -48 -56 432 834
use sg13g2_buf_1  output71
timestamp 1676381911
transform -1 0 21984 0 1 1512
box -48 -56 432 834
use sg13g2_buf_1  output72
timestamp 1676381911
transform -1 0 22368 0 1 1512
box -48 -56 432 834
use sg13g2_buf_1  output73
timestamp 1676381911
transform -1 0 21792 0 -1 3024
box -48 -56 432 834
use sg13g2_buf_1  output74
timestamp 1676381911
transform -1 0 23712 0 -1 3024
box -48 -56 432 834
use sg13g2_buf_1  output75
timestamp 1676381911
transform -1 0 24672 0 1 1512
box -48 -56 432 834
use sg13g2_buf_1  output76
timestamp 1676381911
transform -1 0 24096 0 -1 3024
box -48 -56 432 834
use sg13g2_buf_1  output77
timestamp 1676381911
transform -1 0 25056 0 1 1512
box -48 -56 432 834
use sg13g2_buf_1  output78
timestamp 1676381911
transform -1 0 24480 0 -1 3024
box -48 -56 432 834
use sg13g2_buf_1  output79
timestamp 1676381911
transform -1 0 25440 0 1 1512
box -48 -56 432 834
use sg13g2_buf_1  output80
timestamp 1676381911
transform -1 0 22752 0 1 1512
box -48 -56 432 834
use sg13g2_buf_1  output81
timestamp 1676381911
transform -1 0 22176 0 -1 3024
box -48 -56 432 834
use sg13g2_buf_1  output82
timestamp 1676381911
transform -1 0 23136 0 1 1512
box -48 -56 432 834
use sg13g2_buf_1  output83
timestamp 1676381911
transform -1 0 22560 0 -1 3024
box -48 -56 432 834
use sg13g2_buf_1  output84
timestamp 1676381911
transform -1 0 23520 0 1 1512
box -48 -56 432 834
use sg13g2_buf_1  output85
timestamp 1676381911
transform -1 0 22944 0 -1 3024
box -48 -56 432 834
use sg13g2_buf_1  output86
timestamp 1676381911
transform -1 0 23904 0 1 1512
box -48 -56 432 834
use sg13g2_buf_1  output87
timestamp 1676381911
transform -1 0 23328 0 -1 3024
box -48 -56 432 834
use sg13g2_buf_1  output88
timestamp 1676381911
transform -1 0 24288 0 1 1512
box -48 -56 432 834
use sg13g2_buf_1  output89
timestamp 1676381911
transform -1 0 24864 0 -1 3024
box -48 -56 432 834
use sg13g2_buf_1  output90
timestamp 1676381911
transform -1 0 26784 0 -1 3024
box -48 -56 432 834
use sg13g2_buf_1  output91
timestamp 1676381911
transform -1 0 27744 0 1 1512
box -48 -56 432 834
use sg13g2_buf_1  output92
timestamp 1676381911
transform -1 0 27168 0 -1 3024
box -48 -56 432 834
use sg13g2_buf_1  output93
timestamp 1676381911
transform -1 0 28128 0 1 1512
box -48 -56 432 834
use sg13g2_buf_1  output94
timestamp 1676381911
transform -1 0 27552 0 -1 3024
box -48 -56 432 834
use sg13g2_buf_1  output95
timestamp 1676381911
transform -1 0 28512 0 1 1512
box -48 -56 432 834
use sg13g2_buf_1  output96
timestamp 1676381911
transform -1 0 25824 0 1 1512
box -48 -56 432 834
use sg13g2_buf_1  output97
timestamp 1676381911
transform -1 0 25248 0 -1 3024
box -48 -56 432 834
use sg13g2_buf_1  output98
timestamp 1676381911
transform -1 0 26208 0 1 1512
box -48 -56 432 834
use sg13g2_buf_1  output99
timestamp 1676381911
transform -1 0 25632 0 -1 3024
box -48 -56 432 834
use sg13g2_buf_1  output100
timestamp 1676381911
transform -1 0 26592 0 1 1512
box -48 -56 432 834
use sg13g2_buf_1  output101
timestamp 1676381911
transform -1 0 26016 0 -1 3024
box -48 -56 432 834
use sg13g2_buf_1  output102
timestamp 1676381911
transform -1 0 26976 0 1 1512
box -48 -56 432 834
use sg13g2_buf_1  output103
timestamp 1676381911
transform -1 0 26400 0 -1 3024
box -48 -56 432 834
use sg13g2_buf_1  output104
timestamp 1676381911
transform -1 0 27360 0 1 1512
box -48 -56 432 834
use sg13g2_buf_1  output105
timestamp 1676381911
transform -1 0 2592 0 -1 10584
box -48 -56 432 834
<< labels >>
flabel metal2 s 0 716 90 796 0 FreeSans 320 0 0 0 FrameData[0]
port 0 nsew signal input
flabel metal2 s 0 4076 90 4156 0 FreeSans 320 0 0 0 FrameData[10]
port 1 nsew signal input
flabel metal2 s 0 4412 90 4492 0 FreeSans 320 0 0 0 FrameData[11]
port 2 nsew signal input
flabel metal2 s 0 4748 90 4828 0 FreeSans 320 0 0 0 FrameData[12]
port 3 nsew signal input
flabel metal2 s 0 5084 90 5164 0 FreeSans 320 0 0 0 FrameData[13]
port 4 nsew signal input
flabel metal2 s 0 5420 90 5500 0 FreeSans 320 0 0 0 FrameData[14]
port 5 nsew signal input
flabel metal2 s 0 5756 90 5836 0 FreeSans 320 0 0 0 FrameData[15]
port 6 nsew signal input
flabel metal2 s 0 6092 90 6172 0 FreeSans 320 0 0 0 FrameData[16]
port 7 nsew signal input
flabel metal2 s 0 6428 90 6508 0 FreeSans 320 0 0 0 FrameData[17]
port 8 nsew signal input
flabel metal2 s 0 6764 90 6844 0 FreeSans 320 0 0 0 FrameData[18]
port 9 nsew signal input
flabel metal2 s 0 7100 90 7180 0 FreeSans 320 0 0 0 FrameData[19]
port 10 nsew signal input
flabel metal2 s 0 1052 90 1132 0 FreeSans 320 0 0 0 FrameData[1]
port 11 nsew signal input
flabel metal2 s 0 7436 90 7516 0 FreeSans 320 0 0 0 FrameData[20]
port 12 nsew signal input
flabel metal2 s 0 7772 90 7852 0 FreeSans 320 0 0 0 FrameData[21]
port 13 nsew signal input
flabel metal2 s 0 8108 90 8188 0 FreeSans 320 0 0 0 FrameData[22]
port 14 nsew signal input
flabel metal2 s 0 8444 90 8524 0 FreeSans 320 0 0 0 FrameData[23]
port 15 nsew signal input
flabel metal2 s 0 8780 90 8860 0 FreeSans 320 0 0 0 FrameData[24]
port 16 nsew signal input
flabel metal2 s 0 9116 90 9196 0 FreeSans 320 0 0 0 FrameData[25]
port 17 nsew signal input
flabel metal2 s 0 9452 90 9532 0 FreeSans 320 0 0 0 FrameData[26]
port 18 nsew signal input
flabel metal2 s 0 9788 90 9868 0 FreeSans 320 0 0 0 FrameData[27]
port 19 nsew signal input
flabel metal2 s 0 10124 90 10204 0 FreeSans 320 0 0 0 FrameData[28]
port 20 nsew signal input
flabel metal2 s 0 10460 90 10540 0 FreeSans 320 0 0 0 FrameData[29]
port 21 nsew signal input
flabel metal2 s 0 1388 90 1468 0 FreeSans 320 0 0 0 FrameData[2]
port 22 nsew signal input
flabel metal2 s 0 10796 90 10876 0 FreeSans 320 0 0 0 FrameData[30]
port 23 nsew signal input
flabel metal2 s 0 11132 90 11212 0 FreeSans 320 0 0 0 FrameData[31]
port 24 nsew signal input
flabel metal2 s 0 1724 90 1804 0 FreeSans 320 0 0 0 FrameData[3]
port 25 nsew signal input
flabel metal2 s 0 2060 90 2140 0 FreeSans 320 0 0 0 FrameData[4]
port 26 nsew signal input
flabel metal2 s 0 2396 90 2476 0 FreeSans 320 0 0 0 FrameData[5]
port 27 nsew signal input
flabel metal2 s 0 2732 90 2812 0 FreeSans 320 0 0 0 FrameData[6]
port 28 nsew signal input
flabel metal2 s 0 3068 90 3148 0 FreeSans 320 0 0 0 FrameData[7]
port 29 nsew signal input
flabel metal2 s 0 3404 90 3484 0 FreeSans 320 0 0 0 FrameData[8]
port 30 nsew signal input
flabel metal2 s 0 3740 90 3820 0 FreeSans 320 0 0 0 FrameData[9]
port 31 nsew signal input
flabel metal2 s 39174 716 39264 796 0 FreeSans 320 0 0 0 FrameData_O[0]
port 32 nsew signal output
flabel metal2 s 39174 4076 39264 4156 0 FreeSans 320 0 0 0 FrameData_O[10]
port 33 nsew signal output
flabel metal2 s 39174 4412 39264 4492 0 FreeSans 320 0 0 0 FrameData_O[11]
port 34 nsew signal output
flabel metal2 s 39174 4748 39264 4828 0 FreeSans 320 0 0 0 FrameData_O[12]
port 35 nsew signal output
flabel metal2 s 39174 5084 39264 5164 0 FreeSans 320 0 0 0 FrameData_O[13]
port 36 nsew signal output
flabel metal2 s 39174 5420 39264 5500 0 FreeSans 320 0 0 0 FrameData_O[14]
port 37 nsew signal output
flabel metal2 s 39174 5756 39264 5836 0 FreeSans 320 0 0 0 FrameData_O[15]
port 38 nsew signal output
flabel metal2 s 39174 6092 39264 6172 0 FreeSans 320 0 0 0 FrameData_O[16]
port 39 nsew signal output
flabel metal2 s 39174 6428 39264 6508 0 FreeSans 320 0 0 0 FrameData_O[17]
port 40 nsew signal output
flabel metal2 s 39174 6764 39264 6844 0 FreeSans 320 0 0 0 FrameData_O[18]
port 41 nsew signal output
flabel metal2 s 39174 7100 39264 7180 0 FreeSans 320 0 0 0 FrameData_O[19]
port 42 nsew signal output
flabel metal2 s 39174 1052 39264 1132 0 FreeSans 320 0 0 0 FrameData_O[1]
port 43 nsew signal output
flabel metal2 s 39174 7436 39264 7516 0 FreeSans 320 0 0 0 FrameData_O[20]
port 44 nsew signal output
flabel metal2 s 39174 7772 39264 7852 0 FreeSans 320 0 0 0 FrameData_O[21]
port 45 nsew signal output
flabel metal2 s 39174 8108 39264 8188 0 FreeSans 320 0 0 0 FrameData_O[22]
port 46 nsew signal output
flabel metal2 s 39174 8444 39264 8524 0 FreeSans 320 0 0 0 FrameData_O[23]
port 47 nsew signal output
flabel metal2 s 39174 8780 39264 8860 0 FreeSans 320 0 0 0 FrameData_O[24]
port 48 nsew signal output
flabel metal2 s 39174 9116 39264 9196 0 FreeSans 320 0 0 0 FrameData_O[25]
port 49 nsew signal output
flabel metal2 s 39174 9452 39264 9532 0 FreeSans 320 0 0 0 FrameData_O[26]
port 50 nsew signal output
flabel metal2 s 39174 9788 39264 9868 0 FreeSans 320 0 0 0 FrameData_O[27]
port 51 nsew signal output
flabel metal2 s 39174 10124 39264 10204 0 FreeSans 320 0 0 0 FrameData_O[28]
port 52 nsew signal output
flabel metal2 s 39174 10460 39264 10540 0 FreeSans 320 0 0 0 FrameData_O[29]
port 53 nsew signal output
flabel metal2 s 39174 1388 39264 1468 0 FreeSans 320 0 0 0 FrameData_O[2]
port 54 nsew signal output
flabel metal2 s 39174 10796 39264 10876 0 FreeSans 320 0 0 0 FrameData_O[30]
port 55 nsew signal output
flabel metal2 s 39174 11132 39264 11212 0 FreeSans 320 0 0 0 FrameData_O[31]
port 56 nsew signal output
flabel metal2 s 39174 1724 39264 1804 0 FreeSans 320 0 0 0 FrameData_O[3]
port 57 nsew signal output
flabel metal2 s 39174 2060 39264 2140 0 FreeSans 320 0 0 0 FrameData_O[4]
port 58 nsew signal output
flabel metal2 s 39174 2396 39264 2476 0 FreeSans 320 0 0 0 FrameData_O[5]
port 59 nsew signal output
flabel metal2 s 39174 2732 39264 2812 0 FreeSans 320 0 0 0 FrameData_O[6]
port 60 nsew signal output
flabel metal2 s 39174 3068 39264 3148 0 FreeSans 320 0 0 0 FrameData_O[7]
port 61 nsew signal output
flabel metal2 s 39174 3404 39264 3484 0 FreeSans 320 0 0 0 FrameData_O[8]
port 62 nsew signal output
flabel metal2 s 39174 3740 39264 3820 0 FreeSans 320 0 0 0 FrameData_O[9]
port 63 nsew signal output
flabel metal3 s 27704 0 27784 80 0 FreeSans 320 0 0 0 FrameStrobe[0]
port 64 nsew signal input
flabel metal3 s 29624 0 29704 80 0 FreeSans 320 0 0 0 FrameStrobe[10]
port 65 nsew signal input
flabel metal3 s 29816 0 29896 80 0 FreeSans 320 0 0 0 FrameStrobe[11]
port 66 nsew signal input
flabel metal3 s 30008 0 30088 80 0 FreeSans 320 0 0 0 FrameStrobe[12]
port 67 nsew signal input
flabel metal3 s 30200 0 30280 80 0 FreeSans 320 0 0 0 FrameStrobe[13]
port 68 nsew signal input
flabel metal3 s 30392 0 30472 80 0 FreeSans 320 0 0 0 FrameStrobe[14]
port 69 nsew signal input
flabel metal3 s 30584 0 30664 80 0 FreeSans 320 0 0 0 FrameStrobe[15]
port 70 nsew signal input
flabel metal3 s 30776 0 30856 80 0 FreeSans 320 0 0 0 FrameStrobe[16]
port 71 nsew signal input
flabel metal3 s 30968 0 31048 80 0 FreeSans 320 0 0 0 FrameStrobe[17]
port 72 nsew signal input
flabel metal3 s 31160 0 31240 80 0 FreeSans 320 0 0 0 FrameStrobe[18]
port 73 nsew signal input
flabel metal3 s 31352 0 31432 80 0 FreeSans 320 0 0 0 FrameStrobe[19]
port 74 nsew signal input
flabel metal3 s 27896 0 27976 80 0 FreeSans 320 0 0 0 FrameStrobe[1]
port 75 nsew signal input
flabel metal3 s 28088 0 28168 80 0 FreeSans 320 0 0 0 FrameStrobe[2]
port 76 nsew signal input
flabel metal3 s 28280 0 28360 80 0 FreeSans 320 0 0 0 FrameStrobe[3]
port 77 nsew signal input
flabel metal3 s 28472 0 28552 80 0 FreeSans 320 0 0 0 FrameStrobe[4]
port 78 nsew signal input
flabel metal3 s 28664 0 28744 80 0 FreeSans 320 0 0 0 FrameStrobe[5]
port 79 nsew signal input
flabel metal3 s 28856 0 28936 80 0 FreeSans 320 0 0 0 FrameStrobe[6]
port 80 nsew signal input
flabel metal3 s 29048 0 29128 80 0 FreeSans 320 0 0 0 FrameStrobe[7]
port 81 nsew signal input
flabel metal3 s 29240 0 29320 80 0 FreeSans 320 0 0 0 FrameStrobe[8]
port 82 nsew signal input
flabel metal3 s 29432 0 29512 80 0 FreeSans 320 0 0 0 FrameStrobe[9]
port 83 nsew signal input
flabel metal3 s 3896 12100 3976 12180 0 FreeSans 320 0 0 0 FrameStrobe_O[0]
port 84 nsew signal output
flabel metal3 s 21176 12100 21256 12180 0 FreeSans 320 0 0 0 FrameStrobe_O[10]
port 85 nsew signal output
flabel metal3 s 22904 12100 22984 12180 0 FreeSans 320 0 0 0 FrameStrobe_O[11]
port 86 nsew signal output
flabel metal3 s 24632 12100 24712 12180 0 FreeSans 320 0 0 0 FrameStrobe_O[12]
port 87 nsew signal output
flabel metal3 s 26360 12100 26440 12180 0 FreeSans 320 0 0 0 FrameStrobe_O[13]
port 88 nsew signal output
flabel metal3 s 28088 12100 28168 12180 0 FreeSans 320 0 0 0 FrameStrobe_O[14]
port 89 nsew signal output
flabel metal3 s 29816 12100 29896 12180 0 FreeSans 320 0 0 0 FrameStrobe_O[15]
port 90 nsew signal output
flabel metal3 s 31544 12100 31624 12180 0 FreeSans 320 0 0 0 FrameStrobe_O[16]
port 91 nsew signal output
flabel metal3 s 33272 12100 33352 12180 0 FreeSans 320 0 0 0 FrameStrobe_O[17]
port 92 nsew signal output
flabel metal3 s 35000 12100 35080 12180 0 FreeSans 320 0 0 0 FrameStrobe_O[18]
port 93 nsew signal output
flabel metal3 s 36728 12100 36808 12180 0 FreeSans 320 0 0 0 FrameStrobe_O[19]
port 94 nsew signal output
flabel metal3 s 5624 12100 5704 12180 0 FreeSans 320 0 0 0 FrameStrobe_O[1]
port 95 nsew signal output
flabel metal3 s 7352 12100 7432 12180 0 FreeSans 320 0 0 0 FrameStrobe_O[2]
port 96 nsew signal output
flabel metal3 s 9080 12100 9160 12180 0 FreeSans 320 0 0 0 FrameStrobe_O[3]
port 97 nsew signal output
flabel metal3 s 10808 12100 10888 12180 0 FreeSans 320 0 0 0 FrameStrobe_O[4]
port 98 nsew signal output
flabel metal3 s 12536 12100 12616 12180 0 FreeSans 320 0 0 0 FrameStrobe_O[5]
port 99 nsew signal output
flabel metal3 s 14264 12100 14344 12180 0 FreeSans 320 0 0 0 FrameStrobe_O[6]
port 100 nsew signal output
flabel metal3 s 15992 12100 16072 12180 0 FreeSans 320 0 0 0 FrameStrobe_O[7]
port 101 nsew signal output
flabel metal3 s 17720 12100 17800 12180 0 FreeSans 320 0 0 0 FrameStrobe_O[8]
port 102 nsew signal output
flabel metal3 s 19448 12100 19528 12180 0 FreeSans 320 0 0 0 FrameStrobe_O[9]
port 103 nsew signal output
flabel metal3 s 7544 0 7624 80 0 FreeSans 320 0 0 0 N1END[0]
port 104 nsew signal input
flabel metal3 s 7736 0 7816 80 0 FreeSans 320 0 0 0 N1END[1]
port 105 nsew signal input
flabel metal3 s 7928 0 8008 80 0 FreeSans 320 0 0 0 N1END[2]
port 106 nsew signal input
flabel metal3 s 8120 0 8200 80 0 FreeSans 320 0 0 0 N1END[3]
port 107 nsew signal input
flabel metal3 s 9848 0 9928 80 0 FreeSans 320 0 0 0 N2END[0]
port 108 nsew signal input
flabel metal3 s 10040 0 10120 80 0 FreeSans 320 0 0 0 N2END[1]
port 109 nsew signal input
flabel metal3 s 10232 0 10312 80 0 FreeSans 320 0 0 0 N2END[2]
port 110 nsew signal input
flabel metal3 s 10424 0 10504 80 0 FreeSans 320 0 0 0 N2END[3]
port 111 nsew signal input
flabel metal3 s 10616 0 10696 80 0 FreeSans 320 0 0 0 N2END[4]
port 112 nsew signal input
flabel metal3 s 10808 0 10888 80 0 FreeSans 320 0 0 0 N2END[5]
port 113 nsew signal input
flabel metal3 s 11000 0 11080 80 0 FreeSans 320 0 0 0 N2END[6]
port 114 nsew signal input
flabel metal3 s 11192 0 11272 80 0 FreeSans 320 0 0 0 N2END[7]
port 115 nsew signal input
flabel metal3 s 8312 0 8392 80 0 FreeSans 320 0 0 0 N2MID[0]
port 116 nsew signal input
flabel metal3 s 8504 0 8584 80 0 FreeSans 320 0 0 0 N2MID[1]
port 117 nsew signal input
flabel metal3 s 8696 0 8776 80 0 FreeSans 320 0 0 0 N2MID[2]
port 118 nsew signal input
flabel metal3 s 8888 0 8968 80 0 FreeSans 320 0 0 0 N2MID[3]
port 119 nsew signal input
flabel metal3 s 9080 0 9160 80 0 FreeSans 320 0 0 0 N2MID[4]
port 120 nsew signal input
flabel metal3 s 9272 0 9352 80 0 FreeSans 320 0 0 0 N2MID[5]
port 121 nsew signal input
flabel metal3 s 9464 0 9544 80 0 FreeSans 320 0 0 0 N2MID[6]
port 122 nsew signal input
flabel metal3 s 9656 0 9736 80 0 FreeSans 320 0 0 0 N2MID[7]
port 123 nsew signal input
flabel metal3 s 11384 0 11464 80 0 FreeSans 320 0 0 0 N4END[0]
port 124 nsew signal input
flabel metal3 s 13304 0 13384 80 0 FreeSans 320 0 0 0 N4END[10]
port 125 nsew signal input
flabel metal3 s 13496 0 13576 80 0 FreeSans 320 0 0 0 N4END[11]
port 126 nsew signal input
flabel metal3 s 13688 0 13768 80 0 FreeSans 320 0 0 0 N4END[12]
port 127 nsew signal input
flabel metal3 s 13880 0 13960 80 0 FreeSans 320 0 0 0 N4END[13]
port 128 nsew signal input
flabel metal3 s 14072 0 14152 80 0 FreeSans 320 0 0 0 N4END[14]
port 129 nsew signal input
flabel metal3 s 14264 0 14344 80 0 FreeSans 320 0 0 0 N4END[15]
port 130 nsew signal input
flabel metal3 s 11576 0 11656 80 0 FreeSans 320 0 0 0 N4END[1]
port 131 nsew signal input
flabel metal3 s 11768 0 11848 80 0 FreeSans 320 0 0 0 N4END[2]
port 132 nsew signal input
flabel metal3 s 11960 0 12040 80 0 FreeSans 320 0 0 0 N4END[3]
port 133 nsew signal input
flabel metal3 s 12152 0 12232 80 0 FreeSans 320 0 0 0 N4END[4]
port 134 nsew signal input
flabel metal3 s 12344 0 12424 80 0 FreeSans 320 0 0 0 N4END[5]
port 135 nsew signal input
flabel metal3 s 12536 0 12616 80 0 FreeSans 320 0 0 0 N4END[6]
port 136 nsew signal input
flabel metal3 s 12728 0 12808 80 0 FreeSans 320 0 0 0 N4END[7]
port 137 nsew signal input
flabel metal3 s 12920 0 13000 80 0 FreeSans 320 0 0 0 N4END[8]
port 138 nsew signal input
flabel metal3 s 13112 0 13192 80 0 FreeSans 320 0 0 0 N4END[9]
port 139 nsew signal input
flabel metal3 s 14456 0 14536 80 0 FreeSans 320 0 0 0 NN4END[0]
port 140 nsew signal input
flabel metal3 s 16376 0 16456 80 0 FreeSans 320 0 0 0 NN4END[10]
port 141 nsew signal input
flabel metal3 s 16568 0 16648 80 0 FreeSans 320 0 0 0 NN4END[11]
port 142 nsew signal input
flabel metal3 s 16760 0 16840 80 0 FreeSans 320 0 0 0 NN4END[12]
port 143 nsew signal input
flabel metal3 s 16952 0 17032 80 0 FreeSans 320 0 0 0 NN4END[13]
port 144 nsew signal input
flabel metal3 s 17144 0 17224 80 0 FreeSans 320 0 0 0 NN4END[14]
port 145 nsew signal input
flabel metal3 s 17336 0 17416 80 0 FreeSans 320 0 0 0 NN4END[15]
port 146 nsew signal input
flabel metal3 s 14648 0 14728 80 0 FreeSans 320 0 0 0 NN4END[1]
port 147 nsew signal input
flabel metal3 s 14840 0 14920 80 0 FreeSans 320 0 0 0 NN4END[2]
port 148 nsew signal input
flabel metal3 s 15032 0 15112 80 0 FreeSans 320 0 0 0 NN4END[3]
port 149 nsew signal input
flabel metal3 s 15224 0 15304 80 0 FreeSans 320 0 0 0 NN4END[4]
port 150 nsew signal input
flabel metal3 s 15416 0 15496 80 0 FreeSans 320 0 0 0 NN4END[5]
port 151 nsew signal input
flabel metal3 s 15608 0 15688 80 0 FreeSans 320 0 0 0 NN4END[6]
port 152 nsew signal input
flabel metal3 s 15800 0 15880 80 0 FreeSans 320 0 0 0 NN4END[7]
port 153 nsew signal input
flabel metal3 s 15992 0 16072 80 0 FreeSans 320 0 0 0 NN4END[8]
port 154 nsew signal input
flabel metal3 s 16184 0 16264 80 0 FreeSans 320 0 0 0 NN4END[9]
port 155 nsew signal input
flabel metal3 s 17528 0 17608 80 0 FreeSans 320 0 0 0 S1BEG[0]
port 156 nsew signal output
flabel metal3 s 17720 0 17800 80 0 FreeSans 320 0 0 0 S1BEG[1]
port 157 nsew signal output
flabel metal3 s 17912 0 17992 80 0 FreeSans 320 0 0 0 S1BEG[2]
port 158 nsew signal output
flabel metal3 s 18104 0 18184 80 0 FreeSans 320 0 0 0 S1BEG[3]
port 159 nsew signal output
flabel metal3 s 18296 0 18376 80 0 FreeSans 320 0 0 0 S2BEG[0]
port 160 nsew signal output
flabel metal3 s 18488 0 18568 80 0 FreeSans 320 0 0 0 S2BEG[1]
port 161 nsew signal output
flabel metal3 s 18680 0 18760 80 0 FreeSans 320 0 0 0 S2BEG[2]
port 162 nsew signal output
flabel metal3 s 18872 0 18952 80 0 FreeSans 320 0 0 0 S2BEG[3]
port 163 nsew signal output
flabel metal3 s 19064 0 19144 80 0 FreeSans 320 0 0 0 S2BEG[4]
port 164 nsew signal output
flabel metal3 s 19256 0 19336 80 0 FreeSans 320 0 0 0 S2BEG[5]
port 165 nsew signal output
flabel metal3 s 19448 0 19528 80 0 FreeSans 320 0 0 0 S2BEG[6]
port 166 nsew signal output
flabel metal3 s 19640 0 19720 80 0 FreeSans 320 0 0 0 S2BEG[7]
port 167 nsew signal output
flabel metal3 s 19832 0 19912 80 0 FreeSans 320 0 0 0 S2BEGb[0]
port 168 nsew signal output
flabel metal3 s 20024 0 20104 80 0 FreeSans 320 0 0 0 S2BEGb[1]
port 169 nsew signal output
flabel metal3 s 20216 0 20296 80 0 FreeSans 320 0 0 0 S2BEGb[2]
port 170 nsew signal output
flabel metal3 s 20408 0 20488 80 0 FreeSans 320 0 0 0 S2BEGb[3]
port 171 nsew signal output
flabel metal3 s 20600 0 20680 80 0 FreeSans 320 0 0 0 S2BEGb[4]
port 172 nsew signal output
flabel metal3 s 20792 0 20872 80 0 FreeSans 320 0 0 0 S2BEGb[5]
port 173 nsew signal output
flabel metal3 s 20984 0 21064 80 0 FreeSans 320 0 0 0 S2BEGb[6]
port 174 nsew signal output
flabel metal3 s 21176 0 21256 80 0 FreeSans 320 0 0 0 S2BEGb[7]
port 175 nsew signal output
flabel metal3 s 21368 0 21448 80 0 FreeSans 320 0 0 0 S4BEG[0]
port 176 nsew signal output
flabel metal3 s 23288 0 23368 80 0 FreeSans 320 0 0 0 S4BEG[10]
port 177 nsew signal output
flabel metal3 s 23480 0 23560 80 0 FreeSans 320 0 0 0 S4BEG[11]
port 178 nsew signal output
flabel metal3 s 23672 0 23752 80 0 FreeSans 320 0 0 0 S4BEG[12]
port 179 nsew signal output
flabel metal3 s 23864 0 23944 80 0 FreeSans 320 0 0 0 S4BEG[13]
port 180 nsew signal output
flabel metal3 s 24056 0 24136 80 0 FreeSans 320 0 0 0 S4BEG[14]
port 181 nsew signal output
flabel metal3 s 24248 0 24328 80 0 FreeSans 320 0 0 0 S4BEG[15]
port 182 nsew signal output
flabel metal3 s 21560 0 21640 80 0 FreeSans 320 0 0 0 S4BEG[1]
port 183 nsew signal output
flabel metal3 s 21752 0 21832 80 0 FreeSans 320 0 0 0 S4BEG[2]
port 184 nsew signal output
flabel metal3 s 21944 0 22024 80 0 FreeSans 320 0 0 0 S4BEG[3]
port 185 nsew signal output
flabel metal3 s 22136 0 22216 80 0 FreeSans 320 0 0 0 S4BEG[4]
port 186 nsew signal output
flabel metal3 s 22328 0 22408 80 0 FreeSans 320 0 0 0 S4BEG[5]
port 187 nsew signal output
flabel metal3 s 22520 0 22600 80 0 FreeSans 320 0 0 0 S4BEG[6]
port 188 nsew signal output
flabel metal3 s 22712 0 22792 80 0 FreeSans 320 0 0 0 S4BEG[7]
port 189 nsew signal output
flabel metal3 s 22904 0 22984 80 0 FreeSans 320 0 0 0 S4BEG[8]
port 190 nsew signal output
flabel metal3 s 23096 0 23176 80 0 FreeSans 320 0 0 0 S4BEG[9]
port 191 nsew signal output
flabel metal3 s 24440 0 24520 80 0 FreeSans 320 0 0 0 SS4BEG[0]
port 192 nsew signal output
flabel metal3 s 26360 0 26440 80 0 FreeSans 320 0 0 0 SS4BEG[10]
port 193 nsew signal output
flabel metal3 s 26552 0 26632 80 0 FreeSans 320 0 0 0 SS4BEG[11]
port 194 nsew signal output
flabel metal3 s 26744 0 26824 80 0 FreeSans 320 0 0 0 SS4BEG[12]
port 195 nsew signal output
flabel metal3 s 26936 0 27016 80 0 FreeSans 320 0 0 0 SS4BEG[13]
port 196 nsew signal output
flabel metal3 s 27128 0 27208 80 0 FreeSans 320 0 0 0 SS4BEG[14]
port 197 nsew signal output
flabel metal3 s 27320 0 27400 80 0 FreeSans 320 0 0 0 SS4BEG[15]
port 198 nsew signal output
flabel metal3 s 24632 0 24712 80 0 FreeSans 320 0 0 0 SS4BEG[1]
port 199 nsew signal output
flabel metal3 s 24824 0 24904 80 0 FreeSans 320 0 0 0 SS4BEG[2]
port 200 nsew signal output
flabel metal3 s 25016 0 25096 80 0 FreeSans 320 0 0 0 SS4BEG[3]
port 201 nsew signal output
flabel metal3 s 25208 0 25288 80 0 FreeSans 320 0 0 0 SS4BEG[4]
port 202 nsew signal output
flabel metal3 s 25400 0 25480 80 0 FreeSans 320 0 0 0 SS4BEG[5]
port 203 nsew signal output
flabel metal3 s 25592 0 25672 80 0 FreeSans 320 0 0 0 SS4BEG[6]
port 204 nsew signal output
flabel metal3 s 25784 0 25864 80 0 FreeSans 320 0 0 0 SS4BEG[7]
port 205 nsew signal output
flabel metal3 s 25976 0 26056 80 0 FreeSans 320 0 0 0 SS4BEG[8]
port 206 nsew signal output
flabel metal3 s 26168 0 26248 80 0 FreeSans 320 0 0 0 SS4BEG[9]
port 207 nsew signal output
flabel metal3 s 27512 0 27592 80 0 FreeSans 320 0 0 0 UserCLK
port 208 nsew signal input
flabel metal3 s 2168 12100 2248 12180 0 FreeSans 320 0 0 0 UserCLKo
port 209 nsew signal output
flabel metal5 s 4892 0 5332 12180 0 FreeSans 2560 90 0 0 VGND
port 210 nsew ground bidirectional
flabel metal5 s 4892 0 5332 40 0 FreeSans 320 0 0 0 VGND
port 210 nsew ground bidirectional
flabel metal5 s 4892 12140 5332 12180 0 FreeSans 320 0 0 0 VGND
port 210 nsew ground bidirectional
flabel metal5 s 20012 0 20452 12180 0 FreeSans 2560 90 0 0 VGND
port 210 nsew ground bidirectional
flabel metal5 s 20012 0 20452 40 0 FreeSans 320 0 0 0 VGND
port 210 nsew ground bidirectional
flabel metal5 s 20012 12140 20452 12180 0 FreeSans 320 0 0 0 VGND
port 210 nsew ground bidirectional
flabel metal5 s 35132 0 35572 12180 0 FreeSans 2560 90 0 0 VGND
port 210 nsew ground bidirectional
flabel metal5 s 35132 0 35572 40 0 FreeSans 320 0 0 0 VGND
port 210 nsew ground bidirectional
flabel metal5 s 35132 12140 35572 12180 0 FreeSans 320 0 0 0 VGND
port 210 nsew ground bidirectional
flabel metal5 s 3652 0 4092 12180 0 FreeSans 2560 90 0 0 VPWR
port 211 nsew power bidirectional
flabel metal5 s 3652 0 4092 40 0 FreeSans 320 0 0 0 VPWR
port 211 nsew power bidirectional
flabel metal5 s 3652 12140 4092 12180 0 FreeSans 320 0 0 0 VPWR
port 211 nsew power bidirectional
flabel metal5 s 18772 0 19212 12180 0 FreeSans 2560 90 0 0 VPWR
port 211 nsew power bidirectional
flabel metal5 s 18772 0 19212 40 0 FreeSans 320 0 0 0 VPWR
port 211 nsew power bidirectional
flabel metal5 s 18772 12140 19212 12180 0 FreeSans 320 0 0 0 VPWR
port 211 nsew power bidirectional
flabel metal5 s 33892 0 34332 12180 0 FreeSans 2560 90 0 0 VPWR
port 211 nsew power bidirectional
flabel metal5 s 33892 0 34332 40 0 FreeSans 320 0 0 0 VPWR
port 211 nsew power bidirectional
flabel metal5 s 33892 12140 34332 12180 0 FreeSans 320 0 0 0 VPWR
port 211 nsew power bidirectional
rlabel metal1 19632 10584 19632 10584 0 VGND
rlabel metal1 19632 9828 19632 9828 0 VPWR
rlabel metal2 8096 756 8096 756 0 FrameData[0]
rlabel metal2 128 4116 128 4116 0 FrameData[10]
rlabel metal2 176 4452 176 4452 0 FrameData[11]
rlabel metal2 224 4788 224 4788 0 FrameData[12]
rlabel metal2 752 5124 752 5124 0 FrameData[13]
rlabel metal2 13920 8694 13920 8694 0 FrameData[14]
rlabel metal3 15552 7224 15552 7224 0 FrameData[15]
rlabel metal3 17184 7308 17184 7308 0 FrameData[16]
rlabel metal2 464 6468 464 6468 0 FrameData[17]
rlabel metal2 1472 6804 1472 6804 0 FrameData[18]
rlabel metal3 17280 7812 17280 7812 0 FrameData[19]
rlabel metal2 752 1092 752 1092 0 FrameData[1]
rlabel metal3 13248 8064 13248 8064 0 FrameData[20]
rlabel metal2 11520 7896 11520 7896 0 FrameData[21]
rlabel metal3 15744 8736 15744 8736 0 FrameData[22]
rlabel metal2 1232 8484 1232 8484 0 FrameData[23]
rlabel metal2 128 8820 128 8820 0 FrameData[24]
rlabel metal3 16608 8904 16608 8904 0 FrameData[25]
rlabel metal3 19008 9072 19008 9072 0 FrameData[26]
rlabel metal3 15072 9198 15072 9198 0 FrameData[27]
rlabel metal2 128 10164 128 10164 0 FrameData[28]
rlabel metal2 368 10500 368 10500 0 FrameData[29]
rlabel metal2 704 1428 704 1428 0 FrameData[2]
rlabel metal3 8640 9366 8640 9366 0 FrameData[30]
rlabel metal3 20544 9912 20544 9912 0 FrameData[31]
rlabel metal2 752 1764 752 1764 0 FrameData[3]
rlabel metal2 6512 2100 6512 2100 0 FrameData[4]
rlabel metal2 1808 2436 1808 2436 0 FrameData[5]
rlabel metal2 22752 2898 22752 2898 0 FrameData[6]
rlabel metal2 656 3108 656 3108 0 FrameData[7]
rlabel metal2 320 3444 320 3444 0 FrameData[8]
rlabel metal2 512 3780 512 3780 0 FrameData[9]
rlabel metal3 38304 1218 38304 1218 0 FrameData_O[0]
rlabel metal2 38991 4116 38991 4116 0 FrameData_O[10]
rlabel metal2 38376 4284 38376 4284 0 FrameData_O[11]
rlabel metal2 38439 4788 38439 4788 0 FrameData_O[12]
rlabel metal2 38631 5124 38631 5124 0 FrameData_O[13]
rlabel metal2 38943 5460 38943 5460 0 FrameData_O[14]
rlabel metal2 38631 5796 38631 5796 0 FrameData_O[15]
rlabel metal2 39039 6132 39039 6132 0 FrameData_O[16]
rlabel metal2 38631 6468 38631 6468 0 FrameData_O[17]
rlabel metal2 38895 6804 38895 6804 0 FrameData_O[18]
rlabel metal2 38631 7140 38631 7140 0 FrameData_O[19]
rlabel metal3 37536 1428 37536 1428 0 FrameData_O[1]
rlabel metal2 38631 7476 38631 7476 0 FrameData_O[20]
rlabel metal2 38439 7812 38439 7812 0 FrameData_O[21]
rlabel via2 39183 8148 39183 8148 0 FrameData_O[22]
rlabel metal2 38847 8484 38847 8484 0 FrameData_O[23]
rlabel metal2 38943 8820 38943 8820 0 FrameData_O[24]
rlabel metal2 38439 9156 38439 9156 0 FrameData_O[25]
rlabel metal2 38991 9492 38991 9492 0 FrameData_O[26]
rlabel metal2 38439 9828 38439 9828 0 FrameData_O[27]
rlabel metal2 38304 10122 38304 10122 0 FrameData_O[28]
rlabel metal2 37320 9660 37320 9660 0 FrameData_O[29]
rlabel metal3 38400 1932 38400 1932 0 FrameData_O[2]
rlabel metal2 36360 10416 36360 10416 0 FrameData_O[30]
rlabel metal2 36936 9660 36936 9660 0 FrameData_O[31]
rlabel metal2 38439 1764 38439 1764 0 FrameData_O[3]
rlabel metal2 38631 2100 38631 2100 0 FrameData_O[4]
rlabel metal2 38943 2436 38943 2436 0 FrameData_O[5]
rlabel metal2 38631 2772 38631 2772 0 FrameData_O[6]
rlabel metal2 38559 3108 38559 3108 0 FrameData_O[7]
rlabel metal2 37920 3696 37920 3696 0 FrameData_O[8]
rlabel metal2 38376 3612 38376 3612 0 FrameData_O[9]
rlabel metal3 2688 2898 2688 2898 0 FrameStrobe[0]
rlabel metal2 28752 8988 28752 8988 0 FrameStrobe[10]
rlabel metal2 28800 6468 28800 6468 0 FrameStrobe[11]
rlabel metal2 29088 4956 29088 4956 0 FrameStrobe[12]
rlabel metal3 30240 240 30240 240 0 FrameStrobe[13]
rlabel metal2 29808 3444 29808 3444 0 FrameStrobe[14]
rlabel metal2 30864 3444 30864 3444 0 FrameStrobe[15]
rlabel metal2 31296 3360 31296 3360 0 FrameStrobe[16]
rlabel metal2 31824 4200 31824 4200 0 FrameStrobe[17]
rlabel metal2 31440 4032 31440 4032 0 FrameStrobe[18]
rlabel metal2 31392 4914 31392 4914 0 FrameStrobe[19]
rlabel metal3 27936 198 27936 198 0 FrameStrobe[1]
rlabel metal3 28128 240 28128 240 0 FrameStrobe[2]
rlabel metal3 28320 156 28320 156 0 FrameStrobe[3]
rlabel metal3 17184 9198 17184 9198 0 FrameStrobe[4]
rlabel metal2 29088 7980 29088 7980 0 FrameStrobe[5]
rlabel metal3 28848 8652 28848 8652 0 FrameStrobe[6]
rlabel metal3 29088 1470 29088 1470 0 FrameStrobe[7]
rlabel metal3 24096 9240 24096 9240 0 FrameStrobe[8]
rlabel metal2 27024 9744 27024 9744 0 FrameStrobe[9]
rlabel metal2 3960 10416 3960 10416 0 FrameStrobe_O[0]
rlabel metal2 21240 10416 21240 10416 0 FrameStrobe_O[10]
rlabel metal2 22968 10416 22968 10416 0 FrameStrobe_O[11]
rlabel metal2 24696 10416 24696 10416 0 FrameStrobe_O[12]
rlabel metal2 26424 10416 26424 10416 0 FrameStrobe_O[13]
rlabel metal2 28152 10416 28152 10416 0 FrameStrobe_O[14]
rlabel metal2 29880 10416 29880 10416 0 FrameStrobe_O[15]
rlabel metal2 31608 10416 31608 10416 0 FrameStrobe_O[16]
rlabel metal2 33336 10416 33336 10416 0 FrameStrobe_O[17]
rlabel metal2 35064 10416 35064 10416 0 FrameStrobe_O[18]
rlabel metal2 36792 10416 36792 10416 0 FrameStrobe_O[19]
rlabel metal2 5688 10416 5688 10416 0 FrameStrobe_O[1]
rlabel metal2 7416 10416 7416 10416 0 FrameStrobe_O[2]
rlabel metal2 9144 10416 9144 10416 0 FrameStrobe_O[3]
rlabel metal2 10872 10416 10872 10416 0 FrameStrobe_O[4]
rlabel metal2 12600 10416 12600 10416 0 FrameStrobe_O[5]
rlabel metal2 14328 10416 14328 10416 0 FrameStrobe_O[6]
rlabel metal2 16056 10416 16056 10416 0 FrameStrobe_O[7]
rlabel metal2 17784 10416 17784 10416 0 FrameStrobe_O[8]
rlabel metal2 19512 10416 19512 10416 0 FrameStrobe_O[9]
rlabel metal2 7920 4116 7920 4116 0 N1END[0]
rlabel metal2 8208 4032 8208 4032 0 N1END[1]
rlabel metal2 7824 4956 7824 4956 0 N1END[2]
rlabel metal2 7728 4872 7728 4872 0 N1END[3]
rlabel metal3 9888 1752 9888 1752 0 N2END[0]
rlabel metal2 13008 4116 13008 4116 0 N2END[1]
rlabel metal3 13152 3738 13152 3738 0 N2END[2]
rlabel metal3 10464 2088 10464 2088 0 N2END[3]
rlabel metal2 13440 3402 13440 3402 0 N2END[4]
rlabel metal2 11760 4200 11760 4200 0 N2END[5]
rlabel metal2 11520 4032 11520 4032 0 N2END[6]
rlabel metal2 11568 4116 11568 4116 0 N2END[7]
rlabel metal2 8544 3864 8544 3864 0 N2MID[0]
rlabel metal2 9264 4200 9264 4200 0 N2MID[1]
rlabel metal2 9264 5124 9264 5124 0 N2MID[2]
rlabel metal2 9456 5292 9456 5292 0 N2MID[3]
rlabel metal2 9216 4956 9216 4956 0 N2MID[4]
rlabel metal2 9120 4872 9120 4872 0 N2MID[5]
rlabel metal2 9024 5040 9024 5040 0 N2MID[6]
rlabel metal2 9264 4620 9264 4620 0 N2MID[7]
rlabel metal3 11424 2508 11424 2508 0 N4END[0]
rlabel metal3 13344 744 13344 744 0 N4END[10]
rlabel metal3 13536 240 13536 240 0 N4END[11]
rlabel metal2 15216 3612 15216 3612 0 N4END[12]
rlabel metal2 16032 3360 16032 3360 0 N4END[13]
rlabel metal2 15504 4200 15504 4200 0 N4END[14]
rlabel metal3 14304 240 14304 240 0 N4END[15]
rlabel metal3 14400 3906 14400 3906 0 N4END[1]
rlabel metal3 11808 744 11808 744 0 N4END[2]
rlabel metal3 12000 2508 12000 2508 0 N4END[3]
rlabel metal3 12192 450 12192 450 0 N4END[4]
rlabel metal3 12384 744 12384 744 0 N4END[5]
rlabel metal3 12576 702 12576 702 0 N4END[6]
rlabel metal3 12768 534 12768 534 0 N4END[7]
rlabel metal3 12960 1626 12960 1626 0 N4END[8]
rlabel metal3 13152 786 13152 786 0 N4END[9]
rlabel metal3 14496 240 14496 240 0 NN4END[0]
rlabel metal3 16416 576 16416 576 0 NN4END[10]
rlabel metal3 16608 240 16608 240 0 NN4END[11]
rlabel metal3 16800 408 16800 408 0 NN4END[12]
rlabel metal3 16992 1470 16992 1470 0 NN4END[13]
rlabel metal3 17184 324 17184 324 0 NN4END[14]
rlabel metal3 17376 744 17376 744 0 NN4END[15]
rlabel metal3 14688 282 14688 282 0 NN4END[1]
rlabel metal2 15360 3696 15360 3696 0 NN4END[2]
rlabel via2 15072 72 15072 72 0 NN4END[3]
rlabel metal3 15264 492 15264 492 0 NN4END[4]
rlabel metal3 15456 198 15456 198 0 NN4END[5]
rlabel metal3 15648 618 15648 618 0 NN4END[6]
rlabel metal3 15840 282 15840 282 0 NN4END[7]
rlabel metal3 16032 744 16032 744 0 NN4END[8]
rlabel metal3 16224 366 16224 366 0 NN4END[9]
rlabel metal3 17568 870 17568 870 0 S1BEG[0]
rlabel metal3 17760 1248 17760 1248 0 S1BEG[1]
rlabel metal3 17952 870 17952 870 0 S1BEG[2]
rlabel metal3 18144 1248 18144 1248 0 S1BEG[3]
rlabel metal3 18336 870 18336 870 0 S2BEG[0]
rlabel metal3 18528 1248 18528 1248 0 S2BEG[1]
rlabel metal3 18720 618 18720 618 0 S2BEG[2]
rlabel metal3 18912 660 18912 660 0 S2BEG[3]
rlabel metal3 19104 870 19104 870 0 S2BEG[4]
rlabel metal3 19296 1248 19296 1248 0 S2BEG[5]
rlabel metal3 19488 870 19488 870 0 S2BEG[6]
rlabel metal3 19680 1248 19680 1248 0 S2BEG[7]
rlabel metal3 19872 912 19872 912 0 S2BEGb[0]
rlabel metal3 20064 450 20064 450 0 S2BEGb[1]
rlabel metal3 20256 450 20256 450 0 S2BEGb[2]
rlabel metal3 20448 450 20448 450 0 S2BEGb[3]
rlabel metal3 20640 912 20640 912 0 S2BEGb[4]
rlabel metal3 20832 870 20832 870 0 S2BEGb[5]
rlabel metal3 21024 870 21024 870 0 S2BEGb[6]
rlabel metal3 21216 1038 21216 1038 0 S2BEGb[7]
rlabel metal3 21408 1248 21408 1248 0 S4BEG[0]
rlabel metal3 23328 1248 23328 1248 0 S4BEG[10]
rlabel metal3 23520 828 23520 828 0 S4BEG[11]
rlabel metal3 23712 1248 23712 1248 0 S4BEG[12]
rlabel metal3 23904 912 23904 912 0 S4BEG[13]
rlabel metal3 24096 1248 24096 1248 0 S4BEG[14]
rlabel metal3 24288 828 24288 828 0 S4BEG[15]
rlabel metal3 21600 912 21600 912 0 S4BEG[1]
rlabel metal3 21792 1248 21792 1248 0 S4BEG[2]
rlabel metal3 21984 870 21984 870 0 S4BEG[3]
rlabel metal3 22176 1248 22176 1248 0 S4BEG[4]
rlabel metal3 22368 1038 22368 1038 0 S4BEG[5]
rlabel metal3 22560 1248 22560 1248 0 S4BEG[6]
rlabel metal3 22752 912 22752 912 0 S4BEG[7]
rlabel metal3 22944 1248 22944 1248 0 S4BEG[8]
rlabel metal3 23136 870 23136 870 0 S4BEG[9]
rlabel metal3 24480 1248 24480 1248 0 SS4BEG[0]
rlabel metal3 26400 1248 26400 1248 0 SS4BEG[10]
rlabel metal3 26592 912 26592 912 0 SS4BEG[11]
rlabel metal3 26784 1248 26784 1248 0 SS4BEG[12]
rlabel metal3 26976 828 26976 828 0 SS4BEG[13]
rlabel metal3 27168 1248 27168 1248 0 SS4BEG[14]
rlabel metal3 27360 828 27360 828 0 SS4BEG[15]
rlabel metal3 24672 828 24672 828 0 SS4BEG[1]
rlabel metal3 24864 1248 24864 1248 0 SS4BEG[2]
rlabel metal3 25056 912 25056 912 0 SS4BEG[3]
rlabel metal3 25248 1248 25248 1248 0 SS4BEG[4]
rlabel metal3 25440 828 25440 828 0 SS4BEG[5]
rlabel metal3 25632 1248 25632 1248 0 SS4BEG[6]
rlabel metal3 25824 828 25824 828 0 SS4BEG[7]
rlabel metal3 26016 1248 26016 1248 0 SS4BEG[8]
rlabel metal3 26208 1038 26208 1038 0 SS4BEG[9]
rlabel via3 27552 72 27552 72 0 UserCLK
rlabel metal2 2232 10416 2232 10416 0 UserCLKo
rlabel metal2 37056 1974 37056 1974 0 net1
rlabel metal3 14400 7980 14400 7980 0 net10
rlabel metal2 22968 3948 22968 3948 0 net100
rlabel metal3 22560 3612 22560 3612 0 net101
rlabel metal3 22752 3612 22752 3612 0 net102
rlabel metal3 23520 3990 23520 3990 0 net103
rlabel metal3 21408 3780 21408 3780 0 net104
rlabel metal2 2664 6636 2664 6636 0 net105
rlabel metal2 37824 7098 37824 7098 0 net11
rlabel metal2 34128 1932 34128 1932 0 net12
rlabel metal2 37824 8022 37824 8022 0 net13
rlabel metal2 37440 7812 37440 7812 0 net14
rlabel metal2 37824 8820 37824 8820 0 net15
rlabel metal2 37056 8652 37056 8652 0 net16
rlabel metal3 37632 9198 37632 9198 0 net17
rlabel metal2 37344 9492 37344 9492 0 net18
rlabel metal3 37824 10458 37824 10458 0 net19
rlabel metal2 37440 4158 37440 4158 0 net2
rlabel metal2 37296 10164 37296 10164 0 net20
rlabel metal2 36480 10248 36480 10248 0 net21
rlabel metal2 37056 9534 37056 9534 0 net22
rlabel metal3 33216 3612 33216 3612 0 net23
rlabel metal2 36096 10206 36096 10206 0 net24
rlabel metal2 22632 8568 22632 8568 0 net25
rlabel metal3 37632 3192 37632 3192 0 net26
rlabel metal2 37824 2016 37824 2016 0 net27
rlabel metal3 37536 3318 37536 3318 0 net28
rlabel metal2 37824 2646 37824 2646 0 net29
rlabel metal2 37872 4116 37872 4116 0 net3
rlabel metal3 32352 4074 32352 4074 0 net30
rlabel metal2 36528 4116 36528 4116 0 net31
rlabel metal2 37824 3570 37824 3570 0 net32
rlabel metal2 3576 5628 3576 5628 0 net33
rlabel metal2 21504 10206 21504 10206 0 net34
rlabel metal2 25368 6636 25368 6636 0 net35
rlabel metal2 27144 5124 27144 5124 0 net36
rlabel metal2 27144 3612 27144 3612 0 net37
rlabel metal2 28680 3612 28680 3612 0 net38
rlabel metal2 30504 3612 30504 3612 0 net39
rlabel metal3 37536 6888 37536 6888 0 net4
rlabel metal2 31944 3612 31944 3612 0 net40
rlabel metal2 32904 4284 32904 4284 0 net41
rlabel metal2 35328 10122 35328 10122 0 net42
rlabel metal2 34632 5124 34632 5124 0 net43
rlabel metal2 5880 7056 5880 7056 0 net44
rlabel metal2 7176 8904 7176 8904 0 net45
rlabel metal2 5640 8904 5640 8904 0 net46
rlabel metal2 16392 8904 16392 8904 0 net47
rlabel metal2 20544 10458 20544 10458 0 net48
rlabel metal3 14592 10458 14592 10458 0 net49
rlabel metal2 37776 4956 37776 4956 0 net5
rlabel metal3 20160 9828 20160 9828 0 net50
rlabel metal2 22680 8820 22680 8820 0 net51
rlabel metal2 19872 10122 19872 10122 0 net52
rlabel metal2 16848 1932 16848 1932 0 net53
rlabel metal2 18096 2604 18096 2604 0 net54
rlabel metal2 17520 1932 17520 1932 0 net55
rlabel metal2 16464 2688 16464 2688 0 net56
rlabel metal2 17904 2016 17904 2016 0 net57
rlabel metal3 9024 4536 9024 4536 0 net58
rlabel metal4 17712 1932 17712 1932 0 net59
rlabel metal3 14304 7140 14304 7140 0 net6
rlabel metal2 17568 2352 17568 2352 0 net60
rlabel metal2 15888 1848 15888 1848 0 net61
rlabel metal2 17952 2856 17952 2856 0 net62
rlabel metal2 17808 2100 17808 2100 0 net63
rlabel metal2 19248 2688 19248 2688 0 net64
rlabel metal3 19392 2982 19392 2982 0 net65
rlabel metal2 14592 3150 14592 3150 0 net66
rlabel metal2 20112 1932 20112 1932 0 net67
rlabel metal2 20736 1974 20736 1974 0 net68
rlabel metal2 21024 1848 21024 1848 0 net69
rlabel metal2 37824 5670 37824 5670 0 net7
rlabel metal2 21072 1932 21072 1932 0 net70
rlabel metal2 16320 2184 16320 2184 0 net71
rlabel metal2 17184 1512 17184 1512 0 net72
rlabel metal2 20688 3276 20688 3276 0 net73
rlabel metal2 19824 3696 19824 3696 0 net74
rlabel metal2 20640 4620 20640 4620 0 net75
rlabel metal2 19440 4368 19440 4368 0 net76
rlabel metal2 19224 5040 19224 5040 0 net77
rlabel metal2 18960 2184 18960 2184 0 net78
rlabel metal2 24768 2100 24768 2100 0 net79
rlabel metal2 37440 6510 37440 6510 0 net8
rlabel metal2 22368 2100 22368 2100 0 net80
rlabel metal2 22032 2604 22032 2604 0 net81
rlabel metal2 19968 3066 19968 3066 0 net82
rlabel metal2 20976 4200 20976 4200 0 net83
rlabel metal3 22848 2814 22848 2814 0 net84
rlabel metal2 18144 4578 18144 4578 0 net85
rlabel metal2 19488 3612 19488 3612 0 net86
rlabel metal2 21696 4326 21696 4326 0 net87
rlabel metal3 20928 2856 20928 2856 0 net88
rlabel metal2 22368 3150 22368 3150 0 net89
rlabel metal2 37536 9870 37536 9870 0 net9
rlabel metal3 26688 2742 26688 2742 0 net90
rlabel metal2 27456 2016 27456 2016 0 net91
rlabel metal2 26880 4284 26880 4284 0 net92
rlabel metal2 27768 3948 27768 3948 0 net93
rlabel metal2 27840 2604 27840 2604 0 net94
rlabel metal2 28608 1932 28608 1932 0 net95
rlabel metal2 24120 3192 24120 3192 0 net96
rlabel metal2 23880 4704 23880 4704 0 net97
rlabel metal2 24816 3864 24816 3864 0 net98
rlabel metal2 22464 4662 22464 4662 0 net99
<< properties >>
string FIXED_BBOX 0 0 39264 12180
<< end >>
