module S_CPU_IRQ (CONFIGURED_top,
    Co,
    IRQ_top0,
    IRQ_top1,
    IRQ_top2,
    IRQ_top3,
    UserCLK,
    UserCLKo,
    VPWR,
    VGND,
    FrameData,
    FrameData_O,
    FrameStrobe,
    FrameStrobe_O,
    N1BEG,
    N2BEG,
    N2BEGb,
    N4BEG,
    NN4BEG,
    S1END,
    S2END,
    S2MID,
    S4END,
    SS4END);
 input CONFIGURED_top;
 output Co;
 output IRQ_top0;
 output IRQ_top1;
 output IRQ_top2;
 output IRQ_top3;
 input UserCLK;
 output UserCLKo;
 inout VPWR;
 inout VGND;
 input [31:0] FrameData;
 output [31:0] FrameData_O;
 input [19:0] FrameStrobe;
 output [19:0] FrameStrobe_O;
 output [3:0] N1BEG;
 output [7:0] N2BEG;
 output [7:0] N2BEGb;
 output [15:0] N4BEG;
 output [15:0] NN4BEG;
 input [3:0] S1END;
 input [7:0] S2END;
 input [7:0] S2MID;
 input [15:0] S4END;
 input [15:0] SS4END;

 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire \Inst_S_CPU_IRQ_ConfigMem.Inst_frame0_bit20.Q ;
 wire \Inst_S_CPU_IRQ_ConfigMem.Inst_frame0_bit21.Q ;
 wire \Inst_S_CPU_IRQ_ConfigMem.Inst_frame0_bit22.Q ;
 wire \Inst_S_CPU_IRQ_ConfigMem.Inst_frame0_bit23.Q ;
 wire \Inst_S_CPU_IRQ_ConfigMem.Inst_frame0_bit24.Q ;
 wire \Inst_S_CPU_IRQ_ConfigMem.Inst_frame0_bit25.Q ;
 wire \Inst_S_CPU_IRQ_ConfigMem.Inst_frame0_bit26.Q ;
 wire \Inst_S_CPU_IRQ_ConfigMem.Inst_frame0_bit27.Q ;
 wire \Inst_S_CPU_IRQ_ConfigMem.Inst_frame0_bit28.Q ;
 wire \Inst_S_CPU_IRQ_ConfigMem.Inst_frame0_bit29.Q ;
 wire \Inst_S_CPU_IRQ_ConfigMem.Inst_frame0_bit30.Q ;
 wire \Inst_S_CPU_IRQ_ConfigMem.Inst_frame0_bit31.Q ;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire _000_;
 wire _001_;
 wire _002_;
 wire _003_;
 wire _004_;
 wire _005_;
 wire _006_;
 wire _007_;
 wire _008_;
 wire _009_;
 wire _010_;
 wire _011_;
 wire _012_;
 wire _013_;
 wire _014_;
 wire _015_;
 wire _016_;
 wire _017_;
 wire _018_;
 wire _019_;
 wire _020_;
 wire _021_;
 wire _022_;
 wire _023_;
 wire _024_;
 wire _025_;
 wire _026_;
 wire _027_;
 wire _028_;
 wire _029_;
 wire _030_;
 wire _031_;
 wire _032_;
 wire _033_;
 wire _034_;
 wire _035_;
 wire net5;
 wire net6;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net157;

 sg13g2_mux4_1 _036_ (.S0(\Inst_S_CPU_IRQ_ConfigMem.Inst_frame0_bit20.Q ),
    .A0(net16),
    .A1(net28),
    .A2(net20),
    .A3(net24),
    .S1(\Inst_S_CPU_IRQ_ConfigMem.Inst_frame0_bit21.Q ),
    .X(_000_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _037_ (.A(\Inst_S_CPU_IRQ_ConfigMem.Inst_frame0_bit22.Q ),
    .B(_000_),
    .Y(_001_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _038_ (.A(net36),
    .B_N(\Inst_S_CPU_IRQ_ConfigMem.Inst_frame0_bit20.Q ),
    .Y(_002_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _039_ (.A(\Inst_S_CPU_IRQ_ConfigMem.Inst_frame0_bit20.Q ),
    .B(net32),
    .Y(_003_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _040_ (.A(\Inst_S_CPU_IRQ_ConfigMem.Inst_frame0_bit21.Q ),
    .B(_002_),
    .C(_003_),
    .Y(_004_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _041_ (.A(net44),
    .B_N(\Inst_S_CPU_IRQ_ConfigMem.Inst_frame0_bit20.Q ),
    .Y(_005_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _042_ (.B1(\Inst_S_CPU_IRQ_ConfigMem.Inst_frame0_bit21.Q ),
    .VDD(VPWR),
    .Y(_006_),
    .VSS(VGND),
    .A1(\Inst_S_CPU_IRQ_ConfigMem.Inst_frame0_bit20.Q ),
    .A2(net40));
 sg13g2_o21ai_1 _043_ (.B1(\Inst_S_CPU_IRQ_ConfigMem.Inst_frame0_bit22.Q ),
    .VDD(VPWR),
    .Y(_007_),
    .VSS(VGND),
    .A1(_005_),
    .A2(_006_));
 sg13g2_o21ai_1 _044_ (.B1(net1),
    .VDD(VPWR),
    .Y(_008_),
    .VSS(VGND),
    .A1(_004_),
    .A2(_007_));
 sg13g2_nor2_1 _045_ (.A(_001_),
    .B(_008_),
    .Y(net100),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _046_ (.S0(\Inst_S_CPU_IRQ_ConfigMem.Inst_frame0_bit23.Q ),
    .A0(net17),
    .A1(net29),
    .A2(net21),
    .A3(net25),
    .S1(\Inst_S_CPU_IRQ_ConfigMem.Inst_frame0_bit24.Q ),
    .X(_009_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _047_ (.A(\Inst_S_CPU_IRQ_ConfigMem.Inst_frame0_bit25.Q ),
    .B(_009_),
    .Y(_010_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _048_ (.A(net37),
    .B_N(\Inst_S_CPU_IRQ_ConfigMem.Inst_frame0_bit23.Q ),
    .Y(_011_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _049_ (.A(\Inst_S_CPU_IRQ_ConfigMem.Inst_frame0_bit23.Q ),
    .B(net33),
    .Y(_012_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _050_ (.A(\Inst_S_CPU_IRQ_ConfigMem.Inst_frame0_bit24.Q ),
    .B(_011_),
    .C(_012_),
    .Y(_013_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _051_ (.A(net45),
    .B_N(\Inst_S_CPU_IRQ_ConfigMem.Inst_frame0_bit23.Q ),
    .Y(_014_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _052_ (.B1(\Inst_S_CPU_IRQ_ConfigMem.Inst_frame0_bit24.Q ),
    .VDD(VPWR),
    .Y(_015_),
    .VSS(VGND),
    .A1(\Inst_S_CPU_IRQ_ConfigMem.Inst_frame0_bit23.Q ),
    .A2(net41));
 sg13g2_o21ai_1 _053_ (.B1(\Inst_S_CPU_IRQ_ConfigMem.Inst_frame0_bit25.Q ),
    .VDD(VPWR),
    .Y(_016_),
    .VSS(VGND),
    .A1(_014_),
    .A2(_015_));
 sg13g2_o21ai_1 _054_ (.B1(net1),
    .VDD(VPWR),
    .Y(_017_),
    .VSS(VGND),
    .A1(_013_),
    .A2(_016_));
 sg13g2_nor2_1 _055_ (.A(_010_),
    .B(_017_),
    .Y(net101),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _056_ (.S0(\Inst_S_CPU_IRQ_ConfigMem.Inst_frame0_bit26.Q ),
    .A0(net18),
    .A1(net30),
    .A2(net22),
    .A3(net26),
    .S1(\Inst_S_CPU_IRQ_ConfigMem.Inst_frame0_bit27.Q ),
    .X(_018_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _057_ (.A(\Inst_S_CPU_IRQ_ConfigMem.Inst_frame0_bit28.Q ),
    .B(_018_),
    .Y(_019_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _058_ (.A(net38),
    .B_N(\Inst_S_CPU_IRQ_ConfigMem.Inst_frame0_bit26.Q ),
    .Y(_020_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _059_ (.A(\Inst_S_CPU_IRQ_ConfigMem.Inst_frame0_bit26.Q ),
    .B(net34),
    .Y(_021_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _060_ (.A(\Inst_S_CPU_IRQ_ConfigMem.Inst_frame0_bit27.Q ),
    .B(_020_),
    .C(_021_),
    .Y(_022_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _061_ (.A(net46),
    .B_N(\Inst_S_CPU_IRQ_ConfigMem.Inst_frame0_bit26.Q ),
    .Y(_023_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _062_ (.B1(\Inst_S_CPU_IRQ_ConfigMem.Inst_frame0_bit27.Q ),
    .VDD(VPWR),
    .Y(_024_),
    .VSS(VGND),
    .A1(\Inst_S_CPU_IRQ_ConfigMem.Inst_frame0_bit26.Q ),
    .A2(net42));
 sg13g2_o21ai_1 _063_ (.B1(\Inst_S_CPU_IRQ_ConfigMem.Inst_frame0_bit28.Q ),
    .VDD(VPWR),
    .Y(_025_),
    .VSS(VGND),
    .A1(_023_),
    .A2(_024_));
 sg13g2_o21ai_1 _064_ (.B1(net1),
    .VDD(VPWR),
    .Y(_026_),
    .VSS(VGND),
    .A1(_022_),
    .A2(_025_));
 sg13g2_nor2_1 _065_ (.A(_019_),
    .B(_026_),
    .Y(net102),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _066_ (.S0(\Inst_S_CPU_IRQ_ConfigMem.Inst_frame0_bit29.Q ),
    .A0(net19),
    .A1(net31),
    .A2(net23),
    .A3(net27),
    .S1(\Inst_S_CPU_IRQ_ConfigMem.Inst_frame0_bit30.Q ),
    .X(_027_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _067_ (.A(\Inst_S_CPU_IRQ_ConfigMem.Inst_frame0_bit31.Q ),
    .B(_027_),
    .Y(_028_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _068_ (.A(net39),
    .B_N(\Inst_S_CPU_IRQ_ConfigMem.Inst_frame0_bit29.Q ),
    .Y(_029_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _069_ (.A(\Inst_S_CPU_IRQ_ConfigMem.Inst_frame0_bit29.Q ),
    .B(net35),
    .Y(_030_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _070_ (.A(\Inst_S_CPU_IRQ_ConfigMem.Inst_frame0_bit30.Q ),
    .B(_029_),
    .C(_030_),
    .Y(_031_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _071_ (.A(net47),
    .B_N(\Inst_S_CPU_IRQ_ConfigMem.Inst_frame0_bit29.Q ),
    .Y(_032_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _072_ (.B1(\Inst_S_CPU_IRQ_ConfigMem.Inst_frame0_bit30.Q ),
    .VDD(VPWR),
    .Y(_033_),
    .VSS(VGND),
    .A1(\Inst_S_CPU_IRQ_ConfigMem.Inst_frame0_bit29.Q ),
    .A2(net43));
 sg13g2_o21ai_1 _073_ (.B1(\Inst_S_CPU_IRQ_ConfigMem.Inst_frame0_bit31.Q ),
    .VDD(VPWR),
    .Y(_034_),
    .VSS(VGND),
    .A1(_032_),
    .A2(_033_));
 sg13g2_o21ai_1 _074_ (.B1(net1),
    .VDD(VPWR),
    .Y(_035_),
    .VSS(VGND),
    .A1(_031_),
    .A2(_034_));
 sg13g2_nor2_1 _075_ (.A(_028_),
    .B(_035_),
    .Y(net103),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _076_ (.D(net2),
    .GATE(net5),
    .Q(\Inst_S_CPU_IRQ_ConfigMem.Inst_frame0_bit20.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _077_ (.D(net3),
    .GATE(net6),
    .Q(\Inst_S_CPU_IRQ_ConfigMem.Inst_frame0_bit21.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _078_ (.D(net4),
    .GATE(net6),
    .Q(\Inst_S_CPU_IRQ_ConfigMem.Inst_frame0_bit22.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _079_ (.D(net7),
    .GATE(net5),
    .Q(\Inst_S_CPU_IRQ_ConfigMem.Inst_frame0_bit23.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _080_ (.D(net8),
    .GATE(net5),
    .Q(\Inst_S_CPU_IRQ_ConfigMem.Inst_frame0_bit24.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _081_ (.D(net9),
    .GATE(net5),
    .Q(\Inst_S_CPU_IRQ_ConfigMem.Inst_frame0_bit25.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _082_ (.D(net10),
    .GATE(net5),
    .Q(\Inst_S_CPU_IRQ_ConfigMem.Inst_frame0_bit26.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _083_ (.D(net11),
    .GATE(net5),
    .Q(\Inst_S_CPU_IRQ_ConfigMem.Inst_frame0_bit27.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _084_ (.D(net12),
    .GATE(net5),
    .Q(\Inst_S_CPU_IRQ_ConfigMem.Inst_frame0_bit28.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _085_ (.D(net13),
    .GATE(net6),
    .Q(\Inst_S_CPU_IRQ_ConfigMem.Inst_frame0_bit29.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _086_ (.D(net14),
    .GATE(net6),
    .Q(\Inst_S_CPU_IRQ_ConfigMem.Inst_frame0_bit30.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _087_ (.D(net15),
    .GATE(net6),
    .Q(\Inst_S_CPU_IRQ_ConfigMem.Inst_frame0_bit31.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_antennanp ANTENNA_1 (.VDD(VPWR),
    .VSS(VGND),
    .A(FrameData[10]));
 sg13g2_buf_1 _089_ (.A(FrameData[0]),
    .X(net48),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _090_ (.A(FrameData[1]),
    .X(net59),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _091_ (.A(FrameData[2]),
    .X(net70),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _092_ (.A(FrameData[3]),
    .X(net73),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _093_ (.A(FrameData[4]),
    .X(net74),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _094_ (.A(FrameData[5]),
    .X(net75),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _095_ (.A(FrameData[6]),
    .X(net76),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _096_ (.A(FrameData[7]),
    .X(net77),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _097_ (.A(FrameData[8]),
    .X(net78),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _098_ (.A(FrameData[9]),
    .X(net79),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _099_ (.A(FrameData[10]),
    .X(net49),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _100_ (.A(FrameData[11]),
    .X(net50),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _101_ (.A(FrameData[12]),
    .X(net51),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _102_ (.A(FrameData[13]),
    .X(net52),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _103_ (.A(FrameData[14]),
    .X(net53),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _104_ (.A(FrameData[15]),
    .X(net54),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _105_ (.A(FrameData[16]),
    .X(net55),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _106_ (.A(FrameData[17]),
    .X(net56),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _107_ (.A(FrameData[18]),
    .X(net57),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _108_ (.A(FrameData[19]),
    .X(net58),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _109_ (.A(net2),
    .X(net60),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _110_ (.A(net3),
    .X(net61),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _111_ (.A(net4),
    .X(net62),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _112_ (.A(net7),
    .X(net63),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _113_ (.A(net8),
    .X(net64),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _114_ (.A(net9),
    .X(net65),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _115_ (.A(net10),
    .X(net66),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _116_ (.A(net11),
    .X(net67),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _117_ (.A(net12),
    .X(net68),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _118_ (.A(net13),
    .X(net69),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _119_ (.A(net14),
    .X(net71),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _120_ (.A(net15),
    .X(net72),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _121_ (.A(net5),
    .X(net80),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _122_ (.A(FrameStrobe[1]),
    .X(net91),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _123_ (.A(FrameStrobe[2]),
    .X(net92),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _124_ (.A(FrameStrobe[3]),
    .X(net93),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _125_ (.A(FrameStrobe[4]),
    .X(net94),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _126_ (.A(FrameStrobe[5]),
    .X(net95),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _127_ (.A(FrameStrobe[6]),
    .X(net96),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _128_ (.A(FrameStrobe[7]),
    .X(net97),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _129_ (.A(FrameStrobe[8]),
    .X(net98),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _130_ (.A(FrameStrobe[9]),
    .X(net99),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _131_ (.A(FrameStrobe[10]),
    .X(net81),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _132_ (.A(FrameStrobe[11]),
    .X(net82),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _133_ (.A(FrameStrobe[12]),
    .X(net83),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _134_ (.A(FrameStrobe[13]),
    .X(net84),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _135_ (.A(FrameStrobe[14]),
    .X(net85),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _136_ (.A(FrameStrobe[15]),
    .X(net86),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _137_ (.A(FrameStrobe[16]),
    .X(net87),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _138_ (.A(FrameStrobe[17]),
    .X(net88),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _139_ (.A(FrameStrobe[18]),
    .X(net89),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _140_ (.A(FrameStrobe[19]),
    .X(net90),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _141_ (.A(net19),
    .X(net104),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _142_ (.A(net18),
    .X(net105),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _143_ (.A(net17),
    .X(net106),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _144_ (.A(net16),
    .X(net107),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _145_ (.A(S2MID[7]),
    .X(net108),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _146_ (.A(S2MID[6]),
    .X(net109),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _147_ (.A(S2MID[5]),
    .X(net110),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _148_ (.A(S2MID[4]),
    .X(net111),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _149_ (.A(net31),
    .X(net112),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _150_ (.A(net30),
    .X(net113),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _151_ (.A(net29),
    .X(net114),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _152_ (.A(net28),
    .X(net115),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _153_ (.A(net27),
    .X(net116),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _154_ (.A(net26),
    .X(net117),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _155_ (.A(net25),
    .X(net118),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _156_ (.A(net24),
    .X(net119),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _157_ (.A(net23),
    .X(net120),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _158_ (.A(net22),
    .X(net121),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _159_ (.A(net21),
    .X(net122),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _160_ (.A(net20),
    .X(net123),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _161_ (.A(S4END[15]),
    .X(net124),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _162_ (.A(S4END[14]),
    .X(net131),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _163_ (.A(S4END[13]),
    .X(net132),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _164_ (.A(S4END[12]),
    .X(net133),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _165_ (.A(S4END[11]),
    .X(net134),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _166_ (.A(S4END[10]),
    .X(net135),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _167_ (.A(S4END[9]),
    .X(net136),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _168_ (.A(S4END[8]),
    .X(net137),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _169_ (.A(net39),
    .X(net138),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _170_ (.A(net38),
    .X(net139),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _171_ (.A(net37),
    .X(net125),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _172_ (.A(net36),
    .X(net126),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _173_ (.A(net35),
    .X(net127),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _174_ (.A(net34),
    .X(net128),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _175_ (.A(net33),
    .X(net129),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _176_ (.A(net32),
    .X(net130),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _177_ (.A(SS4END[15]),
    .X(net140),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _178_ (.A(SS4END[14]),
    .X(net147),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _179_ (.A(SS4END[13]),
    .X(net148),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _180_ (.A(SS4END[12]),
    .X(net149),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _181_ (.A(SS4END[11]),
    .X(net150),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _182_ (.A(SS4END[10]),
    .X(net151),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _183_ (.A(SS4END[9]),
    .X(net152),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _184_ (.A(SS4END[8]),
    .X(net153),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _185_ (.A(net47),
    .X(net154),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _186_ (.A(net46),
    .X(net155),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _187_ (.A(net45),
    .X(net141),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _188_ (.A(net44),
    .X(net142),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _189_ (.A(net43),
    .X(net143),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _190_ (.A(net42),
    .X(net144),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _191_ (.A(net41),
    .X(net145),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _192_ (.A(net40),
    .X(net146),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _193_ (.A(UserCLK),
    .X(net156),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout5 (.A(FrameStrobe[0]),
    .X(net5),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout6 (.A(FrameStrobe[0]),
    .X(net6),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input1 (.A(CONFIGURED_top),
    .X(net1),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input2 (.A(FrameData[20]),
    .X(net2),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input3 (.A(FrameData[21]),
    .X(net3),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input4 (.A(FrameData[22]),
    .X(net4),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input5 (.A(FrameData[23]),
    .X(net7),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input6 (.A(FrameData[24]),
    .X(net8),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input7 (.A(FrameData[25]),
    .X(net9),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input8 (.A(FrameData[26]),
    .X(net10),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input9 (.A(FrameData[27]),
    .X(net11),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input10 (.A(FrameData[28]),
    .X(net12),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input11 (.A(FrameData[29]),
    .X(net13),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input12 (.A(FrameData[30]),
    .X(net14),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input13 (.A(FrameData[31]),
    .X(net15),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input14 (.A(S1END[0]),
    .X(net16),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input15 (.A(S1END[1]),
    .X(net17),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input16 (.A(S1END[2]),
    .X(net18),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input17 (.A(S1END[3]),
    .X(net19),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input18 (.A(S2END[0]),
    .X(net20),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input19 (.A(S2END[1]),
    .X(net21),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input20 (.A(S2END[2]),
    .X(net22),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input21 (.A(S2END[3]),
    .X(net23),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input22 (.A(S2END[4]),
    .X(net24),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input23 (.A(S2END[5]),
    .X(net25),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input24 (.A(S2END[6]),
    .X(net26),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input25 (.A(S2END[7]),
    .X(net27),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input26 (.A(S2MID[0]),
    .X(net28),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input27 (.A(S2MID[1]),
    .X(net29),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input28 (.A(S2MID[2]),
    .X(net30),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input29 (.A(S2MID[3]),
    .X(net31),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input30 (.A(S4END[0]),
    .X(net32),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input31 (.A(S4END[1]),
    .X(net33),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input32 (.A(S4END[2]),
    .X(net34),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input33 (.A(S4END[3]),
    .X(net35),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input34 (.A(S4END[4]),
    .X(net36),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input35 (.A(S4END[5]),
    .X(net37),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input36 (.A(S4END[6]),
    .X(net38),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input37 (.A(S4END[7]),
    .X(net39),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input38 (.A(SS4END[0]),
    .X(net40),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input39 (.A(SS4END[1]),
    .X(net41),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input40 (.A(SS4END[2]),
    .X(net42),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input41 (.A(SS4END[3]),
    .X(net43),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input42 (.A(SS4END[4]),
    .X(net44),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input43 (.A(SS4END[5]),
    .X(net45),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input44 (.A(SS4END[6]),
    .X(net46),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input45 (.A(SS4END[7]),
    .X(net47),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output46 (.A(net48),
    .X(FrameData_O[0]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output47 (.A(net49),
    .X(FrameData_O[10]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output48 (.A(net50),
    .X(FrameData_O[11]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output49 (.A(net51),
    .X(FrameData_O[12]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output50 (.A(net52),
    .X(FrameData_O[13]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output51 (.A(net53),
    .X(FrameData_O[14]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output52 (.A(net54),
    .X(FrameData_O[15]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output53 (.A(net55),
    .X(FrameData_O[16]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output54 (.A(net56),
    .X(FrameData_O[17]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output55 (.A(net57),
    .X(FrameData_O[18]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output56 (.A(net58),
    .X(FrameData_O[19]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output57 (.A(net59),
    .X(FrameData_O[1]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output58 (.A(net60),
    .X(FrameData_O[20]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output59 (.A(net61),
    .X(FrameData_O[21]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output60 (.A(net62),
    .X(FrameData_O[22]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output61 (.A(net63),
    .X(FrameData_O[23]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output62 (.A(net64),
    .X(FrameData_O[24]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output63 (.A(net65),
    .X(FrameData_O[25]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output64 (.A(net66),
    .X(FrameData_O[26]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output65 (.A(net67),
    .X(FrameData_O[27]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output66 (.A(net68),
    .X(FrameData_O[28]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output67 (.A(net69),
    .X(FrameData_O[29]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output68 (.A(net70),
    .X(FrameData_O[2]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output69 (.A(net71),
    .X(FrameData_O[30]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output70 (.A(net72),
    .X(FrameData_O[31]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output71 (.A(net73),
    .X(FrameData_O[3]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output72 (.A(net74),
    .X(FrameData_O[4]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output73 (.A(net75),
    .X(FrameData_O[5]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output74 (.A(net76),
    .X(FrameData_O[6]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output75 (.A(net77),
    .X(FrameData_O[7]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output76 (.A(net78),
    .X(FrameData_O[8]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output77 (.A(net79),
    .X(FrameData_O[9]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output78 (.A(net80),
    .X(FrameStrobe_O[0]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output79 (.A(net81),
    .X(FrameStrobe_O[10]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output80 (.A(net82),
    .X(FrameStrobe_O[11]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output81 (.A(net83),
    .X(FrameStrobe_O[12]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output82 (.A(net84),
    .X(FrameStrobe_O[13]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output83 (.A(net85),
    .X(FrameStrobe_O[14]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output84 (.A(net86),
    .X(FrameStrobe_O[15]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output85 (.A(net87),
    .X(FrameStrobe_O[16]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output86 (.A(net88),
    .X(FrameStrobe_O[17]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output87 (.A(net89),
    .X(FrameStrobe_O[18]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output88 (.A(net90),
    .X(FrameStrobe_O[19]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output89 (.A(net91),
    .X(FrameStrobe_O[1]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output90 (.A(net92),
    .X(FrameStrobe_O[2]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output91 (.A(net93),
    .X(FrameStrobe_O[3]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output92 (.A(net94),
    .X(FrameStrobe_O[4]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output93 (.A(net95),
    .X(FrameStrobe_O[5]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output94 (.A(net96),
    .X(FrameStrobe_O[6]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output95 (.A(net97),
    .X(FrameStrobe_O[7]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output96 (.A(net98),
    .X(FrameStrobe_O[8]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output97 (.A(net99),
    .X(FrameStrobe_O[9]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output98 (.A(net100),
    .X(IRQ_top0),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output99 (.A(net101),
    .X(IRQ_top1),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output100 (.A(net102),
    .X(IRQ_top2),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output101 (.A(net103),
    .X(IRQ_top3),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output102 (.A(net104),
    .X(N1BEG[0]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output103 (.A(net105),
    .X(N1BEG[1]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output104 (.A(net106),
    .X(N1BEG[2]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output105 (.A(net107),
    .X(N1BEG[3]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output106 (.A(net108),
    .X(N2BEG[0]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output107 (.A(net109),
    .X(N2BEG[1]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output108 (.A(net110),
    .X(N2BEG[2]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output109 (.A(net111),
    .X(N2BEG[3]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output110 (.A(net112),
    .X(N2BEG[4]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output111 (.A(net113),
    .X(N2BEG[5]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output112 (.A(net114),
    .X(N2BEG[6]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output113 (.A(net115),
    .X(N2BEG[7]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output114 (.A(net116),
    .X(N2BEGb[0]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output115 (.A(net117),
    .X(N2BEGb[1]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output116 (.A(net118),
    .X(N2BEGb[2]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output117 (.A(net119),
    .X(N2BEGb[3]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output118 (.A(net120),
    .X(N2BEGb[4]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output119 (.A(net121),
    .X(N2BEGb[5]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output120 (.A(net122),
    .X(N2BEGb[6]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output121 (.A(net123),
    .X(N2BEGb[7]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output122 (.A(net124),
    .X(N4BEG[0]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output123 (.A(net125),
    .X(N4BEG[10]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output124 (.A(net126),
    .X(N4BEG[11]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output125 (.A(net127),
    .X(N4BEG[12]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output126 (.A(net128),
    .X(N4BEG[13]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output127 (.A(net129),
    .X(N4BEG[14]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output128 (.A(net130),
    .X(N4BEG[15]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output129 (.A(net131),
    .X(N4BEG[1]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output130 (.A(net132),
    .X(N4BEG[2]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output131 (.A(net133),
    .X(N4BEG[3]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output132 (.A(net134),
    .X(N4BEG[4]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output133 (.A(net135),
    .X(N4BEG[5]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output134 (.A(net136),
    .X(N4BEG[6]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output135 (.A(net137),
    .X(N4BEG[7]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output136 (.A(net138),
    .X(N4BEG[8]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output137 (.A(net139),
    .X(N4BEG[9]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output138 (.A(net140),
    .X(NN4BEG[0]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output139 (.A(net141),
    .X(NN4BEG[10]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output140 (.A(net142),
    .X(NN4BEG[11]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output141 (.A(net143),
    .X(NN4BEG[12]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output142 (.A(net144),
    .X(NN4BEG[13]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output143 (.A(net145),
    .X(NN4BEG[14]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output144 (.A(net146),
    .X(NN4BEG[15]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output145 (.A(net147),
    .X(NN4BEG[1]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output146 (.A(net148),
    .X(NN4BEG[2]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output147 (.A(net149),
    .X(NN4BEG[3]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output148 (.A(net150),
    .X(NN4BEG[4]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output149 (.A(net151),
    .X(NN4BEG[5]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output150 (.A(net152),
    .X(NN4BEG[6]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output151 (.A(net153),
    .X(NN4BEG[7]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output152 (.A(net154),
    .X(NN4BEG[8]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output153 (.A(net155),
    .X(NN4BEG[9]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output154 (.A(net156),
    .X(UserCLKo),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_tielo S_CPU_IRQ_155 (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(net157));
 sg13g2_antennanp ANTENNA_2 (.VDD(VPWR),
    .VSS(VGND),
    .A(FrameData[11]));
 sg13g2_antennanp ANTENNA_3 (.VDD(VPWR),
    .VSS(VGND),
    .A(FrameData[18]));
 sg13g2_antennanp ANTENNA_4 (.VDD(VPWR),
    .VSS(VGND),
    .A(FrameData[8]));
 sg13g2_antennanp ANTENNA_5 (.VDD(VPWR),
    .VSS(VGND),
    .A(net63));
 sg13g2_antennanp ANTENNA_6 (.VDD(VPWR),
    .VSS(VGND),
    .A(net64));
 sg13g2_antennanp ANTENNA_7 (.VDD(VPWR),
    .VSS(VGND),
    .A(FrameData[10]));
 sg13g2_antennanp ANTENNA_8 (.VDD(VPWR),
    .VSS(VGND),
    .A(FrameData[11]));
 sg13g2_antennanp ANTENNA_9 (.VDD(VPWR),
    .VSS(VGND),
    .A(FrameData[18]));
 sg13g2_antennanp ANTENNA_10 (.VDD(VPWR),
    .VSS(VGND),
    .A(FrameData[8]));
 sg13g2_antennanp ANTENNA_11 (.VDD(VPWR),
    .VSS(VGND),
    .A(net63));
 sg13g2_antennanp ANTENNA_12 (.VDD(VPWR),
    .VSS(VGND),
    .A(net64));
 sg13g2_antennanp ANTENNA_13 (.VDD(VPWR),
    .VSS(VGND),
    .A(FrameData[10]));
 sg13g2_antennanp ANTENNA_14 (.VDD(VPWR),
    .VSS(VGND),
    .A(FrameData[11]));
 sg13g2_antennanp ANTENNA_15 (.VDD(VPWR),
    .VSS(VGND),
    .A(FrameData[18]));
 sg13g2_antennanp ANTENNA_16 (.VDD(VPWR),
    .VSS(VGND),
    .A(FrameData[8]));
 sg13g2_antennanp ANTENNA_17 (.VDD(VPWR),
    .VSS(VGND),
    .A(net63));
 sg13g2_antennanp ANTENNA_18 (.VDD(VPWR),
    .VSS(VGND),
    .A(net64));
 sg13g2_antennanp ANTENNA_19 (.VDD(VPWR),
    .VSS(VGND),
    .A(FrameData[10]));
 sg13g2_antennanp ANTENNA_20 (.VDD(VPWR),
    .VSS(VGND),
    .A(FrameData[11]));
 sg13g2_antennanp ANTENNA_21 (.VDD(VPWR),
    .VSS(VGND),
    .A(FrameData[18]));
 sg13g2_antennanp ANTENNA_22 (.VDD(VPWR),
    .VSS(VGND),
    .A(FrameData[8]));
 sg13g2_antennanp ANTENNA_23 (.VDD(VPWR),
    .VSS(VGND),
    .A(net63));
 sg13g2_antennanp ANTENNA_24 (.VDD(VPWR),
    .VSS(VGND),
    .A(net64));
 sg13g2_antennanp ANTENNA_25 (.VDD(VPWR),
    .VSS(VGND),
    .A(FrameData[10]));
 sg13g2_antennanp ANTENNA_26 (.VDD(VPWR),
    .VSS(VGND),
    .A(FrameData[11]));
 sg13g2_antennanp ANTENNA_27 (.VDD(VPWR),
    .VSS(VGND),
    .A(FrameData[8]));
 sg13g2_antennanp ANTENNA_28 (.VDD(VPWR),
    .VSS(VGND),
    .A(net63));
 sg13g2_antennanp ANTENNA_29 (.VDD(VPWR),
    .VSS(VGND),
    .A(net64));
 sg13g2_antennanp ANTENNA_30 (.VDD(VPWR),
    .VSS(VGND),
    .A(FrameData[10]));
 sg13g2_antennanp ANTENNA_31 (.VDD(VPWR),
    .VSS(VGND),
    .A(FrameData[11]));
 sg13g2_antennanp ANTENNA_32 (.VDD(VPWR),
    .VSS(VGND),
    .A(FrameData[8]));
 sg13g2_antennanp ANTENNA_33 (.VDD(VPWR),
    .VSS(VGND),
    .A(net63));
 sg13g2_antennanp ANTENNA_34 (.VDD(VPWR),
    .VSS(VGND),
    .A(net64));
 sg13g2_antennanp ANTENNA_35 (.VDD(VPWR),
    .VSS(VGND),
    .A(FrameData[10]));
 sg13g2_antennanp ANTENNA_36 (.VDD(VPWR),
    .VSS(VGND),
    .A(FrameData[11]));
 sg13g2_antennanp ANTENNA_37 (.VDD(VPWR),
    .VSS(VGND),
    .A(FrameData[8]));
 sg13g2_antennanp ANTENNA_38 (.VDD(VPWR),
    .VSS(VGND),
    .A(net63));
 sg13g2_antennanp ANTENNA_39 (.VDD(VPWR),
    .VSS(VGND),
    .A(net64));
 sg13g2_antennanp ANTENNA_40 (.VDD(VPWR),
    .VSS(VGND),
    .A(FrameData[10]));
 sg13g2_antennanp ANTENNA_41 (.VDD(VPWR),
    .VSS(VGND),
    .A(FrameData[11]));
 sg13g2_antennanp ANTENNA_42 (.VDD(VPWR),
    .VSS(VGND),
    .A(FrameData[8]));
 sg13g2_antennanp ANTENNA_43 (.VDD(VPWR),
    .VSS(VGND),
    .A(net63));
 sg13g2_antennanp ANTENNA_44 (.VDD(VPWR),
    .VSS(VGND),
    .A(net64));
 sg13g2_antennanp ANTENNA_45 (.VDD(VPWR),
    .VSS(VGND),
    .A(FrameData[10]));
 sg13g2_antennanp ANTENNA_46 (.VDD(VPWR),
    .VSS(VGND),
    .A(FrameData[11]));
 sg13g2_antennanp ANTENNA_47 (.VDD(VPWR),
    .VSS(VGND),
    .A(FrameData[8]));
 sg13g2_antennanp ANTENNA_48 (.VDD(VPWR),
    .VSS(VGND),
    .A(net63));
 sg13g2_antennanp ANTENNA_49 (.VDD(VPWR),
    .VSS(VGND),
    .A(net64));
 sg13g2_antennanp ANTENNA_50 (.VDD(VPWR),
    .VSS(VGND),
    .A(FrameData[10]));
 sg13g2_antennanp ANTENNA_51 (.VDD(VPWR),
    .VSS(VGND),
    .A(FrameData[11]));
 sg13g2_antennanp ANTENNA_52 (.VDD(VPWR),
    .VSS(VGND),
    .A(FrameData[8]));
 sg13g2_antennanp ANTENNA_53 (.VDD(VPWR),
    .VSS(VGND),
    .A(net63));
 sg13g2_antennanp ANTENNA_54 (.VDD(VPWR),
    .VSS(VGND),
    .A(net64));
 sg13g2_fill_2 FILLER_0_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_0_2 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_25 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_32 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_43 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_50 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_61 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_68 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_79 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_86 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_93 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_100 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_107 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_114 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_121 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_128 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_135 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_142 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_149 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_156 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_163 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_170 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_177 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_184 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_191 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_198 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_205 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_212 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_219 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_226 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_233 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_240 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_247 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_254 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_261 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_268 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_275 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_282 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_289 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_296 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_303 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_310 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_317 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_324 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_331 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_338 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_345 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_352 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_359 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_366 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_373 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_380 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_387 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_394 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_401 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_408 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_415 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_422 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_429 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_0_436 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_0_438 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_63 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_70 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_1_77 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_1_81 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_99 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_106 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_1_117 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_1_123 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_1_127 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_1_137 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_1_142 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_147 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_154 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_161 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_168 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_175 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_182 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_189 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_196 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_203 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_210 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_1_217 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_1_219 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_241 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_248 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_255 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_262 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_269 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_276 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_283 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_290 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_297 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_304 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_311 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_318 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_325 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_332 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_339 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_346 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_353 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_360 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_367 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_374 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_381 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_1_388 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_1_392 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_1_401 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_1_403 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_1_425 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_434 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_1_441 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_1_445 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_63 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_70 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_2_77 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_2_82 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_2_84 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_2_106 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_2_138 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_2_145 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_2_150 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_173 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_180 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_187 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_194 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_201 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_2_208 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_2_251 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_2_253 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_275 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_282 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_289 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_296 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_303 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_310 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_317 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_324 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_331 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_338 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_345 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_352 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_359 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_366 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_373 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_2_380 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_2_390 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_2_395 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_2_397 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_2_415 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_2_417 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_438 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_2_445 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_2_449 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_63 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_70 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_77 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_84 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_91 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_98 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_3_105 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_3_109 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_133 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_3_140 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_3_144 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_150 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_157 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_3_164 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_3_172 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_190 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_197 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_204 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_211 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_3_218 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_247 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_254 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_261 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_268 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_3_275 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_280 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_287 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_294 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_301 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_308 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_315 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_322 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_3_329 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_3_333 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_338 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_345 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_352 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_359 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_366 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_373 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_380 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_391 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_398 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_3_405 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_419 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_430 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_437 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_444 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_63 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_70 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_77 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_84 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_91 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_98 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_105 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_112 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_4_119 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_125 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_132 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_139 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_146 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_153 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_160 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_167 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_174 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_181 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_188 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_195 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_4_202 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_4_225 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_4_229 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_234 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_241 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_248 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_255 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_262 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_4_269 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_4_273 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_292 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_299 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_306 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_313 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_320 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_327 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_334 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_341 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_360 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_367 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_374 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_381 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_388 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_395 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_402 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_409 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_416 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_423 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_430 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_437 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_444 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_63 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_70 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_77 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_84 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_91 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_98 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_105 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_112 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_119 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_126 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_133 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_140 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_147 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_154 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_161 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_168 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_175 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_182 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_189 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_196 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_203 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_210 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_217 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_224 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_231 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_238 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_245 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_252 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_259 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_266 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_273 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_280 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_287 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_294 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_301 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_308 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_315 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_322 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_329 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_336 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_5_343 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_5_347 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_352 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_359 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_366 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_373 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_380 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_387 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_394 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_401 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_408 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_415 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_422 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_429 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_5_436 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_5_450 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_63 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_70 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_77 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_84 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_91 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_98 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_105 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_112 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_119 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_126 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_133 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_140 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_147 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_154 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_161 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_168 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_175 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_182 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_189 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_196 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_203 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_210 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_217 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_224 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_231 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_238 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_245 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_252 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_6_259 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_277 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_6_284 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_6_286 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_6_292 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_302 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_6_309 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_314 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_321 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_328 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_335 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_6_342 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_6_346 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_6_352 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_6_354 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_363 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_6_370 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_6_372 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_377 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_384 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_391 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_398 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_405 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_412 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_6_419 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_425 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_432 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_6_439 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_6_450 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_7_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_31 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_38 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_45 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_52 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_59 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_66 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_73 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_80 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_87 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_94 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_101 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_125 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_132 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_7_139 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_7_143 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_7_148 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_7_158 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_7_160 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_7_166 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_178 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_185 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_192 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_199 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_206 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_7_217 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_222 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_229 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_236 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_243 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_7_250 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_7_252 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_274 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_7_281 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_7_283 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_324 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_331 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_338 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_345 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_7_352 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_7_356 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_361 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_368 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_375 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_7_382 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_7_393 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_7_407 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_415 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_422 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_7_429 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_7_431 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_7_447 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_8 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_15 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_22 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_29 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_36 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_43 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_50 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_57 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_64 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_71 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_78 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_85 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_92 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_8_99 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_8_109 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_8_131 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_185 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_213 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_220 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_227 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_234 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_241 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_248 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_8_255 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_8_257 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_262 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_269 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_276 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_8_283 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_8_307 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_8_311 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_325 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_332 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_339 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_8_346 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_360 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_367 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_8_374 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_8_391 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_8_397 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_8_401 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_410 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_417 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_8_424 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_8_454 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_9_16 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_26 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_33 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_40 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_47 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_54 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_61 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_68 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_75 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_82 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_9_89 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_9_91 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_9_148 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_9_162 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_9_164 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_9_169 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_9_179 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_9_212 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_9_221 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_237 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_244 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_267 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_274 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_281 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_9_288 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_9_290 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_9_295 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_300 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_307 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_314 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_9_321 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_9_351 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_361 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_368 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_375 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_9_382 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_24 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_31 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_38 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_45 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_52 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_59 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_66 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_73 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_10_80 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_10_84 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_273 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_10_280 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_10_309 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_369 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_376 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_383 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_390 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_397 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_10_404 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_10_451 (.VDD(VPWR),
    .VSS(VGND));
 assign Co = net157;
endmodule
