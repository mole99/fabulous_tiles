module S_WARMBOOT (BOOT_top,
    Co,
    RESET_top,
    SLOT_top0,
    SLOT_top1,
    SLOT_top2,
    SLOT_top3,
    UserCLK,
    UserCLKo,
    FrameData,
    FrameData_O,
    FrameStrobe,
    FrameStrobe_O,
    N1BEG,
    N2BEG,
    N2BEGb,
    N4BEG,
    NN4BEG,
    S1END,
    S2END,
    S2MID,
    S4END,
    SS4END);
 output BOOT_top;
 output Co;
 input RESET_top;
 output SLOT_top0;
 output SLOT_top1;
 output SLOT_top2;
 output SLOT_top3;
 input UserCLK;
 output UserCLKo;
 input [31:0] FrameData;
 output [31:0] FrameData_O;
 input [19:0] FrameStrobe;
 output [19:0] FrameStrobe_O;
 output [3:0] N1BEG;
 output [7:0] N2BEG;
 output [7:0] N2BEGb;
 output [15:0] N4BEG;
 output [15:0] NN4BEG;
 input [3:0] S1END;
 input [7:0] S2END;
 input [7:0] S2MID;
 input [15:0] S4END;
 input [15:0] SS4END;

 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire \Inst_S_WARMBOOT_ConfigMem.Inst_frame0_bit13.Q ;
 wire \Inst_S_WARMBOOT_ConfigMem.Inst_frame0_bit14.Q ;
 wire \Inst_S_WARMBOOT_ConfigMem.Inst_frame0_bit15.Q ;
 wire \Inst_S_WARMBOOT_ConfigMem.Inst_frame0_bit16.Q ;
 wire \Inst_S_WARMBOOT_ConfigMem.Inst_frame0_bit17.Q ;
 wire \Inst_S_WARMBOOT_ConfigMem.Inst_frame0_bit18.Q ;
 wire \Inst_S_WARMBOOT_ConfigMem.Inst_frame0_bit19.Q ;
 wire \Inst_S_WARMBOOT_ConfigMem.Inst_frame0_bit20.Q ;
 wire \Inst_S_WARMBOOT_ConfigMem.Inst_frame0_bit21.Q ;
 wire \Inst_S_WARMBOOT_ConfigMem.Inst_frame0_bit22.Q ;
 wire \Inst_S_WARMBOOT_ConfigMem.Inst_frame0_bit23.Q ;
 wire \Inst_S_WARMBOOT_ConfigMem.Inst_frame0_bit24.Q ;
 wire \Inst_S_WARMBOOT_ConfigMem.Inst_frame0_bit25.Q ;
 wire \Inst_S_WARMBOOT_ConfigMem.Inst_frame0_bit26.Q ;
 wire \Inst_S_WARMBOOT_ConfigMem.Inst_frame0_bit27.Q ;
 wire \Inst_S_WARMBOOT_ConfigMem.Inst_frame0_bit28.Q ;
 wire \Inst_S_WARMBOOT_ConfigMem.Inst_frame0_bit29.Q ;
 wire \Inst_S_WARMBOOT_ConfigMem.Inst_frame0_bit30.Q ;
 wire \Inst_S_WARMBOOT_ConfigMem.Inst_frame0_bit31.Q ;
 wire \Inst_S_WARMBOOT_switch_matrix.N1BEG0 ;
 wire \Inst_S_WARMBOOT_switch_matrix.N1BEG1 ;
 wire \Inst_S_WARMBOOT_switch_matrix.N1BEG2 ;
 wire \Inst_S_WARMBOOT_switch_matrix.N1BEG3 ;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire _000_;
 wire _001_;
 wire _002_;
 wire _003_;
 wire _004_;
 wire _005_;
 wire _006_;
 wire _007_;
 wire _008_;
 wire _009_;
 wire _010_;
 wire _011_;
 wire _012_;
 wire _013_;
 wire _014_;
 wire _015_;
 wire _016_;
 wire _017_;
 wire _018_;
 wire _019_;
 wire _020_;
 wire _021_;
 wire _022_;
 wire _023_;
 wire _024_;
 wire _025_;
 wire _026_;
 wire _027_;
 wire _028_;
 wire _029_;
 wire net7;
 wire net8;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net166;

 sky130_fd_sc_hd__inv_1 _030_ (.A(\Inst_S_WARMBOOT_ConfigMem.Inst_frame0_bit31.Q ),
    .Y(_000_));
 sky130_fd_sc_hd__inv_2 _031_ (.A(\Inst_S_WARMBOOT_ConfigMem.Inst_frame0_bit28.Q ),
    .Y(_001_));
 sky130_fd_sc_hd__inv_2 _032_ (.A(\Inst_S_WARMBOOT_ConfigMem.Inst_frame0_bit25.Q ),
    .Y(_002_));
 sky130_fd_sc_hd__inv_2 _033_ (.A(\Inst_S_WARMBOOT_ConfigMem.Inst_frame0_bit22.Q ),
    .Y(_003_));
 sky130_fd_sc_hd__inv_1 _034_ (.A(\Inst_S_WARMBOOT_ConfigMem.Inst_frame0_bit19.Q ),
    .Y(_004_));
 sky130_fd_sc_hd__mux4_1 _035_ (.A0(net43),
    .A1(net47),
    .A2(net51),
    .A3(net55),
    .S0(\Inst_S_WARMBOOT_ConfigMem.Inst_frame0_bit29.Q ),
    .S1(\Inst_S_WARMBOOT_ConfigMem.Inst_frame0_bit30.Q ),
    .X(_005_));
 sky130_fd_sc_hd__nand2b_1 _036_ (.A_N(net39),
    .B(\Inst_S_WARMBOOT_ConfigMem.Inst_frame0_bit29.Q ),
    .Y(_006_));
 sky130_fd_sc_hd__o21ba_1 _037_ (.A1(net27),
    .A2(\Inst_S_WARMBOOT_ConfigMem.Inst_frame0_bit29.Q ),
    .B1_N(\Inst_S_WARMBOOT_ConfigMem.Inst_frame0_bit30.Q ),
    .X(_007_));
 sky130_fd_sc_hd__mux2_1 _038_ (.A0(net31),
    .A1(net35),
    .S(\Inst_S_WARMBOOT_ConfigMem.Inst_frame0_bit29.Q ),
    .X(_008_));
 sky130_fd_sc_hd__a221o_1 _039_ (.A1(_006_),
    .A2(_007_),
    .B1(_008_),
    .B2(\Inst_S_WARMBOOT_ConfigMem.Inst_frame0_bit30.Q ),
    .C1(\Inst_S_WARMBOOT_ConfigMem.Inst_frame0_bit31.Q ),
    .X(_009_));
 sky130_fd_sc_hd__o21a_1 _040_ (.A1(_000_),
    .A2(_005_),
    .B1(_009_),
    .X(net164));
 sky130_fd_sc_hd__mux4_1 _041_ (.A0(net42),
    .A1(net46),
    .A2(net50),
    .A3(net54),
    .S0(\Inst_S_WARMBOOT_ConfigMem.Inst_frame0_bit26.Q ),
    .S1(\Inst_S_WARMBOOT_ConfigMem.Inst_frame0_bit27.Q ),
    .X(_010_));
 sky130_fd_sc_hd__nand2b_1 _042_ (.A_N(net38),
    .B(\Inst_S_WARMBOOT_ConfigMem.Inst_frame0_bit26.Q ),
    .Y(_011_));
 sky130_fd_sc_hd__o21ba_1 _043_ (.A1(net26),
    .A2(\Inst_S_WARMBOOT_ConfigMem.Inst_frame0_bit26.Q ),
    .B1_N(\Inst_S_WARMBOOT_ConfigMem.Inst_frame0_bit27.Q ),
    .X(_012_));
 sky130_fd_sc_hd__mux2_1 _044_ (.A0(net30),
    .A1(net34),
    .S(\Inst_S_WARMBOOT_ConfigMem.Inst_frame0_bit26.Q ),
    .X(_013_));
 sky130_fd_sc_hd__a221o_1 _045_ (.A1(_011_),
    .A2(_012_),
    .B1(_013_),
    .B2(\Inst_S_WARMBOOT_ConfigMem.Inst_frame0_bit27.Q ),
    .C1(\Inst_S_WARMBOOT_ConfigMem.Inst_frame0_bit28.Q ),
    .X(_014_));
 sky130_fd_sc_hd__o21a_1 _046_ (.A1(_001_),
    .A2(_010_),
    .B1(_014_),
    .X(net163));
 sky130_fd_sc_hd__mux4_1 _047_ (.A0(net41),
    .A1(net45),
    .A2(net49),
    .A3(net53),
    .S0(\Inst_S_WARMBOOT_ConfigMem.Inst_frame0_bit23.Q ),
    .S1(\Inst_S_WARMBOOT_ConfigMem.Inst_frame0_bit24.Q ),
    .X(_015_));
 sky130_fd_sc_hd__nand2b_1 _048_ (.A_N(net37),
    .B(\Inst_S_WARMBOOT_ConfigMem.Inst_frame0_bit23.Q ),
    .Y(_016_));
 sky130_fd_sc_hd__o21ba_1 _049_ (.A1(net25),
    .A2(\Inst_S_WARMBOOT_ConfigMem.Inst_frame0_bit23.Q ),
    .B1_N(\Inst_S_WARMBOOT_ConfigMem.Inst_frame0_bit24.Q ),
    .X(_017_));
 sky130_fd_sc_hd__mux2_1 _050_ (.A0(net29),
    .A1(net33),
    .S(\Inst_S_WARMBOOT_ConfigMem.Inst_frame0_bit23.Q ),
    .X(_018_));
 sky130_fd_sc_hd__a221o_1 _051_ (.A1(_016_),
    .A2(_017_),
    .B1(_018_),
    .B2(\Inst_S_WARMBOOT_ConfigMem.Inst_frame0_bit24.Q ),
    .C1(\Inst_S_WARMBOOT_ConfigMem.Inst_frame0_bit25.Q ),
    .X(_019_));
 sky130_fd_sc_hd__o21a_1 _052_ (.A1(_002_),
    .A2(_015_),
    .B1(_019_),
    .X(net162));
 sky130_fd_sc_hd__mux4_1 _053_ (.A0(net40),
    .A1(net44),
    .A2(net48),
    .A3(net52),
    .S0(\Inst_S_WARMBOOT_ConfigMem.Inst_frame0_bit20.Q ),
    .S1(\Inst_S_WARMBOOT_ConfigMem.Inst_frame0_bit21.Q ),
    .X(_020_));
 sky130_fd_sc_hd__nand2b_1 _054_ (.A_N(net36),
    .B(\Inst_S_WARMBOOT_ConfigMem.Inst_frame0_bit20.Q ),
    .Y(_021_));
 sky130_fd_sc_hd__o21ba_1 _055_ (.A1(net24),
    .A2(\Inst_S_WARMBOOT_ConfigMem.Inst_frame0_bit20.Q ),
    .B1_N(\Inst_S_WARMBOOT_ConfigMem.Inst_frame0_bit21.Q ),
    .X(_022_));
 sky130_fd_sc_hd__mux2_1 _056_ (.A0(net28),
    .A1(net32),
    .S(\Inst_S_WARMBOOT_ConfigMem.Inst_frame0_bit20.Q ),
    .X(_023_));
 sky130_fd_sc_hd__a221o_1 _057_ (.A1(_021_),
    .A2(_022_),
    .B1(_023_),
    .B2(\Inst_S_WARMBOOT_ConfigMem.Inst_frame0_bit21.Q ),
    .C1(\Inst_S_WARMBOOT_ConfigMem.Inst_frame0_bit22.Q ),
    .X(_024_));
 sky130_fd_sc_hd__o21a_1 _058_ (.A1(_003_),
    .A2(_020_),
    .B1(_024_),
    .X(net161));
 sky130_fd_sc_hd__mux4_1 _059_ (.A0(net43),
    .A1(net47),
    .A2(net51),
    .A3(net55),
    .S0(\Inst_S_WARMBOOT_ConfigMem.Inst_frame0_bit17.Q ),
    .S1(\Inst_S_WARMBOOT_ConfigMem.Inst_frame0_bit18.Q ),
    .X(_025_));
 sky130_fd_sc_hd__nand2b_1 _060_ (.A_N(net39),
    .B(\Inst_S_WARMBOOT_ConfigMem.Inst_frame0_bit17.Q ),
    .Y(_026_));
 sky130_fd_sc_hd__o21ba_1 _061_ (.A1(net27),
    .A2(\Inst_S_WARMBOOT_ConfigMem.Inst_frame0_bit17.Q ),
    .B1_N(\Inst_S_WARMBOOT_ConfigMem.Inst_frame0_bit18.Q ),
    .X(_027_));
 sky130_fd_sc_hd__mux2_1 _062_ (.A0(net31),
    .A1(net35),
    .S(\Inst_S_WARMBOOT_ConfigMem.Inst_frame0_bit17.Q ),
    .X(_028_));
 sky130_fd_sc_hd__a221o_1 _063_ (.A1(_026_),
    .A2(_027_),
    .B1(_028_),
    .B2(\Inst_S_WARMBOOT_ConfigMem.Inst_frame0_bit18.Q ),
    .C1(\Inst_S_WARMBOOT_ConfigMem.Inst_frame0_bit19.Q ),
    .X(_029_));
 sky130_fd_sc_hd__o21a_1 _064_ (.A1(_004_),
    .A2(_025_),
    .B1(_029_),
    .X(net56));
 sky130_fd_sc_hd__mux2_1 _065_ (.A0(net24),
    .A1(net23),
    .S(\Inst_S_WARMBOOT_ConfigMem.Inst_frame0_bit16.Q ),
    .X(\Inst_S_WARMBOOT_switch_matrix.N1BEG3 ));
 sky130_fd_sc_hd__mux2_1 _066_ (.A0(net25),
    .A1(net23),
    .S(\Inst_S_WARMBOOT_ConfigMem.Inst_frame0_bit15.Q ),
    .X(\Inst_S_WARMBOOT_switch_matrix.N1BEG2 ));
 sky130_fd_sc_hd__mux2_1 _067_ (.A0(net26),
    .A1(net23),
    .S(\Inst_S_WARMBOOT_ConfigMem.Inst_frame0_bit14.Q ),
    .X(\Inst_S_WARMBOOT_switch_matrix.N1BEG1 ));
 sky130_fd_sc_hd__mux2_1 _068_ (.A0(net27),
    .A1(net23),
    .S(\Inst_S_WARMBOOT_ConfigMem.Inst_frame0_bit13.Q ),
    .X(\Inst_S_WARMBOOT_switch_matrix.N1BEG0 ));
 sky130_fd_sc_hd__dlxtp_1 _069_ (.D(net1),
    .GATE(net7),
    .Q(\Inst_S_WARMBOOT_ConfigMem.Inst_frame0_bit13.Q ));
 sky130_fd_sc_hd__dlxtp_1 _070_ (.D(net2),
    .GATE(net7),
    .Q(\Inst_S_WARMBOOT_ConfigMem.Inst_frame0_bit14.Q ));
 sky130_fd_sc_hd__dlxtp_1 _071_ (.D(net3),
    .GATE(net7),
    .Q(\Inst_S_WARMBOOT_ConfigMem.Inst_frame0_bit15.Q ));
 sky130_fd_sc_hd__dlxtp_1 _072_ (.D(net4),
    .GATE(net7),
    .Q(\Inst_S_WARMBOOT_ConfigMem.Inst_frame0_bit16.Q ));
 sky130_fd_sc_hd__dlxtp_1 _073_ (.D(net5),
    .GATE(net8),
    .Q(\Inst_S_WARMBOOT_ConfigMem.Inst_frame0_bit17.Q ));
 sky130_fd_sc_hd__dlxtp_1 _074_ (.D(net6),
    .GATE(net8),
    .Q(\Inst_S_WARMBOOT_ConfigMem.Inst_frame0_bit18.Q ));
 sky130_fd_sc_hd__dlxtp_1 _075_ (.D(net9),
    .GATE(net8),
    .Q(\Inst_S_WARMBOOT_ConfigMem.Inst_frame0_bit19.Q ));
 sky130_fd_sc_hd__dlxtp_1 _076_ (.D(net10),
    .GATE(net8),
    .Q(\Inst_S_WARMBOOT_ConfigMem.Inst_frame0_bit20.Q ));
 sky130_fd_sc_hd__dlxtp_1 _077_ (.D(net11),
    .GATE(net8),
    .Q(\Inst_S_WARMBOOT_ConfigMem.Inst_frame0_bit21.Q ));
 sky130_fd_sc_hd__dlxtp_1 _078_ (.D(net12),
    .GATE(net8),
    .Q(\Inst_S_WARMBOOT_ConfigMem.Inst_frame0_bit22.Q ));
 sky130_fd_sc_hd__dlxtp_1 _079_ (.D(net13),
    .GATE(net8),
    .Q(\Inst_S_WARMBOOT_ConfigMem.Inst_frame0_bit23.Q ));
 sky130_fd_sc_hd__dlxtp_1 _080_ (.D(net14),
    .GATE(net8),
    .Q(\Inst_S_WARMBOOT_ConfigMem.Inst_frame0_bit24.Q ));
 sky130_fd_sc_hd__dlxtp_1 _081_ (.D(net15),
    .GATE(net22),
    .Q(\Inst_S_WARMBOOT_ConfigMem.Inst_frame0_bit25.Q ));
 sky130_fd_sc_hd__dlxtp_1 _082_ (.D(net16),
    .GATE(net7),
    .Q(\Inst_S_WARMBOOT_ConfigMem.Inst_frame0_bit26.Q ));
 sky130_fd_sc_hd__dlxtp_1 _083_ (.D(net17),
    .GATE(net7),
    .Q(\Inst_S_WARMBOOT_ConfigMem.Inst_frame0_bit27.Q ));
 sky130_fd_sc_hd__dlxtp_1 _084_ (.D(net18),
    .GATE(net7),
    .Q(\Inst_S_WARMBOOT_ConfigMem.Inst_frame0_bit28.Q ));
 sky130_fd_sc_hd__dlxtp_1 _085_ (.D(net19),
    .GATE(net7),
    .Q(\Inst_S_WARMBOOT_ConfigMem.Inst_frame0_bit29.Q ));
 sky130_fd_sc_hd__dlxtp_1 _086_ (.D(net20),
    .GATE(net7),
    .Q(\Inst_S_WARMBOOT_ConfigMem.Inst_frame0_bit30.Q ));
 sky130_fd_sc_hd__dlxtp_1 _087_ (.D(net21),
    .GATE(net7),
    .Q(\Inst_S_WARMBOOT_ConfigMem.Inst_frame0_bit31.Q ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1 (.DIODE(FrameData[10]));
 sky130_fd_sc_hd__clkbuf_2 _089_ (.A(FrameData[0]),
    .X(net57));
 sky130_fd_sc_hd__clkbuf_1 _090_ (.A(FrameData[1]),
    .X(net68));
 sky130_fd_sc_hd__clkbuf_2 _091_ (.A(FrameData[2]),
    .X(net79));
 sky130_fd_sc_hd__clkbuf_1 _092_ (.A(FrameData[3]),
    .X(net82));
 sky130_fd_sc_hd__clkbuf_2 _093_ (.A(FrameData[4]),
    .X(net83));
 sky130_fd_sc_hd__clkbuf_2 _094_ (.A(FrameData[5]),
    .X(net84));
 sky130_fd_sc_hd__clkbuf_2 _095_ (.A(FrameData[6]),
    .X(net85));
 sky130_fd_sc_hd__clkbuf_1 _096_ (.A(FrameData[7]),
    .X(net86));
 sky130_fd_sc_hd__buf_1 _097_ (.A(FrameData[8]),
    .X(net87));
 sky130_fd_sc_hd__buf_1 _098_ (.A(FrameData[9]),
    .X(net88));
 sky130_fd_sc_hd__clkbuf_2 _099_ (.A(FrameData[10]),
    .X(net58));
 sky130_fd_sc_hd__clkbuf_1 _100_ (.A(FrameData[11]),
    .X(net59));
 sky130_fd_sc_hd__clkbuf_1 _101_ (.A(FrameData[12]),
    .X(net60));
 sky130_fd_sc_hd__buf_1 _102_ (.A(net1),
    .X(net61));
 sky130_fd_sc_hd__buf_1 _103_ (.A(net2),
    .X(net62));
 sky130_fd_sc_hd__buf_1 _104_ (.A(net3),
    .X(net63));
 sky130_fd_sc_hd__clkbuf_1 _105_ (.A(net4),
    .X(net64));
 sky130_fd_sc_hd__clkbuf_2 _106_ (.A(net5),
    .X(net65));
 sky130_fd_sc_hd__clkbuf_2 _107_ (.A(net6),
    .X(net66));
 sky130_fd_sc_hd__clkbuf_2 _108_ (.A(net9),
    .X(net67));
 sky130_fd_sc_hd__buf_1 _109_ (.A(net10),
    .X(net69));
 sky130_fd_sc_hd__buf_1 _110_ (.A(net11),
    .X(net70));
 sky130_fd_sc_hd__clkbuf_1 _111_ (.A(net12),
    .X(net71));
 sky130_fd_sc_hd__buf_1 _112_ (.A(net13),
    .X(net72));
 sky130_fd_sc_hd__buf_1 _113_ (.A(net14),
    .X(net73));
 sky130_fd_sc_hd__buf_1 _114_ (.A(net15),
    .X(net74));
 sky130_fd_sc_hd__buf_1 _115_ (.A(net16),
    .X(net75));
 sky130_fd_sc_hd__buf_1 _116_ (.A(net17),
    .X(net76));
 sky130_fd_sc_hd__buf_1 _117_ (.A(net18),
    .X(net77));
 sky130_fd_sc_hd__clkbuf_2 _118_ (.A(net19),
    .X(net78));
 sky130_fd_sc_hd__buf_1 _119_ (.A(net20),
    .X(net80));
 sky130_fd_sc_hd__clkbuf_2 _120_ (.A(net21),
    .X(net81));
 sky130_fd_sc_hd__buf_1 _121_ (.A(net8),
    .X(net89));
 sky130_fd_sc_hd__clkbuf_1 _122_ (.A(FrameStrobe[1]),
    .X(net100));
 sky130_fd_sc_hd__clkbuf_1 _123_ (.A(FrameStrobe[2]),
    .X(net101));
 sky130_fd_sc_hd__clkbuf_1 _124_ (.A(FrameStrobe[3]),
    .X(net102));
 sky130_fd_sc_hd__clkbuf_1 _125_ (.A(FrameStrobe[4]),
    .X(net103));
 sky130_fd_sc_hd__clkbuf_1 _126_ (.A(FrameStrobe[5]),
    .X(net104));
 sky130_fd_sc_hd__clkbuf_1 _127_ (.A(FrameStrobe[6]),
    .X(net105));
 sky130_fd_sc_hd__clkbuf_1 _128_ (.A(FrameStrobe[7]),
    .X(net106));
 sky130_fd_sc_hd__clkbuf_1 _129_ (.A(FrameStrobe[8]),
    .X(net107));
 sky130_fd_sc_hd__clkbuf_1 _130_ (.A(FrameStrobe[9]),
    .X(net108));
 sky130_fd_sc_hd__clkbuf_1 _131_ (.A(FrameStrobe[10]),
    .X(net90));
 sky130_fd_sc_hd__clkbuf_1 _132_ (.A(FrameStrobe[11]),
    .X(net91));
 sky130_fd_sc_hd__clkbuf_1 _133_ (.A(FrameStrobe[12]),
    .X(net92));
 sky130_fd_sc_hd__clkbuf_1 _134_ (.A(FrameStrobe[13]),
    .X(net93));
 sky130_fd_sc_hd__clkbuf_1 _135_ (.A(FrameStrobe[14]),
    .X(net94));
 sky130_fd_sc_hd__buf_1 _136_ (.A(FrameStrobe[15]),
    .X(net95));
 sky130_fd_sc_hd__buf_1 _137_ (.A(FrameStrobe[16]),
    .X(net96));
 sky130_fd_sc_hd__clkbuf_1 _138_ (.A(FrameStrobe[17]),
    .X(net97));
 sky130_fd_sc_hd__clkbuf_1 _139_ (.A(FrameStrobe[18]),
    .X(net98));
 sky130_fd_sc_hd__clkbuf_1 _140_ (.A(FrameStrobe[19]),
    .X(net99));
 sky130_fd_sc_hd__buf_1 _141_ (.A(\Inst_S_WARMBOOT_switch_matrix.N1BEG0 ),
    .X(net109));
 sky130_fd_sc_hd__buf_1 _142_ (.A(\Inst_S_WARMBOOT_switch_matrix.N1BEG1 ),
    .X(net110));
 sky130_fd_sc_hd__buf_1 _143_ (.A(\Inst_S_WARMBOOT_switch_matrix.N1BEG2 ),
    .X(net111));
 sky130_fd_sc_hd__buf_1 _144_ (.A(\Inst_S_WARMBOOT_switch_matrix.N1BEG3 ),
    .X(net112));
 sky130_fd_sc_hd__buf_1 _145_ (.A(S2MID[7]),
    .X(net113));
 sky130_fd_sc_hd__clkbuf_1 _146_ (.A(S2MID[6]),
    .X(net114));
 sky130_fd_sc_hd__clkbuf_1 _147_ (.A(S2MID[5]),
    .X(net115));
 sky130_fd_sc_hd__clkbuf_1 _148_ (.A(S2MID[4]),
    .X(net116));
 sky130_fd_sc_hd__clkbuf_1 _149_ (.A(net39),
    .X(net117));
 sky130_fd_sc_hd__buf_1 _150_ (.A(net38),
    .X(net118));
 sky130_fd_sc_hd__buf_1 _151_ (.A(net37),
    .X(net119));
 sky130_fd_sc_hd__buf_1 _152_ (.A(net36),
    .X(net120));
 sky130_fd_sc_hd__clkbuf_1 _153_ (.A(net35),
    .X(net121));
 sky130_fd_sc_hd__buf_1 _154_ (.A(net34),
    .X(net122));
 sky130_fd_sc_hd__buf_1 _155_ (.A(net33),
    .X(net123));
 sky130_fd_sc_hd__buf_1 _156_ (.A(net32),
    .X(net124));
 sky130_fd_sc_hd__clkbuf_1 _157_ (.A(net31),
    .X(net125));
 sky130_fd_sc_hd__buf_1 _158_ (.A(net30),
    .X(net126));
 sky130_fd_sc_hd__buf_1 _159_ (.A(net29),
    .X(net127));
 sky130_fd_sc_hd__buf_1 _160_ (.A(net28),
    .X(net128));
 sky130_fd_sc_hd__clkbuf_1 _161_ (.A(S4END[15]),
    .X(net129));
 sky130_fd_sc_hd__clkbuf_2 _162_ (.A(S4END[14]),
    .X(net136));
 sky130_fd_sc_hd__buf_1 _163_ (.A(S4END[13]),
    .X(net137));
 sky130_fd_sc_hd__clkbuf_2 _164_ (.A(S4END[12]),
    .X(net138));
 sky130_fd_sc_hd__buf_1 _165_ (.A(S4END[11]),
    .X(net139));
 sky130_fd_sc_hd__clkbuf_2 _166_ (.A(S4END[10]),
    .X(net140));
 sky130_fd_sc_hd__buf_1 _167_ (.A(S4END[9]),
    .X(net141));
 sky130_fd_sc_hd__clkbuf_1 _168_ (.A(S4END[8]),
    .X(net142));
 sky130_fd_sc_hd__clkbuf_1 _169_ (.A(net47),
    .X(net143));
 sky130_fd_sc_hd__buf_1 _170_ (.A(net46),
    .X(net144));
 sky130_fd_sc_hd__buf_1 _171_ (.A(net45),
    .X(net130));
 sky130_fd_sc_hd__buf_1 _172_ (.A(net44),
    .X(net131));
 sky130_fd_sc_hd__clkbuf_1 _173_ (.A(net43),
    .X(net132));
 sky130_fd_sc_hd__buf_1 _174_ (.A(net42),
    .X(net133));
 sky130_fd_sc_hd__buf_1 _175_ (.A(net41),
    .X(net134));
 sky130_fd_sc_hd__buf_1 _176_ (.A(net40),
    .X(net135));
 sky130_fd_sc_hd__buf_1 _177_ (.A(SS4END[15]),
    .X(net145));
 sky130_fd_sc_hd__buf_1 _178_ (.A(SS4END[14]),
    .X(net152));
 sky130_fd_sc_hd__buf_1 _179_ (.A(SS4END[13]),
    .X(net153));
 sky130_fd_sc_hd__buf_1 _180_ (.A(SS4END[12]),
    .X(net154));
 sky130_fd_sc_hd__buf_1 _181_ (.A(SS4END[11]),
    .X(net155));
 sky130_fd_sc_hd__buf_1 _182_ (.A(SS4END[10]),
    .X(net156));
 sky130_fd_sc_hd__buf_1 _183_ (.A(SS4END[9]),
    .X(net157));
 sky130_fd_sc_hd__buf_1 _184_ (.A(SS4END[8]),
    .X(net158));
 sky130_fd_sc_hd__buf_1 _185_ (.A(net55),
    .X(net159));
 sky130_fd_sc_hd__clkbuf_1 _186_ (.A(net54),
    .X(net160));
 sky130_fd_sc_hd__buf_1 _187_ (.A(net53),
    .X(net146));
 sky130_fd_sc_hd__clkbuf_1 _188_ (.A(net52),
    .X(net147));
 sky130_fd_sc_hd__buf_1 _189_ (.A(net51),
    .X(net148));
 sky130_fd_sc_hd__clkbuf_1 _190_ (.A(net50),
    .X(net149));
 sky130_fd_sc_hd__buf_1 _191_ (.A(net49),
    .X(net150));
 sky130_fd_sc_hd__clkbuf_1 _192_ (.A(net48),
    .X(net151));
 sky130_fd_sc_hd__buf_2 _193_ (.A(UserCLK),
    .X(net165));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_0_Right_0 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_1_Right_1 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_2_Right_2 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_3_Right_3 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_4_Right_4 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_5_Right_5 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_6_Right_6 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_7_Right_7 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_8_Right_8 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_9_Right_9 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_10_Right_10 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_11_Right_11 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_0_Left_12 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_1_Left_13 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_2_Left_14 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_3_Left_15 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_4_Left_16 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_5_Left_17 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_6_Left_18 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_7_Left_19 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_8_Left_20 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_9_Left_21 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_10_Left_22 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_11_Left_23 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_24 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_25 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_26 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_27 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_28 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_29 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_30 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_31 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_32 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_33 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_34 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_35 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_36 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_37 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_38 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_39 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_40 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_41 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_42 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_43 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_44 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_45 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_46 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_47 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_48 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_49 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_50 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_51 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_52 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_53 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_54 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_55 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_56 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_57 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_58 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_59 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_60 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_61 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_62 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_63 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_64 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_65 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_66 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_67 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_68 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_69 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_70 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_71 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_72 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_73 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_74 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_75 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_76 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_77 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_78 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_79 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_80 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_81 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_82 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_83 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_84 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_85 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_86 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_87 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_88 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_89 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_90 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_91 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_92 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_93 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_94 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_95 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_96 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_97 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_98 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_99 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_121 ();
 sky130_fd_sc_hd__clkbuf_2 fanout7 (.A(net8),
    .X(net7));
 sky130_fd_sc_hd__buf_2 fanout8 (.A(net22),
    .X(net8));
 sky130_fd_sc_hd__buf_1 input1 (.A(FrameData[13]),
    .X(net1));
 sky130_fd_sc_hd__buf_1 input2 (.A(FrameData[14]),
    .X(net2));
 sky130_fd_sc_hd__buf_1 input3 (.A(FrameData[15]),
    .X(net3));
 sky130_fd_sc_hd__buf_1 input4 (.A(FrameData[16]),
    .X(net4));
 sky130_fd_sc_hd__buf_1 input5 (.A(FrameData[17]),
    .X(net5));
 sky130_fd_sc_hd__clkbuf_1 input6 (.A(FrameData[18]),
    .X(net6));
 sky130_fd_sc_hd__buf_1 input7 (.A(FrameData[19]),
    .X(net9));
 sky130_fd_sc_hd__buf_1 input8 (.A(FrameData[20]),
    .X(net10));
 sky130_fd_sc_hd__buf_1 input9 (.A(FrameData[21]),
    .X(net11));
 sky130_fd_sc_hd__buf_1 input10 (.A(FrameData[22]),
    .X(net12));
 sky130_fd_sc_hd__buf_1 input11 (.A(FrameData[23]),
    .X(net13));
 sky130_fd_sc_hd__dlymetal6s2s_1 input12 (.A(FrameData[24]),
    .X(net14));
 sky130_fd_sc_hd__buf_1 input13 (.A(FrameData[25]),
    .X(net15));
 sky130_fd_sc_hd__buf_1 input14 (.A(FrameData[26]),
    .X(net16));
 sky130_fd_sc_hd__clkbuf_1 input15 (.A(FrameData[27]),
    .X(net17));
 sky130_fd_sc_hd__buf_1 input16 (.A(FrameData[28]),
    .X(net18));
 sky130_fd_sc_hd__buf_1 input17 (.A(FrameData[29]),
    .X(net19));
 sky130_fd_sc_hd__buf_1 input18 (.A(FrameData[30]),
    .X(net20));
 sky130_fd_sc_hd__buf_1 input19 (.A(FrameData[31]),
    .X(net21));
 sky130_fd_sc_hd__buf_1 input20 (.A(FrameStrobe[0]),
    .X(net22));
 sky130_fd_sc_hd__dlymetal6s2s_1 input21 (.A(RESET_top),
    .X(net23));
 sky130_fd_sc_hd__buf_1 input22 (.A(S1END[0]),
    .X(net24));
 sky130_fd_sc_hd__buf_1 input23 (.A(S1END[1]),
    .X(net25));
 sky130_fd_sc_hd__clkbuf_1 input24 (.A(S1END[2]),
    .X(net26));
 sky130_fd_sc_hd__buf_1 input25 (.A(S1END[3]),
    .X(net27));
 sky130_fd_sc_hd__buf_1 input26 (.A(S2END[0]),
    .X(net28));
 sky130_fd_sc_hd__buf_1 input27 (.A(S2END[1]),
    .X(net29));
 sky130_fd_sc_hd__clkbuf_1 input28 (.A(S2END[2]),
    .X(net30));
 sky130_fd_sc_hd__buf_1 input29 (.A(S2END[3]),
    .X(net31));
 sky130_fd_sc_hd__buf_1 input30 (.A(S2END[4]),
    .X(net32));
 sky130_fd_sc_hd__buf_1 input31 (.A(S2END[5]),
    .X(net33));
 sky130_fd_sc_hd__clkbuf_1 input32 (.A(S2END[6]),
    .X(net34));
 sky130_fd_sc_hd__buf_1 input33 (.A(S2END[7]),
    .X(net35));
 sky130_fd_sc_hd__buf_1 input34 (.A(S2MID[0]),
    .X(net36));
 sky130_fd_sc_hd__buf_1 input35 (.A(S2MID[1]),
    .X(net37));
 sky130_fd_sc_hd__clkbuf_1 input36 (.A(S2MID[2]),
    .X(net38));
 sky130_fd_sc_hd__clkbuf_1 input37 (.A(S2MID[3]),
    .X(net39));
 sky130_fd_sc_hd__clkbuf_1 input38 (.A(S4END[0]),
    .X(net40));
 sky130_fd_sc_hd__buf_1 input39 (.A(S4END[1]),
    .X(net41));
 sky130_fd_sc_hd__clkbuf_1 input40 (.A(S4END[2]),
    .X(net42));
 sky130_fd_sc_hd__buf_1 input41 (.A(S4END[3]),
    .X(net43));
 sky130_fd_sc_hd__clkbuf_1 input42 (.A(S4END[4]),
    .X(net44));
 sky130_fd_sc_hd__buf_1 input43 (.A(S4END[5]),
    .X(net45));
 sky130_fd_sc_hd__clkbuf_1 input44 (.A(S4END[6]),
    .X(net46));
 sky130_fd_sc_hd__buf_1 input45 (.A(S4END[7]),
    .X(net47));
 sky130_fd_sc_hd__buf_1 input46 (.A(SS4END[0]),
    .X(net48));
 sky130_fd_sc_hd__clkbuf_1 input47 (.A(SS4END[1]),
    .X(net49));
 sky130_fd_sc_hd__buf_1 input48 (.A(SS4END[2]),
    .X(net50));
 sky130_fd_sc_hd__dlymetal6s2s_1 input49 (.A(SS4END[3]),
    .X(net51));
 sky130_fd_sc_hd__buf_1 input50 (.A(SS4END[4]),
    .X(net52));
 sky130_fd_sc_hd__clkbuf_1 input51 (.A(SS4END[5]),
    .X(net53));
 sky130_fd_sc_hd__buf_1 input52 (.A(SS4END[6]),
    .X(net54));
 sky130_fd_sc_hd__clkbuf_2 input53 (.A(SS4END[7]),
    .X(net55));
 sky130_fd_sc_hd__buf_2 output54 (.A(net56),
    .X(BOOT_top));
 sky130_fd_sc_hd__buf_2 output55 (.A(net57),
    .X(FrameData_O[0]));
 sky130_fd_sc_hd__buf_2 output56 (.A(net58),
    .X(FrameData_O[10]));
 sky130_fd_sc_hd__buf_2 output57 (.A(net59),
    .X(FrameData_O[11]));
 sky130_fd_sc_hd__buf_2 output58 (.A(net60),
    .X(FrameData_O[12]));
 sky130_fd_sc_hd__buf_2 output59 (.A(net61),
    .X(FrameData_O[13]));
 sky130_fd_sc_hd__buf_2 output60 (.A(net62),
    .X(FrameData_O[14]));
 sky130_fd_sc_hd__buf_2 output61 (.A(net63),
    .X(FrameData_O[15]));
 sky130_fd_sc_hd__buf_2 output62 (.A(net64),
    .X(FrameData_O[16]));
 sky130_fd_sc_hd__buf_2 output63 (.A(net65),
    .X(FrameData_O[17]));
 sky130_fd_sc_hd__buf_2 output64 (.A(net66),
    .X(FrameData_O[18]));
 sky130_fd_sc_hd__buf_2 output65 (.A(net67),
    .X(FrameData_O[19]));
 sky130_fd_sc_hd__buf_2 output66 (.A(net68),
    .X(FrameData_O[1]));
 sky130_fd_sc_hd__buf_2 output67 (.A(net69),
    .X(FrameData_O[20]));
 sky130_fd_sc_hd__buf_2 output68 (.A(net70),
    .X(FrameData_O[21]));
 sky130_fd_sc_hd__buf_2 output69 (.A(net71),
    .X(FrameData_O[22]));
 sky130_fd_sc_hd__buf_2 output70 (.A(net72),
    .X(FrameData_O[23]));
 sky130_fd_sc_hd__buf_2 output71 (.A(net73),
    .X(FrameData_O[24]));
 sky130_fd_sc_hd__buf_2 output72 (.A(net74),
    .X(FrameData_O[25]));
 sky130_fd_sc_hd__buf_2 output73 (.A(net75),
    .X(FrameData_O[26]));
 sky130_fd_sc_hd__buf_2 output74 (.A(net76),
    .X(FrameData_O[27]));
 sky130_fd_sc_hd__buf_2 output75 (.A(net77),
    .X(FrameData_O[28]));
 sky130_fd_sc_hd__buf_2 output76 (.A(net78),
    .X(FrameData_O[29]));
 sky130_fd_sc_hd__buf_2 output77 (.A(net79),
    .X(FrameData_O[2]));
 sky130_fd_sc_hd__buf_2 output78 (.A(net80),
    .X(FrameData_O[30]));
 sky130_fd_sc_hd__buf_2 output79 (.A(net81),
    .X(FrameData_O[31]));
 sky130_fd_sc_hd__buf_2 output80 (.A(net82),
    .X(FrameData_O[3]));
 sky130_fd_sc_hd__buf_2 output81 (.A(net83),
    .X(FrameData_O[4]));
 sky130_fd_sc_hd__buf_2 output82 (.A(net84),
    .X(FrameData_O[5]));
 sky130_fd_sc_hd__buf_2 output83 (.A(net85),
    .X(FrameData_O[6]));
 sky130_fd_sc_hd__buf_2 output84 (.A(net86),
    .X(FrameData_O[7]));
 sky130_fd_sc_hd__buf_2 output85 (.A(net87),
    .X(FrameData_O[8]));
 sky130_fd_sc_hd__buf_2 output86 (.A(net88),
    .X(FrameData_O[9]));
 sky130_fd_sc_hd__buf_2 output87 (.A(net89),
    .X(FrameStrobe_O[0]));
 sky130_fd_sc_hd__buf_2 output88 (.A(net90),
    .X(FrameStrobe_O[10]));
 sky130_fd_sc_hd__buf_2 output89 (.A(net91),
    .X(FrameStrobe_O[11]));
 sky130_fd_sc_hd__buf_2 output90 (.A(net92),
    .X(FrameStrobe_O[12]));
 sky130_fd_sc_hd__buf_2 output91 (.A(net93),
    .X(FrameStrobe_O[13]));
 sky130_fd_sc_hd__buf_2 output92 (.A(net94),
    .X(FrameStrobe_O[14]));
 sky130_fd_sc_hd__buf_2 output93 (.A(net95),
    .X(FrameStrobe_O[15]));
 sky130_fd_sc_hd__buf_2 output94 (.A(net96),
    .X(FrameStrobe_O[16]));
 sky130_fd_sc_hd__buf_2 output95 (.A(net97),
    .X(FrameStrobe_O[17]));
 sky130_fd_sc_hd__buf_2 output96 (.A(net98),
    .X(FrameStrobe_O[18]));
 sky130_fd_sc_hd__buf_2 output97 (.A(net99),
    .X(FrameStrobe_O[19]));
 sky130_fd_sc_hd__buf_2 output98 (.A(net100),
    .X(FrameStrobe_O[1]));
 sky130_fd_sc_hd__buf_2 output99 (.A(net101),
    .X(FrameStrobe_O[2]));
 sky130_fd_sc_hd__buf_2 output100 (.A(net102),
    .X(FrameStrobe_O[3]));
 sky130_fd_sc_hd__buf_2 output101 (.A(net103),
    .X(FrameStrobe_O[4]));
 sky130_fd_sc_hd__buf_2 output102 (.A(net104),
    .X(FrameStrobe_O[5]));
 sky130_fd_sc_hd__buf_2 output103 (.A(net105),
    .X(FrameStrobe_O[6]));
 sky130_fd_sc_hd__buf_2 output104 (.A(net106),
    .X(FrameStrobe_O[7]));
 sky130_fd_sc_hd__buf_2 output105 (.A(net107),
    .X(FrameStrobe_O[8]));
 sky130_fd_sc_hd__buf_2 output106 (.A(net108),
    .X(FrameStrobe_O[9]));
 sky130_fd_sc_hd__buf_2 output107 (.A(net109),
    .X(N1BEG[0]));
 sky130_fd_sc_hd__buf_2 output108 (.A(net110),
    .X(N1BEG[1]));
 sky130_fd_sc_hd__buf_2 output109 (.A(net111),
    .X(N1BEG[2]));
 sky130_fd_sc_hd__buf_2 output110 (.A(net112),
    .X(N1BEG[3]));
 sky130_fd_sc_hd__buf_2 output111 (.A(net113),
    .X(N2BEG[0]));
 sky130_fd_sc_hd__buf_2 output112 (.A(net114),
    .X(N2BEG[1]));
 sky130_fd_sc_hd__buf_2 output113 (.A(net115),
    .X(N2BEG[2]));
 sky130_fd_sc_hd__buf_2 output114 (.A(net116),
    .X(N2BEG[3]));
 sky130_fd_sc_hd__buf_2 output115 (.A(net117),
    .X(N2BEG[4]));
 sky130_fd_sc_hd__buf_2 output116 (.A(net118),
    .X(N2BEG[5]));
 sky130_fd_sc_hd__buf_2 output117 (.A(net119),
    .X(N2BEG[6]));
 sky130_fd_sc_hd__buf_2 output118 (.A(net120),
    .X(N2BEG[7]));
 sky130_fd_sc_hd__buf_2 output119 (.A(net121),
    .X(N2BEGb[0]));
 sky130_fd_sc_hd__buf_2 output120 (.A(net122),
    .X(N2BEGb[1]));
 sky130_fd_sc_hd__buf_2 output121 (.A(net123),
    .X(N2BEGb[2]));
 sky130_fd_sc_hd__buf_2 output122 (.A(net124),
    .X(N2BEGb[3]));
 sky130_fd_sc_hd__buf_2 output123 (.A(net125),
    .X(N2BEGb[4]));
 sky130_fd_sc_hd__buf_2 output124 (.A(net126),
    .X(N2BEGb[5]));
 sky130_fd_sc_hd__buf_2 output125 (.A(net127),
    .X(N2BEGb[6]));
 sky130_fd_sc_hd__buf_2 output126 (.A(net128),
    .X(N2BEGb[7]));
 sky130_fd_sc_hd__buf_2 output127 (.A(net129),
    .X(N4BEG[0]));
 sky130_fd_sc_hd__buf_2 output128 (.A(net130),
    .X(N4BEG[10]));
 sky130_fd_sc_hd__buf_2 output129 (.A(net131),
    .X(N4BEG[11]));
 sky130_fd_sc_hd__buf_2 output130 (.A(net132),
    .X(N4BEG[12]));
 sky130_fd_sc_hd__buf_2 output131 (.A(net133),
    .X(N4BEG[13]));
 sky130_fd_sc_hd__buf_2 output132 (.A(net134),
    .X(N4BEG[14]));
 sky130_fd_sc_hd__buf_2 output133 (.A(net135),
    .X(N4BEG[15]));
 sky130_fd_sc_hd__buf_2 output134 (.A(net136),
    .X(N4BEG[1]));
 sky130_fd_sc_hd__buf_2 output135 (.A(net137),
    .X(N4BEG[2]));
 sky130_fd_sc_hd__buf_2 output136 (.A(net138),
    .X(N4BEG[3]));
 sky130_fd_sc_hd__buf_2 output137 (.A(net139),
    .X(N4BEG[4]));
 sky130_fd_sc_hd__buf_2 output138 (.A(net140),
    .X(N4BEG[5]));
 sky130_fd_sc_hd__buf_2 output139 (.A(net141),
    .X(N4BEG[6]));
 sky130_fd_sc_hd__buf_2 output140 (.A(net142),
    .X(N4BEG[7]));
 sky130_fd_sc_hd__buf_2 output141 (.A(net143),
    .X(N4BEG[8]));
 sky130_fd_sc_hd__buf_2 output142 (.A(net144),
    .X(N4BEG[9]));
 sky130_fd_sc_hd__buf_2 output143 (.A(net145),
    .X(NN4BEG[0]));
 sky130_fd_sc_hd__buf_2 output144 (.A(net146),
    .X(NN4BEG[10]));
 sky130_fd_sc_hd__buf_2 output145 (.A(net147),
    .X(NN4BEG[11]));
 sky130_fd_sc_hd__buf_2 output146 (.A(net148),
    .X(NN4BEG[12]));
 sky130_fd_sc_hd__buf_2 output147 (.A(net149),
    .X(NN4BEG[13]));
 sky130_fd_sc_hd__buf_2 output148 (.A(net150),
    .X(NN4BEG[14]));
 sky130_fd_sc_hd__buf_2 output149 (.A(net151),
    .X(NN4BEG[15]));
 sky130_fd_sc_hd__buf_2 output150 (.A(net152),
    .X(NN4BEG[1]));
 sky130_fd_sc_hd__buf_2 output151 (.A(net153),
    .X(NN4BEG[2]));
 sky130_fd_sc_hd__buf_2 output152 (.A(net154),
    .X(NN4BEG[3]));
 sky130_fd_sc_hd__buf_2 output153 (.A(net155),
    .X(NN4BEG[4]));
 sky130_fd_sc_hd__buf_2 output154 (.A(net156),
    .X(NN4BEG[5]));
 sky130_fd_sc_hd__buf_2 output155 (.A(net157),
    .X(NN4BEG[6]));
 sky130_fd_sc_hd__buf_2 output156 (.A(net158),
    .X(NN4BEG[7]));
 sky130_fd_sc_hd__buf_2 output157 (.A(net159),
    .X(NN4BEG[8]));
 sky130_fd_sc_hd__buf_2 output158 (.A(net160),
    .X(NN4BEG[9]));
 sky130_fd_sc_hd__buf_2 output159 (.A(net161),
    .X(SLOT_top0));
 sky130_fd_sc_hd__buf_2 output160 (.A(net162),
    .X(SLOT_top1));
 sky130_fd_sc_hd__buf_2 output161 (.A(net163),
    .X(SLOT_top2));
 sky130_fd_sc_hd__buf_2 output162 (.A(net164),
    .X(SLOT_top3));
 sky130_fd_sc_hd__buf_1 output163 (.A(net165),
    .X(UserCLKo));
 sky130_fd_sc_hd__conb_1 S_WARMBOOT_164 (.LO(net166));
 sky130_fd_sc_hd__diode_2 ANTENNA_2 (.DIODE(FrameData[11]));
 sky130_fd_sc_hd__diode_2 ANTENNA_3 (.DIODE(FrameData[1]));
 sky130_fd_sc_hd__diode_2 ANTENNA_4 (.DIODE(FrameData[3]));
 sky130_fd_sc_hd__diode_2 ANTENNA_5 (.DIODE(FrameData[8]));
 sky130_fd_sc_hd__diode_2 ANTENNA_6 (.DIODE(FrameData[9]));
 sky130_fd_sc_hd__diode_2 ANTENNA_7 (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA_8 (.DIODE(FrameStrobe[1]));
 sky130_fd_sc_hd__diode_2 ANTENNA_9 (.DIODE(FrameStrobe[4]));
 sky130_fd_sc_hd__diode_2 ANTENNA_10 (.DIODE(FrameStrobe[5]));
 sky130_fd_sc_hd__diode_2 ANTENNA_11 (.DIODE(net14));
 sky130_fd_sc_hd__diode_2 ANTENNA_12 (.DIODE(net51));
 sky130_fd_sc_hd__diode_2 ANTENNA_13 (.DIODE(net71));
 sky130_fd_sc_hd__decap_6 FILLER_0_13 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_389 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_397 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_219 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_247 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_278 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_289 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_294 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_302 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_312 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_342 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_354 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_367 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_379 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_386 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_52 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_64 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_76 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_117 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_389 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_409 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_30 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_42 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_75 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_81 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_125 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_164 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_173 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_179 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_183 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_292 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_316 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_342 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_354 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_366 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_390 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_397 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_82 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_107 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_122 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_156 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_176 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_187 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_257 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_272 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_284 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_312 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_316 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_328 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_340 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_352 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_356 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_371 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_375 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_387 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_392 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_400 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_412 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_6 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_18 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_30 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_37 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_75 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_86 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_98 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_106 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_273 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_344 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_348 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_355 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_367 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_409 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_9 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_21 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_64 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_76 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_105 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_114 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_171 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_233 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_269 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_291 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_312 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_324 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_336 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_389 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_31 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_43 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_62 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_74 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_86 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_95 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_145 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_167 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_175 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_198 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_231 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_243 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_255 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_320 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_324 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_355 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_359 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_371 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_391 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_400 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_12 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_24 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_80 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_274 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_389 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_396 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_400 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_12 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_24 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_36 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_48 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_75 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_84 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_90 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_189 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_213 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_268 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_293 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_313 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_397 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_21 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_37 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_43 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_59 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_64 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_70 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_76 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_94 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_106 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_115 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_130 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_134 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_148 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_157 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_161 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_174 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_232 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_250 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_256 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_264 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_268 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_280 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_285 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_312 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_324 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_332 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_338 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_342 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_361 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_372 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_385 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_399 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_410 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_19 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_175 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_207 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_222 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_362 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_409 ();
 assign Co = net166;
endmodule
