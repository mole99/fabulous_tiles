magic
tech ihp-sg13g2
magscale 1 2
timestamp 1743692509
<< metal1 >>
rect 1152 9848 45216 9872
rect 1152 9808 3688 9848
rect 3728 9808 3770 9848
rect 3810 9808 3852 9848
rect 3892 9808 3934 9848
rect 3974 9808 4016 9848
rect 4056 9808 18808 9848
rect 18848 9808 18890 9848
rect 18930 9808 18972 9848
rect 19012 9808 19054 9848
rect 19094 9808 19136 9848
rect 19176 9808 33928 9848
rect 33968 9808 34010 9848
rect 34050 9808 34092 9848
rect 34132 9808 34174 9848
rect 34214 9808 34256 9848
rect 34296 9808 45216 9848
rect 1152 9784 45216 9808
rect 2235 9680 2277 9689
rect 2235 9640 2236 9680
rect 2276 9640 2277 9680
rect 2235 9631 2277 9640
rect 10203 9680 10245 9689
rect 10203 9640 10204 9680
rect 10244 9640 10245 9680
rect 10203 9631 10245 9640
rect 11355 9680 11397 9689
rect 11355 9640 11356 9680
rect 11396 9640 11397 9680
rect 11355 9631 11397 9640
rect 12123 9680 12165 9689
rect 12123 9640 12124 9680
rect 12164 9640 12165 9680
rect 12123 9631 12165 9640
rect 12891 9680 12933 9689
rect 12891 9640 12892 9680
rect 12932 9640 12933 9680
rect 12891 9631 12933 9640
rect 13275 9680 13317 9689
rect 13275 9640 13276 9680
rect 13316 9640 13317 9680
rect 13275 9631 13317 9640
rect 14043 9680 14085 9689
rect 14043 9640 14044 9680
rect 14084 9640 14085 9680
rect 14043 9631 14085 9640
rect 14811 9680 14853 9689
rect 14811 9640 14812 9680
rect 14852 9640 14853 9680
rect 14811 9631 14853 9640
rect 15195 9680 15237 9689
rect 15195 9640 15196 9680
rect 15236 9640 15237 9680
rect 15195 9631 15237 9640
rect 15579 9680 15621 9689
rect 15579 9640 15580 9680
rect 15620 9640 15621 9680
rect 15579 9631 15621 9640
rect 15963 9680 16005 9689
rect 15963 9640 15964 9680
rect 16004 9640 16005 9680
rect 15963 9631 16005 9640
rect 16347 9680 16389 9689
rect 16347 9640 16348 9680
rect 16388 9640 16389 9680
rect 16347 9631 16389 9640
rect 16731 9680 16773 9689
rect 16731 9640 16732 9680
rect 16772 9640 16773 9680
rect 16731 9631 16773 9640
rect 17115 9680 17157 9689
rect 17115 9640 17116 9680
rect 17156 9640 17157 9680
rect 17115 9631 17157 9640
rect 17499 9680 17541 9689
rect 17499 9640 17500 9680
rect 17540 9640 17541 9680
rect 17499 9631 17541 9640
rect 17883 9680 17925 9689
rect 17883 9640 17884 9680
rect 17924 9640 17925 9680
rect 17883 9631 17925 9640
rect 18267 9680 18309 9689
rect 18267 9640 18268 9680
rect 18308 9640 18309 9680
rect 18267 9631 18309 9640
rect 18651 9680 18693 9689
rect 18651 9640 18652 9680
rect 18692 9640 18693 9680
rect 18651 9631 18693 9640
rect 19803 9680 19845 9689
rect 19803 9640 19804 9680
rect 19844 9640 19845 9680
rect 19803 9631 19845 9640
rect 20187 9680 20229 9689
rect 20187 9640 20188 9680
rect 20228 9640 20229 9680
rect 20187 9631 20229 9640
rect 20571 9680 20613 9689
rect 20571 9640 20572 9680
rect 20612 9640 20613 9680
rect 20571 9631 20613 9640
rect 21339 9680 21381 9689
rect 21339 9640 21340 9680
rect 21380 9640 21381 9680
rect 21339 9631 21381 9640
rect 25851 9680 25893 9689
rect 25851 9640 25852 9680
rect 25892 9640 25893 9680
rect 25851 9631 25893 9640
rect 27387 9680 27429 9689
rect 27387 9640 27388 9680
rect 27428 9640 27429 9680
rect 27387 9631 27429 9640
rect 31227 9680 31269 9689
rect 31227 9640 31228 9680
rect 31268 9640 31269 9680
rect 31227 9631 31269 9640
rect 31995 9680 32037 9689
rect 31995 9640 31996 9680
rect 32036 9640 32037 9680
rect 31995 9631 32037 9640
rect 34299 9680 34341 9689
rect 34299 9640 34300 9680
rect 34340 9640 34341 9680
rect 34299 9631 34341 9640
rect 34683 9680 34725 9689
rect 34683 9640 34684 9680
rect 34724 9640 34725 9680
rect 34683 9631 34725 9640
rect 35835 9680 35877 9689
rect 35835 9640 35836 9680
rect 35876 9640 35877 9680
rect 35835 9631 35877 9640
rect 42843 9680 42885 9689
rect 42843 9640 42844 9680
rect 42884 9640 42885 9680
rect 42843 9631 42885 9640
rect 43995 9680 44037 9689
rect 43995 9640 43996 9680
rect 44036 9640 44037 9680
rect 43995 9631 44037 9640
rect 44379 9680 44421 9689
rect 44379 9640 44380 9680
rect 44420 9640 44421 9680
rect 44379 9631 44421 9640
rect 44763 9680 44805 9689
rect 44763 9640 44764 9680
rect 44804 9640 44805 9680
rect 44763 9631 44805 9640
rect 10587 9596 10629 9605
rect 10587 9556 10588 9596
rect 10628 9556 10629 9596
rect 10587 9547 10629 9556
rect 11739 9596 11781 9605
rect 11739 9556 11740 9596
rect 11780 9556 11781 9596
rect 11739 9547 11781 9556
rect 12507 9596 12549 9605
rect 12507 9556 12508 9596
rect 12548 9556 12549 9596
rect 12507 9547 12549 9556
rect 13659 9596 13701 9605
rect 13659 9556 13660 9596
rect 13700 9556 13701 9596
rect 13659 9547 13701 9556
rect 14427 9596 14469 9605
rect 14427 9556 14428 9596
rect 14468 9556 14469 9596
rect 14427 9547 14469 9556
rect 19035 9596 19077 9605
rect 19035 9556 19036 9596
rect 19076 9556 19077 9596
rect 19035 9547 19077 9556
rect 28827 9596 28869 9605
rect 28827 9556 28828 9596
rect 28868 9556 28869 9596
rect 28827 9547 28869 9556
rect 31611 9596 31653 9605
rect 31611 9556 31612 9596
rect 31652 9556 31653 9596
rect 31611 9547 31653 9556
rect 32379 9596 32421 9605
rect 32379 9556 32380 9596
rect 32420 9556 32421 9596
rect 32379 9547 32421 9556
rect 33531 9596 33573 9605
rect 33531 9556 33532 9596
rect 33572 9556 33573 9596
rect 33531 9547 33573 9556
rect 35451 9596 35493 9605
rect 35451 9556 35452 9596
rect 35492 9556 35493 9596
rect 35451 9547 35493 9556
rect 1227 9512 1269 9521
rect 1227 9472 1228 9512
rect 1268 9472 1269 9512
rect 1227 9463 1269 9472
rect 1611 9512 1653 9521
rect 1611 9472 1612 9512
rect 1652 9472 1653 9512
rect 1611 9463 1653 9472
rect 1995 9512 2037 9521
rect 1995 9472 1996 9512
rect 2036 9472 2037 9512
rect 1995 9463 2037 9472
rect 2379 9512 2421 9521
rect 2379 9472 2380 9512
rect 2420 9472 2421 9512
rect 2379 9463 2421 9472
rect 2763 9512 2805 9521
rect 2763 9472 2764 9512
rect 2804 9472 2805 9512
rect 2763 9463 2805 9472
rect 3147 9512 3189 9521
rect 3147 9472 3148 9512
rect 3188 9472 3189 9512
rect 3147 9463 3189 9472
rect 9963 9512 10005 9521
rect 9963 9472 9964 9512
rect 10004 9472 10005 9512
rect 9963 9463 10005 9472
rect 10347 9512 10389 9521
rect 10347 9472 10348 9512
rect 10388 9472 10389 9512
rect 10347 9463 10389 9472
rect 10731 9512 10773 9521
rect 10731 9472 10732 9512
rect 10772 9472 10773 9512
rect 10731 9463 10773 9472
rect 11115 9512 11157 9521
rect 11115 9472 11116 9512
rect 11156 9472 11157 9512
rect 11115 9463 11157 9472
rect 11499 9512 11541 9521
rect 11499 9472 11500 9512
rect 11540 9472 11541 9512
rect 11499 9463 11541 9472
rect 11883 9512 11925 9521
rect 11883 9472 11884 9512
rect 11924 9472 11925 9512
rect 11883 9463 11925 9472
rect 12267 9512 12309 9521
rect 12267 9472 12268 9512
rect 12308 9472 12309 9512
rect 12267 9463 12309 9472
rect 12651 9512 12693 9521
rect 12651 9472 12652 9512
rect 12692 9472 12693 9512
rect 12651 9463 12693 9472
rect 13035 9512 13077 9521
rect 13035 9472 13036 9512
rect 13076 9472 13077 9512
rect 13035 9463 13077 9472
rect 13419 9512 13461 9521
rect 13419 9472 13420 9512
rect 13460 9472 13461 9512
rect 13419 9463 13461 9472
rect 13803 9512 13845 9521
rect 13803 9472 13804 9512
rect 13844 9472 13845 9512
rect 13803 9463 13845 9472
rect 14187 9512 14229 9521
rect 14187 9472 14188 9512
rect 14228 9472 14229 9512
rect 14187 9463 14229 9472
rect 14571 9512 14613 9521
rect 14571 9472 14572 9512
rect 14612 9472 14613 9512
rect 14571 9463 14613 9472
rect 14955 9512 14997 9521
rect 14955 9472 14956 9512
rect 14996 9472 14997 9512
rect 14955 9463 14997 9472
rect 15339 9512 15381 9521
rect 15339 9472 15340 9512
rect 15380 9472 15381 9512
rect 15339 9463 15381 9472
rect 15723 9512 15765 9521
rect 15723 9472 15724 9512
rect 15764 9472 15765 9512
rect 15723 9463 15765 9472
rect 16107 9512 16149 9521
rect 16107 9472 16108 9512
rect 16148 9472 16149 9512
rect 16107 9463 16149 9472
rect 16491 9512 16533 9521
rect 16491 9472 16492 9512
rect 16532 9472 16533 9512
rect 16491 9463 16533 9472
rect 16875 9512 16917 9521
rect 16875 9472 16876 9512
rect 16916 9472 16917 9512
rect 16875 9463 16917 9472
rect 17259 9512 17301 9521
rect 17259 9472 17260 9512
rect 17300 9472 17301 9512
rect 17259 9463 17301 9472
rect 17643 9512 17685 9521
rect 17643 9472 17644 9512
rect 17684 9472 17685 9512
rect 17643 9463 17685 9472
rect 18027 9512 18069 9521
rect 18027 9472 18028 9512
rect 18068 9472 18069 9512
rect 18027 9463 18069 9472
rect 18411 9512 18453 9521
rect 18411 9472 18412 9512
rect 18452 9472 18453 9512
rect 18411 9463 18453 9472
rect 18795 9512 18837 9521
rect 18795 9472 18796 9512
rect 18836 9472 18837 9512
rect 18795 9463 18837 9472
rect 19179 9512 19221 9521
rect 19179 9472 19180 9512
rect 19220 9472 19221 9512
rect 19179 9463 19221 9472
rect 19594 9512 19652 9513
rect 19594 9472 19603 9512
rect 19643 9472 19652 9512
rect 19594 9471 19652 9472
rect 19947 9512 19989 9521
rect 19947 9472 19948 9512
rect 19988 9472 19989 9512
rect 19947 9463 19989 9472
rect 20331 9512 20373 9521
rect 20331 9472 20332 9512
rect 20372 9472 20373 9512
rect 20331 9463 20373 9472
rect 20907 9512 20949 9521
rect 20907 9472 20908 9512
rect 20948 9472 20949 9512
rect 20907 9463 20949 9472
rect 21099 9512 21141 9521
rect 21099 9472 21100 9512
rect 21140 9472 21141 9512
rect 21099 9463 21141 9472
rect 21675 9512 21717 9521
rect 21675 9472 21676 9512
rect 21716 9472 21717 9512
rect 21675 9463 21717 9472
rect 21867 9512 21909 9521
rect 21867 9472 21868 9512
rect 21908 9472 21909 9512
rect 21867 9463 21909 9472
rect 22251 9512 22293 9521
rect 22251 9472 22252 9512
rect 22292 9472 22293 9512
rect 22251 9463 22293 9472
rect 22827 9512 22869 9521
rect 22827 9472 22828 9512
rect 22868 9472 22869 9512
rect 22827 9463 22869 9472
rect 23211 9512 23253 9521
rect 23211 9472 23212 9512
rect 23252 9472 23253 9512
rect 23211 9463 23253 9472
rect 23595 9512 23637 9521
rect 23595 9472 23596 9512
rect 23636 9472 23637 9512
rect 23595 9463 23637 9472
rect 24171 9512 24213 9521
rect 24171 9472 24172 9512
rect 24212 9472 24213 9512
rect 24171 9463 24213 9472
rect 24555 9512 24597 9521
rect 24555 9472 24556 9512
rect 24596 9472 24597 9512
rect 24555 9463 24597 9472
rect 24747 9512 24789 9521
rect 24747 9472 24748 9512
rect 24788 9472 24789 9512
rect 24747 9463 24789 9472
rect 25131 9512 25173 9521
rect 25131 9472 25132 9512
rect 25172 9472 25173 9512
rect 25131 9463 25173 9472
rect 25707 9512 25749 9521
rect 25707 9472 25708 9512
rect 25748 9472 25749 9512
rect 25707 9463 25749 9472
rect 26091 9512 26133 9521
rect 26091 9472 26092 9512
rect 26132 9472 26133 9512
rect 26091 9463 26133 9472
rect 26283 9512 26325 9521
rect 26283 9472 26284 9512
rect 26324 9472 26325 9512
rect 26283 9463 26325 9472
rect 26859 9512 26901 9521
rect 26859 9472 26860 9512
rect 26900 9472 26901 9512
rect 26859 9463 26901 9472
rect 27051 9512 27093 9521
rect 27051 9472 27052 9512
rect 27092 9472 27093 9512
rect 27051 9463 27093 9472
rect 27627 9512 27669 9521
rect 27627 9472 27628 9512
rect 27668 9472 27669 9512
rect 27627 9463 27669 9472
rect 28395 9512 28437 9521
rect 28395 9472 28396 9512
rect 28436 9472 28437 9512
rect 28395 9463 28437 9472
rect 28587 9512 28629 9521
rect 28587 9472 28588 9512
rect 28628 9472 28629 9512
rect 28587 9463 28629 9472
rect 29163 9512 29205 9521
rect 29163 9472 29164 9512
rect 29204 9472 29205 9512
rect 29163 9463 29205 9472
rect 29547 9512 29589 9521
rect 29547 9472 29548 9512
rect 29588 9472 29589 9512
rect 29547 9463 29589 9472
rect 29931 9512 29973 9521
rect 29931 9472 29932 9512
rect 29972 9472 29973 9512
rect 29931 9463 29973 9472
rect 30315 9512 30357 9521
rect 30315 9472 30316 9512
rect 30356 9472 30357 9512
rect 30315 9463 30357 9472
rect 31467 9512 31509 9521
rect 31467 9472 31468 9512
rect 31508 9472 31509 9512
rect 31467 9463 31509 9472
rect 31851 9512 31893 9521
rect 31851 9472 31852 9512
rect 31892 9472 31893 9512
rect 31851 9463 31893 9472
rect 32235 9512 32277 9521
rect 32235 9472 32236 9512
rect 32276 9472 32277 9512
rect 32235 9463 32277 9472
rect 32619 9512 32661 9521
rect 32619 9472 32620 9512
rect 32660 9472 32661 9512
rect 32619 9463 32661 9472
rect 33003 9512 33045 9521
rect 33003 9472 33004 9512
rect 33044 9472 33045 9512
rect 33003 9463 33045 9472
rect 33387 9512 33429 9521
rect 33387 9472 33388 9512
rect 33428 9472 33429 9512
rect 33387 9463 33429 9472
rect 33771 9512 33813 9521
rect 33771 9472 33772 9512
rect 33812 9472 33813 9512
rect 33771 9463 33813 9472
rect 34155 9512 34197 9521
rect 34155 9472 34156 9512
rect 34196 9472 34197 9512
rect 34155 9463 34197 9472
rect 34539 9512 34581 9521
rect 34539 9472 34540 9512
rect 34580 9472 34581 9512
rect 34539 9463 34581 9472
rect 34923 9512 34965 9521
rect 34923 9472 34924 9512
rect 34964 9472 34965 9512
rect 34923 9463 34965 9472
rect 35307 9512 35349 9521
rect 35307 9472 35308 9512
rect 35348 9472 35349 9512
rect 35307 9463 35349 9472
rect 35691 9512 35733 9521
rect 35691 9472 35692 9512
rect 35732 9472 35733 9512
rect 35691 9463 35733 9472
rect 36075 9512 36117 9521
rect 36075 9472 36076 9512
rect 36116 9472 36117 9512
rect 36075 9463 36117 9472
rect 42219 9512 42261 9521
rect 42219 9472 42220 9512
rect 42260 9472 42261 9512
rect 42219 9463 42261 9472
rect 42603 9512 42645 9521
rect 42603 9472 42604 9512
rect 42644 9472 42645 9512
rect 42603 9463 42645 9472
rect 43083 9512 43125 9521
rect 43083 9472 43084 9512
rect 43124 9472 43125 9512
rect 43083 9463 43125 9472
rect 43467 9512 43509 9521
rect 43467 9472 43468 9512
rect 43508 9472 43509 9512
rect 43467 9463 43509 9472
rect 43755 9512 43797 9521
rect 43755 9472 43756 9512
rect 43796 9472 43797 9512
rect 43755 9463 43797 9472
rect 44139 9512 44181 9521
rect 44139 9472 44140 9512
rect 44180 9472 44181 9512
rect 44139 9463 44181 9472
rect 44523 9512 44565 9521
rect 44523 9472 44524 9512
rect 44564 9472 44565 9512
rect 44523 9463 44565 9472
rect 44907 9512 44949 9521
rect 44907 9472 44908 9512
rect 44948 9472 44949 9512
rect 44907 9463 44949 9472
rect 2619 9344 2661 9353
rect 2619 9304 2620 9344
rect 2660 9304 2661 9344
rect 2619 9295 2661 9304
rect 3003 9344 3045 9353
rect 3003 9304 3004 9344
rect 3044 9304 3045 9344
rect 3003 9295 3045 9304
rect 10971 9344 11013 9353
rect 10971 9304 10972 9344
rect 11012 9304 11013 9344
rect 10971 9295 11013 9304
rect 19419 9344 19461 9353
rect 19419 9304 19420 9344
rect 19460 9304 19461 9344
rect 19419 9295 19461 9304
rect 22491 9344 22533 9353
rect 22491 9304 22492 9344
rect 22532 9304 22533 9344
rect 22491 9295 22533 9304
rect 23451 9344 23493 9353
rect 23451 9304 23452 9344
rect 23492 9304 23493 9344
rect 23451 9295 23493 9304
rect 23835 9344 23877 9353
rect 23835 9304 23836 9344
rect 23876 9304 23877 9344
rect 23835 9295 23877 9304
rect 24987 9344 25029 9353
rect 24987 9304 24988 9344
rect 25028 9304 25029 9344
rect 24987 9295 25029 9304
rect 25371 9344 25413 9353
rect 25371 9304 25372 9344
rect 25412 9304 25413 9344
rect 25371 9295 25413 9304
rect 26523 9344 26565 9353
rect 26523 9304 26524 9344
rect 26564 9304 26565 9344
rect 26523 9295 26565 9304
rect 27291 9344 27333 9353
rect 27291 9304 27292 9344
rect 27332 9304 27333 9344
rect 27291 9295 27333 9304
rect 32763 9344 32805 9353
rect 32763 9304 32764 9344
rect 32804 9304 32805 9344
rect 32763 9295 32805 9304
rect 33147 9344 33189 9353
rect 33147 9304 33148 9344
rect 33188 9304 33189 9344
rect 33147 9295 33189 9304
rect 35067 9344 35109 9353
rect 35067 9304 35068 9344
rect 35108 9304 35109 9344
rect 35067 9295 35109 9304
rect 45147 9344 45189 9353
rect 45147 9304 45148 9344
rect 45188 9304 45189 9344
rect 45147 9295 45189 9304
rect 1467 9260 1509 9269
rect 1467 9220 1468 9260
rect 1508 9220 1509 9260
rect 1467 9211 1509 9220
rect 1851 9260 1893 9269
rect 1851 9220 1852 9260
rect 1892 9220 1893 9260
rect 1851 9211 1893 9220
rect 3387 9260 3429 9269
rect 3387 9220 3388 9260
rect 3428 9220 3429 9260
rect 3387 9211 3429 9220
rect 20667 9260 20709 9269
rect 20667 9220 20668 9260
rect 20708 9220 20709 9260
rect 20667 9211 20709 9220
rect 21435 9260 21477 9269
rect 21435 9220 21436 9260
rect 21476 9220 21477 9260
rect 21435 9211 21477 9220
rect 22107 9260 22149 9269
rect 22107 9220 22108 9260
rect 22148 9220 22149 9260
rect 22107 9211 22149 9220
rect 22587 9260 22629 9269
rect 22587 9220 22588 9260
rect 22628 9220 22629 9260
rect 22587 9211 22629 9220
rect 23931 9260 23973 9269
rect 23931 9220 23932 9260
rect 23972 9220 23973 9260
rect 23931 9211 23973 9220
rect 24315 9260 24357 9269
rect 24315 9220 24316 9260
rect 24356 9220 24357 9260
rect 24315 9211 24357 9220
rect 25467 9260 25509 9269
rect 25467 9220 25468 9260
rect 25508 9220 25509 9260
rect 25467 9211 25509 9220
rect 26619 9260 26661 9269
rect 26619 9220 26620 9260
rect 26660 9220 26661 9260
rect 26619 9211 26661 9220
rect 28155 9260 28197 9269
rect 28155 9220 28156 9260
rect 28196 9220 28197 9260
rect 28155 9211 28197 9220
rect 28923 9260 28965 9269
rect 28923 9220 28924 9260
rect 28964 9220 28965 9260
rect 28923 9211 28965 9220
rect 29307 9260 29349 9269
rect 29307 9220 29308 9260
rect 29348 9220 29349 9260
rect 29307 9211 29349 9220
rect 29691 9260 29733 9269
rect 29691 9220 29692 9260
rect 29732 9220 29733 9260
rect 29691 9211 29733 9220
rect 30075 9260 30117 9269
rect 30075 9220 30076 9260
rect 30116 9220 30117 9260
rect 30075 9211 30117 9220
rect 33915 9260 33957 9269
rect 33915 9220 33916 9260
rect 33956 9220 33957 9260
rect 33915 9211 33957 9220
rect 41914 9260 41972 9261
rect 41914 9220 41923 9260
rect 41963 9220 41972 9260
rect 41914 9219 41972 9220
rect 42459 9260 42501 9269
rect 42459 9220 42460 9260
rect 42500 9220 42501 9260
rect 42459 9211 42501 9220
rect 43323 9260 43365 9269
rect 43323 9220 43324 9260
rect 43364 9220 43365 9260
rect 43323 9211 43365 9220
rect 43450 9260 43508 9261
rect 43450 9220 43459 9260
rect 43499 9220 43508 9260
rect 43450 9219 43508 9220
rect 1152 9092 45216 9116
rect 1152 9052 4928 9092
rect 4968 9052 5010 9092
rect 5050 9052 5092 9092
rect 5132 9052 5174 9092
rect 5214 9052 5256 9092
rect 5296 9052 20048 9092
rect 20088 9052 20130 9092
rect 20170 9052 20212 9092
rect 20252 9052 20294 9092
rect 20334 9052 20376 9092
rect 20416 9052 35168 9092
rect 35208 9052 35250 9092
rect 35290 9052 35332 9092
rect 35372 9052 35414 9092
rect 35454 9052 35496 9092
rect 35536 9052 45216 9092
rect 1152 9028 45216 9052
rect 1467 8924 1509 8933
rect 1467 8884 1468 8924
rect 1508 8884 1509 8924
rect 1467 8875 1509 8884
rect 9915 8924 9957 8933
rect 9915 8884 9916 8924
rect 9956 8884 9957 8924
rect 9915 8875 9957 8884
rect 10683 8924 10725 8933
rect 10683 8884 10684 8924
rect 10724 8884 10725 8924
rect 10683 8875 10725 8884
rect 11451 8924 11493 8933
rect 11451 8884 11452 8924
rect 11492 8884 11493 8924
rect 11451 8875 11493 8884
rect 11914 8924 11972 8925
rect 11914 8884 11923 8924
rect 11963 8884 11972 8924
rect 11914 8883 11972 8884
rect 12219 8924 12261 8933
rect 12219 8884 12220 8924
rect 12260 8884 12261 8924
rect 12219 8875 12261 8884
rect 12603 8924 12645 8933
rect 12603 8884 12604 8924
rect 12644 8884 12645 8924
rect 12603 8875 12645 8884
rect 12987 8924 13029 8933
rect 12987 8884 12988 8924
rect 13028 8884 13029 8924
rect 12987 8875 13029 8884
rect 13371 8924 13413 8933
rect 13371 8884 13372 8924
rect 13412 8884 13413 8924
rect 13371 8875 13413 8884
rect 13755 8924 13797 8933
rect 13755 8884 13756 8924
rect 13796 8884 13797 8924
rect 13755 8875 13797 8884
rect 14523 8924 14565 8933
rect 14523 8884 14524 8924
rect 14564 8884 14565 8924
rect 14523 8875 14565 8884
rect 15291 8924 15333 8933
rect 15291 8884 15292 8924
rect 15332 8884 15333 8924
rect 15291 8875 15333 8884
rect 15675 8924 15717 8933
rect 15675 8884 15676 8924
rect 15716 8884 15717 8924
rect 15675 8875 15717 8884
rect 16059 8924 16101 8933
rect 16059 8884 16060 8924
rect 16100 8884 16101 8924
rect 16059 8875 16101 8884
rect 16443 8924 16485 8933
rect 16443 8884 16444 8924
rect 16484 8884 16485 8924
rect 16443 8875 16485 8884
rect 16827 8924 16869 8933
rect 16827 8884 16828 8924
rect 16868 8884 16869 8924
rect 16827 8875 16869 8884
rect 17211 8924 17253 8933
rect 17211 8884 17212 8924
rect 17252 8884 17253 8924
rect 17211 8875 17253 8884
rect 17595 8924 17637 8933
rect 17595 8884 17596 8924
rect 17636 8884 17637 8924
rect 17595 8875 17637 8884
rect 17979 8924 18021 8933
rect 17979 8884 17980 8924
rect 18020 8884 18021 8924
rect 17979 8875 18021 8884
rect 18363 8924 18405 8933
rect 18363 8884 18364 8924
rect 18404 8884 18405 8924
rect 18363 8875 18405 8884
rect 18747 8924 18789 8933
rect 18747 8884 18748 8924
rect 18788 8884 18789 8924
rect 18747 8875 18789 8884
rect 19131 8924 19173 8933
rect 19131 8884 19132 8924
rect 19172 8884 19173 8924
rect 19131 8875 19173 8884
rect 19515 8924 19557 8933
rect 19515 8884 19516 8924
rect 19556 8884 19557 8924
rect 19515 8875 19557 8884
rect 20283 8924 20325 8933
rect 20283 8884 20284 8924
rect 20324 8884 20325 8924
rect 20283 8875 20325 8884
rect 21099 8924 21141 8933
rect 21099 8884 21100 8924
rect 21140 8884 21141 8924
rect 21099 8875 21141 8884
rect 32187 8924 32229 8933
rect 32187 8884 32188 8924
rect 32228 8884 32229 8924
rect 32187 8875 32229 8884
rect 32571 8924 32613 8933
rect 32571 8884 32572 8924
rect 32612 8884 32613 8924
rect 32571 8875 32613 8884
rect 32955 8924 32997 8933
rect 32955 8884 32956 8924
rect 32996 8884 32997 8924
rect 32955 8875 32997 8884
rect 33339 8924 33381 8933
rect 33339 8884 33340 8924
rect 33380 8884 33381 8924
rect 33339 8875 33381 8884
rect 33723 8924 33765 8933
rect 33723 8884 33724 8924
rect 33764 8884 33765 8924
rect 33723 8875 33765 8884
rect 34107 8924 34149 8933
rect 34107 8884 34108 8924
rect 34148 8884 34149 8924
rect 34107 8875 34149 8884
rect 34875 8924 34917 8933
rect 34875 8884 34876 8924
rect 34916 8884 34917 8924
rect 34875 8875 34917 8884
rect 43515 8924 43557 8933
rect 43515 8884 43516 8924
rect 43556 8884 43557 8924
rect 43515 8875 43557 8884
rect 44379 8924 44421 8933
rect 44379 8884 44380 8924
rect 44420 8884 44421 8924
rect 44379 8875 44421 8884
rect 10299 8840 10341 8849
rect 10299 8800 10300 8840
rect 10340 8800 10341 8840
rect 10299 8791 10341 8800
rect 20667 8840 20709 8849
rect 20667 8800 20668 8840
rect 20708 8800 20709 8840
rect 20667 8791 20709 8800
rect 21723 8840 21765 8849
rect 21723 8800 21724 8840
rect 21764 8800 21765 8840
rect 21723 8791 21765 8800
rect 23547 8840 23589 8849
rect 23547 8800 23548 8840
rect 23588 8800 23589 8840
rect 23547 8791 23589 8800
rect 25659 8840 25701 8849
rect 25659 8800 25660 8840
rect 25700 8800 25701 8840
rect 25659 8791 25701 8800
rect 28251 8840 28293 8849
rect 28251 8800 28252 8840
rect 28292 8800 28293 8840
rect 28251 8791 28293 8800
rect 29403 8840 29445 8849
rect 29403 8800 29404 8840
rect 29444 8800 29445 8840
rect 29403 8791 29445 8800
rect 34491 8840 34533 8849
rect 34491 8800 34492 8840
rect 34532 8800 34533 8840
rect 34491 8791 34533 8800
rect 42363 8840 42405 8849
rect 42363 8800 42364 8840
rect 42404 8800 42405 8840
rect 42363 8791 42405 8800
rect 42747 8840 42789 8849
rect 42747 8800 42748 8840
rect 42788 8800 42789 8840
rect 42747 8791 42789 8800
rect 11595 8756 11637 8765
rect 11595 8716 11596 8756
rect 11636 8716 11637 8756
rect 27627 8756 27669 8765
rect 11595 8707 11637 8716
rect 11723 8732 11765 8741
rect 11723 8692 11724 8732
rect 11764 8692 11765 8732
rect 27627 8716 27628 8756
rect 27668 8716 27669 8756
rect 27627 8707 27669 8716
rect 27748 8756 27806 8757
rect 27748 8716 27757 8756
rect 27797 8716 27806 8756
rect 27748 8715 27806 8716
rect 28011 8756 28053 8765
rect 28011 8716 28012 8756
rect 28052 8716 28053 8756
rect 28011 8707 28053 8716
rect 11723 8683 11765 8692
rect 1227 8672 1269 8681
rect 1227 8632 1228 8672
rect 1268 8632 1269 8672
rect 1227 8623 1269 8632
rect 1611 8672 1653 8681
rect 1611 8632 1612 8672
rect 1652 8632 1653 8672
rect 1611 8623 1653 8632
rect 1851 8672 1893 8681
rect 1851 8632 1852 8672
rect 1892 8632 1893 8672
rect 1851 8623 1893 8632
rect 1995 8672 2037 8681
rect 1995 8632 1996 8672
rect 2036 8632 2037 8672
rect 1995 8623 2037 8632
rect 2235 8672 2277 8681
rect 2235 8632 2236 8672
rect 2276 8632 2277 8672
rect 2235 8623 2277 8632
rect 2379 8672 2421 8681
rect 2379 8632 2380 8672
rect 2420 8632 2421 8672
rect 2379 8623 2421 8632
rect 2619 8672 2661 8681
rect 2619 8632 2620 8672
rect 2660 8632 2661 8672
rect 2619 8623 2661 8632
rect 9675 8672 9717 8681
rect 9675 8632 9676 8672
rect 9716 8632 9717 8672
rect 9675 8623 9717 8632
rect 10059 8672 10101 8681
rect 10059 8632 10060 8672
rect 10100 8632 10101 8672
rect 10059 8623 10101 8632
rect 10443 8672 10485 8681
rect 10443 8632 10444 8672
rect 10484 8632 10485 8672
rect 10443 8623 10485 8632
rect 10827 8672 10869 8681
rect 10827 8632 10828 8672
rect 10868 8632 10869 8672
rect 10827 8623 10869 8632
rect 11211 8672 11253 8681
rect 11211 8632 11212 8672
rect 11252 8632 11253 8672
rect 11211 8623 11253 8632
rect 12459 8672 12501 8681
rect 12459 8632 12460 8672
rect 12500 8632 12501 8672
rect 12459 8623 12501 8632
rect 12843 8672 12885 8681
rect 12843 8632 12844 8672
rect 12884 8632 12885 8672
rect 12843 8623 12885 8632
rect 13227 8672 13269 8681
rect 13227 8632 13228 8672
rect 13268 8632 13269 8672
rect 13227 8623 13269 8632
rect 13611 8672 13653 8681
rect 13611 8632 13612 8672
rect 13652 8632 13653 8672
rect 13611 8623 13653 8632
rect 13995 8672 14037 8681
rect 13995 8632 13996 8672
rect 14036 8632 14037 8672
rect 13995 8623 14037 8632
rect 14379 8672 14421 8681
rect 14379 8632 14380 8672
rect 14420 8632 14421 8672
rect 14379 8623 14421 8632
rect 14763 8672 14805 8681
rect 14763 8632 14764 8672
rect 14804 8632 14805 8672
rect 14763 8623 14805 8632
rect 14955 8672 14997 8681
rect 14955 8632 14956 8672
rect 14996 8632 14997 8672
rect 14955 8623 14997 8632
rect 15195 8672 15237 8681
rect 15195 8632 15196 8672
rect 15236 8632 15237 8672
rect 15195 8623 15237 8632
rect 15531 8672 15573 8681
rect 15531 8632 15532 8672
rect 15572 8632 15573 8672
rect 15531 8623 15573 8632
rect 15915 8672 15957 8681
rect 15915 8632 15916 8672
rect 15956 8632 15957 8672
rect 15915 8623 15957 8632
rect 16299 8672 16341 8681
rect 16299 8632 16300 8672
rect 16340 8632 16341 8672
rect 16299 8623 16341 8632
rect 16683 8672 16725 8681
rect 16683 8632 16684 8672
rect 16724 8632 16725 8672
rect 16683 8623 16725 8632
rect 17067 8672 17109 8681
rect 17067 8632 17068 8672
rect 17108 8632 17109 8672
rect 17067 8623 17109 8632
rect 17451 8672 17493 8681
rect 17451 8632 17452 8672
rect 17492 8632 17493 8672
rect 17451 8623 17493 8632
rect 17835 8672 17877 8681
rect 17835 8632 17836 8672
rect 17876 8632 17877 8672
rect 17835 8623 17877 8632
rect 18219 8672 18261 8681
rect 18219 8632 18220 8672
rect 18260 8632 18261 8672
rect 18219 8623 18261 8632
rect 18603 8672 18645 8681
rect 18603 8632 18604 8672
rect 18644 8632 18645 8672
rect 18603 8623 18645 8632
rect 18987 8672 19029 8681
rect 18987 8632 18988 8672
rect 19028 8632 19029 8672
rect 18987 8623 19029 8632
rect 19371 8672 19413 8681
rect 19371 8632 19372 8672
rect 19412 8632 19413 8672
rect 19371 8623 19413 8632
rect 19755 8672 19797 8681
rect 19755 8632 19756 8672
rect 19796 8632 19797 8672
rect 19755 8623 19797 8632
rect 19899 8672 19941 8681
rect 19899 8632 19900 8672
rect 19940 8632 19941 8672
rect 19899 8623 19941 8632
rect 20139 8672 20181 8681
rect 20139 8632 20140 8672
rect 20180 8632 20181 8672
rect 20139 8623 20181 8632
rect 20523 8672 20565 8681
rect 20523 8632 20524 8672
rect 20564 8632 20565 8672
rect 20523 8623 20565 8632
rect 20907 8672 20949 8681
rect 20907 8632 20908 8672
rect 20948 8632 20949 8672
rect 20907 8623 20949 8632
rect 21483 8672 21525 8681
rect 21483 8632 21484 8672
rect 21524 8632 21525 8672
rect 21483 8623 21525 8632
rect 22059 8672 22101 8681
rect 22059 8632 22060 8672
rect 22100 8632 22101 8672
rect 22059 8623 22101 8632
rect 23787 8672 23829 8681
rect 23787 8632 23788 8672
rect 23828 8632 23829 8672
rect 23787 8623 23829 8632
rect 25323 8672 25365 8681
rect 25323 8632 25324 8672
rect 25364 8632 25365 8672
rect 25323 8623 25365 8632
rect 25899 8672 25941 8681
rect 25899 8632 25900 8672
rect 25940 8632 25941 8672
rect 25899 8623 25941 8632
rect 26091 8672 26133 8681
rect 26091 8632 26092 8672
rect 26132 8632 26133 8672
rect 26091 8623 26133 8632
rect 26427 8672 26469 8681
rect 26427 8632 26428 8672
rect 26468 8632 26469 8672
rect 26427 8623 26469 8632
rect 26667 8672 26709 8681
rect 26667 8632 26668 8672
rect 26708 8632 26709 8672
rect 26667 8623 26709 8632
rect 26811 8672 26853 8681
rect 26811 8632 26812 8672
rect 26852 8632 26853 8672
rect 26811 8623 26853 8632
rect 27051 8672 27093 8681
rect 27051 8632 27052 8672
rect 27092 8632 27093 8672
rect 27051 8623 27093 8632
rect 28491 8672 28533 8681
rect 28491 8632 28492 8672
rect 28532 8632 28533 8672
rect 28491 8623 28533 8632
rect 29163 8672 29205 8681
rect 29163 8632 29164 8672
rect 29204 8632 29205 8672
rect 29163 8623 29205 8632
rect 29739 8672 29781 8681
rect 29739 8632 29740 8672
rect 29780 8632 29781 8672
rect 29739 8623 29781 8632
rect 32427 8672 32469 8681
rect 32427 8632 32428 8672
rect 32468 8632 32469 8672
rect 32427 8623 32469 8632
rect 32811 8672 32853 8681
rect 32811 8632 32812 8672
rect 32852 8632 32853 8672
rect 32811 8623 32853 8632
rect 33195 8672 33237 8681
rect 33195 8632 33196 8672
rect 33236 8632 33237 8672
rect 33195 8623 33237 8632
rect 33579 8672 33621 8681
rect 33579 8632 33580 8672
rect 33620 8632 33621 8672
rect 33579 8623 33621 8632
rect 33963 8672 34005 8681
rect 33963 8632 33964 8672
rect 34004 8632 34005 8672
rect 33963 8623 34005 8632
rect 34347 8672 34389 8681
rect 34347 8632 34348 8672
rect 34388 8632 34389 8672
rect 34347 8623 34389 8632
rect 34731 8672 34773 8681
rect 34731 8632 34732 8672
rect 34772 8632 34773 8672
rect 34731 8623 34773 8632
rect 35115 8672 35157 8681
rect 35115 8632 35116 8672
rect 35156 8632 35157 8672
rect 35115 8623 35157 8632
rect 42603 8672 42645 8681
rect 42603 8632 42604 8672
rect 42644 8632 42645 8672
rect 42603 8623 42645 8632
rect 42987 8672 43029 8681
rect 42987 8632 42988 8672
rect 43028 8632 43029 8672
rect 42987 8623 43029 8632
rect 43131 8672 43173 8681
rect 43131 8632 43132 8672
rect 43172 8632 43173 8672
rect 43131 8623 43173 8632
rect 43371 8672 43413 8681
rect 43371 8632 43372 8672
rect 43412 8632 43413 8672
rect 43371 8623 43413 8632
rect 43755 8672 43797 8681
rect 43755 8632 43756 8672
rect 43796 8632 43797 8672
rect 43755 8623 43797 8632
rect 44139 8672 44181 8681
rect 44139 8632 44140 8672
rect 44180 8632 44181 8672
rect 44139 8623 44181 8632
rect 44523 8672 44565 8681
rect 44523 8632 44524 8672
rect 44564 8632 44565 8672
rect 44523 8623 44565 8632
rect 44907 8672 44949 8681
rect 44907 8632 44908 8672
rect 44948 8632 44949 8672
rect 44907 8623 44949 8632
rect 11067 8588 11109 8597
rect 11067 8548 11068 8588
rect 11108 8548 11109 8588
rect 11067 8539 11109 8548
rect 21819 8588 21861 8597
rect 21819 8548 21820 8588
rect 21860 8548 21861 8588
rect 21819 8539 21861 8548
rect 25563 8588 25605 8597
rect 25563 8548 25564 8588
rect 25604 8548 25605 8588
rect 25563 8539 25605 8548
rect 26331 8588 26373 8597
rect 26331 8548 26332 8588
rect 26372 8548 26373 8588
rect 26331 8539 26373 8548
rect 14139 8504 14181 8513
rect 14139 8464 14140 8504
rect 14180 8464 14181 8504
rect 14139 8455 14181 8464
rect 27339 8504 27381 8513
rect 27339 8464 27340 8504
rect 27380 8464 27381 8504
rect 27339 8455 27381 8464
rect 29499 8504 29541 8513
rect 29499 8464 29500 8504
rect 29540 8464 29541 8504
rect 29499 8455 29541 8464
rect 44763 8504 44805 8513
rect 44763 8464 44764 8504
rect 44804 8464 44805 8504
rect 44763 8455 44805 8464
rect 45147 8504 45189 8513
rect 45147 8464 45148 8504
rect 45188 8464 45189 8504
rect 45147 8455 45189 8464
rect 1152 8336 45216 8360
rect 1152 8296 3688 8336
rect 3728 8296 3770 8336
rect 3810 8296 3852 8336
rect 3892 8296 3934 8336
rect 3974 8296 4016 8336
rect 4056 8296 18808 8336
rect 18848 8296 18890 8336
rect 18930 8296 18972 8336
rect 19012 8296 19054 8336
rect 19094 8296 19136 8336
rect 19176 8296 33928 8336
rect 33968 8296 34010 8336
rect 34050 8296 34092 8336
rect 34132 8296 34174 8336
rect 34214 8296 34256 8336
rect 34296 8296 45216 8336
rect 1152 8272 45216 8296
rect 17883 8168 17925 8177
rect 17883 8128 17884 8168
rect 17924 8128 17925 8168
rect 17883 8119 17925 8128
rect 22875 8168 22917 8177
rect 22875 8128 22876 8168
rect 22916 8128 22917 8168
rect 22875 8119 22917 8128
rect 28251 8168 28293 8177
rect 28251 8128 28252 8168
rect 28292 8128 28293 8168
rect 28251 8119 28293 8128
rect 28635 8168 28677 8177
rect 28635 8128 28636 8168
rect 28676 8128 28677 8168
rect 28635 8119 28677 8128
rect 32091 8168 32133 8177
rect 32091 8128 32092 8168
rect 32132 8128 32133 8168
rect 32091 8119 32133 8128
rect 34491 8168 34533 8177
rect 34491 8128 34492 8168
rect 34532 8128 34533 8168
rect 34491 8119 34533 8128
rect 34971 8168 35013 8177
rect 34971 8128 34972 8168
rect 35012 8128 35013 8168
rect 34971 8119 35013 8128
rect 36699 8168 36741 8177
rect 36699 8128 36700 8168
rect 36740 8128 36741 8168
rect 36699 8119 36741 8128
rect 42747 8168 42789 8177
rect 42747 8128 42748 8168
rect 42788 8128 42789 8168
rect 42747 8119 42789 8128
rect 43131 8168 43173 8177
rect 43131 8128 43132 8168
rect 43172 8128 43173 8168
rect 43131 8119 43173 8128
rect 43899 8168 43941 8177
rect 43899 8128 43900 8168
rect 43940 8128 43941 8168
rect 43899 8119 43941 8128
rect 24843 8084 24885 8093
rect 24843 8044 24844 8084
rect 24884 8044 24885 8084
rect 24843 8035 24885 8044
rect 34875 8084 34917 8093
rect 34875 8044 34876 8084
rect 34916 8044 34917 8084
rect 34875 8035 34917 8044
rect 1227 8000 1269 8009
rect 1227 7960 1228 8000
rect 1268 7960 1269 8000
rect 1227 7951 1269 7960
rect 1611 8000 1653 8009
rect 1611 7960 1612 8000
rect 1652 7960 1653 8000
rect 1611 7951 1653 7960
rect 2475 8000 2517 8009
rect 2475 7960 2476 8000
rect 2516 7960 2517 8000
rect 2475 7951 2517 7960
rect 2715 8000 2757 8009
rect 2715 7960 2716 8000
rect 2756 7960 2757 8000
rect 2715 7951 2757 7960
rect 2859 8000 2901 8009
rect 2859 7960 2860 8000
rect 2900 7960 2901 8000
rect 2859 7951 2901 7960
rect 3243 8000 3285 8009
rect 3243 7960 3244 8000
rect 3284 7960 3285 8000
rect 3243 7951 3285 7960
rect 3483 8000 3525 8009
rect 3483 7960 3484 8000
rect 3524 7960 3525 8000
rect 3483 7951 3525 7960
rect 3627 8000 3669 8009
rect 3627 7960 3628 8000
rect 3668 7960 3669 8000
rect 3627 7951 3669 7960
rect 4011 8000 4053 8009
rect 4011 7960 4012 8000
rect 4052 7960 4053 8000
rect 4011 7951 4053 7960
rect 4395 8000 4437 8009
rect 4395 7960 4396 8000
rect 4436 7960 4437 8000
rect 4395 7951 4437 7960
rect 10251 8000 10293 8009
rect 10251 7960 10252 8000
rect 10292 7960 10293 8000
rect 10251 7951 10293 7960
rect 14475 8000 14517 8009
rect 14475 7960 14476 8000
rect 14516 7960 14517 8000
rect 14475 7951 14517 7960
rect 16971 8000 17013 8009
rect 16971 7960 16972 8000
rect 17012 7960 17013 8000
rect 16971 7951 17013 7960
rect 18123 8000 18165 8009
rect 18123 7960 18124 8000
rect 18164 7960 18165 8000
rect 18123 7951 18165 7960
rect 22635 8000 22677 8009
rect 22635 7960 22636 8000
rect 22676 7960 22677 8000
rect 22635 7951 22677 7960
rect 23019 8000 23061 8009
rect 23019 7960 23020 8000
rect 23060 7960 23061 8000
rect 23019 7951 23061 7960
rect 26091 8000 26133 8009
rect 26091 7960 26092 8000
rect 26132 7960 26133 8000
rect 26091 7951 26133 7960
rect 26859 8000 26901 8009
rect 26859 7960 26860 8000
rect 26900 7960 26901 8000
rect 26859 7951 26901 7960
rect 28491 8000 28533 8009
rect 28491 7960 28492 8000
rect 28532 7960 28533 8000
rect 28491 7951 28533 7960
rect 28875 8000 28917 8009
rect 28875 7960 28876 8000
rect 28916 7960 28917 8000
rect 28875 7951 28917 7960
rect 29451 8000 29493 8009
rect 29451 7960 29452 8000
rect 29492 7960 29493 8000
rect 29451 7951 29493 7960
rect 31563 8000 31605 8009
rect 31563 7960 31564 8000
rect 31604 7960 31605 8000
rect 31563 7951 31605 7960
rect 31851 8000 31893 8009
rect 31851 7960 31852 8000
rect 31892 7960 31893 8000
rect 31851 7951 31893 7960
rect 32427 8000 32469 8009
rect 32427 7960 32428 8000
rect 32468 7960 32469 8000
rect 32427 7951 32469 7960
rect 32715 8000 32757 8009
rect 32715 7960 32716 8000
rect 32756 7960 32757 8000
rect 32715 7951 32757 7960
rect 33195 8000 33237 8009
rect 33195 7960 33196 8000
rect 33236 7960 33237 8000
rect 33195 7951 33237 7960
rect 33483 8000 33525 8009
rect 33483 7960 33484 8000
rect 33524 7960 33525 8000
rect 33483 7951 33525 7960
rect 33867 8000 33909 8009
rect 33867 7960 33868 8000
rect 33908 7960 33909 8000
rect 33867 7951 33909 7960
rect 34251 8000 34293 8009
rect 34251 7960 34252 8000
rect 34292 7960 34293 8000
rect 34251 7951 34293 7960
rect 34635 8000 34677 8009
rect 34635 7960 34636 8000
rect 34676 7960 34677 8000
rect 34635 7951 34677 7960
rect 35211 8000 35253 8009
rect 35211 7960 35212 8000
rect 35252 7960 35253 8000
rect 35211 7951 35253 7960
rect 36490 8000 36548 8001
rect 36490 7960 36499 8000
rect 36539 7960 36548 8000
rect 36490 7959 36548 7960
rect 41835 8000 41877 8009
rect 41835 7960 41836 8000
rect 41876 7960 41877 8000
rect 41835 7951 41877 7960
rect 41979 8000 42021 8009
rect 41979 7960 41980 8000
rect 42020 7960 42021 8000
rect 41979 7951 42021 7960
rect 42219 8000 42261 8009
rect 42219 7960 42220 8000
rect 42260 7960 42261 8000
rect 42219 7951 42261 7960
rect 42603 8000 42645 8009
rect 42603 7960 42604 8000
rect 42644 7960 42645 8000
rect 42603 7951 42645 7960
rect 42987 8000 43029 8009
rect 42987 7960 42988 8000
rect 43028 7960 43029 8000
rect 42987 7951 43029 7960
rect 43371 8000 43413 8009
rect 43371 7960 43372 8000
rect 43412 7960 43413 8000
rect 43371 7951 43413 7960
rect 43755 8000 43797 8009
rect 43755 7960 43756 8000
rect 43796 7960 43797 8000
rect 43755 7951 43797 7960
rect 44139 8000 44181 8009
rect 44139 7960 44140 8000
rect 44180 7960 44181 8000
rect 44139 7951 44181 7960
rect 44523 8000 44565 8009
rect 44523 7960 44524 8000
rect 44564 7960 44565 8000
rect 44523 7951 44565 7960
rect 44907 8000 44949 8009
rect 44907 7960 44908 8000
rect 44948 7960 44949 8000
rect 44907 7951 44949 7960
rect 9754 7916 9812 7917
rect 9754 7876 9763 7916
rect 9803 7876 9812 7916
rect 9754 7875 9812 7876
rect 9867 7916 9909 7925
rect 9867 7876 9868 7916
rect 9908 7876 9909 7916
rect 9867 7867 9909 7876
rect 10347 7916 10389 7925
rect 10347 7876 10348 7916
rect 10388 7876 10389 7916
rect 10347 7867 10389 7876
rect 10819 7916 10877 7917
rect 10819 7876 10828 7916
rect 10868 7876 10877 7916
rect 10819 7875 10877 7876
rect 11307 7916 11365 7917
rect 11307 7876 11316 7916
rect 11356 7876 11365 7916
rect 11307 7875 11365 7876
rect 11787 7916 11829 7925
rect 11787 7876 11788 7916
rect 11828 7876 11829 7916
rect 11787 7867 11829 7876
rect 12058 7916 12116 7917
rect 12058 7876 12067 7916
rect 12107 7876 12116 7916
rect 12058 7875 12116 7876
rect 12603 7916 12645 7925
rect 12603 7876 12604 7916
rect 12644 7876 12645 7916
rect 12603 7867 12645 7876
rect 12747 7916 12789 7925
rect 12747 7876 12748 7916
rect 12788 7876 12789 7916
rect 12747 7867 12789 7876
rect 14859 7916 14901 7925
rect 14859 7876 14860 7916
rect 14900 7876 14901 7916
rect 14859 7867 14901 7876
rect 16099 7916 16157 7917
rect 16099 7876 16108 7916
rect 16148 7876 16157 7916
rect 16099 7875 16157 7876
rect 23403 7916 23445 7925
rect 23403 7876 23404 7916
rect 23444 7876 23445 7916
rect 23403 7867 23445 7876
rect 24643 7916 24701 7917
rect 24643 7876 24652 7916
rect 24692 7876 24701 7916
rect 24643 7875 24701 7876
rect 26362 7916 26420 7917
rect 26362 7876 26371 7916
rect 26411 7876 26420 7916
rect 26362 7875 26420 7876
rect 26475 7916 26517 7925
rect 26475 7876 26476 7916
rect 26516 7876 26517 7916
rect 26475 7867 26517 7876
rect 26955 7916 26997 7925
rect 26955 7876 26956 7916
rect 26996 7876 26997 7916
rect 26955 7867 26997 7876
rect 27427 7916 27485 7917
rect 27427 7876 27436 7916
rect 27476 7876 27485 7916
rect 27427 7875 27485 7876
rect 27946 7916 28004 7917
rect 27946 7876 27955 7916
rect 27995 7876 28004 7916
rect 27946 7875 28004 7876
rect 1851 7832 1893 7841
rect 1851 7792 1852 7832
rect 1892 7792 1893 7832
rect 1851 7783 1893 7792
rect 3099 7832 3141 7841
rect 3099 7792 3100 7832
rect 3140 7792 3141 7832
rect 3099 7783 3141 7792
rect 12171 7832 12213 7841
rect 12171 7792 12172 7832
rect 12212 7792 12213 7832
rect 12171 7783 12213 7792
rect 41595 7832 41637 7841
rect 41595 7792 41596 7832
rect 41636 7792 41637 7832
rect 41595 7783 41637 7792
rect 43515 7832 43557 7841
rect 43515 7792 43516 7832
rect 43556 7792 43557 7832
rect 43515 7783 43557 7792
rect 1467 7748 1509 7757
rect 1467 7708 1468 7748
rect 1508 7708 1509 7748
rect 1467 7699 1509 7708
rect 3867 7748 3909 7757
rect 3867 7708 3868 7748
rect 3908 7708 3909 7748
rect 3867 7699 3909 7708
rect 4251 7748 4293 7757
rect 4251 7708 4252 7748
rect 4292 7708 4293 7748
rect 4251 7699 4293 7708
rect 4635 7748 4677 7757
rect 4635 7708 4636 7748
rect 4676 7708 4677 7748
rect 4635 7699 4677 7708
rect 11499 7748 11541 7757
rect 11499 7708 11500 7748
rect 11540 7708 11541 7748
rect 11499 7699 11541 7708
rect 12507 7748 12549 7757
rect 12507 7708 12508 7748
rect 12548 7708 12549 7748
rect 12507 7699 12549 7708
rect 14715 7748 14757 7757
rect 14715 7708 14716 7748
rect 14756 7708 14757 7748
rect 14715 7699 14757 7708
rect 16299 7748 16341 7757
rect 16299 7708 16300 7748
rect 16340 7708 16341 7748
rect 16299 7699 16341 7708
rect 17211 7748 17253 7757
rect 17211 7708 17212 7748
rect 17252 7708 17253 7748
rect 17211 7699 17253 7708
rect 23259 7748 23301 7757
rect 23259 7708 23260 7748
rect 23300 7708 23301 7748
rect 23259 7699 23301 7708
rect 25851 7748 25893 7757
rect 25851 7708 25852 7748
rect 25892 7708 25893 7748
rect 25851 7699 25893 7708
rect 28107 7748 28149 7757
rect 28107 7708 28108 7748
rect 28148 7708 28149 7748
rect 28107 7699 28149 7708
rect 29691 7748 29733 7757
rect 29691 7708 29692 7748
rect 29732 7708 29733 7748
rect 29691 7699 29733 7708
rect 31642 7748 31700 7749
rect 31642 7708 31651 7748
rect 31691 7708 31700 7748
rect 31642 7707 31700 7708
rect 32410 7748 32468 7749
rect 32410 7708 32419 7748
rect 32459 7708 32468 7748
rect 32410 7707 32468 7708
rect 32955 7748 32997 7757
rect 32955 7708 32956 7748
rect 32996 7708 32997 7748
rect 32955 7699 32997 7708
rect 33178 7748 33236 7749
rect 33178 7708 33187 7748
rect 33227 7708 33236 7748
rect 33178 7707 33236 7708
rect 33723 7748 33765 7757
rect 33723 7708 33724 7748
rect 33764 7708 33765 7748
rect 33723 7699 33765 7708
rect 34107 7748 34149 7757
rect 34107 7708 34108 7748
rect 34148 7708 34149 7748
rect 34107 7699 34149 7708
rect 36250 7748 36308 7749
rect 36250 7708 36259 7748
rect 36299 7708 36308 7748
rect 36250 7707 36308 7708
rect 36826 7748 36884 7749
rect 36826 7708 36835 7748
rect 36875 7708 36884 7748
rect 36826 7707 36884 7708
rect 42363 7748 42405 7757
rect 42363 7708 42364 7748
rect 42404 7708 42405 7748
rect 42363 7699 42405 7708
rect 44763 7748 44805 7757
rect 44763 7708 44764 7748
rect 44804 7708 44805 7748
rect 44763 7699 44805 7708
rect 45147 7748 45189 7757
rect 45147 7708 45148 7748
rect 45188 7708 45189 7748
rect 45147 7699 45189 7708
rect 1152 7580 45216 7604
rect 1152 7540 4928 7580
rect 4968 7540 5010 7580
rect 5050 7540 5092 7580
rect 5132 7540 5174 7580
rect 5214 7540 5256 7580
rect 5296 7540 20048 7580
rect 20088 7540 20130 7580
rect 20170 7540 20212 7580
rect 20252 7540 20294 7580
rect 20334 7540 20376 7580
rect 20416 7540 35168 7580
rect 35208 7540 35250 7580
rect 35290 7540 35332 7580
rect 35372 7540 35414 7580
rect 35454 7540 35496 7580
rect 35536 7540 45216 7580
rect 1152 7516 45216 7540
rect 11770 7412 11828 7413
rect 11770 7372 11779 7412
rect 11819 7372 11828 7412
rect 11770 7371 11828 7372
rect 12538 7412 12596 7413
rect 12538 7372 12547 7412
rect 12587 7372 12596 7412
rect 12538 7371 12596 7372
rect 28011 7412 28053 7421
rect 28011 7372 28012 7412
rect 28052 7372 28053 7412
rect 28011 7363 28053 7372
rect 33082 7412 33140 7413
rect 33082 7372 33091 7412
rect 33131 7372 33140 7412
rect 33082 7371 33140 7372
rect 33370 7412 33428 7413
rect 33370 7372 33379 7412
rect 33419 7372 33428 7412
rect 33370 7371 33428 7372
rect 33946 7412 34004 7413
rect 33946 7372 33955 7412
rect 33995 7372 34004 7412
rect 33946 7371 34004 7372
rect 34522 7412 34580 7413
rect 34522 7372 34531 7412
rect 34571 7372 34580 7412
rect 34522 7371 34580 7372
rect 35098 7412 35156 7413
rect 35098 7372 35107 7412
rect 35147 7372 35156 7412
rect 35098 7371 35156 7372
rect 35674 7412 35732 7413
rect 35674 7372 35683 7412
rect 35723 7372 35732 7412
rect 35674 7371 35732 7372
rect 36154 7412 36212 7413
rect 36154 7372 36163 7412
rect 36203 7372 36212 7412
rect 36154 7371 36212 7372
rect 44026 7412 44084 7413
rect 44026 7372 44035 7412
rect 44075 7372 44084 7412
rect 44026 7371 44084 7372
rect 44619 7412 44661 7421
rect 44619 7372 44620 7412
rect 44660 7372 44661 7412
rect 44619 7363 44661 7372
rect 10539 7328 10581 7337
rect 10539 7288 10540 7328
rect 10580 7288 10581 7328
rect 10539 7279 10581 7288
rect 12651 7328 12693 7337
rect 12651 7288 12652 7328
rect 12692 7288 12693 7328
rect 12651 7279 12693 7288
rect 29163 7328 29205 7337
rect 29163 7288 29164 7328
rect 29204 7288 29205 7328
rect 29163 7279 29205 7288
rect 36747 7328 36789 7337
rect 36747 7288 36748 7328
rect 36788 7288 36789 7328
rect 36747 7279 36789 7288
rect 37611 7328 37653 7337
rect 37611 7288 37612 7328
rect 37652 7288 37653 7328
rect 37611 7279 37653 7288
rect 10155 7244 10197 7253
rect 10155 7204 10156 7244
rect 10196 7204 10197 7244
rect 10155 7195 10197 7204
rect 10426 7244 10484 7245
rect 10426 7204 10435 7244
rect 10475 7204 10484 7244
rect 11866 7244 11924 7245
rect 10426 7203 10484 7204
rect 11707 7233 11749 7242
rect 11707 7193 11708 7233
rect 11748 7193 11749 7233
rect 11866 7204 11875 7244
rect 11915 7204 11924 7244
rect 11866 7203 11924 7204
rect 11991 7244 12033 7253
rect 12442 7244 12500 7245
rect 11991 7204 11992 7244
rect 12032 7204 12033 7244
rect 11991 7195 12033 7204
rect 12123 7235 12165 7244
rect 12123 7195 12124 7235
rect 12164 7195 12165 7235
rect 11707 7184 11749 7193
rect 12123 7186 12165 7195
rect 12256 7233 12298 7242
rect 12256 7193 12257 7233
rect 12297 7193 12298 7233
rect 12442 7204 12451 7244
rect 12491 7204 12500 7244
rect 12442 7203 12500 7204
rect 12758 7244 12800 7253
rect 12758 7204 12759 7244
rect 12799 7204 12800 7244
rect 12758 7195 12800 7204
rect 13035 7244 13077 7253
rect 13035 7204 13036 7244
rect 13076 7204 13077 7244
rect 13035 7195 13077 7204
rect 14859 7244 14901 7253
rect 23307 7244 23349 7253
rect 26266 7244 26324 7245
rect 14859 7204 14860 7244
rect 14900 7204 14901 7244
rect 14859 7195 14901 7204
rect 16107 7235 16149 7244
rect 16107 7195 16108 7235
rect 16148 7195 16149 7235
rect 23307 7204 23308 7244
rect 23348 7204 23349 7244
rect 23307 7195 23349 7204
rect 24555 7235 24597 7244
rect 24555 7195 24556 7235
rect 24596 7195 24597 7235
rect 26266 7204 26275 7244
rect 26315 7204 26324 7244
rect 26266 7203 26324 7204
rect 26384 7244 26426 7253
rect 26384 7204 26385 7244
rect 26425 7204 26426 7244
rect 26384 7195 26426 7204
rect 26763 7244 26805 7253
rect 30603 7244 30645 7253
rect 26763 7204 26764 7244
rect 26804 7204 26805 7244
rect 26763 7195 26805 7204
rect 27339 7235 27381 7244
rect 27339 7195 27340 7235
rect 27380 7195 27381 7235
rect 12256 7184 12298 7193
rect 16107 7186 16149 7195
rect 24555 7186 24597 7195
rect 27339 7186 27381 7195
rect 27819 7235 27861 7244
rect 27819 7195 27820 7235
rect 27860 7195 27861 7235
rect 27819 7186 27861 7195
rect 29355 7235 29397 7244
rect 29355 7195 29356 7235
rect 29396 7195 29397 7235
rect 30603 7204 30604 7244
rect 30644 7204 30645 7244
rect 30603 7195 30645 7204
rect 32715 7244 32757 7253
rect 32715 7204 32716 7244
rect 32756 7204 32757 7244
rect 32715 7195 32757 7204
rect 33003 7244 33045 7253
rect 33003 7204 33004 7244
rect 33044 7204 33045 7244
rect 33003 7195 33045 7204
rect 33579 7244 33621 7253
rect 33579 7204 33580 7244
rect 33620 7204 33621 7244
rect 33579 7195 33621 7204
rect 37899 7244 37941 7253
rect 37899 7204 37900 7244
rect 37940 7204 37941 7244
rect 37899 7195 37941 7204
rect 29355 7186 29397 7195
rect 1227 7160 1269 7169
rect 1227 7120 1228 7160
rect 1268 7120 1269 7160
rect 1227 7111 1269 7120
rect 1611 7160 1653 7169
rect 1611 7120 1612 7160
rect 1652 7120 1653 7160
rect 1611 7111 1653 7120
rect 1851 7160 1893 7169
rect 1851 7120 1852 7160
rect 1892 7120 1893 7160
rect 1851 7111 1893 7120
rect 9675 7160 9717 7169
rect 9675 7120 9676 7160
rect 9716 7120 9717 7160
rect 9675 7111 9717 7120
rect 11115 7160 11157 7169
rect 11115 7120 11116 7160
rect 11156 7120 11157 7160
rect 11115 7111 11157 7120
rect 11355 7160 11397 7169
rect 11355 7120 11356 7160
rect 11396 7120 11397 7160
rect 11355 7111 11397 7120
rect 12891 7160 12933 7169
rect 12891 7120 12892 7160
rect 12932 7120 12933 7160
rect 12891 7111 12933 7120
rect 21675 7160 21717 7169
rect 21675 7120 21676 7160
rect 21716 7120 21717 7160
rect 21675 7111 21717 7120
rect 26859 7160 26901 7169
rect 26859 7120 26860 7160
rect 26900 7120 26901 7160
rect 26859 7111 26901 7120
rect 28395 7160 28437 7169
rect 28395 7120 28396 7160
rect 28436 7120 28437 7160
rect 28395 7111 28437 7120
rect 32331 7160 32373 7169
rect 32331 7120 32332 7160
rect 32372 7120 32373 7160
rect 32331 7111 32373 7120
rect 34155 7160 34197 7169
rect 34155 7120 34156 7160
rect 34196 7120 34197 7160
rect 34155 7111 34197 7120
rect 34731 7160 34773 7169
rect 34731 7120 34732 7160
rect 34772 7120 34773 7160
rect 34731 7111 34773 7120
rect 35307 7160 35349 7169
rect 35307 7120 35308 7160
rect 35348 7120 35349 7160
rect 35307 7111 35349 7120
rect 35883 7160 35925 7169
rect 35883 7120 35884 7160
rect 35924 7120 35925 7160
rect 35883 7111 35925 7120
rect 36459 7160 36501 7169
rect 36459 7120 36460 7160
rect 36500 7120 36501 7160
rect 36459 7111 36501 7120
rect 37035 7160 37077 7169
rect 37035 7120 37036 7160
rect 37076 7120 37077 7160
rect 37035 7111 37077 7120
rect 37323 7160 37365 7169
rect 37323 7120 37324 7160
rect 37364 7120 37365 7160
rect 37323 7111 37365 7120
rect 41931 7160 41973 7169
rect 41931 7120 41932 7160
rect 41972 7120 41973 7160
rect 41931 7111 41973 7120
rect 42315 7160 42357 7169
rect 42315 7120 42316 7160
rect 42356 7120 42357 7160
rect 42315 7111 42357 7120
rect 42699 7160 42741 7169
rect 42699 7120 42700 7160
rect 42740 7120 42741 7160
rect 42699 7111 42741 7120
rect 43083 7160 43125 7169
rect 43083 7120 43084 7160
rect 43124 7120 43125 7160
rect 43083 7111 43125 7120
rect 43467 7160 43509 7169
rect 43467 7120 43468 7160
rect 43508 7120 43509 7160
rect 43467 7111 43509 7120
rect 43755 7160 43797 7169
rect 43755 7120 43756 7160
rect 43796 7120 43797 7160
rect 43755 7111 43797 7120
rect 44043 7160 44085 7169
rect 44043 7120 44044 7160
rect 44084 7120 44085 7160
rect 44043 7111 44085 7120
rect 44235 7160 44277 7169
rect 44235 7120 44236 7160
rect 44276 7120 44277 7160
rect 44235 7111 44277 7120
rect 44715 7160 44757 7169
rect 44715 7120 44716 7160
rect 44756 7120 44757 7160
rect 44715 7111 44757 7120
rect 44907 7160 44949 7169
rect 44907 7120 44908 7160
rect 44948 7120 44949 7160
rect 44907 7111 44949 7120
rect 1467 7076 1509 7085
rect 1467 7036 1468 7076
rect 1508 7036 1509 7076
rect 1467 7027 1509 7036
rect 9915 7076 9957 7085
rect 9915 7036 9916 7076
rect 9956 7036 9957 7076
rect 9915 7027 9957 7036
rect 10827 7076 10869 7085
rect 10827 7036 10828 7076
rect 10868 7036 10869 7076
rect 10827 7027 10869 7036
rect 28155 7076 28197 7085
rect 28155 7036 28156 7076
rect 28196 7036 28197 7076
rect 28155 7027 28197 7036
rect 42843 7076 42885 7085
rect 42843 7036 42844 7076
rect 42884 7036 42885 7076
rect 42843 7027 42885 7036
rect 16299 6992 16341 7001
rect 16299 6952 16300 6992
rect 16340 6952 16341 6992
rect 16299 6943 16341 6952
rect 21915 6992 21957 7001
rect 21915 6952 21916 6992
rect 21956 6952 21957 6992
rect 21915 6943 21957 6952
rect 24747 6992 24789 7001
rect 24747 6952 24748 6992
rect 24788 6952 24789 6992
rect 24747 6943 24789 6952
rect 32571 6992 32613 7001
rect 32571 6952 32572 6992
rect 32612 6952 32613 6992
rect 32571 6943 32613 6952
rect 41691 6992 41733 7001
rect 41691 6952 41692 6992
rect 41732 6952 41733 6992
rect 41691 6943 41733 6952
rect 42075 6992 42117 7001
rect 42075 6952 42076 6992
rect 42116 6952 42117 6992
rect 42075 6943 42117 6952
rect 42459 6992 42501 7001
rect 42459 6952 42460 6992
rect 42500 6952 42501 6992
rect 42459 6943 42501 6952
rect 43227 6992 43269 7001
rect 43227 6952 43228 6992
rect 43268 6952 43269 6992
rect 43227 6943 43269 6952
rect 44475 6992 44517 7001
rect 44475 6952 44476 6992
rect 44516 6952 44517 6992
rect 44475 6943 44517 6952
rect 45147 6992 45189 7001
rect 45147 6952 45148 6992
rect 45188 6952 45189 6992
rect 45147 6943 45189 6952
rect 1152 6824 45216 6848
rect 1152 6784 3688 6824
rect 3728 6784 3770 6824
rect 3810 6784 3852 6824
rect 3892 6784 3934 6824
rect 3974 6784 4016 6824
rect 4056 6784 18808 6824
rect 18848 6784 18890 6824
rect 18930 6784 18972 6824
rect 19012 6784 19054 6824
rect 19094 6784 19136 6824
rect 19176 6784 33928 6824
rect 33968 6784 34010 6824
rect 34050 6784 34092 6824
rect 34132 6784 34174 6824
rect 34214 6784 34256 6824
rect 34296 6784 45216 6824
rect 1152 6760 45216 6784
rect 7947 6656 7989 6665
rect 7947 6616 7948 6656
rect 7988 6616 7989 6656
rect 7947 6607 7989 6616
rect 11242 6656 11300 6657
rect 11242 6616 11251 6656
rect 11291 6616 11300 6656
rect 11242 6615 11300 6616
rect 1467 6572 1509 6581
rect 1467 6532 1468 6572
rect 1508 6532 1509 6572
rect 1467 6523 1509 6532
rect 12171 6572 12213 6581
rect 12171 6532 12172 6572
rect 12212 6532 12213 6572
rect 12171 6523 12213 6532
rect 1227 6488 1269 6497
rect 1227 6448 1228 6488
rect 1268 6448 1269 6488
rect 1227 6439 1269 6448
rect 1611 6488 1653 6497
rect 1611 6448 1612 6488
rect 1652 6448 1653 6488
rect 1611 6439 1653 6448
rect 6123 6488 6165 6497
rect 6123 6448 6124 6488
rect 6164 6448 6165 6488
rect 6123 6439 6165 6448
rect 9003 6488 9045 6497
rect 9003 6448 9004 6488
rect 9044 6448 9045 6488
rect 9003 6439 9045 6448
rect 9963 6488 10005 6497
rect 9963 6448 9964 6488
rect 10004 6448 10005 6488
rect 9963 6439 10005 6448
rect 17163 6488 17205 6497
rect 17163 6448 17164 6488
rect 17204 6448 17205 6488
rect 17163 6439 17205 6448
rect 44523 6488 44565 6497
rect 44523 6448 44524 6488
rect 44564 6448 44565 6488
rect 44523 6439 44565 6448
rect 6507 6404 6549 6413
rect 6507 6364 6508 6404
rect 6548 6364 6549 6404
rect 6507 6355 6549 6364
rect 7755 6404 7813 6405
rect 7755 6364 7764 6404
rect 7804 6364 7813 6404
rect 7755 6363 7813 6364
rect 9466 6404 9524 6405
rect 9466 6364 9475 6404
rect 9515 6364 9524 6404
rect 9466 6363 9524 6364
rect 9579 6404 9621 6413
rect 9579 6364 9580 6404
rect 9620 6364 9621 6404
rect 9579 6355 9621 6364
rect 10059 6404 10101 6413
rect 10059 6364 10060 6404
rect 10100 6364 10101 6404
rect 10059 6355 10101 6364
rect 10531 6404 10589 6405
rect 10531 6364 10540 6404
rect 10580 6364 10589 6404
rect 10531 6363 10589 6364
rect 11050 6404 11108 6405
rect 11050 6364 11059 6404
rect 11099 6364 11108 6404
rect 11050 6363 11108 6364
rect 11499 6404 11541 6413
rect 11499 6364 11500 6404
rect 11540 6364 11541 6404
rect 11499 6355 11541 6364
rect 11770 6404 11828 6405
rect 11770 6364 11779 6404
rect 11819 6364 11828 6404
rect 11770 6363 11828 6364
rect 11883 6320 11925 6329
rect 11883 6280 11884 6320
rect 11924 6280 11925 6320
rect 11883 6271 11925 6280
rect 44907 6320 44949 6329
rect 44907 6280 44908 6320
rect 44948 6280 44949 6320
rect 44907 6271 44949 6280
rect 1851 6236 1893 6245
rect 1851 6196 1852 6236
rect 1892 6196 1893 6236
rect 1851 6187 1893 6196
rect 6363 6236 6405 6245
rect 6363 6196 6364 6236
rect 6404 6196 6405 6236
rect 6363 6187 6405 6196
rect 9243 6236 9285 6245
rect 9243 6196 9244 6236
rect 9284 6196 9285 6236
rect 9243 6187 9285 6196
rect 16923 6236 16965 6245
rect 16923 6196 16924 6236
rect 16964 6196 16965 6236
rect 16923 6187 16965 6196
rect 43642 6236 43700 6237
rect 43642 6196 43651 6236
rect 43691 6196 43700 6236
rect 43642 6195 43700 6196
rect 43930 6236 43988 6237
rect 43930 6196 43939 6236
rect 43979 6196 43988 6236
rect 43930 6195 43988 6196
rect 44218 6236 44276 6237
rect 44218 6196 44227 6236
rect 44267 6196 44276 6236
rect 44218 6195 44276 6196
rect 44763 6236 44805 6245
rect 44763 6196 44764 6236
rect 44804 6196 44805 6236
rect 44763 6187 44805 6196
rect 1152 6068 45216 6092
rect 1152 6028 4928 6068
rect 4968 6028 5010 6068
rect 5050 6028 5092 6068
rect 5132 6028 5174 6068
rect 5214 6028 5256 6068
rect 5296 6028 20048 6068
rect 20088 6028 20130 6068
rect 20170 6028 20212 6068
rect 20252 6028 20294 6068
rect 20334 6028 20376 6068
rect 20416 6028 35168 6068
rect 35208 6028 35250 6068
rect 35290 6028 35332 6068
rect 35372 6028 35414 6068
rect 35454 6028 35496 6068
rect 35536 6028 45216 6068
rect 1152 6004 45216 6028
rect 11115 5900 11157 5909
rect 11115 5860 11116 5900
rect 11156 5860 11157 5900
rect 11115 5851 11157 5860
rect 13179 5900 13221 5909
rect 13179 5860 13180 5900
rect 13220 5860 13221 5900
rect 13179 5851 13221 5860
rect 43738 5900 43796 5901
rect 43738 5860 43747 5900
rect 43787 5860 43796 5900
rect 43738 5859 43796 5860
rect 44218 5900 44276 5901
rect 44218 5860 44227 5900
rect 44267 5860 44276 5900
rect 44218 5859 44276 5860
rect 9370 5732 9428 5733
rect 9370 5692 9379 5732
rect 9419 5692 9428 5732
rect 9370 5691 9428 5692
rect 9483 5732 9525 5741
rect 9483 5692 9484 5732
rect 9524 5692 9525 5732
rect 9483 5683 9525 5692
rect 9867 5732 9909 5741
rect 13323 5732 13365 5741
rect 9867 5692 9868 5732
rect 9908 5692 9909 5732
rect 9867 5683 9909 5692
rect 10443 5723 10485 5732
rect 10443 5683 10444 5723
rect 10484 5683 10485 5723
rect 10443 5674 10485 5683
rect 10923 5723 10965 5732
rect 10923 5683 10924 5723
rect 10964 5683 10965 5723
rect 13323 5692 13324 5732
rect 13364 5692 13365 5732
rect 13323 5683 13365 5692
rect 10923 5674 10965 5683
rect 1227 5648 1269 5657
rect 1227 5608 1228 5648
rect 1268 5608 1269 5648
rect 1227 5599 1269 5608
rect 1611 5648 1653 5657
rect 1611 5608 1612 5648
rect 1652 5608 1653 5648
rect 1611 5599 1653 5608
rect 1995 5648 2037 5657
rect 1995 5608 1996 5648
rect 2036 5608 2037 5648
rect 1995 5599 2037 5608
rect 9963 5648 10005 5657
rect 9963 5608 9964 5648
rect 10004 5608 10005 5648
rect 9963 5599 10005 5608
rect 11307 5648 11349 5657
rect 11307 5608 11308 5648
rect 11348 5608 11349 5648
rect 11307 5599 11349 5608
rect 11547 5648 11589 5657
rect 11547 5608 11548 5648
rect 11588 5608 11589 5648
rect 11547 5599 11589 5608
rect 43659 5648 43701 5657
rect 43659 5608 43660 5648
rect 43700 5608 43701 5648
rect 43659 5599 43701 5608
rect 44043 5648 44085 5657
rect 44043 5608 44044 5648
rect 44084 5608 44085 5648
rect 44043 5599 44085 5608
rect 44523 5648 44565 5657
rect 44523 5608 44524 5648
rect 44564 5608 44565 5648
rect 44523 5599 44565 5608
rect 44907 5648 44949 5657
rect 44907 5608 44908 5648
rect 44948 5608 44949 5648
rect 44907 5599 44949 5608
rect 45147 5648 45189 5657
rect 45147 5608 45148 5648
rect 45188 5608 45189 5648
rect 45147 5599 45189 5608
rect 1467 5480 1509 5489
rect 1467 5440 1468 5480
rect 1508 5440 1509 5480
rect 1467 5431 1509 5440
rect 1851 5480 1893 5489
rect 1851 5440 1852 5480
rect 1892 5440 1893 5480
rect 1851 5431 1893 5440
rect 2235 5480 2277 5489
rect 2235 5440 2236 5480
rect 2276 5440 2277 5480
rect 2235 5431 2277 5440
rect 44763 5480 44805 5489
rect 44763 5440 44764 5480
rect 44804 5440 44805 5480
rect 44763 5431 44805 5440
rect 1152 5312 45216 5336
rect 1152 5272 3688 5312
rect 3728 5272 3770 5312
rect 3810 5272 3852 5312
rect 3892 5272 3934 5312
rect 3974 5272 4016 5312
rect 4056 5272 18808 5312
rect 18848 5272 18890 5312
rect 18930 5272 18972 5312
rect 19012 5272 19054 5312
rect 19094 5272 19136 5312
rect 19176 5272 33928 5312
rect 33968 5272 34010 5312
rect 34050 5272 34092 5312
rect 34132 5272 34174 5312
rect 34214 5272 34256 5312
rect 34296 5272 45216 5312
rect 1152 5248 45216 5272
rect 32955 5144 32997 5153
rect 32955 5104 32956 5144
rect 32996 5104 32997 5144
rect 32955 5095 32997 5104
rect 42843 5144 42885 5153
rect 42843 5104 42844 5144
rect 42884 5104 42885 5144
rect 42843 5095 42885 5104
rect 45147 5144 45189 5153
rect 45147 5104 45148 5144
rect 45188 5104 45189 5144
rect 45147 5095 45189 5104
rect 30987 4976 31029 4985
rect 30987 4936 30988 4976
rect 31028 4936 31029 4976
rect 30987 4927 31029 4936
rect 33195 4976 33237 4985
rect 33195 4936 33196 4976
rect 33236 4936 33237 4976
rect 33195 4927 33237 4936
rect 43083 4976 43125 4985
rect 43083 4936 43084 4976
rect 43124 4936 43125 4976
rect 43083 4927 43125 4936
rect 44523 4976 44565 4985
rect 44523 4936 44524 4976
rect 44564 4936 44565 4976
rect 44523 4927 44565 4936
rect 44907 4976 44949 4985
rect 44907 4936 44908 4976
rect 44948 4936 44949 4976
rect 44907 4927 44949 4936
rect 31371 4892 31413 4901
rect 31371 4852 31372 4892
rect 31412 4852 31413 4892
rect 31371 4843 31413 4852
rect 32611 4892 32669 4893
rect 32611 4852 32620 4892
rect 32660 4852 32669 4892
rect 32611 4851 32669 4852
rect 44235 4892 44277 4901
rect 44235 4852 44236 4892
rect 44276 4852 44277 4892
rect 44235 4843 44277 4852
rect 31227 4724 31269 4733
rect 31227 4684 31228 4724
rect 31268 4684 31269 4724
rect 31227 4675 31269 4684
rect 32811 4724 32853 4733
rect 32811 4684 32812 4724
rect 32852 4684 32853 4724
rect 32811 4675 32853 4684
rect 43450 4724 43508 4725
rect 43450 4684 43459 4724
rect 43499 4684 43508 4724
rect 43450 4683 43508 4684
rect 43642 4724 43700 4725
rect 43642 4684 43651 4724
rect 43691 4684 43700 4724
rect 43642 4683 43700 4684
rect 43930 4724 43988 4725
rect 43930 4684 43939 4724
rect 43979 4684 43988 4724
rect 43930 4683 43988 4684
rect 44763 4724 44805 4733
rect 44763 4684 44764 4724
rect 44804 4684 44805 4724
rect 44763 4675 44805 4684
rect 1152 4556 45216 4580
rect 1152 4516 4928 4556
rect 4968 4516 5010 4556
rect 5050 4516 5092 4556
rect 5132 4516 5174 4556
rect 5214 4516 5256 4556
rect 5296 4516 20048 4556
rect 20088 4516 20130 4556
rect 20170 4516 20212 4556
rect 20252 4516 20294 4556
rect 20334 4516 20376 4556
rect 20416 4516 35168 4556
rect 35208 4516 35250 4556
rect 35290 4516 35332 4556
rect 35372 4516 35414 4556
rect 35454 4516 35496 4556
rect 35536 4516 45216 4556
rect 1152 4492 45216 4516
rect 19995 4388 20037 4397
rect 19995 4348 19996 4388
rect 20036 4348 20037 4388
rect 19995 4339 20037 4348
rect 33483 4388 33525 4397
rect 33483 4348 33484 4388
rect 33524 4348 33525 4388
rect 33483 4339 33525 4348
rect 43930 4388 43988 4389
rect 43930 4348 43939 4388
rect 43979 4348 43988 4388
rect 43930 4347 43988 4348
rect 44602 4388 44660 4389
rect 44602 4348 44611 4388
rect 44651 4348 44660 4388
rect 44602 4347 44660 4348
rect 24027 4304 24069 4313
rect 24027 4264 24028 4304
rect 24068 4264 24069 4304
rect 24027 4255 24069 4264
rect 25611 4304 25653 4313
rect 25611 4264 25612 4304
rect 25652 4264 25653 4304
rect 25611 4255 25653 4264
rect 27099 4304 27141 4313
rect 27099 4264 27100 4304
rect 27140 4264 27141 4304
rect 27099 4255 27141 4264
rect 31467 4304 31509 4313
rect 31467 4264 31468 4304
rect 31508 4264 31509 4304
rect 31467 4255 31509 4264
rect 33963 4304 34005 4313
rect 33963 4264 33964 4304
rect 34004 4264 34005 4304
rect 33963 4255 34005 4264
rect 41979 4304 42021 4313
rect 41979 4264 41980 4304
rect 42020 4264 42021 4304
rect 41979 4255 42021 4264
rect 42747 4304 42789 4313
rect 42747 4264 42748 4304
rect 42788 4264 42789 4304
rect 42747 4255 42789 4264
rect 45147 4304 45189 4313
rect 45147 4264 45148 4304
rect 45188 4264 45189 4304
rect 45147 4255 45189 4264
rect 9675 4220 9717 4229
rect 9675 4180 9676 4220
rect 9716 4180 9717 4220
rect 9675 4171 9717 4180
rect 9776 4220 9834 4221
rect 9776 4180 9785 4220
rect 9825 4180 9834 4220
rect 9776 4179 9834 4180
rect 10059 4220 10101 4229
rect 10059 4180 10060 4220
rect 10100 4180 10101 4220
rect 10059 4171 10101 4180
rect 18027 4220 18069 4229
rect 22923 4220 22965 4229
rect 18027 4180 18028 4220
rect 18068 4180 18069 4220
rect 18027 4171 18069 4180
rect 19275 4211 19317 4220
rect 19275 4171 19276 4211
rect 19316 4171 19317 4211
rect 19275 4162 19317 4171
rect 21675 4211 21717 4220
rect 21675 4171 21676 4211
rect 21716 4171 21717 4211
rect 22923 4180 22924 4220
rect 22964 4180 22965 4220
rect 22923 4171 22965 4180
rect 24171 4220 24213 4229
rect 25899 4220 25941 4229
rect 24171 4180 24172 4220
rect 24212 4180 24213 4220
rect 24171 4171 24213 4180
rect 25419 4211 25461 4220
rect 25419 4171 25420 4211
rect 25460 4171 25461 4211
rect 25899 4180 25900 4220
rect 25940 4180 25941 4220
rect 25899 4171 25941 4180
rect 26146 4220 26204 4221
rect 26146 4180 26155 4220
rect 26195 4180 26204 4220
rect 26146 4179 26204 4180
rect 26268 4220 26326 4221
rect 26268 4180 26277 4220
rect 26317 4180 26326 4220
rect 26268 4179 26326 4180
rect 30027 4220 30069 4229
rect 31738 4220 31796 4221
rect 30027 4180 30028 4220
rect 30068 4180 30069 4220
rect 30027 4171 30069 4180
rect 31275 4211 31317 4220
rect 31275 4171 31276 4211
rect 31316 4171 31317 4211
rect 31738 4180 31747 4220
rect 31787 4180 31796 4220
rect 31738 4179 31796 4180
rect 31851 4220 31893 4229
rect 31851 4180 31852 4220
rect 31892 4180 31893 4220
rect 31851 4171 31893 4180
rect 32235 4220 32277 4229
rect 34064 4220 34122 4221
rect 32235 4180 32236 4220
rect 32276 4180 32277 4220
rect 32235 4171 32277 4180
rect 32811 4211 32853 4220
rect 32811 4171 32812 4211
rect 32852 4171 32853 4211
rect 21675 4162 21717 4171
rect 25419 4162 25461 4171
rect 31275 4162 31317 4171
rect 32811 4162 32853 4171
rect 33291 4211 33333 4220
rect 33291 4171 33292 4211
rect 33332 4171 33333 4211
rect 34064 4180 34073 4220
rect 34113 4180 34122 4220
rect 34064 4179 34122 4180
rect 34347 4220 34389 4229
rect 34347 4180 34348 4220
rect 34388 4180 34389 4220
rect 34347 4171 34389 4180
rect 33291 4162 33333 4171
rect 17643 4136 17685 4145
rect 17643 4096 17644 4136
rect 17684 4096 17685 4136
rect 17643 4087 17685 4096
rect 17883 4136 17925 4145
rect 17883 4096 17884 4136
rect 17924 4096 17925 4136
rect 17883 4087 17925 4096
rect 19707 4136 19749 4145
rect 19707 4096 19708 4136
rect 19748 4096 19749 4136
rect 19707 4087 19749 4096
rect 20331 4136 20373 4145
rect 20331 4096 20332 4136
rect 20372 4096 20373 4136
rect 20331 4087 20373 4096
rect 21099 4136 21141 4145
rect 21099 4096 21100 4136
rect 21140 4096 21141 4136
rect 21099 4087 21141 4096
rect 21339 4136 21381 4145
rect 21339 4096 21340 4136
rect 21380 4096 21381 4136
rect 21339 4087 21381 4096
rect 23787 4136 23829 4145
rect 23787 4096 23788 4136
rect 23828 4096 23829 4136
rect 23787 4087 23829 4096
rect 26763 4136 26805 4145
rect 26763 4096 26764 4136
rect 26804 4096 26805 4136
rect 26763 4087 26805 4096
rect 27339 4136 27381 4145
rect 27339 4096 27340 4136
rect 27380 4096 27381 4136
rect 27339 4087 27381 4096
rect 32331 4136 32373 4145
rect 32331 4096 32332 4136
rect 32372 4096 32373 4136
rect 32331 4087 32373 4096
rect 38379 4136 38421 4145
rect 38379 4096 38380 4136
rect 38420 4096 38421 4136
rect 38379 4087 38421 4096
rect 38571 4136 38613 4145
rect 38571 4096 38572 4136
rect 38612 4096 38613 4136
rect 38571 4087 38613 4096
rect 42219 4136 42261 4145
rect 42219 4096 42220 4136
rect 42260 4096 42261 4136
rect 42219 4087 42261 4096
rect 42603 4136 42645 4145
rect 42603 4096 42604 4136
rect 42644 4096 42645 4136
rect 42603 4087 42645 4096
rect 42987 4136 43029 4145
rect 42987 4096 42988 4136
rect 43028 4096 43029 4136
rect 42987 4087 43029 4096
rect 43371 4136 43413 4145
rect 43371 4096 43372 4136
rect 43412 4096 43413 4136
rect 43371 4087 43413 4096
rect 43755 4136 43797 4145
rect 43755 4096 43756 4136
rect 43796 4096 43797 4136
rect 43755 4087 43797 4096
rect 44235 4136 44277 4145
rect 44235 4096 44236 4136
rect 44276 4096 44277 4136
rect 44235 4087 44277 4096
rect 44619 4136 44661 4145
rect 44619 4096 44620 4136
rect 44660 4096 44661 4136
rect 44619 4087 44661 4096
rect 44907 4136 44949 4145
rect 44907 4096 44908 4136
rect 44948 4096 44949 4136
rect 44907 4087 44949 4096
rect 26571 4052 26613 4061
rect 26571 4012 26572 4052
rect 26612 4012 26613 4052
rect 26571 4003 26613 4012
rect 44475 4052 44517 4061
rect 44475 4012 44476 4052
rect 44516 4012 44517 4052
rect 44475 4003 44517 4012
rect 9387 3968 9429 3977
rect 9387 3928 9388 3968
rect 9428 3928 9429 3968
rect 9387 3919 9429 3928
rect 19467 3968 19509 3977
rect 19467 3928 19468 3968
rect 19508 3928 19509 3968
rect 19467 3919 19509 3928
rect 20091 3968 20133 3977
rect 20091 3928 20092 3968
rect 20132 3928 20133 3968
rect 20091 3919 20133 3928
rect 21483 3968 21525 3977
rect 21483 3928 21484 3968
rect 21524 3928 21525 3968
rect 21483 3919 21525 3928
rect 27003 3968 27045 3977
rect 27003 3928 27004 3968
rect 27044 3928 27045 3968
rect 27003 3919 27045 3928
rect 33675 3968 33717 3977
rect 33675 3928 33676 3968
rect 33716 3928 33717 3968
rect 33675 3919 33717 3928
rect 38811 3968 38853 3977
rect 38811 3928 38812 3968
rect 38852 3928 38853 3968
rect 38811 3919 38853 3928
rect 42363 3968 42405 3977
rect 42363 3928 42364 3968
rect 42404 3928 42405 3968
rect 42363 3919 42405 3928
rect 43131 3968 43173 3977
rect 43131 3928 43132 3968
rect 43172 3928 43173 3968
rect 43131 3919 43173 3928
rect 43515 3968 43557 3977
rect 43515 3928 43516 3968
rect 43556 3928 43557 3968
rect 43515 3919 43557 3928
rect 1152 3800 45216 3824
rect 1152 3760 3688 3800
rect 3728 3760 3770 3800
rect 3810 3760 3852 3800
rect 3892 3760 3934 3800
rect 3974 3760 4016 3800
rect 4056 3760 18808 3800
rect 18848 3760 18890 3800
rect 18930 3760 18972 3800
rect 19012 3760 19054 3800
rect 19094 3760 19136 3800
rect 19176 3760 33928 3800
rect 33968 3760 34010 3800
rect 34050 3760 34092 3800
rect 34132 3760 34174 3800
rect 34214 3760 34256 3800
rect 34296 3760 45216 3800
rect 1152 3736 45216 3760
rect 9243 3632 9285 3641
rect 9243 3592 9244 3632
rect 9284 3592 9285 3632
rect 9243 3583 9285 3592
rect 9627 3632 9669 3641
rect 9627 3592 9628 3632
rect 9668 3592 9669 3632
rect 9627 3583 9669 3592
rect 11211 3632 11253 3641
rect 11211 3592 11212 3632
rect 11252 3592 11253 3632
rect 11211 3583 11253 3592
rect 12027 3632 12069 3641
rect 12027 3592 12028 3632
rect 12068 3592 12069 3632
rect 12027 3583 12069 3592
rect 13611 3632 13653 3641
rect 13611 3592 13612 3632
rect 13652 3592 13653 3632
rect 13611 3583 13653 3592
rect 18171 3632 18213 3641
rect 18171 3592 18172 3632
rect 18212 3592 18213 3632
rect 18171 3583 18213 3592
rect 32571 3632 32613 3641
rect 32571 3592 32572 3632
rect 32612 3592 32613 3632
rect 32571 3583 32613 3592
rect 42747 3632 42789 3641
rect 42747 3592 42748 3632
rect 42788 3592 42789 3632
rect 42747 3583 42789 3592
rect 43899 3632 43941 3641
rect 43899 3592 43900 3632
rect 43940 3592 43941 3632
rect 43899 3583 43941 3592
rect 45147 3632 45189 3641
rect 45147 3592 45148 3632
rect 45188 3592 45189 3632
rect 45147 3583 45189 3592
rect 17787 3548 17829 3557
rect 17787 3508 17788 3548
rect 17828 3508 17829 3548
rect 17787 3499 17829 3508
rect 21099 3548 21141 3557
rect 21099 3508 21100 3548
rect 21140 3508 21141 3548
rect 21099 3499 21141 3508
rect 26859 3548 26901 3557
rect 26859 3508 26860 3548
rect 26900 3508 26901 3548
rect 26859 3499 26901 3508
rect 27867 3548 27909 3557
rect 27867 3508 27868 3548
rect 27908 3508 27909 3548
rect 27867 3499 27909 3508
rect 29451 3548 29493 3557
rect 29451 3508 29452 3548
rect 29492 3508 29493 3548
rect 29451 3499 29493 3508
rect 32955 3548 32997 3557
rect 32955 3508 32956 3548
rect 32996 3508 32997 3548
rect 32955 3499 32997 3508
rect 42267 3548 42309 3557
rect 42267 3508 42268 3548
rect 42308 3508 42309 3548
rect 42267 3499 42309 3508
rect 43131 3548 43173 3557
rect 43131 3508 43132 3548
rect 43172 3508 43173 3548
rect 43131 3499 43173 3508
rect 9003 3464 9045 3473
rect 9003 3424 9004 3464
rect 9044 3424 9045 3464
rect 9003 3415 9045 3424
rect 9387 3464 9429 3473
rect 9387 3424 9388 3464
rect 9428 3424 9429 3464
rect 9387 3415 9429 3424
rect 11787 3464 11829 3473
rect 11787 3424 11788 3464
rect 11828 3424 11829 3464
rect 11787 3415 11829 3424
rect 15435 3464 15477 3473
rect 15435 3424 15436 3464
rect 15476 3424 15477 3464
rect 15435 3415 15477 3424
rect 15771 3464 15813 3473
rect 15771 3424 15772 3464
rect 15812 3424 15813 3464
rect 15771 3415 15813 3424
rect 16011 3464 16053 3473
rect 16011 3424 16012 3464
rect 16052 3424 16053 3464
rect 16011 3415 16053 3424
rect 18027 3464 18069 3473
rect 18027 3424 18028 3464
rect 18068 3424 18069 3464
rect 18027 3415 18069 3424
rect 18411 3464 18453 3473
rect 18411 3424 18412 3464
rect 18452 3424 18453 3464
rect 18411 3415 18453 3424
rect 18795 3464 18837 3473
rect 18795 3424 18796 3464
rect 18836 3424 18837 3464
rect 18795 3415 18837 3424
rect 19563 3464 19605 3473
rect 19563 3424 19564 3464
rect 19604 3424 19605 3464
rect 19563 3415 19605 3424
rect 27003 3464 27045 3473
rect 27003 3424 27004 3464
rect 27044 3424 27045 3464
rect 27003 3415 27045 3424
rect 27243 3464 27285 3473
rect 27243 3424 27244 3464
rect 27284 3424 27285 3464
rect 27243 3415 27285 3424
rect 27627 3464 27669 3473
rect 27627 3424 27628 3464
rect 27668 3424 27669 3464
rect 27627 3415 27669 3424
rect 30219 3464 30261 3473
rect 30219 3424 30220 3464
rect 30260 3424 30261 3464
rect 30219 3415 30261 3424
rect 31179 3464 31221 3473
rect 31179 3424 31180 3464
rect 31220 3424 31221 3464
rect 31179 3415 31221 3424
rect 32811 3464 32853 3473
rect 32811 3424 32812 3464
rect 32852 3424 32853 3464
rect 32811 3415 32853 3424
rect 33195 3464 33237 3473
rect 33195 3424 33196 3464
rect 33236 3424 33237 3464
rect 33195 3415 33237 3424
rect 33579 3464 33621 3473
rect 33579 3424 33580 3464
rect 33620 3424 33621 3464
rect 33579 3415 33621 3424
rect 37515 3464 37557 3473
rect 37515 3424 37516 3464
rect 37556 3424 37557 3464
rect 37515 3415 37557 3424
rect 37803 3464 37845 3473
rect 37803 3424 37804 3464
rect 37844 3424 37845 3464
rect 37803 3415 37845 3424
rect 38187 3464 38229 3473
rect 38187 3424 38188 3464
rect 38228 3424 38229 3464
rect 38187 3415 38229 3424
rect 38571 3464 38613 3473
rect 38571 3424 38572 3464
rect 38612 3424 38613 3464
rect 38571 3415 38613 3424
rect 39051 3464 39093 3473
rect 39051 3424 39052 3464
rect 39092 3424 39093 3464
rect 39051 3415 39093 3424
rect 39339 3464 39381 3473
rect 39339 3424 39340 3464
rect 39380 3424 39381 3464
rect 39339 3415 39381 3424
rect 39723 3464 39765 3473
rect 39723 3424 39724 3464
rect 39764 3424 39765 3464
rect 39723 3415 39765 3424
rect 42507 3464 42549 3473
rect 42507 3424 42508 3464
rect 42548 3424 42549 3464
rect 42507 3415 42549 3424
rect 42987 3464 43029 3473
rect 42987 3424 42988 3464
rect 43028 3424 43029 3464
rect 42987 3415 43029 3424
rect 43371 3464 43413 3473
rect 43371 3424 43372 3464
rect 43412 3424 43413 3464
rect 43371 3415 43413 3424
rect 43755 3464 43797 3473
rect 43755 3424 43756 3464
rect 43796 3424 43797 3464
rect 43755 3415 43797 3424
rect 44139 3464 44181 3473
rect 44139 3424 44140 3464
rect 44180 3424 44181 3464
rect 44139 3415 44181 3424
rect 44523 3464 44565 3473
rect 44523 3424 44524 3464
rect 44564 3424 44565 3464
rect 44523 3415 44565 3424
rect 44907 3464 44949 3473
rect 44907 3424 44908 3464
rect 44948 3424 44949 3464
rect 44907 3415 44949 3424
rect 9771 3380 9813 3389
rect 9771 3340 9772 3380
rect 9812 3340 9813 3380
rect 9771 3331 9813 3340
rect 11011 3380 11069 3381
rect 11011 3340 11020 3380
rect 11060 3340 11069 3380
rect 11011 3339 11069 3340
rect 12171 3380 12213 3389
rect 12171 3340 12172 3380
rect 12212 3340 12213 3380
rect 12171 3331 12213 3340
rect 13411 3380 13469 3381
rect 13411 3340 13420 3380
rect 13460 3340 13469 3380
rect 13411 3339 13469 3340
rect 13803 3380 13845 3389
rect 13803 3340 13804 3380
rect 13844 3340 13845 3380
rect 13803 3331 13845 3340
rect 15043 3380 15101 3381
rect 15043 3340 15052 3380
rect 15092 3340 15101 3380
rect 15043 3339 15101 3340
rect 16203 3380 16245 3389
rect 16203 3340 16204 3380
rect 16244 3340 16245 3380
rect 16203 3331 16245 3340
rect 17443 3380 17501 3381
rect 17443 3340 17452 3380
rect 17492 3340 17501 3380
rect 17443 3339 17501 3340
rect 19066 3380 19124 3381
rect 19066 3340 19075 3380
rect 19115 3340 19124 3380
rect 19066 3339 19124 3340
rect 19168 3380 19226 3381
rect 19168 3340 19177 3380
rect 19217 3340 19226 3380
rect 19168 3339 19226 3340
rect 19659 3380 19701 3389
rect 19659 3340 19660 3380
rect 19700 3340 19701 3380
rect 19659 3331 19701 3340
rect 20131 3380 20189 3381
rect 20131 3340 20140 3380
rect 20180 3340 20189 3380
rect 20131 3339 20189 3340
rect 20619 3380 20677 3381
rect 21771 3380 21813 3389
rect 20619 3340 20628 3380
rect 20668 3340 20677 3380
rect 20619 3339 20677 3340
rect 21483 3371 21525 3380
rect 21483 3331 21484 3371
rect 21524 3331 21525 3371
rect 21771 3340 21772 3380
rect 21812 3340 21813 3380
rect 21771 3331 21813 3340
rect 24267 3380 24309 3389
rect 24267 3340 24268 3380
rect 24308 3340 24309 3380
rect 24267 3331 24309 3340
rect 25507 3380 25565 3381
rect 25507 3340 25516 3380
rect 25556 3340 25565 3380
rect 25507 3339 25565 3340
rect 26187 3380 26229 3389
rect 26187 3340 26188 3380
rect 26228 3340 26229 3380
rect 26187 3331 26229 3340
rect 26434 3380 26492 3381
rect 26434 3340 26443 3380
rect 26483 3340 26492 3380
rect 26434 3339 26492 3340
rect 26555 3380 26613 3381
rect 26555 3340 26564 3380
rect 26604 3340 26613 3380
rect 26555 3339 26613 3340
rect 28011 3380 28053 3389
rect 28011 3340 28012 3380
rect 28052 3340 28053 3380
rect 28011 3331 28053 3340
rect 29251 3380 29309 3381
rect 29251 3340 29260 3380
rect 29300 3340 29309 3380
rect 29251 3339 29309 3340
rect 30682 3380 30740 3381
rect 30682 3340 30691 3380
rect 30731 3340 30740 3380
rect 30682 3339 30740 3340
rect 30795 3380 30837 3389
rect 30795 3340 30796 3380
rect 30836 3340 30837 3380
rect 30795 3331 30837 3340
rect 31275 3380 31317 3389
rect 31275 3340 31276 3380
rect 31316 3340 31317 3380
rect 31275 3331 31317 3340
rect 31747 3380 31805 3381
rect 31747 3340 31756 3380
rect 31796 3340 31805 3380
rect 31747 3339 31805 3340
rect 32266 3380 32324 3381
rect 32266 3340 32275 3380
rect 32315 3340 32324 3380
rect 32266 3339 32324 3340
rect 32458 3380 32516 3381
rect 32458 3340 32467 3380
rect 32507 3340 32516 3380
rect 32458 3339 32516 3340
rect 21483 3322 21525 3331
rect 15675 3296 15717 3305
rect 15675 3256 15676 3296
rect 15716 3256 15717 3296
rect 15675 3247 15717 3256
rect 21387 3296 21429 3305
rect 21387 3256 21388 3296
rect 21428 3256 21429 3296
rect 21387 3247 21429 3256
rect 25707 3296 25749 3305
rect 25707 3256 25708 3296
rect 25748 3256 25749 3296
rect 25707 3247 25749 3256
rect 33339 3296 33381 3305
rect 33339 3256 33340 3296
rect 33380 3256 33381 3296
rect 33339 3247 33381 3256
rect 38427 3296 38469 3305
rect 38427 3256 38428 3296
rect 38468 3256 38469 3296
rect 38427 3247 38469 3256
rect 39579 3296 39621 3305
rect 39579 3256 39580 3296
rect 39620 3256 39621 3296
rect 39579 3247 39621 3256
rect 43515 3296 43557 3305
rect 43515 3256 43516 3296
rect 43556 3256 43557 3296
rect 43515 3247 43557 3256
rect 44763 3296 44805 3305
rect 44763 3256 44764 3296
rect 44804 3256 44805 3296
rect 44763 3247 44805 3256
rect 15243 3212 15285 3221
rect 15243 3172 15244 3212
rect 15284 3172 15285 3212
rect 15243 3163 15285 3172
rect 17643 3212 17685 3221
rect 17643 3172 17644 3212
rect 17684 3172 17685 3212
rect 17643 3163 17685 3172
rect 18555 3212 18597 3221
rect 18555 3172 18556 3212
rect 18596 3172 18597 3212
rect 18555 3163 18597 3172
rect 20811 3212 20853 3221
rect 20811 3172 20812 3212
rect 20852 3172 20853 3212
rect 20811 3163 20853 3172
rect 30459 3212 30501 3221
rect 30459 3172 30460 3212
rect 30500 3172 30501 3212
rect 30459 3163 30501 3172
rect 37018 3212 37076 3213
rect 37018 3172 37027 3212
rect 37067 3172 37076 3212
rect 37018 3171 37076 3172
rect 37306 3212 37364 3213
rect 37306 3172 37315 3212
rect 37355 3172 37364 3212
rect 37306 3171 37364 3172
rect 37594 3212 37652 3213
rect 37594 3172 37603 3212
rect 37643 3172 37652 3212
rect 37594 3171 37652 3172
rect 38043 3212 38085 3221
rect 38043 3172 38044 3212
rect 38084 3172 38085 3212
rect 38043 3163 38085 3172
rect 39034 3212 39092 3213
rect 39034 3172 39043 3212
rect 39083 3172 39092 3212
rect 39034 3171 39092 3172
rect 39963 3212 40005 3221
rect 39963 3172 39964 3212
rect 40004 3172 40005 3212
rect 39963 3163 40005 3172
rect 1152 3044 45216 3068
rect 1152 3004 4928 3044
rect 4968 3004 5010 3044
rect 5050 3004 5092 3044
rect 5132 3004 5174 3044
rect 5214 3004 5256 3044
rect 5296 3004 20048 3044
rect 20088 3004 20130 3044
rect 20170 3004 20212 3044
rect 20252 3004 20294 3044
rect 20334 3004 20376 3044
rect 20416 3004 35168 3044
rect 35208 3004 35250 3044
rect 35290 3004 35332 3044
rect 35372 3004 35414 3044
rect 35454 3004 35496 3044
rect 35536 3004 45216 3044
rect 1152 2980 45216 3004
rect 9195 2876 9237 2885
rect 9195 2836 9196 2876
rect 9236 2836 9237 2876
rect 9195 2827 9237 2836
rect 10923 2876 10965 2885
rect 10923 2836 10924 2876
rect 10964 2836 10965 2876
rect 10923 2827 10965 2836
rect 14043 2876 14085 2885
rect 14043 2836 14044 2876
rect 14084 2836 14085 2876
rect 14043 2827 14085 2836
rect 20187 2876 20229 2885
rect 20187 2836 20188 2876
rect 20228 2836 20229 2876
rect 20187 2827 20229 2836
rect 24507 2876 24549 2885
rect 24507 2836 24508 2876
rect 24548 2836 24549 2876
rect 24507 2827 24549 2836
rect 45147 2876 45189 2885
rect 45147 2836 45148 2876
rect 45188 2836 45189 2876
rect 45147 2827 45189 2836
rect 15915 2792 15957 2801
rect 15915 2752 15916 2792
rect 15956 2752 15957 2792
rect 15915 2743 15957 2752
rect 31803 2792 31845 2801
rect 31803 2752 31804 2792
rect 31844 2752 31845 2792
rect 31803 2743 31845 2752
rect 37515 2792 37557 2801
rect 37515 2752 37516 2792
rect 37556 2752 37557 2792
rect 37515 2743 37557 2752
rect 37803 2792 37845 2801
rect 37803 2752 37804 2792
rect 37844 2752 37845 2792
rect 37803 2743 37845 2752
rect 38091 2792 38133 2801
rect 38091 2752 38092 2792
rect 38132 2752 38133 2792
rect 38091 2743 38133 2752
rect 38379 2792 38421 2801
rect 38379 2752 38380 2792
rect 38420 2752 38421 2792
rect 38379 2743 38421 2752
rect 38667 2792 38709 2801
rect 38667 2752 38668 2792
rect 38708 2752 38709 2792
rect 38667 2743 38709 2752
rect 7755 2708 7797 2717
rect 9483 2708 9525 2717
rect 15531 2708 15573 2717
rect 7755 2668 7756 2708
rect 7796 2668 7797 2708
rect 7755 2659 7797 2668
rect 9003 2699 9045 2708
rect 9003 2659 9004 2699
rect 9044 2659 9045 2699
rect 9483 2668 9484 2708
rect 9524 2668 9525 2708
rect 9483 2659 9525 2668
rect 10731 2699 10773 2708
rect 10731 2659 10732 2699
rect 10772 2659 10773 2699
rect 15531 2668 15532 2708
rect 15572 2668 15573 2708
rect 15531 2659 15573 2668
rect 15802 2708 15860 2709
rect 15802 2668 15811 2708
rect 15851 2668 15860 2708
rect 15802 2667 15860 2668
rect 18202 2708 18260 2709
rect 18202 2668 18211 2708
rect 18251 2668 18260 2708
rect 18202 2667 18260 2668
rect 18315 2708 18357 2717
rect 18315 2668 18316 2708
rect 18356 2668 18357 2708
rect 18315 2659 18357 2668
rect 18699 2708 18741 2717
rect 19978 2708 20036 2709
rect 18699 2668 18700 2708
rect 18740 2668 18741 2708
rect 18699 2659 18741 2668
rect 19275 2699 19317 2708
rect 19275 2659 19276 2699
rect 19316 2659 19317 2699
rect 9003 2650 9045 2659
rect 10731 2650 10773 2659
rect 19275 2650 19317 2659
rect 19755 2699 19797 2708
rect 19755 2659 19756 2699
rect 19796 2659 19797 2699
rect 19978 2668 19987 2708
rect 20027 2668 20036 2708
rect 19978 2667 20036 2668
rect 19755 2650 19797 2659
rect 7371 2624 7413 2633
rect 7371 2584 7372 2624
rect 7412 2584 7413 2624
rect 7371 2575 7413 2584
rect 13803 2624 13845 2633
rect 13803 2584 13804 2624
rect 13844 2584 13845 2624
rect 13803 2575 13845 2584
rect 18795 2624 18837 2633
rect 18795 2584 18796 2624
rect 18836 2584 18837 2624
rect 18795 2575 18837 2584
rect 20427 2624 20469 2633
rect 20427 2584 20428 2624
rect 20468 2584 20469 2624
rect 20427 2575 20469 2584
rect 24267 2624 24309 2633
rect 24267 2584 24268 2624
rect 24308 2584 24309 2624
rect 24267 2575 24309 2584
rect 31275 2624 31317 2633
rect 31275 2584 31276 2624
rect 31316 2584 31317 2624
rect 31275 2575 31317 2584
rect 31659 2624 31701 2633
rect 31659 2584 31660 2624
rect 31700 2584 31701 2624
rect 31659 2575 31701 2584
rect 32043 2624 32085 2633
rect 32043 2584 32044 2624
rect 32084 2584 32085 2624
rect 32043 2575 32085 2584
rect 36363 2624 36405 2633
rect 36363 2584 36364 2624
rect 36404 2584 36405 2624
rect 36363 2575 36405 2584
rect 39243 2624 39285 2633
rect 39243 2584 39244 2624
rect 39284 2584 39285 2624
rect 39243 2575 39285 2584
rect 39531 2624 39573 2633
rect 39531 2584 39532 2624
rect 39572 2584 39573 2624
rect 39531 2575 39573 2584
rect 39723 2624 39765 2633
rect 39723 2584 39724 2624
rect 39764 2584 39765 2624
rect 39723 2575 39765 2584
rect 40107 2624 40149 2633
rect 40107 2584 40108 2624
rect 40148 2584 40149 2624
rect 40107 2575 40149 2584
rect 40491 2624 40533 2633
rect 40491 2584 40492 2624
rect 40532 2584 40533 2624
rect 40491 2575 40533 2584
rect 40875 2624 40917 2633
rect 40875 2584 40876 2624
rect 40916 2584 40917 2624
rect 40875 2575 40917 2584
rect 41163 2624 41205 2633
rect 41163 2584 41164 2624
rect 41204 2584 41205 2624
rect 41163 2575 41205 2584
rect 43083 2624 43125 2633
rect 43083 2584 43084 2624
rect 43124 2584 43125 2624
rect 43083 2575 43125 2584
rect 44139 2624 44181 2633
rect 44139 2584 44140 2624
rect 44180 2584 44181 2624
rect 44139 2575 44181 2584
rect 44379 2624 44421 2633
rect 44379 2584 44380 2624
rect 44420 2584 44421 2624
rect 44379 2575 44421 2584
rect 44523 2624 44565 2633
rect 44523 2584 44524 2624
rect 44564 2584 44565 2624
rect 44523 2575 44565 2584
rect 44907 2624 44949 2633
rect 44907 2584 44908 2624
rect 44948 2584 44949 2624
rect 44907 2575 44949 2584
rect 39963 2540 40005 2549
rect 39963 2500 39964 2540
rect 40004 2500 40005 2540
rect 39963 2491 40005 2500
rect 44763 2540 44805 2549
rect 44763 2500 44764 2540
rect 44804 2500 44805 2540
rect 44763 2491 44805 2500
rect 7611 2456 7653 2465
rect 7611 2416 7612 2456
rect 7652 2416 7653 2456
rect 7611 2407 7653 2416
rect 16203 2456 16245 2465
rect 16203 2416 16204 2456
rect 16244 2416 16245 2456
rect 16203 2407 16245 2416
rect 31035 2456 31077 2465
rect 31035 2416 31036 2456
rect 31076 2416 31077 2456
rect 31035 2407 31077 2416
rect 31419 2456 31461 2465
rect 31419 2416 31420 2456
rect 31460 2416 31461 2456
rect 31419 2407 31461 2416
rect 36603 2456 36645 2465
rect 36603 2416 36604 2456
rect 36644 2416 36645 2456
rect 36603 2407 36645 2416
rect 40347 2456 40389 2465
rect 40347 2416 40348 2456
rect 40388 2416 40389 2456
rect 40347 2407 40389 2416
rect 40731 2456 40773 2465
rect 40731 2416 40732 2456
rect 40772 2416 40773 2456
rect 40731 2407 40773 2416
rect 42843 2456 42885 2465
rect 42843 2416 42844 2456
rect 42884 2416 42885 2456
rect 42843 2407 42885 2416
rect 1152 2288 45216 2312
rect 1152 2248 3688 2288
rect 3728 2248 3770 2288
rect 3810 2248 3852 2288
rect 3892 2248 3934 2288
rect 3974 2248 4016 2288
rect 4056 2248 18808 2288
rect 18848 2248 18890 2288
rect 18930 2248 18972 2288
rect 19012 2248 19054 2288
rect 19094 2248 19136 2288
rect 19176 2248 33928 2288
rect 33968 2248 34010 2288
rect 34050 2248 34092 2288
rect 34132 2248 34174 2288
rect 34214 2248 34256 2288
rect 34296 2248 45216 2288
rect 1152 2224 45216 2248
rect 4251 2120 4293 2129
rect 4251 2080 4252 2120
rect 4292 2080 4293 2120
rect 4251 2071 4293 2080
rect 9627 2120 9669 2129
rect 9627 2080 9628 2120
rect 9668 2080 9669 2120
rect 9627 2071 9669 2080
rect 45147 2120 45189 2129
rect 45147 2080 45148 2120
rect 45188 2080 45189 2120
rect 45147 2071 45189 2080
rect 2715 2036 2757 2045
rect 2715 1996 2716 2036
rect 2756 1996 2757 2036
rect 2715 1987 2757 1996
rect 43227 2036 43269 2045
rect 43227 1996 43228 2036
rect 43268 1996 43269 2036
rect 43227 1987 43269 1996
rect 2475 1952 2517 1961
rect 2475 1912 2476 1952
rect 2516 1912 2517 1952
rect 2475 1903 2517 1912
rect 4011 1952 4053 1961
rect 4011 1912 4012 1952
rect 4052 1912 4053 1952
rect 4011 1903 4053 1912
rect 5739 1952 5781 1961
rect 5739 1912 5740 1952
rect 5780 1912 5781 1952
rect 5739 1903 5781 1912
rect 7275 1952 7317 1961
rect 7275 1912 7276 1952
rect 7316 1912 7317 1952
rect 7275 1903 7317 1912
rect 8811 1952 8853 1961
rect 8811 1912 8812 1952
rect 8852 1912 8853 1952
rect 8811 1903 8853 1912
rect 9387 1952 9429 1961
rect 9387 1912 9388 1952
rect 9428 1912 9429 1952
rect 9387 1903 9429 1912
rect 10347 1952 10389 1961
rect 10347 1912 10348 1952
rect 10388 1912 10389 1952
rect 10347 1903 10389 1912
rect 11883 1952 11925 1961
rect 11883 1912 11884 1952
rect 11924 1912 11925 1952
rect 11883 1903 11925 1912
rect 18795 1952 18837 1961
rect 18795 1912 18796 1952
rect 18836 1912 18837 1952
rect 18795 1903 18837 1912
rect 39243 1952 39285 1961
rect 39243 1912 39244 1952
rect 39284 1912 39285 1952
rect 39243 1903 39285 1912
rect 40107 1952 40149 1961
rect 40107 1912 40108 1952
rect 40148 1912 40149 1952
rect 40107 1903 40149 1912
rect 42987 1952 43029 1961
rect 42987 1912 42988 1952
rect 43028 1912 43029 1952
rect 42987 1903 43029 1912
rect 43371 1952 43413 1961
rect 43371 1912 43372 1952
rect 43412 1912 43413 1952
rect 43371 1903 43413 1912
rect 43755 1952 43797 1961
rect 43755 1912 43756 1952
rect 43796 1912 43797 1952
rect 43755 1903 43797 1912
rect 44139 1952 44181 1961
rect 44139 1912 44140 1952
rect 44180 1912 44181 1952
rect 44139 1903 44181 1912
rect 44523 1952 44565 1961
rect 44523 1912 44524 1952
rect 44564 1912 44565 1952
rect 44523 1903 44565 1912
rect 44907 1952 44949 1961
rect 44907 1912 44908 1952
rect 44948 1912 44949 1952
rect 44907 1903 44949 1912
rect 40299 1868 40341 1877
rect 40299 1828 40300 1868
rect 40340 1828 40341 1868
rect 40299 1819 40341 1828
rect 43995 1784 44037 1793
rect 43995 1744 43996 1784
rect 44036 1744 44037 1784
rect 43995 1735 44037 1744
rect 5499 1700 5541 1709
rect 5499 1660 5500 1700
rect 5540 1660 5541 1700
rect 5499 1651 5541 1660
rect 7035 1700 7077 1709
rect 7035 1660 7036 1700
rect 7076 1660 7077 1700
rect 7035 1651 7077 1660
rect 8571 1700 8613 1709
rect 8571 1660 8572 1700
rect 8612 1660 8613 1700
rect 8571 1651 8613 1660
rect 10107 1700 10149 1709
rect 10107 1660 10108 1700
rect 10148 1660 10149 1700
rect 10107 1651 10149 1660
rect 11643 1700 11685 1709
rect 11643 1660 11644 1700
rect 11684 1660 11685 1700
rect 11643 1651 11685 1660
rect 18555 1700 18597 1709
rect 18555 1660 18556 1700
rect 18596 1660 18597 1700
rect 18555 1651 18597 1660
rect 39147 1700 39189 1709
rect 39147 1660 39148 1700
rect 39188 1660 39189 1700
rect 39147 1651 39189 1660
rect 39418 1700 39476 1701
rect 39418 1660 39427 1700
rect 39467 1660 39476 1700
rect 39418 1659 39476 1660
rect 39706 1700 39764 1701
rect 39706 1660 39715 1700
rect 39755 1660 39764 1700
rect 39706 1659 39764 1660
rect 40570 1700 40628 1701
rect 40570 1660 40579 1700
rect 40619 1660 40628 1700
rect 40570 1659 40628 1660
rect 43611 1700 43653 1709
rect 43611 1660 43612 1700
rect 43652 1660 43653 1700
rect 43611 1651 43653 1660
rect 44379 1700 44421 1709
rect 44379 1660 44380 1700
rect 44420 1660 44421 1700
rect 44379 1651 44421 1660
rect 44763 1700 44805 1709
rect 44763 1660 44764 1700
rect 44804 1660 44805 1700
rect 44763 1651 44805 1660
rect 1152 1532 45216 1556
rect 1152 1492 4928 1532
rect 4968 1492 5010 1532
rect 5050 1492 5092 1532
rect 5132 1492 5174 1532
rect 5214 1492 5256 1532
rect 5296 1492 20048 1532
rect 20088 1492 20130 1532
rect 20170 1492 20212 1532
rect 20252 1492 20294 1532
rect 20334 1492 20376 1532
rect 20416 1492 35168 1532
rect 35208 1492 35250 1532
rect 35290 1492 35332 1532
rect 35372 1492 35414 1532
rect 35454 1492 35496 1532
rect 35536 1492 45216 1532
rect 1152 1468 45216 1492
<< via1 >>
rect 3688 9808 3728 9848
rect 3770 9808 3810 9848
rect 3852 9808 3892 9848
rect 3934 9808 3974 9848
rect 4016 9808 4056 9848
rect 18808 9808 18848 9848
rect 18890 9808 18930 9848
rect 18972 9808 19012 9848
rect 19054 9808 19094 9848
rect 19136 9808 19176 9848
rect 33928 9808 33968 9848
rect 34010 9808 34050 9848
rect 34092 9808 34132 9848
rect 34174 9808 34214 9848
rect 34256 9808 34296 9848
rect 2236 9640 2276 9680
rect 10204 9640 10244 9680
rect 11356 9640 11396 9680
rect 12124 9640 12164 9680
rect 12892 9640 12932 9680
rect 13276 9640 13316 9680
rect 14044 9640 14084 9680
rect 14812 9640 14852 9680
rect 15196 9640 15236 9680
rect 15580 9640 15620 9680
rect 15964 9640 16004 9680
rect 16348 9640 16388 9680
rect 16732 9640 16772 9680
rect 17116 9640 17156 9680
rect 17500 9640 17540 9680
rect 17884 9640 17924 9680
rect 18268 9640 18308 9680
rect 18652 9640 18692 9680
rect 19804 9640 19844 9680
rect 20188 9640 20228 9680
rect 20572 9640 20612 9680
rect 21340 9640 21380 9680
rect 25852 9640 25892 9680
rect 27388 9640 27428 9680
rect 31228 9640 31268 9680
rect 31996 9640 32036 9680
rect 34300 9640 34340 9680
rect 34684 9640 34724 9680
rect 35836 9640 35876 9680
rect 42844 9640 42884 9680
rect 43996 9640 44036 9680
rect 44380 9640 44420 9680
rect 44764 9640 44804 9680
rect 10588 9556 10628 9596
rect 11740 9556 11780 9596
rect 12508 9556 12548 9596
rect 13660 9556 13700 9596
rect 14428 9556 14468 9596
rect 19036 9556 19076 9596
rect 28828 9556 28868 9596
rect 31612 9556 31652 9596
rect 32380 9556 32420 9596
rect 33532 9556 33572 9596
rect 35452 9556 35492 9596
rect 1228 9472 1268 9512
rect 1612 9472 1652 9512
rect 1996 9472 2036 9512
rect 2380 9472 2420 9512
rect 2764 9472 2804 9512
rect 3148 9472 3188 9512
rect 9964 9472 10004 9512
rect 10348 9472 10388 9512
rect 10732 9472 10772 9512
rect 11116 9472 11156 9512
rect 11500 9472 11540 9512
rect 11884 9472 11924 9512
rect 12268 9472 12308 9512
rect 12652 9472 12692 9512
rect 13036 9472 13076 9512
rect 13420 9472 13460 9512
rect 13804 9472 13844 9512
rect 14188 9472 14228 9512
rect 14572 9472 14612 9512
rect 14956 9472 14996 9512
rect 15340 9472 15380 9512
rect 15724 9472 15764 9512
rect 16108 9472 16148 9512
rect 16492 9472 16532 9512
rect 16876 9472 16916 9512
rect 17260 9472 17300 9512
rect 17644 9472 17684 9512
rect 18028 9472 18068 9512
rect 18412 9472 18452 9512
rect 18796 9472 18836 9512
rect 19180 9472 19220 9512
rect 19603 9472 19643 9512
rect 19948 9472 19988 9512
rect 20332 9472 20372 9512
rect 20908 9472 20948 9512
rect 21100 9472 21140 9512
rect 21676 9472 21716 9512
rect 21868 9472 21908 9512
rect 22252 9472 22292 9512
rect 22828 9472 22868 9512
rect 23212 9472 23252 9512
rect 23596 9472 23636 9512
rect 24172 9472 24212 9512
rect 24556 9472 24596 9512
rect 24748 9472 24788 9512
rect 25132 9472 25172 9512
rect 25708 9472 25748 9512
rect 26092 9472 26132 9512
rect 26284 9472 26324 9512
rect 26860 9472 26900 9512
rect 27052 9472 27092 9512
rect 27628 9472 27668 9512
rect 28396 9472 28436 9512
rect 28588 9472 28628 9512
rect 29164 9472 29204 9512
rect 29548 9472 29588 9512
rect 29932 9472 29972 9512
rect 30316 9472 30356 9512
rect 31468 9472 31508 9512
rect 31852 9472 31892 9512
rect 32236 9472 32276 9512
rect 32620 9472 32660 9512
rect 33004 9472 33044 9512
rect 33388 9472 33428 9512
rect 33772 9472 33812 9512
rect 34156 9472 34196 9512
rect 34540 9472 34580 9512
rect 34924 9472 34964 9512
rect 35308 9472 35348 9512
rect 35692 9472 35732 9512
rect 36076 9472 36116 9512
rect 42220 9472 42260 9512
rect 42604 9472 42644 9512
rect 43084 9472 43124 9512
rect 43468 9472 43508 9512
rect 43756 9472 43796 9512
rect 44140 9472 44180 9512
rect 44524 9472 44564 9512
rect 44908 9472 44948 9512
rect 2620 9304 2660 9344
rect 3004 9304 3044 9344
rect 10972 9304 11012 9344
rect 19420 9304 19460 9344
rect 22492 9304 22532 9344
rect 23452 9304 23492 9344
rect 23836 9304 23876 9344
rect 24988 9304 25028 9344
rect 25372 9304 25412 9344
rect 26524 9304 26564 9344
rect 27292 9304 27332 9344
rect 32764 9304 32804 9344
rect 33148 9304 33188 9344
rect 35068 9304 35108 9344
rect 45148 9304 45188 9344
rect 1468 9220 1508 9260
rect 1852 9220 1892 9260
rect 3388 9220 3428 9260
rect 20668 9220 20708 9260
rect 21436 9220 21476 9260
rect 22108 9220 22148 9260
rect 22588 9220 22628 9260
rect 23932 9220 23972 9260
rect 24316 9220 24356 9260
rect 25468 9220 25508 9260
rect 26620 9220 26660 9260
rect 28156 9220 28196 9260
rect 28924 9220 28964 9260
rect 29308 9220 29348 9260
rect 29692 9220 29732 9260
rect 30076 9220 30116 9260
rect 33916 9220 33956 9260
rect 41923 9220 41963 9260
rect 42460 9220 42500 9260
rect 43324 9220 43364 9260
rect 43459 9220 43499 9260
rect 4928 9052 4968 9092
rect 5010 9052 5050 9092
rect 5092 9052 5132 9092
rect 5174 9052 5214 9092
rect 5256 9052 5296 9092
rect 20048 9052 20088 9092
rect 20130 9052 20170 9092
rect 20212 9052 20252 9092
rect 20294 9052 20334 9092
rect 20376 9052 20416 9092
rect 35168 9052 35208 9092
rect 35250 9052 35290 9092
rect 35332 9052 35372 9092
rect 35414 9052 35454 9092
rect 35496 9052 35536 9092
rect 1468 8884 1508 8924
rect 9916 8884 9956 8924
rect 10684 8884 10724 8924
rect 11452 8884 11492 8924
rect 11923 8884 11963 8924
rect 12220 8884 12260 8924
rect 12604 8884 12644 8924
rect 12988 8884 13028 8924
rect 13372 8884 13412 8924
rect 13756 8884 13796 8924
rect 14524 8884 14564 8924
rect 15292 8884 15332 8924
rect 15676 8884 15716 8924
rect 16060 8884 16100 8924
rect 16444 8884 16484 8924
rect 16828 8884 16868 8924
rect 17212 8884 17252 8924
rect 17596 8884 17636 8924
rect 17980 8884 18020 8924
rect 18364 8884 18404 8924
rect 18748 8884 18788 8924
rect 19132 8884 19172 8924
rect 19516 8884 19556 8924
rect 20284 8884 20324 8924
rect 21100 8884 21140 8924
rect 32188 8884 32228 8924
rect 32572 8884 32612 8924
rect 32956 8884 32996 8924
rect 33340 8884 33380 8924
rect 33724 8884 33764 8924
rect 34108 8884 34148 8924
rect 34876 8884 34916 8924
rect 43516 8884 43556 8924
rect 44380 8884 44420 8924
rect 10300 8800 10340 8840
rect 20668 8800 20708 8840
rect 21724 8800 21764 8840
rect 23548 8800 23588 8840
rect 25660 8800 25700 8840
rect 28252 8800 28292 8840
rect 29404 8800 29444 8840
rect 34492 8800 34532 8840
rect 42364 8800 42404 8840
rect 42748 8800 42788 8840
rect 11596 8716 11636 8756
rect 11724 8692 11764 8732
rect 27628 8716 27668 8756
rect 27757 8716 27797 8756
rect 28012 8716 28052 8756
rect 1228 8632 1268 8672
rect 1612 8632 1652 8672
rect 1852 8632 1892 8672
rect 1996 8632 2036 8672
rect 2236 8632 2276 8672
rect 2380 8632 2420 8672
rect 2620 8632 2660 8672
rect 9676 8632 9716 8672
rect 10060 8632 10100 8672
rect 10444 8632 10484 8672
rect 10828 8632 10868 8672
rect 11212 8632 11252 8672
rect 12460 8632 12500 8672
rect 12844 8632 12884 8672
rect 13228 8632 13268 8672
rect 13612 8632 13652 8672
rect 13996 8632 14036 8672
rect 14380 8632 14420 8672
rect 14764 8632 14804 8672
rect 14956 8632 14996 8672
rect 15196 8632 15236 8672
rect 15532 8632 15572 8672
rect 15916 8632 15956 8672
rect 16300 8632 16340 8672
rect 16684 8632 16724 8672
rect 17068 8632 17108 8672
rect 17452 8632 17492 8672
rect 17836 8632 17876 8672
rect 18220 8632 18260 8672
rect 18604 8632 18644 8672
rect 18988 8632 19028 8672
rect 19372 8632 19412 8672
rect 19756 8632 19796 8672
rect 19900 8632 19940 8672
rect 20140 8632 20180 8672
rect 20524 8632 20564 8672
rect 20908 8632 20948 8672
rect 21484 8632 21524 8672
rect 22060 8632 22100 8672
rect 23788 8632 23828 8672
rect 25324 8632 25364 8672
rect 25900 8632 25940 8672
rect 26092 8632 26132 8672
rect 26428 8632 26468 8672
rect 26668 8632 26708 8672
rect 26812 8632 26852 8672
rect 27052 8632 27092 8672
rect 28492 8632 28532 8672
rect 29164 8632 29204 8672
rect 29740 8632 29780 8672
rect 32428 8632 32468 8672
rect 32812 8632 32852 8672
rect 33196 8632 33236 8672
rect 33580 8632 33620 8672
rect 33964 8632 34004 8672
rect 34348 8632 34388 8672
rect 34732 8632 34772 8672
rect 35116 8632 35156 8672
rect 42604 8632 42644 8672
rect 42988 8632 43028 8672
rect 43132 8632 43172 8672
rect 43372 8632 43412 8672
rect 43756 8632 43796 8672
rect 44140 8632 44180 8672
rect 44524 8632 44564 8672
rect 44908 8632 44948 8672
rect 11068 8548 11108 8588
rect 21820 8548 21860 8588
rect 25564 8548 25604 8588
rect 26332 8548 26372 8588
rect 14140 8464 14180 8504
rect 27340 8464 27380 8504
rect 29500 8464 29540 8504
rect 44764 8464 44804 8504
rect 45148 8464 45188 8504
rect 3688 8296 3728 8336
rect 3770 8296 3810 8336
rect 3852 8296 3892 8336
rect 3934 8296 3974 8336
rect 4016 8296 4056 8336
rect 18808 8296 18848 8336
rect 18890 8296 18930 8336
rect 18972 8296 19012 8336
rect 19054 8296 19094 8336
rect 19136 8296 19176 8336
rect 33928 8296 33968 8336
rect 34010 8296 34050 8336
rect 34092 8296 34132 8336
rect 34174 8296 34214 8336
rect 34256 8296 34296 8336
rect 17884 8128 17924 8168
rect 22876 8128 22916 8168
rect 28252 8128 28292 8168
rect 28636 8128 28676 8168
rect 32092 8128 32132 8168
rect 34492 8128 34532 8168
rect 34972 8128 35012 8168
rect 36700 8128 36740 8168
rect 42748 8128 42788 8168
rect 43132 8128 43172 8168
rect 43900 8128 43940 8168
rect 24844 8044 24884 8084
rect 34876 8044 34916 8084
rect 1228 7960 1268 8000
rect 1612 7960 1652 8000
rect 2476 7960 2516 8000
rect 2716 7960 2756 8000
rect 2860 7960 2900 8000
rect 3244 7960 3284 8000
rect 3484 7960 3524 8000
rect 3628 7960 3668 8000
rect 4012 7960 4052 8000
rect 4396 7960 4436 8000
rect 10252 7960 10292 8000
rect 14476 7960 14516 8000
rect 16972 7960 17012 8000
rect 18124 7960 18164 8000
rect 22636 7960 22676 8000
rect 23020 7960 23060 8000
rect 26092 7960 26132 8000
rect 26860 7960 26900 8000
rect 28492 7960 28532 8000
rect 28876 7960 28916 8000
rect 29452 7960 29492 8000
rect 31564 7960 31604 8000
rect 31852 7960 31892 8000
rect 32428 7960 32468 8000
rect 32716 7960 32756 8000
rect 33196 7960 33236 8000
rect 33484 7960 33524 8000
rect 33868 7960 33908 8000
rect 34252 7960 34292 8000
rect 34636 7960 34676 8000
rect 35212 7960 35252 8000
rect 36499 7960 36539 8000
rect 41836 7960 41876 8000
rect 41980 7960 42020 8000
rect 42220 7960 42260 8000
rect 42604 7960 42644 8000
rect 42988 7960 43028 8000
rect 43372 7960 43412 8000
rect 43756 7960 43796 8000
rect 44140 7960 44180 8000
rect 44524 7960 44564 8000
rect 44908 7960 44948 8000
rect 9763 7876 9803 7916
rect 9868 7876 9908 7916
rect 10348 7876 10388 7916
rect 10828 7876 10868 7916
rect 11316 7876 11356 7916
rect 11788 7876 11828 7916
rect 12067 7876 12107 7916
rect 12604 7876 12644 7916
rect 12748 7876 12788 7916
rect 14860 7876 14900 7916
rect 16108 7876 16148 7916
rect 23404 7876 23444 7916
rect 24652 7876 24692 7916
rect 26371 7876 26411 7916
rect 26476 7876 26516 7916
rect 26956 7876 26996 7916
rect 27436 7876 27476 7916
rect 27955 7876 27995 7916
rect 1852 7792 1892 7832
rect 3100 7792 3140 7832
rect 12172 7792 12212 7832
rect 41596 7792 41636 7832
rect 43516 7792 43556 7832
rect 1468 7708 1508 7748
rect 3868 7708 3908 7748
rect 4252 7708 4292 7748
rect 4636 7708 4676 7748
rect 11500 7708 11540 7748
rect 12508 7708 12548 7748
rect 14716 7708 14756 7748
rect 16300 7708 16340 7748
rect 17212 7708 17252 7748
rect 23260 7708 23300 7748
rect 25852 7708 25892 7748
rect 28108 7708 28148 7748
rect 29692 7708 29732 7748
rect 31651 7708 31691 7748
rect 32419 7708 32459 7748
rect 32956 7708 32996 7748
rect 33187 7708 33227 7748
rect 33724 7708 33764 7748
rect 34108 7708 34148 7748
rect 36259 7708 36299 7748
rect 36835 7708 36875 7748
rect 42364 7708 42404 7748
rect 44764 7708 44804 7748
rect 45148 7708 45188 7748
rect 4928 7540 4968 7580
rect 5010 7540 5050 7580
rect 5092 7540 5132 7580
rect 5174 7540 5214 7580
rect 5256 7540 5296 7580
rect 20048 7540 20088 7580
rect 20130 7540 20170 7580
rect 20212 7540 20252 7580
rect 20294 7540 20334 7580
rect 20376 7540 20416 7580
rect 35168 7540 35208 7580
rect 35250 7540 35290 7580
rect 35332 7540 35372 7580
rect 35414 7540 35454 7580
rect 35496 7540 35536 7580
rect 11779 7372 11819 7412
rect 12547 7372 12587 7412
rect 28012 7372 28052 7412
rect 33091 7372 33131 7412
rect 33379 7372 33419 7412
rect 33955 7372 33995 7412
rect 34531 7372 34571 7412
rect 35107 7372 35147 7412
rect 35683 7372 35723 7412
rect 36163 7372 36203 7412
rect 44035 7372 44075 7412
rect 44620 7372 44660 7412
rect 10540 7288 10580 7328
rect 12652 7288 12692 7328
rect 29164 7288 29204 7328
rect 36748 7288 36788 7328
rect 37612 7288 37652 7328
rect 10156 7204 10196 7244
rect 10435 7204 10475 7244
rect 11708 7193 11748 7233
rect 11875 7204 11915 7244
rect 11992 7204 12032 7244
rect 12124 7195 12164 7235
rect 12257 7193 12297 7233
rect 12451 7204 12491 7244
rect 12759 7204 12799 7244
rect 13036 7204 13076 7244
rect 14860 7204 14900 7244
rect 16108 7195 16148 7235
rect 23308 7204 23348 7244
rect 24556 7195 24596 7235
rect 26275 7204 26315 7244
rect 26385 7204 26425 7244
rect 26764 7204 26804 7244
rect 27340 7195 27380 7235
rect 27820 7195 27860 7235
rect 29356 7195 29396 7235
rect 30604 7204 30644 7244
rect 32716 7204 32756 7244
rect 33004 7204 33044 7244
rect 33580 7204 33620 7244
rect 37900 7204 37940 7244
rect 1228 7120 1268 7160
rect 1612 7120 1652 7160
rect 1852 7120 1892 7160
rect 9676 7120 9716 7160
rect 11116 7120 11156 7160
rect 11356 7120 11396 7160
rect 12892 7120 12932 7160
rect 21676 7120 21716 7160
rect 26860 7120 26900 7160
rect 28396 7120 28436 7160
rect 32332 7120 32372 7160
rect 34156 7120 34196 7160
rect 34732 7120 34772 7160
rect 35308 7120 35348 7160
rect 35884 7120 35924 7160
rect 36460 7120 36500 7160
rect 37036 7120 37076 7160
rect 37324 7120 37364 7160
rect 41932 7120 41972 7160
rect 42316 7120 42356 7160
rect 42700 7120 42740 7160
rect 43084 7120 43124 7160
rect 43468 7120 43508 7160
rect 43756 7120 43796 7160
rect 44044 7120 44084 7160
rect 44236 7120 44276 7160
rect 44716 7120 44756 7160
rect 44908 7120 44948 7160
rect 1468 7036 1508 7076
rect 9916 7036 9956 7076
rect 10828 7036 10868 7076
rect 28156 7036 28196 7076
rect 42844 7036 42884 7076
rect 16300 6952 16340 6992
rect 21916 6952 21956 6992
rect 24748 6952 24788 6992
rect 32572 6952 32612 6992
rect 41692 6952 41732 6992
rect 42076 6952 42116 6992
rect 42460 6952 42500 6992
rect 43228 6952 43268 6992
rect 44476 6952 44516 6992
rect 45148 6952 45188 6992
rect 3688 6784 3728 6824
rect 3770 6784 3810 6824
rect 3852 6784 3892 6824
rect 3934 6784 3974 6824
rect 4016 6784 4056 6824
rect 18808 6784 18848 6824
rect 18890 6784 18930 6824
rect 18972 6784 19012 6824
rect 19054 6784 19094 6824
rect 19136 6784 19176 6824
rect 33928 6784 33968 6824
rect 34010 6784 34050 6824
rect 34092 6784 34132 6824
rect 34174 6784 34214 6824
rect 34256 6784 34296 6824
rect 7948 6616 7988 6656
rect 11251 6616 11291 6656
rect 1468 6532 1508 6572
rect 12172 6532 12212 6572
rect 1228 6448 1268 6488
rect 1612 6448 1652 6488
rect 6124 6448 6164 6488
rect 9004 6448 9044 6488
rect 9964 6448 10004 6488
rect 17164 6448 17204 6488
rect 44524 6448 44564 6488
rect 6508 6364 6548 6404
rect 7764 6364 7804 6404
rect 9475 6364 9515 6404
rect 9580 6364 9620 6404
rect 10060 6364 10100 6404
rect 10540 6364 10580 6404
rect 11059 6364 11099 6404
rect 11500 6364 11540 6404
rect 11779 6364 11819 6404
rect 11884 6280 11924 6320
rect 44908 6280 44948 6320
rect 1852 6196 1892 6236
rect 6364 6196 6404 6236
rect 9244 6196 9284 6236
rect 16924 6196 16964 6236
rect 43651 6196 43691 6236
rect 43939 6196 43979 6236
rect 44227 6196 44267 6236
rect 44764 6196 44804 6236
rect 4928 6028 4968 6068
rect 5010 6028 5050 6068
rect 5092 6028 5132 6068
rect 5174 6028 5214 6068
rect 5256 6028 5296 6068
rect 20048 6028 20088 6068
rect 20130 6028 20170 6068
rect 20212 6028 20252 6068
rect 20294 6028 20334 6068
rect 20376 6028 20416 6068
rect 35168 6028 35208 6068
rect 35250 6028 35290 6068
rect 35332 6028 35372 6068
rect 35414 6028 35454 6068
rect 35496 6028 35536 6068
rect 11116 5860 11156 5900
rect 13180 5860 13220 5900
rect 43747 5860 43787 5900
rect 44227 5860 44267 5900
rect 9379 5692 9419 5732
rect 9484 5692 9524 5732
rect 9868 5692 9908 5732
rect 10444 5683 10484 5723
rect 10924 5683 10964 5723
rect 13324 5692 13364 5732
rect 1228 5608 1268 5648
rect 1612 5608 1652 5648
rect 1996 5608 2036 5648
rect 9964 5608 10004 5648
rect 11308 5608 11348 5648
rect 11548 5608 11588 5648
rect 43660 5608 43700 5648
rect 44044 5608 44084 5648
rect 44524 5608 44564 5648
rect 44908 5608 44948 5648
rect 45148 5608 45188 5648
rect 1468 5440 1508 5480
rect 1852 5440 1892 5480
rect 2236 5440 2276 5480
rect 44764 5440 44804 5480
rect 3688 5272 3728 5312
rect 3770 5272 3810 5312
rect 3852 5272 3892 5312
rect 3934 5272 3974 5312
rect 4016 5272 4056 5312
rect 18808 5272 18848 5312
rect 18890 5272 18930 5312
rect 18972 5272 19012 5312
rect 19054 5272 19094 5312
rect 19136 5272 19176 5312
rect 33928 5272 33968 5312
rect 34010 5272 34050 5312
rect 34092 5272 34132 5312
rect 34174 5272 34214 5312
rect 34256 5272 34296 5312
rect 32956 5104 32996 5144
rect 42844 5104 42884 5144
rect 45148 5104 45188 5144
rect 30988 4936 31028 4976
rect 33196 4936 33236 4976
rect 43084 4936 43124 4976
rect 44524 4936 44564 4976
rect 44908 4936 44948 4976
rect 31372 4852 31412 4892
rect 32620 4852 32660 4892
rect 44236 4852 44276 4892
rect 31228 4684 31268 4724
rect 32812 4684 32852 4724
rect 43459 4684 43499 4724
rect 43651 4684 43691 4724
rect 43939 4684 43979 4724
rect 44764 4684 44804 4724
rect 4928 4516 4968 4556
rect 5010 4516 5050 4556
rect 5092 4516 5132 4556
rect 5174 4516 5214 4556
rect 5256 4516 5296 4556
rect 20048 4516 20088 4556
rect 20130 4516 20170 4556
rect 20212 4516 20252 4556
rect 20294 4516 20334 4556
rect 20376 4516 20416 4556
rect 35168 4516 35208 4556
rect 35250 4516 35290 4556
rect 35332 4516 35372 4556
rect 35414 4516 35454 4556
rect 35496 4516 35536 4556
rect 19996 4348 20036 4388
rect 33484 4348 33524 4388
rect 43939 4348 43979 4388
rect 44611 4348 44651 4388
rect 24028 4264 24068 4304
rect 25612 4264 25652 4304
rect 27100 4264 27140 4304
rect 31468 4264 31508 4304
rect 33964 4264 34004 4304
rect 41980 4264 42020 4304
rect 42748 4264 42788 4304
rect 45148 4264 45188 4304
rect 9676 4180 9716 4220
rect 9785 4180 9825 4220
rect 10060 4180 10100 4220
rect 18028 4180 18068 4220
rect 19276 4171 19316 4211
rect 21676 4171 21716 4211
rect 22924 4180 22964 4220
rect 24172 4180 24212 4220
rect 25420 4171 25460 4211
rect 25900 4180 25940 4220
rect 26155 4180 26195 4220
rect 26277 4180 26317 4220
rect 30028 4180 30068 4220
rect 31276 4171 31316 4211
rect 31747 4180 31787 4220
rect 31852 4180 31892 4220
rect 32236 4180 32276 4220
rect 32812 4171 32852 4211
rect 33292 4171 33332 4211
rect 34073 4180 34113 4220
rect 34348 4180 34388 4220
rect 17644 4096 17684 4136
rect 17884 4096 17924 4136
rect 19708 4096 19748 4136
rect 20332 4096 20372 4136
rect 21100 4096 21140 4136
rect 21340 4096 21380 4136
rect 23788 4096 23828 4136
rect 26764 4096 26804 4136
rect 27340 4096 27380 4136
rect 32332 4096 32372 4136
rect 38380 4096 38420 4136
rect 38572 4096 38612 4136
rect 42220 4096 42260 4136
rect 42604 4096 42644 4136
rect 42988 4096 43028 4136
rect 43372 4096 43412 4136
rect 43756 4096 43796 4136
rect 44236 4096 44276 4136
rect 44620 4096 44660 4136
rect 44908 4096 44948 4136
rect 26572 4012 26612 4052
rect 44476 4012 44516 4052
rect 9388 3928 9428 3968
rect 19468 3928 19508 3968
rect 20092 3928 20132 3968
rect 21484 3928 21524 3968
rect 27004 3928 27044 3968
rect 33676 3928 33716 3968
rect 38812 3928 38852 3968
rect 42364 3928 42404 3968
rect 43132 3928 43172 3968
rect 43516 3928 43556 3968
rect 3688 3760 3728 3800
rect 3770 3760 3810 3800
rect 3852 3760 3892 3800
rect 3934 3760 3974 3800
rect 4016 3760 4056 3800
rect 18808 3760 18848 3800
rect 18890 3760 18930 3800
rect 18972 3760 19012 3800
rect 19054 3760 19094 3800
rect 19136 3760 19176 3800
rect 33928 3760 33968 3800
rect 34010 3760 34050 3800
rect 34092 3760 34132 3800
rect 34174 3760 34214 3800
rect 34256 3760 34296 3800
rect 9244 3592 9284 3632
rect 9628 3592 9668 3632
rect 11212 3592 11252 3632
rect 12028 3592 12068 3632
rect 13612 3592 13652 3632
rect 18172 3592 18212 3632
rect 32572 3592 32612 3632
rect 42748 3592 42788 3632
rect 43900 3592 43940 3632
rect 45148 3592 45188 3632
rect 17788 3508 17828 3548
rect 21100 3508 21140 3548
rect 26860 3508 26900 3548
rect 27868 3508 27908 3548
rect 29452 3508 29492 3548
rect 32956 3508 32996 3548
rect 42268 3508 42308 3548
rect 43132 3508 43172 3548
rect 9004 3424 9044 3464
rect 9388 3424 9428 3464
rect 11788 3424 11828 3464
rect 15436 3424 15476 3464
rect 15772 3424 15812 3464
rect 16012 3424 16052 3464
rect 18028 3424 18068 3464
rect 18412 3424 18452 3464
rect 18796 3424 18836 3464
rect 19564 3424 19604 3464
rect 27004 3424 27044 3464
rect 27244 3424 27284 3464
rect 27628 3424 27668 3464
rect 30220 3424 30260 3464
rect 31180 3424 31220 3464
rect 32812 3424 32852 3464
rect 33196 3424 33236 3464
rect 33580 3424 33620 3464
rect 37516 3424 37556 3464
rect 37804 3424 37844 3464
rect 38188 3424 38228 3464
rect 38572 3424 38612 3464
rect 39052 3424 39092 3464
rect 39340 3424 39380 3464
rect 39724 3424 39764 3464
rect 42508 3424 42548 3464
rect 42988 3424 43028 3464
rect 43372 3424 43412 3464
rect 43756 3424 43796 3464
rect 44140 3424 44180 3464
rect 44524 3424 44564 3464
rect 44908 3424 44948 3464
rect 9772 3340 9812 3380
rect 11020 3340 11060 3380
rect 12172 3340 12212 3380
rect 13420 3340 13460 3380
rect 13804 3340 13844 3380
rect 15052 3340 15092 3380
rect 16204 3340 16244 3380
rect 17452 3340 17492 3380
rect 19075 3340 19115 3380
rect 19177 3340 19217 3380
rect 19660 3340 19700 3380
rect 20140 3340 20180 3380
rect 20628 3340 20668 3380
rect 21484 3331 21524 3371
rect 21772 3340 21812 3380
rect 24268 3340 24308 3380
rect 25516 3340 25556 3380
rect 26188 3340 26228 3380
rect 26443 3340 26483 3380
rect 26564 3340 26604 3380
rect 28012 3340 28052 3380
rect 29260 3340 29300 3380
rect 30691 3340 30731 3380
rect 30796 3340 30836 3380
rect 31276 3340 31316 3380
rect 31756 3340 31796 3380
rect 32275 3340 32315 3380
rect 32467 3340 32507 3380
rect 15676 3256 15716 3296
rect 21388 3256 21428 3296
rect 25708 3256 25748 3296
rect 33340 3256 33380 3296
rect 38428 3256 38468 3296
rect 39580 3256 39620 3296
rect 43516 3256 43556 3296
rect 44764 3256 44804 3296
rect 15244 3172 15284 3212
rect 17644 3172 17684 3212
rect 18556 3172 18596 3212
rect 20812 3172 20852 3212
rect 30460 3172 30500 3212
rect 37027 3172 37067 3212
rect 37315 3172 37355 3212
rect 37603 3172 37643 3212
rect 38044 3172 38084 3212
rect 39043 3172 39083 3212
rect 39964 3172 40004 3212
rect 4928 3004 4968 3044
rect 5010 3004 5050 3044
rect 5092 3004 5132 3044
rect 5174 3004 5214 3044
rect 5256 3004 5296 3044
rect 20048 3004 20088 3044
rect 20130 3004 20170 3044
rect 20212 3004 20252 3044
rect 20294 3004 20334 3044
rect 20376 3004 20416 3044
rect 35168 3004 35208 3044
rect 35250 3004 35290 3044
rect 35332 3004 35372 3044
rect 35414 3004 35454 3044
rect 35496 3004 35536 3044
rect 9196 2836 9236 2876
rect 10924 2836 10964 2876
rect 14044 2836 14084 2876
rect 20188 2836 20228 2876
rect 24508 2836 24548 2876
rect 45148 2836 45188 2876
rect 15916 2752 15956 2792
rect 31804 2752 31844 2792
rect 37516 2752 37556 2792
rect 37804 2752 37844 2792
rect 38092 2752 38132 2792
rect 38380 2752 38420 2792
rect 38668 2752 38708 2792
rect 7756 2668 7796 2708
rect 9004 2659 9044 2699
rect 9484 2668 9524 2708
rect 10732 2659 10772 2699
rect 15532 2668 15572 2708
rect 15811 2668 15851 2708
rect 18211 2668 18251 2708
rect 18316 2668 18356 2708
rect 18700 2668 18740 2708
rect 19276 2659 19316 2699
rect 19756 2659 19796 2699
rect 19987 2668 20027 2708
rect 7372 2584 7412 2624
rect 13804 2584 13844 2624
rect 18796 2584 18836 2624
rect 20428 2584 20468 2624
rect 24268 2584 24308 2624
rect 31276 2584 31316 2624
rect 31660 2584 31700 2624
rect 32044 2584 32084 2624
rect 36364 2584 36404 2624
rect 39244 2584 39284 2624
rect 39532 2584 39572 2624
rect 39724 2584 39764 2624
rect 40108 2584 40148 2624
rect 40492 2584 40532 2624
rect 40876 2584 40916 2624
rect 41164 2584 41204 2624
rect 43084 2584 43124 2624
rect 44140 2584 44180 2624
rect 44380 2584 44420 2624
rect 44524 2584 44564 2624
rect 44908 2584 44948 2624
rect 39964 2500 40004 2540
rect 44764 2500 44804 2540
rect 7612 2416 7652 2456
rect 16204 2416 16244 2456
rect 31036 2416 31076 2456
rect 31420 2416 31460 2456
rect 36604 2416 36644 2456
rect 40348 2416 40388 2456
rect 40732 2416 40772 2456
rect 42844 2416 42884 2456
rect 3688 2248 3728 2288
rect 3770 2248 3810 2288
rect 3852 2248 3892 2288
rect 3934 2248 3974 2288
rect 4016 2248 4056 2288
rect 18808 2248 18848 2288
rect 18890 2248 18930 2288
rect 18972 2248 19012 2288
rect 19054 2248 19094 2288
rect 19136 2248 19176 2288
rect 33928 2248 33968 2288
rect 34010 2248 34050 2288
rect 34092 2248 34132 2288
rect 34174 2248 34214 2288
rect 34256 2248 34296 2288
rect 4252 2080 4292 2120
rect 9628 2080 9668 2120
rect 45148 2080 45188 2120
rect 2716 1996 2756 2036
rect 43228 1996 43268 2036
rect 2476 1912 2516 1952
rect 4012 1912 4052 1952
rect 5740 1912 5780 1952
rect 7276 1912 7316 1952
rect 8812 1912 8852 1952
rect 9388 1912 9428 1952
rect 10348 1912 10388 1952
rect 11884 1912 11924 1952
rect 18796 1912 18836 1952
rect 39244 1912 39284 1952
rect 40108 1912 40148 1952
rect 42988 1912 43028 1952
rect 43372 1912 43412 1952
rect 43756 1912 43796 1952
rect 44140 1912 44180 1952
rect 44524 1912 44564 1952
rect 44908 1912 44948 1952
rect 40300 1828 40340 1868
rect 43996 1744 44036 1784
rect 5500 1660 5540 1700
rect 7036 1660 7076 1700
rect 8572 1660 8612 1700
rect 10108 1660 10148 1700
rect 11644 1660 11684 1700
rect 18556 1660 18596 1700
rect 39148 1660 39188 1700
rect 39427 1660 39467 1700
rect 39715 1660 39755 1700
rect 40579 1660 40619 1700
rect 43612 1660 43652 1700
rect 44380 1660 44420 1700
rect 44764 1660 44804 1700
rect 4928 1492 4968 1532
rect 5010 1492 5050 1532
rect 5092 1492 5132 1532
rect 5174 1492 5214 1532
rect 5256 1492 5296 1532
rect 20048 1492 20088 1532
rect 20130 1492 20170 1532
rect 20212 1492 20252 1532
rect 20294 1492 20334 1532
rect 20376 1492 20416 1532
rect 35168 1492 35208 1532
rect 35250 1492 35290 1532
rect 35332 1492 35372 1532
rect 35414 1492 35454 1532
rect 35496 1492 35536 1532
<< metal2 >>
rect 2467 11740 2476 11780
rect 2516 11740 26764 11780
rect 26804 11740 26813 11780
rect 2947 11656 2956 11696
rect 2996 11656 26956 11696
rect 26996 11656 27005 11696
rect 0 11024 90 11044
rect 46278 11024 46368 11044
rect 0 10984 1324 11024
rect 1364 10984 1373 11024
rect 43171 10984 43180 11024
rect 43220 10984 46368 11024
rect 0 10964 90 10984
rect 46278 10964 46368 10984
rect 0 10688 90 10708
rect 46278 10688 46368 10708
rect 0 10648 1132 10688
rect 1172 10648 1181 10688
rect 44035 10648 44044 10688
rect 44084 10648 46368 10688
rect 0 10628 90 10648
rect 46278 10628 46368 10648
rect 0 10352 90 10372
rect 46278 10352 46368 10372
rect 0 10312 1420 10352
rect 1460 10312 1469 10352
rect 44419 10312 44428 10352
rect 44468 10312 46368 10352
rect 0 10292 90 10312
rect 46278 10292 46368 10312
rect 19555 10228 19564 10268
rect 19604 10228 27244 10268
rect 27284 10228 27293 10268
rect 22828 10144 23156 10184
rect 22828 10100 22868 10144
rect 23116 10100 23156 10144
rect 24460 10144 26036 10184
rect 18595 10060 18604 10100
rect 18644 10060 19028 10100
rect 19171 10060 19180 10100
rect 19220 10060 22868 10100
rect 22924 10060 23060 10100
rect 23116 10060 24172 10100
rect 24212 10060 24221 10100
rect 0 10016 90 10036
rect 18988 10016 19028 10060
rect 22924 10016 22964 10060
rect 0 9976 980 10016
rect 1315 9976 1324 10016
rect 1364 9976 3148 10016
rect 3188 9976 3197 10016
rect 9763 9976 9772 10016
rect 9812 9976 15532 10016
rect 15572 9976 15581 10016
rect 18403 9976 18412 10016
rect 18452 9976 18892 10016
rect 18932 9976 18941 10016
rect 18988 9976 19892 10016
rect 20131 9976 20140 10016
rect 20180 9976 22964 10016
rect 23020 10016 23060 10060
rect 24460 10016 24500 10144
rect 25996 10100 26036 10144
rect 25027 10060 25036 10100
rect 25076 10060 25900 10100
rect 25940 10060 25949 10100
rect 25996 10060 28204 10100
rect 28244 10060 28253 10100
rect 29827 10060 29836 10100
rect 29876 10060 42988 10100
rect 43028 10060 43037 10100
rect 46278 10016 46368 10036
rect 23020 9976 24500 10016
rect 24547 9976 24556 10016
rect 24596 9976 42892 10016
rect 42932 9976 42941 10016
rect 44515 9976 44524 10016
rect 44564 9976 46368 10016
rect 0 9956 90 9976
rect 940 9848 980 9976
rect 19852 9932 19892 9976
rect 46278 9956 46368 9976
rect 7843 9892 7852 9932
rect 7892 9892 10060 9932
rect 10100 9892 10109 9932
rect 13411 9892 13420 9932
rect 13460 9892 16108 9932
rect 16148 9892 16157 9932
rect 16291 9892 16300 9932
rect 16340 9892 19564 9932
rect 19604 9892 19613 9932
rect 19852 9892 42316 9932
rect 42356 9892 42365 9932
rect 940 9808 2132 9848
rect 3679 9808 3688 9848
rect 3728 9808 3770 9848
rect 3810 9808 3852 9848
rect 3892 9808 3934 9848
rect 3974 9808 4016 9848
rect 4056 9808 4065 9848
rect 18799 9808 18808 9848
rect 18848 9808 18890 9848
rect 18930 9808 18972 9848
rect 19012 9808 19054 9848
rect 19094 9808 19136 9848
rect 19176 9808 19185 9848
rect 19948 9808 23252 9848
rect 27235 9808 27244 9848
rect 27284 9808 28972 9848
rect 29012 9808 29021 9848
rect 29251 9808 29260 9848
rect 29300 9808 30356 9848
rect 33919 9808 33928 9848
rect 33968 9808 34010 9848
rect 34050 9808 34092 9848
rect 34132 9808 34174 9848
rect 34214 9808 34256 9848
rect 34296 9808 34305 9848
rect 40483 9808 40492 9848
rect 40532 9808 44140 9848
rect 44180 9808 44189 9848
rect 0 9680 90 9700
rect 0 9640 2036 9680
rect 0 9620 90 9640
rect 1411 9556 1420 9596
rect 1460 9556 1748 9596
rect 1097 9472 1228 9512
rect 1268 9472 1277 9512
rect 1603 9472 1612 9512
rect 1652 9472 1661 9512
rect 0 9344 90 9364
rect 1612 9344 1652 9472
rect 1708 9428 1748 9556
rect 1996 9512 2036 9640
rect 2092 9512 2132 9808
rect 2860 9724 16300 9764
rect 16340 9724 16349 9764
rect 18403 9724 18412 9764
rect 18452 9724 18644 9764
rect 2860 9680 2900 9724
rect 18604 9680 18644 9724
rect 2227 9640 2236 9680
rect 2276 9640 2900 9680
rect 10195 9640 10204 9680
rect 10244 9640 11212 9680
rect 11252 9640 11261 9680
rect 11347 9640 11356 9680
rect 11396 9640 11980 9680
rect 12020 9640 12029 9680
rect 12115 9640 12124 9680
rect 12164 9640 12748 9680
rect 12788 9640 12797 9680
rect 12883 9640 12892 9680
rect 12932 9640 13172 9680
rect 13267 9640 13276 9680
rect 13316 9640 13900 9680
rect 13940 9640 13949 9680
rect 14035 9640 14044 9680
rect 14084 9640 14668 9680
rect 14708 9640 14717 9680
rect 14803 9640 14812 9680
rect 14852 9640 15052 9680
rect 15092 9640 15101 9680
rect 15187 9640 15196 9680
rect 15236 9640 15436 9680
rect 15476 9640 15485 9680
rect 15571 9640 15580 9680
rect 15620 9640 15820 9680
rect 15860 9640 15869 9680
rect 15955 9640 15964 9680
rect 16004 9640 16204 9680
rect 16244 9640 16253 9680
rect 16339 9640 16348 9680
rect 16388 9640 16588 9680
rect 16628 9640 16637 9680
rect 16723 9640 16732 9680
rect 16772 9640 16972 9680
rect 17012 9640 17021 9680
rect 17107 9640 17116 9680
rect 17156 9640 17356 9680
rect 17396 9640 17405 9680
rect 17491 9640 17500 9680
rect 17540 9640 17740 9680
rect 17780 9640 17789 9680
rect 17875 9640 17884 9680
rect 17924 9640 18124 9680
rect 18164 9640 18173 9680
rect 18259 9640 18268 9680
rect 18308 9640 18508 9680
rect 18548 9640 18557 9680
rect 18604 9640 18652 9680
rect 18692 9640 18701 9680
rect 19673 9640 19756 9680
rect 19796 9640 19804 9680
rect 19844 9640 19853 9680
rect 13132 9596 13172 9640
rect 10579 9556 10588 9596
rect 10628 9556 11404 9596
rect 11444 9556 11453 9596
rect 11731 9556 11740 9596
rect 11780 9556 12364 9596
rect 12404 9556 12413 9596
rect 12499 9556 12508 9596
rect 12548 9556 12940 9596
rect 12980 9556 12989 9596
rect 13132 9556 13516 9596
rect 13556 9556 13565 9596
rect 13651 9556 13660 9596
rect 13700 9556 14284 9596
rect 14324 9556 14333 9596
rect 14419 9556 14428 9596
rect 14468 9556 14860 9596
rect 14900 9556 14909 9596
rect 19027 9556 19036 9596
rect 19076 9556 19372 9596
rect 19412 9556 19421 9596
rect 19948 9512 19988 9808
rect 23212 9764 23252 9808
rect 23212 9724 26092 9764
rect 26132 9724 26141 9764
rect 26371 9724 26380 9764
rect 26420 9724 26956 9764
rect 26996 9724 27005 9764
rect 28867 9724 28876 9764
rect 28916 9724 29972 9764
rect 20179 9640 20188 9680
rect 20228 9640 20428 9680
rect 20468 9640 20477 9680
rect 20563 9640 20572 9680
rect 20612 9640 20812 9680
rect 20852 9640 20861 9680
rect 21331 9640 21340 9680
rect 21380 9640 24364 9680
rect 24404 9640 24413 9680
rect 24643 9640 24652 9680
rect 24692 9640 25172 9680
rect 25315 9640 25324 9680
rect 25364 9640 25852 9680
rect 25892 9640 25901 9680
rect 26179 9640 26188 9680
rect 26228 9640 27092 9680
rect 27305 9640 27388 9680
rect 27428 9640 27436 9680
rect 27476 9640 27485 9680
rect 28483 9640 28492 9680
rect 28532 9640 28724 9680
rect 20908 9556 21196 9596
rect 21236 9556 21245 9596
rect 21571 9556 21580 9596
rect 21620 9556 21629 9596
rect 21676 9556 21964 9596
rect 22004 9556 22013 9596
rect 22147 9556 22156 9596
rect 22196 9556 22205 9596
rect 23212 9556 23692 9596
rect 23732 9556 23741 9596
rect 24259 9556 24268 9596
rect 24308 9556 24317 9596
rect 24451 9556 24460 9596
rect 24500 9556 24788 9596
rect 20908 9512 20948 9556
rect 21580 9512 21620 9556
rect 21676 9512 21716 9556
rect 22156 9512 22196 9556
rect 23212 9512 23252 9556
rect 24268 9512 24308 9556
rect 24748 9512 24788 9556
rect 25132 9512 25172 9640
rect 25411 9556 25420 9596
rect 25460 9556 26324 9596
rect 26284 9512 26324 9556
rect 27052 9512 27092 9640
rect 28291 9556 28300 9596
rect 28340 9556 28628 9596
rect 28588 9512 28628 9556
rect 28684 9512 28724 9640
rect 28819 9556 28828 9596
rect 28868 9556 29876 9596
rect 1987 9472 1996 9512
rect 2036 9472 2045 9512
rect 2092 9472 2380 9512
rect 2420 9472 2429 9512
rect 2755 9472 2764 9512
rect 2804 9472 2813 9512
rect 3017 9472 3148 9512
rect 3188 9472 3197 9512
rect 9955 9472 9964 9512
rect 10004 9472 10013 9512
rect 10339 9472 10348 9512
rect 10388 9472 10397 9512
rect 10601 9472 10732 9512
rect 10772 9472 10781 9512
rect 10985 9472 11116 9512
rect 11156 9472 11165 9512
rect 11369 9472 11500 9512
rect 11540 9472 11549 9512
rect 11753 9472 11884 9512
rect 11924 9472 11933 9512
rect 12259 9472 12268 9512
rect 12308 9472 12460 9512
rect 12500 9472 12509 9512
rect 12643 9472 12652 9512
rect 12692 9472 12823 9512
rect 13027 9472 13036 9512
rect 13076 9472 13085 9512
rect 13411 9472 13420 9512
rect 13460 9472 13612 9512
rect 13652 9472 13661 9512
rect 13795 9472 13804 9512
rect 13844 9472 13996 9512
rect 14036 9472 14045 9512
rect 14179 9472 14188 9512
rect 14228 9472 14359 9512
rect 14441 9472 14572 9512
rect 14612 9472 14621 9512
rect 14825 9472 14956 9512
rect 14996 9472 15005 9512
rect 15209 9472 15340 9512
rect 15380 9472 15389 9512
rect 15715 9472 15724 9512
rect 15764 9472 15773 9512
rect 16099 9472 16108 9512
rect 16148 9472 16204 9512
rect 16244 9472 16279 9512
rect 16361 9472 16492 9512
rect 16532 9472 16541 9512
rect 16745 9472 16876 9512
rect 16916 9472 16925 9512
rect 17129 9472 17260 9512
rect 17300 9472 17309 9512
rect 17513 9472 17644 9512
rect 17684 9472 17693 9512
rect 17897 9472 18028 9512
rect 18068 9472 18077 9512
rect 18281 9472 18412 9512
rect 18452 9472 18461 9512
rect 18595 9472 18604 9512
rect 18644 9472 18796 9512
rect 18836 9472 18845 9512
rect 19049 9472 19084 9512
rect 19124 9472 19180 9512
rect 19220 9472 19229 9512
rect 19594 9472 19603 9512
rect 19643 9472 19700 9512
rect 19939 9472 19948 9512
rect 19988 9472 19997 9512
rect 20131 9472 20140 9512
rect 20180 9472 20332 9512
rect 20372 9472 20381 9512
rect 20899 9472 20908 9512
rect 20948 9472 20957 9512
rect 21091 9472 21100 9512
rect 21140 9472 21620 9512
rect 21667 9472 21676 9512
rect 21716 9472 21725 9512
rect 21859 9472 21868 9512
rect 21908 9472 22196 9512
rect 22243 9472 22252 9512
rect 22292 9472 22348 9512
rect 22388 9472 22423 9512
rect 22531 9472 22540 9512
rect 22580 9472 22828 9512
rect 22868 9472 22877 9512
rect 23203 9472 23212 9512
rect 23252 9472 23261 9512
rect 23587 9472 23596 9512
rect 23636 9472 23884 9512
rect 23924 9472 23933 9512
rect 24041 9472 24076 9512
rect 24116 9472 24172 9512
rect 24212 9472 24221 9512
rect 24268 9472 24556 9512
rect 24596 9472 24605 9512
rect 24739 9472 24748 9512
rect 24788 9472 24797 9512
rect 25123 9472 25132 9512
rect 25172 9472 25181 9512
rect 25699 9472 25708 9512
rect 25748 9472 25757 9512
rect 25891 9472 25900 9512
rect 25940 9472 26092 9512
rect 26132 9472 26141 9512
rect 26275 9472 26284 9512
rect 26324 9472 26333 9512
rect 26851 9472 26860 9512
rect 26900 9472 26909 9512
rect 27043 9472 27052 9512
rect 27092 9472 27101 9512
rect 27148 9472 27628 9512
rect 27668 9472 27677 9512
rect 28099 9472 28108 9512
rect 28148 9472 28396 9512
rect 28436 9472 28445 9512
rect 28579 9472 28588 9512
rect 28628 9472 28637 9512
rect 28684 9472 29164 9512
rect 29204 9472 29213 9512
rect 29539 9472 29548 9512
rect 29588 9472 29597 9512
rect 2764 9428 2804 9472
rect 1708 9388 2804 9428
rect 2860 9388 7892 9428
rect 2860 9344 2900 9388
rect 0 9304 1652 9344
rect 2611 9304 2620 9344
rect 2660 9304 2900 9344
rect 2995 9304 3004 9344
rect 3044 9304 6124 9344
rect 6164 9304 6173 9344
rect 0 9284 90 9304
rect 7852 9260 7892 9388
rect 9964 9344 10004 9472
rect 10348 9428 10388 9472
rect 10348 9388 12844 9428
rect 12884 9388 12893 9428
rect 13036 9344 13076 9472
rect 15724 9428 15764 9472
rect 19660 9428 19700 9472
rect 25708 9428 25748 9472
rect 26860 9428 26900 9472
rect 27148 9428 27188 9472
rect 29548 9428 29588 9472
rect 15724 9388 17836 9428
rect 17876 9388 17885 9428
rect 19660 9388 19756 9428
rect 19796 9388 19805 9428
rect 19939 9388 19948 9428
rect 19988 9388 19997 9428
rect 22348 9388 24556 9428
rect 24596 9388 24605 9428
rect 24835 9388 24844 9428
rect 24884 9388 25748 9428
rect 25795 9388 25804 9428
rect 25844 9388 26900 9428
rect 26947 9388 26956 9428
rect 26996 9388 27188 9428
rect 27331 9388 27340 9428
rect 27380 9388 27476 9428
rect 28675 9388 28684 9428
rect 28724 9388 29588 9428
rect 29836 9428 29876 9556
rect 29932 9512 29972 9724
rect 30316 9512 30356 9808
rect 32620 9724 40340 9764
rect 41827 9724 41836 9764
rect 41876 9724 43796 9764
rect 31171 9640 31180 9680
rect 31220 9640 31228 9680
rect 31268 9640 31351 9680
rect 31555 9640 31564 9680
rect 31604 9640 31996 9680
rect 32036 9640 32045 9680
rect 31363 9556 31372 9596
rect 31412 9556 31612 9596
rect 31652 9556 31661 9596
rect 31747 9556 31756 9596
rect 31796 9556 32380 9596
rect 32420 9556 32429 9596
rect 32620 9512 32660 9724
rect 33475 9640 33484 9680
rect 33524 9640 34300 9680
rect 34340 9640 34349 9680
rect 34601 9640 34684 9680
rect 34724 9640 34732 9680
rect 34772 9640 34781 9680
rect 35011 9640 35020 9680
rect 35060 9640 35836 9680
rect 35876 9640 35885 9680
rect 32707 9556 32716 9596
rect 32756 9556 33532 9596
rect 33572 9556 33581 9596
rect 35395 9556 35404 9596
rect 35444 9556 35452 9596
rect 35492 9556 35575 9596
rect 40300 9512 40340 9724
rect 42835 9640 42844 9680
rect 42884 9640 43084 9680
rect 43124 9640 43133 9680
rect 43756 9596 43796 9724
rect 46278 9680 46368 9700
rect 43913 9640 43996 9680
rect 44036 9640 44044 9680
rect 44084 9640 44093 9680
rect 44297 9640 44380 9680
rect 44420 9640 44428 9680
rect 44468 9640 44477 9680
rect 44755 9640 44764 9680
rect 44804 9640 46368 9680
rect 46278 9620 46368 9640
rect 40387 9556 40396 9596
rect 40436 9556 43124 9596
rect 43084 9512 43124 9556
rect 43180 9556 43564 9596
rect 43604 9556 43613 9596
rect 43756 9556 43892 9596
rect 29923 9472 29932 9512
rect 29972 9472 29981 9512
rect 30307 9472 30316 9512
rect 30356 9472 30365 9512
rect 31337 9472 31468 9512
rect 31508 9472 31517 9512
rect 31651 9472 31660 9512
rect 31700 9472 31852 9512
rect 31892 9472 31901 9512
rect 32105 9472 32236 9512
rect 32276 9472 32285 9512
rect 32611 9472 32620 9512
rect 32660 9472 32669 9512
rect 32969 9472 33004 9512
rect 33044 9472 33100 9512
rect 33140 9472 33149 9512
rect 33257 9472 33388 9512
rect 33428 9472 33437 9512
rect 33641 9472 33772 9512
rect 33812 9472 33821 9512
rect 34025 9472 34156 9512
rect 34196 9472 34205 9512
rect 34531 9472 34540 9512
rect 34580 9472 34732 9512
rect 34772 9472 34781 9512
rect 34915 9472 34924 9512
rect 34964 9472 35020 9512
rect 35060 9472 35095 9512
rect 35212 9472 35308 9512
rect 35348 9472 35357 9512
rect 35561 9472 35692 9512
rect 35732 9472 35741 9512
rect 36067 9472 36076 9512
rect 36116 9472 38860 9512
rect 38900 9472 38909 9512
rect 40300 9472 41644 9512
rect 41684 9472 41693 9512
rect 42089 9472 42220 9512
rect 42260 9472 42269 9512
rect 42473 9472 42604 9512
rect 42644 9472 42653 9512
rect 43075 9472 43084 9512
rect 43124 9472 43133 9512
rect 29836 9388 31412 9428
rect 19948 9344 19988 9388
rect 22348 9344 22388 9388
rect 27436 9344 27476 9388
rect 9964 9304 10828 9344
rect 10868 9304 10877 9344
rect 10963 9304 10972 9344
rect 11012 9304 11788 9344
rect 11828 9304 11837 9344
rect 13036 9304 13364 9344
rect 19289 9304 19372 9344
rect 19412 9304 19420 9344
rect 19460 9304 19469 9344
rect 19555 9304 19564 9344
rect 19604 9304 19988 9344
rect 20044 9304 22388 9344
rect 22483 9304 22492 9344
rect 22532 9304 23308 9344
rect 23348 9304 23357 9344
rect 23443 9304 23452 9344
rect 23492 9304 23692 9344
rect 23732 9304 23741 9344
rect 23827 9304 23836 9344
rect 23876 9304 24884 9344
rect 24979 9304 24988 9344
rect 25028 9304 25036 9344
rect 25076 9304 25159 9344
rect 25363 9304 25372 9344
rect 25412 9304 25708 9344
rect 25748 9304 25757 9344
rect 26393 9304 26476 9344
rect 26516 9304 26524 9344
rect 26564 9304 26573 9344
rect 26851 9304 26860 9344
rect 26900 9304 27292 9344
rect 27332 9304 27341 9344
rect 27436 9304 30260 9344
rect 13324 9260 13364 9304
rect 20044 9260 20084 9304
rect 1459 9220 1468 9260
rect 1508 9220 1708 9260
rect 1748 9220 1757 9260
rect 1843 9220 1852 9260
rect 1892 9220 1901 9260
rect 3379 9220 3388 9260
rect 3428 9220 7084 9260
rect 7124 9220 7133 9260
rect 7852 9220 10924 9260
rect 10964 9220 10973 9260
rect 13324 9220 14284 9260
rect 14324 9220 14333 9260
rect 14659 9220 14668 9260
rect 14708 9220 17452 9260
rect 17492 9220 17501 9260
rect 19996 9220 20084 9260
rect 20659 9220 20668 9260
rect 20708 9220 20716 9260
rect 20756 9220 20839 9260
rect 21187 9220 21196 9260
rect 21236 9220 21436 9260
rect 21476 9220 21485 9260
rect 22099 9220 22108 9260
rect 22148 9220 22484 9260
rect 22531 9220 22540 9260
rect 22580 9220 22588 9260
rect 22628 9220 22711 9260
rect 23587 9220 23596 9260
rect 23636 9220 23932 9260
rect 23972 9220 23981 9260
rect 24307 9220 24316 9260
rect 24356 9220 24364 9260
rect 24404 9220 24487 9260
rect 1852 9176 1892 9220
rect 19996 9176 20036 9220
rect 1852 9136 15092 9176
rect 16195 9136 16204 9176
rect 16244 9136 19372 9176
rect 19412 9136 19421 9176
rect 19948 9136 20036 9176
rect 15052 9092 15092 9136
rect 19948 9092 19988 9136
rect 22444 9092 22484 9220
rect 24844 9176 24884 9304
rect 25123 9220 25132 9260
rect 25172 9220 25468 9260
rect 25508 9220 25517 9260
rect 26611 9220 26620 9260
rect 26660 9220 26956 9260
rect 26996 9220 27005 9260
rect 27139 9220 27148 9260
rect 27188 9220 28156 9260
rect 28196 9220 28205 9260
rect 28300 9220 28924 9260
rect 28964 9220 28973 9260
rect 29155 9220 29164 9260
rect 29204 9220 29308 9260
rect 29348 9220 29357 9260
rect 29452 9220 29692 9260
rect 29732 9220 29741 9260
rect 29827 9220 29836 9260
rect 29876 9220 30076 9260
rect 30116 9220 30125 9260
rect 28300 9176 28340 9220
rect 29452 9176 29492 9220
rect 24163 9136 24172 9176
rect 24212 9136 24788 9176
rect 24844 9136 26380 9176
rect 26420 9136 26429 9176
rect 26659 9136 26668 9176
rect 26708 9136 28340 9176
rect 28579 9136 28588 9176
rect 28628 9136 29492 9176
rect 24748 9092 24788 9136
rect 30220 9092 30260 9304
rect 31372 9260 31412 9388
rect 31939 9304 31948 9344
rect 31988 9304 32764 9344
rect 32804 9304 32813 9344
rect 33100 9304 33148 9344
rect 33188 9304 33197 9344
rect 33379 9304 33388 9344
rect 33428 9304 33772 9344
rect 33812 9304 33821 9344
rect 34531 9304 34540 9344
rect 34580 9304 35068 9344
rect 35108 9304 35117 9344
rect 33100 9260 33140 9304
rect 31372 9220 32044 9260
rect 32084 9220 32093 9260
rect 32323 9220 32332 9260
rect 32372 9220 33140 9260
rect 33187 9220 33196 9260
rect 33236 9220 33916 9260
rect 33956 9220 33965 9260
rect 35212 9176 35252 9472
rect 43180 9428 43220 9556
rect 43852 9512 43892 9556
rect 43459 9472 43468 9512
rect 43508 9472 43756 9512
rect 43796 9472 43805 9512
rect 43852 9472 44140 9512
rect 44180 9472 44189 9512
rect 44515 9472 44524 9512
rect 44564 9472 44573 9512
rect 44777 9472 44908 9512
rect 44948 9472 44957 9512
rect 37795 9388 37804 9428
rect 37844 9388 43220 9428
rect 44524 9344 44564 9472
rect 46278 9344 46368 9364
rect 37699 9304 37708 9344
rect 37748 9304 44564 9344
rect 45139 9304 45148 9344
rect 45188 9304 46368 9344
rect 46278 9284 46368 9304
rect 35779 9220 35788 9260
rect 35828 9220 40492 9260
rect 40532 9220 40541 9260
rect 41827 9220 41836 9260
rect 41876 9220 41923 9260
rect 41963 9220 42007 9260
rect 42451 9220 42460 9260
rect 42500 9220 42740 9260
rect 34531 9136 34540 9176
rect 34580 9136 35252 9176
rect 35971 9136 35980 9176
rect 36020 9136 37612 9176
rect 37652 9136 37661 9176
rect 37891 9136 37900 9176
rect 37940 9136 42220 9176
rect 42260 9136 42269 9176
rect 42700 9092 42740 9220
rect 43276 9220 43324 9260
rect 43364 9220 43373 9260
rect 43450 9220 43459 9260
rect 43508 9220 43639 9260
rect 43276 9176 43316 9220
rect 43276 9136 46196 9176
rect 4919 9052 4928 9092
rect 4968 9052 5010 9092
rect 5050 9052 5092 9092
rect 5132 9052 5174 9092
rect 5214 9052 5256 9092
rect 5296 9052 5305 9092
rect 10051 9052 10060 9092
rect 10100 9052 11884 9092
rect 11924 9052 11933 9092
rect 15052 9052 19796 9092
rect 0 9008 90 9028
rect 0 8968 1228 9008
rect 1268 8968 1277 9008
rect 12259 8968 12268 9008
rect 12308 8968 16684 9008
rect 16724 8968 16733 9008
rect 16867 8968 16876 9008
rect 16916 8968 19660 9008
rect 19700 8968 19709 9008
rect 0 8948 90 8968
rect 19756 8924 19796 9052
rect 19852 9052 19988 9092
rect 20039 9052 20048 9092
rect 20088 9052 20130 9092
rect 20170 9052 20212 9092
rect 20252 9052 20294 9092
rect 20334 9052 20376 9092
rect 20416 9052 20425 9092
rect 22444 9052 23116 9092
rect 23156 9052 23165 9092
rect 24748 9052 26764 9092
rect 26804 9052 26813 9092
rect 27043 9052 27052 9092
rect 27092 9052 30164 9092
rect 30220 9052 31892 9092
rect 35159 9052 35168 9092
rect 35208 9052 35250 9092
rect 35290 9052 35332 9092
rect 35372 9052 35414 9092
rect 35454 9052 35496 9092
rect 35536 9052 35545 9092
rect 35587 9052 35596 9092
rect 35636 9052 40108 9092
rect 40148 9052 40157 9092
rect 42700 9052 46100 9092
rect 19852 9008 19892 9052
rect 30124 9008 30164 9052
rect 31852 9008 31892 9052
rect 19843 8968 19852 9008
rect 19892 8968 19901 9008
rect 20803 8968 20812 9008
rect 20852 8968 28396 9008
rect 28436 8968 28445 9008
rect 28492 8968 29164 9008
rect 29204 8968 29213 9008
rect 30124 8968 31756 9008
rect 31796 8968 31805 9008
rect 31852 8968 42988 9008
rect 43028 8968 43037 9008
rect 28492 8924 28532 8968
rect 1459 8884 1468 8924
rect 1508 8884 7852 8924
rect 7892 8884 7901 8924
rect 9907 8884 9916 8924
rect 9956 8884 10540 8924
rect 10580 8884 10589 8924
rect 10675 8884 10684 8924
rect 10724 8884 11020 8924
rect 11060 8884 11069 8924
rect 11443 8884 11452 8924
rect 11492 8884 11596 8924
rect 11636 8884 11645 8924
rect 11801 8884 11884 8924
rect 11963 8884 11981 8924
rect 12163 8884 12172 8924
rect 12212 8884 12220 8924
rect 12260 8884 12343 8924
rect 12547 8884 12556 8924
rect 12596 8884 12604 8924
rect 12644 8884 12727 8924
rect 12979 8884 12988 8924
rect 13028 8884 13036 8924
rect 13076 8884 13159 8924
rect 13315 8884 13324 8924
rect 13364 8884 13372 8924
rect 13412 8884 13495 8924
rect 13699 8884 13708 8924
rect 13748 8884 13756 8924
rect 13796 8884 13879 8924
rect 14467 8884 14476 8924
rect 14516 8884 14524 8924
rect 14564 8884 14647 8924
rect 15235 8884 15244 8924
rect 15284 8884 15292 8924
rect 15332 8884 15415 8924
rect 15619 8884 15628 8924
rect 15668 8884 15676 8924
rect 15716 8884 15799 8924
rect 16003 8884 16012 8924
rect 16052 8884 16060 8924
rect 16100 8884 16183 8924
rect 16387 8884 16396 8924
rect 16436 8884 16444 8924
rect 16484 8884 16567 8924
rect 16771 8884 16780 8924
rect 16820 8884 16828 8924
rect 16868 8884 16951 8924
rect 17155 8884 17164 8924
rect 17204 8884 17212 8924
rect 17252 8884 17335 8924
rect 17539 8884 17548 8924
rect 17588 8884 17596 8924
rect 17636 8884 17719 8924
rect 17923 8884 17932 8924
rect 17972 8884 17980 8924
rect 18020 8884 18103 8924
rect 18307 8884 18316 8924
rect 18356 8884 18364 8924
rect 18404 8884 18487 8924
rect 18691 8884 18700 8924
rect 18740 8884 18748 8924
rect 18788 8884 18871 8924
rect 19123 8884 19132 8924
rect 19172 8884 19276 8924
rect 19316 8884 19325 8924
rect 19459 8884 19468 8924
rect 19508 8884 19516 8924
rect 19556 8884 19639 8924
rect 19756 8884 20044 8924
rect 20084 8884 20093 8924
rect 20275 8884 20284 8924
rect 20324 8884 20524 8924
rect 20564 8884 20573 8924
rect 20969 8884 21004 8924
rect 21044 8884 21100 8924
rect 21140 8884 21149 8924
rect 21283 8884 21292 8924
rect 21332 8884 28532 8924
rect 28675 8884 28684 8924
rect 28724 8884 31948 8924
rect 31988 8884 31997 8924
rect 32131 8884 32140 8924
rect 32180 8884 32188 8924
rect 32228 8884 32311 8924
rect 32515 8884 32524 8924
rect 32564 8884 32572 8924
rect 32612 8884 32695 8924
rect 32899 8884 32908 8924
rect 32948 8884 32956 8924
rect 32996 8884 33079 8924
rect 33283 8884 33292 8924
rect 33332 8884 33340 8924
rect 33380 8884 33463 8924
rect 33667 8884 33676 8924
rect 33716 8884 33724 8924
rect 33764 8884 33847 8924
rect 34099 8884 34108 8924
rect 34148 8884 34348 8924
rect 34388 8884 34397 8924
rect 34819 8884 34828 8924
rect 34868 8884 34876 8924
rect 34916 8884 34999 8924
rect 37219 8884 37228 8924
rect 37268 8884 37900 8924
rect 37940 8884 37949 8924
rect 38476 8884 43516 8924
rect 43556 8884 43565 8924
rect 44371 8884 44380 8924
rect 44420 8884 44524 8924
rect 44564 8884 44573 8924
rect 1123 8800 1132 8840
rect 1172 8800 2420 8840
rect 10291 8800 10300 8840
rect 10340 8800 10964 8840
rect 19747 8800 19756 8840
rect 19796 8800 20428 8840
rect 20468 8800 20477 8840
rect 20611 8800 20620 8840
rect 20660 8800 20668 8840
rect 20708 8800 20791 8840
rect 21715 8800 21724 8840
rect 21764 8800 22388 8840
rect 22819 8800 22828 8840
rect 22868 8800 23548 8840
rect 23588 8800 23597 8840
rect 23971 8800 23980 8840
rect 24020 8800 25660 8840
rect 25700 8800 25709 8840
rect 25891 8800 25900 8840
rect 25940 8800 28052 8840
rect 28195 8800 28204 8840
rect 28244 8800 28252 8840
rect 28292 8800 28375 8840
rect 29395 8800 29404 8840
rect 29444 8800 29740 8840
rect 29780 8800 29789 8840
rect 32611 8800 32620 8840
rect 32660 8800 34388 8840
rect 34435 8800 34444 8840
rect 34484 8800 34492 8840
rect 34532 8800 34615 8840
rect 34723 8800 34732 8840
rect 34772 8800 38380 8840
rect 38420 8800 38429 8840
rect 556 8716 2036 8756
rect 0 8672 90 8692
rect 556 8672 596 8716
rect 1996 8672 2036 8716
rect 2380 8672 2420 8800
rect 10924 8756 10964 8800
rect 9667 8716 9676 8756
rect 9716 8716 10484 8756
rect 10924 8716 11348 8756
rect 11465 8716 11596 8756
rect 11636 8716 11645 8756
rect 10444 8672 10484 8716
rect 0 8632 596 8672
rect 643 8632 652 8672
rect 692 8632 1228 8672
rect 1268 8632 1277 8672
rect 1603 8632 1612 8672
rect 1652 8632 1661 8672
rect 1721 8632 1804 8672
rect 1844 8632 1852 8672
rect 1892 8632 1901 8672
rect 1987 8632 1996 8672
rect 2036 8632 2045 8672
rect 2105 8632 2188 8672
rect 2228 8632 2236 8672
rect 2276 8632 2285 8672
rect 2371 8632 2380 8672
rect 2420 8632 2429 8672
rect 2611 8632 2620 8672
rect 2660 8632 9004 8672
rect 9044 8632 9053 8672
rect 9641 8632 9676 8672
rect 9716 8632 9772 8672
rect 9812 8632 9821 8672
rect 10051 8632 10060 8672
rect 10100 8632 10156 8672
rect 10196 8632 10231 8672
rect 10435 8632 10444 8672
rect 10484 8632 10493 8672
rect 10819 8632 10828 8672
rect 10868 8632 10877 8672
rect 11081 8632 11212 8672
rect 11252 8632 11261 8672
rect 0 8612 90 8632
rect 0 8336 90 8356
rect 1612 8336 1652 8632
rect 10828 8504 10868 8632
rect 11308 8588 11348 8716
rect 11692 8692 11724 8732
rect 11764 8692 11773 8732
rect 11971 8716 11980 8756
rect 12020 8716 12884 8756
rect 12931 8716 12940 8756
rect 12980 8716 13652 8756
rect 11692 8672 11732 8692
rect 12844 8672 12884 8716
rect 13612 8672 13652 8716
rect 18988 8716 19852 8756
rect 19892 8716 19901 8756
rect 20140 8716 21292 8756
rect 21332 8716 21341 8756
rect 18988 8672 19028 8716
rect 20140 8672 20180 8716
rect 22348 8672 22388 8800
rect 28012 8756 28052 8800
rect 25987 8716 25996 8756
rect 26036 8716 26045 8756
rect 26179 8716 26188 8756
rect 26228 8716 26237 8756
rect 26755 8716 26764 8756
rect 26804 8716 26813 8756
rect 27497 8716 27628 8756
rect 27668 8716 27677 8756
rect 27748 8716 27757 8756
rect 27797 8716 27956 8756
rect 28003 8716 28012 8756
rect 28052 8716 28061 8756
rect 28492 8716 29836 8756
rect 29876 8716 29885 8756
rect 32428 8716 33100 8756
rect 33140 8716 33149 8756
rect 33196 8716 33484 8756
rect 33524 8716 33533 8756
rect 33580 8716 34252 8756
rect 34292 8716 34301 8756
rect 25996 8672 26036 8716
rect 26188 8672 26228 8716
rect 26764 8672 26804 8716
rect 27916 8672 27956 8716
rect 28492 8672 28532 8716
rect 32428 8672 32468 8716
rect 33196 8672 33236 8716
rect 33580 8672 33620 8716
rect 34348 8672 34388 8800
rect 38476 8756 38516 8884
rect 46060 8840 46100 9052
rect 46156 8924 46196 9136
rect 46278 9008 46368 9028
rect 46252 8948 46368 9008
rect 46252 8924 46292 8948
rect 46156 8884 46292 8924
rect 38659 8800 38668 8840
rect 38708 8800 41932 8840
rect 41972 8800 41981 8840
rect 42307 8800 42316 8840
rect 42356 8800 42364 8840
rect 42404 8800 42487 8840
rect 42691 8800 42700 8840
rect 42740 8800 42748 8840
rect 42788 8800 42871 8840
rect 43075 8800 43084 8840
rect 43124 8800 43412 8840
rect 46060 8800 46196 8840
rect 34444 8716 38516 8756
rect 39043 8716 39052 8756
rect 39092 8716 40300 8756
rect 40340 8716 40349 8756
rect 42883 8716 42892 8756
rect 42932 8716 43124 8756
rect 11395 8632 11404 8672
rect 11444 8632 11732 8672
rect 11884 8632 12268 8672
rect 12308 8632 12317 8672
rect 12451 8632 12460 8672
rect 12500 8632 12509 8672
rect 12835 8632 12844 8672
rect 12884 8632 12893 8672
rect 13097 8632 13228 8672
rect 13268 8632 13277 8672
rect 13603 8632 13612 8672
rect 13652 8632 13661 8672
rect 13987 8632 13996 8672
rect 14036 8632 14188 8672
rect 14228 8632 14237 8672
rect 14371 8632 14380 8672
rect 14420 8632 14551 8672
rect 14633 8632 14764 8672
rect 14804 8632 14813 8672
rect 14860 8632 14956 8672
rect 14996 8632 15005 8672
rect 15113 8632 15196 8672
rect 15236 8632 15244 8672
rect 15284 8632 15293 8672
rect 15401 8632 15532 8672
rect 15572 8632 15581 8672
rect 15785 8632 15916 8672
rect 15956 8632 15965 8672
rect 16291 8632 16300 8672
rect 16340 8632 16349 8672
rect 16553 8632 16684 8672
rect 16724 8632 16733 8672
rect 17059 8632 17068 8672
rect 17108 8632 17396 8672
rect 17443 8632 17452 8672
rect 17492 8632 17548 8672
rect 17588 8632 17623 8672
rect 17705 8632 17740 8672
rect 17780 8632 17836 8672
rect 17876 8632 17885 8672
rect 18089 8632 18220 8672
rect 18260 8632 18269 8672
rect 18473 8632 18604 8672
rect 18644 8632 18653 8672
rect 18979 8632 18988 8672
rect 19028 8632 19037 8672
rect 19171 8632 19180 8672
rect 19220 8632 19372 8672
rect 19412 8632 19421 8672
rect 19625 8632 19756 8672
rect 19796 8632 19805 8672
rect 19891 8632 19900 8672
rect 19940 8632 19948 8672
rect 19988 8632 20071 8672
rect 20131 8632 20140 8672
rect 20180 8632 20189 8672
rect 20236 8632 20524 8672
rect 20564 8632 20573 8672
rect 20777 8632 20908 8672
rect 20948 8632 20957 8672
rect 21353 8632 21388 8672
rect 21428 8632 21484 8672
rect 21524 8632 21533 8672
rect 21763 8632 21772 8672
rect 21812 8632 22060 8672
rect 22100 8632 22109 8672
rect 22348 8632 23308 8672
rect 23348 8632 23357 8672
rect 23491 8632 23500 8672
rect 23540 8632 23788 8672
rect 23828 8632 23837 8672
rect 25193 8632 25228 8672
rect 25268 8632 25324 8672
rect 25364 8632 25373 8672
rect 25603 8632 25612 8672
rect 25652 8632 25900 8672
rect 25940 8632 25949 8672
rect 25996 8632 26092 8672
rect 26132 8632 26141 8672
rect 26188 8632 26428 8672
rect 26468 8632 26477 8672
rect 26537 8632 26668 8672
rect 26708 8632 26717 8672
rect 26764 8632 26812 8672
rect 26852 8632 26861 8672
rect 27043 8632 27052 8672
rect 27092 8632 27223 8672
rect 27916 8632 28012 8672
rect 28052 8632 28061 8672
rect 28483 8632 28492 8672
rect 28532 8632 28541 8672
rect 29033 8632 29068 8672
rect 29108 8632 29164 8672
rect 29204 8632 29213 8672
rect 29443 8632 29452 8672
rect 29492 8632 29740 8672
rect 29780 8632 29789 8672
rect 30307 8632 30316 8672
rect 30356 8632 31564 8672
rect 31604 8632 31613 8672
rect 32419 8632 32428 8672
rect 32468 8632 32477 8672
rect 32803 8632 32812 8672
rect 32852 8632 32861 8672
rect 33187 8632 33196 8672
rect 33236 8632 33245 8672
rect 33571 8632 33580 8672
rect 33620 8632 33629 8672
rect 33955 8632 33964 8672
rect 34004 8632 34292 8672
rect 34339 8632 34348 8672
rect 34388 8632 34397 8672
rect 11884 8588 11924 8632
rect 12460 8588 12500 8632
rect 14860 8588 14900 8632
rect 11011 8548 11020 8588
rect 11060 8548 11068 8588
rect 11108 8548 11191 8588
rect 11308 8548 11924 8588
rect 11971 8548 11980 8588
rect 12020 8548 12500 8588
rect 12547 8548 12556 8588
rect 12596 8548 14612 8588
rect 14851 8548 14860 8588
rect 14900 8548 14909 8588
rect 14572 8504 14612 8548
rect 16300 8504 16340 8632
rect 17356 8588 17396 8632
rect 20236 8588 20276 8632
rect 28492 8588 28532 8632
rect 32812 8588 32852 8632
rect 34252 8588 34292 8632
rect 34444 8588 34484 8716
rect 43084 8672 43124 8716
rect 43372 8672 43412 8800
rect 43555 8716 43564 8756
rect 43604 8716 44564 8756
rect 44524 8672 44564 8716
rect 46156 8672 46196 8800
rect 46278 8672 46368 8692
rect 34601 8632 34732 8672
rect 34772 8632 34781 8672
rect 34828 8632 35116 8672
rect 35156 8632 35165 8672
rect 35299 8632 35308 8672
rect 35348 8632 38956 8672
rect 38996 8632 39005 8672
rect 41731 8632 41740 8672
rect 41780 8632 42604 8672
rect 42644 8632 42653 8672
rect 42857 8632 42988 8672
rect 43028 8632 43037 8672
rect 43084 8632 43132 8672
rect 43172 8632 43181 8672
rect 43363 8632 43372 8672
rect 43412 8632 43421 8672
rect 43468 8632 43756 8672
rect 43796 8632 43805 8672
rect 44009 8632 44140 8672
rect 44180 8632 44189 8672
rect 44515 8632 44524 8672
rect 44564 8632 44573 8672
rect 44777 8632 44908 8672
rect 44948 8632 44957 8672
rect 46156 8632 46368 8672
rect 34828 8588 34868 8632
rect 43468 8588 43508 8632
rect 46278 8612 46368 8632
rect 17347 8548 17356 8588
rect 17396 8548 17405 8588
rect 20076 8548 20140 8588
rect 20180 8548 20276 8588
rect 21571 8548 21580 8588
rect 21620 8548 21820 8588
rect 21860 8548 21869 8588
rect 21964 8548 24940 8588
rect 24980 8548 24989 8588
rect 25555 8548 25564 8588
rect 25604 8548 25804 8588
rect 25844 8548 25853 8588
rect 26323 8548 26332 8588
rect 26372 8548 26764 8588
rect 26804 8548 26813 8588
rect 27427 8548 27436 8588
rect 27476 8548 28532 8588
rect 28588 8548 29684 8588
rect 32812 8548 33484 8588
rect 33524 8548 33533 8588
rect 34252 8548 34484 8588
rect 34540 8548 34868 8588
rect 34915 8548 34924 8588
rect 34964 8548 40780 8588
rect 40820 8548 40829 8588
rect 42883 8548 42892 8588
rect 42932 8548 43508 8588
rect 21964 8504 22004 8548
rect 28588 8504 28628 8548
rect 29644 8504 29684 8548
rect 34540 8504 34580 8548
rect 10339 8464 10348 8504
rect 10388 8464 12076 8504
rect 12116 8464 12125 8504
rect 13891 8464 13900 8504
rect 13940 8464 14140 8504
rect 14180 8464 14189 8504
rect 14572 8464 16340 8504
rect 18115 8464 18124 8504
rect 18164 8464 22004 8504
rect 22051 8464 22060 8504
rect 22100 8464 25228 8504
rect 25268 8464 25277 8504
rect 27209 8464 27340 8504
rect 27380 8464 27389 8504
rect 27523 8464 27532 8504
rect 27572 8464 28628 8504
rect 28867 8464 28876 8504
rect 28916 8464 29500 8504
rect 29540 8464 29549 8504
rect 29644 8464 33580 8504
rect 33620 8464 33629 8504
rect 33763 8464 33772 8504
rect 33812 8464 34580 8504
rect 35011 8464 35020 8504
rect 35060 8464 43220 8504
rect 44755 8464 44764 8504
rect 44804 8464 45044 8504
rect 45139 8464 45148 8504
rect 45188 8464 45772 8504
rect 45812 8464 45821 8504
rect 0 8296 1652 8336
rect 3532 8380 12364 8420
rect 12404 8380 12413 8420
rect 14563 8380 14572 8420
rect 14612 8380 42740 8420
rect 0 8276 90 8296
rect 3532 8252 3572 8380
rect 3679 8296 3688 8336
rect 3728 8296 3770 8336
rect 3810 8296 3852 8336
rect 3892 8296 3934 8336
rect 3974 8296 4016 8336
rect 4056 8296 4065 8336
rect 4387 8296 4396 8336
rect 4436 8296 11116 8336
rect 11156 8296 11165 8336
rect 11299 8296 11308 8336
rect 11348 8296 18508 8336
rect 18548 8296 18557 8336
rect 18799 8296 18808 8336
rect 18848 8296 18890 8336
rect 18930 8296 18972 8336
rect 19012 8296 19054 8336
rect 19094 8296 19136 8336
rect 19176 8296 19185 8336
rect 22435 8296 22444 8336
rect 22484 8296 22636 8336
rect 22676 8296 22685 8336
rect 27715 8296 27724 8336
rect 27764 8296 28780 8336
rect 28820 8296 28829 8336
rect 30019 8296 30028 8336
rect 30068 8296 33812 8336
rect 33919 8296 33928 8336
rect 33968 8296 34010 8336
rect 34050 8296 34092 8336
rect 34132 8296 34174 8336
rect 34214 8296 34256 8336
rect 34296 8296 34305 8336
rect 34627 8296 34636 8336
rect 34676 8296 35980 8336
rect 36020 8296 36029 8336
rect 38851 8296 38860 8336
rect 38900 8296 41972 8336
rect 33772 8252 33812 8296
rect 3148 8212 3572 8252
rect 7843 8212 7852 8252
rect 7892 8212 12844 8252
rect 12884 8212 12893 8252
rect 17443 8212 17452 8252
rect 17492 8212 18644 8252
rect 26083 8212 26092 8252
rect 26132 8212 33580 8252
rect 33620 8212 33629 8252
rect 33772 8212 40436 8252
rect 0 8000 90 8020
rect 0 7960 652 8000
rect 692 7960 701 8000
rect 1097 7960 1228 8000
rect 1268 7960 1277 8000
rect 1603 7960 1612 8000
rect 1652 7960 1661 8000
rect 2345 7960 2476 8000
rect 2516 7960 2525 8000
rect 2707 7960 2716 8000
rect 2756 7960 2804 8000
rect 2851 7960 2860 8000
rect 2900 7960 2956 8000
rect 2996 7960 3031 8000
rect 0 7940 90 7960
rect 1612 7832 1652 7960
rect 2764 7916 2804 7960
rect 3148 7916 3188 8212
rect 18604 8168 18644 8212
rect 4396 8128 12460 8168
rect 12500 8128 12509 8168
rect 15139 8128 15148 8168
rect 15188 8128 17108 8168
rect 17827 8128 17836 8168
rect 17876 8128 17884 8168
rect 17924 8128 18007 8168
rect 18604 8128 20140 8168
rect 20180 8128 20189 8168
rect 22793 8128 22876 8168
rect 22916 8128 22924 8168
rect 22964 8128 22973 8168
rect 28121 8128 28204 8168
rect 28244 8128 28252 8168
rect 28292 8128 28301 8168
rect 28387 8128 28396 8168
rect 28436 8128 28636 8168
rect 28676 8128 28685 8168
rect 28771 8128 28780 8168
rect 28820 8128 29012 8168
rect 32083 8128 32092 8168
rect 32132 8128 33772 8168
rect 33812 8128 33821 8168
rect 34409 8128 34492 8168
rect 34532 8128 34540 8168
rect 34580 8128 34589 8168
rect 34723 8128 34732 8168
rect 34772 8128 34972 8168
rect 35012 8128 35021 8168
rect 36691 8128 36700 8168
rect 36740 8128 38668 8168
rect 38708 8128 38717 8168
rect 3628 8044 4300 8084
rect 4340 8044 4349 8084
rect 3628 8000 3668 8044
rect 4396 8000 4436 8128
rect 17068 8084 17108 8128
rect 9868 8044 10444 8084
rect 10484 8044 10493 8084
rect 10732 8044 12884 8084
rect 14659 8044 14668 8084
rect 14708 8044 17012 8084
rect 17068 8044 22060 8084
rect 22100 8044 22109 8084
rect 24835 8044 24844 8084
rect 24884 8044 25900 8084
rect 25940 8044 25949 8084
rect 26860 8044 28916 8084
rect 9868 8000 9908 8044
rect 3235 7960 3244 8000
rect 3284 7960 3415 8000
rect 3475 7960 3484 8000
rect 3524 7960 3572 8000
rect 3619 7960 3628 8000
rect 3668 7960 3677 8000
rect 3881 7960 4012 8000
rect 4052 7960 4061 8000
rect 4387 7960 4396 8000
rect 4436 7960 4445 8000
rect 9763 7960 9772 8000
rect 9812 7960 9908 8000
rect 10147 7960 10156 8000
rect 10196 7960 10252 8000
rect 10292 7960 10540 8000
rect 10580 7960 10589 8000
rect 2764 7876 3188 7916
rect 3532 7916 3572 7960
rect 9868 7916 9908 7960
rect 3532 7876 7948 7916
rect 7988 7876 7997 7916
rect 9379 7876 9388 7916
rect 9428 7876 9763 7916
rect 9803 7876 9812 7916
rect 9859 7876 9868 7916
rect 9908 7876 9917 7916
rect 10217 7876 10348 7916
rect 10388 7876 10397 7916
rect 10732 7832 10772 8044
rect 11299 7960 11308 8000
rect 11348 7960 12788 8000
rect 844 7792 1652 7832
rect 1843 7792 1852 7832
rect 1892 7792 2956 7832
rect 2996 7792 3005 7832
rect 3091 7792 3100 7832
rect 3140 7792 10772 7832
rect 10828 7916 10868 7925
rect 12748 7916 12788 7960
rect 10915 7876 10924 7916
rect 10964 7876 11316 7916
rect 11356 7876 11365 7916
rect 11657 7876 11788 7916
rect 11828 7876 11837 7916
rect 11945 7876 12067 7916
rect 12116 7876 12125 7916
rect 12259 7876 12268 7916
rect 12308 7876 12604 7916
rect 12644 7876 12653 7916
rect 12739 7876 12748 7916
rect 12788 7876 12797 7916
rect 10828 7832 10868 7876
rect 12844 7832 12884 8044
rect 16972 8000 17012 8044
rect 26860 8000 26900 8044
rect 28876 8000 28916 8044
rect 14345 7960 14476 8000
rect 14516 7960 14525 8000
rect 16963 7960 16972 8000
rect 17012 7960 17021 8000
rect 17993 7960 18124 8000
rect 18164 7960 18173 8000
rect 21667 7960 21676 8000
rect 21716 7960 22636 8000
rect 22676 7960 22685 8000
rect 23011 7960 23020 8000
rect 23060 7960 23069 8000
rect 26083 7960 26092 8000
rect 26132 7960 26516 8000
rect 26729 7960 26860 8000
rect 26900 7960 26909 8000
rect 27532 7960 28492 8000
rect 28532 7960 28541 8000
rect 28867 7960 28876 8000
rect 28916 7960 28925 8000
rect 14476 7916 14516 7960
rect 16108 7916 16148 7925
rect 23020 7916 23060 7960
rect 24652 7916 24692 7925
rect 26476 7916 26516 7960
rect 27436 7916 27476 7925
rect 14476 7876 14860 7916
rect 14900 7876 14909 7916
rect 15977 7876 16108 7916
rect 16148 7876 16157 7916
rect 18499 7876 18508 7916
rect 18548 7876 23404 7916
rect 23444 7876 23453 7916
rect 24521 7876 24652 7916
rect 24692 7876 24701 7916
rect 26179 7876 26188 7916
rect 26228 7876 26371 7916
rect 26411 7876 26420 7916
rect 26467 7876 26476 7916
rect 26516 7876 26647 7916
rect 26755 7876 26764 7916
rect 26804 7876 26956 7916
rect 26996 7876 27005 7916
rect 27305 7876 27436 7916
rect 27476 7876 27485 7916
rect 16108 7867 16148 7876
rect 24652 7867 24692 7876
rect 27436 7867 27476 7876
rect 10828 7792 11116 7832
rect 11156 7792 12172 7832
rect 12212 7792 12799 7832
rect 12844 7792 15340 7832
rect 15380 7792 15389 7832
rect 16195 7792 16204 7832
rect 16244 7792 22444 7832
rect 22484 7792 22493 7832
rect 24844 7792 26092 7832
rect 26132 7792 26141 7832
rect 0 7664 90 7684
rect 844 7664 884 7792
rect 12759 7748 12799 7792
rect 24844 7748 24884 7792
rect 27532 7748 27572 7960
rect 28972 7916 29012 8128
rect 31852 8044 33580 8084
rect 33620 8044 33629 8084
rect 34867 8044 34876 8084
rect 34916 8044 35692 8084
rect 35732 8044 35741 8084
rect 31852 8000 31892 8044
rect 40396 8000 40436 8212
rect 41932 8168 41972 8296
rect 42700 8252 42740 8380
rect 43180 8252 43220 8464
rect 45004 8336 45044 8464
rect 46278 8336 46368 8356
rect 45004 8296 46368 8336
rect 46278 8276 46368 8296
rect 42700 8212 42932 8252
rect 43180 8212 43268 8252
rect 42892 8168 42932 8212
rect 43228 8168 43268 8212
rect 41932 8128 42748 8168
rect 42788 8128 42797 8168
rect 42892 8128 43132 8168
rect 43172 8128 43181 8168
rect 43228 8128 43900 8168
rect 43940 8128 43949 8168
rect 41731 8044 41740 8084
rect 41780 8044 41972 8084
rect 42019 8044 42028 8084
rect 42068 8044 44180 8084
rect 41932 8000 41972 8044
rect 44140 8000 44180 8044
rect 46278 8000 46368 8020
rect 29059 7960 29068 8000
rect 29108 7960 29452 8000
rect 29492 7960 29501 8000
rect 31171 7960 31180 8000
rect 31220 7960 31564 8000
rect 31604 7960 31613 8000
rect 31843 7960 31852 8000
rect 31892 7960 31901 8000
rect 32419 7960 32428 8000
rect 32468 7960 32716 8000
rect 32756 7960 32765 8000
rect 33187 7960 33196 8000
rect 33236 7960 33484 8000
rect 33524 7960 33533 8000
rect 33763 7960 33772 8000
rect 33812 7960 33868 8000
rect 33908 7960 33943 8000
rect 34121 7960 34252 8000
rect 34292 7960 34301 8000
rect 34627 7960 34636 8000
rect 34676 7960 34924 8000
rect 34964 7960 34973 8000
rect 35203 7960 35212 8000
rect 35252 7960 36076 8000
rect 36116 7960 36125 8000
rect 36490 7960 36499 8000
rect 36539 7960 36596 8000
rect 40396 7960 41836 8000
rect 41876 7960 41885 8000
rect 41932 7960 41980 8000
rect 42020 7960 42029 8000
rect 42211 7960 42220 8000
rect 42260 7960 42269 8000
rect 42316 7960 42604 8000
rect 42644 7960 42653 8000
rect 42979 7960 42988 8000
rect 43028 7960 43316 8000
rect 43363 7960 43372 8000
rect 43412 7960 43421 8000
rect 43747 7960 43756 8000
rect 43796 7960 43805 8000
rect 44131 7960 44140 8000
rect 44180 7960 44189 8000
rect 44393 7960 44524 8000
rect 44564 7960 44573 8000
rect 44777 7960 44908 8000
rect 44948 7960 44957 8000
rect 45763 7960 45772 8000
rect 45812 7960 46368 8000
rect 27946 7876 27955 7916
rect 27995 7876 28780 7916
rect 28820 7876 28829 7916
rect 28972 7876 33004 7916
rect 33044 7876 33053 7916
rect 27907 7792 27916 7832
rect 27956 7792 36460 7832
rect 36500 7792 36509 7832
rect 36556 7748 36596 7960
rect 42220 7916 42260 7960
rect 36643 7876 36652 7916
rect 36692 7876 42260 7916
rect 42316 7832 42356 7960
rect 43276 7916 43316 7960
rect 43267 7876 43276 7916
rect 43316 7876 43325 7916
rect 43372 7832 43412 7960
rect 36739 7792 36748 7832
rect 36788 7792 41596 7832
rect 41636 7792 41645 7832
rect 42028 7792 42356 7832
rect 43180 7792 43412 7832
rect 43459 7792 43468 7832
rect 43508 7792 43516 7832
rect 43556 7792 43639 7832
rect 42028 7748 42068 7792
rect 1459 7708 1468 7748
rect 1508 7708 1517 7748
rect 3859 7708 3868 7748
rect 3908 7708 4148 7748
rect 4243 7708 4252 7748
rect 4292 7708 4396 7748
rect 4436 7708 4445 7748
rect 4627 7708 4636 7748
rect 4676 7708 10868 7748
rect 11491 7708 11500 7748
rect 11540 7708 11692 7748
rect 11732 7708 11741 7748
rect 12355 7708 12364 7748
rect 12404 7708 12508 7748
rect 12548 7708 12557 7748
rect 12759 7708 12844 7748
rect 12884 7708 12893 7748
rect 14707 7708 14716 7748
rect 14756 7708 15820 7748
rect 15860 7708 15869 7748
rect 16291 7708 16300 7748
rect 16340 7708 16349 7748
rect 17155 7708 17164 7748
rect 17204 7708 17212 7748
rect 17252 7708 17335 7748
rect 19651 7708 19660 7748
rect 19700 7708 23156 7748
rect 23251 7708 23260 7748
rect 23300 7708 24884 7748
rect 24940 7708 25852 7748
rect 25892 7708 25901 7748
rect 26371 7708 26380 7748
rect 26420 7708 27572 7748
rect 27619 7708 27628 7748
rect 27668 7708 28108 7748
rect 28148 7708 28157 7748
rect 29683 7708 29692 7748
rect 29732 7708 31412 7748
rect 31642 7708 31651 7748
rect 31691 7708 32419 7748
rect 32459 7708 32468 7748
rect 32873 7708 32956 7748
rect 32996 7708 33004 7748
rect 33044 7708 33053 7748
rect 33178 7708 33187 7748
rect 33236 7708 33367 7748
rect 33715 7708 33724 7748
rect 33764 7708 33964 7748
rect 34004 7708 34013 7748
rect 34099 7708 34108 7748
rect 34148 7708 35980 7748
rect 36020 7708 36029 7748
rect 36137 7708 36259 7748
rect 36308 7708 36835 7748
rect 36875 7708 36884 7748
rect 37123 7708 37132 7748
rect 37172 7708 42068 7748
rect 42115 7708 42124 7748
rect 42164 7708 42364 7748
rect 42404 7708 42413 7748
rect 0 7624 884 7664
rect 0 7604 90 7624
rect 1468 7496 1508 7708
rect 4108 7664 4148 7708
rect 10828 7664 10868 7708
rect 16300 7664 16340 7708
rect 23116 7664 23156 7708
rect 24940 7664 24980 7708
rect 4108 7624 10732 7664
rect 10772 7624 10781 7664
rect 10828 7624 11980 7664
rect 12020 7624 12029 7664
rect 12547 7624 12556 7664
rect 12596 7624 16340 7664
rect 18403 7624 18412 7664
rect 18452 7624 23060 7664
rect 23116 7624 24980 7664
rect 25699 7624 25708 7664
rect 25748 7624 27052 7664
rect 27092 7624 27101 7664
rect 27235 7624 27244 7664
rect 27284 7624 29204 7664
rect 23020 7580 23060 7624
rect 4919 7540 4928 7580
rect 4968 7540 5010 7580
rect 5050 7540 5092 7580
rect 5132 7540 5174 7580
rect 5214 7540 5256 7580
rect 5296 7540 5305 7580
rect 7852 7540 12172 7580
rect 12212 7540 12221 7580
rect 20039 7540 20048 7580
rect 20088 7540 20130 7580
rect 20170 7540 20212 7580
rect 20252 7540 20294 7580
rect 20334 7540 20376 7580
rect 20416 7540 20425 7580
rect 23020 7540 27916 7580
rect 27956 7540 27965 7580
rect 7852 7496 7892 7540
rect 29164 7496 29204 7624
rect 31372 7580 31412 7708
rect 43180 7664 43220 7792
rect 31459 7624 31468 7664
rect 31508 7624 33236 7664
rect 33283 7624 33292 7664
rect 33332 7624 43220 7664
rect 33196 7580 33236 7624
rect 31372 7540 33100 7580
rect 33140 7540 33149 7580
rect 33196 7540 35020 7580
rect 35060 7540 35069 7580
rect 35159 7540 35168 7580
rect 35208 7540 35250 7580
rect 35290 7540 35332 7580
rect 35372 7540 35414 7580
rect 35454 7540 35496 7580
rect 35536 7540 35545 7580
rect 35587 7540 35596 7580
rect 35636 7540 42028 7580
rect 42068 7540 42077 7580
rect 43756 7496 43796 7960
rect 46278 7940 46368 7960
rect 44755 7708 44764 7748
rect 44804 7708 45044 7748
rect 45139 7708 45148 7748
rect 45188 7708 45964 7748
rect 46004 7708 46013 7748
rect 45004 7664 45044 7708
rect 46278 7664 46368 7684
rect 45004 7624 46368 7664
rect 46278 7604 46368 7624
rect 1468 7456 7892 7496
rect 7939 7456 7948 7496
rect 7988 7456 11500 7496
rect 11540 7456 11549 7496
rect 12508 7456 12556 7496
rect 12596 7456 12605 7496
rect 12835 7456 12844 7496
rect 12884 7456 28876 7496
rect 28916 7456 28925 7496
rect 29164 7456 43796 7496
rect 12508 7412 12548 7456
rect 4003 7372 4012 7412
rect 4052 7372 11596 7412
rect 11636 7372 11645 7412
rect 11770 7372 11779 7412
rect 11819 7372 11828 7412
rect 12259 7372 12268 7412
rect 12308 7372 12317 7412
rect 12508 7372 12547 7412
rect 12587 7372 12596 7412
rect 12940 7372 13132 7412
rect 13172 7372 13181 7412
rect 20131 7372 20140 7412
rect 20180 7372 22156 7412
rect 22196 7372 22205 7412
rect 27881 7372 28012 7412
rect 28052 7372 28061 7412
rect 28195 7372 28204 7412
rect 28244 7372 31468 7412
rect 31508 7372 31517 7412
rect 33082 7372 33091 7412
rect 33131 7372 33379 7412
rect 33419 7372 33955 7412
rect 33995 7372 34531 7412
rect 34571 7372 35107 7412
rect 35147 7372 35683 7412
rect 35723 7372 36163 7412
rect 36203 7372 36212 7412
rect 36355 7372 36364 7412
rect 36404 7372 40300 7412
rect 40340 7372 40349 7412
rect 44026 7372 44035 7412
rect 44075 7372 44620 7412
rect 44660 7372 44669 7412
rect 0 7328 90 7348
rect 11788 7328 11828 7372
rect 0 7288 1228 7328
rect 1268 7288 1277 7328
rect 2947 7288 2956 7328
rect 2996 7288 9964 7328
rect 10004 7288 10013 7328
rect 10147 7288 10156 7328
rect 10196 7288 10205 7328
rect 10409 7288 10540 7328
rect 10580 7288 10589 7328
rect 10636 7288 11828 7328
rect 11875 7288 11884 7328
rect 11924 7288 12020 7328
rect 0 7268 90 7288
rect 10156 7244 10196 7288
rect 10636 7244 10676 7288
rect 11980 7244 12020 7288
rect 12124 7288 12172 7328
rect 12212 7288 12221 7328
rect 8035 7204 8044 7244
rect 8084 7204 10100 7244
rect 10147 7204 10156 7244
rect 10196 7204 10243 7244
rect 10313 7204 10435 7244
rect 10484 7204 10493 7244
rect 10540 7204 10676 7244
rect 10060 7160 10100 7204
rect 10540 7160 10580 7204
rect 11692 7193 11708 7233
rect 11748 7193 11757 7233
rect 11866 7204 11875 7244
rect 11915 7204 11924 7244
rect 11980 7204 11992 7244
rect 12032 7204 12041 7244
rect 12124 7235 12164 7288
rect 1219 7120 1228 7160
rect 1268 7120 1277 7160
rect 1324 7120 1612 7160
rect 1652 7120 1661 7160
rect 1843 7120 1852 7160
rect 1892 7120 7892 7160
rect 9667 7120 9676 7160
rect 9716 7120 9964 7160
rect 10004 7120 10013 7160
rect 10060 7120 10580 7160
rect 10985 7120 11116 7160
rect 11156 7120 11165 7160
rect 11347 7120 11356 7160
rect 11396 7120 11500 7160
rect 11540 7120 11549 7160
rect 0 6992 90 7012
rect 1228 6992 1268 7120
rect 0 6952 1268 6992
rect 0 6932 90 6952
rect 0 6656 90 6676
rect 1324 6656 1364 7120
rect 1459 7036 1468 7076
rect 1508 7036 2900 7076
rect 2860 6740 2900 7036
rect 7852 6992 7892 7120
rect 11692 7076 11732 7193
rect 11884 7160 11924 7204
rect 12268 7233 12308 7372
rect 12940 7328 12980 7372
rect 46278 7328 46368 7348
rect 12643 7288 12652 7328
rect 12692 7288 12980 7328
rect 13027 7288 13036 7328
rect 13076 7288 23212 7328
rect 23252 7288 23261 7328
rect 26275 7288 26284 7328
rect 26324 7288 26420 7328
rect 26380 7244 26420 7288
rect 26764 7288 27148 7328
rect 27188 7288 27197 7328
rect 27340 7288 28396 7328
rect 28436 7288 28445 7328
rect 29155 7288 29164 7328
rect 29204 7288 29213 7328
rect 29356 7288 32140 7328
rect 32180 7288 32189 7328
rect 33763 7288 33772 7328
rect 33812 7288 36748 7328
rect 36788 7288 37612 7328
rect 37652 7288 37661 7328
rect 38659 7288 38668 7328
rect 38708 7288 44908 7328
rect 44948 7288 44957 7328
rect 45955 7288 45964 7328
rect 46004 7288 46368 7328
rect 26764 7244 26804 7288
rect 27340 7244 27380 7288
rect 29164 7244 29204 7288
rect 12124 7186 12164 7195
rect 12248 7193 12257 7233
rect 12297 7193 12308 7233
rect 12442 7204 12451 7244
rect 12500 7204 12631 7244
rect 12748 7204 12759 7244
rect 12799 7204 12835 7244
rect 12931 7204 12940 7244
rect 12980 7204 13036 7244
rect 13076 7204 13111 7244
rect 14729 7204 14860 7244
rect 14900 7204 14909 7244
rect 15977 7204 16108 7244
rect 16148 7204 17204 7244
rect 22627 7204 22636 7244
rect 22676 7204 23308 7244
rect 23348 7204 23357 7244
rect 24556 7235 24652 7244
rect 12748 7160 12788 7204
rect 16108 7186 16148 7195
rect 17164 7160 17204 7204
rect 24596 7204 24652 7235
rect 24692 7204 24756 7244
rect 26153 7204 26188 7244
rect 26228 7204 26275 7244
rect 26315 7204 26333 7244
rect 26376 7204 26385 7244
rect 26425 7204 26434 7244
rect 26755 7204 26764 7244
rect 26804 7204 26813 7244
rect 27043 7204 27052 7244
rect 27092 7235 27380 7244
rect 27092 7204 27340 7235
rect 24556 7160 24596 7195
rect 27340 7186 27380 7195
rect 27820 7235 28780 7244
rect 27860 7204 28780 7235
rect 28820 7204 29204 7244
rect 29356 7235 29396 7288
rect 46278 7268 46368 7288
rect 27820 7186 27860 7195
rect 29443 7204 29452 7244
rect 29492 7204 30604 7244
rect 30644 7204 30653 7244
rect 31171 7204 31180 7244
rect 31220 7204 32716 7244
rect 32756 7204 33004 7244
rect 33044 7204 33053 7244
rect 33187 7204 33196 7244
rect 33236 7204 33580 7244
rect 33620 7204 34196 7244
rect 34243 7204 34252 7244
rect 34292 7204 37708 7244
rect 37748 7204 37757 7244
rect 37804 7204 37900 7244
rect 37940 7204 37949 7244
rect 42019 7204 42028 7244
rect 42068 7204 42452 7244
rect 29356 7186 29396 7195
rect 34156 7160 34196 7204
rect 37804 7160 37844 7204
rect 42412 7160 42452 7204
rect 11837 7120 11884 7160
rect 11924 7120 11933 7160
rect 12739 7120 12748 7160
rect 12788 7120 12797 7160
rect 12883 7120 12892 7160
rect 12932 7120 12980 7160
rect 17155 7120 17164 7160
rect 17204 7120 21676 7160
rect 21716 7120 24596 7160
rect 26371 7120 26380 7160
rect 26420 7120 26860 7160
rect 26900 7120 26909 7160
rect 28265 7120 28396 7160
rect 28436 7120 28445 7160
rect 32323 7120 32332 7160
rect 32372 7120 32381 7160
rect 34147 7120 34156 7160
rect 34196 7120 34732 7160
rect 34772 7120 35308 7160
rect 35348 7120 35884 7160
rect 35924 7120 36460 7160
rect 36500 7120 37036 7160
rect 37076 7120 37324 7160
rect 37364 7120 37844 7160
rect 38083 7120 38092 7160
rect 38132 7120 41932 7160
rect 41972 7120 41981 7160
rect 42115 7120 42124 7160
rect 42164 7120 42316 7160
rect 42356 7120 42365 7160
rect 42412 7120 42700 7160
rect 42740 7120 42749 7160
rect 42953 7120 43084 7160
rect 43124 7120 43133 7160
rect 43337 7120 43468 7160
rect 43508 7120 43517 7160
rect 43651 7120 43660 7160
rect 43700 7120 43756 7160
rect 43796 7120 44044 7160
rect 44084 7120 44093 7160
rect 44227 7120 44236 7160
rect 44276 7120 44407 7160
rect 44707 7120 44716 7160
rect 44756 7120 44908 7160
rect 44948 7120 44957 7160
rect 12940 7076 12980 7120
rect 32332 7076 32372 7120
rect 9907 7036 9916 7076
rect 9956 7036 10060 7076
rect 10100 7036 10109 7076
rect 10819 7036 10828 7076
rect 10868 7036 11404 7076
rect 11444 7036 11453 7076
rect 11692 7036 12460 7076
rect 12500 7036 12509 7076
rect 12931 7036 12940 7076
rect 12980 7036 12989 7076
rect 13036 7036 28156 7076
rect 28196 7036 28205 7076
rect 32332 7036 33140 7076
rect 13036 6992 13076 7036
rect 33100 6992 33140 7036
rect 37324 7036 42844 7076
rect 42884 7036 42893 7076
rect 7852 6952 12596 6992
rect 12643 6952 12652 6992
rect 12692 6952 13076 6992
rect 13123 6952 13132 6992
rect 13172 6952 16300 6992
rect 16340 6952 16349 6992
rect 21667 6952 21676 6992
rect 21716 6952 21916 6992
rect 21956 6952 21965 6992
rect 24739 6952 24748 6992
rect 24788 6952 26188 6992
rect 26228 6952 26237 6992
rect 32489 6952 32572 6992
rect 32612 6952 32620 6992
rect 32660 6952 32669 6992
rect 33100 6952 36172 6992
rect 36212 6952 36221 6992
rect 12556 6908 12596 6952
rect 37324 6908 37364 7036
rect 46278 6992 46368 7012
rect 41683 6952 41692 6992
rect 41732 6952 41780 6992
rect 41827 6952 41836 6992
rect 41876 6952 42076 6992
rect 42116 6952 42125 6992
rect 42220 6952 42460 6992
rect 42500 6952 42509 6992
rect 42595 6952 42604 6992
rect 42644 6952 43228 6992
rect 43268 6952 43351 6992
rect 44467 6952 44476 6992
rect 44516 6952 45044 6992
rect 45139 6952 45148 6992
rect 45188 6952 46368 6992
rect 10243 6868 10252 6908
rect 10292 6868 11788 6908
rect 11828 6868 11837 6908
rect 12556 6868 14476 6908
rect 14516 6868 14525 6908
rect 18019 6868 18028 6908
rect 18068 6868 37364 6908
rect 41740 6908 41780 6952
rect 41740 6868 41876 6908
rect 3679 6784 3688 6824
rect 3728 6784 3770 6824
rect 3810 6784 3852 6824
rect 3892 6784 3934 6824
rect 3974 6784 4016 6824
rect 4056 6784 4065 6824
rect 9955 6784 9964 6824
rect 10004 6784 17780 6824
rect 18799 6784 18808 6824
rect 18848 6784 18890 6824
rect 18930 6784 18972 6824
rect 19012 6784 19054 6824
rect 19094 6784 19136 6824
rect 19176 6784 19185 6824
rect 33919 6784 33928 6824
rect 33968 6784 34010 6824
rect 34050 6784 34092 6824
rect 34132 6784 34174 6824
rect 34214 6784 34256 6824
rect 34296 6784 34305 6824
rect 34915 6784 34924 6824
rect 34964 6784 41740 6824
rect 41780 6784 41789 6824
rect 2860 6700 10004 6740
rect 10051 6700 10060 6740
rect 10100 6700 13076 6740
rect 9964 6656 10004 6700
rect 0 6616 1364 6656
rect 7939 6616 7948 6656
rect 7988 6616 9388 6656
rect 9428 6616 9437 6656
rect 9964 6616 11116 6656
rect 11156 6616 11165 6656
rect 11242 6616 11251 6656
rect 11291 6616 12844 6656
rect 12884 6616 12893 6656
rect 0 6596 90 6616
rect 13036 6572 13076 6700
rect 17740 6656 17780 6784
rect 41836 6740 41876 6868
rect 18211 6700 18220 6740
rect 18260 6700 41876 6740
rect 17740 6616 22540 6656
rect 22580 6616 22589 6656
rect 30787 6616 30796 6656
rect 30836 6616 42124 6656
rect 42164 6616 42173 6656
rect 1459 6532 1468 6572
rect 1508 6532 11828 6572
rect 11875 6532 11884 6572
rect 11924 6532 12172 6572
rect 12212 6532 12221 6572
rect 13036 6532 23596 6572
rect 23636 6532 23645 6572
rect 30211 6532 30220 6572
rect 30260 6532 42028 6572
rect 42068 6532 42077 6572
rect 11788 6488 11828 6532
rect 42220 6488 42260 6952
rect 45004 6656 45044 6952
rect 46278 6932 46368 6952
rect 46278 6656 46368 6676
rect 45004 6616 46368 6656
rect 46278 6596 46368 6616
rect 1219 6448 1228 6488
rect 1268 6448 1277 6488
rect 1603 6448 1612 6488
rect 1652 6448 1661 6488
rect 5993 6448 6124 6488
rect 6164 6448 6548 6488
rect 8995 6448 9004 6488
rect 9044 6448 9908 6488
rect 9955 6448 9964 6488
rect 10004 6448 10135 6488
rect 11788 6448 14860 6488
rect 14900 6448 14909 6488
rect 17033 6448 17164 6488
rect 17204 6448 17213 6488
rect 19843 6448 19852 6488
rect 19892 6448 42260 6488
rect 42307 6448 42316 6488
rect 42356 6448 44524 6488
rect 44564 6448 44573 6488
rect 0 6320 90 6340
rect 1228 6320 1268 6448
rect 0 6280 1268 6320
rect 0 6260 90 6280
rect 0 5984 90 6004
rect 1612 5984 1652 6448
rect 6508 6404 6548 6448
rect 9868 6404 9908 6448
rect 10540 6404 10580 6413
rect 6499 6364 6508 6404
rect 6548 6364 6557 6404
rect 7755 6364 7764 6404
rect 7804 6364 8908 6404
rect 8948 6364 8957 6404
rect 9466 6364 9475 6404
rect 9515 6364 9524 6404
rect 9571 6364 9580 6404
rect 9620 6364 9751 6404
rect 9868 6364 10060 6404
rect 10100 6364 10109 6404
rect 11050 6364 11059 6404
rect 11099 6364 11212 6404
rect 11252 6364 11261 6404
rect 11491 6364 11500 6404
rect 11540 6364 11549 6404
rect 11657 6364 11779 6404
rect 11828 6364 11837 6404
rect 15811 6364 15820 6404
rect 15860 6364 17452 6404
rect 17492 6364 17501 6404
rect 17635 6364 17644 6404
rect 17684 6364 21772 6404
rect 21812 6364 21821 6404
rect 30979 6364 30988 6404
rect 31028 6364 37996 6404
rect 38036 6364 38045 6404
rect 38179 6364 38188 6404
rect 38228 6364 43220 6404
rect 9484 6320 9524 6364
rect 10540 6320 10580 6364
rect 11500 6320 11540 6364
rect 43180 6320 43220 6364
rect 46278 6320 46368 6340
rect 2860 6280 8084 6320
rect 9484 6280 10252 6320
rect 10292 6280 10301 6320
rect 10380 6280 10444 6320
rect 10484 6280 11444 6320
rect 11491 6280 11500 6320
rect 11540 6280 11587 6320
rect 11683 6280 11692 6320
rect 11732 6280 11884 6320
rect 11924 6280 11933 6320
rect 11980 6280 25132 6320
rect 25172 6280 25181 6320
rect 30403 6280 30412 6320
rect 30452 6280 43084 6320
rect 43124 6280 43133 6320
rect 43180 6280 43468 6320
rect 43508 6280 43517 6320
rect 44236 6280 44908 6320
rect 44948 6280 44957 6320
rect 45187 6280 45196 6320
rect 45236 6280 46368 6320
rect 2860 6236 2900 6280
rect 1843 6196 1852 6236
rect 1892 6196 2900 6236
rect 6355 6196 6364 6236
rect 6404 6196 7988 6236
rect 4919 6028 4928 6068
rect 4968 6028 5010 6068
rect 5050 6028 5092 6068
rect 5132 6028 5174 6068
rect 5214 6028 5256 6068
rect 5296 6028 5305 6068
rect 0 5944 1652 5984
rect 7948 5984 7988 6196
rect 8044 6068 8084 6280
rect 11404 6236 11444 6280
rect 11980 6236 12020 6280
rect 44236 6236 44276 6280
rect 46278 6260 46368 6280
rect 9235 6196 9244 6236
rect 9284 6196 10636 6236
rect 10676 6196 10685 6236
rect 11395 6196 11404 6236
rect 11444 6196 12020 6236
rect 16867 6196 16876 6236
rect 16916 6196 16924 6236
rect 16964 6196 17047 6236
rect 17164 6196 42316 6236
rect 42356 6196 42365 6236
rect 43529 6196 43651 6236
rect 43700 6196 43939 6236
rect 43979 6196 44227 6236
rect 44267 6196 44276 6236
rect 44755 6196 44764 6236
rect 44804 6196 46196 6236
rect 17164 6068 17204 6196
rect 46156 6152 46196 6196
rect 17443 6112 17452 6152
rect 17492 6112 44236 6152
rect 44276 6112 44285 6152
rect 46156 6112 46252 6152
rect 46292 6112 46301 6152
rect 8044 6028 13804 6068
rect 13844 6028 13853 6068
rect 14083 6028 14092 6068
rect 14132 6028 17204 6068
rect 20039 6028 20048 6068
rect 20088 6028 20130 6068
rect 20170 6028 20212 6068
rect 20252 6028 20294 6068
rect 20334 6028 20376 6068
rect 20416 6028 20425 6068
rect 30595 6028 30604 6068
rect 30644 6028 35060 6068
rect 35159 6028 35168 6068
rect 35208 6028 35250 6068
rect 35290 6028 35332 6068
rect 35372 6028 35414 6068
rect 35454 6028 35496 6068
rect 35536 6028 35545 6068
rect 35020 5984 35060 6028
rect 46278 5984 46368 6004
rect 7948 5944 34924 5984
rect 34964 5944 34973 5984
rect 35020 5944 38188 5984
rect 38228 5944 38237 5984
rect 46243 5944 46252 5984
rect 46292 5944 46368 5984
rect 0 5924 90 5944
rect 46278 5924 46368 5944
rect 11107 5860 11116 5900
rect 11156 5860 11788 5900
rect 11828 5860 11837 5900
rect 12739 5860 12748 5900
rect 12788 5860 13180 5900
rect 13220 5860 13229 5900
rect 18595 5860 18604 5900
rect 18644 5860 42604 5900
rect 42644 5860 42653 5900
rect 43738 5860 43747 5900
rect 43787 5860 44227 5900
rect 44267 5860 44276 5900
rect 9341 5776 9388 5816
rect 9428 5776 9437 5816
rect 9484 5776 9580 5816
rect 9620 5776 9772 5816
rect 9812 5776 21580 5816
rect 21620 5776 21629 5816
rect 21763 5776 21772 5816
rect 21812 5776 41836 5816
rect 41876 5776 41885 5816
rect 9388 5732 9428 5776
rect 9484 5732 9524 5776
rect 9370 5692 9379 5732
rect 9419 5692 9428 5732
rect 9475 5692 9484 5732
rect 9524 5692 9533 5732
rect 9833 5692 9868 5732
rect 9908 5692 9964 5732
rect 10004 5692 10013 5732
rect 10313 5692 10444 5732
rect 10484 5692 10493 5732
rect 10793 5692 10924 5732
rect 10964 5692 10973 5732
rect 13193 5692 13324 5732
rect 13364 5692 13373 5732
rect 23020 5692 44948 5732
rect 10444 5674 10484 5683
rect 10924 5674 10964 5683
rect 0 5648 90 5668
rect 23020 5648 23060 5692
rect 44908 5648 44948 5692
rect 46278 5648 46368 5668
rect 0 5608 1228 5648
rect 1268 5608 1277 5648
rect 1603 5608 1612 5648
rect 1652 5608 1661 5648
rect 1865 5608 1996 5648
rect 2036 5608 2045 5648
rect 9929 5608 9964 5648
rect 10004 5608 10060 5648
rect 10100 5608 10109 5648
rect 11273 5608 11308 5648
rect 11348 5608 11404 5648
rect 11444 5608 11453 5648
rect 11539 5608 11548 5648
rect 11588 5608 12556 5648
rect 12596 5608 12605 5648
rect 15235 5608 15244 5648
rect 15284 5608 23060 5648
rect 43529 5608 43660 5648
rect 43700 5608 43709 5648
rect 43939 5608 43948 5648
rect 43988 5608 44044 5648
rect 44084 5608 44119 5648
rect 44515 5608 44524 5648
rect 44564 5608 44573 5648
rect 44899 5608 44908 5648
rect 44948 5608 44957 5648
rect 45065 5608 45148 5648
rect 45188 5608 45196 5648
rect 45236 5608 45245 5648
rect 45379 5608 45388 5648
rect 45428 5608 46368 5648
rect 0 5588 90 5608
rect 1612 5564 1652 5608
rect 44524 5564 44564 5608
rect 46278 5588 46368 5608
rect 844 5524 1652 5564
rect 24067 5524 24076 5564
rect 24116 5524 44564 5564
rect 0 5312 90 5332
rect 844 5312 884 5524
rect 1459 5440 1468 5480
rect 1508 5440 1748 5480
rect 1843 5440 1852 5480
rect 1892 5440 2132 5480
rect 2227 5440 2236 5480
rect 2276 5440 5740 5480
rect 5780 5440 5789 5480
rect 44755 5440 44764 5480
rect 44804 5440 45044 5480
rect 0 5272 884 5312
rect 0 5252 90 5272
rect 1708 5228 1748 5440
rect 2092 5396 2132 5440
rect 2092 5356 21868 5396
rect 21908 5356 21917 5396
rect 45004 5312 45044 5440
rect 46278 5312 46368 5332
rect 3679 5272 3688 5312
rect 3728 5272 3770 5312
rect 3810 5272 3852 5312
rect 3892 5272 3934 5312
rect 3974 5272 4016 5312
rect 4056 5272 4065 5312
rect 18799 5272 18808 5312
rect 18848 5272 18890 5312
rect 18930 5272 18972 5312
rect 19012 5272 19054 5312
rect 19094 5272 19136 5312
rect 19176 5272 19185 5312
rect 33919 5272 33928 5312
rect 33968 5272 34010 5312
rect 34050 5272 34092 5312
rect 34132 5272 34174 5312
rect 34214 5272 34256 5312
rect 34296 5272 34305 5312
rect 45004 5272 46368 5312
rect 46278 5252 46368 5272
rect 1708 5188 24268 5228
rect 24308 5188 24317 5228
rect 33283 5188 33292 5228
rect 33332 5188 42892 5228
rect 42932 5188 42941 5228
rect 20899 5104 20908 5144
rect 20948 5104 32956 5144
rect 32996 5104 33005 5144
rect 41635 5104 41644 5144
rect 41684 5104 42844 5144
rect 42884 5104 42893 5144
rect 45139 5104 45148 5144
rect 45188 5104 45388 5144
rect 45428 5104 45437 5144
rect 1699 5020 1708 5060
rect 1748 5020 23060 5060
rect 0 4976 90 4996
rect 23020 4976 23060 5020
rect 31468 5020 32756 5060
rect 35971 5020 35980 5060
rect 36020 5020 44564 5060
rect 0 4936 1996 4976
rect 2036 4936 2045 4976
rect 23020 4936 30988 4976
rect 31028 4936 31037 4976
rect 0 4916 90 4936
rect 30988 4892 31028 4936
rect 17827 4852 17836 4892
rect 17876 4852 23060 4892
rect 30988 4852 31372 4892
rect 31412 4852 31421 4892
rect 23020 4808 23060 4852
rect 31468 4808 31508 5020
rect 32620 4892 32660 4901
rect 32131 4852 32140 4892
rect 32180 4852 32620 4892
rect 32716 4892 32756 5020
rect 44524 4976 44564 5020
rect 46278 4976 46368 4996
rect 32899 4936 32908 4976
rect 32948 4936 33196 4976
rect 33236 4936 33245 4976
rect 43075 4936 43084 4976
rect 43124 4936 43133 4976
rect 44515 4936 44524 4976
rect 44564 4936 44573 4976
rect 44899 4936 44908 4976
rect 44948 4936 44957 4976
rect 45763 4936 45772 4976
rect 45812 4936 46368 4976
rect 43084 4892 43124 4936
rect 32716 4852 43124 4892
rect 43171 4852 43180 4892
rect 43220 4852 43660 4892
rect 43700 4852 44236 4892
rect 44276 4852 44285 4892
rect 32620 4843 32660 4852
rect 44908 4808 44948 4936
rect 46278 4916 46368 4936
rect 23020 4768 31508 4808
rect 32716 4768 33140 4808
rect 39139 4768 39148 4808
rect 39188 4768 44948 4808
rect 32716 4724 32756 4768
rect 33100 4724 33140 4768
rect 31219 4684 31228 4724
rect 31268 4684 32756 4724
rect 32803 4684 32812 4724
rect 32852 4684 32861 4724
rect 33100 4684 39052 4724
rect 39092 4684 39101 4724
rect 43450 4684 43459 4724
rect 43499 4684 43651 4724
rect 43691 4684 43939 4724
rect 43988 4684 43997 4724
rect 44755 4684 44764 4724
rect 44804 4684 45044 4724
rect 0 4640 90 4660
rect 32812 4640 32852 4684
rect 45004 4640 45044 4684
rect 46278 4640 46368 4660
rect 0 4600 23060 4640
rect 32812 4600 34348 4640
rect 34388 4600 34397 4640
rect 45004 4600 46368 4640
rect 0 4580 90 4600
rect 23020 4556 23060 4600
rect 46278 4580 46368 4600
rect 4919 4516 4928 4556
rect 4968 4516 5010 4556
rect 5050 4516 5092 4556
rect 5132 4516 5174 4556
rect 5214 4516 5256 4556
rect 5296 4516 5305 4556
rect 20039 4516 20048 4556
rect 20088 4516 20130 4556
rect 20170 4516 20212 4556
rect 20252 4516 20294 4556
rect 20334 4516 20376 4556
rect 20416 4516 20425 4556
rect 23020 4516 33772 4556
rect 33812 4516 33821 4556
rect 35159 4516 35168 4556
rect 35208 4516 35250 4556
rect 35290 4516 35332 4556
rect 35372 4516 35414 4556
rect 35454 4516 35496 4556
rect 35536 4516 35545 4556
rect 32035 4432 32044 4472
rect 32084 4432 32428 4472
rect 32468 4432 32908 4472
rect 32948 4432 32957 4472
rect 33379 4432 33388 4472
rect 33428 4432 33908 4472
rect 33868 4388 33908 4432
rect 19747 4348 19756 4388
rect 19796 4348 19996 4388
rect 20036 4348 20045 4388
rect 21379 4348 21388 4388
rect 21428 4348 21908 4388
rect 0 4304 90 4324
rect 21868 4304 21908 4348
rect 23788 4348 24212 4388
rect 23788 4304 23828 4348
rect 24172 4304 24212 4348
rect 31372 4348 33196 4388
rect 33236 4348 33245 4388
rect 33475 4348 33484 4388
rect 33524 4348 33533 4388
rect 33868 4348 34100 4388
rect 31372 4304 31412 4348
rect 33484 4304 33524 4348
rect 34060 4304 34100 4348
rect 40108 4348 42164 4388
rect 43817 4348 43939 4388
rect 43988 4348 44611 4388
rect 44651 4348 44660 4388
rect 40108 4304 40148 4348
rect 42124 4304 42164 4348
rect 46278 4304 46368 4324
rect 0 4264 19412 4304
rect 0 4244 90 4264
rect 19372 4220 19412 4264
rect 20188 4264 21812 4304
rect 21868 4264 23828 4304
rect 23945 4264 24028 4304
rect 24068 4264 24076 4304
rect 24116 4264 24125 4304
rect 24172 4264 25556 4304
rect 25603 4264 25612 4304
rect 25652 4264 25940 4304
rect 26275 4264 26284 4304
rect 26324 4264 26516 4304
rect 27043 4264 27052 4304
rect 27092 4264 27100 4304
rect 27140 4264 27223 4304
rect 27340 4264 31412 4304
rect 31459 4264 31468 4304
rect 31508 4264 32332 4304
rect 32372 4264 33044 4304
rect 33484 4264 33964 4304
rect 34004 4264 34013 4304
rect 34060 4264 40148 4304
rect 40195 4264 40204 4304
rect 40244 4264 41980 4304
rect 42020 4264 42029 4304
rect 42124 4264 42748 4304
rect 42788 4264 42797 4304
rect 45139 4264 45148 4304
rect 45188 4264 45772 4304
rect 45812 4264 45821 4304
rect 45955 4264 45964 4304
rect 46004 4264 46368 4304
rect 20188 4220 20228 4264
rect 7267 4180 7276 4220
rect 7316 4180 9676 4220
rect 9716 4180 9725 4220
rect 9772 4180 9785 4220
rect 9825 4180 9859 4220
rect 9929 4180 10060 4220
rect 10100 4180 10109 4220
rect 17644 4180 18028 4220
rect 18068 4180 18077 4220
rect 19145 4180 19276 4220
rect 19316 4180 19325 4220
rect 19372 4180 20228 4220
rect 20332 4180 21580 4220
rect 21620 4180 21629 4220
rect 21676 4211 21716 4220
rect 0 3968 90 3988
rect 9676 3968 9716 4180
rect 9772 4136 9812 4180
rect 17644 4136 17684 4180
rect 19276 4162 19316 4171
rect 20332 4136 20372 4180
rect 21676 4136 21716 4171
rect 9763 4096 9772 4136
rect 9812 4096 9821 4136
rect 11971 4096 11980 4136
rect 12020 4096 17644 4136
rect 17684 4096 17693 4136
rect 17801 4096 17884 4136
rect 17924 4096 17932 4136
rect 17972 4096 17981 4136
rect 19577 4096 19660 4136
rect 19700 4096 19708 4136
rect 19748 4096 19757 4136
rect 19843 4096 19852 4136
rect 19892 4096 20332 4136
rect 20372 4096 20381 4136
rect 20969 4096 21100 4136
rect 21140 4096 21149 4136
rect 21331 4096 21340 4136
rect 21380 4096 21484 4136
rect 21524 4096 21533 4136
rect 21629 4096 21676 4136
rect 21716 4096 21725 4136
rect 21772 4052 21812 4264
rect 21955 4180 21964 4220
rect 22004 4180 22924 4220
rect 22964 4180 22973 4220
rect 24163 4180 24172 4220
rect 24212 4180 24221 4220
rect 25289 4180 25420 4220
rect 25460 4180 25469 4220
rect 24172 4136 24212 4180
rect 25420 4162 25460 4171
rect 21859 4096 21868 4136
rect 21908 4096 23788 4136
rect 23828 4096 24212 4136
rect 25516 4136 25556 4264
rect 25900 4220 25940 4264
rect 26476 4220 26516 4264
rect 27340 4220 27380 4264
rect 33004 4220 33044 4264
rect 46278 4244 46368 4264
rect 25891 4180 25900 4220
rect 25940 4180 25949 4220
rect 26033 4180 26092 4220
rect 26132 4180 26155 4220
rect 26195 4180 26213 4220
rect 26268 4180 26277 4220
rect 26317 4180 26420 4220
rect 26476 4180 27380 4220
rect 29897 4180 30028 4220
rect 30068 4180 30077 4220
rect 30499 4180 30508 4220
rect 30548 4211 31316 4220
rect 30548 4180 31276 4211
rect 26380 4136 26420 4180
rect 31363 4180 31372 4220
rect 31412 4180 31747 4220
rect 31787 4180 31796 4220
rect 31843 4180 31852 4220
rect 31892 4180 32023 4220
rect 32227 4180 32236 4220
rect 32276 4180 32524 4220
rect 32564 4180 32573 4220
rect 32812 4211 32852 4220
rect 31276 4136 31316 4171
rect 33004 4211 33332 4220
rect 33004 4180 33292 4211
rect 25516 4096 26188 4136
rect 26228 4096 26237 4136
rect 26380 4096 26516 4136
rect 26563 4096 26572 4136
rect 26612 4096 26764 4136
rect 26804 4096 26813 4136
rect 26956 4096 27340 4136
rect 27380 4096 27389 4136
rect 27907 4096 27916 4136
rect 27956 4096 31180 4136
rect 31220 4096 31229 4136
rect 31276 4096 32140 4136
rect 32180 4096 32189 4136
rect 32297 4096 32332 4136
rect 32372 4096 32428 4136
rect 32468 4096 32477 4136
rect 13123 4012 13132 4052
rect 13172 4012 21620 4052
rect 21772 4012 26284 4052
rect 26324 4012 26333 4052
rect 0 3928 2900 3968
rect 9379 3928 9388 3968
rect 9428 3928 9437 3968
rect 9676 3928 15628 3968
rect 15668 3928 19180 3968
rect 19220 3928 19229 3968
rect 19459 3928 19468 3968
rect 19508 3928 19756 3968
rect 19796 3928 19805 3968
rect 19852 3928 20092 3968
rect 20132 3928 20141 3968
rect 21353 3928 21484 3968
rect 21524 3928 21533 3968
rect 0 3908 90 3928
rect 0 3632 90 3652
rect 0 3592 652 3632
rect 692 3592 701 3632
rect 0 3572 90 3592
rect 0 3296 90 3316
rect 0 3256 1324 3296
rect 1364 3256 1373 3296
rect 0 3236 90 3256
rect 0 2960 90 2980
rect 2860 2960 2900 3928
rect 3679 3760 3688 3800
rect 3728 3760 3770 3800
rect 3810 3760 3852 3800
rect 3892 3760 3934 3800
rect 3974 3760 4016 3800
rect 4056 3760 4065 3800
rect 9161 3592 9244 3632
rect 9284 3592 9292 3632
rect 9332 3592 9341 3632
rect 9388 3464 9428 3928
rect 19852 3884 19892 3928
rect 16483 3844 16492 3884
rect 16532 3844 19892 3884
rect 21580 3884 21620 4012
rect 26476 3968 26516 4096
rect 26956 4052 26996 4096
rect 32812 4052 32852 4171
rect 33571 4180 33580 4220
rect 33620 4180 34073 4220
rect 34113 4180 34122 4220
rect 34339 4180 34348 4220
rect 34388 4180 34519 4220
rect 40291 4180 40300 4220
rect 40340 4180 44372 4220
rect 33292 4162 33332 4171
rect 38249 4096 38380 4136
rect 38420 4096 38572 4136
rect 38612 4096 38621 4136
rect 38851 4096 38860 4136
rect 38900 4096 42220 4136
rect 42260 4096 42269 4136
rect 42595 4096 42604 4136
rect 42644 4096 42653 4136
rect 42857 4096 42988 4136
rect 43028 4096 43037 4136
rect 43363 4096 43372 4136
rect 43412 4096 43468 4136
rect 43508 4096 43543 4136
rect 43625 4096 43756 4136
rect 43796 4096 43805 4136
rect 44227 4096 44236 4136
rect 44276 4096 44285 4136
rect 42604 4052 42644 4096
rect 44236 4052 44276 4096
rect 26563 4012 26572 4052
rect 26612 4012 26996 4052
rect 27427 4012 27436 4052
rect 27476 4012 28588 4052
rect 28628 4012 28637 4052
rect 29731 4012 29740 4052
rect 29780 4012 32908 4052
rect 32948 4012 33012 4052
rect 33475 4012 33484 4052
rect 33524 4012 40436 4052
rect 41443 4012 41452 4052
rect 41492 4012 42644 4052
rect 42892 4012 44276 4052
rect 40396 3968 40436 4012
rect 21763 3928 21772 3968
rect 21812 3928 26572 3968
rect 26612 3928 26676 3968
rect 26995 3928 27004 3968
rect 27044 3928 31660 3968
rect 31700 3928 31709 3968
rect 32419 3928 32428 3968
rect 32468 3928 33676 3968
rect 33716 3928 33725 3968
rect 34243 3928 34252 3968
rect 34292 3928 38668 3968
rect 38708 3928 38717 3968
rect 38803 3928 38812 3968
rect 38852 3928 40300 3968
rect 40340 3928 40349 3968
rect 40396 3928 42364 3968
rect 42404 3928 42413 3968
rect 42892 3884 42932 4012
rect 44332 3968 44372 4180
rect 44611 4096 44620 4136
rect 44660 4096 44908 4136
rect 44948 4096 44957 4136
rect 44467 4012 44476 4052
rect 44516 4012 45428 4052
rect 45388 3968 45428 4012
rect 46278 3968 46368 3988
rect 43049 3928 43132 3968
rect 43172 3928 43180 3968
rect 43220 3928 43229 3968
rect 43276 3928 43516 3968
rect 43556 3928 43565 3968
rect 44332 3928 44948 3968
rect 45388 3928 46368 3968
rect 43276 3884 43316 3928
rect 21580 3844 33140 3884
rect 33187 3844 33196 3884
rect 33236 3844 42932 3884
rect 42979 3844 42988 3884
rect 43028 3844 43316 3884
rect 33100 3800 33140 3844
rect 18799 3760 18808 3800
rect 18848 3760 18890 3800
rect 18930 3760 18972 3800
rect 19012 3760 19054 3800
rect 19094 3760 19136 3800
rect 19176 3760 19185 3800
rect 19651 3760 19660 3800
rect 19700 3760 25036 3800
rect 25076 3760 25085 3800
rect 25507 3760 25516 3800
rect 25556 3760 33004 3800
rect 33044 3760 33053 3800
rect 33100 3760 33716 3800
rect 33919 3760 33928 3800
rect 33968 3760 34010 3800
rect 34050 3760 34092 3800
rect 34132 3760 34174 3800
rect 34214 3760 34256 3800
rect 34296 3760 34305 3800
rect 38947 3760 38956 3800
rect 38996 3760 43220 3800
rect 33676 3716 33716 3760
rect 17731 3676 17740 3716
rect 17780 3676 21388 3716
rect 21428 3676 21437 3716
rect 21571 3676 21580 3716
rect 21620 3676 25748 3716
rect 25795 3676 25804 3716
rect 25844 3676 31852 3716
rect 31892 3676 31901 3716
rect 32515 3676 32524 3716
rect 32564 3676 32756 3716
rect 32899 3676 32908 3716
rect 32948 3676 33620 3716
rect 33676 3676 43084 3716
rect 43124 3676 43133 3716
rect 9545 3592 9628 3632
rect 9668 3592 9676 3632
rect 9716 3592 9725 3632
rect 10915 3592 10924 3632
rect 10964 3592 11212 3632
rect 11252 3592 11261 3632
rect 12019 3592 12028 3632
rect 12068 3592 13132 3632
rect 13172 3592 13181 3632
rect 13315 3592 13324 3632
rect 13364 3592 13612 3632
rect 13652 3592 13661 3632
rect 13987 3592 13996 3632
rect 14036 3592 15860 3632
rect 17251 3592 17260 3632
rect 17300 3592 18172 3632
rect 18212 3592 18221 3632
rect 18316 3592 19276 3632
rect 19316 3592 21676 3632
rect 21716 3592 21725 3632
rect 23299 3592 23308 3632
rect 23348 3592 25612 3632
rect 25652 3592 25661 3632
rect 15820 3548 15860 3592
rect 18316 3548 18356 3592
rect 25708 3548 25748 3676
rect 32716 3632 32756 3676
rect 26179 3592 26188 3632
rect 26228 3592 32572 3632
rect 32612 3592 32621 3632
rect 32716 3592 33140 3632
rect 33100 3548 33140 3592
rect 15043 3508 15052 3548
rect 15092 3508 15572 3548
rect 15820 3508 17788 3548
rect 17828 3508 17837 3548
rect 17932 3508 18356 3548
rect 18787 3508 18796 3548
rect 18836 3508 21100 3548
rect 21140 3508 21149 3548
rect 21571 3508 21580 3548
rect 21620 3508 25036 3548
rect 25076 3508 25085 3548
rect 25219 3508 25228 3548
rect 25268 3508 25652 3548
rect 25708 3508 26668 3548
rect 26708 3508 26717 3548
rect 26851 3508 26860 3548
rect 26900 3508 27284 3548
rect 27859 3508 27868 3548
rect 27908 3508 28684 3548
rect 28724 3508 28733 3548
rect 29443 3508 29452 3548
rect 29492 3508 31372 3548
rect 31412 3508 31421 3548
rect 32803 3508 32812 3548
rect 32852 3508 32956 3548
rect 32996 3508 33005 3548
rect 33100 3508 33236 3548
rect 15532 3464 15572 3508
rect 17932 3464 17972 3508
rect 25612 3464 25652 3508
rect 27244 3464 27284 3508
rect 30796 3464 30836 3508
rect 33196 3464 33236 3508
rect 33580 3464 33620 3676
rect 43180 3632 43220 3760
rect 38563 3592 38572 3632
rect 38612 3592 42748 3632
rect 42788 3592 42797 3632
rect 43180 3592 43900 3632
rect 43940 3592 43949 3632
rect 34435 3508 34444 3548
rect 34484 3508 41740 3548
rect 41780 3508 41789 3548
rect 41923 3508 41932 3548
rect 41972 3508 42268 3548
rect 42308 3508 42317 3548
rect 42412 3508 43132 3548
rect 43172 3508 43181 3548
rect 43660 3508 44180 3548
rect 42412 3464 42452 3508
rect 8873 3424 9004 3464
rect 9044 3424 9053 3464
rect 9379 3424 9388 3464
rect 9428 3424 9437 3464
rect 11587 3424 11596 3464
rect 11636 3424 11788 3464
rect 11828 3424 12212 3464
rect 9004 3380 9044 3424
rect 11020 3380 11060 3389
rect 12172 3380 12212 3424
rect 13420 3424 15092 3464
rect 15305 3424 15436 3464
rect 15476 3424 15485 3464
rect 15532 3424 15772 3464
rect 15812 3424 15821 3464
rect 16003 3424 16012 3464
rect 16052 3424 16204 3464
rect 16244 3424 16253 3464
rect 17452 3424 17972 3464
rect 18019 3424 18028 3464
rect 18068 3424 18220 3464
rect 18260 3424 18269 3464
rect 18403 3424 18412 3464
rect 18452 3424 18461 3464
rect 18787 3424 18796 3464
rect 18836 3424 19372 3464
rect 19412 3424 19421 3464
rect 19555 3424 19564 3464
rect 19604 3424 19852 3464
rect 19892 3424 19901 3464
rect 20140 3424 20524 3464
rect 20564 3424 21388 3464
rect 21428 3424 21437 3464
rect 21955 3424 21964 3464
rect 22004 3424 22828 3464
rect 22868 3424 22877 3464
rect 25612 3424 27004 3464
rect 27044 3424 27053 3464
rect 27235 3424 27244 3464
rect 27284 3424 27293 3464
rect 27497 3424 27628 3464
rect 27668 3424 27677 3464
rect 30019 3424 30028 3464
rect 30068 3424 30220 3464
rect 30260 3424 30269 3464
rect 30700 3424 30836 3464
rect 30883 3424 30892 3464
rect 30932 3424 31180 3464
rect 31220 3424 31229 3464
rect 31843 3424 31852 3464
rect 31892 3424 32812 3464
rect 32852 3424 32861 3464
rect 33187 3424 33196 3464
rect 33236 3424 33245 3464
rect 33571 3424 33580 3464
rect 33620 3424 33629 3464
rect 37507 3424 37516 3464
rect 37556 3424 37804 3464
rect 37844 3424 37853 3464
rect 38057 3424 38188 3464
rect 38228 3424 38572 3464
rect 38612 3424 38621 3464
rect 39043 3424 39052 3464
rect 39092 3424 39340 3464
rect 39380 3424 39389 3464
rect 39523 3424 39532 3464
rect 39572 3424 39724 3464
rect 39764 3424 39773 3464
rect 40099 3424 40108 3464
rect 40148 3424 42452 3464
rect 42499 3424 42508 3464
rect 42548 3424 42557 3464
rect 42857 3424 42988 3464
rect 43028 3424 43037 3464
rect 43241 3424 43372 3464
rect 43412 3424 43421 3464
rect 13420 3380 13460 3424
rect 15052 3380 15092 3424
rect 15436 3380 15476 3424
rect 17452 3380 17492 3424
rect 9004 3340 9772 3380
rect 9812 3340 9821 3380
rect 12163 3340 12172 3380
rect 12212 3340 12221 3380
rect 13673 3340 13804 3380
rect 13844 3340 13853 3380
rect 14921 3340 15052 3380
rect 15092 3340 15101 3380
rect 15436 3340 16204 3380
rect 16244 3340 16253 3380
rect 11020 3296 11060 3340
rect 13420 3296 13460 3340
rect 15052 3331 15092 3340
rect 17452 3331 17492 3340
rect 18412 3296 18452 3424
rect 20140 3380 20180 3424
rect 25516 3380 25556 3389
rect 27628 3380 27668 3424
rect 29260 3380 29300 3389
rect 30700 3380 30740 3424
rect 31756 3380 31796 3389
rect 42508 3380 42548 3424
rect 43660 3380 43700 3508
rect 44140 3464 44180 3508
rect 44908 3464 44948 3928
rect 46278 3908 46368 3928
rect 46278 3632 46368 3652
rect 45139 3592 45148 3632
rect 45188 3592 45964 3632
rect 46004 3592 46013 3632
rect 46147 3592 46156 3632
rect 46196 3592 46368 3632
rect 46278 3572 46368 3592
rect 43747 3424 43756 3464
rect 43796 3424 43805 3464
rect 44131 3424 44140 3464
rect 44180 3424 44189 3464
rect 44393 3424 44524 3464
rect 44564 3424 44573 3464
rect 44899 3424 44908 3464
rect 44948 3424 44957 3464
rect 18499 3340 18508 3380
rect 18548 3340 19075 3380
rect 19115 3340 19124 3380
rect 19168 3340 19177 3380
rect 19217 3340 19508 3380
rect 19651 3340 19660 3380
rect 19700 3340 19831 3380
rect 19180 3296 19220 3340
rect 10723 3256 10732 3296
rect 10772 3256 13460 3296
rect 15667 3256 15676 3296
rect 15716 3256 16300 3296
rect 16340 3256 16349 3296
rect 18412 3256 19220 3296
rect 15235 3172 15244 3212
rect 15284 3172 15532 3212
rect 15572 3172 15581 3212
rect 17513 3172 17644 3212
rect 17684 3172 18412 3212
rect 18452 3172 18461 3212
rect 18547 3172 18556 3212
rect 18596 3172 18605 3212
rect 18556 3128 18596 3172
rect 14275 3088 14284 3128
rect 14324 3088 18596 3128
rect 4919 3004 4928 3044
rect 4968 3004 5010 3044
rect 5050 3004 5092 3044
rect 5132 3004 5174 3044
rect 5214 3004 5256 3044
rect 5296 3004 5305 3044
rect 19468 2960 19508 3340
rect 20140 3331 20180 3340
rect 20236 3340 20628 3380
rect 20668 3340 20677 3380
rect 21353 3340 21484 3380
rect 21524 3340 21533 3380
rect 21641 3340 21772 3380
rect 21812 3340 21821 3380
rect 24137 3340 24268 3380
rect 24308 3340 24317 3380
rect 24652 3340 25420 3380
rect 25460 3340 25516 3380
rect 20236 3212 20276 3340
rect 21484 3322 21524 3331
rect 24652 3296 24692 3340
rect 25516 3331 25556 3340
rect 25804 3340 26188 3380
rect 26228 3340 26237 3380
rect 26380 3340 26443 3380
rect 26483 3340 26492 3380
rect 26555 3340 26564 3380
rect 26612 3340 26743 3380
rect 27628 3340 28012 3380
rect 28052 3340 28061 3380
rect 29300 3340 30508 3380
rect 30548 3340 30557 3380
rect 30682 3340 30691 3380
rect 30731 3340 30740 3380
rect 30787 3340 30796 3380
rect 30836 3340 30967 3380
rect 31267 3340 31276 3380
rect 31316 3340 31325 3380
rect 31625 3340 31756 3380
rect 31796 3340 31805 3380
rect 32201 3340 32275 3380
rect 32315 3340 32332 3380
rect 32372 3340 32381 3380
rect 32458 3340 32467 3380
rect 32507 3340 33580 3380
rect 33620 3340 33629 3380
rect 37804 3340 42548 3380
rect 43075 3340 43084 3380
rect 43124 3340 43700 3380
rect 25804 3296 25844 3340
rect 26380 3296 26420 3340
rect 29260 3296 29300 3340
rect 31276 3296 31316 3340
rect 31756 3331 31796 3340
rect 21379 3256 21388 3296
rect 21428 3256 21437 3296
rect 21571 3256 21580 3296
rect 21620 3256 24692 3296
rect 25699 3256 25708 3296
rect 25748 3256 25844 3296
rect 25891 3256 25900 3296
rect 25940 3256 26612 3296
rect 26659 3256 26668 3296
rect 26708 3256 29300 3296
rect 30316 3256 31276 3296
rect 31316 3256 31325 3296
rect 31852 3256 33044 3296
rect 33091 3256 33100 3296
rect 33140 3256 33340 3296
rect 33380 3256 33389 3296
rect 33580 3256 37228 3296
rect 37268 3256 37277 3296
rect 21388 3212 21428 3256
rect 26572 3212 26612 3256
rect 19747 3172 19756 3212
rect 19796 3172 20276 3212
rect 20803 3172 20812 3212
rect 20852 3172 21428 3212
rect 21667 3172 21676 3212
rect 21716 3172 26476 3212
rect 26516 3172 26525 3212
rect 26572 3172 30220 3212
rect 30260 3172 30269 3212
rect 30316 3128 30356 3256
rect 31852 3212 31892 3256
rect 30451 3172 30460 3212
rect 30500 3172 31892 3212
rect 33004 3212 33044 3256
rect 33580 3212 33620 3256
rect 33004 3172 33620 3212
rect 33667 3172 33676 3212
rect 33716 3172 36844 3212
rect 36884 3172 36893 3212
rect 37018 3172 37027 3212
rect 37067 3172 37315 3212
rect 37355 3172 37603 3212
rect 37652 3172 37661 3212
rect 37804 3128 37844 3340
rect 38419 3256 38428 3296
rect 38468 3256 38860 3296
rect 38900 3256 38909 3296
rect 39571 3256 39580 3296
rect 39620 3256 41644 3296
rect 41684 3256 41693 3296
rect 41827 3256 41836 3296
rect 41876 3256 43516 3296
rect 43556 3256 43565 3296
rect 38035 3172 38044 3212
rect 38084 3172 38420 3212
rect 38921 3172 39043 3212
rect 39092 3172 39101 3212
rect 39955 3172 39964 3212
rect 40004 3172 41740 3212
rect 41780 3172 41789 3212
rect 19555 3088 19564 3128
rect 19604 3088 24172 3128
rect 24212 3088 24221 3128
rect 24451 3088 24460 3128
rect 24500 3088 30356 3128
rect 31555 3088 31564 3128
rect 31604 3088 37844 3128
rect 38380 3128 38420 3172
rect 38380 3088 39724 3128
rect 39764 3088 39773 3128
rect 20039 3004 20048 3044
rect 20088 3004 20130 3044
rect 20170 3004 20212 3044
rect 20252 3004 20294 3044
rect 20334 3004 20376 3044
rect 20416 3004 20425 3044
rect 20524 3004 25324 3044
rect 25364 3004 25373 3044
rect 25603 3004 25612 3044
rect 25652 3004 27916 3044
rect 27956 3004 27965 3044
rect 28012 3004 33004 3044
rect 33044 3004 33053 3044
rect 35159 3004 35168 3044
rect 35208 3004 35250 3044
rect 35290 3004 35332 3044
rect 35372 3004 35414 3044
rect 35454 3004 35496 3044
rect 35536 3004 35545 3044
rect 36835 3004 36844 3044
rect 36884 3004 42892 3044
rect 42932 3004 42941 3044
rect 20524 2960 20564 3004
rect 28012 2960 28052 3004
rect 43756 2960 43796 3424
rect 46278 3296 46368 3316
rect 44755 3256 44764 3296
rect 44804 3256 46368 3296
rect 46278 3236 46368 3256
rect 46278 2960 46368 2980
rect 0 2920 1420 2960
rect 1460 2920 1469 2960
rect 2860 2920 19372 2960
rect 19412 2920 19421 2960
rect 19468 2920 20564 2960
rect 21580 2920 28052 2960
rect 28483 2920 28492 2960
rect 28532 2920 43796 2960
rect 45475 2920 45484 2960
rect 45524 2920 46368 2960
rect 0 2900 90 2920
rect 21580 2876 21620 2920
rect 46278 2900 46368 2920
rect 9187 2836 9196 2876
rect 9236 2836 10060 2876
rect 10100 2836 10109 2876
rect 10915 2836 10924 2876
rect 10964 2836 11500 2876
rect 11540 2836 11549 2876
rect 13961 2836 14044 2876
rect 14084 2836 14092 2876
rect 14132 2836 14141 2876
rect 14275 2836 14284 2876
rect 14324 2836 19988 2876
rect 20179 2836 20188 2876
rect 20228 2836 20620 2876
rect 20660 2836 20669 2876
rect 21283 2836 21292 2876
rect 21332 2836 21620 2876
rect 24499 2836 24508 2876
rect 24548 2836 39148 2876
rect 39188 2836 39197 2876
rect 39619 2836 39628 2876
rect 39668 2836 44524 2876
rect 44564 2836 44573 2876
rect 45139 2836 45148 2876
rect 45188 2836 46156 2876
rect 46196 2836 46205 2876
rect 19948 2792 19988 2836
rect 7075 2752 7084 2792
rect 7124 2752 9524 2792
rect 15619 2752 15628 2792
rect 15668 2752 15916 2792
rect 15956 2752 15965 2792
rect 18316 2752 19660 2792
rect 19700 2752 19709 2792
rect 19948 2752 31804 2792
rect 31844 2752 31853 2792
rect 32140 2752 37516 2792
rect 37556 2752 37612 2792
rect 37652 2752 37804 2792
rect 37844 2752 38092 2792
rect 38132 2752 38380 2792
rect 38420 2752 38668 2792
rect 38708 2752 38717 2792
rect 39715 2752 39724 2792
rect 39764 2752 44564 2792
rect 9484 2708 9524 2752
rect 18316 2708 18356 2752
rect 7747 2668 7756 2708
rect 7796 2668 7805 2708
rect 8899 2668 8908 2708
rect 8948 2699 9079 2708
rect 8948 2668 9004 2699
rect 0 2624 90 2644
rect 7756 2624 7796 2668
rect 0 2584 3188 2624
rect 5731 2584 5740 2624
rect 5780 2584 7372 2624
rect 7412 2584 7796 2624
rect 9044 2668 9079 2699
rect 9324 2668 9388 2708
rect 9428 2668 9484 2708
rect 9524 2668 9533 2708
rect 10601 2668 10732 2708
rect 10772 2668 10781 2708
rect 15401 2668 15532 2708
rect 15572 2668 15581 2708
rect 15802 2668 15811 2708
rect 15851 2668 17300 2708
rect 17635 2668 17644 2708
rect 17684 2668 18211 2708
rect 18251 2668 18260 2708
rect 18307 2668 18316 2708
rect 18356 2668 18365 2708
rect 18569 2668 18700 2708
rect 18740 2668 18749 2708
rect 19145 2668 19276 2708
rect 19316 2668 19325 2708
rect 19625 2668 19756 2708
rect 19796 2668 19805 2708
rect 19978 2668 19987 2708
rect 20027 2668 21484 2708
rect 21524 2668 21533 2708
rect 31267 2668 31276 2708
rect 31316 2668 31700 2708
rect 31747 2668 31756 2708
rect 31796 2668 31805 2708
rect 9004 2624 9044 2659
rect 10732 2624 10772 2659
rect 17260 2624 17300 2668
rect 18316 2624 18356 2668
rect 19276 2650 19316 2659
rect 19756 2650 19796 2659
rect 31660 2624 31700 2668
rect 31756 2624 31796 2668
rect 9004 2584 10772 2624
rect 13673 2584 13804 2624
rect 13844 2584 13853 2624
rect 17260 2584 18356 2624
rect 18665 2584 18796 2624
rect 18836 2584 18845 2624
rect 20393 2584 20428 2624
rect 20468 2584 20524 2624
rect 20564 2584 20573 2624
rect 24137 2584 24268 2624
rect 24308 2584 24317 2624
rect 31145 2584 31180 2624
rect 31220 2584 31276 2624
rect 31316 2584 31325 2624
rect 31651 2584 31660 2624
rect 31700 2584 31709 2624
rect 31756 2584 32044 2624
rect 32084 2584 32093 2624
rect 0 2564 90 2584
rect 3148 2540 3188 2584
rect 32140 2540 32180 2752
rect 40003 2668 40012 2708
rect 40052 2668 43124 2708
rect 43084 2624 43124 2668
rect 44524 2624 44564 2752
rect 46278 2624 46368 2644
rect 36233 2584 36364 2624
rect 36404 2584 36413 2624
rect 39113 2584 39148 2624
rect 39188 2584 39244 2624
rect 39284 2584 39293 2624
rect 39427 2584 39436 2624
rect 39476 2584 39532 2624
rect 39572 2584 39607 2624
rect 39715 2584 39724 2624
rect 39764 2584 39895 2624
rect 40099 2584 40108 2624
rect 40148 2584 40279 2624
rect 40361 2584 40492 2624
rect 40532 2584 40876 2624
rect 40916 2584 41164 2624
rect 41204 2584 41213 2624
rect 43075 2584 43084 2624
rect 43124 2584 43133 2624
rect 43180 2584 44140 2624
rect 44180 2584 44189 2624
rect 44249 2584 44332 2624
rect 44372 2584 44380 2624
rect 44420 2584 44429 2624
rect 44515 2584 44524 2624
rect 44564 2584 44573 2624
rect 44777 2584 44908 2624
rect 44948 2584 44957 2624
rect 45772 2584 46368 2624
rect 43180 2540 43220 2584
rect 45772 2540 45812 2584
rect 46278 2564 46368 2584
rect 3148 2500 32180 2540
rect 39955 2500 39964 2540
rect 40004 2500 43220 2540
rect 43363 2500 43372 2540
rect 43412 2500 44468 2540
rect 44755 2500 44764 2540
rect 44804 2500 45812 2540
rect 7603 2416 7612 2456
rect 7652 2416 13132 2456
rect 13172 2416 13181 2456
rect 16073 2416 16204 2456
rect 16244 2416 16253 2456
rect 19180 2416 19412 2456
rect 19843 2416 19852 2456
rect 19892 2416 22388 2456
rect 27043 2416 27052 2456
rect 27092 2416 31036 2456
rect 31076 2416 31085 2456
rect 31180 2416 31420 2456
rect 31460 2416 31469 2456
rect 36595 2416 36604 2456
rect 36644 2416 39380 2456
rect 40339 2416 40348 2456
rect 40388 2416 40588 2456
rect 40628 2416 40637 2456
rect 40723 2416 40732 2456
rect 40772 2416 41972 2456
rect 42019 2416 42028 2456
rect 42068 2416 42844 2456
rect 42884 2416 42893 2456
rect 19180 2372 19220 2416
rect 3532 2332 19220 2372
rect 0 2288 90 2308
rect 3532 2288 3572 2332
rect 19372 2288 19412 2416
rect 22348 2372 22388 2416
rect 31180 2372 31220 2416
rect 22348 2332 31220 2372
rect 39340 2372 39380 2416
rect 41932 2372 41972 2416
rect 44428 2372 44468 2500
rect 39340 2332 39628 2372
rect 39668 2332 39677 2372
rect 41932 2332 44372 2372
rect 44428 2332 46292 2372
rect 0 2248 3572 2288
rect 3679 2248 3688 2288
rect 3728 2248 3770 2288
rect 3810 2248 3852 2288
rect 3892 2248 3934 2288
rect 3974 2248 4016 2288
rect 4056 2248 4065 2288
rect 8707 2248 8716 2288
rect 8756 2248 18604 2288
rect 18644 2248 18653 2288
rect 18799 2248 18808 2288
rect 18848 2248 18890 2288
rect 18930 2248 18972 2288
rect 19012 2248 19054 2288
rect 19094 2248 19136 2288
rect 19176 2248 19185 2288
rect 19372 2248 32044 2288
rect 32084 2248 32093 2288
rect 33919 2248 33928 2288
rect 33968 2248 34010 2288
rect 34050 2248 34092 2288
rect 34132 2248 34174 2288
rect 34214 2248 34256 2288
rect 34296 2248 34305 2288
rect 37900 2248 43084 2288
rect 43124 2248 43133 2288
rect 0 2228 90 2248
rect 8812 2164 11404 2204
rect 11444 2164 11453 2204
rect 16195 2164 16204 2204
rect 16244 2164 30220 2204
rect 30260 2164 30269 2204
rect 8812 2120 8852 2164
rect 4243 2080 4252 2120
rect 4292 2080 7180 2120
rect 7220 2080 7229 2120
rect 8620 2080 8852 2120
rect 9545 2080 9628 2120
rect 9668 2080 9676 2120
rect 9716 2080 9725 2120
rect 10348 2080 26860 2120
rect 26900 2080 26909 2120
rect 27628 2080 32428 2120
rect 32468 2080 32477 2120
rect 8620 2036 8660 2080
rect 2707 1996 2716 2036
rect 2756 1996 8660 2036
rect 0 1952 90 1972
rect 10348 1952 10388 2080
rect 27628 2036 27668 2080
rect 13036 1996 27668 2036
rect 27724 1996 36364 2036
rect 36404 1996 36413 2036
rect 0 1912 1268 1952
rect 2345 1912 2380 1952
rect 2420 1912 2476 1952
rect 2516 1912 2525 1952
rect 3881 1912 3916 1952
rect 3956 1912 4012 1952
rect 4052 1912 4061 1952
rect 5731 1912 5740 1952
rect 5780 1912 7220 1952
rect 7267 1912 7276 1952
rect 7316 1912 8620 1952
rect 8660 1912 8669 1952
rect 8803 1912 8812 1952
rect 8852 1912 8861 1952
rect 9257 1912 9388 1952
rect 9428 1912 9437 1952
rect 10339 1912 10348 1952
rect 10388 1912 10397 1952
rect 11753 1912 11884 1952
rect 11924 1912 11933 1952
rect 0 1892 90 1912
rect 0 1616 90 1636
rect 1228 1616 1268 1912
rect 7180 1868 7220 1912
rect 8812 1868 8852 1912
rect 13036 1868 13076 1996
rect 27724 1952 27764 1996
rect 37900 1952 37940 2248
rect 44332 2204 44372 2332
rect 46252 2308 46292 2332
rect 46252 2248 46368 2308
rect 46278 2228 46368 2248
rect 40579 2164 40588 2204
rect 40628 2164 44180 2204
rect 44332 2164 44948 2204
rect 44140 2120 44180 2164
rect 13219 1912 13228 1952
rect 13268 1912 18604 1952
rect 18644 1912 18653 1952
rect 18787 1912 18796 1952
rect 18836 1912 21196 1952
rect 21236 1912 21245 1952
rect 23107 1912 23116 1952
rect 23156 1912 27764 1952
rect 30019 1912 30028 1952
rect 30068 1912 37940 1952
rect 38284 2080 43948 2120
rect 43988 2080 43997 2120
rect 44140 2080 44276 2120
rect 7180 1828 8044 1868
rect 8084 1828 8093 1868
rect 8812 1828 13076 1868
rect 13123 1828 13132 1868
rect 13172 1828 22924 1868
rect 22964 1828 22973 1868
rect 38284 1784 38324 2080
rect 43219 1996 43228 2036
rect 43268 1996 43372 2036
rect 43412 1996 43421 2036
rect 44236 1952 44276 2080
rect 44323 1996 44332 2036
rect 44372 1996 44852 2036
rect 39084 1912 39148 1952
rect 39188 1912 39244 1952
rect 39284 1912 39724 1952
rect 39764 1912 40108 1952
rect 40148 1912 40157 1952
rect 40291 1912 40300 1952
rect 40340 1912 42988 1952
rect 43028 1912 43037 1952
rect 43180 1912 43372 1952
rect 43412 1912 43421 1952
rect 43747 1912 43756 1952
rect 43796 1912 43805 1952
rect 44131 1912 44140 1952
rect 44180 1912 44276 1952
rect 44515 1912 44524 1952
rect 44564 1912 44573 1952
rect 40108 1868 40148 1912
rect 43180 1868 43220 1912
rect 40108 1828 40300 1868
rect 40340 1828 40349 1868
rect 41635 1828 41644 1868
rect 41684 1828 43220 1868
rect 43756 1784 43796 1912
rect 44524 1868 44564 1912
rect 43843 1828 43852 1868
rect 43892 1828 44564 1868
rect 44812 1868 44852 1996
rect 44908 1952 44948 2164
rect 45139 2080 45148 2120
rect 45188 2080 45484 2120
rect 45524 2080 45533 2120
rect 46278 1952 46368 1972
rect 44899 1912 44908 1952
rect 44948 1912 44957 1952
rect 45388 1912 46368 1952
rect 45388 1868 45428 1912
rect 46278 1892 46368 1912
rect 44812 1828 45428 1868
rect 1315 1744 1324 1784
rect 1364 1744 23020 1784
rect 23060 1744 23069 1784
rect 30211 1744 30220 1784
rect 30260 1744 38324 1784
rect 41731 1744 41740 1784
rect 41780 1744 43796 1784
rect 43987 1744 43996 1784
rect 44036 1744 45676 1784
rect 45716 1744 45725 1784
rect 5369 1660 5452 1700
rect 5492 1660 5500 1700
rect 5540 1660 5549 1700
rect 6905 1660 6988 1700
rect 7028 1660 7036 1700
rect 7076 1660 7085 1700
rect 8441 1660 8524 1700
rect 8564 1660 8572 1700
rect 8612 1660 8621 1700
rect 9977 1660 10060 1700
rect 10100 1660 10108 1700
rect 10148 1660 10157 1700
rect 11513 1660 11596 1700
rect 11636 1660 11644 1700
rect 11684 1660 11693 1700
rect 16003 1660 16012 1700
rect 16052 1660 18556 1700
rect 18596 1660 18605 1700
rect 18691 1660 18700 1700
rect 18740 1660 27052 1700
rect 27092 1660 27101 1700
rect 28012 1660 39148 1700
rect 39188 1660 39197 1700
rect 39305 1660 39427 1700
rect 39476 1660 39715 1700
rect 39755 1660 40108 1700
rect 40148 1660 40579 1700
rect 40619 1660 40628 1700
rect 43603 1660 43612 1700
rect 43652 1660 44276 1700
rect 44371 1660 44380 1700
rect 44420 1660 44620 1700
rect 44660 1660 44669 1700
rect 44755 1660 44764 1700
rect 44804 1660 44813 1700
rect 28012 1616 28052 1660
rect 0 1576 460 1616
rect 500 1576 509 1616
rect 1228 1576 7220 1616
rect 14755 1576 14764 1616
rect 14804 1576 19852 1616
rect 19892 1576 19901 1616
rect 19948 1576 28052 1616
rect 32227 1576 32236 1616
rect 32276 1576 42028 1616
rect 42068 1576 42077 1616
rect 0 1556 90 1576
rect 7180 1532 7220 1576
rect 19948 1532 19988 1576
rect 44236 1532 44276 1660
rect 44764 1616 44804 1660
rect 46278 1616 46368 1636
rect 44764 1576 46368 1616
rect 46278 1556 46368 1576
rect 4919 1492 4928 1532
rect 4968 1492 5010 1532
rect 5050 1492 5092 1532
rect 5132 1492 5174 1532
rect 5214 1492 5256 1532
rect 5296 1492 5305 1532
rect 7180 1492 19988 1532
rect 20039 1492 20048 1532
rect 20088 1492 20130 1532
rect 20170 1492 20212 1532
rect 20252 1492 20294 1532
rect 20334 1492 20376 1532
rect 20416 1492 20425 1532
rect 35159 1492 35168 1532
rect 35208 1492 35250 1532
rect 35290 1492 35332 1532
rect 35372 1492 35414 1532
rect 35454 1492 35496 1532
rect 35536 1492 35545 1532
rect 38851 1492 38860 1532
rect 38900 1492 43756 1532
rect 43796 1492 43805 1532
rect 44236 1492 46196 1532
rect 46156 1448 46196 1492
rect 46156 1408 46252 1448
rect 46292 1408 46301 1448
rect 0 1280 90 1300
rect 46278 1280 46368 1300
rect 0 1240 39052 1280
rect 39092 1240 39101 1280
rect 46243 1240 46252 1280
rect 46292 1240 46368 1280
rect 0 1220 90 1240
rect 46278 1220 46368 1240
rect 0 944 90 964
rect 46278 944 46368 964
rect 0 904 39532 944
rect 39572 904 39581 944
rect 45667 904 45676 944
rect 45716 904 46368 944
rect 0 884 90 904
rect 46278 884 46368 904
rect 0 608 90 628
rect 46278 608 46368 628
rect 0 568 39436 608
rect 39476 568 39485 608
rect 44611 568 44620 608
rect 44660 568 46368 608
rect 0 548 90 568
rect 46278 548 46368 568
rect 23875 316 23884 356
rect 23924 316 41452 356
rect 41492 316 41501 356
rect 22339 232 22348 272
rect 22388 232 43660 272
rect 43700 232 43709 272
rect 19267 148 19276 188
rect 19316 148 43468 188
rect 43508 148 43517 188
rect 13123 64 13132 104
rect 13172 64 42988 104
rect 43028 64 43037 104
<< via2 >>
rect 2476 11740 2516 11780
rect 26764 11740 26804 11780
rect 2956 11656 2996 11696
rect 26956 11656 26996 11696
rect 1324 10984 1364 11024
rect 43180 10984 43220 11024
rect 1132 10648 1172 10688
rect 44044 10648 44084 10688
rect 1420 10312 1460 10352
rect 44428 10312 44468 10352
rect 19564 10228 19604 10268
rect 27244 10228 27284 10268
rect 18604 10060 18644 10100
rect 19180 10060 19220 10100
rect 24172 10060 24212 10100
rect 1324 9976 1364 10016
rect 3148 9976 3188 10016
rect 9772 9976 9812 10016
rect 15532 9976 15572 10016
rect 18412 9976 18452 10016
rect 18892 9976 18932 10016
rect 20140 9976 20180 10016
rect 25036 10060 25076 10100
rect 25900 10060 25940 10100
rect 28204 10060 28244 10100
rect 29836 10060 29876 10100
rect 42988 10060 43028 10100
rect 24556 9976 24596 10016
rect 42892 9976 42932 10016
rect 44524 9976 44564 10016
rect 7852 9892 7892 9932
rect 10060 9892 10100 9932
rect 13420 9892 13460 9932
rect 16108 9892 16148 9932
rect 16300 9892 16340 9932
rect 19564 9892 19604 9932
rect 42316 9892 42356 9932
rect 3688 9808 3728 9848
rect 3770 9808 3810 9848
rect 3852 9808 3892 9848
rect 3934 9808 3974 9848
rect 4016 9808 4056 9848
rect 18808 9808 18848 9848
rect 18890 9808 18930 9848
rect 18972 9808 19012 9848
rect 19054 9808 19094 9848
rect 19136 9808 19176 9848
rect 27244 9808 27284 9848
rect 28972 9808 29012 9848
rect 29260 9808 29300 9848
rect 33928 9808 33968 9848
rect 34010 9808 34050 9848
rect 34092 9808 34132 9848
rect 34174 9808 34214 9848
rect 34256 9808 34296 9848
rect 40492 9808 40532 9848
rect 44140 9808 44180 9848
rect 1420 9556 1460 9596
rect 1228 9472 1268 9512
rect 16300 9724 16340 9764
rect 18412 9724 18452 9764
rect 11212 9640 11252 9680
rect 11980 9640 12020 9680
rect 12748 9640 12788 9680
rect 13900 9640 13940 9680
rect 14668 9640 14708 9680
rect 15052 9640 15092 9680
rect 15436 9640 15476 9680
rect 15820 9640 15860 9680
rect 16204 9640 16244 9680
rect 16588 9640 16628 9680
rect 16972 9640 17012 9680
rect 17356 9640 17396 9680
rect 17740 9640 17780 9680
rect 18124 9640 18164 9680
rect 18508 9640 18548 9680
rect 19756 9640 19796 9680
rect 11404 9556 11444 9596
rect 12364 9556 12404 9596
rect 12940 9556 12980 9596
rect 13516 9556 13556 9596
rect 14284 9556 14324 9596
rect 14860 9556 14900 9596
rect 19372 9556 19412 9596
rect 26092 9724 26132 9764
rect 26380 9724 26420 9764
rect 26956 9724 26996 9764
rect 28876 9724 28916 9764
rect 20428 9640 20468 9680
rect 20812 9640 20852 9680
rect 24364 9640 24404 9680
rect 24652 9640 24692 9680
rect 25324 9640 25364 9680
rect 26188 9640 26228 9680
rect 27436 9640 27476 9680
rect 28492 9640 28532 9680
rect 21196 9556 21236 9596
rect 21580 9556 21620 9596
rect 21964 9556 22004 9596
rect 22156 9556 22196 9596
rect 23692 9556 23732 9596
rect 24268 9556 24308 9596
rect 24460 9556 24500 9596
rect 25420 9556 25460 9596
rect 28300 9556 28340 9596
rect 3148 9472 3188 9512
rect 10732 9472 10772 9512
rect 11116 9472 11156 9512
rect 11500 9472 11540 9512
rect 11884 9472 11924 9512
rect 12460 9472 12500 9512
rect 12652 9472 12692 9512
rect 13612 9472 13652 9512
rect 13996 9472 14036 9512
rect 14188 9472 14228 9512
rect 14572 9472 14612 9512
rect 14956 9472 14996 9512
rect 15340 9472 15380 9512
rect 16204 9472 16244 9512
rect 16492 9472 16532 9512
rect 16876 9472 16916 9512
rect 17260 9472 17300 9512
rect 17644 9472 17684 9512
rect 18028 9472 18068 9512
rect 18412 9472 18452 9512
rect 18604 9472 18644 9512
rect 19084 9472 19124 9512
rect 20140 9472 20180 9512
rect 22348 9472 22388 9512
rect 22540 9472 22580 9512
rect 23884 9472 23924 9512
rect 24076 9472 24116 9512
rect 25900 9472 25940 9512
rect 28108 9472 28148 9512
rect 6124 9304 6164 9344
rect 12844 9388 12884 9428
rect 17836 9388 17876 9428
rect 19756 9388 19796 9428
rect 19948 9388 19988 9428
rect 24556 9388 24596 9428
rect 24844 9388 24884 9428
rect 25804 9388 25844 9428
rect 26956 9388 26996 9428
rect 27340 9388 27380 9428
rect 28684 9388 28724 9428
rect 41836 9724 41876 9764
rect 31180 9640 31220 9680
rect 31564 9640 31604 9680
rect 31372 9556 31412 9596
rect 31756 9556 31796 9596
rect 33484 9640 33524 9680
rect 34732 9640 34772 9680
rect 35020 9640 35060 9680
rect 32716 9556 32756 9596
rect 35404 9556 35444 9596
rect 43084 9640 43124 9680
rect 44044 9640 44084 9680
rect 44428 9640 44468 9680
rect 40396 9556 40436 9596
rect 43564 9556 43604 9596
rect 31468 9472 31508 9512
rect 31660 9472 31700 9512
rect 32236 9472 32276 9512
rect 33100 9472 33140 9512
rect 33388 9472 33428 9512
rect 33772 9472 33812 9512
rect 34156 9472 34196 9512
rect 34732 9472 34772 9512
rect 35020 9472 35060 9512
rect 35692 9472 35732 9512
rect 38860 9472 38900 9512
rect 41644 9472 41684 9512
rect 42220 9472 42260 9512
rect 42604 9472 42644 9512
rect 10828 9304 10868 9344
rect 11788 9304 11828 9344
rect 19372 9304 19412 9344
rect 19564 9304 19604 9344
rect 23308 9304 23348 9344
rect 23692 9304 23732 9344
rect 25036 9304 25076 9344
rect 25708 9304 25748 9344
rect 26476 9304 26516 9344
rect 26860 9304 26900 9344
rect 1708 9220 1748 9260
rect 7084 9220 7124 9260
rect 10924 9220 10964 9260
rect 14284 9220 14324 9260
rect 14668 9220 14708 9260
rect 17452 9220 17492 9260
rect 20716 9220 20756 9260
rect 21196 9220 21236 9260
rect 22540 9220 22580 9260
rect 23596 9220 23636 9260
rect 24364 9220 24404 9260
rect 16204 9136 16244 9176
rect 19372 9136 19412 9176
rect 25132 9220 25172 9260
rect 26956 9220 26996 9260
rect 27148 9220 27188 9260
rect 29164 9220 29204 9260
rect 29836 9220 29876 9260
rect 24172 9136 24212 9176
rect 26380 9136 26420 9176
rect 26668 9136 26708 9176
rect 28588 9136 28628 9176
rect 31948 9304 31988 9344
rect 33388 9304 33428 9344
rect 33772 9304 33812 9344
rect 34540 9304 34580 9344
rect 32044 9220 32084 9260
rect 32332 9220 32372 9260
rect 33196 9220 33236 9260
rect 44908 9472 44948 9512
rect 37804 9388 37844 9428
rect 37708 9304 37748 9344
rect 35788 9220 35828 9260
rect 40492 9220 40532 9260
rect 41836 9220 41876 9260
rect 34540 9136 34580 9176
rect 35980 9136 36020 9176
rect 37612 9136 37652 9176
rect 37900 9136 37940 9176
rect 42220 9136 42260 9176
rect 43468 9220 43499 9260
rect 43499 9220 43508 9260
rect 4928 9052 4968 9092
rect 5010 9052 5050 9092
rect 5092 9052 5132 9092
rect 5174 9052 5214 9092
rect 5256 9052 5296 9092
rect 10060 9052 10100 9092
rect 11884 9052 11924 9092
rect 1228 8968 1268 9008
rect 12268 8968 12308 9008
rect 16684 8968 16724 9008
rect 16876 8968 16916 9008
rect 19660 8968 19700 9008
rect 20048 9052 20088 9092
rect 20130 9052 20170 9092
rect 20212 9052 20252 9092
rect 20294 9052 20334 9092
rect 20376 9052 20416 9092
rect 23116 9052 23156 9092
rect 26764 9052 26804 9092
rect 27052 9052 27092 9092
rect 35168 9052 35208 9092
rect 35250 9052 35290 9092
rect 35332 9052 35372 9092
rect 35414 9052 35454 9092
rect 35496 9052 35536 9092
rect 35596 9052 35636 9092
rect 40108 9052 40148 9092
rect 19852 8968 19892 9008
rect 20812 8968 20852 9008
rect 28396 8968 28436 9008
rect 29164 8968 29204 9008
rect 31756 8968 31796 9008
rect 42988 8968 43028 9008
rect 7852 8884 7892 8924
rect 10540 8884 10580 8924
rect 11020 8884 11060 8924
rect 11596 8884 11636 8924
rect 11884 8884 11923 8924
rect 11923 8884 11924 8924
rect 12172 8884 12212 8924
rect 12556 8884 12596 8924
rect 13036 8884 13076 8924
rect 13324 8884 13364 8924
rect 13708 8884 13748 8924
rect 14476 8884 14516 8924
rect 15244 8884 15284 8924
rect 15628 8884 15668 8924
rect 16012 8884 16052 8924
rect 16396 8884 16436 8924
rect 16780 8884 16820 8924
rect 17164 8884 17204 8924
rect 17548 8884 17588 8924
rect 17932 8884 17972 8924
rect 18316 8884 18356 8924
rect 18700 8884 18740 8924
rect 19276 8884 19316 8924
rect 19468 8884 19508 8924
rect 20044 8884 20084 8924
rect 20524 8884 20564 8924
rect 21004 8884 21044 8924
rect 21292 8884 21332 8924
rect 28684 8884 28724 8924
rect 31948 8884 31988 8924
rect 32140 8884 32180 8924
rect 32524 8884 32564 8924
rect 32908 8884 32948 8924
rect 33292 8884 33332 8924
rect 33676 8884 33716 8924
rect 34348 8884 34388 8924
rect 34828 8884 34868 8924
rect 37228 8884 37268 8924
rect 37900 8884 37940 8924
rect 44524 8884 44564 8924
rect 1132 8800 1172 8840
rect 19756 8800 19796 8840
rect 20428 8800 20468 8840
rect 20620 8800 20660 8840
rect 22828 8800 22868 8840
rect 23980 8800 24020 8840
rect 25900 8800 25940 8840
rect 28204 8800 28244 8840
rect 29740 8800 29780 8840
rect 32620 8800 32660 8840
rect 34444 8800 34484 8840
rect 34732 8800 34772 8840
rect 38380 8800 38420 8840
rect 9676 8716 9716 8756
rect 11596 8716 11636 8756
rect 652 8632 692 8672
rect 1804 8632 1844 8672
rect 2188 8632 2228 8672
rect 9004 8632 9044 8672
rect 9772 8632 9812 8672
rect 10156 8632 10196 8672
rect 11212 8632 11252 8672
rect 11980 8716 12020 8756
rect 12940 8716 12980 8756
rect 19852 8716 19892 8756
rect 21292 8716 21332 8756
rect 25996 8716 26036 8756
rect 26188 8716 26228 8756
rect 26764 8716 26804 8756
rect 27628 8716 27668 8756
rect 29836 8716 29876 8756
rect 33100 8716 33140 8756
rect 33484 8716 33524 8756
rect 34252 8716 34292 8756
rect 38668 8800 38708 8840
rect 41932 8800 41972 8840
rect 42316 8800 42356 8840
rect 42700 8800 42740 8840
rect 43084 8800 43124 8840
rect 39052 8716 39092 8756
rect 40300 8716 40340 8756
rect 42892 8716 42932 8756
rect 11404 8632 11444 8672
rect 12268 8632 12308 8672
rect 13228 8632 13268 8672
rect 14188 8632 14228 8672
rect 14380 8632 14420 8672
rect 14764 8632 14804 8672
rect 15244 8632 15284 8672
rect 15532 8632 15572 8672
rect 15916 8632 15956 8672
rect 16684 8632 16724 8672
rect 17548 8632 17588 8672
rect 17740 8632 17780 8672
rect 18220 8632 18260 8672
rect 18604 8632 18644 8672
rect 19180 8632 19220 8672
rect 19756 8632 19796 8672
rect 19948 8632 19988 8672
rect 20908 8632 20948 8672
rect 21388 8632 21428 8672
rect 21772 8632 21812 8672
rect 23308 8632 23348 8672
rect 23500 8632 23540 8672
rect 25228 8632 25268 8672
rect 25612 8632 25652 8672
rect 26668 8632 26708 8672
rect 27052 8632 27092 8672
rect 28012 8632 28052 8672
rect 29068 8632 29108 8672
rect 29452 8632 29492 8672
rect 30316 8632 30356 8672
rect 31564 8632 31604 8672
rect 11020 8548 11060 8588
rect 11980 8548 12020 8588
rect 12556 8548 12596 8588
rect 14860 8548 14900 8588
rect 43564 8716 43604 8756
rect 34732 8632 34772 8672
rect 35308 8632 35348 8672
rect 38956 8632 38996 8672
rect 41740 8632 41780 8672
rect 42988 8632 43028 8672
rect 44140 8632 44180 8672
rect 44908 8632 44948 8672
rect 17356 8548 17396 8588
rect 20140 8548 20180 8588
rect 21580 8548 21620 8588
rect 24940 8548 24980 8588
rect 25804 8548 25844 8588
rect 26764 8548 26804 8588
rect 27436 8548 27476 8588
rect 33484 8548 33524 8588
rect 34924 8548 34964 8588
rect 40780 8548 40820 8588
rect 42892 8548 42932 8588
rect 10348 8464 10388 8504
rect 12076 8464 12116 8504
rect 13900 8464 13940 8504
rect 18124 8464 18164 8504
rect 22060 8464 22100 8504
rect 25228 8464 25268 8504
rect 27340 8464 27380 8504
rect 27532 8464 27572 8504
rect 28876 8464 28916 8504
rect 33580 8464 33620 8504
rect 33772 8464 33812 8504
rect 35020 8464 35060 8504
rect 45772 8464 45812 8504
rect 12364 8380 12404 8420
rect 14572 8380 14612 8420
rect 3688 8296 3728 8336
rect 3770 8296 3810 8336
rect 3852 8296 3892 8336
rect 3934 8296 3974 8336
rect 4016 8296 4056 8336
rect 4396 8296 4436 8336
rect 11116 8296 11156 8336
rect 11308 8296 11348 8336
rect 18508 8296 18548 8336
rect 18808 8296 18848 8336
rect 18890 8296 18930 8336
rect 18972 8296 19012 8336
rect 19054 8296 19094 8336
rect 19136 8296 19176 8336
rect 22444 8296 22484 8336
rect 22636 8296 22676 8336
rect 27724 8296 27764 8336
rect 28780 8296 28820 8336
rect 30028 8296 30068 8336
rect 33928 8296 33968 8336
rect 34010 8296 34050 8336
rect 34092 8296 34132 8336
rect 34174 8296 34214 8336
rect 34256 8296 34296 8336
rect 34636 8296 34676 8336
rect 35980 8296 36020 8336
rect 38860 8296 38900 8336
rect 7852 8212 7892 8252
rect 12844 8212 12884 8252
rect 17452 8212 17492 8252
rect 26092 8212 26132 8252
rect 33580 8212 33620 8252
rect 652 7960 692 8000
rect 1228 7960 1268 8000
rect 2476 7960 2516 8000
rect 2956 7960 2996 8000
rect 12460 8128 12500 8168
rect 15148 8128 15188 8168
rect 17836 8128 17876 8168
rect 20140 8128 20180 8168
rect 22924 8128 22964 8168
rect 28204 8128 28244 8168
rect 28396 8128 28436 8168
rect 28780 8128 28820 8168
rect 33772 8128 33812 8168
rect 34540 8128 34580 8168
rect 34732 8128 34772 8168
rect 38668 8128 38708 8168
rect 4300 8044 4340 8084
rect 10444 8044 10484 8084
rect 14668 8044 14708 8084
rect 22060 8044 22100 8084
rect 25900 8044 25940 8084
rect 3244 7960 3284 8000
rect 4012 7960 4052 8000
rect 9772 7960 9812 8000
rect 10156 7960 10196 8000
rect 10540 7960 10580 8000
rect 7948 7876 7988 7916
rect 9388 7876 9428 7916
rect 10348 7876 10388 7916
rect 11308 7960 11348 8000
rect 2956 7792 2996 7832
rect 10924 7876 10964 7916
rect 11788 7876 11828 7916
rect 12076 7876 12107 7916
rect 12107 7876 12116 7916
rect 12268 7876 12308 7916
rect 14476 7960 14516 8000
rect 18124 7960 18164 8000
rect 21676 7960 21716 8000
rect 22636 7960 22676 8000
rect 26860 7960 26900 8000
rect 16108 7876 16148 7916
rect 18508 7876 18548 7916
rect 24652 7876 24692 7916
rect 26188 7876 26228 7916
rect 26476 7876 26516 7916
rect 26764 7876 26804 7916
rect 27436 7876 27476 7916
rect 11116 7792 11156 7832
rect 15340 7792 15380 7832
rect 16204 7792 16244 7832
rect 22444 7792 22484 7832
rect 26092 7792 26132 7832
rect 33580 8044 33620 8084
rect 35692 8044 35732 8084
rect 41740 8044 41780 8084
rect 42028 8044 42068 8084
rect 29068 7960 29108 8000
rect 29452 7960 29492 8000
rect 31180 7960 31220 8000
rect 33772 7960 33812 8000
rect 34252 7960 34292 8000
rect 34924 7960 34964 8000
rect 36076 7960 36116 8000
rect 44524 7960 44564 8000
rect 44908 7960 44948 8000
rect 45772 7960 45812 8000
rect 28780 7876 28820 7916
rect 33004 7876 33044 7916
rect 27916 7792 27956 7832
rect 36460 7792 36500 7832
rect 36652 7876 36692 7916
rect 43276 7876 43316 7916
rect 36748 7792 36788 7832
rect 43468 7792 43508 7832
rect 4396 7708 4436 7748
rect 11692 7708 11732 7748
rect 12364 7708 12404 7748
rect 12844 7708 12884 7748
rect 15820 7708 15860 7748
rect 17164 7708 17204 7748
rect 19660 7708 19700 7748
rect 26380 7708 26420 7748
rect 27628 7708 27668 7748
rect 33004 7708 33044 7748
rect 33196 7708 33227 7748
rect 33227 7708 33236 7748
rect 33964 7708 34004 7748
rect 35980 7708 36020 7748
rect 36268 7708 36299 7748
rect 36299 7708 36308 7748
rect 37132 7708 37172 7748
rect 42124 7708 42164 7748
rect 10732 7624 10772 7664
rect 11980 7624 12020 7664
rect 12556 7624 12596 7664
rect 18412 7624 18452 7664
rect 25708 7624 25748 7664
rect 27052 7624 27092 7664
rect 27244 7624 27284 7664
rect 4928 7540 4968 7580
rect 5010 7540 5050 7580
rect 5092 7540 5132 7580
rect 5174 7540 5214 7580
rect 5256 7540 5296 7580
rect 12172 7540 12212 7580
rect 20048 7540 20088 7580
rect 20130 7540 20170 7580
rect 20212 7540 20252 7580
rect 20294 7540 20334 7580
rect 20376 7540 20416 7580
rect 27916 7540 27956 7580
rect 31468 7624 31508 7664
rect 33292 7624 33332 7664
rect 33100 7540 33140 7580
rect 35020 7540 35060 7580
rect 35168 7540 35208 7580
rect 35250 7540 35290 7580
rect 35332 7540 35372 7580
rect 35414 7540 35454 7580
rect 35496 7540 35536 7580
rect 35596 7540 35636 7580
rect 42028 7540 42068 7580
rect 45964 7708 46004 7748
rect 7948 7456 7988 7496
rect 11500 7456 11540 7496
rect 12556 7456 12596 7496
rect 12844 7456 12884 7496
rect 28876 7456 28916 7496
rect 4012 7372 4052 7412
rect 11596 7372 11636 7412
rect 12268 7372 12308 7412
rect 13132 7372 13172 7412
rect 20140 7372 20180 7412
rect 22156 7372 22196 7412
rect 28012 7372 28052 7412
rect 28204 7372 28244 7412
rect 31468 7372 31508 7412
rect 36364 7372 36404 7412
rect 40300 7372 40340 7412
rect 1228 7288 1268 7328
rect 2956 7288 2996 7328
rect 9964 7288 10004 7328
rect 10156 7288 10196 7328
rect 10540 7288 10580 7328
rect 11884 7288 11924 7328
rect 12172 7288 12212 7328
rect 8044 7204 8084 7244
rect 10444 7204 10475 7244
rect 10475 7204 10484 7244
rect 9964 7120 10004 7160
rect 11116 7120 11156 7160
rect 11500 7120 11540 7160
rect 13036 7288 13076 7328
rect 23212 7288 23252 7328
rect 26284 7288 26324 7328
rect 27148 7288 27188 7328
rect 28396 7288 28436 7328
rect 32140 7288 32180 7328
rect 33772 7288 33812 7328
rect 38668 7288 38708 7328
rect 44908 7288 44948 7328
rect 45964 7288 46004 7328
rect 12460 7204 12491 7244
rect 12491 7204 12500 7244
rect 12940 7204 12980 7244
rect 14860 7204 14900 7244
rect 16108 7235 16148 7244
rect 16108 7204 16148 7235
rect 22636 7204 22676 7244
rect 24652 7204 24692 7244
rect 26188 7204 26228 7244
rect 27052 7204 27092 7244
rect 28780 7204 28820 7244
rect 29452 7204 29492 7244
rect 31180 7204 31220 7244
rect 33196 7204 33236 7244
rect 34252 7204 34292 7244
rect 37708 7204 37748 7244
rect 42028 7204 42068 7244
rect 11884 7120 11924 7160
rect 12748 7120 12788 7160
rect 17164 7120 17204 7160
rect 26380 7120 26420 7160
rect 28396 7120 28436 7160
rect 38092 7120 38132 7160
rect 42124 7120 42164 7160
rect 43084 7120 43124 7160
rect 43468 7120 43508 7160
rect 43660 7120 43700 7160
rect 44236 7120 44276 7160
rect 10060 7036 10100 7076
rect 11404 7036 11444 7076
rect 12460 7036 12500 7076
rect 12940 7036 12980 7076
rect 12652 6952 12692 6992
rect 13132 6952 13172 6992
rect 21676 6952 21716 6992
rect 26188 6952 26228 6992
rect 32620 6952 32660 6992
rect 36172 6952 36212 6992
rect 41836 6952 41876 6992
rect 42604 6952 42644 6992
rect 10252 6868 10292 6908
rect 11788 6868 11828 6908
rect 14476 6868 14516 6908
rect 18028 6868 18068 6908
rect 3688 6784 3728 6824
rect 3770 6784 3810 6824
rect 3852 6784 3892 6824
rect 3934 6784 3974 6824
rect 4016 6784 4056 6824
rect 9964 6784 10004 6824
rect 18808 6784 18848 6824
rect 18890 6784 18930 6824
rect 18972 6784 19012 6824
rect 19054 6784 19094 6824
rect 19136 6784 19176 6824
rect 33928 6784 33968 6824
rect 34010 6784 34050 6824
rect 34092 6784 34132 6824
rect 34174 6784 34214 6824
rect 34256 6784 34296 6824
rect 34924 6784 34964 6824
rect 41740 6784 41780 6824
rect 10060 6700 10100 6740
rect 9388 6616 9428 6656
rect 11116 6616 11156 6656
rect 12844 6616 12884 6656
rect 18220 6700 18260 6740
rect 22540 6616 22580 6656
rect 30796 6616 30836 6656
rect 42124 6616 42164 6656
rect 11884 6532 11924 6572
rect 23596 6532 23636 6572
rect 30220 6532 30260 6572
rect 42028 6532 42068 6572
rect 6124 6448 6164 6488
rect 9964 6448 10004 6488
rect 14860 6448 14900 6488
rect 17164 6448 17204 6488
rect 19852 6448 19892 6488
rect 42316 6448 42356 6488
rect 8908 6364 8948 6404
rect 9580 6364 9620 6404
rect 10060 6364 10100 6404
rect 11212 6364 11252 6404
rect 11788 6364 11819 6404
rect 11819 6364 11828 6404
rect 15820 6364 15860 6404
rect 17452 6364 17492 6404
rect 17644 6364 17684 6404
rect 21772 6364 21812 6404
rect 30988 6364 31028 6404
rect 37996 6364 38036 6404
rect 38188 6364 38228 6404
rect 10252 6280 10292 6320
rect 10444 6280 10484 6320
rect 11500 6280 11540 6320
rect 11692 6280 11732 6320
rect 25132 6280 25172 6320
rect 30412 6280 30452 6320
rect 43084 6280 43124 6320
rect 43468 6280 43508 6320
rect 45196 6280 45236 6320
rect 4928 6028 4968 6068
rect 5010 6028 5050 6068
rect 5092 6028 5132 6068
rect 5174 6028 5214 6068
rect 5256 6028 5296 6068
rect 10636 6196 10676 6236
rect 11404 6196 11444 6236
rect 16876 6196 16916 6236
rect 42316 6196 42356 6236
rect 43660 6196 43691 6236
rect 43691 6196 43700 6236
rect 17452 6112 17492 6152
rect 44236 6112 44276 6152
rect 46252 6112 46292 6152
rect 13804 6028 13844 6068
rect 14092 6028 14132 6068
rect 20048 6028 20088 6068
rect 20130 6028 20170 6068
rect 20212 6028 20252 6068
rect 20294 6028 20334 6068
rect 20376 6028 20416 6068
rect 30604 6028 30644 6068
rect 35168 6028 35208 6068
rect 35250 6028 35290 6068
rect 35332 6028 35372 6068
rect 35414 6028 35454 6068
rect 35496 6028 35536 6068
rect 34924 5944 34964 5984
rect 38188 5944 38228 5984
rect 46252 5944 46292 5984
rect 11788 5860 11828 5900
rect 12748 5860 12788 5900
rect 18604 5860 18644 5900
rect 42604 5860 42644 5900
rect 9388 5776 9428 5816
rect 9580 5776 9620 5816
rect 9772 5776 9812 5816
rect 21580 5776 21620 5816
rect 21772 5776 21812 5816
rect 41836 5776 41876 5816
rect 9964 5692 10004 5732
rect 10444 5723 10484 5732
rect 10444 5692 10484 5723
rect 10924 5723 10964 5732
rect 10924 5692 10964 5723
rect 13324 5692 13364 5732
rect 1996 5608 2036 5648
rect 10060 5608 10100 5648
rect 11404 5608 11444 5648
rect 12556 5608 12596 5648
rect 15244 5608 15284 5648
rect 43660 5608 43700 5648
rect 43948 5608 43988 5648
rect 45196 5608 45236 5648
rect 45388 5608 45428 5648
rect 24076 5524 24116 5564
rect 5740 5440 5780 5480
rect 21868 5356 21908 5396
rect 3688 5272 3728 5312
rect 3770 5272 3810 5312
rect 3852 5272 3892 5312
rect 3934 5272 3974 5312
rect 4016 5272 4056 5312
rect 18808 5272 18848 5312
rect 18890 5272 18930 5312
rect 18972 5272 19012 5312
rect 19054 5272 19094 5312
rect 19136 5272 19176 5312
rect 33928 5272 33968 5312
rect 34010 5272 34050 5312
rect 34092 5272 34132 5312
rect 34174 5272 34214 5312
rect 34256 5272 34296 5312
rect 24268 5188 24308 5228
rect 33292 5188 33332 5228
rect 42892 5188 42932 5228
rect 20908 5104 20948 5144
rect 41644 5104 41684 5144
rect 45388 5104 45428 5144
rect 1708 5020 1748 5060
rect 35980 5020 36020 5060
rect 1996 4936 2036 4976
rect 17836 4852 17876 4892
rect 32140 4852 32180 4892
rect 32908 4936 32948 4976
rect 45772 4936 45812 4976
rect 43180 4852 43220 4892
rect 43660 4852 43700 4892
rect 39148 4768 39188 4808
rect 39052 4684 39092 4724
rect 43948 4684 43979 4724
rect 43979 4684 43988 4724
rect 34348 4600 34388 4640
rect 4928 4516 4968 4556
rect 5010 4516 5050 4556
rect 5092 4516 5132 4556
rect 5174 4516 5214 4556
rect 5256 4516 5296 4556
rect 20048 4516 20088 4556
rect 20130 4516 20170 4556
rect 20212 4516 20252 4556
rect 20294 4516 20334 4556
rect 20376 4516 20416 4556
rect 33772 4516 33812 4556
rect 35168 4516 35208 4556
rect 35250 4516 35290 4556
rect 35332 4516 35372 4556
rect 35414 4516 35454 4556
rect 35496 4516 35536 4556
rect 32044 4432 32084 4472
rect 32428 4432 32468 4472
rect 32908 4432 32948 4472
rect 33388 4432 33428 4472
rect 19756 4348 19796 4388
rect 21388 4348 21428 4388
rect 33196 4348 33236 4388
rect 43948 4348 43979 4388
rect 43979 4348 43988 4388
rect 24076 4264 24116 4304
rect 26284 4264 26324 4304
rect 27052 4264 27092 4304
rect 32332 4264 32372 4304
rect 40204 4264 40244 4304
rect 45772 4264 45812 4304
rect 45964 4264 46004 4304
rect 7276 4180 7316 4220
rect 10060 4180 10100 4220
rect 19276 4211 19316 4220
rect 19276 4180 19316 4211
rect 21580 4180 21620 4220
rect 9772 4096 9812 4136
rect 11980 4096 12020 4136
rect 17932 4096 17972 4136
rect 19660 4096 19700 4136
rect 19852 4096 19892 4136
rect 21100 4096 21140 4136
rect 21484 4096 21524 4136
rect 21676 4096 21716 4136
rect 21964 4180 22004 4220
rect 25420 4211 25460 4220
rect 25420 4180 25460 4211
rect 21868 4096 21908 4136
rect 26092 4180 26132 4220
rect 30028 4180 30068 4220
rect 30508 4180 30548 4220
rect 31372 4180 31412 4220
rect 31852 4180 31892 4220
rect 32524 4180 32564 4220
rect 26188 4096 26228 4136
rect 26572 4096 26612 4136
rect 27916 4096 27956 4136
rect 31180 4096 31220 4136
rect 32140 4096 32180 4136
rect 32428 4096 32468 4136
rect 13132 4012 13172 4052
rect 26284 4012 26324 4052
rect 15628 3928 15668 3968
rect 19180 3928 19220 3968
rect 19756 3928 19796 3968
rect 21484 3928 21524 3968
rect 652 3592 692 3632
rect 1324 3256 1364 3296
rect 3688 3760 3728 3800
rect 3770 3760 3810 3800
rect 3852 3760 3892 3800
rect 3934 3760 3974 3800
rect 4016 3760 4056 3800
rect 9292 3592 9332 3632
rect 16492 3844 16532 3884
rect 33580 4180 33620 4220
rect 34348 4180 34388 4220
rect 40300 4180 40340 4220
rect 38380 4096 38420 4136
rect 38860 4096 38900 4136
rect 42988 4096 43028 4136
rect 43468 4096 43508 4136
rect 43756 4096 43796 4136
rect 27436 4012 27476 4052
rect 28588 4012 28628 4052
rect 29740 4012 29780 4052
rect 32908 4012 32948 4052
rect 33484 4012 33524 4052
rect 41452 4012 41492 4052
rect 21772 3928 21812 3968
rect 26572 3928 26612 3968
rect 31660 3928 31700 3968
rect 32428 3928 32468 3968
rect 34252 3928 34292 3968
rect 38668 3928 38708 3968
rect 40300 3928 40340 3968
rect 43180 3928 43220 3968
rect 33196 3844 33236 3884
rect 42988 3844 43028 3884
rect 18808 3760 18848 3800
rect 18890 3760 18930 3800
rect 18972 3760 19012 3800
rect 19054 3760 19094 3800
rect 19136 3760 19176 3800
rect 19660 3760 19700 3800
rect 25036 3760 25076 3800
rect 25516 3760 25556 3800
rect 33004 3760 33044 3800
rect 33928 3760 33968 3800
rect 34010 3760 34050 3800
rect 34092 3760 34132 3800
rect 34174 3760 34214 3800
rect 34256 3760 34296 3800
rect 38956 3760 38996 3800
rect 17740 3676 17780 3716
rect 21388 3676 21428 3716
rect 21580 3676 21620 3716
rect 25804 3676 25844 3716
rect 31852 3676 31892 3716
rect 32524 3676 32564 3716
rect 32908 3676 32948 3716
rect 43084 3676 43124 3716
rect 9676 3592 9716 3632
rect 10924 3592 10964 3632
rect 13132 3592 13172 3632
rect 13324 3592 13364 3632
rect 13996 3592 14036 3632
rect 17260 3592 17300 3632
rect 19276 3592 19316 3632
rect 21676 3592 21716 3632
rect 23308 3592 23348 3632
rect 25612 3592 25652 3632
rect 26188 3592 26228 3632
rect 15052 3508 15092 3548
rect 18796 3508 18836 3548
rect 21580 3508 21620 3548
rect 25036 3508 25076 3548
rect 25228 3508 25268 3548
rect 26668 3508 26708 3548
rect 28684 3508 28724 3548
rect 31372 3508 31412 3548
rect 32812 3508 32852 3548
rect 38572 3592 38612 3632
rect 34444 3508 34484 3548
rect 41740 3508 41780 3548
rect 41932 3508 41972 3548
rect 9004 3424 9044 3464
rect 11596 3424 11636 3464
rect 15436 3424 15476 3464
rect 16204 3424 16244 3464
rect 18220 3424 18260 3464
rect 19372 3424 19412 3464
rect 19852 3424 19892 3464
rect 20524 3424 20564 3464
rect 21388 3424 21428 3464
rect 21964 3424 22004 3464
rect 22828 3424 22868 3464
rect 27628 3424 27668 3464
rect 30028 3424 30068 3464
rect 30892 3424 30932 3464
rect 31180 3424 31220 3464
rect 31852 3424 31892 3464
rect 38188 3424 38228 3464
rect 39532 3424 39572 3464
rect 40108 3424 40148 3464
rect 42988 3424 43028 3464
rect 43372 3424 43412 3464
rect 13804 3340 13844 3380
rect 15052 3340 15092 3380
rect 45964 3592 46004 3632
rect 46156 3592 46196 3632
rect 44524 3424 44564 3464
rect 18508 3340 18548 3380
rect 19660 3340 19700 3380
rect 10732 3256 10772 3296
rect 16300 3256 16340 3296
rect 15532 3172 15572 3212
rect 17644 3172 17684 3212
rect 18412 3172 18452 3212
rect 14284 3088 14324 3128
rect 4928 3004 4968 3044
rect 5010 3004 5050 3044
rect 5092 3004 5132 3044
rect 5174 3004 5214 3044
rect 5256 3004 5296 3044
rect 21484 3371 21524 3380
rect 21484 3340 21524 3371
rect 21772 3340 21812 3380
rect 24268 3340 24308 3380
rect 25420 3340 25460 3380
rect 26572 3340 26604 3380
rect 26604 3340 26612 3380
rect 30508 3340 30548 3380
rect 30796 3340 30836 3380
rect 31756 3340 31796 3380
rect 32332 3340 32372 3380
rect 33580 3340 33620 3380
rect 43084 3340 43124 3380
rect 21580 3256 21620 3296
rect 25900 3256 25940 3296
rect 26668 3256 26708 3296
rect 31276 3256 31316 3296
rect 33100 3256 33140 3296
rect 37228 3256 37268 3296
rect 19756 3172 19796 3212
rect 21676 3172 21716 3212
rect 26476 3172 26516 3212
rect 30220 3172 30260 3212
rect 33676 3172 33716 3212
rect 36844 3172 36884 3212
rect 37612 3172 37643 3212
rect 37643 3172 37652 3212
rect 38860 3256 38900 3296
rect 41644 3256 41684 3296
rect 41836 3256 41876 3296
rect 39052 3172 39083 3212
rect 39083 3172 39092 3212
rect 41740 3172 41780 3212
rect 19564 3088 19604 3128
rect 24172 3088 24212 3128
rect 24460 3088 24500 3128
rect 31564 3088 31604 3128
rect 39724 3088 39764 3128
rect 20048 3004 20088 3044
rect 20130 3004 20170 3044
rect 20212 3004 20252 3044
rect 20294 3004 20334 3044
rect 20376 3004 20416 3044
rect 25324 3004 25364 3044
rect 25612 3004 25652 3044
rect 27916 3004 27956 3044
rect 33004 3004 33044 3044
rect 35168 3004 35208 3044
rect 35250 3004 35290 3044
rect 35332 3004 35372 3044
rect 35414 3004 35454 3044
rect 35496 3004 35536 3044
rect 36844 3004 36884 3044
rect 42892 3004 42932 3044
rect 1420 2920 1460 2960
rect 19372 2920 19412 2960
rect 28492 2920 28532 2960
rect 45484 2920 45524 2960
rect 10060 2836 10100 2876
rect 11500 2836 11540 2876
rect 14092 2836 14132 2876
rect 14284 2836 14324 2876
rect 20620 2836 20660 2876
rect 21292 2836 21332 2876
rect 39148 2836 39188 2876
rect 39628 2836 39668 2876
rect 44524 2836 44564 2876
rect 46156 2836 46196 2876
rect 7084 2752 7124 2792
rect 15628 2752 15668 2792
rect 19660 2752 19700 2792
rect 37612 2752 37652 2792
rect 39724 2752 39764 2792
rect 8908 2668 8948 2708
rect 5740 2584 5780 2624
rect 9388 2668 9428 2708
rect 10732 2699 10772 2708
rect 10732 2668 10772 2699
rect 15532 2668 15572 2708
rect 17644 2668 17684 2708
rect 18700 2668 18740 2708
rect 19276 2699 19316 2708
rect 19276 2668 19316 2699
rect 19756 2699 19796 2708
rect 19756 2668 19796 2699
rect 21484 2668 21524 2708
rect 31276 2668 31316 2708
rect 31756 2668 31796 2708
rect 13804 2584 13844 2624
rect 18796 2584 18836 2624
rect 20524 2584 20564 2624
rect 24268 2584 24308 2624
rect 31180 2584 31220 2624
rect 40012 2668 40052 2708
rect 36364 2584 36404 2624
rect 39148 2584 39188 2624
rect 39436 2584 39476 2624
rect 39724 2584 39764 2624
rect 40108 2584 40148 2624
rect 40492 2584 40532 2624
rect 44332 2584 44372 2624
rect 44908 2584 44948 2624
rect 43372 2500 43412 2540
rect 13132 2416 13172 2456
rect 16204 2416 16244 2456
rect 19852 2416 19892 2456
rect 27052 2416 27092 2456
rect 40588 2416 40628 2456
rect 42028 2416 42068 2456
rect 39628 2332 39668 2372
rect 3688 2248 3728 2288
rect 3770 2248 3810 2288
rect 3852 2248 3892 2288
rect 3934 2248 3974 2288
rect 4016 2248 4056 2288
rect 8716 2248 8756 2288
rect 18604 2248 18644 2288
rect 18808 2248 18848 2288
rect 18890 2248 18930 2288
rect 18972 2248 19012 2288
rect 19054 2248 19094 2288
rect 19136 2248 19176 2288
rect 32044 2248 32084 2288
rect 33928 2248 33968 2288
rect 34010 2248 34050 2288
rect 34092 2248 34132 2288
rect 34174 2248 34214 2288
rect 34256 2248 34296 2288
rect 43084 2248 43124 2288
rect 11404 2164 11444 2204
rect 16204 2164 16244 2204
rect 30220 2164 30260 2204
rect 7180 2080 7220 2120
rect 9676 2080 9716 2120
rect 26860 2080 26900 2120
rect 32428 2080 32468 2120
rect 36364 1996 36404 2036
rect 2380 1912 2420 1952
rect 3916 1912 3956 1952
rect 8620 1912 8660 1952
rect 9388 1912 9428 1952
rect 11884 1912 11924 1952
rect 40588 2164 40628 2204
rect 13228 1912 13268 1952
rect 18604 1912 18644 1952
rect 18796 1912 18836 1952
rect 21196 1912 21236 1952
rect 23116 1912 23156 1952
rect 30028 1912 30068 1952
rect 43948 2080 43988 2120
rect 8044 1828 8084 1868
rect 13132 1828 13172 1868
rect 22924 1828 22964 1868
rect 43372 1996 43412 2036
rect 44332 1996 44372 2036
rect 39148 1912 39188 1952
rect 39724 1912 39764 1952
rect 40300 1912 40340 1952
rect 41644 1828 41684 1868
rect 43852 1828 43892 1868
rect 45484 2080 45524 2120
rect 1324 1744 1364 1784
rect 23020 1744 23060 1784
rect 30220 1744 30260 1784
rect 41740 1744 41780 1784
rect 45676 1744 45716 1784
rect 5452 1660 5492 1700
rect 6988 1660 7028 1700
rect 8524 1660 8564 1700
rect 10060 1660 10100 1700
rect 11596 1660 11636 1700
rect 16012 1660 16052 1700
rect 18700 1660 18740 1700
rect 27052 1660 27092 1700
rect 39436 1660 39467 1700
rect 39467 1660 39476 1700
rect 40108 1660 40148 1700
rect 44620 1660 44660 1700
rect 460 1576 500 1616
rect 14764 1576 14804 1616
rect 19852 1576 19892 1616
rect 32236 1576 32276 1616
rect 42028 1576 42068 1616
rect 4928 1492 4968 1532
rect 5010 1492 5050 1532
rect 5092 1492 5132 1532
rect 5174 1492 5214 1532
rect 5256 1492 5296 1532
rect 20048 1492 20088 1532
rect 20130 1492 20170 1532
rect 20212 1492 20252 1532
rect 20294 1492 20334 1532
rect 20376 1492 20416 1532
rect 35168 1492 35208 1532
rect 35250 1492 35290 1532
rect 35332 1492 35372 1532
rect 35414 1492 35454 1532
rect 35496 1492 35536 1532
rect 38860 1492 38900 1532
rect 43756 1492 43796 1532
rect 46252 1408 46292 1448
rect 39052 1240 39092 1280
rect 46252 1240 46292 1280
rect 39532 904 39572 944
rect 45676 904 45716 944
rect 39436 568 39476 608
rect 44620 568 44660 608
rect 23884 316 23924 356
rect 41452 316 41492 356
rect 22348 232 22388 272
rect 43660 232 43700 272
rect 19276 148 19316 188
rect 43468 148 43508 188
rect 13132 64 13172 104
rect 42988 64 43028 104
<< metal3 >>
rect 2476 11780 2516 11789
rect 1324 11024 1364 11033
rect 1132 10688 1172 10697
rect 1132 8840 1172 10648
rect 1324 10016 1364 10984
rect 1324 9967 1364 9976
rect 1420 10352 1460 10361
rect 1420 9596 1460 10312
rect 1420 9547 1460 9556
rect 1228 9512 1268 9521
rect 1228 9008 1268 9472
rect 1228 8959 1268 8968
rect 1708 9260 1748 9269
rect 1132 8791 1172 8800
rect 652 8672 692 8681
rect 652 8000 692 8632
rect 652 7951 692 7960
rect 1228 8000 1268 8009
rect 1228 7328 1268 7960
rect 1228 7279 1268 7288
rect 1708 5060 1748 9220
rect 1708 5011 1748 5020
rect 1804 8672 1844 8681
rect 652 3632 692 3641
rect 652 3497 692 3592
rect 460 3464 500 3473
rect 460 1616 500 3424
rect 1804 3380 1844 8632
rect 2188 8672 2228 8681
rect 1996 5648 2036 5657
rect 1996 4976 2036 5608
rect 1996 4927 2036 4936
rect 2188 4220 2228 8632
rect 2476 8000 2516 11740
rect 4300 11780 4340 11789
rect 11000 11764 11080 11844
rect 11192 11764 11272 11844
rect 11384 11764 11464 11844
rect 11576 11764 11656 11844
rect 11768 11764 11848 11844
rect 11960 11764 12040 11844
rect 12152 11764 12232 11844
rect 12344 11764 12424 11844
rect 12536 11764 12616 11844
rect 12728 11764 12808 11844
rect 12920 11764 13000 11844
rect 13112 11764 13192 11844
rect 13304 11764 13384 11844
rect 13496 11764 13576 11844
rect 13688 11764 13768 11844
rect 13880 11764 13960 11844
rect 14072 11764 14152 11844
rect 14264 11764 14344 11844
rect 14456 11764 14536 11844
rect 14648 11764 14728 11844
rect 14840 11764 14920 11844
rect 15032 11764 15112 11844
rect 15224 11764 15304 11844
rect 15416 11764 15496 11844
rect 15608 11764 15688 11844
rect 15800 11764 15880 11844
rect 15992 11764 16072 11844
rect 16184 11764 16264 11844
rect 16376 11764 16456 11844
rect 16568 11764 16648 11844
rect 16760 11764 16840 11844
rect 16952 11764 17032 11844
rect 17144 11764 17224 11844
rect 17336 11764 17416 11844
rect 17528 11764 17608 11844
rect 17720 11764 17800 11844
rect 17912 11764 17992 11844
rect 18104 11764 18184 11844
rect 18296 11764 18376 11844
rect 18488 11764 18568 11844
rect 18680 11764 18760 11844
rect 18872 11764 18952 11844
rect 19064 11764 19144 11844
rect 19256 11764 19336 11844
rect 19448 11764 19528 11844
rect 19640 11764 19720 11844
rect 19832 11764 19912 11844
rect 20024 11764 20104 11844
rect 20216 11764 20296 11844
rect 20408 11764 20488 11844
rect 20600 11764 20680 11844
rect 20792 11764 20872 11844
rect 20984 11764 21064 11844
rect 21176 11764 21256 11844
rect 21368 11764 21448 11844
rect 21560 11764 21640 11844
rect 21752 11764 21832 11844
rect 21944 11764 22024 11844
rect 22136 11764 22216 11844
rect 22328 11764 22408 11844
rect 22520 11764 22600 11844
rect 22712 11764 22792 11844
rect 22904 11764 22984 11844
rect 23096 11764 23176 11844
rect 23288 11780 23368 11844
rect 23288 11764 23308 11780
rect 2476 7951 2516 7960
rect 2956 11696 2996 11705
rect 2956 8000 2996 11656
rect 3148 10016 3188 10025
rect 3148 9512 3188 9976
rect 3688 9848 4056 9857
rect 3728 9808 3770 9848
rect 3810 9808 3852 9848
rect 3892 9808 3934 9848
rect 3974 9808 4016 9848
rect 3688 9799 4056 9808
rect 3148 9463 3188 9472
rect 3688 8336 4056 8345
rect 3728 8296 3770 8336
rect 3810 8296 3852 8336
rect 3892 8296 3934 8336
rect 3974 8296 4016 8336
rect 3688 8287 4056 8296
rect 2956 7951 2996 7960
rect 3244 8252 3284 8261
rect 3244 8000 3284 8212
rect 4300 8084 4340 11740
rect 9772 10016 9812 10025
rect 7852 9932 7892 9941
rect 6124 9344 6164 9353
rect 4928 9092 5296 9101
rect 4968 9052 5010 9092
rect 5050 9052 5092 9092
rect 5132 9052 5174 9092
rect 5214 9052 5256 9092
rect 4928 9043 5296 9052
rect 4300 8035 4340 8044
rect 4396 8336 4436 8345
rect 3244 7951 3284 7960
rect 4012 8000 4052 8009
rect 2956 7832 2996 7841
rect 2956 7328 2996 7792
rect 4012 7412 4052 7960
rect 4396 7748 4436 8296
rect 4396 7699 4436 7708
rect 4928 7580 5296 7589
rect 4968 7540 5010 7580
rect 5050 7540 5092 7580
rect 5132 7540 5174 7580
rect 5214 7540 5256 7580
rect 4928 7531 5296 7540
rect 4012 7363 4052 7372
rect 2956 7279 2996 7288
rect 3688 6824 4056 6833
rect 3728 6784 3770 6824
rect 3810 6784 3852 6824
rect 3892 6784 3934 6824
rect 3974 6784 4016 6824
rect 3688 6775 4056 6784
rect 6124 6488 6164 9304
rect 6124 6439 6164 6448
rect 7084 9260 7124 9269
rect 4928 6068 5296 6077
rect 4968 6028 5010 6068
rect 5050 6028 5092 6068
rect 5132 6028 5174 6068
rect 5214 6028 5256 6068
rect 4928 6019 5296 6028
rect 5740 5480 5780 5489
rect 3688 5312 4056 5321
rect 3728 5272 3770 5312
rect 3810 5272 3852 5312
rect 3892 5272 3934 5312
rect 3974 5272 4016 5312
rect 3688 5263 4056 5272
rect 4928 4556 5296 4565
rect 4968 4516 5010 4556
rect 5050 4516 5092 4556
rect 5132 4516 5174 4556
rect 5214 4516 5256 4556
rect 4928 4507 5296 4516
rect 2188 4171 2228 4180
rect 3688 3800 4056 3809
rect 3728 3760 3770 3800
rect 3810 3760 3852 3800
rect 3892 3760 3934 3800
rect 3974 3760 4016 3800
rect 3688 3751 4056 3760
rect 1804 3331 1844 3340
rect 1324 3296 1364 3305
rect 1324 1784 1364 3256
rect 4928 3044 5296 3053
rect 4968 3004 5010 3044
rect 5050 3004 5092 3044
rect 5132 3004 5174 3044
rect 5214 3004 5256 3044
rect 4928 2995 5296 3004
rect 1420 2960 1460 2969
rect 1420 2624 1460 2920
rect 1420 2575 1460 2584
rect 5740 2624 5780 5440
rect 7084 2792 7124 9220
rect 7852 8924 7892 9892
rect 7852 8875 7892 8884
rect 9292 9260 9332 9269
rect 9004 8672 9044 8681
rect 7852 8252 7892 8261
rect 7852 8117 7892 8212
rect 7948 7916 7988 7925
rect 7948 7496 7988 7876
rect 7948 7447 7988 7456
rect 8044 7244 8084 7253
rect 7084 2743 7124 2752
rect 7276 4220 7316 4229
rect 5740 2575 5780 2584
rect 3688 2288 4056 2297
rect 3728 2248 3770 2288
rect 3810 2248 3852 2288
rect 3892 2248 3934 2288
rect 3974 2248 4016 2288
rect 3688 2239 4056 2248
rect 7180 2120 7220 2129
rect 7276 2120 7316 4180
rect 7220 2080 7316 2120
rect 7180 2071 7220 2080
rect 1324 1735 1364 1744
rect 2380 1952 2420 1961
rect 460 1567 500 1576
rect 2380 80 2420 1912
rect 3916 1952 3956 1961
rect 3916 80 3956 1912
rect 8044 1868 8084 7204
rect 8908 6404 8948 6413
rect 8908 2708 8948 6364
rect 9004 3464 9044 8632
rect 9292 3632 9332 9220
rect 9676 8756 9716 8765
rect 9388 7916 9428 7925
rect 9388 6656 9428 7876
rect 9388 5816 9428 6616
rect 9388 5767 9428 5776
rect 9580 6404 9620 6413
rect 9580 5816 9620 6364
rect 9580 5767 9620 5776
rect 9292 3583 9332 3592
rect 9676 3632 9716 8716
rect 9772 8672 9812 9976
rect 10060 9932 10100 9941
rect 10060 9797 10100 9892
rect 10156 9764 10196 9773
rect 9772 8000 9812 8632
rect 9772 7951 9812 7960
rect 9868 9176 9908 9185
rect 9772 5816 9812 5825
rect 9772 4136 9812 5776
rect 9772 4087 9812 4096
rect 9676 3583 9716 3592
rect 9004 3415 9044 3424
rect 9868 2900 9908 9136
rect 10060 9092 10100 9101
rect 9964 7328 10004 7423
rect 9964 7279 10004 7288
rect 9964 7160 10004 7169
rect 9964 6824 10004 7120
rect 10060 7076 10100 9052
rect 10156 8672 10196 9724
rect 10732 9512 10772 9521
rect 10540 8924 10580 8933
rect 10540 8756 10580 8884
rect 10540 8707 10580 8716
rect 10156 8000 10196 8632
rect 10156 7951 10196 7960
rect 10348 8504 10388 8513
rect 10348 7916 10388 8464
rect 10348 7867 10388 7876
rect 10444 8084 10484 8093
rect 10060 7027 10100 7036
rect 10156 7328 10196 7337
rect 10156 6908 10196 7288
rect 10444 7244 10484 8044
rect 10540 8000 10580 8009
rect 10540 7328 10580 7960
rect 10732 7664 10772 9472
rect 10732 7615 10772 7624
rect 10828 9344 10868 9353
rect 10540 7279 10580 7288
rect 10444 7195 10484 7204
rect 10252 6908 10292 6917
rect 10156 6868 10252 6908
rect 9964 6488 10004 6784
rect 9964 5732 10004 6448
rect 9964 5683 10004 5692
rect 10060 6740 10100 6749
rect 10060 6404 10100 6700
rect 10060 5648 10100 6364
rect 10252 6320 10292 6868
rect 10252 6271 10292 6280
rect 10444 6320 10484 6329
rect 10444 5732 10484 6280
rect 10636 6236 10676 6245
rect 10636 6101 10676 6196
rect 10444 5683 10484 5692
rect 10060 5599 10100 5608
rect 10828 5060 10868 9304
rect 10924 9260 10964 9269
rect 10924 8168 10964 9220
rect 11020 8924 11060 11764
rect 11212 9680 11252 11764
rect 11212 9631 11252 9640
rect 11404 9596 11444 11764
rect 11404 9547 11444 9556
rect 11020 8875 11060 8884
rect 11116 9512 11156 9521
rect 11020 8588 11060 8597
rect 11020 8453 11060 8548
rect 11116 8336 11156 9472
rect 11500 9512 11540 9521
rect 11212 8672 11252 8681
rect 11212 8537 11252 8632
rect 11404 8672 11444 8681
rect 11116 8287 11156 8296
rect 11308 8336 11348 8345
rect 11308 8168 11348 8296
rect 10924 8128 11348 8168
rect 11308 8000 11348 8009
rect 10828 5011 10868 5020
rect 10924 7916 10964 7925
rect 10924 5732 10964 7876
rect 11116 7832 11156 7841
rect 11116 7160 11156 7792
rect 11116 7111 11156 7120
rect 11212 7664 11252 7673
rect 11116 6656 11156 6665
rect 11116 6404 11156 6616
rect 11116 6355 11156 6364
rect 11212 6404 11252 7624
rect 11212 6355 11252 6364
rect 9676 2860 9908 2900
rect 10060 4220 10100 4229
rect 10060 2876 10100 4180
rect 10924 3632 10964 5692
rect 10924 3583 10964 3592
rect 8908 2659 8948 2668
rect 9388 2708 9428 2717
rect 8716 2288 8756 2297
rect 8620 2248 8716 2288
rect 8620 1952 8660 2248
rect 8716 2239 8756 2248
rect 8620 1903 8660 1912
rect 9388 1952 9428 2668
rect 9676 2120 9716 2860
rect 10060 2827 10100 2836
rect 10732 3296 10772 3305
rect 10732 2708 10772 3256
rect 11308 2900 11348 7960
rect 11404 7076 11444 8632
rect 11500 7496 11540 9472
rect 11596 8924 11636 11764
rect 11788 9344 11828 11764
rect 11884 10016 11924 10025
rect 11884 9512 11924 9976
rect 11980 9680 12020 11764
rect 11980 9631 12020 9640
rect 11884 9463 11924 9472
rect 11788 9295 11828 9304
rect 11884 9092 11924 9101
rect 11924 9052 12020 9092
rect 11884 9043 11924 9052
rect 11596 8875 11636 8884
rect 11884 8924 11924 8933
rect 11596 8756 11636 8765
rect 11596 7664 11636 8716
rect 11788 7916 11828 7925
rect 11596 7615 11636 7624
rect 11692 7748 11732 7757
rect 11500 7447 11540 7456
rect 11596 7496 11636 7505
rect 11596 7412 11636 7456
rect 11596 7361 11636 7372
rect 11404 7027 11444 7036
rect 11500 7160 11540 7169
rect 11500 7025 11540 7120
rect 11596 6404 11636 6413
rect 11500 6320 11540 6329
rect 11404 6236 11444 6245
rect 11404 5648 11444 6196
rect 11404 5599 11444 5608
rect 11308 2860 11444 2900
rect 10732 2659 10772 2668
rect 11404 2204 11444 2860
rect 11500 2876 11540 6280
rect 11596 3464 11636 6364
rect 11692 6320 11732 7708
rect 11788 6992 11828 7876
rect 11884 7328 11924 8884
rect 11980 8756 12020 9052
rect 12172 8924 12212 11764
rect 12364 9596 12404 11764
rect 12364 9547 12404 9556
rect 12460 9512 12500 9521
rect 12460 9377 12500 9472
rect 12172 8875 12212 8884
rect 12268 9008 12308 9017
rect 11980 8707 12020 8716
rect 12076 8840 12116 8849
rect 11980 8588 12020 8597
rect 11980 7664 12020 8548
rect 12076 8504 12116 8800
rect 12268 8672 12308 8968
rect 12556 8924 12596 11764
rect 12748 9680 12788 11764
rect 12940 11444 12980 11764
rect 12940 11404 13076 11444
rect 12748 9631 12788 9640
rect 12844 9848 12884 9857
rect 12556 8875 12596 8884
rect 12652 9512 12692 9521
rect 12268 8623 12308 8632
rect 12556 8588 12596 8597
rect 12076 7916 12116 8464
rect 12364 8548 12556 8588
rect 12364 8420 12404 8548
rect 12556 8539 12596 8548
rect 12364 8371 12404 8380
rect 12460 8168 12500 8177
rect 12076 7867 12116 7876
rect 12268 7916 12308 7925
rect 11980 7615 12020 7624
rect 12172 7580 12212 7589
rect 12172 7445 12212 7540
rect 12268 7412 12308 7876
rect 12268 7363 12308 7372
rect 12364 7748 12404 7757
rect 11884 7279 11924 7288
rect 11980 7328 12020 7337
rect 11788 6908 11828 6952
rect 11788 6828 11828 6868
rect 11884 7160 11924 7169
rect 11884 6908 11924 7120
rect 11884 6859 11924 6868
rect 11884 6572 11924 6581
rect 11692 6271 11732 6280
rect 11788 6404 11828 6413
rect 11788 5900 11828 6364
rect 11788 5851 11828 5860
rect 11596 3415 11636 3424
rect 11500 2827 11540 2836
rect 11404 2155 11444 2164
rect 9676 2071 9716 2080
rect 9388 1903 9428 1912
rect 11884 1952 11924 6532
rect 11980 4136 12020 7288
rect 12172 7328 12212 7339
rect 12172 7244 12212 7288
rect 12364 7244 12404 7708
rect 12460 7412 12500 8128
rect 12556 7664 12596 7673
rect 12556 7496 12596 7624
rect 12556 7447 12596 7456
rect 12460 7363 12500 7372
rect 12556 7328 12596 7337
rect 12460 7244 12500 7253
rect 12364 7204 12460 7244
rect 12172 7195 12212 7204
rect 12460 7195 12500 7204
rect 12460 7076 12500 7085
rect 12460 6941 12500 7036
rect 12556 5648 12596 7288
rect 12652 6992 12692 9472
rect 12844 9428 12884 9808
rect 12940 9596 12980 9605
rect 12940 9461 12980 9556
rect 12844 9379 12884 9388
rect 13036 8924 13076 11404
rect 13132 9596 13172 11764
rect 13132 9547 13172 9556
rect 13036 8875 13076 8884
rect 13324 8924 13364 11764
rect 13420 9932 13460 9941
rect 13420 9512 13460 9892
rect 13516 9596 13556 11764
rect 13516 9547 13556 9556
rect 13420 9463 13460 9472
rect 13612 9512 13652 9521
rect 13612 9377 13652 9472
rect 13324 8875 13364 8884
rect 13708 8924 13748 11764
rect 13900 9680 13940 11764
rect 13900 9631 13940 9640
rect 13996 9512 14036 9521
rect 13708 8875 13748 8884
rect 13900 9092 13940 9101
rect 12940 8756 12980 8765
rect 12748 8716 12940 8756
rect 12748 7328 12788 8716
rect 12940 8707 12980 8716
rect 13228 8672 13268 8681
rect 12844 8252 12884 8261
rect 12844 8117 12884 8212
rect 12844 7748 12884 7757
rect 12844 7496 12884 7708
rect 12844 7447 12884 7456
rect 13036 7496 13076 7505
rect 12748 7279 12788 7288
rect 13036 7328 13076 7456
rect 13036 7279 13076 7288
rect 13132 7412 13172 7421
rect 12940 7244 12980 7253
rect 12844 7204 12940 7244
rect 12652 6943 12692 6952
rect 12748 7160 12788 7169
rect 12748 6908 12788 7120
rect 12748 5900 12788 6868
rect 12844 6656 12884 7204
rect 12940 7195 12980 7204
rect 13132 7244 13172 7372
rect 13132 7195 13172 7204
rect 12940 7076 12980 7085
rect 12940 6941 12980 7036
rect 13132 6992 13172 7001
rect 13132 6857 13172 6952
rect 12844 6607 12884 6616
rect 12748 5851 12788 5860
rect 12556 5599 12596 5608
rect 11980 4087 12020 4096
rect 13132 4052 13172 4061
rect 13132 3632 13172 4012
rect 13132 3583 13172 3592
rect 11884 1903 11924 1912
rect 13132 2456 13172 2465
rect 8044 1819 8084 1828
rect 13132 1868 13172 2416
rect 13228 1952 13268 8632
rect 13900 8504 13940 9052
rect 13900 8455 13940 8464
rect 13804 6068 13844 6077
rect 13324 5732 13364 5741
rect 13324 3632 13364 5692
rect 13324 3583 13364 3592
rect 13804 3380 13844 6028
rect 13996 3632 14036 9472
rect 14092 9092 14132 11764
rect 14284 9596 14324 11764
rect 14284 9547 14324 9556
rect 14092 9043 14132 9052
rect 14188 9512 14228 9521
rect 14188 8924 14228 9472
rect 14092 8884 14228 8924
rect 14284 9260 14324 9269
rect 14092 7748 14132 8884
rect 14092 7699 14132 7708
rect 14188 8672 14228 8681
rect 13996 3583 14036 3592
rect 14092 6068 14132 6077
rect 13804 2624 13844 3340
rect 14092 2876 14132 6028
rect 14188 2900 14228 8632
rect 14284 3128 14324 9220
rect 14476 8924 14516 11764
rect 14668 9680 14708 11764
rect 14668 9631 14708 9640
rect 14860 9596 14900 11764
rect 14860 9547 14900 9556
rect 14956 9680 14996 9689
rect 14476 8875 14516 8884
rect 14572 9512 14612 9521
rect 14380 8672 14420 8681
rect 14380 6236 14420 8632
rect 14572 8420 14612 9472
rect 14668 9512 14708 9521
rect 14668 9260 14708 9472
rect 14956 9512 14996 9640
rect 15052 9680 15092 11764
rect 15052 9631 15092 9640
rect 15148 9848 15188 9857
rect 14956 9463 14996 9472
rect 14668 9211 14708 9220
rect 14572 8371 14612 8380
rect 14764 8672 14804 8681
rect 14668 8084 14708 8093
rect 14476 8000 14516 8009
rect 14476 6908 14516 7960
rect 14476 6859 14516 6868
rect 14380 6187 14420 6196
rect 14284 3079 14324 3088
rect 14188 2876 14324 2900
rect 14188 2860 14284 2876
rect 14092 2827 14132 2836
rect 14284 2827 14324 2836
rect 13804 2575 13844 2584
rect 13228 1903 13268 1912
rect 13132 1819 13172 1828
rect 5452 1700 5492 1709
rect 4928 1532 5296 1541
rect 4968 1492 5010 1532
rect 5050 1492 5092 1532
rect 5132 1492 5174 1532
rect 5214 1492 5256 1532
rect 4928 1483 5296 1492
rect 5452 80 5492 1660
rect 6988 1700 7028 1709
rect 6988 80 7028 1660
rect 8524 1700 8564 1709
rect 8524 80 8564 1660
rect 10060 1700 10100 1709
rect 10060 80 10100 1660
rect 11596 1700 11636 1709
rect 11596 80 11636 1660
rect 13132 104 13172 113
rect 2360 0 2440 80
rect 3896 0 3976 80
rect 5432 0 5512 80
rect 6968 0 7048 80
rect 8504 0 8584 80
rect 10040 0 10120 80
rect 11576 0 11656 80
rect 13112 64 13132 80
rect 14668 80 14708 8044
rect 14764 1616 14804 8632
rect 15052 8672 15092 8681
rect 14860 8588 14900 8597
rect 14860 7244 14900 8548
rect 14860 6488 14900 7204
rect 14860 6439 14900 6448
rect 15052 3548 15092 8632
rect 15148 8168 15188 9808
rect 15244 8924 15284 11764
rect 15436 9680 15476 11764
rect 15436 9631 15476 9640
rect 15532 10016 15572 10025
rect 15244 8875 15284 8884
rect 15340 9512 15380 9521
rect 15148 8119 15188 8128
rect 15244 8672 15284 8681
rect 15244 5648 15284 8632
rect 15340 7832 15380 9472
rect 15532 9512 15572 9976
rect 15532 9463 15572 9472
rect 15628 8924 15668 11764
rect 15820 9680 15860 11764
rect 15820 9631 15860 9640
rect 15628 8875 15668 8884
rect 16012 8924 16052 11764
rect 16012 8875 16052 8884
rect 16108 9932 16148 9941
rect 16108 8756 16148 9892
rect 16204 9680 16244 11764
rect 16300 9932 16340 9941
rect 16300 9764 16340 9892
rect 16300 9715 16340 9724
rect 16204 9631 16244 9640
rect 16204 9512 16244 9521
rect 16204 9176 16244 9472
rect 16204 9127 16244 9136
rect 16396 8924 16436 11764
rect 16588 9680 16628 11764
rect 16588 9631 16628 9640
rect 16396 8875 16436 8884
rect 16492 9512 16532 9521
rect 16012 8716 16148 8756
rect 15532 8672 15572 8681
rect 15532 7916 15572 8632
rect 15532 7867 15572 7876
rect 15916 8672 15956 8681
rect 15340 7783 15380 7792
rect 15916 7832 15956 8632
rect 15916 7783 15956 7792
rect 15820 7748 15860 7757
rect 15244 5599 15284 5608
rect 15436 7580 15476 7589
rect 15052 3499 15092 3508
rect 15436 3464 15476 7540
rect 15820 6404 15860 7708
rect 15820 6355 15860 6364
rect 15436 3415 15476 3424
rect 15628 3968 15668 3977
rect 15052 3380 15092 3391
rect 15052 3296 15092 3340
rect 15052 3247 15092 3256
rect 15532 3212 15572 3221
rect 15532 2708 15572 3172
rect 15628 2792 15668 3928
rect 15628 2743 15668 2752
rect 15532 2659 15572 2668
rect 16012 1700 16052 8716
rect 16204 8252 16244 8261
rect 16108 7916 16148 7925
rect 16108 7244 16148 7876
rect 16204 7832 16244 8212
rect 16204 7783 16244 7792
rect 16300 8000 16340 8009
rect 16108 7195 16148 7204
rect 16204 3464 16244 3473
rect 16204 2456 16244 3424
rect 16300 3296 16340 7960
rect 16492 3884 16532 9472
rect 16684 9008 16724 9017
rect 16684 8672 16724 8968
rect 16780 8924 16820 11764
rect 16972 9680 17012 11764
rect 16972 9631 17012 9640
rect 16876 9512 16916 9521
rect 16876 9008 16916 9472
rect 16876 8959 16916 8968
rect 16780 8875 16820 8884
rect 17164 8924 17204 11764
rect 17356 9680 17396 11764
rect 17356 9631 17396 9640
rect 17164 8875 17204 8884
rect 17260 9512 17300 9521
rect 16684 8623 16724 8632
rect 17164 7748 17204 7757
rect 17164 7160 17204 7708
rect 17164 6488 17204 7120
rect 17164 6439 17204 6448
rect 16492 3835 16532 3844
rect 16876 6236 16916 6245
rect 16300 3247 16340 3256
rect 16876 3296 16916 6196
rect 17260 3632 17300 9472
rect 17452 9260 17492 9269
rect 17356 8588 17396 8597
rect 17356 6488 17396 8548
rect 17452 8252 17492 9220
rect 17548 8924 17588 11764
rect 17740 9680 17780 11764
rect 17740 9631 17780 9640
rect 17548 8875 17588 8884
rect 17644 9512 17684 9521
rect 17548 8756 17588 8767
rect 17548 8672 17588 8716
rect 17548 8623 17588 8632
rect 17452 8203 17492 8212
rect 17356 6439 17396 6448
rect 17452 6404 17492 6413
rect 17452 6152 17492 6364
rect 17644 6404 17684 9472
rect 17836 9428 17876 9437
rect 17644 6355 17684 6364
rect 17740 8672 17780 8681
rect 17452 6103 17492 6112
rect 17740 3716 17780 8632
rect 17836 8168 17876 9388
rect 17932 8924 17972 11764
rect 18124 9680 18164 11764
rect 18124 9631 18164 9640
rect 17932 8875 17972 8884
rect 18028 9512 18068 9521
rect 17836 8119 17876 8128
rect 17932 7664 17972 7673
rect 17740 3667 17780 3676
rect 17836 4892 17876 4901
rect 17260 3583 17300 3592
rect 16876 3247 16916 3256
rect 17644 3212 17684 3221
rect 17644 2708 17684 3172
rect 17644 2659 17684 2668
rect 17836 2456 17876 4852
rect 17932 4136 17972 7624
rect 18028 6908 18068 9472
rect 18316 8924 18356 11764
rect 18412 10016 18452 10025
rect 18412 9764 18452 9976
rect 18412 9715 18452 9724
rect 18508 9680 18548 11764
rect 18508 9631 18548 9640
rect 18604 10100 18644 10109
rect 18316 8875 18356 8884
rect 18412 9512 18452 9521
rect 18220 8672 18260 8681
rect 18124 8504 18164 8513
rect 18124 8000 18164 8464
rect 18124 7951 18164 7960
rect 18028 6859 18068 6868
rect 18220 6740 18260 8632
rect 18412 7664 18452 9472
rect 18604 9512 18644 10060
rect 18604 9463 18644 9472
rect 18700 8924 18740 11764
rect 18892 10016 18932 11764
rect 19084 10268 19124 11764
rect 19276 10352 19316 11764
rect 19276 10312 19412 10352
rect 19084 10228 19316 10268
rect 18892 9967 18932 9976
rect 19180 10100 19220 10109
rect 19180 9965 19220 10060
rect 18808 9848 19176 9857
rect 18848 9808 18890 9848
rect 18930 9808 18972 9848
rect 19012 9808 19054 9848
rect 19094 9808 19136 9848
rect 18808 9799 19176 9808
rect 19180 9680 19220 9689
rect 19084 9596 19124 9607
rect 19084 9512 19124 9556
rect 19084 9463 19124 9472
rect 19180 9344 19220 9640
rect 19180 9295 19220 9304
rect 18700 8875 18740 8884
rect 19180 8924 19220 8933
rect 18604 8672 18644 8681
rect 18508 8336 18548 8345
rect 18508 7916 18548 8296
rect 18508 7867 18548 7876
rect 18412 7615 18452 7624
rect 18220 6691 18260 6700
rect 18604 5900 18644 8632
rect 19180 8672 19220 8884
rect 19276 8924 19316 10228
rect 19372 9596 19412 10312
rect 19372 9547 19412 9556
rect 19372 9428 19412 9437
rect 19372 9344 19412 9388
rect 19372 9293 19412 9304
rect 19372 9176 19412 9185
rect 19372 9008 19412 9136
rect 19372 8959 19412 8968
rect 19276 8875 19316 8884
rect 19468 8924 19508 11764
rect 19564 10268 19604 10277
rect 19564 9932 19604 10228
rect 19564 9883 19604 9892
rect 19564 9680 19604 9689
rect 19564 9512 19604 9640
rect 19564 9463 19604 9472
rect 19660 9428 19700 11764
rect 19852 10520 19892 11764
rect 19852 10471 19892 10480
rect 20044 10184 20084 11764
rect 19756 10144 20084 10184
rect 19756 9680 19796 10144
rect 20044 10016 20084 10025
rect 20140 10016 20180 10025
rect 20084 9976 20140 10016
rect 20044 9967 20084 9976
rect 20140 9967 20180 9976
rect 19756 9631 19796 9640
rect 19852 9680 19892 9689
rect 20044 9680 20084 9689
rect 19892 9640 20044 9680
rect 19852 9631 19892 9640
rect 20044 9631 20084 9640
rect 20140 9512 20180 9521
rect 19948 9472 20140 9512
rect 19660 9379 19700 9388
rect 19756 9428 19796 9437
rect 19564 9344 19604 9353
rect 19564 9092 19604 9304
rect 19564 9043 19604 9052
rect 19468 8875 19508 8884
rect 19660 9008 19700 9017
rect 19180 8623 19220 8632
rect 18808 8336 19176 8345
rect 18848 8296 18890 8336
rect 18930 8296 18972 8336
rect 19012 8296 19054 8336
rect 19094 8296 19136 8336
rect 18808 8287 19176 8296
rect 19660 7748 19700 8968
rect 19756 8840 19796 9388
rect 19948 9428 19988 9472
rect 20140 9463 20180 9472
rect 19948 9379 19988 9388
rect 20236 9344 20276 11764
rect 20428 9680 20468 11764
rect 20428 9631 20468 9640
rect 20236 9304 20564 9344
rect 20048 9092 20416 9101
rect 20088 9052 20130 9092
rect 20170 9052 20212 9092
rect 20252 9052 20294 9092
rect 20334 9052 20376 9092
rect 20048 9043 20416 9052
rect 19852 9008 19892 9019
rect 19852 8924 19892 8968
rect 19852 8875 19892 8884
rect 20044 8924 20084 8933
rect 20044 8840 20084 8884
rect 20524 8924 20564 9304
rect 20524 8875 20564 8884
rect 20236 8840 20276 8849
rect 20044 8800 20236 8840
rect 19756 8791 19796 8800
rect 20236 8791 20276 8800
rect 20428 8840 20468 8849
rect 19852 8756 19892 8765
rect 19660 7699 19700 7708
rect 19756 8672 19796 8681
rect 19756 7160 19796 8632
rect 19756 7111 19796 7120
rect 18808 6824 19176 6833
rect 18848 6784 18890 6824
rect 18930 6784 18972 6824
rect 19012 6784 19054 6824
rect 19094 6784 19136 6824
rect 18808 6775 19176 6784
rect 19852 6488 19892 8716
rect 19948 8672 19988 8767
rect 19948 8623 19988 8632
rect 20140 8588 20180 8597
rect 20140 8453 20180 8548
rect 20140 8168 20180 8177
rect 20140 8033 20180 8128
rect 20428 7748 20468 8800
rect 20620 8840 20660 11764
rect 20812 9680 20852 11764
rect 20812 9631 20852 9640
rect 20620 8791 20660 8800
rect 20716 9260 20756 9269
rect 20428 7708 20660 7748
rect 20048 7580 20416 7589
rect 20088 7540 20130 7580
rect 20170 7540 20212 7580
rect 20252 7540 20294 7580
rect 20334 7540 20376 7580
rect 20048 7531 20416 7540
rect 20140 7412 20180 7421
rect 20140 7277 20180 7372
rect 19852 6439 19892 6448
rect 20048 6068 20416 6077
rect 20088 6028 20130 6068
rect 20170 6028 20212 6068
rect 20252 6028 20294 6068
rect 20334 6028 20376 6068
rect 20048 6019 20416 6028
rect 18604 5851 18644 5860
rect 18808 5312 19176 5321
rect 18848 5272 18890 5312
rect 18930 5272 18972 5312
rect 19012 5272 19054 5312
rect 19094 5272 19136 5312
rect 18808 5263 19176 5272
rect 20048 4556 20416 4565
rect 20088 4516 20130 4556
rect 20170 4516 20212 4556
rect 20252 4516 20294 4556
rect 20334 4516 20376 4556
rect 20048 4507 20416 4516
rect 19756 4388 19796 4397
rect 19756 4253 19796 4348
rect 17932 4087 17972 4096
rect 19276 4220 19316 4229
rect 19180 3968 19220 4063
rect 19180 3919 19220 3928
rect 18808 3800 19176 3809
rect 18848 3760 18890 3800
rect 18930 3760 18972 3800
rect 19012 3760 19054 3800
rect 19094 3760 19136 3800
rect 18808 3751 19176 3760
rect 19276 3632 19316 4180
rect 19276 3583 19316 3592
rect 19660 4136 19700 4145
rect 19660 3800 19700 4096
rect 19852 4136 19892 4145
rect 18796 3548 18836 3557
rect 18700 3508 18796 3548
rect 18220 3464 18260 3473
rect 18220 3212 18260 3424
rect 18508 3380 18548 3389
rect 18220 3163 18260 3172
rect 18412 3340 18508 3380
rect 18412 3212 18452 3340
rect 18508 3331 18548 3340
rect 18412 3163 18452 3172
rect 18700 2876 18740 3508
rect 18796 3499 18836 3508
rect 19372 3548 19412 3557
rect 19372 3464 19412 3508
rect 19276 3424 19372 3464
rect 16204 2407 16244 2416
rect 17740 2416 17876 2456
rect 18604 2836 18740 2876
rect 18796 3212 18836 3221
rect 16012 1651 16052 1660
rect 16204 2204 16244 2213
rect 14764 1567 14804 1576
rect 16204 80 16244 2164
rect 17740 80 17780 2416
rect 18604 2288 18644 2836
rect 18604 2239 18644 2248
rect 18700 2708 18740 2717
rect 18700 2036 18740 2668
rect 18796 2624 18836 3172
rect 19276 2708 19316 3424
rect 19372 3413 19412 3424
rect 19660 3380 19700 3760
rect 19660 3331 19700 3340
rect 19756 3968 19796 3977
rect 19756 3212 19796 3928
rect 19852 3464 19892 4096
rect 19852 3415 19892 3424
rect 20524 3464 20564 3473
rect 19564 3128 19604 3137
rect 19372 2960 19412 2969
rect 19564 2960 19604 3088
rect 19412 2920 19604 2960
rect 19372 2911 19412 2920
rect 19276 2659 19316 2668
rect 19660 2792 19700 2801
rect 19660 2657 19700 2752
rect 19756 2708 19796 3172
rect 20048 3044 20416 3053
rect 20088 3004 20130 3044
rect 20170 3004 20212 3044
rect 20252 3004 20294 3044
rect 20334 3004 20376 3044
rect 20048 2995 20416 3004
rect 19756 2659 19796 2668
rect 18796 2575 18836 2584
rect 20524 2624 20564 3424
rect 20620 2876 20660 7708
rect 20620 2827 20660 2836
rect 20716 2792 20756 9220
rect 20812 9008 20852 9017
rect 20812 8873 20852 8968
rect 21004 8924 21044 11764
rect 21004 8875 21044 8884
rect 21100 9848 21140 9857
rect 20908 8672 20948 8681
rect 20908 5144 20948 8632
rect 20908 5095 20948 5104
rect 21100 4304 21140 9808
rect 21196 9596 21236 11764
rect 21196 9547 21236 9556
rect 20716 2743 20756 2752
rect 20812 4136 20852 4145
rect 20524 2575 20564 2584
rect 19852 2456 19892 2465
rect 18808 2288 19176 2297
rect 18848 2248 18890 2288
rect 18930 2248 18972 2288
rect 19012 2248 19054 2288
rect 19094 2248 19136 2288
rect 18808 2239 19176 2248
rect 18700 1996 18836 2036
rect 18604 1952 18644 1961
rect 18796 1952 18836 1996
rect 18644 1912 18740 1952
rect 18604 1903 18644 1912
rect 18700 1700 18740 1912
rect 18796 1903 18836 1912
rect 18700 1651 18740 1660
rect 19852 1616 19892 2416
rect 19852 1567 19892 1576
rect 20048 1532 20416 1541
rect 20088 1492 20130 1532
rect 20170 1492 20212 1532
rect 20252 1492 20294 1532
rect 20334 1492 20376 1532
rect 20048 1483 20416 1492
rect 19276 188 19316 197
rect 19276 80 19316 148
rect 20812 80 20852 4096
rect 21100 4136 21140 4264
rect 21100 4087 21140 4096
rect 21196 9260 21236 9269
rect 21196 1952 21236 9220
rect 21292 8924 21332 9019
rect 21292 8875 21332 8884
rect 21292 8756 21332 8765
rect 21292 2876 21332 8716
rect 21388 8672 21428 11764
rect 21580 9596 21620 11764
rect 21580 9547 21620 9556
rect 21676 8840 21716 8849
rect 21388 8623 21428 8632
rect 21484 8672 21524 8681
rect 21388 4388 21428 4397
rect 21388 3716 21428 4348
rect 21484 4136 21524 8632
rect 21580 8588 21620 8597
rect 21580 5816 21620 8548
rect 21676 8000 21716 8800
rect 21772 8672 21812 11764
rect 21964 9596 22004 11764
rect 21964 9547 22004 9556
rect 22156 9596 22196 11764
rect 22156 9547 22196 9556
rect 22348 9512 22388 11764
rect 22348 9463 22388 9472
rect 22540 9512 22580 11764
rect 22732 9932 22772 11764
rect 22924 10016 22964 11764
rect 23116 10184 23156 11764
rect 23348 11764 23368 11780
rect 23480 11764 23560 11844
rect 23672 11764 23752 11844
rect 23864 11764 23944 11844
rect 24056 11764 24136 11844
rect 24248 11764 24328 11844
rect 24440 11764 24520 11844
rect 24632 11764 24712 11844
rect 24824 11764 24904 11844
rect 25016 11764 25096 11844
rect 25208 11764 25288 11844
rect 25400 11764 25480 11844
rect 25592 11764 25672 11844
rect 25784 11764 25864 11844
rect 25976 11764 26056 11844
rect 26168 11764 26248 11844
rect 26360 11764 26440 11844
rect 26552 11764 26632 11844
rect 26744 11780 26824 11844
rect 26744 11764 26764 11780
rect 23308 11731 23348 11740
rect 23116 10144 23252 10184
rect 22540 9463 22580 9472
rect 22636 9892 22772 9932
rect 22828 9976 22964 10016
rect 22540 9260 22580 9269
rect 21772 8623 21812 8632
rect 22156 9092 22196 9101
rect 22060 8504 22100 8513
rect 22060 8084 22100 8464
rect 22060 8035 22100 8044
rect 21676 7951 21716 7960
rect 22156 7412 22196 9052
rect 22444 8336 22484 8345
rect 22444 7832 22484 8296
rect 22444 7783 22484 7792
rect 22156 7363 22196 7372
rect 21580 5767 21620 5776
rect 21676 6992 21716 7001
rect 21484 4087 21524 4096
rect 21580 4220 21620 4229
rect 21388 3667 21428 3676
rect 21484 3968 21524 3977
rect 21484 3716 21524 3928
rect 21484 3667 21524 3676
rect 21580 3716 21620 4180
rect 21580 3667 21620 3676
rect 21676 4136 21716 6952
rect 22540 6656 22580 9220
rect 22636 8336 22676 9892
rect 22828 9092 22868 9976
rect 22828 9043 22868 9052
rect 22924 9344 22964 9353
rect 22636 8287 22676 8296
rect 22828 8840 22868 8849
rect 22636 8000 22676 8009
rect 22636 7244 22676 7960
rect 22636 7195 22676 7204
rect 22540 6607 22580 6616
rect 21772 6404 21812 6413
rect 21772 5816 21812 6364
rect 21772 5767 21812 5776
rect 21676 3632 21716 4096
rect 21868 5396 21908 5405
rect 21868 4136 21908 5356
rect 21964 4304 22004 4313
rect 21964 4220 22004 4264
rect 21964 4169 22004 4180
rect 21868 4087 21908 4096
rect 21772 3968 21812 3977
rect 21772 3833 21812 3928
rect 21580 3548 21620 3557
rect 21388 3508 21580 3548
rect 21388 3464 21428 3508
rect 21580 3499 21620 3508
rect 21388 3415 21428 3424
rect 21292 2827 21332 2836
rect 21484 3380 21524 3389
rect 21484 2708 21524 3340
rect 21580 3296 21620 3305
rect 21580 3161 21620 3256
rect 21676 3212 21716 3592
rect 21772 3716 21812 3725
rect 21772 3380 21812 3676
rect 21772 3331 21812 3340
rect 21964 3464 22004 3473
rect 21676 3163 21716 3172
rect 21964 3212 22004 3424
rect 22828 3464 22868 8800
rect 22924 8168 22964 9304
rect 23116 9092 23156 9101
rect 23116 9008 23156 9052
rect 23116 8957 23156 8968
rect 22924 8119 22964 8128
rect 23212 7328 23252 10144
rect 23308 9344 23348 9353
rect 23308 8840 23348 9304
rect 23308 8791 23348 8800
rect 23212 7279 23252 7288
rect 23308 8672 23348 8681
rect 23308 3632 23348 8632
rect 23500 8672 23540 11764
rect 23692 9596 23732 11764
rect 23692 9547 23732 9556
rect 23884 9512 23924 11764
rect 23884 9463 23924 9472
rect 23980 9680 24020 9689
rect 23692 9344 23732 9353
rect 23500 8623 23540 8632
rect 23596 9260 23636 9269
rect 23596 6572 23636 9220
rect 23692 9092 23732 9304
rect 23692 9043 23732 9052
rect 23980 8840 24020 9640
rect 24076 9512 24116 11764
rect 24076 9463 24116 9472
rect 24172 10100 24212 10109
rect 24172 9176 24212 10060
rect 24268 9596 24308 11764
rect 24268 9547 24308 9556
rect 24364 9680 24404 9689
rect 24364 9545 24404 9640
rect 24460 9596 24500 11764
rect 24460 9547 24500 9556
rect 24556 10016 24596 10025
rect 24556 9428 24596 9976
rect 24652 9680 24692 11764
rect 24652 9631 24692 9640
rect 24556 9379 24596 9388
rect 24844 9428 24884 11764
rect 25036 10100 25076 11764
rect 25036 10051 25076 10060
rect 24844 9379 24884 9388
rect 25036 9344 25076 9353
rect 24172 9127 24212 9136
rect 24364 9260 24404 9269
rect 23980 8791 24020 8800
rect 23596 6523 23636 6532
rect 24076 5564 24116 5573
rect 24076 4304 24116 5524
rect 24076 4255 24116 4264
rect 24268 5228 24308 5237
rect 23308 3583 23348 3592
rect 22828 3415 22868 3424
rect 21964 3163 22004 3172
rect 24268 3380 24308 5188
rect 24364 3548 24404 9220
rect 24364 3499 24404 3508
rect 24460 9092 24500 9101
rect 24172 3128 24212 3137
rect 24172 2993 24212 3088
rect 21484 2659 21524 2668
rect 24268 2624 24308 3340
rect 24460 3128 24500 9052
rect 25036 9092 25076 9304
rect 25036 9043 25076 9052
rect 25132 9260 25172 9269
rect 25036 8924 25076 8933
rect 24940 8672 24980 8683
rect 24940 8588 24980 8632
rect 24940 8539 24980 8548
rect 24652 7916 24692 7925
rect 24652 7244 24692 7876
rect 24652 7195 24692 7204
rect 25036 3800 25076 8884
rect 25132 6320 25172 9220
rect 25228 8672 25268 11764
rect 25228 8623 25268 8632
rect 25324 9680 25364 9689
rect 25132 6271 25172 6280
rect 25228 8504 25268 8513
rect 25036 3751 25076 3760
rect 25036 3548 25076 3557
rect 25036 3413 25076 3508
rect 25228 3548 25268 8464
rect 25228 3499 25268 3508
rect 24460 3079 24500 3088
rect 25324 3044 25364 9640
rect 25420 9596 25460 11764
rect 25420 9547 25460 9556
rect 25612 8672 25652 11764
rect 25804 9428 25844 11764
rect 25900 10100 25940 10109
rect 25900 9512 25940 10060
rect 25900 9463 25940 9472
rect 25804 9379 25844 9388
rect 25612 8623 25652 8632
rect 25708 9344 25748 9353
rect 25708 7664 25748 9304
rect 25900 8840 25940 8849
rect 25708 7615 25748 7624
rect 25804 8588 25844 8597
rect 25420 4220 25460 4229
rect 25420 3380 25460 4180
rect 25420 3331 25460 3340
rect 25516 3800 25556 3809
rect 25324 2995 25364 3004
rect 25516 2900 25556 3760
rect 25804 3716 25844 8548
rect 25900 8084 25940 8800
rect 25996 8756 26036 11764
rect 26092 9764 26132 9773
rect 26092 8756 26132 9724
rect 26188 9680 26228 11764
rect 26380 9764 26420 11764
rect 26380 9715 26420 9724
rect 26188 9631 26228 9640
rect 26284 9680 26324 9689
rect 26188 8756 26228 8765
rect 26092 8716 26188 8756
rect 25996 8707 26036 8716
rect 26188 8707 26228 8716
rect 25900 8035 25940 8044
rect 26092 8252 26132 8261
rect 26092 7832 26132 8212
rect 26092 7783 26132 7792
rect 26188 7916 26228 7925
rect 26188 7244 26228 7876
rect 26188 6992 26228 7204
rect 26188 6943 26228 6952
rect 26284 7328 26324 9640
rect 26476 9344 26516 9353
rect 26284 6824 26324 7288
rect 26380 9176 26420 9185
rect 26380 7748 26420 9136
rect 26476 7916 26516 9304
rect 26572 8672 26612 11764
rect 26804 11764 26824 11780
rect 26936 11764 27016 11844
rect 27128 11764 27208 11844
rect 27320 11764 27400 11844
rect 27512 11764 27592 11844
rect 27704 11764 27784 11844
rect 27896 11764 27976 11844
rect 28088 11764 28168 11844
rect 28280 11764 28360 11844
rect 28472 11764 28552 11844
rect 28664 11764 28744 11844
rect 28856 11764 28936 11844
rect 29048 11764 29128 11844
rect 29240 11764 29320 11844
rect 29432 11764 29512 11844
rect 29624 11780 29704 11844
rect 29624 11764 29644 11780
rect 26764 11731 26804 11740
rect 26956 11696 26996 11764
rect 26956 11647 26996 11656
rect 26956 9764 26996 9773
rect 26956 9428 26996 9724
rect 27148 9596 27188 11764
rect 27244 10268 27284 10277
rect 27244 9848 27284 10228
rect 27244 9799 27284 9808
rect 27148 9556 27284 9596
rect 26956 9379 26996 9388
rect 26860 9344 26900 9353
rect 26572 8623 26612 8632
rect 26668 9176 26708 9185
rect 26668 8672 26708 9136
rect 26764 9092 26804 9101
rect 26764 8756 26804 9052
rect 26764 8707 26804 8716
rect 26668 7916 26708 8632
rect 26764 8588 26804 8597
rect 26764 8453 26804 8548
rect 26860 8000 26900 9304
rect 26860 7951 26900 7960
rect 26956 9260 26996 9269
rect 26764 7916 26804 7925
rect 26668 7876 26764 7916
rect 26476 7867 26516 7876
rect 26764 7867 26804 7876
rect 26380 7160 26420 7708
rect 26380 7111 26420 7120
rect 26092 6784 26324 6824
rect 26092 4220 26132 6784
rect 26092 4171 26132 4180
rect 26284 4304 26324 4313
rect 25804 3667 25844 3676
rect 26188 4136 26228 4145
rect 25612 3632 25652 3641
rect 25612 3296 25652 3592
rect 26188 3632 26228 4096
rect 26284 4052 26324 4264
rect 26572 4136 26612 4145
rect 26284 4003 26324 4012
rect 26476 4096 26572 4136
rect 26188 3583 26228 3592
rect 25900 3296 25940 3305
rect 25612 3256 25900 3296
rect 25900 3247 25940 3256
rect 26476 3212 26516 4096
rect 26572 4087 26612 4096
rect 26572 3968 26612 3977
rect 26572 3380 26612 3928
rect 26668 3548 26708 3557
rect 26956 3548 26996 9220
rect 27148 9260 27188 9269
rect 27052 9092 27092 9101
rect 27052 8957 27092 9052
rect 27148 8924 27188 9220
rect 27148 8875 27188 8884
rect 27052 8840 27092 8849
rect 27052 8672 27092 8800
rect 27092 8632 27188 8672
rect 27052 8623 27092 8632
rect 27052 7664 27092 7673
rect 27052 7244 27092 7624
rect 27148 7328 27188 8632
rect 27244 7664 27284 9556
rect 27340 9428 27380 11764
rect 27436 10352 27476 10361
rect 27436 9680 27476 10312
rect 27436 9631 27476 9640
rect 27340 9379 27380 9388
rect 27436 8588 27476 8597
rect 27244 7615 27284 7624
rect 27340 8504 27380 8513
rect 27148 7279 27188 7288
rect 27052 7195 27092 7204
rect 27052 5060 27092 5069
rect 27052 4304 27092 5020
rect 27052 4255 27092 4264
rect 26708 3508 26996 3548
rect 26668 3499 26708 3508
rect 26572 3331 26612 3340
rect 26668 3296 26708 3305
rect 26668 3212 26708 3256
rect 26516 3172 26708 3212
rect 26956 3296 26996 3305
rect 26476 3163 26516 3172
rect 25612 3128 25652 3137
rect 25612 3044 25652 3088
rect 25612 2993 25652 3004
rect 24268 2575 24308 2584
rect 25420 2860 25556 2900
rect 26860 2960 26900 2969
rect 21196 1903 21236 1912
rect 23116 1952 23156 1961
rect 22924 1868 22964 1879
rect 22924 1784 22964 1828
rect 22924 1735 22964 1744
rect 23020 1784 23060 1793
rect 23116 1784 23156 1912
rect 23060 1744 23156 1784
rect 23020 1735 23060 1744
rect 23884 356 23924 365
rect 22348 272 22388 281
rect 22348 80 22388 232
rect 23884 80 23924 316
rect 25420 80 25460 2860
rect 26860 2120 26900 2920
rect 26860 2071 26900 2080
rect 26956 80 26996 3256
rect 27340 2960 27380 8464
rect 27436 7916 27476 8548
rect 27532 8504 27572 11764
rect 27532 8455 27572 8464
rect 27628 8756 27668 8765
rect 27436 7867 27476 7876
rect 27628 7748 27668 8716
rect 27724 8336 27764 11764
rect 27916 9344 27956 11764
rect 28108 9512 28148 11764
rect 28108 9463 28148 9472
rect 28204 10100 28244 10109
rect 27916 9304 28148 9344
rect 27724 8287 27764 8296
rect 28012 8672 28052 8681
rect 27628 7699 27668 7708
rect 27916 7832 27956 7841
rect 27916 7580 27956 7792
rect 27916 7531 27956 7540
rect 28012 7412 28052 8632
rect 28108 7412 28148 9304
rect 28204 8840 28244 10060
rect 28300 9596 28340 11764
rect 28492 9680 28532 11764
rect 28492 9631 28532 9640
rect 28300 9547 28340 9556
rect 28684 9428 28724 11764
rect 28876 9764 28916 11764
rect 28876 9715 28916 9724
rect 28972 9848 29012 9857
rect 28684 9379 28724 9388
rect 28588 9176 28628 9185
rect 28204 8791 28244 8800
rect 28396 9008 28436 9017
rect 28204 8168 28244 8177
rect 28204 8033 28244 8128
rect 28396 8168 28436 8968
rect 28396 8119 28436 8128
rect 28204 7412 28244 7421
rect 28108 7372 28204 7412
rect 28012 7363 28052 7372
rect 28204 7363 28244 7372
rect 28396 7328 28436 7337
rect 28396 7160 28436 7288
rect 28396 7111 28436 7120
rect 27916 4136 27956 4145
rect 27436 4052 27476 4061
rect 27436 3548 27476 4012
rect 27436 3499 27476 3508
rect 27628 3464 27668 3475
rect 27628 3380 27668 3424
rect 27628 3331 27668 3340
rect 27916 3044 27956 4096
rect 28588 4052 28628 9136
rect 28588 4003 28628 4012
rect 28684 8924 28724 8933
rect 28684 3548 28724 8884
rect 28876 8504 28916 8513
rect 28780 8336 28820 8345
rect 28780 8168 28820 8296
rect 28780 8119 28820 8128
rect 28780 7916 28820 7925
rect 28780 7244 28820 7876
rect 28876 7496 28916 8464
rect 28972 8000 29012 9808
rect 29068 8672 29108 11764
rect 29260 9848 29300 11764
rect 29260 9799 29300 9808
rect 29164 9260 29204 9269
rect 29164 9008 29204 9220
rect 29164 8959 29204 8968
rect 29068 8623 29108 8632
rect 29452 8672 29492 11764
rect 29684 11764 29704 11780
rect 29816 11764 29896 11844
rect 30008 11764 30088 11844
rect 30200 11764 30280 11844
rect 30392 11764 30472 11844
rect 30584 11764 30664 11844
rect 30776 11764 30856 11844
rect 30968 11764 31048 11844
rect 31160 11764 31240 11844
rect 31352 11764 31432 11844
rect 31544 11764 31624 11844
rect 31736 11764 31816 11844
rect 31928 11764 32008 11844
rect 32120 11764 32200 11844
rect 32312 11764 32392 11844
rect 32504 11764 32584 11844
rect 32696 11764 32776 11844
rect 32888 11764 32968 11844
rect 33080 11764 33160 11844
rect 33272 11764 33352 11844
rect 33464 11764 33544 11844
rect 33656 11764 33736 11844
rect 33848 11764 33928 11844
rect 34040 11764 34120 11844
rect 34232 11764 34312 11844
rect 34424 11764 34504 11844
rect 34616 11764 34696 11844
rect 34808 11764 34888 11844
rect 35000 11764 35080 11844
rect 41740 11780 41780 11789
rect 29644 11731 29684 11740
rect 29836 10100 29876 11764
rect 29836 10051 29876 10060
rect 29836 9260 29876 9269
rect 29452 8623 29492 8632
rect 29740 8840 29780 8849
rect 29068 8000 29108 8009
rect 28972 7960 29068 8000
rect 29068 7951 29108 7960
rect 29452 8000 29492 8009
rect 28876 7447 28916 7456
rect 28780 7195 28820 7204
rect 29452 7244 29492 7960
rect 29452 7195 29492 7204
rect 29740 4052 29780 8800
rect 29836 8756 29876 9220
rect 29836 8707 29876 8716
rect 30028 8336 30068 11764
rect 30028 8287 30068 8296
rect 30220 6572 30260 11764
rect 30316 8672 30356 8683
rect 30316 8588 30356 8632
rect 30316 8539 30356 8548
rect 30220 6523 30260 6532
rect 30412 6320 30452 11764
rect 30412 6271 30452 6280
rect 30604 6068 30644 11764
rect 30796 6656 30836 11764
rect 30796 6607 30836 6616
rect 30892 9008 30932 9017
rect 30604 6019 30644 6028
rect 29740 4003 29780 4012
rect 30028 4220 30068 4229
rect 28684 3499 28724 3508
rect 30028 3464 30068 4180
rect 30028 3415 30068 3424
rect 30508 4220 30548 4229
rect 30508 3380 30548 4180
rect 30892 3464 30932 8968
rect 30988 6404 31028 11764
rect 31180 9680 31220 11764
rect 31180 9631 31220 9640
rect 31372 9596 31412 11764
rect 31564 9680 31604 11764
rect 31564 9631 31604 9640
rect 31372 9547 31412 9556
rect 31756 9596 31796 11764
rect 31756 9547 31796 9556
rect 31468 9512 31508 9521
rect 31468 8420 31508 9472
rect 31660 9512 31700 9521
rect 31468 8371 31508 8380
rect 31564 8672 31604 8681
rect 30988 6355 31028 6364
rect 31180 8000 31220 8009
rect 31180 7244 31220 7960
rect 31468 7664 31508 7673
rect 31468 7412 31508 7624
rect 31468 7363 31508 7372
rect 31180 4136 31220 7204
rect 31180 4087 31220 4096
rect 31372 4220 31412 4229
rect 31372 3548 31412 4180
rect 31564 4220 31604 8632
rect 31564 4171 31604 4180
rect 31660 3968 31700 9472
rect 31948 9344 31988 11764
rect 31948 9295 31988 9304
rect 32044 9260 32084 9269
rect 31660 3919 31700 3928
rect 31756 9008 31796 9017
rect 31372 3499 31412 3508
rect 30892 3415 30932 3424
rect 31180 3464 31220 3473
rect 30508 3331 30548 3340
rect 30796 3380 30836 3389
rect 30220 3212 30260 3221
rect 30796 3212 30836 3340
rect 30260 3172 30836 3212
rect 30220 3163 30260 3172
rect 27916 2995 27956 3004
rect 27340 2911 27380 2920
rect 28492 2960 28532 2969
rect 27052 2456 27092 2465
rect 27052 1700 27092 2416
rect 27052 1651 27092 1660
rect 28492 80 28532 2920
rect 31180 2624 31220 3424
rect 31756 3380 31796 8968
rect 31948 8924 31988 8933
rect 31948 8789 31988 8884
rect 32044 4472 32084 9220
rect 32140 8924 32180 11764
rect 32140 8875 32180 8884
rect 32236 9512 32276 9521
rect 32044 4423 32084 4432
rect 32140 7328 32180 7337
rect 32140 4892 32180 7288
rect 31852 4220 31892 4229
rect 31852 3716 31892 4180
rect 32140 4136 32180 4852
rect 32140 4087 32180 4096
rect 31852 3464 31892 3676
rect 31852 3415 31892 3424
rect 32044 4052 32084 4061
rect 31276 3296 31316 3305
rect 31276 2708 31316 3256
rect 31276 2659 31316 2668
rect 31564 3128 31604 3137
rect 31180 2575 31220 2584
rect 30220 2204 30260 2213
rect 30220 2069 30260 2164
rect 30028 1952 30068 1961
rect 30028 80 30068 1912
rect 30220 1784 30260 1793
rect 30220 1649 30260 1744
rect 31564 80 31604 3088
rect 31756 2708 31796 3340
rect 31756 2659 31796 2668
rect 32044 2288 32084 4012
rect 32044 2239 32084 2248
rect 32236 1616 32276 9472
rect 32332 9260 32372 11764
rect 32332 9211 32372 9220
rect 32524 8924 32564 11764
rect 32716 9596 32756 11764
rect 32716 9547 32756 9556
rect 32524 8875 32564 8884
rect 32908 8924 32948 11764
rect 33100 11444 33140 11764
rect 33100 11404 33236 11444
rect 33100 9512 33140 9521
rect 33100 9092 33140 9472
rect 33196 9260 33236 11404
rect 33196 9211 33236 9220
rect 33100 9052 33236 9092
rect 32908 8875 32948 8884
rect 32620 8840 32660 8849
rect 32620 6992 32660 8800
rect 33100 8756 33140 8765
rect 33100 8672 33140 8716
rect 33196 8672 33236 9052
rect 33292 8924 33332 11764
rect 33484 9680 33524 11764
rect 33484 9631 33524 9640
rect 33388 9512 33428 9521
rect 33388 9344 33428 9472
rect 33388 9295 33428 9304
rect 33292 8875 33332 8884
rect 33484 9008 33524 9017
rect 33484 8756 33524 8968
rect 33676 8924 33716 11764
rect 33868 10016 33908 11764
rect 34060 10016 34100 11764
rect 34252 10184 34292 11764
rect 34252 10135 34292 10144
rect 34060 9976 34388 10016
rect 33868 9967 33908 9976
rect 33928 9848 34296 9857
rect 33968 9808 34010 9848
rect 34050 9808 34092 9848
rect 34132 9808 34174 9848
rect 34214 9808 34256 9848
rect 33928 9799 34296 9808
rect 33772 9512 33812 9607
rect 33772 9463 33812 9472
rect 34156 9512 34196 9521
rect 33676 8875 33716 8884
rect 33772 9344 33812 9353
rect 33484 8707 33524 8716
rect 33388 8672 33428 8681
rect 33772 8672 33812 9304
rect 33196 8632 33332 8672
rect 33100 8621 33140 8632
rect 33292 8252 33332 8632
rect 33292 8203 33332 8212
rect 33004 8084 33044 8093
rect 33004 7916 33044 8044
rect 33004 7867 33044 7876
rect 33292 8084 33332 8093
rect 32620 6943 32660 6952
rect 33004 7748 33044 7757
rect 32812 6488 32852 6497
rect 32428 4472 32468 4481
rect 32332 4304 32372 4313
rect 32332 3380 32372 4264
rect 32428 4136 32468 4432
rect 32428 4087 32468 4096
rect 32524 4220 32564 4229
rect 32332 3331 32372 3340
rect 32428 3968 32468 3977
rect 32428 2120 32468 3928
rect 32524 3716 32564 4180
rect 32524 3667 32564 3676
rect 32812 3548 32852 6448
rect 32908 4976 32948 4985
rect 32908 4472 32948 4936
rect 32908 4423 32948 4432
rect 33004 4220 33044 7708
rect 33196 7748 33236 7757
rect 33100 7580 33140 7589
rect 33100 7445 33140 7540
rect 33196 7244 33236 7708
rect 33292 7664 33332 8044
rect 33292 7615 33332 7624
rect 33196 4388 33236 7204
rect 33196 4339 33236 4348
rect 33292 5228 33332 5237
rect 33004 4171 33044 4180
rect 33196 4220 33236 4229
rect 32908 4052 32948 4061
rect 32908 3716 32948 4012
rect 33004 3884 33044 3893
rect 33004 3800 33044 3844
rect 33196 3884 33236 4180
rect 33196 3835 33236 3844
rect 33004 3749 33044 3760
rect 32908 3667 32948 3676
rect 32812 3499 32852 3508
rect 33100 3296 33140 3305
rect 33004 3256 33100 3296
rect 33004 3044 33044 3256
rect 33100 3247 33140 3256
rect 33004 2995 33044 3004
rect 33292 2900 33332 5188
rect 33388 4472 33428 8632
rect 33676 8632 33812 8672
rect 33388 4423 33428 4432
rect 33484 8588 33524 8597
rect 33484 4052 33524 8548
rect 33580 8504 33620 8599
rect 33580 8455 33620 8464
rect 33580 8252 33620 8347
rect 33580 8203 33620 8212
rect 33580 8084 33620 8093
rect 33580 7949 33620 8044
rect 33484 4003 33524 4012
rect 33580 4220 33620 4229
rect 33580 3380 33620 4180
rect 33580 3331 33620 3340
rect 33676 3212 33716 8632
rect 33772 8504 33812 8513
rect 34156 8504 34196 9472
rect 34348 8924 34388 9976
rect 34348 8875 34388 8884
rect 34444 8840 34484 11764
rect 34540 10184 34580 10193
rect 34540 9344 34580 10144
rect 34636 9596 34676 11764
rect 34732 10016 34772 10025
rect 34732 9680 34772 9976
rect 34732 9631 34772 9640
rect 34636 9547 34676 9556
rect 34540 9295 34580 9304
rect 34732 9512 34772 9521
rect 34444 8791 34484 8800
rect 34540 9176 34580 9185
rect 34252 8756 34292 8765
rect 34252 8672 34292 8716
rect 34252 8621 34292 8632
rect 34156 8464 34484 8504
rect 33772 8168 33812 8464
rect 33928 8336 34296 8345
rect 33968 8296 34010 8336
rect 34050 8296 34092 8336
rect 34132 8296 34174 8336
rect 34214 8296 34256 8336
rect 33928 8287 34296 8296
rect 33772 8119 33812 8128
rect 34348 8168 34388 8177
rect 33772 8000 33812 8009
rect 33772 7328 33812 7960
rect 34252 8000 34292 8009
rect 33964 7748 34004 7757
rect 33964 7412 34004 7708
rect 33964 7363 34004 7372
rect 33772 4556 33812 7288
rect 34252 7244 34292 7960
rect 34252 7195 34292 7204
rect 33928 6824 34296 6833
rect 33968 6784 34010 6824
rect 34050 6784 34092 6824
rect 34132 6784 34174 6824
rect 34214 6784 34256 6824
rect 33928 6775 34296 6784
rect 33928 5312 34296 5321
rect 33968 5272 34010 5312
rect 34050 5272 34092 5312
rect 34132 5272 34174 5312
rect 34214 5272 34256 5312
rect 33928 5263 34296 5272
rect 34348 4808 34388 8128
rect 33772 4507 33812 4516
rect 34252 4768 34388 4808
rect 34252 3968 34292 4768
rect 34348 4640 34388 4649
rect 34348 4220 34388 4600
rect 34348 4171 34388 4180
rect 34252 3919 34292 3928
rect 33928 3800 34296 3809
rect 33968 3760 34010 3800
rect 34050 3760 34092 3800
rect 34132 3760 34174 3800
rect 34214 3760 34256 3800
rect 33928 3751 34296 3760
rect 34444 3548 34484 8464
rect 34540 8168 34580 9136
rect 34732 8840 34772 9472
rect 34828 8924 34868 11764
rect 35020 9680 35060 11764
rect 35020 9631 35060 9640
rect 40492 9848 40532 9857
rect 35404 9596 35444 9605
rect 40396 9596 40436 9605
rect 34828 8875 34868 8884
rect 35020 9512 35060 9521
rect 34732 8791 34772 8800
rect 34732 8672 34772 8681
rect 34540 8119 34580 8128
rect 34636 8336 34676 8345
rect 34636 7580 34676 8296
rect 34732 8168 34772 8632
rect 34732 8119 34772 8128
rect 34924 8588 34964 8597
rect 34636 7531 34676 7540
rect 34828 8084 34868 8093
rect 34828 5396 34868 8044
rect 34924 8000 34964 8548
rect 35020 8504 35060 9472
rect 35404 9461 35444 9556
rect 40300 9556 40396 9596
rect 35692 9512 35732 9521
rect 35168 9092 35536 9101
rect 35208 9052 35250 9092
rect 35290 9052 35332 9092
rect 35372 9052 35414 9092
rect 35454 9052 35496 9092
rect 35168 9043 35536 9052
rect 35596 9092 35636 9103
rect 35596 9008 35636 9052
rect 35596 8959 35636 8968
rect 35308 8672 35348 8681
rect 35308 8537 35348 8632
rect 35020 8455 35060 8464
rect 35692 8084 35732 9472
rect 38860 9512 38900 9521
rect 37804 9428 37844 9437
rect 37708 9344 37748 9353
rect 37612 9304 37708 9344
rect 35788 9260 35828 9269
rect 35788 8252 35828 9220
rect 35980 9176 36020 9185
rect 35980 8336 36020 9136
rect 37612 9176 37652 9304
rect 37708 9295 37748 9304
rect 37612 9127 37652 9136
rect 37228 8924 37268 8933
rect 35980 8287 36020 8296
rect 36652 8504 36692 8513
rect 35788 8203 35828 8212
rect 35692 8035 35732 8044
rect 34924 7951 34964 7960
rect 36076 8000 36116 8009
rect 35980 7748 36020 7757
rect 35020 7580 35060 7591
rect 35020 7496 35060 7540
rect 35168 7580 35536 7589
rect 35208 7540 35250 7580
rect 35290 7540 35332 7580
rect 35372 7540 35414 7580
rect 35454 7540 35496 7580
rect 35168 7531 35536 7540
rect 35596 7580 35636 7589
rect 35020 7447 35060 7456
rect 34924 6824 34964 6833
rect 34924 5984 34964 6784
rect 35168 6068 35536 6077
rect 35208 6028 35250 6068
rect 35290 6028 35332 6068
rect 35372 6028 35414 6068
rect 35454 6028 35496 6068
rect 35168 6019 35536 6028
rect 34924 5935 34964 5944
rect 34828 5347 34868 5356
rect 35168 4556 35536 4565
rect 35208 4516 35250 4556
rect 35290 4516 35332 4556
rect 35372 4516 35414 4556
rect 35454 4516 35496 4556
rect 35168 4507 35536 4516
rect 34444 3499 34484 3508
rect 33676 3163 33716 3172
rect 35168 3044 35536 3053
rect 35208 3004 35250 3044
rect 35290 3004 35332 3044
rect 35372 3004 35414 3044
rect 35454 3004 35496 3044
rect 35168 2995 35536 3004
rect 35596 2900 35636 7540
rect 35980 5060 36020 7708
rect 35980 5011 36020 5020
rect 32428 2071 32468 2080
rect 33196 2860 33332 2900
rect 34636 2860 35636 2900
rect 32236 1567 32276 1576
rect 33196 440 33236 2860
rect 33928 2288 34296 2297
rect 33968 2248 34010 2288
rect 34050 2248 34092 2288
rect 34132 2248 34174 2288
rect 34214 2248 34256 2288
rect 33928 2239 34296 2248
rect 33100 400 33236 440
rect 33100 80 33140 400
rect 34636 80 34676 2860
rect 35168 1532 35536 1541
rect 35208 1492 35250 1532
rect 35290 1492 35332 1532
rect 35372 1492 35414 1532
rect 35454 1492 35496 1532
rect 35168 1483 35536 1492
rect 36076 1196 36116 7960
rect 36652 7916 36692 8464
rect 36652 7867 36692 7876
rect 36460 7832 36500 7841
rect 36268 7748 36308 7757
rect 36460 7748 36500 7792
rect 36748 7832 36788 7841
rect 36748 7748 36788 7792
rect 36460 7708 36788 7748
rect 37132 7748 37172 7757
rect 36076 1147 36116 1156
rect 36172 6992 36212 7001
rect 36172 80 36212 6952
rect 36268 3632 36308 7708
rect 37132 7496 37172 7708
rect 37132 7447 37172 7456
rect 36364 7412 36404 7421
rect 36364 7277 36404 7372
rect 36268 3583 36308 3592
rect 37228 3296 37268 8884
rect 37804 8924 37844 9388
rect 37804 8875 37844 8884
rect 37900 9176 37940 9185
rect 37900 8924 37940 9136
rect 37900 8875 37940 8884
rect 38380 8840 38420 8849
rect 38668 8840 38708 8849
rect 38420 8800 38668 8840
rect 38380 8791 38420 8800
rect 38668 8791 38708 8800
rect 38572 8420 38612 8429
rect 37228 3247 37268 3256
rect 37708 7244 37748 7253
rect 36844 3212 36884 3221
rect 36844 3044 36884 3172
rect 36844 2995 36884 3004
rect 37612 3212 37652 3221
rect 37612 2792 37652 3172
rect 37612 2743 37652 2752
rect 36364 2624 36404 2633
rect 36364 2036 36404 2584
rect 36364 1987 36404 1996
rect 37708 80 37748 7204
rect 38092 7160 38132 7169
rect 37996 6404 38036 6413
rect 38092 6404 38132 7120
rect 38036 6364 38132 6404
rect 38188 6404 38228 6413
rect 37996 6355 38036 6364
rect 38188 5984 38228 6364
rect 38188 5935 38228 5944
rect 38380 4136 38420 4147
rect 38380 4052 38420 4096
rect 38380 4003 38420 4012
rect 38572 3632 38612 8380
rect 38860 8336 38900 9472
rect 40204 9512 40244 9521
rect 40108 9092 40148 9101
rect 39052 8756 39092 8765
rect 38860 8287 38900 8296
rect 38956 8672 38996 8681
rect 38668 8168 38708 8177
rect 38668 7328 38708 8128
rect 38668 7279 38708 7288
rect 38860 4136 38900 4145
rect 38668 3968 38708 3977
rect 38668 3833 38708 3928
rect 38860 3884 38900 4096
rect 38860 3835 38900 3844
rect 38956 3800 38996 8632
rect 39052 4724 39092 8716
rect 39052 4675 39092 4684
rect 39148 4808 39188 4817
rect 38956 3751 38996 3760
rect 38572 3583 38612 3592
rect 38188 3464 38228 3473
rect 38188 3329 38228 3424
rect 38860 3296 38900 3305
rect 38860 1532 38900 3256
rect 38860 1483 38900 1492
rect 39052 3212 39092 3221
rect 39052 1280 39092 3172
rect 39148 2876 39188 4768
rect 39148 2827 39188 2836
rect 39532 3464 39572 3473
rect 39148 2624 39188 2633
rect 39148 1952 39188 2584
rect 39148 1903 39188 1912
rect 39436 2624 39476 2633
rect 39052 1231 39092 1240
rect 39436 1700 39476 2584
rect 39244 1196 39284 1205
rect 39244 80 39284 1156
rect 39436 608 39476 1660
rect 39532 944 39572 3424
rect 40108 3464 40148 9052
rect 40204 4304 40244 9472
rect 40300 8756 40340 9556
rect 40396 9547 40436 9556
rect 40492 9260 40532 9808
rect 40492 9211 40532 9220
rect 41644 9512 41684 9521
rect 40300 8707 40340 8716
rect 40780 8588 40820 8597
rect 40204 4255 40244 4264
rect 40300 7412 40340 7421
rect 40300 4220 40340 7372
rect 40300 4171 40340 4180
rect 40108 3415 40148 3424
rect 40300 3968 40340 3977
rect 39724 3128 39764 3137
rect 39628 2876 39668 2885
rect 39628 2372 39668 2836
rect 39724 2792 39764 3088
rect 39724 2743 39764 2752
rect 40012 2708 40052 2717
rect 39628 2323 39668 2332
rect 39724 2624 39764 2633
rect 39724 1952 39764 2584
rect 40012 2204 40052 2668
rect 40012 2155 40052 2164
rect 40108 2624 40148 2633
rect 39724 1903 39764 1912
rect 40108 1700 40148 2584
rect 40300 1952 40340 3928
rect 40492 2624 40532 2633
rect 40492 2489 40532 2584
rect 40588 2456 40628 2465
rect 40588 2204 40628 2416
rect 40588 2155 40628 2164
rect 40300 1903 40340 1912
rect 40108 1651 40148 1660
rect 39532 895 39572 904
rect 39436 559 39476 568
rect 40780 80 40820 8548
rect 41644 5144 41684 9472
rect 41740 8672 41780 11740
rect 43180 11024 43220 11033
rect 43084 10984 43180 11024
rect 42988 10100 43028 10109
rect 42892 10016 42932 10025
rect 42316 9932 42356 9941
rect 41740 8623 41780 8632
rect 41836 9764 41876 9773
rect 41836 9260 41876 9724
rect 41740 8084 41780 8093
rect 41740 7916 41780 8044
rect 41740 7867 41780 7876
rect 41836 7664 41876 9220
rect 42220 9512 42260 9521
rect 42220 9176 42260 9472
rect 42220 9127 42260 9136
rect 41740 7624 41876 7664
rect 41932 8840 41972 8849
rect 41740 6824 41780 7624
rect 41740 6775 41780 6784
rect 41836 6992 41876 7001
rect 41836 5816 41876 6952
rect 41836 5767 41876 5776
rect 41644 5095 41684 5104
rect 41452 4052 41492 4061
rect 41452 356 41492 4012
rect 41740 3548 41780 3557
rect 41932 3548 41972 8800
rect 42316 8840 42356 9892
rect 42604 9512 42644 9521
rect 42604 9176 42644 9472
rect 42604 9127 42644 9136
rect 42700 9428 42740 9437
rect 42316 8791 42356 8800
rect 42700 8840 42740 9388
rect 42700 8791 42740 8800
rect 42892 8756 42932 9976
rect 42988 9428 43028 10060
rect 43084 9680 43124 10984
rect 43180 10975 43220 10984
rect 43084 9631 43124 9640
rect 44044 10688 44084 10697
rect 44044 9680 44084 10648
rect 44428 10352 44468 10361
rect 44044 9631 44084 9640
rect 44140 9848 44180 9857
rect 43564 9596 43604 9605
rect 42988 9388 43124 9428
rect 42892 8707 42932 8716
rect 42988 9008 43028 9017
rect 42988 8672 43028 8968
rect 43084 8840 43124 9388
rect 43468 9260 43508 9269
rect 43468 9125 43508 9220
rect 43084 8791 43124 8800
rect 43564 8756 43604 9556
rect 43564 8707 43604 8716
rect 42988 8623 43028 8632
rect 44140 8672 44180 9808
rect 44428 9680 44468 10312
rect 44428 9631 44468 9640
rect 44524 10016 44564 10025
rect 44524 8924 44564 9976
rect 44908 9512 44948 9521
rect 44908 9344 44948 9472
rect 44908 9295 44948 9304
rect 44524 8875 44564 8884
rect 44140 8623 44180 8632
rect 44908 8756 44948 8767
rect 44908 8672 44948 8716
rect 44908 8623 44948 8632
rect 42892 8588 42932 8597
rect 42028 8084 42068 8093
rect 42028 7580 42068 8044
rect 42124 7748 42164 7757
rect 42124 7613 42164 7708
rect 42028 7531 42068 7540
rect 42028 7244 42068 7253
rect 42028 6572 42068 7204
rect 42124 7160 42164 7169
rect 42124 6656 42164 7120
rect 42124 6607 42164 6616
rect 42604 6992 42644 7001
rect 42028 6523 42068 6532
rect 42316 6488 42356 6497
rect 42316 6236 42356 6448
rect 42316 6187 42356 6196
rect 42604 5900 42644 6952
rect 42604 5851 42644 5860
rect 41780 3508 41876 3548
rect 41740 3499 41780 3508
rect 41644 3296 41684 3305
rect 41644 1868 41684 3256
rect 41836 3296 41876 3508
rect 41932 3499 41972 3508
rect 42316 5396 42356 5405
rect 41836 3247 41876 3256
rect 41644 1819 41684 1828
rect 41740 3212 41780 3221
rect 41740 1784 41780 3172
rect 41740 1735 41780 1744
rect 42028 2456 42068 2465
rect 42028 1616 42068 2416
rect 42028 1567 42068 1576
rect 41452 307 41492 316
rect 42316 80 42356 5356
rect 42892 5228 42932 8548
rect 45772 8504 45812 8513
rect 44524 8000 44564 8009
rect 43276 7916 43316 7925
rect 43084 7160 43124 7169
rect 43084 6320 43124 7120
rect 43084 6271 43124 6280
rect 42892 5179 42932 5188
rect 43180 4892 43220 4901
rect 43084 4852 43180 4892
rect 42988 4136 43028 4145
rect 42988 4001 43028 4096
rect 42988 3884 43028 3893
rect 42892 3844 42988 3884
rect 42892 3044 42932 3844
rect 42988 3835 43028 3844
rect 43084 3716 43124 4852
rect 43180 4843 43220 4852
rect 43180 3968 43220 3977
rect 43180 3833 43220 3928
rect 43084 3667 43124 3676
rect 42892 2995 42932 3004
rect 42988 3464 43028 3473
rect 42988 104 43028 3424
rect 43084 3380 43124 3389
rect 43084 2288 43124 3340
rect 43084 2239 43124 2248
rect 13172 64 13192 80
rect 13112 0 13192 64
rect 14648 0 14728 80
rect 16184 0 16264 80
rect 17720 0 17800 80
rect 19256 0 19336 80
rect 20792 0 20872 80
rect 22328 0 22408 80
rect 23864 0 23944 80
rect 25400 0 25480 80
rect 26936 0 27016 80
rect 28472 0 28552 80
rect 30008 0 30088 80
rect 31544 0 31624 80
rect 33080 0 33160 80
rect 34616 0 34696 80
rect 36152 0 36232 80
rect 37688 0 37768 80
rect 39224 0 39304 80
rect 40760 0 40840 80
rect 42296 0 42376 80
rect 42988 55 43028 64
rect 43276 60 43316 7876
rect 43468 7832 43508 7841
rect 43468 7697 43508 7792
rect 44524 7664 44564 7960
rect 44908 8000 44948 8009
rect 44908 7865 44948 7960
rect 45772 8000 45812 8464
rect 45772 7951 45812 7960
rect 44524 7615 44564 7624
rect 45964 7748 46004 7757
rect 44908 7328 44948 7337
rect 43468 7160 43508 7169
rect 43468 6320 43508 7120
rect 43468 6271 43508 6280
rect 43660 7160 43700 7169
rect 43660 6236 43700 7120
rect 43660 5648 43700 6196
rect 44236 7160 44276 7169
rect 44236 6152 44276 7120
rect 44236 6103 44276 6112
rect 43660 4892 43700 5608
rect 43660 4843 43700 4852
rect 43948 5648 43988 5657
rect 43948 4724 43988 5608
rect 43948 4388 43988 4684
rect 43468 4136 43508 4145
rect 43372 3464 43412 3473
rect 43372 3296 43412 3424
rect 43372 3247 43412 3256
rect 43372 2540 43412 2549
rect 43372 2036 43412 2500
rect 43372 1987 43412 1996
rect 43468 188 43508 4096
rect 43756 4136 43796 4145
rect 43756 2900 43796 4096
rect 43660 2860 43796 2900
rect 43660 272 43700 2860
rect 43948 2120 43988 4348
rect 44524 3464 44564 3473
rect 44524 2876 44564 3424
rect 44524 2827 44564 2836
rect 43948 2071 43988 2080
rect 44332 2624 44372 2633
rect 44332 2036 44372 2584
rect 44908 2624 44948 7288
rect 45964 7328 46004 7708
rect 45964 7279 46004 7288
rect 45196 6320 45236 6329
rect 45196 5648 45236 6280
rect 46252 6152 46292 6161
rect 46252 5984 46292 6112
rect 46252 5935 46292 5944
rect 45196 5599 45236 5608
rect 45388 5648 45428 5657
rect 45388 5144 45428 5608
rect 45388 5095 45428 5104
rect 45772 4976 45812 4985
rect 45772 4304 45812 4936
rect 45772 4255 45812 4264
rect 45964 4304 46004 4313
rect 45964 3632 46004 4264
rect 45964 3583 46004 3592
rect 46156 3632 46196 3641
rect 44908 2575 44948 2584
rect 45484 2960 45524 2969
rect 45484 2120 45524 2920
rect 46156 2876 46196 3592
rect 46156 2827 46196 2836
rect 45484 2071 45524 2080
rect 44332 1987 44372 1996
rect 43852 1868 43892 1877
rect 43756 1532 43796 1541
rect 43852 1532 43892 1828
rect 45676 1784 45716 1793
rect 43796 1492 43892 1532
rect 44620 1700 44660 1709
rect 43756 1483 43796 1492
rect 44620 608 44660 1660
rect 45676 944 45716 1744
rect 46252 1448 46292 1457
rect 46252 1280 46292 1408
rect 46252 1231 46292 1240
rect 45676 895 45716 904
rect 44620 559 44660 568
rect 43660 223 43700 232
rect 43468 139 43508 148
rect 43660 104 43700 113
rect 43852 104 43892 113
rect 43660 60 43700 64
rect 43276 20 43700 60
rect 43832 64 43852 80
rect 43892 64 43912 80
rect 43832 0 43912 64
<< via3 >>
rect 652 3592 692 3632
rect 460 3424 500 3464
rect 4300 11740 4340 11780
rect 3688 9808 3728 9848
rect 3770 9808 3810 9848
rect 3852 9808 3892 9848
rect 3934 9808 3974 9848
rect 4016 9808 4056 9848
rect 3688 8296 3728 8336
rect 3770 8296 3810 8336
rect 3852 8296 3892 8336
rect 3934 8296 3974 8336
rect 4016 8296 4056 8336
rect 3244 8212 3284 8252
rect 4928 9052 4968 9092
rect 5010 9052 5050 9092
rect 5092 9052 5132 9092
rect 5174 9052 5214 9092
rect 5256 9052 5296 9092
rect 4928 7540 4968 7580
rect 5010 7540 5050 7580
rect 5092 7540 5132 7580
rect 5174 7540 5214 7580
rect 5256 7540 5296 7580
rect 3688 6784 3728 6824
rect 3770 6784 3810 6824
rect 3852 6784 3892 6824
rect 3934 6784 3974 6824
rect 4016 6784 4056 6824
rect 4928 6028 4968 6068
rect 5010 6028 5050 6068
rect 5092 6028 5132 6068
rect 5174 6028 5214 6068
rect 5256 6028 5296 6068
rect 3688 5272 3728 5312
rect 3770 5272 3810 5312
rect 3852 5272 3892 5312
rect 3934 5272 3974 5312
rect 4016 5272 4056 5312
rect 4928 4516 4968 4556
rect 5010 4516 5050 4556
rect 5092 4516 5132 4556
rect 5174 4516 5214 4556
rect 5256 4516 5296 4556
rect 2188 4180 2228 4220
rect 3688 3760 3728 3800
rect 3770 3760 3810 3800
rect 3852 3760 3892 3800
rect 3934 3760 3974 3800
rect 4016 3760 4056 3800
rect 1804 3340 1844 3380
rect 4928 3004 4968 3044
rect 5010 3004 5050 3044
rect 5092 3004 5132 3044
rect 5174 3004 5214 3044
rect 5256 3004 5296 3044
rect 1420 2584 1460 2624
rect 9292 9220 9332 9260
rect 7852 8212 7892 8252
rect 3688 2248 3728 2288
rect 3770 2248 3810 2288
rect 3852 2248 3892 2288
rect 3934 2248 3974 2288
rect 4016 2248 4056 2288
rect 10060 9892 10100 9932
rect 10156 9724 10196 9764
rect 9868 9136 9908 9176
rect 9964 7288 10004 7328
rect 10540 8716 10580 8756
rect 10636 6196 10676 6236
rect 11020 8548 11060 8588
rect 11212 8632 11252 8672
rect 10828 5020 10868 5060
rect 11212 7624 11252 7664
rect 11116 6364 11156 6404
rect 11884 9976 11924 10016
rect 11596 7624 11636 7664
rect 11596 7456 11636 7496
rect 11500 7120 11540 7160
rect 11596 6364 11636 6404
rect 12460 9472 12500 9512
rect 12076 8800 12116 8840
rect 12844 9808 12884 9848
rect 12172 7540 12212 7580
rect 11980 7288 12020 7328
rect 11788 6952 11828 6992
rect 11884 6868 11924 6908
rect 12172 7204 12212 7244
rect 12556 7624 12596 7664
rect 12460 7372 12500 7412
rect 12556 7288 12596 7328
rect 12460 7036 12500 7076
rect 12940 9556 12980 9596
rect 13132 9556 13172 9596
rect 13420 9472 13460 9512
rect 13612 9472 13652 9512
rect 13900 9052 13940 9092
rect 12844 8212 12884 8252
rect 13036 7456 13076 7496
rect 12748 7288 12788 7328
rect 12748 6868 12788 6908
rect 13132 7204 13172 7244
rect 12940 7036 12980 7076
rect 13132 6952 13172 6992
rect 14092 9052 14132 9092
rect 14092 7708 14132 7748
rect 14956 9640 14996 9680
rect 14668 9472 14708 9512
rect 15148 9808 15188 9848
rect 14380 6196 14420 6236
rect 4928 1492 4968 1532
rect 5010 1492 5050 1532
rect 5092 1492 5132 1532
rect 5174 1492 5214 1532
rect 5256 1492 5296 1532
rect 15052 8632 15092 8672
rect 15532 9472 15572 9512
rect 15532 7876 15572 7916
rect 15916 7792 15956 7832
rect 15436 7540 15476 7580
rect 15052 3256 15092 3296
rect 16204 8212 16244 8252
rect 16300 7960 16340 8000
rect 17548 8716 17588 8756
rect 17356 6448 17396 6488
rect 17932 7624 17972 7664
rect 16876 3256 16916 3296
rect 19180 10060 19220 10100
rect 18808 9808 18848 9848
rect 18890 9808 18930 9848
rect 18972 9808 19012 9848
rect 19054 9808 19094 9848
rect 19136 9808 19176 9848
rect 19180 9640 19220 9680
rect 19084 9556 19124 9596
rect 19180 9304 19220 9344
rect 19180 8884 19220 8924
rect 19372 9388 19412 9428
rect 19372 8968 19412 9008
rect 19564 9640 19604 9680
rect 19564 9472 19604 9512
rect 19852 10480 19892 10520
rect 20044 9976 20084 10016
rect 19852 9640 19892 9680
rect 20044 9640 20084 9680
rect 19660 9388 19700 9428
rect 19564 9052 19604 9092
rect 18808 8296 18848 8336
rect 18890 8296 18930 8336
rect 18972 8296 19012 8336
rect 19054 8296 19094 8336
rect 19136 8296 19176 8336
rect 20048 9052 20088 9092
rect 20130 9052 20170 9092
rect 20212 9052 20252 9092
rect 20294 9052 20334 9092
rect 20376 9052 20416 9092
rect 19852 8884 19892 8924
rect 20236 8800 20276 8840
rect 19756 7120 19796 7160
rect 18808 6784 18848 6824
rect 18890 6784 18930 6824
rect 18972 6784 19012 6824
rect 19054 6784 19094 6824
rect 19136 6784 19176 6824
rect 19948 8632 19988 8672
rect 20140 8548 20180 8588
rect 20140 8128 20180 8168
rect 20048 7540 20088 7580
rect 20130 7540 20170 7580
rect 20212 7540 20252 7580
rect 20294 7540 20334 7580
rect 20376 7540 20416 7580
rect 20140 7372 20180 7412
rect 20048 6028 20088 6068
rect 20130 6028 20170 6068
rect 20212 6028 20252 6068
rect 20294 6028 20334 6068
rect 20376 6028 20416 6068
rect 18808 5272 18848 5312
rect 18890 5272 18930 5312
rect 18972 5272 19012 5312
rect 19054 5272 19094 5312
rect 19136 5272 19176 5312
rect 20048 4516 20088 4556
rect 20130 4516 20170 4556
rect 20212 4516 20252 4556
rect 20294 4516 20334 4556
rect 20376 4516 20416 4556
rect 19756 4348 19796 4388
rect 19180 3928 19220 3968
rect 18808 3760 18848 3800
rect 18890 3760 18930 3800
rect 18972 3760 19012 3800
rect 19054 3760 19094 3800
rect 19136 3760 19176 3800
rect 18220 3172 18260 3212
rect 19372 3508 19412 3548
rect 18796 3172 18836 3212
rect 19660 2752 19700 2792
rect 20048 3004 20088 3044
rect 20130 3004 20170 3044
rect 20212 3004 20252 3044
rect 20294 3004 20334 3044
rect 20376 3004 20416 3044
rect 20812 8968 20852 9008
rect 21100 9808 21140 9848
rect 21100 4264 21140 4304
rect 20716 2752 20756 2792
rect 20812 4096 20852 4136
rect 18808 2248 18848 2288
rect 18890 2248 18930 2288
rect 18972 2248 19012 2288
rect 19054 2248 19094 2288
rect 19136 2248 19176 2288
rect 20048 1492 20088 1532
rect 20130 1492 20170 1532
rect 20212 1492 20252 1532
rect 20294 1492 20334 1532
rect 20376 1492 20416 1532
rect 21292 8884 21332 8924
rect 21676 8800 21716 8840
rect 21484 8632 21524 8672
rect 23308 11740 23348 11780
rect 22156 9052 22196 9092
rect 21484 3676 21524 3716
rect 22828 9052 22868 9092
rect 22924 9304 22964 9344
rect 21964 4264 22004 4304
rect 21772 3928 21812 3968
rect 21580 3256 21620 3296
rect 21772 3676 21812 3716
rect 23116 8968 23156 9008
rect 23308 8800 23348 8840
rect 23980 9640 24020 9680
rect 23692 9052 23732 9092
rect 24364 9640 24404 9680
rect 21964 3172 22004 3212
rect 24364 3508 24404 3548
rect 24460 9052 24500 9092
rect 24172 3088 24212 3128
rect 25036 9052 25076 9092
rect 25036 8884 25076 8924
rect 24940 8632 24980 8672
rect 25036 3508 25076 3548
rect 26284 9640 26324 9680
rect 26572 8632 26612 8672
rect 26764 8548 26804 8588
rect 27052 9052 27092 9092
rect 27148 8884 27188 8924
rect 27052 8800 27092 8840
rect 27436 10312 27476 10352
rect 27052 5020 27092 5060
rect 26956 3256 26996 3296
rect 25612 3088 25652 3128
rect 26860 2920 26900 2960
rect 22924 1744 22964 1784
rect 28204 8128 28244 8168
rect 27436 3508 27476 3548
rect 27628 3340 27668 3380
rect 29644 11740 29684 11780
rect 30316 8548 30356 8588
rect 30892 8968 30932 9008
rect 30028 4180 30068 4220
rect 31468 8380 31508 8420
rect 31564 4180 31604 4220
rect 27340 2920 27380 2960
rect 31948 8884 31988 8924
rect 32044 4012 32084 4052
rect 30220 2164 30260 2204
rect 30220 1744 30260 1784
rect 33100 8632 33140 8672
rect 33484 8968 33524 9008
rect 33868 9976 33908 10016
rect 34252 10144 34292 10184
rect 33928 9808 33968 9848
rect 34010 9808 34050 9848
rect 34092 9808 34132 9848
rect 34174 9808 34214 9848
rect 34256 9808 34296 9848
rect 33772 9472 33812 9512
rect 33292 8212 33332 8252
rect 33388 8632 33428 8672
rect 33004 8044 33044 8084
rect 33292 8044 33332 8084
rect 32812 6448 32852 6488
rect 32524 4180 32564 4220
rect 33100 7540 33140 7580
rect 33004 4180 33044 4220
rect 33196 4180 33236 4220
rect 33004 3844 33044 3884
rect 33580 8464 33620 8504
rect 33580 8212 33620 8252
rect 33580 8044 33620 8084
rect 34540 10144 34580 10184
rect 34732 9976 34772 10016
rect 34636 9556 34676 9596
rect 34252 8632 34292 8672
rect 33928 8296 33968 8336
rect 34010 8296 34050 8336
rect 34092 8296 34132 8336
rect 34174 8296 34214 8336
rect 34256 8296 34296 8336
rect 34348 8128 34388 8168
rect 33964 7372 34004 7412
rect 33928 6784 33968 6824
rect 34010 6784 34050 6824
rect 34092 6784 34132 6824
rect 34174 6784 34214 6824
rect 34256 6784 34296 6824
rect 33928 5272 33968 5312
rect 34010 5272 34050 5312
rect 34092 5272 34132 5312
rect 34174 5272 34214 5312
rect 34256 5272 34296 5312
rect 33928 3760 33968 3800
rect 34010 3760 34050 3800
rect 34092 3760 34132 3800
rect 34174 3760 34214 3800
rect 34256 3760 34296 3800
rect 41740 11740 41780 11780
rect 35404 9556 35444 9596
rect 34636 7540 34676 7580
rect 34828 8044 34868 8084
rect 35168 9052 35208 9092
rect 35250 9052 35290 9092
rect 35332 9052 35372 9092
rect 35414 9052 35454 9092
rect 35496 9052 35536 9092
rect 35596 8968 35636 9008
rect 35308 8632 35348 8672
rect 36652 8464 36692 8504
rect 35788 8212 35828 8252
rect 35168 7540 35208 7580
rect 35250 7540 35290 7580
rect 35332 7540 35372 7580
rect 35414 7540 35454 7580
rect 35496 7540 35536 7580
rect 35020 7456 35060 7496
rect 35168 6028 35208 6068
rect 35250 6028 35290 6068
rect 35332 6028 35372 6068
rect 35414 6028 35454 6068
rect 35496 6028 35536 6068
rect 34828 5356 34868 5396
rect 35168 4516 35208 4556
rect 35250 4516 35290 4556
rect 35332 4516 35372 4556
rect 35414 4516 35454 4556
rect 35496 4516 35536 4556
rect 35168 3004 35208 3044
rect 35250 3004 35290 3044
rect 35332 3004 35372 3044
rect 35414 3004 35454 3044
rect 35496 3004 35536 3044
rect 33928 2248 33968 2288
rect 34010 2248 34050 2288
rect 34092 2248 34132 2288
rect 34174 2248 34214 2288
rect 34256 2248 34296 2288
rect 35168 1492 35208 1532
rect 35250 1492 35290 1532
rect 35332 1492 35372 1532
rect 35414 1492 35454 1532
rect 35496 1492 35536 1532
rect 36076 1156 36116 1196
rect 37132 7456 37172 7496
rect 36364 7372 36404 7412
rect 36268 3592 36308 3632
rect 37804 8884 37844 8924
rect 38572 8380 38612 8420
rect 38380 4012 38420 4052
rect 40204 9472 40244 9512
rect 38668 3928 38708 3968
rect 38860 3844 38900 3884
rect 38188 3424 38228 3464
rect 39244 1156 39284 1196
rect 40012 2164 40052 2204
rect 40492 2584 40532 2624
rect 41740 7876 41780 7916
rect 42604 9136 42644 9176
rect 42700 9388 42740 9428
rect 43468 9220 43508 9260
rect 44908 9304 44948 9344
rect 44908 8716 44948 8756
rect 42124 7708 42164 7748
rect 42316 5356 42356 5396
rect 42988 4096 43028 4136
rect 43180 3928 43220 3968
rect 43468 7792 43508 7832
rect 44908 7960 44948 8000
rect 44524 7624 44564 7664
rect 43372 3256 43412 3296
rect 43660 64 43700 104
rect 43852 64 43892 104
<< metal4 >>
rect 4291 11740 4300 11780
rect 4340 11740 23308 11780
rect 23348 11740 23357 11780
rect 29635 11740 29644 11780
rect 29684 11740 41740 11780
rect 41780 11740 41789 11780
rect 19757 10480 19852 10520
rect 19892 10480 19901 10520
rect 19459 10312 19468 10352
rect 19508 10312 27436 10352
rect 27476 10312 27485 10352
rect 19747 10228 19756 10268
rect 19796 10228 20084 10268
rect 19171 10060 19180 10100
rect 19220 10060 19229 10100
rect 19180 10016 19220 10060
rect 20044 10016 20084 10228
rect 34243 10144 34252 10184
rect 34292 10144 34540 10184
rect 34580 10144 34589 10184
rect 11875 9976 11884 10016
rect 11924 9976 19220 10016
rect 20035 9976 20044 10016
rect 20084 9976 20093 10016
rect 33859 9976 33868 10016
rect 33908 9976 34732 10016
rect 34772 9976 34781 10016
rect 10051 9892 10060 9932
rect 10100 9892 19660 9932
rect 19700 9892 19709 9932
rect 3679 9808 3688 9848
rect 3728 9808 3770 9848
rect 3810 9808 3852 9848
rect 3892 9808 3934 9848
rect 3974 9808 4016 9848
rect 4056 9808 4065 9848
rect 12835 9808 12844 9848
rect 12884 9808 15148 9848
rect 15188 9808 15197 9848
rect 18799 9808 18808 9848
rect 18848 9808 18890 9848
rect 18930 9808 18972 9848
rect 19012 9808 19054 9848
rect 19094 9808 19136 9848
rect 19176 9808 19185 9848
rect 20044 9808 21100 9848
rect 21140 9808 21149 9848
rect 33919 9808 33928 9848
rect 33968 9808 34010 9848
rect 34050 9808 34092 9848
rect 34132 9808 34174 9848
rect 34214 9808 34256 9848
rect 34296 9808 34305 9848
rect 20044 9764 20084 9808
rect 10147 9724 10156 9764
rect 10196 9724 19468 9764
rect 19508 9724 19517 9764
rect 19651 9724 19660 9764
rect 19700 9724 20084 9764
rect 14947 9640 14956 9680
rect 14996 9640 19180 9680
rect 19220 9640 19229 9680
rect 19555 9640 19564 9680
rect 19604 9640 19852 9680
rect 19892 9640 19901 9680
rect 20035 9640 20044 9680
rect 20084 9640 23980 9680
rect 24020 9640 24029 9680
rect 24355 9640 24364 9680
rect 24404 9640 26284 9680
rect 26324 9640 26333 9680
rect 12931 9556 12940 9596
rect 12980 9556 13132 9596
rect 13172 9556 13181 9596
rect 19075 9556 19084 9596
rect 19124 9556 19756 9596
rect 19796 9556 19805 9596
rect 34627 9556 34636 9596
rect 34676 9556 35404 9596
rect 35444 9556 35453 9596
rect 12451 9472 12460 9512
rect 12500 9472 13420 9512
rect 13460 9472 13469 9512
rect 13603 9472 13612 9512
rect 13652 9472 14668 9512
rect 14708 9472 14717 9512
rect 15523 9472 15532 9512
rect 15572 9472 19564 9512
rect 19604 9472 19613 9512
rect 33763 9472 33772 9512
rect 33812 9472 40204 9512
rect 40244 9472 40253 9512
rect 19363 9388 19372 9428
rect 19412 9388 19660 9428
rect 19700 9388 19709 9428
rect 19996 9388 42700 9428
rect 42740 9388 42749 9428
rect 19996 9344 20036 9388
rect 19171 9304 19180 9344
rect 19220 9304 20036 9344
rect 22915 9304 22924 9344
rect 22964 9304 44908 9344
rect 44948 9304 44957 9344
rect 9283 9220 9292 9260
rect 9332 9220 43468 9260
rect 43508 9220 43517 9260
rect 9859 9136 9868 9176
rect 9908 9136 42604 9176
rect 42644 9136 42653 9176
rect 4919 9052 4928 9092
rect 4968 9052 5010 9092
rect 5050 9052 5092 9092
rect 5132 9052 5174 9092
rect 5214 9052 5256 9092
rect 5296 9052 5305 9092
rect 13891 9052 13900 9092
rect 13940 9052 14092 9092
rect 14132 9052 14141 9092
rect 19555 9052 19564 9092
rect 19604 9052 19756 9092
rect 19796 9052 19805 9092
rect 20039 9052 20048 9092
rect 20088 9052 20130 9092
rect 20170 9052 20212 9092
rect 20252 9052 20294 9092
rect 20334 9052 20376 9092
rect 20416 9052 20425 9092
rect 22147 9052 22156 9092
rect 22196 9052 22828 9092
rect 22868 9052 22877 9092
rect 23683 9052 23692 9092
rect 23732 9052 24460 9092
rect 24500 9052 24509 9092
rect 25027 9052 25036 9092
rect 25076 9052 27052 9092
rect 27092 9052 27101 9092
rect 35159 9052 35168 9092
rect 35208 9052 35250 9092
rect 35290 9052 35332 9092
rect 35372 9052 35414 9092
rect 35454 9052 35496 9092
rect 35536 9052 35545 9092
rect 19363 8968 19372 9008
rect 19412 8968 20812 9008
rect 20852 8968 20861 9008
rect 23107 8968 23116 9008
rect 23156 8968 30892 9008
rect 30932 8968 30941 9008
rect 33475 8968 33484 9008
rect 33524 8968 35596 9008
rect 35636 8968 35645 9008
rect 19171 8884 19180 8924
rect 19220 8884 19852 8924
rect 19892 8884 19901 8924
rect 20140 8884 21292 8924
rect 21332 8884 21341 8924
rect 25027 8884 25036 8924
rect 25076 8884 27148 8924
rect 27188 8884 27197 8924
rect 31939 8884 31948 8924
rect 31988 8884 37804 8924
rect 37844 8884 37853 8924
rect 12067 8800 12076 8840
rect 12116 8800 17684 8840
rect 17644 8756 17684 8800
rect 20140 8756 20180 8884
rect 20227 8800 20236 8840
rect 20276 8800 21676 8840
rect 21716 8800 21725 8840
rect 23299 8800 23308 8840
rect 23348 8800 27052 8840
rect 27092 8800 27101 8840
rect 10531 8716 10540 8756
rect 10580 8716 17548 8756
rect 17588 8716 17597 8756
rect 17644 8716 20180 8756
rect 23020 8716 44908 8756
rect 44948 8716 44957 8756
rect 23020 8672 23060 8716
rect 11203 8632 11212 8672
rect 11252 8632 15052 8672
rect 15092 8632 15101 8672
rect 19843 8632 19852 8672
rect 19892 8632 19948 8672
rect 19988 8632 19997 8672
rect 21475 8632 21484 8672
rect 21524 8632 23060 8672
rect 24931 8632 24940 8672
rect 24980 8632 26572 8672
rect 26612 8632 26621 8672
rect 33091 8632 33100 8672
rect 33140 8632 33388 8672
rect 33428 8632 33437 8672
rect 34243 8632 34252 8672
rect 34292 8632 35308 8672
rect 35348 8632 35357 8672
rect 11011 8548 11020 8588
rect 11060 8548 20140 8588
rect 20180 8548 20189 8588
rect 26755 8548 26764 8588
rect 26804 8548 30316 8588
rect 30356 8548 30365 8588
rect 33571 8464 33580 8504
rect 33620 8464 36652 8504
rect 36692 8464 36701 8504
rect 31459 8380 31468 8420
rect 31508 8380 38572 8420
rect 38612 8380 38621 8420
rect 3679 8296 3688 8336
rect 3728 8296 3770 8336
rect 3810 8296 3852 8336
rect 3892 8296 3934 8336
rect 3974 8296 4016 8336
rect 4056 8296 4065 8336
rect 18799 8296 18808 8336
rect 18848 8296 18890 8336
rect 18930 8296 18972 8336
rect 19012 8296 19054 8336
rect 19094 8296 19136 8336
rect 19176 8296 19185 8336
rect 33919 8296 33928 8336
rect 33968 8296 34010 8336
rect 34050 8296 34092 8336
rect 34132 8296 34174 8336
rect 34214 8296 34256 8336
rect 34296 8296 34305 8336
rect 3235 8212 3244 8252
rect 3284 8212 7852 8252
rect 7892 8212 7901 8252
rect 12835 8212 12844 8252
rect 12884 8212 16204 8252
rect 16244 8212 16253 8252
rect 33283 8212 33292 8252
rect 33332 8212 33341 8252
rect 33571 8212 33580 8252
rect 33620 8212 35788 8252
rect 35828 8212 35837 8252
rect 33292 8168 33332 8212
rect 20131 8128 20140 8168
rect 20180 8128 28204 8168
rect 28244 8128 28253 8168
rect 33292 8128 34348 8168
rect 34388 8128 34397 8168
rect 32995 8044 33004 8084
rect 33044 8044 33292 8084
rect 33332 8044 33341 8084
rect 33571 8044 33580 8084
rect 33620 8044 34828 8084
rect 34868 8044 34877 8084
rect 16291 7960 16300 8000
rect 16340 7960 44908 8000
rect 44948 7960 44957 8000
rect 15523 7876 15532 7916
rect 15572 7876 41740 7916
rect 41780 7876 41789 7916
rect 15907 7792 15916 7832
rect 15956 7792 43468 7832
rect 43508 7792 43517 7832
rect 14083 7708 14092 7748
rect 14132 7708 42124 7748
rect 42164 7708 42173 7748
rect 11203 7624 11212 7664
rect 11252 7624 11596 7664
rect 11636 7624 12556 7664
rect 12596 7624 12605 7664
rect 17923 7624 17932 7664
rect 17972 7624 44524 7664
rect 44564 7624 44573 7664
rect 4919 7540 4928 7580
rect 4968 7540 5010 7580
rect 5050 7540 5092 7580
rect 5132 7540 5174 7580
rect 5214 7540 5256 7580
rect 5296 7540 5305 7580
rect 12163 7540 12172 7580
rect 12212 7540 15436 7580
rect 15476 7540 15485 7580
rect 20039 7540 20048 7580
rect 20088 7540 20130 7580
rect 20170 7540 20212 7580
rect 20252 7540 20294 7580
rect 20334 7540 20376 7580
rect 20416 7540 20425 7580
rect 33091 7540 33100 7580
rect 33140 7540 34636 7580
rect 34676 7540 34685 7580
rect 35159 7540 35168 7580
rect 35208 7540 35250 7580
rect 35290 7540 35332 7580
rect 35372 7540 35414 7580
rect 35454 7540 35496 7580
rect 35536 7540 35545 7580
rect 11587 7456 11596 7496
rect 11636 7456 13036 7496
rect 13076 7456 13085 7496
rect 35011 7456 35020 7496
rect 35060 7456 37132 7496
rect 37172 7456 37181 7496
rect 12451 7372 12460 7412
rect 12500 7372 20140 7412
rect 20180 7372 20189 7412
rect 33955 7372 33964 7412
rect 34004 7372 36364 7412
rect 36404 7372 36413 7412
rect 9955 7288 9964 7328
rect 10004 7288 11980 7328
rect 12020 7288 12029 7328
rect 12547 7288 12556 7328
rect 12596 7288 12748 7328
rect 12788 7288 12797 7328
rect 12163 7204 12172 7244
rect 12212 7204 13132 7244
rect 13172 7204 13181 7244
rect 11491 7120 11500 7160
rect 11540 7120 19756 7160
rect 19796 7120 19805 7160
rect 12451 7036 12460 7076
rect 12500 7036 12940 7076
rect 12980 7036 12989 7076
rect 11779 6952 11788 6992
rect 11828 6952 13132 6992
rect 13172 6952 13181 6992
rect 11875 6868 11884 6908
rect 11924 6868 12748 6908
rect 12788 6868 12797 6908
rect 3679 6784 3688 6824
rect 3728 6784 3770 6824
rect 3810 6784 3852 6824
rect 3892 6784 3934 6824
rect 3974 6784 4016 6824
rect 4056 6784 4065 6824
rect 18799 6784 18808 6824
rect 18848 6784 18890 6824
rect 18930 6784 18972 6824
rect 19012 6784 19054 6824
rect 19094 6784 19136 6824
rect 19176 6784 19185 6824
rect 33919 6784 33928 6824
rect 33968 6784 34010 6824
rect 34050 6784 34092 6824
rect 34132 6784 34174 6824
rect 34214 6784 34256 6824
rect 34296 6784 34305 6824
rect 17347 6448 17356 6488
rect 17396 6448 32812 6488
rect 32852 6448 32861 6488
rect 11107 6364 11116 6404
rect 11156 6364 11596 6404
rect 11636 6364 11645 6404
rect 10627 6196 10636 6236
rect 10676 6196 14380 6236
rect 14420 6196 14429 6236
rect 4919 6028 4928 6068
rect 4968 6028 5010 6068
rect 5050 6028 5092 6068
rect 5132 6028 5174 6068
rect 5214 6028 5256 6068
rect 5296 6028 5305 6068
rect 20039 6028 20048 6068
rect 20088 6028 20130 6068
rect 20170 6028 20212 6068
rect 20252 6028 20294 6068
rect 20334 6028 20376 6068
rect 20416 6028 20425 6068
rect 35159 6028 35168 6068
rect 35208 6028 35250 6068
rect 35290 6028 35332 6068
rect 35372 6028 35414 6068
rect 35454 6028 35496 6068
rect 35536 6028 35545 6068
rect 34819 5356 34828 5396
rect 34868 5356 42316 5396
rect 42356 5356 42365 5396
rect 3679 5272 3688 5312
rect 3728 5272 3770 5312
rect 3810 5272 3852 5312
rect 3892 5272 3934 5312
rect 3974 5272 4016 5312
rect 4056 5272 4065 5312
rect 18799 5272 18808 5312
rect 18848 5272 18890 5312
rect 18930 5272 18972 5312
rect 19012 5272 19054 5312
rect 19094 5272 19136 5312
rect 19176 5272 19185 5312
rect 33919 5272 33928 5312
rect 33968 5272 34010 5312
rect 34050 5272 34092 5312
rect 34132 5272 34174 5312
rect 34214 5272 34256 5312
rect 34296 5272 34305 5312
rect 10819 5020 10828 5060
rect 10868 5020 27052 5060
rect 27092 5020 27101 5060
rect 4919 4516 4928 4556
rect 4968 4516 5010 4556
rect 5050 4516 5092 4556
rect 5132 4516 5174 4556
rect 5214 4516 5256 4556
rect 5296 4516 5305 4556
rect 20039 4516 20048 4556
rect 20088 4516 20130 4556
rect 20170 4516 20212 4556
rect 20252 4516 20294 4556
rect 20334 4516 20376 4556
rect 20416 4516 20425 4556
rect 35159 4516 35168 4556
rect 35208 4516 35250 4556
rect 35290 4516 35332 4556
rect 35372 4516 35414 4556
rect 35454 4516 35496 4556
rect 35536 4516 35545 4556
rect 19661 4348 19756 4388
rect 19796 4348 19805 4388
rect 21091 4264 21100 4304
rect 21140 4264 21964 4304
rect 22004 4264 22013 4304
rect 2179 4180 2188 4220
rect 2228 4180 30028 4220
rect 30068 4180 30077 4220
rect 31555 4180 31564 4220
rect 31604 4180 32524 4220
rect 32564 4180 32573 4220
rect 32995 4180 33004 4220
rect 33044 4180 33196 4220
rect 33236 4180 33245 4220
rect 20803 4096 20812 4136
rect 20852 4096 42988 4136
rect 43028 4096 43037 4136
rect 32035 4012 32044 4052
rect 32084 4012 38380 4052
rect 38420 4012 38429 4052
rect 19171 3928 19180 3968
rect 19220 3928 21772 3968
rect 21812 3928 21821 3968
rect 38659 3928 38668 3968
rect 38708 3928 43180 3968
rect 43220 3928 43229 3968
rect 32995 3844 33004 3884
rect 33044 3844 38860 3884
rect 38900 3844 38909 3884
rect 3679 3760 3688 3800
rect 3728 3760 3770 3800
rect 3810 3760 3852 3800
rect 3892 3760 3934 3800
rect 3974 3760 4016 3800
rect 4056 3760 4065 3800
rect 18799 3760 18808 3800
rect 18848 3760 18890 3800
rect 18930 3760 18972 3800
rect 19012 3760 19054 3800
rect 19094 3760 19136 3800
rect 19176 3760 19185 3800
rect 33919 3760 33928 3800
rect 33968 3760 34010 3800
rect 34050 3760 34092 3800
rect 34132 3760 34174 3800
rect 34214 3760 34256 3800
rect 34296 3760 34305 3800
rect 21475 3676 21484 3716
rect 21524 3676 21772 3716
rect 21812 3676 21821 3716
rect 643 3592 652 3632
rect 692 3592 36268 3632
rect 36308 3592 36317 3632
rect 19363 3508 19372 3548
rect 19412 3508 24364 3548
rect 24404 3508 24413 3548
rect 25027 3508 25036 3548
rect 25076 3508 27436 3548
rect 27476 3508 27485 3548
rect 451 3424 460 3464
rect 500 3424 38188 3464
rect 38228 3424 38237 3464
rect 1795 3340 1804 3380
rect 1844 3340 27628 3380
rect 27668 3340 27677 3380
rect 15043 3256 15052 3296
rect 15092 3256 16876 3296
rect 16916 3256 21580 3296
rect 21620 3256 21629 3296
rect 26947 3256 26956 3296
rect 26996 3256 43372 3296
rect 43412 3256 43421 3296
rect 18211 3172 18220 3212
rect 18260 3172 18796 3212
rect 18836 3172 21964 3212
rect 22004 3172 22013 3212
rect 24163 3088 24172 3128
rect 24212 3088 25612 3128
rect 25652 3088 25661 3128
rect 4919 3004 4928 3044
rect 4968 3004 5010 3044
rect 5050 3004 5092 3044
rect 5132 3004 5174 3044
rect 5214 3004 5256 3044
rect 5296 3004 5305 3044
rect 20039 3004 20048 3044
rect 20088 3004 20130 3044
rect 20170 3004 20212 3044
rect 20252 3004 20294 3044
rect 20334 3004 20376 3044
rect 20416 3004 20425 3044
rect 35159 3004 35168 3044
rect 35208 3004 35250 3044
rect 35290 3004 35332 3044
rect 35372 3004 35414 3044
rect 35454 3004 35496 3044
rect 35536 3004 35545 3044
rect 26851 2920 26860 2960
rect 26900 2920 27340 2960
rect 27380 2920 27389 2960
rect 19651 2752 19660 2792
rect 19700 2752 20716 2792
rect 20756 2752 20765 2792
rect 1411 2584 1420 2624
rect 1460 2584 40492 2624
rect 40532 2584 40541 2624
rect 3679 2248 3688 2288
rect 3728 2248 3770 2288
rect 3810 2248 3852 2288
rect 3892 2248 3934 2288
rect 3974 2248 4016 2288
rect 4056 2248 4065 2288
rect 18799 2248 18808 2288
rect 18848 2248 18890 2288
rect 18930 2248 18972 2288
rect 19012 2248 19054 2288
rect 19094 2248 19136 2288
rect 19176 2248 19185 2288
rect 33919 2248 33928 2288
rect 33968 2248 34010 2288
rect 34050 2248 34092 2288
rect 34132 2248 34174 2288
rect 34214 2248 34256 2288
rect 34296 2248 34305 2288
rect 30211 2164 30220 2204
rect 30260 2164 40012 2204
rect 40052 2164 40061 2204
rect 22915 1744 22924 1784
rect 22964 1744 30220 1784
rect 30260 1744 30269 1784
rect 4919 1492 4928 1532
rect 4968 1492 5010 1532
rect 5050 1492 5092 1532
rect 5132 1492 5174 1532
rect 5214 1492 5256 1532
rect 5296 1492 5305 1532
rect 20039 1492 20048 1532
rect 20088 1492 20130 1532
rect 20170 1492 20212 1532
rect 20252 1492 20294 1532
rect 20334 1492 20376 1532
rect 20416 1492 20425 1532
rect 35159 1492 35168 1532
rect 35208 1492 35250 1532
rect 35290 1492 35332 1532
rect 35372 1492 35414 1532
rect 35454 1492 35496 1532
rect 35536 1492 35545 1532
rect 36067 1156 36076 1196
rect 36116 1156 39244 1196
rect 39284 1156 39293 1196
rect 43651 64 43660 104
rect 43700 64 43852 104
rect 43892 64 43901 104
<< via4 >>
rect 19852 10480 19892 10520
rect 19468 10312 19508 10352
rect 19756 10228 19796 10268
rect 19660 9892 19700 9932
rect 3688 9808 3728 9848
rect 3770 9808 3810 9848
rect 3852 9808 3892 9848
rect 3934 9808 3974 9848
rect 4016 9808 4056 9848
rect 18808 9808 18848 9848
rect 18890 9808 18930 9848
rect 18972 9808 19012 9848
rect 19054 9808 19094 9848
rect 19136 9808 19176 9848
rect 33928 9808 33968 9848
rect 34010 9808 34050 9848
rect 34092 9808 34132 9848
rect 34174 9808 34214 9848
rect 34256 9808 34296 9848
rect 19468 9724 19508 9764
rect 19660 9724 19700 9764
rect 19756 9556 19796 9596
rect 4928 9052 4968 9092
rect 5010 9052 5050 9092
rect 5092 9052 5132 9092
rect 5174 9052 5214 9092
rect 5256 9052 5296 9092
rect 19756 9052 19796 9092
rect 20048 9052 20088 9092
rect 20130 9052 20170 9092
rect 20212 9052 20252 9092
rect 20294 9052 20334 9092
rect 20376 9052 20416 9092
rect 35168 9052 35208 9092
rect 35250 9052 35290 9092
rect 35332 9052 35372 9092
rect 35414 9052 35454 9092
rect 35496 9052 35536 9092
rect 19852 8632 19892 8672
rect 3688 8296 3728 8336
rect 3770 8296 3810 8336
rect 3852 8296 3892 8336
rect 3934 8296 3974 8336
rect 4016 8296 4056 8336
rect 18808 8296 18848 8336
rect 18890 8296 18930 8336
rect 18972 8296 19012 8336
rect 19054 8296 19094 8336
rect 19136 8296 19176 8336
rect 33928 8296 33968 8336
rect 34010 8296 34050 8336
rect 34092 8296 34132 8336
rect 34174 8296 34214 8336
rect 34256 8296 34296 8336
rect 4928 7540 4968 7580
rect 5010 7540 5050 7580
rect 5092 7540 5132 7580
rect 5174 7540 5214 7580
rect 5256 7540 5296 7580
rect 20048 7540 20088 7580
rect 20130 7540 20170 7580
rect 20212 7540 20252 7580
rect 20294 7540 20334 7580
rect 20376 7540 20416 7580
rect 35168 7540 35208 7580
rect 35250 7540 35290 7580
rect 35332 7540 35372 7580
rect 35414 7540 35454 7580
rect 35496 7540 35536 7580
rect 3688 6784 3728 6824
rect 3770 6784 3810 6824
rect 3852 6784 3892 6824
rect 3934 6784 3974 6824
rect 4016 6784 4056 6824
rect 18808 6784 18848 6824
rect 18890 6784 18930 6824
rect 18972 6784 19012 6824
rect 19054 6784 19094 6824
rect 19136 6784 19176 6824
rect 33928 6784 33968 6824
rect 34010 6784 34050 6824
rect 34092 6784 34132 6824
rect 34174 6784 34214 6824
rect 34256 6784 34296 6824
rect 4928 6028 4968 6068
rect 5010 6028 5050 6068
rect 5092 6028 5132 6068
rect 5174 6028 5214 6068
rect 5256 6028 5296 6068
rect 20048 6028 20088 6068
rect 20130 6028 20170 6068
rect 20212 6028 20252 6068
rect 20294 6028 20334 6068
rect 20376 6028 20416 6068
rect 35168 6028 35208 6068
rect 35250 6028 35290 6068
rect 35332 6028 35372 6068
rect 35414 6028 35454 6068
rect 35496 6028 35536 6068
rect 3688 5272 3728 5312
rect 3770 5272 3810 5312
rect 3852 5272 3892 5312
rect 3934 5272 3974 5312
rect 4016 5272 4056 5312
rect 18808 5272 18848 5312
rect 18890 5272 18930 5312
rect 18972 5272 19012 5312
rect 19054 5272 19094 5312
rect 19136 5272 19176 5312
rect 33928 5272 33968 5312
rect 34010 5272 34050 5312
rect 34092 5272 34132 5312
rect 34174 5272 34214 5312
rect 34256 5272 34296 5312
rect 4928 4516 4968 4556
rect 5010 4516 5050 4556
rect 5092 4516 5132 4556
rect 5174 4516 5214 4556
rect 5256 4516 5296 4556
rect 20048 4516 20088 4556
rect 20130 4516 20170 4556
rect 20212 4516 20252 4556
rect 20294 4516 20334 4556
rect 20376 4516 20416 4556
rect 35168 4516 35208 4556
rect 35250 4516 35290 4556
rect 35332 4516 35372 4556
rect 35414 4516 35454 4556
rect 35496 4516 35536 4556
rect 19756 4348 19796 4388
rect 3688 3760 3728 3800
rect 3770 3760 3810 3800
rect 3852 3760 3892 3800
rect 3934 3760 3974 3800
rect 4016 3760 4056 3800
rect 18808 3760 18848 3800
rect 18890 3760 18930 3800
rect 18972 3760 19012 3800
rect 19054 3760 19094 3800
rect 19136 3760 19176 3800
rect 33928 3760 33968 3800
rect 34010 3760 34050 3800
rect 34092 3760 34132 3800
rect 34174 3760 34214 3800
rect 34256 3760 34296 3800
rect 4928 3004 4968 3044
rect 5010 3004 5050 3044
rect 5092 3004 5132 3044
rect 5174 3004 5214 3044
rect 5256 3004 5296 3044
rect 20048 3004 20088 3044
rect 20130 3004 20170 3044
rect 20212 3004 20252 3044
rect 20294 3004 20334 3044
rect 20376 3004 20416 3044
rect 35168 3004 35208 3044
rect 35250 3004 35290 3044
rect 35332 3004 35372 3044
rect 35414 3004 35454 3044
rect 35496 3004 35536 3044
rect 3688 2248 3728 2288
rect 3770 2248 3810 2288
rect 3852 2248 3892 2288
rect 3934 2248 3974 2288
rect 4016 2248 4056 2288
rect 18808 2248 18848 2288
rect 18890 2248 18930 2288
rect 18972 2248 19012 2288
rect 19054 2248 19094 2288
rect 19136 2248 19176 2288
rect 33928 2248 33968 2288
rect 34010 2248 34050 2288
rect 34092 2248 34132 2288
rect 34174 2248 34214 2288
rect 34256 2248 34296 2288
rect 4928 1492 4968 1532
rect 5010 1492 5050 1532
rect 5092 1492 5132 1532
rect 5174 1492 5214 1532
rect 5256 1492 5296 1532
rect 20048 1492 20088 1532
rect 20130 1492 20170 1532
rect 20212 1492 20252 1532
rect 20294 1492 20334 1532
rect 20376 1492 20416 1532
rect 35168 1492 35208 1532
rect 35250 1492 35290 1532
rect 35332 1492 35372 1532
rect 35414 1492 35454 1532
rect 35496 1492 35536 1532
<< metal5 >>
rect 3652 9848 4092 11844
rect 3652 9808 3688 9848
rect 3728 9808 3770 9848
rect 3810 9808 3852 9848
rect 3892 9808 3934 9848
rect 3974 9808 4016 9848
rect 4056 9808 4092 9848
rect 3652 8336 4092 9808
rect 3652 8296 3688 8336
rect 3728 8296 3770 8336
rect 3810 8296 3852 8336
rect 3892 8296 3934 8336
rect 3974 8296 4016 8336
rect 4056 8296 4092 8336
rect 3652 6824 4092 8296
rect 3652 6784 3688 6824
rect 3728 6784 3770 6824
rect 3810 6784 3852 6824
rect 3892 6784 3934 6824
rect 3974 6784 4016 6824
rect 4056 6784 4092 6824
rect 3652 5312 4092 6784
rect 3652 5272 3688 5312
rect 3728 5272 3770 5312
rect 3810 5272 3852 5312
rect 3892 5272 3934 5312
rect 3974 5272 4016 5312
rect 4056 5272 4092 5312
rect 3652 3800 4092 5272
rect 3652 3760 3688 3800
rect 3728 3760 3770 3800
rect 3810 3760 3852 3800
rect 3892 3760 3934 3800
rect 3974 3760 4016 3800
rect 4056 3760 4092 3800
rect 3652 2288 4092 3760
rect 3652 2248 3688 2288
rect 3728 2248 3770 2288
rect 3810 2248 3852 2288
rect 3892 2248 3934 2288
rect 3974 2248 4016 2288
rect 4056 2248 4092 2288
rect 3652 0 4092 2248
rect 4892 9092 5332 11844
rect 4892 9052 4928 9092
rect 4968 9052 5010 9092
rect 5050 9052 5092 9092
rect 5132 9052 5174 9092
rect 5214 9052 5256 9092
rect 5296 9052 5332 9092
rect 4892 7580 5332 9052
rect 4892 7540 4928 7580
rect 4968 7540 5010 7580
rect 5050 7540 5092 7580
rect 5132 7540 5174 7580
rect 5214 7540 5256 7580
rect 5296 7540 5332 7580
rect 4892 6068 5332 7540
rect 4892 6028 4928 6068
rect 4968 6028 5010 6068
rect 5050 6028 5092 6068
rect 5132 6028 5174 6068
rect 5214 6028 5256 6068
rect 5296 6028 5332 6068
rect 4892 4556 5332 6028
rect 4892 4516 4928 4556
rect 4968 4516 5010 4556
rect 5050 4516 5092 4556
rect 5132 4516 5174 4556
rect 5214 4516 5256 4556
rect 5296 4516 5332 4556
rect 4892 3044 5332 4516
rect 4892 3004 4928 3044
rect 4968 3004 5010 3044
rect 5050 3004 5092 3044
rect 5132 3004 5174 3044
rect 5214 3004 5256 3044
rect 5296 3004 5332 3044
rect 4892 1532 5332 3004
rect 4892 1492 4928 1532
rect 4968 1492 5010 1532
rect 5050 1492 5092 1532
rect 5132 1492 5174 1532
rect 5214 1492 5256 1532
rect 5296 1492 5332 1532
rect 4892 0 5332 1492
rect 18772 9848 19212 11844
rect 19852 10520 19892 10529
rect 18772 9808 18808 9848
rect 18848 9808 18890 9848
rect 18930 9808 18972 9848
rect 19012 9808 19054 9848
rect 19094 9808 19136 9848
rect 19176 9808 19212 9848
rect 18772 8336 19212 9808
rect 19468 10352 19508 10361
rect 19468 9764 19508 10312
rect 19756 10268 19796 10277
rect 19468 9715 19508 9724
rect 19660 9932 19700 9941
rect 19660 9764 19700 9892
rect 19660 9715 19700 9724
rect 19756 9596 19796 10228
rect 19756 9547 19796 9556
rect 18772 8296 18808 8336
rect 18848 8296 18890 8336
rect 18930 8296 18972 8336
rect 19012 8296 19054 8336
rect 19094 8296 19136 8336
rect 19176 8296 19212 8336
rect 18772 6824 19212 8296
rect 18772 6784 18808 6824
rect 18848 6784 18890 6824
rect 18930 6784 18972 6824
rect 19012 6784 19054 6824
rect 19094 6784 19136 6824
rect 19176 6784 19212 6824
rect 18772 5312 19212 6784
rect 18772 5272 18808 5312
rect 18848 5272 18890 5312
rect 18930 5272 18972 5312
rect 19012 5272 19054 5312
rect 19094 5272 19136 5312
rect 19176 5272 19212 5312
rect 18772 3800 19212 5272
rect 19756 9092 19796 9101
rect 19756 4388 19796 9052
rect 19852 8672 19892 10480
rect 19852 8623 19892 8632
rect 20012 9092 20452 11844
rect 20012 9052 20048 9092
rect 20088 9052 20130 9092
rect 20170 9052 20212 9092
rect 20252 9052 20294 9092
rect 20334 9052 20376 9092
rect 20416 9052 20452 9092
rect 19756 4339 19796 4348
rect 20012 7580 20452 9052
rect 20012 7540 20048 7580
rect 20088 7540 20130 7580
rect 20170 7540 20212 7580
rect 20252 7540 20294 7580
rect 20334 7540 20376 7580
rect 20416 7540 20452 7580
rect 20012 6068 20452 7540
rect 20012 6028 20048 6068
rect 20088 6028 20130 6068
rect 20170 6028 20212 6068
rect 20252 6028 20294 6068
rect 20334 6028 20376 6068
rect 20416 6028 20452 6068
rect 20012 4556 20452 6028
rect 20012 4516 20048 4556
rect 20088 4516 20130 4556
rect 20170 4516 20212 4556
rect 20252 4516 20294 4556
rect 20334 4516 20376 4556
rect 20416 4516 20452 4556
rect 18772 3760 18808 3800
rect 18848 3760 18890 3800
rect 18930 3760 18972 3800
rect 19012 3760 19054 3800
rect 19094 3760 19136 3800
rect 19176 3760 19212 3800
rect 18772 2288 19212 3760
rect 18772 2248 18808 2288
rect 18848 2248 18890 2288
rect 18930 2248 18972 2288
rect 19012 2248 19054 2288
rect 19094 2248 19136 2288
rect 19176 2248 19212 2288
rect 18772 0 19212 2248
rect 20012 3044 20452 4516
rect 20012 3004 20048 3044
rect 20088 3004 20130 3044
rect 20170 3004 20212 3044
rect 20252 3004 20294 3044
rect 20334 3004 20376 3044
rect 20416 3004 20452 3044
rect 20012 1532 20452 3004
rect 20012 1492 20048 1532
rect 20088 1492 20130 1532
rect 20170 1492 20212 1532
rect 20252 1492 20294 1532
rect 20334 1492 20376 1532
rect 20416 1492 20452 1532
rect 20012 0 20452 1492
rect 33892 9848 34332 11844
rect 33892 9808 33928 9848
rect 33968 9808 34010 9848
rect 34050 9808 34092 9848
rect 34132 9808 34174 9848
rect 34214 9808 34256 9848
rect 34296 9808 34332 9848
rect 33892 8336 34332 9808
rect 33892 8296 33928 8336
rect 33968 8296 34010 8336
rect 34050 8296 34092 8336
rect 34132 8296 34174 8336
rect 34214 8296 34256 8336
rect 34296 8296 34332 8336
rect 33892 6824 34332 8296
rect 33892 6784 33928 6824
rect 33968 6784 34010 6824
rect 34050 6784 34092 6824
rect 34132 6784 34174 6824
rect 34214 6784 34256 6824
rect 34296 6784 34332 6824
rect 33892 5312 34332 6784
rect 33892 5272 33928 5312
rect 33968 5272 34010 5312
rect 34050 5272 34092 5312
rect 34132 5272 34174 5312
rect 34214 5272 34256 5312
rect 34296 5272 34332 5312
rect 33892 3800 34332 5272
rect 33892 3760 33928 3800
rect 33968 3760 34010 3800
rect 34050 3760 34092 3800
rect 34132 3760 34174 3800
rect 34214 3760 34256 3800
rect 34296 3760 34332 3800
rect 33892 2288 34332 3760
rect 33892 2248 33928 2288
rect 33968 2248 34010 2288
rect 34050 2248 34092 2288
rect 34132 2248 34174 2288
rect 34214 2248 34256 2288
rect 34296 2248 34332 2288
rect 33892 0 34332 2248
rect 35132 9092 35572 11844
rect 35132 9052 35168 9092
rect 35208 9052 35250 9092
rect 35290 9052 35332 9092
rect 35372 9052 35414 9092
rect 35454 9052 35496 9092
rect 35536 9052 35572 9092
rect 35132 7580 35572 9052
rect 35132 7540 35168 7580
rect 35208 7540 35250 7580
rect 35290 7540 35332 7580
rect 35372 7540 35414 7580
rect 35454 7540 35496 7580
rect 35536 7540 35572 7580
rect 35132 6068 35572 7540
rect 35132 6028 35168 6068
rect 35208 6028 35250 6068
rect 35290 6028 35332 6068
rect 35372 6028 35414 6068
rect 35454 6028 35496 6068
rect 35536 6028 35572 6068
rect 35132 4556 35572 6028
rect 35132 4516 35168 4556
rect 35208 4516 35250 4556
rect 35290 4516 35332 4556
rect 35372 4516 35414 4556
rect 35454 4516 35496 4556
rect 35536 4516 35572 4556
rect 35132 3044 35572 4516
rect 35132 3004 35168 3044
rect 35208 3004 35250 3044
rect 35290 3004 35332 3044
rect 35372 3004 35414 3044
rect 35454 3004 35496 3044
rect 35536 3004 35572 3044
rect 35132 1532 35572 3004
rect 35132 1492 35168 1532
rect 35208 1492 35250 1532
rect 35290 1492 35332 1532
rect 35372 1492 35414 1532
rect 35454 1492 35496 1532
rect 35536 1492 35572 1532
rect 35132 0 35572 1492
use sg13g2_inv_1  _016_
timestamp 1676382929
transform -1 0 13440 0 -1 6048
box -48 -56 336 834
use sg13g2_inv_1  _017_
timestamp 1676382929
transform -1 0 12864 0 1 7560
box -48 -56 336 834
use sg13g2_mux4_1  _018_
timestamp 1677257233
transform 1 0 9312 0 1 6048
box -48 -56 2064 834
use sg13g2_inv_1  _019_
timestamp 1676382929
transform -1 0 13152 0 -1 7560
box -48 -56 336 834
use sg13g2_mux2_1  _020_
timestamp 1677247768
transform 1 0 9984 0 -1 7560
box -48 -56 1008 834
use sg13g2_nand2b_1  _021_
timestamp 1676567195
transform 1 0 11520 0 -1 9072
box -48 -56 528 834
use sg13g2_mux2_1  _022_
timestamp 1677247768
transform 1 0 11616 0 1 7560
box -48 -56 1008 834
use sg13g2_a21oi_1  _023_
timestamp 1683973020
transform -1 0 12864 0 -1 7560
box -48 -56 528 834
use sg13g2_a221oi_1  _024_
timestamp 1685197497
transform -1 0 12384 0 -1 7560
box -48 -56 816 834
use sg13g2_mux4_1  _025_
timestamp 1677257233
transform 1 0 9600 0 1 7560
box -48 -56 2064 834
use sg13g2_mux4_1  _026_
timestamp 1677257233
transform 1 0 9216 0 -1 6048
box -48 -56 2064 834
use sg13g2_mux2_1  _027_
timestamp 1677247768
transform 1 0 11328 0 1 6048
box -48 -56 1008 834
use sg13g2_mux4_1  _028_
timestamp 1677257233
transform 1 0 26208 0 1 7560
box -48 -56 2064 834
use sg13g2_mux4_1  _029_
timestamp 1677257233
transform 1 0 26112 0 -1 7560
box -48 -56 2064 834
use sg13g2_mux2_1  _030_
timestamp 1677247768
transform -1 0 28224 0 -1 9072
box -48 -56 1008 834
use sg13g2_mux4_1  _031_
timestamp 1677257233
transform 1 0 31584 0 -1 4536
box -48 -56 2064 834
use sg13g2_mux4_1  _032_
timestamp 1677257233
transform 1 0 30528 0 1 3024
box -48 -56 2064 834
use sg13g2_mux2_1  _033_
timestamp 1677247768
transform -1 0 34560 0 -1 4536
box -48 -56 1008 834
use sg13g2_mux4_1  _034_
timestamp 1677257233
transform 1 0 18912 0 1 3024
box -48 -56 2064 834
use sg13g2_mux4_1  _035_
timestamp 1677257233
transform 1 0 18048 0 -1 3024
box -48 -56 2064 834
use sg13g2_mux2_1  _036_
timestamp 1677247768
transform -1 0 21984 0 1 3024
box -48 -56 1008 834
use sg13g2_mux2_1  _037_
timestamp 1677247768
transform 1 0 15360 0 -1 3024
box -48 -56 1008 834
use sg13g2_mux2_1  _038_
timestamp 1677247768
transform 1 0 26016 0 1 3024
box -48 -56 1008 834
use sg13g2_mux2_1  _039_
timestamp 1677247768
transform 1 0 25728 0 -1 4536
box -48 -56 1008 834
use sg13g2_mux2_1  _040_
timestamp 1677247768
transform -1 0 10272 0 -1 4536
box -48 -56 1008 834
use sg13g2_dlhq_1  _041_
timestamp 1678805552
transform 1 0 7680 0 -1 3024
box -50 -56 1692 834
use sg13g2_dlhq_1  _042_
timestamp 1678805552
transform 1 0 24096 0 -1 4536
box -50 -56 1692 834
use sg13g2_dlhq_1  _043_
timestamp 1678805552
transform 1 0 24192 0 1 3024
box -50 -56 1692 834
use sg13g2_dlhq_1  _044_
timestamp 1678805552
transform 1 0 13728 0 1 3024
box -50 -56 1692 834
use sg13g2_dlhq_1  _045_
timestamp 1678805552
transform 1 0 14784 0 -1 7560
box -50 -56 1692 834
use sg13g2_dlhq_1  _046_
timestamp 1678805552
transform 1 0 14784 0 1 7560
box -50 -56 1692 834
use sg13g2_dlhq_1  _047_
timestamp 1678805552
transform 1 0 12096 0 1 3024
box -50 -56 1692 834
use sg13g2_dlhq_1  _048_
timestamp 1678805552
transform 1 0 16128 0 1 3024
box -50 -56 1692 834
use sg13g2_dlhq_1  _049_
timestamp 1678805552
transform 1 0 17952 0 -1 4536
box -50 -56 1692 834
use sg13g2_dlhq_1  _050_
timestamp 1678805552
transform -1 0 23040 0 -1 4536
box -50 -56 1692 834
use sg13g2_dlhq_1  _051_
timestamp 1678805552
transform 1 0 27936 0 1 3024
box -50 -56 1692 834
use sg13g2_dlhq_1  _052_
timestamp 1678805552
transform 1 0 29952 0 -1 4536
box -50 -56 1692 834
use sg13g2_dlhq_1  _053_
timestamp 1678805552
transform 1 0 31296 0 1 4536
box -50 -56 1692 834
use sg13g2_dlhq_1  _054_
timestamp 1678805552
transform 1 0 23232 0 -1 7560
box -50 -56 1692 834
use sg13g2_dlhq_1  _055_
timestamp 1678805552
transform -1 0 30720 0 -1 7560
box -50 -56 1692 834
use sg13g2_dlhq_1  _056_
timestamp 1678805552
transform 1 0 23328 0 1 7560
box -50 -56 1692 834
use sg13g2_dlhq_1  _057_
timestamp 1678805552
transform 1 0 6432 0 1 6048
box -50 -56 1692 834
use sg13g2_dlhq_1  _058_
timestamp 1678805552
transform 1 0 9696 0 1 3024
box -50 -56 1692 834
use sg13g2_dlhq_1  _059_
timestamp 1678805552
transform 1 0 9408 0 -1 3024
box -50 -56 1692 834
use sg13g2_buf_1  _061_
timestamp 1676381911
transform 1 0 40032 0 -1 3024
box -48 -56 432 834
use sg13g2_buf_1  _062_
timestamp 1676381911
transform 1 0 39648 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  _063_
timestamp 1676381911
transform 1 0 39264 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  _064_
timestamp 1676381911
transform 1 0 38112 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  _065_
timestamp 1676381911
transform 1 0 39648 0 -1 3024
box -48 -56 432 834
use sg13g2_buf_1  _066_
timestamp 1676381911
transform 1 0 38496 0 -1 4536
box -48 -56 432 834
use sg13g2_buf_1  _067_
timestamp 1676381911
transform 1 0 37728 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  _068_
timestamp 1676381911
transform 1 0 40416 0 -1 3024
box -48 -56 432 834
use sg13g2_buf_1  _069_
timestamp 1676381911
transform 1 0 36288 0 -1 3024
box -48 -56 432 834
use sg13g2_buf_1  _070_
timestamp 1676381911
transform 1 0 36384 0 1 7560
box -48 -56 432 834
use sg13g2_buf_1  _071_
timestamp 1676381911
transform 1 0 32640 0 1 7560
box -48 -56 432 834
use sg13g2_buf_1  _072_
timestamp 1676381911
transform 1 0 33408 0 1 7560
box -48 -56 432 834
use sg13g2_buf_1  _073_
timestamp 1676381911
transform 1 0 33792 0 1 7560
box -48 -56 432 834
use sg13g2_buf_1  _074_
timestamp 1676381911
transform 1 0 7296 0 -1 3024
box -48 -56 432 834
use sg13g2_buf_1  _075_
timestamp 1676381911
transform 1 0 23712 0 -1 4536
box -48 -56 432 834
use sg13g2_buf_1  _076_
timestamp 1676381911
transform 1 0 24192 0 -1 3024
box -48 -56 432 834
use sg13g2_buf_1  _077_
timestamp 1676381911
transform 1 0 13728 0 -1 3024
box -48 -56 432 834
use sg13g2_buf_1  _078_
timestamp 1676381911
transform 1 0 14880 0 -1 9072
box -48 -56 432 834
use sg13g2_buf_1  _079_
timestamp 1676381911
transform 1 0 14400 0 1 7560
box -48 -56 432 834
use sg13g2_buf_1  _080_
timestamp 1676381911
transform 1 0 11712 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  _081_
timestamp 1676381911
transform 1 0 15360 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  _082_
timestamp 1676381911
transform 1 0 17568 0 -1 4536
box -48 -56 432 834
use sg13g2_buf_1  _083_
timestamp 1676381911
transform 1 0 21024 0 -1 4536
box -48 -56 432 834
use sg13g2_buf_1  _084_
timestamp 1676381911
transform 1 0 27552 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  _085_
timestamp 1676381911
transform 1 0 30144 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  _086_
timestamp 1676381911
transform 1 0 30912 0 1 4536
box -48 -56 432 834
use sg13g2_buf_1  _087_
timestamp 1676381911
transform 1 0 22560 0 1 7560
box -48 -56 432 834
use sg13g2_buf_1  _088_
timestamp 1676381911
transform 1 0 29376 0 1 7560
box -48 -56 432 834
use sg13g2_buf_1  _089_
timestamp 1676381911
transform 1 0 22944 0 1 7560
box -48 -56 432 834
use sg13g2_buf_1  _090_
timestamp 1676381911
transform 1 0 6048 0 1 6048
box -48 -56 432 834
use sg13g2_buf_1  _091_
timestamp 1676381911
transform 1 0 8928 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  _092_
timestamp 1676381911
transform 1 0 9312 0 1 1512
box -48 -56 432 834
use sg13g2_buf_1  _093_
timestamp 1676381911
transform 1 0 26688 0 -1 4536
box -48 -56 432 834
use sg13g2_buf_1  _094_
timestamp 1676381911
transform -1 0 43200 0 -1 3024
box -48 -56 432 834
use sg13g2_buf_1  _095_
timestamp 1676381911
transform -1 0 43200 0 1 4536
box -48 -56 432 834
use sg13g2_buf_1  _096_
timestamp 1676381911
transform -1 0 43488 0 -1 4536
box -48 -56 432 834
use sg13g2_buf_1  _097_
timestamp 1676381911
transform -1 0 43104 0 -1 4536
box -48 -56 432 834
use sg13g2_buf_1  _098_
timestamp 1676381911
transform -1 0 43872 0 -1 4536
box -48 -56 432 834
use sg13g2_buf_1  _099_
timestamp 1676381911
transform -1 0 42720 0 -1 4536
box -48 -56 432 834
use sg13g2_buf_1  _100_
timestamp 1676381911
transform -1 0 42336 0 -1 4536
box -48 -56 432 834
use sg13g2_buf_1  _101_
timestamp 1676381911
transform -1 0 43488 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  _102_
timestamp 1676381911
transform -1 0 43872 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  _103_
timestamp 1676381911
transform -1 0 44256 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  _104_
timestamp 1676381911
transform -1 0 42624 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  _105_
timestamp 1676381911
transform -1 0 43872 0 -1 9072
box -48 -56 432 834
use sg13g2_buf_1  _106_
timestamp 1676381911
transform -1 0 44256 0 1 7560
box -48 -56 432 834
use sg13g2_buf_1  _107_
timestamp 1676381911
transform 1 0 32256 0 -1 7560
box -48 -56 432 834
use sg13g2_buf_1  _108_
timestamp 1676381911
transform 1 0 34176 0 1 7560
box -48 -56 432 834
use sg13g2_buf_1  _109_
timestamp 1676381911
transform -1 0 35328 0 1 7560
box -48 -56 432 834
use sg13g2_buf_1  _110_
timestamp 1676381911
transform 1 0 34560 0 1 7560
box -48 -56 432 834
use sg13g2_buf_1  _111_
timestamp 1676381911
transform 1 0 31776 0 1 7560
box -48 -56 432 834
use sg13g2_buf_1  _112_
timestamp 1676381911
transform -1 0 43104 0 1 7560
box -48 -56 432 834
use sg13g2_buf_1  _113_
timestamp 1676381911
transform 1 0 9312 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  _114_
timestamp 1676381911
transform -1 0 27456 0 -1 4536
box -48 -56 432 834
use sg13g2_buf_1  _115_
timestamp 1676381911
transform -1 0 27360 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  _116_
timestamp 1676381911
transform -1 0 16128 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  _117_
timestamp 1676381911
transform 1 0 3552 0 1 7560
box -48 -56 432 834
use sg13g2_buf_1  _118_
timestamp 1676381911
transform 1 0 3936 0 1 7560
box -48 -56 432 834
use sg13g2_buf_1  _119_
timestamp 1676381911
transform 1 0 4320 0 1 7560
box -48 -56 432 834
use sg13g2_buf_1  _120_
timestamp 1676381911
transform 1 0 3168 0 1 7560
box -48 -56 432 834
use sg13g2_buf_1  _121_
timestamp 1676381911
transform 1 0 9600 0 -1 7560
box -48 -56 432 834
use sg13g2_buf_1  _122_
timestamp 1676381911
transform -1 0 27168 0 -1 9072
box -48 -56 432 834
use sg13g2_buf_1  _123_
timestamp 1676381911
transform -1 0 31392 0 -1 3024
box -48 -56 432 834
use sg13g2_buf_1  _124_
timestamp 1676381911
transform -1 0 18912 0 1 1512
box -48 -56 432 834
use sg13g2_buf_1  _125_
timestamp 1676381911
transform 1 0 11232 0 -1 6048
box -48 -56 432 834
use sg13g2_buf_1  _126_
timestamp 1676381911
transform -1 0 28512 0 -1 7560
box -48 -56 432 834
use sg13g2_buf_1  _127_
timestamp 1676381911
transform -1 0 32160 0 -1 3024
box -48 -56 432 834
use sg13g2_buf_1  _128_
timestamp 1676381911
transform -1 0 18912 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  _129_
timestamp 1676381911
transform 1 0 8928 0 1 6048
box -48 -56 432 834
use sg13g2_buf_1  _130_
timestamp 1676381911
transform -1 0 28608 0 1 7560
box -48 -56 432 834
use sg13g2_buf_1  _131_
timestamp 1676381911
transform -1 0 31776 0 -1 3024
box -48 -56 432 834
use sg13g2_buf_1  _132_
timestamp 1676381911
transform -1 0 18144 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  _133_
timestamp 1676381911
transform -1 0 42720 0 1 7560
box -48 -56 432 834
use sg13g2_buf_1  _134_
timestamp 1676381911
transform -1 0 43488 0 1 7560
box -48 -56 432 834
use sg13g2_buf_1  _135_
timestamp 1676381911
transform -1 0 42336 0 1 7560
box -48 -56 432 834
use sg13g2_buf_1  _136_
timestamp 1676381911
transform -1 0 43104 0 -1 9072
box -48 -56 432 834
use sg13g2_buf_1  _137_
timestamp 1676381911
transform -1 0 43872 0 1 7560
box -48 -56 432 834
use sg13g2_buf_1  _138_
timestamp 1676381911
transform 1 0 2784 0 1 7560
box -48 -56 432 834
use sg13g2_buf_1  _139_
timestamp 1676381911
transform 1 0 2400 0 1 7560
box -48 -56 432 834
use sg13g2_buf_1  _140_
timestamp 1676381911
transform -1 0 18240 0 1 7560
box -48 -56 432 834
use sg13g2_buf_1  _141_
timestamp 1676381911
transform 1 0 9984 0 -1 9072
box -48 -56 432 834
use sg13g2_buf_1  _142_
timestamp 1676381911
transform -1 0 28992 0 1 7560
box -48 -56 432 834
use sg13g2_buf_1  _143_
timestamp 1676381911
transform -1 0 33312 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  _144_
timestamp 1676381911
transform -1 0 20448 0 -1 4536
box -48 -56 432 834
use sg13g2_buf_1  _145_
timestamp 1676381911
transform 1 0 9600 0 -1 9072
box -48 -56 432 834
use sg13g2_buf_1  _146_
timestamp 1676381911
transform -1 0 26208 0 1 7560
box -48 -56 432 834
use sg13g2_buf_1  _147_
timestamp 1676381911
transform -1 0 32928 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  _148_
timestamp 1676381911
transform -1 0 18528 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  _149_
timestamp 1676381911
transform -1 0 42048 0 -1 7560
box -48 -56 432 834
use sg13g2_buf_1  _150_
timestamp 1676381911
transform -1 0 42432 0 -1 7560
box -48 -56 432 834
use sg13g2_buf_1  _151_
timestamp 1676381911
transform -1 0 43584 0 -1 7560
box -48 -56 432 834
use sg13g2_buf_1  _152_
timestamp 1676381911
transform -1 0 43200 0 -1 7560
box -48 -56 432 834
use sg13g2_buf_1  _153_
timestamp 1676381911
transform -1 0 42816 0 -1 7560
box -48 -56 432 834
use sg13g2_buf_1  _154_
timestamp 1676381911
transform -1 0 41952 0 1 7560
box -48 -56 432 834
use sg13g2_buf_1  _155_
timestamp 1676381911
transform -1 0 43488 0 -1 9072
box -48 -56 432 834
use sg13g2_buf_1  _156_
timestamp 1676381911
transform -1 0 42720 0 -1 9072
box -48 -56 432 834
use sg13g2_buf_1  _157_
timestamp 1676381911
transform 1 0 11040 0 -1 7560
box -48 -56 432 834
use sg13g2_buf_1  _158_
timestamp 1676381911
transform -1 0 28608 0 -1 9072
box -48 -56 432 834
use sg13g2_buf_1  _159_
timestamp 1676381911
transform -1 0 33696 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  _160_
timestamp 1676381911
transform -1 0 20544 0 -1 3024
box -48 -56 432 834
use sg13g2_buf_1  _161_
timestamp 1676381911
transform 1 0 10752 0 -1 9072
box -48 -56 432 834
use sg13g2_buf_1  _162_
timestamp 1676381911
transform -1 0 26784 0 -1 9072
box -48 -56 432 834
use sg13g2_buf_1  _163_
timestamp 1676381911
transform -1 0 33312 0 1 4536
box -48 -56 432 834
use sg13g2_buf_1  _164_
timestamp 1676381911
transform 1 0 19680 0 -1 4536
box -48 -56 432 834
use sg13g2_buf_1  _165_
timestamp 1676381911
transform -1 0 43104 0 1 3024
box -48 -56 432 834
use sg13g2_antennanp  ANTENNA_1
timestamp 1679999689
transform 1 0 36096 0 -1 7560
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_2
timestamp 1679999689
transform 1 0 37824 0 -1 7560
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_3
timestamp 1679999689
transform 1 0 37536 0 -1 7560
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_4
timestamp 1679999689
transform 1 0 38976 0 1 3024
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_5
timestamp 1679999689
transform 1 0 38496 0 1 3024
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_6
timestamp 1679999689
transform -1 0 38496 0 -1 4536
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_7
timestamp 1679999689
transform 1 0 37152 0 1 3024
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_8
timestamp 1679999689
transform 1 0 36768 0 1 7560
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_9
timestamp 1679999689
transform 1 0 44160 0 1 6048
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_10
timestamp 1679999689
transform 1 0 41856 0 1 9072
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_11
timestamp 1679999689
transform 1 0 31488 0 1 7560
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_12
timestamp 1679999689
transform 1 0 37248 0 -1 7560
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_13
timestamp 1679999689
transform 1 0 36672 0 -1 7560
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_14
timestamp 1679999689
transform 1 0 40224 0 1 1512
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_15
timestamp 1679999689
transform 1 0 36864 0 1 3024
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_16
timestamp 1679999689
transform 1 0 36096 0 1 7560
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_17
timestamp 1679999689
transform 1 0 43872 0 -1 4536
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_18
timestamp 1679999689
transform 1 0 43872 0 1 6048
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_19
timestamp 1679999689
transform 1 0 43392 0 1 9072
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_20
timestamp 1679999689
transform 1 0 39648 0 1 1512
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_21
timestamp 1679999689
transform 1 0 35520 0 -1 7560
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_22
timestamp 1679999689
transform 1 0 36960 0 -1 7560
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_23
timestamp 1679999689
transform 1 0 38592 0 -1 3024
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_24
timestamp 1679999689
transform 1 0 43296 0 1 4536
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_25
timestamp 1679999689
transform -1 0 44160 0 -1 7560
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_26
timestamp 1679999689
transform 1 0 40512 0 1 1512
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_27
timestamp 1679999689
transform 1 0 34944 0 -1 7560
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_28
timestamp 1679999689
transform 1 0 36384 0 -1 7560
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_29
timestamp 1679999689
transform 1 0 38304 0 -1 3024
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_30
timestamp 1679999689
transform 1 0 43872 0 1 4536
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_31
timestamp 1679999689
transform -1 0 43872 0 -1 7560
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_32
timestamp 1679999689
transform 1 0 34368 0 -1 7560
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_33
timestamp 1679999689
transform 1 0 35808 0 -1 7560
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_34
timestamp 1679999689
transform 1 0 38016 0 -1 3024
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_35
timestamp 1679999689
transform 1 0 43584 0 1 4536
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_36
timestamp 1679999689
transform 1 0 43584 0 1 6048
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_37
timestamp 1679999689
transform 1 0 33792 0 -1 7560
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_38
timestamp 1679999689
transform 1 0 35232 0 -1 7560
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_39
timestamp 1679999689
transform 1 0 37728 0 -1 3024
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_40
timestamp 1679999689
transform -1 0 44160 0 -1 6048
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_41
timestamp 1679999689
transform 1 0 43584 0 -1 6048
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_42
timestamp 1679999689
transform 1 0 33216 0 -1 7560
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_43
timestamp 1679999689
transform 1 0 34656 0 -1 7560
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_44
timestamp 1679999689
transform 1 0 37440 0 -1 3024
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_45
timestamp 1679999689
transform 1 0 44544 0 -1 4536
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_46
timestamp 1679999689
transform 1 0 44160 0 1 4536
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_47
timestamp 1679999689
transform 1 0 32928 0 -1 7560
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_48
timestamp 1679999689
transform 1 0 34080 0 -1 7560
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_49
timestamp 1679999689
transform -1 0 40224 0 1 1512
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_50
timestamp 1679999689
transform 1 0 37440 0 1 3024
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_51
timestamp 1679999689
transform 1 0 44160 0 -1 6048
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_52
timestamp 1679999689
transform 1 0 39360 0 1 1512
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_53
timestamp 1679999689
transform 1 0 32640 0 -1 7560
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_54
timestamp 1679999689
transform 1 0 33504 0 -1 7560
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_55
timestamp 1679999689
transform -1 0 39360 0 1 1512
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_56
timestamp 1679999689
transform 1 0 41088 0 -1 3024
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_57
timestamp 1679999689
transform 1 0 44832 0 1 6048
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_58
timestamp 1679999689
transform -1 0 39648 0 -1 3024
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_59
timestamp 1679999689
transform 1 0 32352 0 1 7560
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_60
timestamp 1679999689
transform 1 0 33120 0 1 7560
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_61
timestamp 1679999689
transform -1 0 39360 0 -1 3024
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_62
timestamp 1679999689
transform 1 0 40800 0 -1 3024
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_63
timestamp 1679999689
transform -1 0 44832 0 -1 7560
box -48 -56 336 834
use sg13g2_buf_1  fanout7
timestamp 1676381911
transform -1 0 17280 0 1 6048
box -48 -56 432 834
use sg13g2_buf_1  fanout8
timestamp 1676381911
transform 1 0 21600 0 -1 7560
box -48 -56 432 834
use sg13g2_buf_1  fanout9
timestamp 1676381911
transform 1 0 16896 0 1 7560
box -48 -56 432 834
use sg13g2_decap_8  FILLER_0_0
timestamp 1679581782
transform 1 0 1152 0 1 1512
box -48 -56 720 834
use sg13g2_decap_4  FILLER_0_7
timestamp 1679577901
transform 1 0 1824 0 1 1512
box -48 -56 432 834
use sg13g2_fill_2  FILLER_0_11
timestamp 1677580104
transform 1 0 2208 0 1 1512
box -48 -56 240 834
use sg13g2_decap_8  FILLER_0_17
timestamp 1679581782
transform 1 0 2784 0 1 1512
box -48 -56 720 834
use sg13g2_decap_4  FILLER_0_24
timestamp 1679577901
transform 1 0 3456 0 1 1512
box -48 -56 432 834
use sg13g2_fill_1  FILLER_0_28
timestamp 1677579658
transform 1 0 3840 0 1 1512
box -48 -56 144 834
use sg13g2_decap_8  FILLER_0_33
timestamp 1679581782
transform 1 0 4320 0 1 1512
box -48 -56 720 834
use sg13g2_decap_4  FILLER_0_40
timestamp 1679577901
transform 1 0 4992 0 1 1512
box -48 -56 432 834
use sg13g2_fill_1  FILLER_0_44
timestamp 1677579658
transform 1 0 5376 0 1 1512
box -48 -56 144 834
use sg13g2_decap_8  FILLER_0_49
timestamp 1679581782
transform 1 0 5856 0 1 1512
box -48 -56 720 834
use sg13g2_decap_4  FILLER_0_56
timestamp 1679577901
transform 1 0 6528 0 1 1512
box -48 -56 432 834
use sg13g2_fill_1  FILLER_0_60
timestamp 1677579658
transform 1 0 6912 0 1 1512
box -48 -56 144 834
use sg13g2_decap_8  FILLER_0_65
timestamp 1679581782
transform 1 0 7392 0 1 1512
box -48 -56 720 834
use sg13g2_decap_4  FILLER_0_72
timestamp 1679577901
transform 1 0 8064 0 1 1512
box -48 -56 432 834
use sg13g2_fill_1  FILLER_0_76
timestamp 1677579658
transform 1 0 8448 0 1 1512
box -48 -56 144 834
use sg13g2_decap_4  FILLER_0_81
timestamp 1679577901
transform 1 0 8928 0 1 1512
box -48 -56 432 834
use sg13g2_decap_4  FILLER_0_89
timestamp 1679577901
transform 1 0 9696 0 1 1512
box -48 -56 432 834
use sg13g2_decap_8  FILLER_0_97
timestamp 1679581782
transform 1 0 10464 0 1 1512
box -48 -56 720 834
use sg13g2_decap_4  FILLER_0_104
timestamp 1679577901
transform 1 0 11136 0 1 1512
box -48 -56 432 834
use sg13g2_fill_1  FILLER_0_108
timestamp 1677579658
transform 1 0 11520 0 1 1512
box -48 -56 144 834
use sg13g2_decap_8  FILLER_0_113
timestamp 1679581782
transform 1 0 12000 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_120
timestamp 1679581782
transform 1 0 12672 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_127
timestamp 1679581782
transform 1 0 13344 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_134
timestamp 1679581782
transform 1 0 14016 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_141
timestamp 1679581782
transform 1 0 14688 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_148
timestamp 1679581782
transform 1 0 15360 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_155
timestamp 1679581782
transform 1 0 16032 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_162
timestamp 1679581782
transform 1 0 16704 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_169
timestamp 1679581782
transform 1 0 17376 0 1 1512
box -48 -56 720 834
use sg13g2_decap_4  FILLER_0_176
timestamp 1679577901
transform 1 0 18048 0 1 1512
box -48 -56 432 834
use sg13g2_fill_1  FILLER_0_180
timestamp 1677579658
transform 1 0 18432 0 1 1512
box -48 -56 144 834
use sg13g2_decap_8  FILLER_0_185
timestamp 1679581782
transform 1 0 18912 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_192
timestamp 1679581782
transform 1 0 19584 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_199
timestamp 1679581782
transform 1 0 20256 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_206
timestamp 1679581782
transform 1 0 20928 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_213
timestamp 1679581782
transform 1 0 21600 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_220
timestamp 1679581782
transform 1 0 22272 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_227
timestamp 1679581782
transform 1 0 22944 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_234
timestamp 1679581782
transform 1 0 23616 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_241
timestamp 1679581782
transform 1 0 24288 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_248
timestamp 1679581782
transform 1 0 24960 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_255
timestamp 1679581782
transform 1 0 25632 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_262
timestamp 1679581782
transform 1 0 26304 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_269
timestamp 1679581782
transform 1 0 26976 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_276
timestamp 1679581782
transform 1 0 27648 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_283
timestamp 1679581782
transform 1 0 28320 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_290
timestamp 1679581782
transform 1 0 28992 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_297
timestamp 1679581782
transform 1 0 29664 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_304
timestamp 1679581782
transform 1 0 30336 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_311
timestamp 1679581782
transform 1 0 31008 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_318
timestamp 1679581782
transform 1 0 31680 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_325
timestamp 1679581782
transform 1 0 32352 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_332
timestamp 1679581782
transform 1 0 33024 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_339
timestamp 1679581782
transform 1 0 33696 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_346
timestamp 1679581782
transform 1 0 34368 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_353
timestamp 1679581782
transform 1 0 35040 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_360
timestamp 1679581782
transform 1 0 35712 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_367
timestamp 1679581782
transform 1 0 36384 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_374
timestamp 1679581782
transform 1 0 37056 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_381
timestamp 1679581782
transform 1 0 37728 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_388
timestamp 1679581782
transform 1 0 38400 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_413
timestamp 1679581782
transform 1 0 40800 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_420
timestamp 1679581782
transform 1 0 41472 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_427
timestamp 1679581782
transform 1 0 42144 0 1 1512
box -48 -56 720 834
use sg13g2_fill_1  FILLER_0_434
timestamp 1677579658
transform 1 0 42816 0 1 1512
box -48 -56 144 834
use sg13g2_decap_8  FILLER_1_0
timestamp 1679581782
transform 1 0 1152 0 -1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_7
timestamp 1679581782
transform 1 0 1824 0 -1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_14
timestamp 1679581782
transform 1 0 2496 0 -1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_21
timestamp 1679581782
transform 1 0 3168 0 -1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_28
timestamp 1679581782
transform 1 0 3840 0 -1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_35
timestamp 1679581782
transform 1 0 4512 0 -1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_42
timestamp 1679581782
transform 1 0 5184 0 -1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_49
timestamp 1679581782
transform 1 0 5856 0 -1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_56
timestamp 1679581782
transform 1 0 6528 0 -1 3024
box -48 -56 720 834
use sg13g2_fill_1  FILLER_1_63
timestamp 1677579658
transform 1 0 7200 0 -1 3024
box -48 -56 144 834
use sg13g2_fill_1  FILLER_1_85
timestamp 1677579658
transform 1 0 9312 0 -1 3024
box -48 -56 144 834
use sg13g2_decap_8  FILLER_1_103
timestamp 1679581782
transform 1 0 11040 0 -1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_110
timestamp 1679581782
transform 1 0 11712 0 -1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_117
timestamp 1679581782
transform 1 0 12384 0 -1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_124
timestamp 1679581782
transform 1 0 13056 0 -1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_135
timestamp 1679581782
transform 1 0 14112 0 -1 3024
box -48 -56 720 834
use sg13g2_decap_4  FILLER_1_142
timestamp 1679577901
transform 1 0 14784 0 -1 3024
box -48 -56 432 834
use sg13g2_fill_2  FILLER_1_146
timestamp 1677580104
transform 1 0 15168 0 -1 3024
box -48 -56 240 834
use sg13g2_decap_8  FILLER_1_158
timestamp 1679581782
transform 1 0 16320 0 -1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_165
timestamp 1679581782
transform 1 0 16992 0 -1 3024
box -48 -56 720 834
use sg13g2_decap_4  FILLER_1_172
timestamp 1679577901
transform 1 0 17664 0 -1 3024
box -48 -56 432 834
use sg13g2_fill_1  FILLER_1_197
timestamp 1677579658
transform 1 0 20064 0 -1 3024
box -48 -56 144 834
use sg13g2_decap_8  FILLER_1_202
timestamp 1679581782
transform 1 0 20544 0 -1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_209
timestamp 1679581782
transform 1 0 21216 0 -1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_216
timestamp 1679581782
transform 1 0 21888 0 -1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_223
timestamp 1679581782
transform 1 0 22560 0 -1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_230
timestamp 1679581782
transform 1 0 23232 0 -1 3024
box -48 -56 720 834
use sg13g2_fill_2  FILLER_1_237
timestamp 1677580104
transform 1 0 23904 0 -1 3024
box -48 -56 240 834
use sg13g2_fill_1  FILLER_1_239
timestamp 1677579658
transform 1 0 24096 0 -1 3024
box -48 -56 144 834
use sg13g2_decap_8  FILLER_1_244
timestamp 1679581782
transform 1 0 24576 0 -1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_251
timestamp 1679581782
transform 1 0 25248 0 -1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_258
timestamp 1679581782
transform 1 0 25920 0 -1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_265
timestamp 1679581782
transform 1 0 26592 0 -1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_272
timestamp 1679581782
transform 1 0 27264 0 -1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_279
timestamp 1679581782
transform 1 0 27936 0 -1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_286
timestamp 1679581782
transform 1 0 28608 0 -1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_293
timestamp 1679581782
transform 1 0 29280 0 -1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_300
timestamp 1679581782
transform 1 0 29952 0 -1 3024
box -48 -56 720 834
use sg13g2_decap_4  FILLER_1_307
timestamp 1679577901
transform 1 0 30624 0 -1 3024
box -48 -56 432 834
use sg13g2_decap_8  FILLER_1_323
timestamp 1679581782
transform 1 0 32160 0 -1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_330
timestamp 1679581782
transform 1 0 32832 0 -1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_337
timestamp 1679581782
transform 1 0 33504 0 -1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_344
timestamp 1679581782
transform 1 0 34176 0 -1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_351
timestamp 1679581782
transform 1 0 34848 0 -1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_358
timestamp 1679581782
transform 1 0 35520 0 -1 3024
box -48 -56 720 834
use sg13g2_fill_1  FILLER_1_365
timestamp 1677579658
transform 1 0 36192 0 -1 3024
box -48 -56 144 834
use sg13g2_decap_8  FILLER_1_370
timestamp 1679581782
transform 1 0 36672 0 -1 3024
box -48 -56 720 834
use sg13g2_fill_1  FILLER_1_377
timestamp 1677579658
transform 1 0 37344 0 -1 3024
box -48 -56 144 834
use sg13g2_fill_2  FILLER_1_393
timestamp 1677580104
transform 1 0 38880 0 -1 3024
box -48 -56 240 834
use sg13g2_decap_8  FILLER_1_419
timestamp 1679581782
transform 1 0 41376 0 -1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_426
timestamp 1679581782
transform 1 0 42048 0 -1 3024
box -48 -56 720 834
use sg13g2_fill_1  FILLER_1_433
timestamp 1677579658
transform 1 0 42720 0 -1 3024
box -48 -56 144 834
use sg13g2_decap_8  FILLER_1_438
timestamp 1679581782
transform 1 0 43200 0 -1 3024
box -48 -56 720 834
use sg13g2_fill_2  FILLER_1_445
timestamp 1677580104
transform 1 0 43872 0 -1 3024
box -48 -56 240 834
use sg13g2_decap_8  FILLER_2_0
timestamp 1679581782
transform 1 0 1152 0 1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_7
timestamp 1679581782
transform 1 0 1824 0 1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_14
timestamp 1679581782
transform 1 0 2496 0 1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_21
timestamp 1679581782
transform 1 0 3168 0 1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_28
timestamp 1679581782
transform 1 0 3840 0 1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_35
timestamp 1679581782
transform 1 0 4512 0 1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_42
timestamp 1679581782
transform 1 0 5184 0 1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_49
timestamp 1679581782
transform 1 0 5856 0 1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_56
timestamp 1679581782
transform 1 0 6528 0 1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_63
timestamp 1679581782
transform 1 0 7200 0 1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_70
timestamp 1679581782
transform 1 0 7872 0 1 3024
box -48 -56 720 834
use sg13g2_decap_4  FILLER_2_77
timestamp 1679577901
transform 1 0 8544 0 1 3024
box -48 -56 432 834
use sg13g2_decap_4  FILLER_2_106
timestamp 1679577901
transform 1 0 11328 0 1 3024
box -48 -56 432 834
use sg13g2_fill_1  FILLER_2_206
timestamp 1677579658
transform 1 0 20928 0 1 3024
box -48 -56 144 834
use sg13g2_decap_8  FILLER_2_217
timestamp 1679581782
transform 1 0 21984 0 1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_224
timestamp 1679581782
transform 1 0 22656 0 1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_231
timestamp 1679581782
transform 1 0 23328 0 1 3024
box -48 -56 720 834
use sg13g2_fill_2  FILLER_2_238
timestamp 1677580104
transform 1 0 24000 0 1 3024
box -48 -56 240 834
use sg13g2_fill_2  FILLER_2_257
timestamp 1677580104
transform 1 0 25824 0 1 3024
box -48 -56 240 834
use sg13g2_fill_2  FILLER_2_273
timestamp 1677580104
transform 1 0 27360 0 1 3024
box -48 -56 240 834
use sg13g2_decap_4  FILLER_2_296
timestamp 1679577901
transform 1 0 29568 0 1 3024
box -48 -56 432 834
use sg13g2_fill_2  FILLER_2_300
timestamp 1677580104
transform 1 0 29952 0 1 3024
box -48 -56 240 834
use sg13g2_decap_8  FILLER_2_339
timestamp 1679581782
transform 1 0 33696 0 1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_346
timestamp 1679581782
transform 1 0 34368 0 1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_353
timestamp 1679581782
transform 1 0 35040 0 1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_360
timestamp 1679581782
transform 1 0 35712 0 1 3024
box -48 -56 720 834
use sg13g2_decap_4  FILLER_2_367
timestamp 1679577901
transform 1 0 36384 0 1 3024
box -48 -56 432 834
use sg13g2_fill_1  FILLER_2_371
timestamp 1677579658
transform 1 0 36768 0 1 3024
box -48 -56 144 834
use sg13g2_fill_2  FILLER_2_392
timestamp 1677580104
transform 1 0 38784 0 1 3024
box -48 -56 240 834
use sg13g2_decap_8  FILLER_2_405
timestamp 1679581782
transform 1 0 40032 0 1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_412
timestamp 1679581782
transform 1 0 40704 0 1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_419
timestamp 1679581782
transform 1 0 41376 0 1 3024
box -48 -56 720 834
use sg13g2_fill_2  FILLER_2_426
timestamp 1677580104
transform 1 0 42048 0 1 3024
box -48 -56 240 834
use sg13g2_fill_1  FILLER_2_432
timestamp 1677579658
transform 1 0 42624 0 1 3024
box -48 -56 144 834
use sg13g2_fill_2  FILLER_2_449
timestamp 1677580104
transform 1 0 44256 0 1 3024
box -48 -56 240 834
use sg13g2_decap_8  FILLER_3_0
timestamp 1679581782
transform 1 0 1152 0 -1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_7
timestamp 1679581782
transform 1 0 1824 0 -1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_14
timestamp 1679581782
transform 1 0 2496 0 -1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_21
timestamp 1679581782
transform 1 0 3168 0 -1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_28
timestamp 1679581782
transform 1 0 3840 0 -1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_35
timestamp 1679581782
transform 1 0 4512 0 -1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_42
timestamp 1679581782
transform 1 0 5184 0 -1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_49
timestamp 1679581782
transform 1 0 5856 0 -1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_56
timestamp 1679581782
transform 1 0 6528 0 -1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_63
timestamp 1679581782
transform 1 0 7200 0 -1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_70
timestamp 1679581782
transform 1 0 7872 0 -1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_77
timestamp 1679581782
transform 1 0 8544 0 -1 4536
box -48 -56 720 834
use sg13g2_fill_1  FILLER_3_84
timestamp 1677579658
transform 1 0 9216 0 -1 4536
box -48 -56 144 834
use sg13g2_decap_8  FILLER_3_95
timestamp 1679581782
transform 1 0 10272 0 -1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_102
timestamp 1679581782
transform 1 0 10944 0 -1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_109
timestamp 1679581782
transform 1 0 11616 0 -1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_116
timestamp 1679581782
transform 1 0 12288 0 -1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_123
timestamp 1679581782
transform 1 0 12960 0 -1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_130
timestamp 1679581782
transform 1 0 13632 0 -1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_137
timestamp 1679581782
transform 1 0 14304 0 -1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_144
timestamp 1679581782
transform 1 0 14976 0 -1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_151
timestamp 1679581782
transform 1 0 15648 0 -1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_158
timestamp 1679581782
transform 1 0 16320 0 -1 4536
box -48 -56 720 834
use sg13g2_decap_4  FILLER_3_165
timestamp 1679577901
transform 1 0 16992 0 -1 4536
box -48 -56 432 834
use sg13g2_fill_2  FILLER_3_169
timestamp 1677580104
transform 1 0 17376 0 -1 4536
box -48 -56 240 834
use sg13g2_fill_1  FILLER_3_192
timestamp 1677579658
transform 1 0 19584 0 -1 4536
box -48 -56 144 834
use sg13g2_decap_4  FILLER_3_201
timestamp 1679577901
transform 1 0 20448 0 -1 4536
box -48 -56 432 834
use sg13g2_fill_2  FILLER_3_205
timestamp 1677580104
transform 1 0 20832 0 -1 4536
box -48 -56 240 834
use sg13g2_decap_8  FILLER_3_228
timestamp 1679581782
transform 1 0 23040 0 -1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_274
timestamp 1679581782
transform 1 0 27456 0 -1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_281
timestamp 1679581782
transform 1 0 28128 0 -1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_288
timestamp 1679581782
transform 1 0 28800 0 -1 4536
box -48 -56 720 834
use sg13g2_decap_4  FILLER_3_295
timestamp 1679577901
transform 1 0 29472 0 -1 4536
box -48 -56 432 834
use sg13g2_fill_1  FILLER_3_299
timestamp 1677579658
transform 1 0 29856 0 -1 4536
box -48 -56 144 834
use sg13g2_decap_8  FILLER_3_348
timestamp 1679581782
transform 1 0 34560 0 -1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_355
timestamp 1679581782
transform 1 0 35232 0 -1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_362
timestamp 1679581782
transform 1 0 35904 0 -1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_369
timestamp 1679581782
transform 1 0 36576 0 -1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_376
timestamp 1679581782
transform 1 0 37248 0 -1 4536
box -48 -56 720 834
use sg13g2_fill_2  FILLER_3_383
timestamp 1677580104
transform 1 0 37920 0 -1 4536
box -48 -56 240 834
use sg13g2_fill_1  FILLER_3_385
timestamp 1677579658
transform 1 0 38112 0 -1 4536
box -48 -56 144 834
use sg13g2_decap_8  FILLER_3_393
timestamp 1679581782
transform 1 0 38880 0 -1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_400
timestamp 1679581782
transform 1 0 39552 0 -1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_407
timestamp 1679581782
transform 1 0 40224 0 -1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_414
timestamp 1679581782
transform 1 0 40896 0 -1 4536
box -48 -56 720 834
use sg13g2_decap_4  FILLER_3_421
timestamp 1679577901
transform 1 0 41568 0 -1 4536
box -48 -56 432 834
use sg13g2_decap_8  FILLER_4_0
timestamp 1679581782
transform 1 0 1152 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_7
timestamp 1679581782
transform 1 0 1824 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_14
timestamp 1679581782
transform 1 0 2496 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_21
timestamp 1679581782
transform 1 0 3168 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_28
timestamp 1679581782
transform 1 0 3840 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_35
timestamp 1679581782
transform 1 0 4512 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_42
timestamp 1679581782
transform 1 0 5184 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_49
timestamp 1679581782
transform 1 0 5856 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_56
timestamp 1679581782
transform 1 0 6528 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_63
timestamp 1679581782
transform 1 0 7200 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_70
timestamp 1679581782
transform 1 0 7872 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_77
timestamp 1679581782
transform 1 0 8544 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_84
timestamp 1679581782
transform 1 0 9216 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_91
timestamp 1679581782
transform 1 0 9888 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_98
timestamp 1679581782
transform 1 0 10560 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_105
timestamp 1679581782
transform 1 0 11232 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_112
timestamp 1679581782
transform 1 0 11904 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_119
timestamp 1679581782
transform 1 0 12576 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_126
timestamp 1679581782
transform 1 0 13248 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_133
timestamp 1679581782
transform 1 0 13920 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_140
timestamp 1679581782
transform 1 0 14592 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_147
timestamp 1679581782
transform 1 0 15264 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_154
timestamp 1679581782
transform 1 0 15936 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_161
timestamp 1679581782
transform 1 0 16608 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_168
timestamp 1679581782
transform 1 0 17280 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_175
timestamp 1679581782
transform 1 0 17952 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_182
timestamp 1679581782
transform 1 0 18624 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_189
timestamp 1679581782
transform 1 0 19296 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_196
timestamp 1679581782
transform 1 0 19968 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_203
timestamp 1679581782
transform 1 0 20640 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_210
timestamp 1679581782
transform 1 0 21312 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_217
timestamp 1679581782
transform 1 0 21984 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_224
timestamp 1679581782
transform 1 0 22656 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_231
timestamp 1679581782
transform 1 0 23328 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_238
timestamp 1679581782
transform 1 0 24000 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_245
timestamp 1679581782
transform 1 0 24672 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_252
timestamp 1679581782
transform 1 0 25344 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_259
timestamp 1679581782
transform 1 0 26016 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_266
timestamp 1679581782
transform 1 0 26688 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_273
timestamp 1679581782
transform 1 0 27360 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_280
timestamp 1679581782
transform 1 0 28032 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_287
timestamp 1679581782
transform 1 0 28704 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_294
timestamp 1679581782
transform 1 0 29376 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_301
timestamp 1679581782
transform 1 0 30048 0 1 4536
box -48 -56 720 834
use sg13g2_fill_2  FILLER_4_308
timestamp 1677580104
transform 1 0 30720 0 1 4536
box -48 -56 240 834
use sg13g2_decap_8  FILLER_4_335
timestamp 1679581782
transform 1 0 33312 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_342
timestamp 1679581782
transform 1 0 33984 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_349
timestamp 1679581782
transform 1 0 34656 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_356
timestamp 1679581782
transform 1 0 35328 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_363
timestamp 1679581782
transform 1 0 36000 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_370
timestamp 1679581782
transform 1 0 36672 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_377
timestamp 1679581782
transform 1 0 37344 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_384
timestamp 1679581782
transform 1 0 38016 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_391
timestamp 1679581782
transform 1 0 38688 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_398
timestamp 1679581782
transform 1 0 39360 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_405
timestamp 1679581782
transform 1 0 40032 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_412
timestamp 1679581782
transform 1 0 40704 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_419
timestamp 1679581782
transform 1 0 41376 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_426
timestamp 1679581782
transform 1 0 42048 0 1 4536
box -48 -56 720 834
use sg13g2_fill_1  FILLER_4_433
timestamp 1677579658
transform 1 0 42720 0 1 4536
box -48 -56 144 834
use sg13g2_fill_1  FILLER_4_438
timestamp 1677579658
transform 1 0 43200 0 1 4536
box -48 -56 144 834
use sg13g2_decap_8  FILLER_5_12
timestamp 1679581782
transform 1 0 2304 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_19
timestamp 1679581782
transform 1 0 2976 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_26
timestamp 1679581782
transform 1 0 3648 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_33
timestamp 1679581782
transform 1 0 4320 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_40
timestamp 1679581782
transform 1 0 4992 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_47
timestamp 1679581782
transform 1 0 5664 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_54
timestamp 1679581782
transform 1 0 6336 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_61
timestamp 1679581782
transform 1 0 7008 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_68
timestamp 1679581782
transform 1 0 7680 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_75
timestamp 1679581782
transform 1 0 8352 0 -1 6048
box -48 -56 720 834
use sg13g2_fill_2  FILLER_5_82
timestamp 1677580104
transform 1 0 9024 0 -1 6048
box -48 -56 240 834
use sg13g2_decap_8  FILLER_5_109
timestamp 1679581782
transform 1 0 11616 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_116
timestamp 1679581782
transform 1 0 12288 0 -1 6048
box -48 -56 720 834
use sg13g2_fill_2  FILLER_5_123
timestamp 1677580104
transform 1 0 12960 0 -1 6048
box -48 -56 240 834
use sg13g2_decap_8  FILLER_5_128
timestamp 1679581782
transform 1 0 13440 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_135
timestamp 1679581782
transform 1 0 14112 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_142
timestamp 1679581782
transform 1 0 14784 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_149
timestamp 1679581782
transform 1 0 15456 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_156
timestamp 1679581782
transform 1 0 16128 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_163
timestamp 1679581782
transform 1 0 16800 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_170
timestamp 1679581782
transform 1 0 17472 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_177
timestamp 1679581782
transform 1 0 18144 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_184
timestamp 1679581782
transform 1 0 18816 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_191
timestamp 1679581782
transform 1 0 19488 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_198
timestamp 1679581782
transform 1 0 20160 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_205
timestamp 1679581782
transform 1 0 20832 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_212
timestamp 1679581782
transform 1 0 21504 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_219
timestamp 1679581782
transform 1 0 22176 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_226
timestamp 1679581782
transform 1 0 22848 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_233
timestamp 1679581782
transform 1 0 23520 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_240
timestamp 1679581782
transform 1 0 24192 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_247
timestamp 1679581782
transform 1 0 24864 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_254
timestamp 1679581782
transform 1 0 25536 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_261
timestamp 1679581782
transform 1 0 26208 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_268
timestamp 1679581782
transform 1 0 26880 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_275
timestamp 1679581782
transform 1 0 27552 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_282
timestamp 1679581782
transform 1 0 28224 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_289
timestamp 1679581782
transform 1 0 28896 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_296
timestamp 1679581782
transform 1 0 29568 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_303
timestamp 1679581782
transform 1 0 30240 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_310
timestamp 1679581782
transform 1 0 30912 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_317
timestamp 1679581782
transform 1 0 31584 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_324
timestamp 1679581782
transform 1 0 32256 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_331
timestamp 1679581782
transform 1 0 32928 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_338
timestamp 1679581782
transform 1 0 33600 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_345
timestamp 1679581782
transform 1 0 34272 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_352
timestamp 1679581782
transform 1 0 34944 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_359
timestamp 1679581782
transform 1 0 35616 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_366
timestamp 1679581782
transform 1 0 36288 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_373
timestamp 1679581782
transform 1 0 36960 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_380
timestamp 1679581782
transform 1 0 37632 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_387
timestamp 1679581782
transform 1 0 38304 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_394
timestamp 1679581782
transform 1 0 38976 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_401
timestamp 1679581782
transform 1 0 39648 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_408
timestamp 1679581782
transform 1 0 40320 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_415
timestamp 1679581782
transform 1 0 40992 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_422
timestamp 1679581782
transform 1 0 41664 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_429
timestamp 1679581782
transform 1 0 42336 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_4  FILLER_5_436
timestamp 1679577901
transform 1 0 43008 0 -1 6048
box -48 -56 432 834
use sg13g2_fill_2  FILLER_5_440
timestamp 1677580104
transform 1 0 43392 0 -1 6048
box -48 -56 240 834
use sg13g2_decap_8  FILLER_6_8
timestamp 1679581782
transform 1 0 1920 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_15
timestamp 1679581782
transform 1 0 2592 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_22
timestamp 1679581782
transform 1 0 3264 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_29
timestamp 1679581782
transform 1 0 3936 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_36
timestamp 1679581782
transform 1 0 4608 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_43
timestamp 1679581782
transform 1 0 5280 0 1 6048
box -48 -56 720 834
use sg13g2_fill_1  FILLER_6_50
timestamp 1677579658
transform 1 0 5952 0 1 6048
box -48 -56 144 834
use sg13g2_decap_8  FILLER_6_72
timestamp 1679581782
transform 1 0 8064 0 1 6048
box -48 -56 720 834
use sg13g2_fill_2  FILLER_6_79
timestamp 1677580104
transform 1 0 8736 0 1 6048
box -48 -56 240 834
use sg13g2_decap_8  FILLER_6_116
timestamp 1679581782
transform 1 0 12288 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_123
timestamp 1679581782
transform 1 0 12960 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_130
timestamp 1679581782
transform 1 0 13632 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_137
timestamp 1679581782
transform 1 0 14304 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_144
timestamp 1679581782
transform 1 0 14976 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_151
timestamp 1679581782
transform 1 0 15648 0 1 6048
box -48 -56 720 834
use sg13g2_decap_4  FILLER_6_158
timestamp 1679577901
transform 1 0 16320 0 1 6048
box -48 -56 432 834
use sg13g2_fill_2  FILLER_6_162
timestamp 1677580104
transform 1 0 16704 0 1 6048
box -48 -56 240 834
use sg13g2_decap_8  FILLER_6_168
timestamp 1679581782
transform 1 0 17280 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_175
timestamp 1679581782
transform 1 0 17952 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_182
timestamp 1679581782
transform 1 0 18624 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_189
timestamp 1679581782
transform 1 0 19296 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_196
timestamp 1679581782
transform 1 0 19968 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_203
timestamp 1679581782
transform 1 0 20640 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_210
timestamp 1679581782
transform 1 0 21312 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_217
timestamp 1679581782
transform 1 0 21984 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_224
timestamp 1679581782
transform 1 0 22656 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_231
timestamp 1679581782
transform 1 0 23328 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_238
timestamp 1679581782
transform 1 0 24000 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_245
timestamp 1679581782
transform 1 0 24672 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_252
timestamp 1679581782
transform 1 0 25344 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_259
timestamp 1679581782
transform 1 0 26016 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_266
timestamp 1679581782
transform 1 0 26688 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_273
timestamp 1679581782
transform 1 0 27360 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_280
timestamp 1679581782
transform 1 0 28032 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_287
timestamp 1679581782
transform 1 0 28704 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_294
timestamp 1679581782
transform 1 0 29376 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_301
timestamp 1679581782
transform 1 0 30048 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_308
timestamp 1679581782
transform 1 0 30720 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_315
timestamp 1679581782
transform 1 0 31392 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_322
timestamp 1679581782
transform 1 0 32064 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_329
timestamp 1679581782
transform 1 0 32736 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_336
timestamp 1679581782
transform 1 0 33408 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_343
timestamp 1679581782
transform 1 0 34080 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_350
timestamp 1679581782
transform 1 0 34752 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_357
timestamp 1679581782
transform 1 0 35424 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_364
timestamp 1679581782
transform 1 0 36096 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_371
timestamp 1679581782
transform 1 0 36768 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_378
timestamp 1679581782
transform 1 0 37440 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_385
timestamp 1679581782
transform 1 0 38112 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_392
timestamp 1679581782
transform 1 0 38784 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_399
timestamp 1679581782
transform 1 0 39456 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_406
timestamp 1679581782
transform 1 0 40128 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_413
timestamp 1679581782
transform 1 0 40800 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_420
timestamp 1679581782
transform 1 0 41472 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_427
timestamp 1679581782
transform 1 0 42144 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_434
timestamp 1679581782
transform 1 0 42816 0 1 6048
box -48 -56 720 834
use sg13g2_fill_1  FILLER_6_441
timestamp 1677579658
transform 1 0 43488 0 1 6048
box -48 -56 144 834
use sg13g2_fill_1  FILLER_6_458
timestamp 1677579658
transform 1 0 45120 0 1 6048
box -48 -56 144 834
use sg13g2_decap_8  FILLER_7_8
timestamp 1679581782
transform 1 0 1920 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_15
timestamp 1679581782
transform 1 0 2592 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_22
timestamp 1679581782
transform 1 0 3264 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_29
timestamp 1679581782
transform 1 0 3936 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_36
timestamp 1679581782
transform 1 0 4608 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_43
timestamp 1679581782
transform 1 0 5280 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_50
timestamp 1679581782
transform 1 0 5952 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_57
timestamp 1679581782
transform 1 0 6624 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_64
timestamp 1679581782
transform 1 0 7296 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_71
timestamp 1679581782
transform 1 0 7968 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_78
timestamp 1679581782
transform 1 0 8640 0 -1 7560
box -48 -56 720 834
use sg13g2_fill_2  FILLER_7_85
timestamp 1677580104
transform 1 0 9312 0 -1 7560
box -48 -56 240 834
use sg13g2_fill_1  FILLER_7_87
timestamp 1677579658
transform 1 0 9504 0 -1 7560
box -48 -56 144 834
use sg13g2_fill_1  FILLER_7_102
timestamp 1677579658
transform 1 0 10944 0 -1 7560
box -48 -56 144 834
use sg13g2_fill_2  FILLER_7_107
timestamp 1677580104
transform 1 0 11424 0 -1 7560
box -48 -56 240 834
use sg13g2_decap_8  FILLER_7_125
timestamp 1679581782
transform 1 0 13152 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_132
timestamp 1679581782
transform 1 0 13824 0 -1 7560
box -48 -56 720 834
use sg13g2_fill_2  FILLER_7_139
timestamp 1677580104
transform 1 0 14496 0 -1 7560
box -48 -56 240 834
use sg13g2_fill_1  FILLER_7_141
timestamp 1677579658
transform 1 0 14688 0 -1 7560
box -48 -56 144 834
use sg13g2_decap_8  FILLER_7_159
timestamp 1679581782
transform 1 0 16416 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_166
timestamp 1679581782
transform 1 0 17088 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_173
timestamp 1679581782
transform 1 0 17760 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_180
timestamp 1679581782
transform 1 0 18432 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_187
timestamp 1679581782
transform 1 0 19104 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_194
timestamp 1679581782
transform 1 0 19776 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_201
timestamp 1679581782
transform 1 0 20448 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_4  FILLER_7_208
timestamp 1679577901
transform 1 0 21120 0 -1 7560
box -48 -56 432 834
use sg13g2_fill_1  FILLER_7_212
timestamp 1677579658
transform 1 0 21504 0 -1 7560
box -48 -56 144 834
use sg13g2_decap_8  FILLER_7_217
timestamp 1679581782
transform 1 0 21984 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_4  FILLER_7_224
timestamp 1679577901
transform 1 0 22656 0 -1 7560
box -48 -56 432 834
use sg13g2_fill_2  FILLER_7_228
timestamp 1677580104
transform 1 0 23040 0 -1 7560
box -48 -56 240 834
use sg13g2_decap_8  FILLER_7_247
timestamp 1679581782
transform 1 0 24864 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_4  FILLER_7_254
timestamp 1679577901
transform 1 0 25536 0 -1 7560
box -48 -56 432 834
use sg13g2_fill_2  FILLER_7_258
timestamp 1677580104
transform 1 0 25920 0 -1 7560
box -48 -56 240 834
use sg13g2_decap_4  FILLER_7_285
timestamp 1679577901
transform 1 0 28512 0 -1 7560
box -48 -56 432 834
use sg13g2_fill_2  FILLER_7_289
timestamp 1677580104
transform 1 0 28896 0 -1 7560
box -48 -56 240 834
use sg13g2_decap_8  FILLER_7_308
timestamp 1679581782
transform 1 0 30720 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_315
timestamp 1679581782
transform 1 0 31392 0 -1 7560
box -48 -56 720 834
use sg13g2_fill_2  FILLER_7_322
timestamp 1677580104
transform 1 0 32064 0 -1 7560
box -48 -56 240 834
use sg13g2_decap_8  FILLER_7_385
timestamp 1679581782
transform 1 0 38112 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_392
timestamp 1679581782
transform 1 0 38784 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_399
timestamp 1679581782
transform 1 0 39456 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_406
timestamp 1679581782
transform 1 0 40128 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_413
timestamp 1679581782
transform 1 0 40800 0 -1 7560
box -48 -56 720 834
use sg13g2_fill_2  FILLER_7_420
timestamp 1677580104
transform 1 0 41472 0 -1 7560
box -48 -56 240 834
use sg13g2_decap_4  FILLER_8_8
timestamp 1679577901
transform 1 0 1920 0 1 7560
box -48 -56 432 834
use sg13g2_fill_1  FILLER_8_12
timestamp 1677579658
transform 1 0 2304 0 1 7560
box -48 -56 144 834
use sg13g2_decap_8  FILLER_8_37
timestamp 1679581782
transform 1 0 4704 0 1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_44
timestamp 1679581782
transform 1 0 5376 0 1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_51
timestamp 1679581782
transform 1 0 6048 0 1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_58
timestamp 1679581782
transform 1 0 6720 0 1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_65
timestamp 1679581782
transform 1 0 7392 0 1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_72
timestamp 1679581782
transform 1 0 8064 0 1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_79
timestamp 1679581782
transform 1 0 8736 0 1 7560
box -48 -56 720 834
use sg13g2_fill_2  FILLER_8_86
timestamp 1677580104
transform 1 0 9408 0 1 7560
box -48 -56 240 834
use sg13g2_decap_8  FILLER_8_122
timestamp 1679581782
transform 1 0 12864 0 1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_129
timestamp 1679581782
transform 1 0 13536 0 1 7560
box -48 -56 720 834
use sg13g2_fill_2  FILLER_8_136
timestamp 1677580104
transform 1 0 14208 0 1 7560
box -48 -56 240 834
use sg13g2_decap_4  FILLER_8_159
timestamp 1679577901
transform 1 0 16416 0 1 7560
box -48 -56 432 834
use sg13g2_fill_1  FILLER_8_163
timestamp 1677579658
transform 1 0 16800 0 1 7560
box -48 -56 144 834
use sg13g2_decap_4  FILLER_8_168
timestamp 1679577901
transform 1 0 17280 0 1 7560
box -48 -56 432 834
use sg13g2_fill_2  FILLER_8_172
timestamp 1677580104
transform 1 0 17664 0 1 7560
box -48 -56 240 834
use sg13g2_decap_8  FILLER_8_178
timestamp 1679581782
transform 1 0 18240 0 1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_185
timestamp 1679581782
transform 1 0 18912 0 1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_192
timestamp 1679581782
transform 1 0 19584 0 1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_199
timestamp 1679581782
transform 1 0 20256 0 1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_206
timestamp 1679581782
transform 1 0 20928 0 1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_213
timestamp 1679581782
transform 1 0 21600 0 1 7560
box -48 -56 720 834
use sg13g2_fill_2  FILLER_8_220
timestamp 1677580104
transform 1 0 22272 0 1 7560
box -48 -56 240 834
use sg13g2_fill_1  FILLER_8_222
timestamp 1677579658
transform 1 0 22464 0 1 7560
box -48 -56 144 834
use sg13g2_decap_8  FILLER_8_248
timestamp 1679581782
transform 1 0 24960 0 1 7560
box -48 -56 720 834
use sg13g2_fill_2  FILLER_8_255
timestamp 1677580104
transform 1 0 25632 0 1 7560
box -48 -56 240 834
use sg13g2_decap_4  FILLER_8_290
timestamp 1679577901
transform 1 0 28992 0 1 7560
box -48 -56 432 834
use sg13g2_decap_8  FILLER_8_298
timestamp 1679581782
transform 1 0 29760 0 1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_305
timestamp 1679581782
transform 1 0 30432 0 1 7560
box -48 -56 720 834
use sg13g2_decap_4  FILLER_8_312
timestamp 1679577901
transform 1 0 31104 0 1 7560
box -48 -56 432 834
use sg13g2_fill_2  FILLER_8_323
timestamp 1677580104
transform 1 0 32160 0 1 7560
box -48 -56 240 834
use sg13g2_fill_1  FILLER_8_332
timestamp 1677579658
transform 1 0 33024 0 1 7560
box -48 -56 144 834
use sg13g2_decap_8  FILLER_8_356
timestamp 1679581782
transform 1 0 35328 0 1 7560
box -48 -56 720 834
use sg13g2_fill_1  FILLER_8_363
timestamp 1677579658
transform 1 0 36000 0 1 7560
box -48 -56 144 834
use sg13g2_decap_8  FILLER_8_374
timestamp 1679581782
transform 1 0 37056 0 1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_381
timestamp 1679581782
transform 1 0 37728 0 1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_388
timestamp 1679581782
transform 1 0 38400 0 1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_395
timestamp 1679581782
transform 1 0 39072 0 1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_402
timestamp 1679581782
transform 1 0 39744 0 1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_409
timestamp 1679581782
transform 1 0 40416 0 1 7560
box -48 -56 720 834
use sg13g2_decap_4  FILLER_8_416
timestamp 1679577901
transform 1 0 41088 0 1 7560
box -48 -56 432 834
use sg13g2_fill_1  FILLER_8_420
timestamp 1677579658
transform 1 0 41472 0 1 7560
box -48 -56 144 834
use sg13g2_fill_2  FILLER_8_449
timestamp 1677580104
transform 1 0 44256 0 1 7560
box -48 -56 240 834
use sg13g2_decap_8  FILLER_9_16
timestamp 1679581782
transform 1 0 2688 0 -1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_23
timestamp 1679581782
transform 1 0 3360 0 -1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_30
timestamp 1679581782
transform 1 0 4032 0 -1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_37
timestamp 1679581782
transform 1 0 4704 0 -1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_44
timestamp 1679581782
transform 1 0 5376 0 -1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_51
timestamp 1679581782
transform 1 0 6048 0 -1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_58
timestamp 1679581782
transform 1 0 6720 0 -1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_65
timestamp 1679581782
transform 1 0 7392 0 -1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_72
timestamp 1679581782
transform 1 0 8064 0 -1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_79
timestamp 1679581782
transform 1 0 8736 0 -1 9072
box -48 -56 720 834
use sg13g2_fill_2  FILLER_9_86
timestamp 1677580104
transform 1 0 9408 0 -1 9072
box -48 -56 240 834
use sg13g2_fill_2  FILLER_9_113
timestamp 1677580104
transform 1 0 12000 0 -1 9072
box -48 -56 240 834
use sg13g2_decap_8  FILLER_9_219
timestamp 1679581782
transform 1 0 22176 0 -1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_226
timestamp 1679581782
transform 1 0 22848 0 -1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_237
timestamp 1679581782
transform 1 0 23904 0 -1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_244
timestamp 1679581782
transform 1 0 24576 0 -1 9072
box -48 -56 720 834
use sg13g2_fill_1  FILLER_9_271
timestamp 1677579658
transform 1 0 27168 0 -1 9072
box -48 -56 144 834
use sg13g2_decap_4  FILLER_9_286
timestamp 1679577901
transform 1 0 28608 0 -1 9072
box -48 -56 432 834
use sg13g2_fill_1  FILLER_9_290
timestamp 1677579658
transform 1 0 28992 0 -1 9072
box -48 -56 144 834
use sg13g2_decap_8  FILLER_9_299
timestamp 1679581782
transform 1 0 29856 0 -1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_306
timestamp 1679581782
transform 1 0 30528 0 -1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_313
timestamp 1679581782
transform 1 0 31200 0 -1 9072
box -48 -56 720 834
use sg13g2_fill_2  FILLER_9_320
timestamp 1677580104
transform 1 0 31872 0 -1 9072
box -48 -56 240 834
use sg13g2_fill_1  FILLER_9_322
timestamp 1677579658
transform 1 0 32064 0 -1 9072
box -48 -56 144 834
use sg13g2_decap_8  FILLER_9_355
timestamp 1679581782
transform 1 0 35232 0 -1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_362
timestamp 1679581782
transform 1 0 35904 0 -1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_369
timestamp 1679581782
transform 1 0 36576 0 -1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_376
timestamp 1679581782
transform 1 0 37248 0 -1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_383
timestamp 1679581782
transform 1 0 37920 0 -1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_390
timestamp 1679581782
transform 1 0 38592 0 -1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_397
timestamp 1679581782
transform 1 0 39264 0 -1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_404
timestamp 1679581782
transform 1 0 39936 0 -1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_411
timestamp 1679581782
transform 1 0 40608 0 -1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_418
timestamp 1679581782
transform 1 0 41280 0 -1 9072
box -48 -56 720 834
use sg13g2_decap_4  FILLER_9_425
timestamp 1679577901
transform 1 0 41952 0 -1 9072
box -48 -56 432 834
use sg13g2_fill_2  FILLER_9_445
timestamp 1677580104
transform 1 0 43872 0 -1 9072
box -48 -56 240 834
use sg13g2_decap_8  FILLER_10_24
timestamp 1679581782
transform 1 0 3456 0 1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_31
timestamp 1679581782
transform 1 0 4128 0 1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_38
timestamp 1679581782
transform 1 0 4800 0 1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_45
timestamp 1679581782
transform 1 0 5472 0 1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_52
timestamp 1679581782
transform 1 0 6144 0 1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_59
timestamp 1679581782
transform 1 0 6816 0 1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_66
timestamp 1679581782
transform 1 0 7488 0 1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_73
timestamp 1679581782
transform 1 0 8160 0 1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_80
timestamp 1679581782
transform 1 0 8832 0 1 9072
box -48 -56 720 834
use sg13g2_decap_4  FILLER_10_87
timestamp 1679577901
transform 1 0 9504 0 1 9072
box -48 -56 432 834
use sg13g2_fill_2  FILLER_10_227
timestamp 1677580104
transform 1 0 22944 0 1 9072
box -48 -56 240 834
use sg13g2_decap_4  FILLER_10_277
timestamp 1679577901
transform 1 0 27744 0 1 9072
box -48 -56 432 834
use sg13g2_decap_8  FILLER_10_305
timestamp 1679581782
transform 1 0 30432 0 1 9072
box -48 -56 720 834
use sg13g2_fill_1  FILLER_10_312
timestamp 1677579658
transform 1 0 31104 0 1 9072
box -48 -56 144 834
use sg13g2_decap_8  FILLER_10_365
timestamp 1679581782
transform 1 0 36192 0 1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_372
timestamp 1679581782
transform 1 0 36864 0 1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_379
timestamp 1679581782
transform 1 0 37536 0 1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_386
timestamp 1679581782
transform 1 0 38208 0 1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_393
timestamp 1679581782
transform 1 0 38880 0 1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_400
timestamp 1679581782
transform 1 0 39552 0 1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_407
timestamp 1679581782
transform 1 0 40224 0 1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_414
timestamp 1679581782
transform 1 0 40896 0 1 9072
box -48 -56 720 834
use sg13g2_fill_2  FILLER_10_421
timestamp 1677580104
transform 1 0 41568 0 1 9072
box -48 -56 240 834
use sg13g2_fill_1  FILLER_10_423
timestamp 1677579658
transform 1 0 41760 0 1 9072
box -48 -56 144 834
use sg13g2_fill_1  FILLER_10_435
timestamp 1677579658
transform 1 0 42912 0 1 9072
box -48 -56 144 834
use sg13g2_buf_1  input1
timestamp 1676381911
transform 1 0 2400 0 1 1512
box -48 -56 432 834
use sg13g2_buf_1  input2
timestamp 1676381911
transform 1 0 1920 0 -1 6048
box -48 -56 432 834
use sg13g2_buf_1  input3
timestamp 1676381911
transform 1 0 1536 0 -1 6048
box -48 -56 432 834
use sg13g2_buf_1  input4
timestamp 1676381911
transform 1 0 1152 0 -1 6048
box -48 -56 432 834
use sg13g2_buf_1  input5
timestamp 1676381911
transform 1 0 1536 0 1 6048
box -48 -56 432 834
use sg13g2_buf_1  input6
timestamp 1676381911
transform 1 0 1152 0 1 6048
box -48 -56 432 834
use sg13g2_buf_1  input7
timestamp 1676381911
transform 1 0 1536 0 -1 7560
box -48 -56 432 834
use sg13g2_buf_1  input8
timestamp 1676381911
transform 1 0 1152 0 -1 7560
box -48 -56 432 834
use sg13g2_buf_1  input9
timestamp 1676381911
transform 1 0 1152 0 1 7560
box -48 -56 432 834
use sg13g2_buf_1  input10
timestamp 1676381911
transform 1 0 1536 0 1 7560
box -48 -56 432 834
use sg13g2_buf_1  input11
timestamp 1676381911
transform 1 0 1152 0 -1 9072
box -48 -56 432 834
use sg13g2_buf_1  input12
timestamp 1676381911
transform 1 0 1536 0 -1 9072
box -48 -56 432 834
use sg13g2_buf_1  input13
timestamp 1676381911
transform 1 0 1920 0 -1 9072
box -48 -56 432 834
use sg13g2_buf_1  input14
timestamp 1676381911
transform 1 0 1152 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  input15
timestamp 1676381911
transform 1 0 1536 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  input16
timestamp 1676381911
transform 1 0 1920 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  input17
timestamp 1676381911
transform 1 0 2304 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  input18
timestamp 1676381911
transform 1 0 2688 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  input19
timestamp 1676381911
transform 1 0 2304 0 -1 9072
box -48 -56 432 834
use sg13g2_buf_1  input20
timestamp 1676381911
transform 1 0 3072 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  input21
timestamp 1676381911
transform 1 0 3936 0 1 1512
box -48 -56 432 834
use sg13g2_buf_1  input22
timestamp 1676381911
transform -1 0 21024 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  input23
timestamp 1676381911
transform 1 0 21408 0 -1 9072
box -48 -56 432 834
use sg13g2_buf_1  input24
timestamp 1676381911
transform 1 0 21024 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  input25
timestamp 1676381911
transform -1 0 22176 0 -1 9072
box -48 -56 432 834
use sg13g2_buf_1  input26
timestamp 1676381911
transform -1 0 23904 0 -1 9072
box -48 -56 432 834
use sg13g2_buf_1  input27
timestamp 1676381911
transform 1 0 23136 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  input28
timestamp 1676381911
transform 1 0 23520 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  input29
timestamp 1676381911
transform -1 0 24288 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  input30
timestamp 1676381911
transform -1 0 24672 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  input31
timestamp 1676381911
transform 1 0 24672 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  input32
timestamp 1676381911
transform 1 0 25056 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  input33
timestamp 1676381911
transform -1 0 25824 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  input34
timestamp 1676381911
transform -1 0 21792 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  input35
timestamp 1676381911
transform 1 0 21792 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  input36
timestamp 1676381911
transform 1 0 22176 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  input37
timestamp 1676381911
transform -1 0 22944 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  input38
timestamp 1676381911
transform -1 0 26208 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  input39
timestamp 1676381911
transform 1 0 25248 0 -1 9072
box -48 -56 432 834
use sg13g2_buf_1  input40
timestamp 1676381911
transform 1 0 26208 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  input41
timestamp 1676381911
transform -1 0 26016 0 -1 9072
box -48 -56 432 834
use sg13g2_buf_1  input42
timestamp 1676381911
transform -1 0 26976 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  input43
timestamp 1676381911
transform 1 0 26016 0 -1 9072
box -48 -56 432 834
use sg13g2_buf_1  input44
timestamp 1676381911
transform 1 0 26976 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  input45
timestamp 1676381911
transform -1 0 27744 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  input46
timestamp 1676381911
transform -1 0 28512 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  input47
timestamp 1676381911
transform 1 0 28512 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  input48
timestamp 1676381911
transform -1 0 29280 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  input49
timestamp 1676381911
transform -1 0 29664 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  input50
timestamp 1676381911
transform -1 0 30048 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  input51
timestamp 1676381911
transform 1 0 29088 0 -1 9072
box -48 -56 432 834
use sg13g2_buf_1  input52
timestamp 1676381911
transform -1 0 30432 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  input53
timestamp 1676381911
transform -1 0 29856 0 -1 9072
box -48 -56 432 834
use sg13g2_buf_1  output54
timestamp 1676381911
transform -1 0 5856 0 1 1512
box -48 -56 432 834
use sg13g2_buf_1  output55
timestamp 1676381911
transform 1 0 44064 0 1 1512
box -48 -56 432 834
use sg13g2_buf_1  output56
timestamp 1676381911
transform 1 0 44160 0 -1 4536
box -48 -56 432 834
use sg13g2_buf_1  output57
timestamp 1676381911
transform 1 0 44832 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  output58
timestamp 1676381911
transform 1 0 44448 0 1 4536
box -48 -56 432 834
use sg13g2_buf_1  output59
timestamp 1676381911
transform 1 0 44832 0 -1 4536
box -48 -56 432 834
use sg13g2_buf_1  output60
timestamp 1676381911
transform 1 0 44448 0 -1 6048
box -48 -56 432 834
use sg13g2_buf_1  output61
timestamp 1676381911
transform 1 0 44832 0 1 4536
box -48 -56 432 834
use sg13g2_buf_1  output62
timestamp 1676381911
transform 1 0 44448 0 1 6048
box -48 -56 432 834
use sg13g2_buf_1  output63
timestamp 1676381911
transform 1 0 44832 0 -1 6048
box -48 -56 432 834
use sg13g2_buf_1  output64
timestamp 1676381911
transform 1 0 44160 0 -1 7560
box -48 -56 432 834
use sg13g2_buf_1  output65
timestamp 1676381911
transform 1 0 44832 0 -1 7560
box -48 -56 432 834
use sg13g2_buf_1  output66
timestamp 1676381911
transform 1 0 43680 0 1 1512
box -48 -56 432 834
use sg13g2_buf_1  output67
timestamp 1676381911
transform 1 0 44832 0 1 7560
box -48 -56 432 834
use sg13g2_buf_1  output68
timestamp 1676381911
transform 1 0 44448 0 1 7560
box -48 -56 432 834
use sg13g2_buf_1  output69
timestamp 1676381911
transform 1 0 44832 0 -1 9072
box -48 -56 432 834
use sg13g2_buf_1  output70
timestamp 1676381911
transform 1 0 44448 0 -1 9072
box -48 -56 432 834
use sg13g2_buf_1  output71
timestamp 1676381911
transform 1 0 42144 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  output72
timestamp 1676381911
transform 1 0 43008 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  output73
timestamp 1676381911
transform 1 0 44832 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  output74
timestamp 1676381911
transform 1 0 44448 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  output75
timestamp 1676381911
transform 1 0 44064 0 -1 9072
box -48 -56 432 834
use sg13g2_buf_1  output76
timestamp 1676381911
transform 1 0 44064 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  output77
timestamp 1676381911
transform 1 0 43296 0 1 1512
box -48 -56 432 834
use sg13g2_buf_1  output78
timestamp 1676381911
transform 1 0 43680 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  output79
timestamp 1676381911
transform 1 0 42528 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  output80
timestamp 1676381911
transform 1 0 44448 0 1 1512
box -48 -56 432 834
use sg13g2_buf_1  output81
timestamp 1676381911
transform 1 0 44064 0 -1 3024
box -48 -56 432 834
use sg13g2_buf_1  output82
timestamp 1676381911
transform 1 0 42912 0 1 1512
box -48 -56 432 834
use sg13g2_buf_1  output83
timestamp 1676381911
transform 1 0 44448 0 -1 3024
box -48 -56 432 834
use sg13g2_buf_1  output84
timestamp 1676381911
transform 1 0 44832 0 1 1512
box -48 -56 432 834
use sg13g2_buf_1  output85
timestamp 1676381911
transform 1 0 44448 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  output86
timestamp 1676381911
transform 1 0 44832 0 -1 3024
box -48 -56 432 834
use sg13g2_buf_1  output87
timestamp 1676381911
transform -1 0 31968 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  output88
timestamp 1676381911
transform -1 0 33696 0 -1 9072
box -48 -56 432 834
use sg13g2_buf_1  output89
timestamp 1676381911
transform -1 0 34656 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  output90
timestamp 1676381911
transform -1 0 34080 0 -1 9072
box -48 -56 432 834
use sg13g2_buf_1  output91
timestamp 1676381911
transform -1 0 35040 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  output92
timestamp 1676381911
transform -1 0 34464 0 -1 9072
box -48 -56 432 834
use sg13g2_buf_1  output93
timestamp 1676381911
transform -1 0 35424 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  output94
timestamp 1676381911
transform -1 0 34848 0 -1 9072
box -48 -56 432 834
use sg13g2_buf_1  output95
timestamp 1676381911
transform -1 0 35808 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  output96
timestamp 1676381911
transform -1 0 35232 0 -1 9072
box -48 -56 432 834
use sg13g2_buf_1  output97
timestamp 1676381911
transform -1 0 36192 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  output98
timestamp 1676381911
transform -1 0 32352 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  output99
timestamp 1676381911
transform -1 0 32736 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  output100
timestamp 1676381911
transform -1 0 33120 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  output101
timestamp 1676381911
transform -1 0 32544 0 -1 9072
box -48 -56 432 834
use sg13g2_buf_1  output102
timestamp 1676381911
transform -1 0 33504 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  output103
timestamp 1676381911
transform -1 0 32928 0 -1 9072
box -48 -56 432 834
use sg13g2_buf_1  output104
timestamp 1676381911
transform -1 0 33888 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  output105
timestamp 1676381911
transform -1 0 33312 0 -1 9072
box -48 -56 432 834
use sg13g2_buf_1  output106
timestamp 1676381911
transform -1 0 34272 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  output107
timestamp 1676381911
transform 1 0 10368 0 -1 9072
box -48 -56 432 834
use sg13g2_buf_1  output108
timestamp 1676381911
transform 1 0 9888 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  output109
timestamp 1676381911
transform 1 0 10272 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  output110
timestamp 1676381911
transform 1 0 11136 0 -1 9072
box -48 -56 432 834
use sg13g2_buf_1  output111
timestamp 1676381911
transform 1 0 10656 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  output112
timestamp 1676381911
transform 1 0 11040 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  output113
timestamp 1676381911
transform -1 0 12576 0 -1 9072
box -48 -56 432 834
use sg13g2_buf_1  output114
timestamp 1676381911
transform 1 0 11424 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  output115
timestamp 1676381911
transform -1 0 12960 0 -1 9072
box -48 -56 432 834
use sg13g2_buf_1  output116
timestamp 1676381911
transform 1 0 11808 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  output117
timestamp 1676381911
transform -1 0 13344 0 -1 9072
box -48 -56 432 834
use sg13g2_buf_1  output118
timestamp 1676381911
transform 1 0 12192 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  output119
timestamp 1676381911
transform -1 0 13728 0 -1 9072
box -48 -56 432 834
use sg13g2_buf_1  output120
timestamp 1676381911
transform 1 0 12576 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  output121
timestamp 1676381911
transform -1 0 14112 0 -1 9072
box -48 -56 432 834
use sg13g2_buf_1  output122
timestamp 1676381911
transform 1 0 12960 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  output123
timestamp 1676381911
transform -1 0 14496 0 -1 9072
box -48 -56 432 834
use sg13g2_buf_1  output124
timestamp 1676381911
transform 1 0 13344 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  output125
timestamp 1676381911
transform -1 0 14880 0 -1 9072
box -48 -56 432 834
use sg13g2_buf_1  output126
timestamp 1676381911
transform 1 0 13728 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  output127
timestamp 1676381911
transform 1 0 14112 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  output128
timestamp 1676381911
transform -1 0 17184 0 -1 9072
box -48 -56 432 834
use sg13g2_buf_1  output129
timestamp 1676381911
transform 1 0 16416 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  output130
timestamp 1676381911
transform -1 0 17568 0 -1 9072
box -48 -56 432 834
use sg13g2_buf_1  output131
timestamp 1676381911
transform 1 0 16800 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  output132
timestamp 1676381911
transform -1 0 17952 0 -1 9072
box -48 -56 432 834
use sg13g2_buf_1  output133
timestamp 1676381911
transform 1 0 17184 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  output134
timestamp 1676381911
transform 1 0 14496 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  output135
timestamp 1676381911
transform -1 0 15648 0 -1 9072
box -48 -56 432 834
use sg13g2_buf_1  output136
timestamp 1676381911
transform 1 0 14880 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  output137
timestamp 1676381911
transform -1 0 16032 0 -1 9072
box -48 -56 432 834
use sg13g2_buf_1  output138
timestamp 1676381911
transform 1 0 15264 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  output139
timestamp 1676381911
transform -1 0 16416 0 -1 9072
box -48 -56 432 834
use sg13g2_buf_1  output140
timestamp 1676381911
transform 1 0 15648 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  output141
timestamp 1676381911
transform -1 0 16800 0 -1 9072
box -48 -56 432 834
use sg13g2_buf_1  output142
timestamp 1676381911
transform 1 0 16032 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  output143
timestamp 1676381911
transform -1 0 18336 0 -1 9072
box -48 -56 432 834
use sg13g2_buf_1  output144
timestamp 1676381911
transform -1 0 20256 0 -1 9072
box -48 -56 432 834
use sg13g2_buf_1  output145
timestamp 1676381911
transform 1 0 19488 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  output146
timestamp 1676381911
transform -1 0 20640 0 -1 9072
box -48 -56 432 834
use sg13g2_buf_1  output147
timestamp 1676381911
transform 1 0 19872 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  output148
timestamp 1676381911
transform -1 0 21024 0 -1 9072
box -48 -56 432 834
use sg13g2_buf_1  output149
timestamp 1676381911
transform 1 0 20256 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  output150
timestamp 1676381911
transform 1 0 17568 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  output151
timestamp 1676381911
transform -1 0 18720 0 -1 9072
box -48 -56 432 834
use sg13g2_buf_1  output152
timestamp 1676381911
transform 1 0 17952 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  output153
timestamp 1676381911
transform -1 0 19104 0 -1 9072
box -48 -56 432 834
use sg13g2_buf_1  output154
timestamp 1676381911
transform 1 0 18336 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  output155
timestamp 1676381911
transform -1 0 19488 0 -1 9072
box -48 -56 432 834
use sg13g2_buf_1  output156
timestamp 1676381911
transform 1 0 18720 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  output157
timestamp 1676381911
transform -1 0 19872 0 -1 9072
box -48 -56 432 834
use sg13g2_buf_1  output158
timestamp 1676381911
transform 1 0 19104 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  output159
timestamp 1676381911
transform -1 0 7392 0 1 1512
box -48 -56 432 834
use sg13g2_buf_1  output160
timestamp 1676381911
transform -1 0 8928 0 1 1512
box -48 -56 432 834
use sg13g2_buf_1  output161
timestamp 1676381911
transform -1 0 10464 0 1 1512
box -48 -56 432 834
use sg13g2_buf_1  output162
timestamp 1676381911
transform -1 0 12000 0 1 1512
box -48 -56 432 834
use sg13g2_buf_1  output163
timestamp 1676381911
transform -1 0 31584 0 1 9072
box -48 -56 432 834
use sg13g2_tielo  S_WARMBOOT_164
timestamp 1680000637
transform -1 0 21408 0 -1 9072
box -48 -56 432 834
<< labels >>
flabel metal3 s 5432 0 5512 80 0 FreeSans 320 0 0 0 BOOT_top
port 0 nsew signal output
flabel metal3 s 2360 0 2440 80 0 FreeSans 320 0 0 0 CONFIGURED_top
port 1 nsew signal input
flabel metal3 s 20984 11764 21064 11844 0 FreeSans 320 0 0 0 Co
port 2 nsew signal output
flabel metal2 s 0 548 90 628 0 FreeSans 320 0 0 0 FrameData[0]
port 3 nsew signal input
flabel metal2 s 0 3908 90 3988 0 FreeSans 320 0 0 0 FrameData[10]
port 4 nsew signal input
flabel metal2 s 0 4244 90 4324 0 FreeSans 320 0 0 0 FrameData[11]
port 5 nsew signal input
flabel metal2 s 0 4580 90 4660 0 FreeSans 320 0 0 0 FrameData[12]
port 6 nsew signal input
flabel metal2 s 0 4916 90 4996 0 FreeSans 320 0 0 0 FrameData[13]
port 7 nsew signal input
flabel metal2 s 0 5252 90 5332 0 FreeSans 320 0 0 0 FrameData[14]
port 8 nsew signal input
flabel metal2 s 0 5588 90 5668 0 FreeSans 320 0 0 0 FrameData[15]
port 9 nsew signal input
flabel metal2 s 0 5924 90 6004 0 FreeSans 320 0 0 0 FrameData[16]
port 10 nsew signal input
flabel metal2 s 0 6260 90 6340 0 FreeSans 320 0 0 0 FrameData[17]
port 11 nsew signal input
flabel metal2 s 0 6596 90 6676 0 FreeSans 320 0 0 0 FrameData[18]
port 12 nsew signal input
flabel metal2 s 0 6932 90 7012 0 FreeSans 320 0 0 0 FrameData[19]
port 13 nsew signal input
flabel metal2 s 0 884 90 964 0 FreeSans 320 0 0 0 FrameData[1]
port 14 nsew signal input
flabel metal2 s 0 7268 90 7348 0 FreeSans 320 0 0 0 FrameData[20]
port 15 nsew signal input
flabel metal2 s 0 7604 90 7684 0 FreeSans 320 0 0 0 FrameData[21]
port 16 nsew signal input
flabel metal2 s 0 7940 90 8020 0 FreeSans 320 0 0 0 FrameData[22]
port 17 nsew signal input
flabel metal2 s 0 8276 90 8356 0 FreeSans 320 0 0 0 FrameData[23]
port 18 nsew signal input
flabel metal2 s 0 8612 90 8692 0 FreeSans 320 0 0 0 FrameData[24]
port 19 nsew signal input
flabel metal2 s 0 8948 90 9028 0 FreeSans 320 0 0 0 FrameData[25]
port 20 nsew signal input
flabel metal2 s 0 9284 90 9364 0 FreeSans 320 0 0 0 FrameData[26]
port 21 nsew signal input
flabel metal2 s 0 9620 90 9700 0 FreeSans 320 0 0 0 FrameData[27]
port 22 nsew signal input
flabel metal2 s 0 9956 90 10036 0 FreeSans 320 0 0 0 FrameData[28]
port 23 nsew signal input
flabel metal2 s 0 10292 90 10372 0 FreeSans 320 0 0 0 FrameData[29]
port 24 nsew signal input
flabel metal2 s 0 1220 90 1300 0 FreeSans 320 0 0 0 FrameData[2]
port 25 nsew signal input
flabel metal2 s 0 10628 90 10708 0 FreeSans 320 0 0 0 FrameData[30]
port 26 nsew signal input
flabel metal2 s 0 10964 90 11044 0 FreeSans 320 0 0 0 FrameData[31]
port 27 nsew signal input
flabel metal2 s 0 1556 90 1636 0 FreeSans 320 0 0 0 FrameData[3]
port 28 nsew signal input
flabel metal2 s 0 1892 90 1972 0 FreeSans 320 0 0 0 FrameData[4]
port 29 nsew signal input
flabel metal2 s 0 2228 90 2308 0 FreeSans 320 0 0 0 FrameData[5]
port 30 nsew signal input
flabel metal2 s 0 2564 90 2644 0 FreeSans 320 0 0 0 FrameData[6]
port 31 nsew signal input
flabel metal2 s 0 2900 90 2980 0 FreeSans 320 0 0 0 FrameData[7]
port 32 nsew signal input
flabel metal2 s 0 3236 90 3316 0 FreeSans 320 0 0 0 FrameData[8]
port 33 nsew signal input
flabel metal2 s 0 3572 90 3652 0 FreeSans 320 0 0 0 FrameData[9]
port 34 nsew signal input
flabel metal2 s 46278 548 46368 628 0 FreeSans 320 0 0 0 FrameData_O[0]
port 35 nsew signal output
flabel metal2 s 46278 3908 46368 3988 0 FreeSans 320 0 0 0 FrameData_O[10]
port 36 nsew signal output
flabel metal2 s 46278 4244 46368 4324 0 FreeSans 320 0 0 0 FrameData_O[11]
port 37 nsew signal output
flabel metal2 s 46278 4580 46368 4660 0 FreeSans 320 0 0 0 FrameData_O[12]
port 38 nsew signal output
flabel metal2 s 46278 4916 46368 4996 0 FreeSans 320 0 0 0 FrameData_O[13]
port 39 nsew signal output
flabel metal2 s 46278 5252 46368 5332 0 FreeSans 320 0 0 0 FrameData_O[14]
port 40 nsew signal output
flabel metal2 s 46278 5588 46368 5668 0 FreeSans 320 0 0 0 FrameData_O[15]
port 41 nsew signal output
flabel metal2 s 46278 5924 46368 6004 0 FreeSans 320 0 0 0 FrameData_O[16]
port 42 nsew signal output
flabel metal2 s 46278 6260 46368 6340 0 FreeSans 320 0 0 0 FrameData_O[17]
port 43 nsew signal output
flabel metal2 s 46278 6596 46368 6676 0 FreeSans 320 0 0 0 FrameData_O[18]
port 44 nsew signal output
flabel metal2 s 46278 6932 46368 7012 0 FreeSans 320 0 0 0 FrameData_O[19]
port 45 nsew signal output
flabel metal2 s 46278 884 46368 964 0 FreeSans 320 0 0 0 FrameData_O[1]
port 46 nsew signal output
flabel metal2 s 46278 7268 46368 7348 0 FreeSans 320 0 0 0 FrameData_O[20]
port 47 nsew signal output
flabel metal2 s 46278 7604 46368 7684 0 FreeSans 320 0 0 0 FrameData_O[21]
port 48 nsew signal output
flabel metal2 s 46278 7940 46368 8020 0 FreeSans 320 0 0 0 FrameData_O[22]
port 49 nsew signal output
flabel metal2 s 46278 8276 46368 8356 0 FreeSans 320 0 0 0 FrameData_O[23]
port 50 nsew signal output
flabel metal2 s 46278 8612 46368 8692 0 FreeSans 320 0 0 0 FrameData_O[24]
port 51 nsew signal output
flabel metal2 s 46278 8948 46368 9028 0 FreeSans 320 0 0 0 FrameData_O[25]
port 52 nsew signal output
flabel metal2 s 46278 9284 46368 9364 0 FreeSans 320 0 0 0 FrameData_O[26]
port 53 nsew signal output
flabel metal2 s 46278 9620 46368 9700 0 FreeSans 320 0 0 0 FrameData_O[27]
port 54 nsew signal output
flabel metal2 s 46278 9956 46368 10036 0 FreeSans 320 0 0 0 FrameData_O[28]
port 55 nsew signal output
flabel metal2 s 46278 10292 46368 10372 0 FreeSans 320 0 0 0 FrameData_O[29]
port 56 nsew signal output
flabel metal2 s 46278 1220 46368 1300 0 FreeSans 320 0 0 0 FrameData_O[2]
port 57 nsew signal output
flabel metal2 s 46278 10628 46368 10708 0 FreeSans 320 0 0 0 FrameData_O[30]
port 58 nsew signal output
flabel metal2 s 46278 10964 46368 11044 0 FreeSans 320 0 0 0 FrameData_O[31]
port 59 nsew signal output
flabel metal2 s 46278 1556 46368 1636 0 FreeSans 320 0 0 0 FrameData_O[3]
port 60 nsew signal output
flabel metal2 s 46278 1892 46368 1972 0 FreeSans 320 0 0 0 FrameData_O[4]
port 61 nsew signal output
flabel metal2 s 46278 2228 46368 2308 0 FreeSans 320 0 0 0 FrameData_O[5]
port 62 nsew signal output
flabel metal2 s 46278 2564 46368 2644 0 FreeSans 320 0 0 0 FrameData_O[6]
port 63 nsew signal output
flabel metal2 s 46278 2900 46368 2980 0 FreeSans 320 0 0 0 FrameData_O[7]
port 64 nsew signal output
flabel metal2 s 46278 3236 46368 3316 0 FreeSans 320 0 0 0 FrameData_O[8]
port 65 nsew signal output
flabel metal2 s 46278 3572 46368 3652 0 FreeSans 320 0 0 0 FrameData_O[9]
port 66 nsew signal output
flabel metal3 s 14648 0 14728 80 0 FreeSans 320 0 0 0 FrameStrobe[0]
port 67 nsew signal input
flabel metal3 s 30008 0 30088 80 0 FreeSans 320 0 0 0 FrameStrobe[10]
port 68 nsew signal input
flabel metal3 s 31544 0 31624 80 0 FreeSans 320 0 0 0 FrameStrobe[11]
port 69 nsew signal input
flabel metal3 s 33080 0 33160 80 0 FreeSans 320 0 0 0 FrameStrobe[12]
port 70 nsew signal input
flabel metal3 s 34616 0 34696 80 0 FreeSans 320 0 0 0 FrameStrobe[13]
port 71 nsew signal input
flabel metal3 s 36152 0 36232 80 0 FreeSans 320 0 0 0 FrameStrobe[14]
port 72 nsew signal input
flabel metal3 s 37688 0 37768 80 0 FreeSans 320 0 0 0 FrameStrobe[15]
port 73 nsew signal input
flabel metal3 s 39224 0 39304 80 0 FreeSans 320 0 0 0 FrameStrobe[16]
port 74 nsew signal input
flabel metal3 s 40760 0 40840 80 0 FreeSans 320 0 0 0 FrameStrobe[17]
port 75 nsew signal input
flabel metal3 s 42296 0 42376 80 0 FreeSans 320 0 0 0 FrameStrobe[18]
port 76 nsew signal input
flabel metal3 s 43832 0 43912 80 0 FreeSans 320 0 0 0 FrameStrobe[19]
port 77 nsew signal input
flabel metal3 s 16184 0 16264 80 0 FreeSans 320 0 0 0 FrameStrobe[1]
port 78 nsew signal input
flabel metal3 s 17720 0 17800 80 0 FreeSans 320 0 0 0 FrameStrobe[2]
port 79 nsew signal input
flabel metal3 s 19256 0 19336 80 0 FreeSans 320 0 0 0 FrameStrobe[3]
port 80 nsew signal input
flabel metal3 s 20792 0 20872 80 0 FreeSans 320 0 0 0 FrameStrobe[4]
port 81 nsew signal input
flabel metal3 s 22328 0 22408 80 0 FreeSans 320 0 0 0 FrameStrobe[5]
port 82 nsew signal input
flabel metal3 s 23864 0 23944 80 0 FreeSans 320 0 0 0 FrameStrobe[6]
port 83 nsew signal input
flabel metal3 s 25400 0 25480 80 0 FreeSans 320 0 0 0 FrameStrobe[7]
port 84 nsew signal input
flabel metal3 s 26936 0 27016 80 0 FreeSans 320 0 0 0 FrameStrobe[8]
port 85 nsew signal input
flabel metal3 s 28472 0 28552 80 0 FreeSans 320 0 0 0 FrameStrobe[9]
port 86 nsew signal input
flabel metal3 s 31352 11764 31432 11844 0 FreeSans 320 0 0 0 FrameStrobe_O[0]
port 87 nsew signal output
flabel metal3 s 33272 11764 33352 11844 0 FreeSans 320 0 0 0 FrameStrobe_O[10]
port 88 nsew signal output
flabel metal3 s 33464 11764 33544 11844 0 FreeSans 320 0 0 0 FrameStrobe_O[11]
port 89 nsew signal output
flabel metal3 s 33656 11764 33736 11844 0 FreeSans 320 0 0 0 FrameStrobe_O[12]
port 90 nsew signal output
flabel metal3 s 33848 11764 33928 11844 0 FreeSans 320 0 0 0 FrameStrobe_O[13]
port 91 nsew signal output
flabel metal3 s 34040 11764 34120 11844 0 FreeSans 320 0 0 0 FrameStrobe_O[14]
port 92 nsew signal output
flabel metal3 s 34232 11764 34312 11844 0 FreeSans 320 0 0 0 FrameStrobe_O[15]
port 93 nsew signal output
flabel metal3 s 34424 11764 34504 11844 0 FreeSans 320 0 0 0 FrameStrobe_O[16]
port 94 nsew signal output
flabel metal3 s 34616 11764 34696 11844 0 FreeSans 320 0 0 0 FrameStrobe_O[17]
port 95 nsew signal output
flabel metal3 s 34808 11764 34888 11844 0 FreeSans 320 0 0 0 FrameStrobe_O[18]
port 96 nsew signal output
flabel metal3 s 35000 11764 35080 11844 0 FreeSans 320 0 0 0 FrameStrobe_O[19]
port 97 nsew signal output
flabel metal3 s 31544 11764 31624 11844 0 FreeSans 320 0 0 0 FrameStrobe_O[1]
port 98 nsew signal output
flabel metal3 s 31736 11764 31816 11844 0 FreeSans 320 0 0 0 FrameStrobe_O[2]
port 99 nsew signal output
flabel metal3 s 31928 11764 32008 11844 0 FreeSans 320 0 0 0 FrameStrobe_O[3]
port 100 nsew signal output
flabel metal3 s 32120 11764 32200 11844 0 FreeSans 320 0 0 0 FrameStrobe_O[4]
port 101 nsew signal output
flabel metal3 s 32312 11764 32392 11844 0 FreeSans 320 0 0 0 FrameStrobe_O[5]
port 102 nsew signal output
flabel metal3 s 32504 11764 32584 11844 0 FreeSans 320 0 0 0 FrameStrobe_O[6]
port 103 nsew signal output
flabel metal3 s 32696 11764 32776 11844 0 FreeSans 320 0 0 0 FrameStrobe_O[7]
port 104 nsew signal output
flabel metal3 s 32888 11764 32968 11844 0 FreeSans 320 0 0 0 FrameStrobe_O[8]
port 105 nsew signal output
flabel metal3 s 33080 11764 33160 11844 0 FreeSans 320 0 0 0 FrameStrobe_O[9]
port 106 nsew signal output
flabel metal3 s 11000 11764 11080 11844 0 FreeSans 320 0 0 0 N1BEG[0]
port 107 nsew signal output
flabel metal3 s 11192 11764 11272 11844 0 FreeSans 320 0 0 0 N1BEG[1]
port 108 nsew signal output
flabel metal3 s 11384 11764 11464 11844 0 FreeSans 320 0 0 0 N1BEG[2]
port 109 nsew signal output
flabel metal3 s 11576 11764 11656 11844 0 FreeSans 320 0 0 0 N1BEG[3]
port 110 nsew signal output
flabel metal3 s 11768 11764 11848 11844 0 FreeSans 320 0 0 0 N2BEG[0]
port 111 nsew signal output
flabel metal3 s 11960 11764 12040 11844 0 FreeSans 320 0 0 0 N2BEG[1]
port 112 nsew signal output
flabel metal3 s 12152 11764 12232 11844 0 FreeSans 320 0 0 0 N2BEG[2]
port 113 nsew signal output
flabel metal3 s 12344 11764 12424 11844 0 FreeSans 320 0 0 0 N2BEG[3]
port 114 nsew signal output
flabel metal3 s 12536 11764 12616 11844 0 FreeSans 320 0 0 0 N2BEG[4]
port 115 nsew signal output
flabel metal3 s 12728 11764 12808 11844 0 FreeSans 320 0 0 0 N2BEG[5]
port 116 nsew signal output
flabel metal3 s 12920 11764 13000 11844 0 FreeSans 320 0 0 0 N2BEG[6]
port 117 nsew signal output
flabel metal3 s 13112 11764 13192 11844 0 FreeSans 320 0 0 0 N2BEG[7]
port 118 nsew signal output
flabel metal3 s 13304 11764 13384 11844 0 FreeSans 320 0 0 0 N2BEGb[0]
port 119 nsew signal output
flabel metal3 s 13496 11764 13576 11844 0 FreeSans 320 0 0 0 N2BEGb[1]
port 120 nsew signal output
flabel metal3 s 13688 11764 13768 11844 0 FreeSans 320 0 0 0 N2BEGb[2]
port 121 nsew signal output
flabel metal3 s 13880 11764 13960 11844 0 FreeSans 320 0 0 0 N2BEGb[3]
port 122 nsew signal output
flabel metal3 s 14072 11764 14152 11844 0 FreeSans 320 0 0 0 N2BEGb[4]
port 123 nsew signal output
flabel metal3 s 14264 11764 14344 11844 0 FreeSans 320 0 0 0 N2BEGb[5]
port 124 nsew signal output
flabel metal3 s 14456 11764 14536 11844 0 FreeSans 320 0 0 0 N2BEGb[6]
port 125 nsew signal output
flabel metal3 s 14648 11764 14728 11844 0 FreeSans 320 0 0 0 N2BEGb[7]
port 126 nsew signal output
flabel metal3 s 14840 11764 14920 11844 0 FreeSans 320 0 0 0 N4BEG[0]
port 127 nsew signal output
flabel metal3 s 16760 11764 16840 11844 0 FreeSans 320 0 0 0 N4BEG[10]
port 128 nsew signal output
flabel metal3 s 16952 11764 17032 11844 0 FreeSans 320 0 0 0 N4BEG[11]
port 129 nsew signal output
flabel metal3 s 17144 11764 17224 11844 0 FreeSans 320 0 0 0 N4BEG[12]
port 130 nsew signal output
flabel metal3 s 17336 11764 17416 11844 0 FreeSans 320 0 0 0 N4BEG[13]
port 131 nsew signal output
flabel metal3 s 17528 11764 17608 11844 0 FreeSans 320 0 0 0 N4BEG[14]
port 132 nsew signal output
flabel metal3 s 17720 11764 17800 11844 0 FreeSans 320 0 0 0 N4BEG[15]
port 133 nsew signal output
flabel metal3 s 15032 11764 15112 11844 0 FreeSans 320 0 0 0 N4BEG[1]
port 134 nsew signal output
flabel metal3 s 15224 11764 15304 11844 0 FreeSans 320 0 0 0 N4BEG[2]
port 135 nsew signal output
flabel metal3 s 15416 11764 15496 11844 0 FreeSans 320 0 0 0 N4BEG[3]
port 136 nsew signal output
flabel metal3 s 15608 11764 15688 11844 0 FreeSans 320 0 0 0 N4BEG[4]
port 137 nsew signal output
flabel metal3 s 15800 11764 15880 11844 0 FreeSans 320 0 0 0 N4BEG[5]
port 138 nsew signal output
flabel metal3 s 15992 11764 16072 11844 0 FreeSans 320 0 0 0 N4BEG[6]
port 139 nsew signal output
flabel metal3 s 16184 11764 16264 11844 0 FreeSans 320 0 0 0 N4BEG[7]
port 140 nsew signal output
flabel metal3 s 16376 11764 16456 11844 0 FreeSans 320 0 0 0 N4BEG[8]
port 141 nsew signal output
flabel metal3 s 16568 11764 16648 11844 0 FreeSans 320 0 0 0 N4BEG[9]
port 142 nsew signal output
flabel metal3 s 17912 11764 17992 11844 0 FreeSans 320 0 0 0 NN4BEG[0]
port 143 nsew signal output
flabel metal3 s 19832 11764 19912 11844 0 FreeSans 320 0 0 0 NN4BEG[10]
port 144 nsew signal output
flabel metal3 s 20024 11764 20104 11844 0 FreeSans 320 0 0 0 NN4BEG[11]
port 145 nsew signal output
flabel metal3 s 20216 11764 20296 11844 0 FreeSans 320 0 0 0 NN4BEG[12]
port 146 nsew signal output
flabel metal3 s 20408 11764 20488 11844 0 FreeSans 320 0 0 0 NN4BEG[13]
port 147 nsew signal output
flabel metal3 s 20600 11764 20680 11844 0 FreeSans 320 0 0 0 NN4BEG[14]
port 148 nsew signal output
flabel metal3 s 20792 11764 20872 11844 0 FreeSans 320 0 0 0 NN4BEG[15]
port 149 nsew signal output
flabel metal3 s 18104 11764 18184 11844 0 FreeSans 320 0 0 0 NN4BEG[1]
port 150 nsew signal output
flabel metal3 s 18296 11764 18376 11844 0 FreeSans 320 0 0 0 NN4BEG[2]
port 151 nsew signal output
flabel metal3 s 18488 11764 18568 11844 0 FreeSans 320 0 0 0 NN4BEG[3]
port 152 nsew signal output
flabel metal3 s 18680 11764 18760 11844 0 FreeSans 320 0 0 0 NN4BEG[4]
port 153 nsew signal output
flabel metal3 s 18872 11764 18952 11844 0 FreeSans 320 0 0 0 NN4BEG[5]
port 154 nsew signal output
flabel metal3 s 19064 11764 19144 11844 0 FreeSans 320 0 0 0 NN4BEG[6]
port 155 nsew signal output
flabel metal3 s 19256 11764 19336 11844 0 FreeSans 320 0 0 0 NN4BEG[7]
port 156 nsew signal output
flabel metal3 s 19448 11764 19528 11844 0 FreeSans 320 0 0 0 NN4BEG[8]
port 157 nsew signal output
flabel metal3 s 19640 11764 19720 11844 0 FreeSans 320 0 0 0 NN4BEG[9]
port 158 nsew signal output
flabel metal3 s 3896 0 3976 80 0 FreeSans 320 0 0 0 RESET_top
port 159 nsew signal input
flabel metal3 s 21176 11764 21256 11844 0 FreeSans 320 0 0 0 S1END[0]
port 160 nsew signal input
flabel metal3 s 21368 11764 21448 11844 0 FreeSans 320 0 0 0 S1END[1]
port 161 nsew signal input
flabel metal3 s 21560 11764 21640 11844 0 FreeSans 320 0 0 0 S1END[2]
port 162 nsew signal input
flabel metal3 s 21752 11764 21832 11844 0 FreeSans 320 0 0 0 S1END[3]
port 163 nsew signal input
flabel metal3 s 23480 11764 23560 11844 0 FreeSans 320 0 0 0 S2END[0]
port 164 nsew signal input
flabel metal3 s 23672 11764 23752 11844 0 FreeSans 320 0 0 0 S2END[1]
port 165 nsew signal input
flabel metal3 s 23864 11764 23944 11844 0 FreeSans 320 0 0 0 S2END[2]
port 166 nsew signal input
flabel metal3 s 24056 11764 24136 11844 0 FreeSans 320 0 0 0 S2END[3]
port 167 nsew signal input
flabel metal3 s 24248 11764 24328 11844 0 FreeSans 320 0 0 0 S2END[4]
port 168 nsew signal input
flabel metal3 s 24440 11764 24520 11844 0 FreeSans 320 0 0 0 S2END[5]
port 169 nsew signal input
flabel metal3 s 24632 11764 24712 11844 0 FreeSans 320 0 0 0 S2END[6]
port 170 nsew signal input
flabel metal3 s 24824 11764 24904 11844 0 FreeSans 320 0 0 0 S2END[7]
port 171 nsew signal input
flabel metal3 s 21944 11764 22024 11844 0 FreeSans 320 0 0 0 S2MID[0]
port 172 nsew signal input
flabel metal3 s 22136 11764 22216 11844 0 FreeSans 320 0 0 0 S2MID[1]
port 173 nsew signal input
flabel metal3 s 22328 11764 22408 11844 0 FreeSans 320 0 0 0 S2MID[2]
port 174 nsew signal input
flabel metal3 s 22520 11764 22600 11844 0 FreeSans 320 0 0 0 S2MID[3]
port 175 nsew signal input
flabel metal3 s 22712 11764 22792 11844 0 FreeSans 320 0 0 0 S2MID[4]
port 176 nsew signal input
flabel metal3 s 22904 11764 22984 11844 0 FreeSans 320 0 0 0 S2MID[5]
port 177 nsew signal input
flabel metal3 s 23096 11764 23176 11844 0 FreeSans 320 0 0 0 S2MID[6]
port 178 nsew signal input
flabel metal3 s 23288 11764 23368 11844 0 FreeSans 320 0 0 0 S2MID[7]
port 179 nsew signal input
flabel metal3 s 25016 11764 25096 11844 0 FreeSans 320 0 0 0 S4END[0]
port 180 nsew signal input
flabel metal3 s 26936 11764 27016 11844 0 FreeSans 320 0 0 0 S4END[10]
port 181 nsew signal input
flabel metal3 s 27128 11764 27208 11844 0 FreeSans 320 0 0 0 S4END[11]
port 182 nsew signal input
flabel metal3 s 27320 11764 27400 11844 0 FreeSans 320 0 0 0 S4END[12]
port 183 nsew signal input
flabel metal3 s 27512 11764 27592 11844 0 FreeSans 320 0 0 0 S4END[13]
port 184 nsew signal input
flabel metal3 s 27704 11764 27784 11844 0 FreeSans 320 0 0 0 S4END[14]
port 185 nsew signal input
flabel metal3 s 27896 11764 27976 11844 0 FreeSans 320 0 0 0 S4END[15]
port 186 nsew signal input
flabel metal3 s 25208 11764 25288 11844 0 FreeSans 320 0 0 0 S4END[1]
port 187 nsew signal input
flabel metal3 s 25400 11764 25480 11844 0 FreeSans 320 0 0 0 S4END[2]
port 188 nsew signal input
flabel metal3 s 25592 11764 25672 11844 0 FreeSans 320 0 0 0 S4END[3]
port 189 nsew signal input
flabel metal3 s 25784 11764 25864 11844 0 FreeSans 320 0 0 0 S4END[4]
port 190 nsew signal input
flabel metal3 s 25976 11764 26056 11844 0 FreeSans 320 0 0 0 S4END[5]
port 191 nsew signal input
flabel metal3 s 26168 11764 26248 11844 0 FreeSans 320 0 0 0 S4END[6]
port 192 nsew signal input
flabel metal3 s 26360 11764 26440 11844 0 FreeSans 320 0 0 0 S4END[7]
port 193 nsew signal input
flabel metal3 s 26552 11764 26632 11844 0 FreeSans 320 0 0 0 S4END[8]
port 194 nsew signal input
flabel metal3 s 26744 11764 26824 11844 0 FreeSans 320 0 0 0 S4END[9]
port 195 nsew signal input
flabel metal3 s 6968 0 7048 80 0 FreeSans 320 0 0 0 SLOT_top0
port 196 nsew signal output
flabel metal3 s 8504 0 8584 80 0 FreeSans 320 0 0 0 SLOT_top1
port 197 nsew signal output
flabel metal3 s 10040 0 10120 80 0 FreeSans 320 0 0 0 SLOT_top2
port 198 nsew signal output
flabel metal3 s 11576 0 11656 80 0 FreeSans 320 0 0 0 SLOT_top3
port 199 nsew signal output
flabel metal3 s 28088 11764 28168 11844 0 FreeSans 320 0 0 0 SS4END[0]
port 200 nsew signal input
flabel metal3 s 30008 11764 30088 11844 0 FreeSans 320 0 0 0 SS4END[10]
port 201 nsew signal input
flabel metal3 s 30200 11764 30280 11844 0 FreeSans 320 0 0 0 SS4END[11]
port 202 nsew signal input
flabel metal3 s 30392 11764 30472 11844 0 FreeSans 320 0 0 0 SS4END[12]
port 203 nsew signal input
flabel metal3 s 30584 11764 30664 11844 0 FreeSans 320 0 0 0 SS4END[13]
port 204 nsew signal input
flabel metal3 s 30776 11764 30856 11844 0 FreeSans 320 0 0 0 SS4END[14]
port 205 nsew signal input
flabel metal3 s 30968 11764 31048 11844 0 FreeSans 320 0 0 0 SS4END[15]
port 206 nsew signal input
flabel metal3 s 28280 11764 28360 11844 0 FreeSans 320 0 0 0 SS4END[1]
port 207 nsew signal input
flabel metal3 s 28472 11764 28552 11844 0 FreeSans 320 0 0 0 SS4END[2]
port 208 nsew signal input
flabel metal3 s 28664 11764 28744 11844 0 FreeSans 320 0 0 0 SS4END[3]
port 209 nsew signal input
flabel metal3 s 28856 11764 28936 11844 0 FreeSans 320 0 0 0 SS4END[4]
port 210 nsew signal input
flabel metal3 s 29048 11764 29128 11844 0 FreeSans 320 0 0 0 SS4END[5]
port 211 nsew signal input
flabel metal3 s 29240 11764 29320 11844 0 FreeSans 320 0 0 0 SS4END[6]
port 212 nsew signal input
flabel metal3 s 29432 11764 29512 11844 0 FreeSans 320 0 0 0 SS4END[7]
port 213 nsew signal input
flabel metal3 s 29624 11764 29704 11844 0 FreeSans 320 0 0 0 SS4END[8]
port 214 nsew signal input
flabel metal3 s 29816 11764 29896 11844 0 FreeSans 320 0 0 0 SS4END[9]
port 215 nsew signal input
flabel metal3 s 13112 0 13192 80 0 FreeSans 320 0 0 0 UserCLK
port 216 nsew signal input
flabel metal3 s 31160 11764 31240 11844 0 FreeSans 320 0 0 0 UserCLKo
port 217 nsew signal output
flabel metal5 s 4892 0 5332 11844 0 FreeSans 2560 90 0 0 VGND
port 218 nsew ground bidirectional
flabel metal5 s 4892 0 5332 40 0 FreeSans 320 0 0 0 VGND
port 218 nsew ground bidirectional
flabel metal5 s 4892 11804 5332 11844 0 FreeSans 320 0 0 0 VGND
port 218 nsew ground bidirectional
flabel metal5 s 20012 0 20452 11844 0 FreeSans 2560 90 0 0 VGND
port 218 nsew ground bidirectional
flabel metal5 s 20012 0 20452 40 0 FreeSans 320 0 0 0 VGND
port 218 nsew ground bidirectional
flabel metal5 s 20012 11804 20452 11844 0 FreeSans 320 0 0 0 VGND
port 218 nsew ground bidirectional
flabel metal5 s 35132 0 35572 11844 0 FreeSans 2560 90 0 0 VGND
port 218 nsew ground bidirectional
flabel metal5 s 35132 0 35572 40 0 FreeSans 320 0 0 0 VGND
port 218 nsew ground bidirectional
flabel metal5 s 35132 11804 35572 11844 0 FreeSans 320 0 0 0 VGND
port 218 nsew ground bidirectional
flabel metal5 s 3652 0 4092 11844 0 FreeSans 2560 90 0 0 VPWR
port 219 nsew power bidirectional
flabel metal5 s 3652 0 4092 40 0 FreeSans 320 0 0 0 VPWR
port 219 nsew power bidirectional
flabel metal5 s 3652 11804 4092 11844 0 FreeSans 320 0 0 0 VPWR
port 219 nsew power bidirectional
flabel metal5 s 18772 0 19212 11844 0 FreeSans 2560 90 0 0 VPWR
port 219 nsew power bidirectional
flabel metal5 s 18772 0 19212 40 0 FreeSans 320 0 0 0 VPWR
port 219 nsew power bidirectional
flabel metal5 s 18772 11804 19212 11844 0 FreeSans 320 0 0 0 VPWR
port 219 nsew power bidirectional
flabel metal5 s 33892 0 34332 11844 0 FreeSans 2560 90 0 0 VPWR
port 219 nsew power bidirectional
flabel metal5 s 33892 0 34332 40 0 FreeSans 320 0 0 0 VPWR
port 219 nsew power bidirectional
flabel metal5 s 33892 11804 34332 11844 0 FreeSans 320 0 0 0 VPWR
port 219 nsew power bidirectional
rlabel metal1 23184 9072 23184 9072 0 VGND
rlabel metal1 23184 9828 23184 9828 0 VPWR
rlabel metal3 5472 870 5472 870 0 BOOT_top
rlabel metal3 2400 996 2400 996 0 CONFIGURED_top
rlabel metal3 39456 1134 39456 1134 0 FrameData[0]
rlabel metal3 19488 2940 19488 2940 0 FrameData[10]
rlabel metal2 19392 4242 19392 4242 0 FrameData[11]
rlabel metal2 33840 7980 33840 7980 0 FrameData[12]
rlabel metal2 1040 4956 1040 4956 0 FrameData[13]
rlabel metal2 464 5292 464 5292 0 FrameData[14]
rlabel metal2 656 5628 656 5628 0 FrameData[15]
rlabel metal2 848 5964 848 5964 0 FrameData[16]
rlabel metal2 656 6300 656 6300 0 FrameData[17]
rlabel metal2 704 6636 704 6636 0 FrameData[18]
rlabel metal2 656 6972 656 6972 0 FrameData[19]
rlabel metal2 39648 3444 39648 3444 0 FrameData[1]
rlabel metal2 656 7308 656 7308 0 FrameData[20]
rlabel metal2 464 7644 464 7644 0 FrameData[21]
rlabel metal2 368 7980 368 7980 0 FrameData[22]
rlabel metal2 848 8316 848 8316 0 FrameData[23]
rlabel metal2 320 8652 320 8652 0 FrameData[24]
rlabel metal2 656 8988 656 8988 0 FrameData[25]
rlabel metal2 848 9324 848 9324 0 FrameData[26]
rlabel metal2 1040 9660 1040 9660 0 FrameData[27]
rlabel metal2 512 9996 512 9996 0 FrameData[28]
rlabel metal2 752 10332 752 10332 0 FrameData[29]
rlabel metal2 39216 3444 39216 3444 0 FrameData[2]
rlabel metal2 608 10668 608 10668 0 FrameData[30]
rlabel metal2 704 11004 704 11004 0 FrameData[31]
rlabel metal2 272 1596 272 1596 0 FrameData[3]
rlabel metal2 656 1932 656 1932 0 FrameData[4]
rlabel metal2 1808 2268 1808 2268 0 FrameData[5]
rlabel metal2 1616 2604 1616 2604 0 FrameData[6]
rlabel metal2 752 2940 752 2940 0 FrameData[7]
rlabel metal2 704 3276 704 3276 0 FrameData[8]
rlabel metal2 368 3612 368 3612 0 FrameData[9]
rlabel metal2 45471 588 45471 588 0 FrameData_O[0]
rlabel metal2 45855 3948 45855 3948 0 FrameData_O[10]
rlabel metal2 45576 3612 45576 3612 0 FrameData_O[11]
rlabel metal2 45663 4620 45663 4620 0 FrameData_O[12]
rlabel metal2 45480 4284 45480 4284 0 FrameData_O[13]
rlabel metal2 45663 5292 45663 5292 0 FrameData_O[14]
rlabel metal2 45288 5124 45288 5124 0 FrameData_O[15]
rlabel via2 46287 5964 46287 5964 0 FrameData_O[16]
rlabel metal2 45192 5628 45192 5628 0 FrameData_O[17]
rlabel metal2 45663 6636 45663 6636 0 FrameData_O[18]
rlabel metal2 45735 6972 45735 6972 0 FrameData_O[19]
rlabel metal2 45999 924 45999 924 0 FrameData_O[1]
rlabel metal2 46143 7308 46143 7308 0 FrameData_O[20]
rlabel metal2 45663 7644 45663 7644 0 FrameData_O[21]
rlabel metal2 46047 7980 46047 7980 0 FrameData_O[22]
rlabel metal2 45663 8316 45663 8316 0 FrameData_O[23]
rlabel metal2 46239 8652 46239 8652 0 FrameData_O[24]
rlabel metal2 46287 8988 46287 8988 0 FrameData_O[25]
rlabel metal2 45735 9324 45735 9324 0 FrameData_O[26]
rlabel metal2 45543 9660 45543 9660 0 FrameData_O[27]
rlabel metal2 44472 8904 44472 8904 0 FrameData_O[28]
rlabel metal2 44424 9660 44424 9660 0 FrameData_O[29]
rlabel via2 46287 1260 46287 1260 0 FrameData_O[2]
rlabel metal2 44040 9660 44040 9660 0 FrameData_O[30]
rlabel metal2 44751 11004 44751 11004 0 FrameData_O[31]
rlabel metal2 45543 1596 45543 1596 0 FrameData_O[3]
rlabel metal2 45855 1932 45855 1932 0 FrameData_O[4]
rlabel metal2 43320 2016 43320 2016 0 FrameData_O[5]
rlabel metal2 46047 2604 46047 2604 0 FrameData_O[6]
rlabel metal2 45903 2940 45903 2940 0 FrameData_O[7]
rlabel metal2 45543 3276 45543 3276 0 FrameData_O[8]
rlabel metal2 46239 3612 46239 3612 0 FrameData_O[9]
rlabel metal2 15840 8064 15840 8064 0 FrameStrobe[0]
rlabel metal2 43680 3444 43680 3444 0 FrameStrobe[10]
rlabel metal2 37824 3234 37824 3234 0 FrameStrobe[11]
rlabel metal2 43488 8610 43488 8610 0 FrameStrobe[12]
rlabel metal2 44160 8022 44160 8022 0 FrameStrobe[13]
rlabel metal3 36192 3516 36192 3516 0 FrameStrobe[14]
rlabel metal2 36000 7224 36000 7224 0 FrameStrobe[15]
rlabel metal3 39264 618 39264 618 0 FrameStrobe[16]
rlabel metal2 37872 8568 37872 8568 0 FrameStrobe[17]
rlabel metal4 34224 8064 34224 8064 0 FrameStrobe[18]
rlabel metal2 43296 7938 43296 7938 0 FrameStrobe[19]
rlabel metal3 16224 1122 16224 1122 0 FrameStrobe[1]
rlabel metal3 17760 1248 17760 1248 0 FrameStrobe[2]
rlabel metal3 19296 114 19296 114 0 FrameStrobe[3]
rlabel metal3 20832 2088 20832 2088 0 FrameStrobe[4]
rlabel metal3 22368 156 22368 156 0 FrameStrobe[5]
rlabel metal2 42048 4032 42048 4032 0 FrameStrobe[6]
rlabel metal3 25440 1470 25440 1470 0 FrameStrobe[7]
rlabel metal3 43392 3360 43392 3360 0 FrameStrobe[8]
rlabel metal2 43776 3192 43776 3192 0 FrameStrobe[9]
rlabel metal2 31512 9576 31512 9576 0 FrameStrobe_O[0]
rlabel metal2 33336 8904 33336 8904 0 FrameStrobe_O[10]
rlabel metal2 33912 9660 33912 9660 0 FrameStrobe_O[11]
rlabel metal2 33720 8904 33720 8904 0 FrameStrobe_O[12]
rlabel metal2 34728 9660 34728 9660 0 FrameStrobe_O[13]
rlabel metal2 34248 8904 34248 8904 0 FrameStrobe_O[14]
rlabel metal2 34824 9324 34824 9324 0 FrameStrobe_O[15]
rlabel metal2 34488 8820 34488 8820 0 FrameStrobe_O[16]
rlabel metal2 35448 9576 35448 9576 0 FrameStrobe_O[17]
rlabel metal2 34872 8904 34872 8904 0 FrameStrobe_O[18]
rlabel metal2 35448 9660 35448 9660 0 FrameStrobe_O[19]
rlabel metal2 31800 9660 31800 9660 0 FrameStrobe_O[1]
rlabel metal2 32088 9576 32088 9576 0 FrameStrobe_O[2]
rlabel metal2 32376 9324 32376 9324 0 FrameStrobe_O[3]
rlabel metal2 32184 8904 32184 8904 0 FrameStrobe_O[4]
rlabel metal2 33144 9324 33144 9324 0 FrameStrobe_O[5]
rlabel metal2 32568 8904 32568 8904 0 FrameStrobe_O[6]
rlabel metal3 32736 10680 32736 10680 0 FrameStrobe_O[7]
rlabel metal2 32952 8904 32952 8904 0 FrameStrobe_O[8]
rlabel metal2 33576 9240 33576 9240 0 FrameStrobe_O[9]
rlabel metal2 9648 2856 9648 2856 0 Inst_S_WARMBOOT_ConfigMem.Inst_frame0_bit13.Q
rlabel metal2 25920 4242 25920 4242 0 Inst_S_WARMBOOT_ConfigMem.Inst_frame0_bit14.Q
rlabel metal2 26016 3360 26016 3360 0 Inst_S_WARMBOOT_ConfigMem.Inst_frame0_bit15.Q
rlabel metal2 15408 3192 15408 3192 0 Inst_S_WARMBOOT_ConfigMem.Inst_frame0_bit16.Q
rlabel metal2 14736 6972 14736 6972 0 Inst_S_WARMBOOT_ConfigMem.Inst_frame0_bit17.Q
rlabel via1 12552 7392 12552 7392 0 Inst_S_WARMBOOT_ConfigMem.Inst_frame0_bit18.Q
rlabel metal2 13488 3612 13488 3612 0 Inst_S_WARMBOOT_ConfigMem.Inst_frame0_bit19.Q
rlabel metal2 17952 2688 17952 2688 0 Inst_S_WARMBOOT_ConfigMem.Inst_frame0_bit20.Q
rlabel metal2 19632 3948 19632 3948 0 Inst_S_WARMBOOT_ConfigMem.Inst_frame0_bit21.Q
rlabel metal3 21792 3528 21792 3528 0 Inst_S_WARMBOOT_ConfigMem.Inst_frame0_bit22.Q
rlabel metal2 30720 3402 30720 3402 0 Inst_S_WARMBOOT_ConfigMem.Inst_frame0_bit23.Q
rlabel metal2 33024 4242 33024 4242 0 Inst_S_WARMBOOT_ConfigMem.Inst_frame0_bit24.Q
rlabel metal3 34368 4410 34368 4410 0 Inst_S_WARMBOOT_ConfigMem.Inst_frame0_bit25.Q
rlabel metal2 26256 7224 26256 7224 0 Inst_S_WARMBOOT_ConfigMem.Inst_frame0_bit26.Q
rlabel metal2 28512 7224 28512 7224 0 Inst_S_WARMBOOT_ConfigMem.Inst_frame0_bit27.Q
rlabel metal2 25392 8064 25392 8064 0 Inst_S_WARMBOOT_ConfigMem.Inst_frame0_bit28.Q
rlabel metal2 9408 5754 9408 5754 0 Inst_S_WARMBOOT_ConfigMem.Inst_frame0_bit29.Q
rlabel metal3 10944 6804 10944 6804 0 Inst_S_WARMBOOT_ConfigMem.Inst_frame0_bit30.Q
rlabel metal2 11232 2856 11232 2856 0 Inst_S_WARMBOOT_ConfigMem.Inst_frame0_bit31.Q
rlabel metal2 9408 3696 9408 3696 0 Inst_S_WARMBOOT_switch_matrix.N1BEG0
rlabel metal2 27168 4116 27168 4116 0 Inst_S_WARMBOOT_switch_matrix.N1BEG1
rlabel metal2 27264 3486 27264 3486 0 Inst_S_WARMBOOT_switch_matrix.N1BEG2
rlabel metal2 16128 3444 16128 3444 0 Inst_S_WARMBOOT_switch_matrix.N1BEG3
rlabel metal2 10872 8904 10872 8904 0 N1BEG[0]
rlabel metal2 10728 9660 10728 9660 0 N1BEG[1]
rlabel metal2 11016 9576 11016 9576 0 N1BEG[2]
rlabel metal2 11544 8904 11544 8904 0 N1BEG[3]
rlabel metal2 11400 9324 11400 9324 0 N2BEG[0]
rlabel metal2 11688 9660 11688 9660 0 N2BEG[1]
rlabel metal2 12216 8904 12216 8904 0 N2BEG[2]
rlabel metal2 12072 9576 12072 9576 0 N2BEG[3]
rlabel metal2 12600 8904 12600 8904 0 N2BEG[4]
rlabel metal2 12456 9660 12456 9660 0 N2BEG[5]
rlabel metal2 13032 8904 13032 8904 0 N2BEG[6]
rlabel metal3 13152 10680 13152 10680 0 N2BEG[7]
rlabel metal2 13368 8904 13368 8904 0 N2BEGb[0]
rlabel metal3 13536 10680 13536 10680 0 N2BEGb[1]
rlabel metal2 13752 8904 13752 8904 0 N2BEGb[2]
rlabel metal2 13608 9660 13608 9660 0 N2BEGb[3]
rlabel metal2 14040 8484 14040 8484 0 N2BEGb[4]
rlabel metal2 13992 9576 13992 9576 0 N2BEGb[5]
rlabel metal2 14520 8904 14520 8904 0 N2BEGb[6]
rlabel metal2 14376 9660 14376 9660 0 N2BEGb[7]
rlabel metal2 14664 9576 14664 9576 0 N4BEG[0]
rlabel metal2 16824 8904 16824 8904 0 N4BEG[10]
rlabel metal2 16872 9660 16872 9660 0 N4BEG[11]
rlabel metal2 17208 8904 17208 8904 0 N4BEG[12]
rlabel metal2 17256 9660 17256 9660 0 N4BEG[13]
rlabel metal2 17592 8904 17592 8904 0 N4BEG[14]
rlabel metal2 17640 9660 17640 9660 0 N4BEG[15]
rlabel metal2 14952 9660 14952 9660 0 N4BEG[1]
rlabel metal2 15288 8904 15288 8904 0 N4BEG[2]
rlabel metal2 15336 9660 15336 9660 0 N4BEG[3]
rlabel metal2 15672 8904 15672 8904 0 N4BEG[4]
rlabel metal2 15720 9660 15720 9660 0 N4BEG[5]
rlabel metal2 16056 8904 16056 8904 0 N4BEG[6]
rlabel metal2 16104 9660 16104 9660 0 N4BEG[7]
rlabel metal2 16440 8904 16440 8904 0 N4BEG[8]
rlabel metal2 16488 9660 16488 9660 0 N4BEG[9]
rlabel metal2 17976 8904 17976 8904 0 NN4BEG[0]
rlabel metal2 19944 8652 19944 8652 0 NN4BEG[10]
rlabel metal2 19800 9660 19800 9660 0 NN4BEG[11]
rlabel metal2 20424 8904 20424 8904 0 NN4BEG[12]
rlabel metal2 20328 9660 20328 9660 0 NN4BEG[13]
rlabel metal2 20664 8820 20664 8820 0 NN4BEG[14]
rlabel metal2 20712 9660 20712 9660 0 NN4BEG[15]
rlabel metal2 18024 9660 18024 9660 0 NN4BEG[1]
rlabel metal2 18360 8904 18360 8904 0 NN4BEG[2]
rlabel metal2 18408 9660 18408 9660 0 NN4BEG[3]
rlabel metal2 18744 8904 18744 8904 0 NN4BEG[4]
rlabel metal2 18648 9660 18648 9660 0 NN4BEG[5]
rlabel metal2 19224 8904 19224 8904 0 NN4BEG[6]
rlabel metal3 19344 10332 19344 10332 0 NN4BEG[7]
rlabel metal2 19512 8904 19512 8904 0 NN4BEG[8]
rlabel metal2 19416 9324 19416 9324 0 NN4BEG[9]
rlabel metal3 3936 996 3936 996 0 RESET_top
rlabel metal3 21216 10680 21216 10680 0 S1END[0]
rlabel metal3 21408 10218 21408 10218 0 S1END[1]
rlabel metal3 21600 10680 21600 10680 0 S1END[2]
rlabel metal3 21792 10218 21792 10218 0 S1END[3]
rlabel metal3 23520 10218 23520 10218 0 S2END[0]
rlabel metal3 23712 10680 23712 10680 0 S2END[1]
rlabel metal3 23904 10638 23904 10638 0 S2END[2]
rlabel metal3 24096 10638 24096 10638 0 S2END[3]
rlabel metal3 24288 10680 24288 10680 0 S2END[4]
rlabel metal3 24480 10680 24480 10680 0 S2END[5]
rlabel metal3 24672 10722 24672 10722 0 S2END[6]
rlabel metal3 24864 10596 24864 10596 0 S2END[7]
rlabel metal3 21984 10680 21984 10680 0 S2MID[0]
rlabel metal3 22176 10680 22176 10680 0 S2MID[1]
rlabel metal3 22368 10638 22368 10638 0 S2MID[2]
rlabel metal3 22560 10638 22560 10638 0 S2MID[3]
rlabel metal3 22752 10848 22752 10848 0 S2MID[4]
rlabel metal3 22944 10890 22944 10890 0 S2MID[5]
rlabel metal3 4032 7686 4032 7686 0 S2MID[6]
rlabel metal3 4320 9912 4320 9912 0 S2MID[7]
rlabel metal3 25056 10932 25056 10932 0 S4END[0]
rlabel metal2 2928 7980 2928 7980 0 S4END[10]
rlabel metal2 43776 7728 43776 7728 0 S4END[11]
rlabel metal3 43008 8820 43008 8820 0 S4END[12]
rlabel metal2 42240 7938 42240 7938 0 S4END[13]
rlabel metal2 43392 7896 43392 7896 0 S4END[14]
rlabel metal2 33216 7602 33216 7602 0 S4END[15]
rlabel metal3 25248 10218 25248 10218 0 S4END[1]
rlabel metal3 25440 10680 25440 10680 0 S4END[2]
rlabel metal3 25632 10218 25632 10218 0 S4END[3]
rlabel metal3 25824 10596 25824 10596 0 S4END[4]
rlabel metal3 26016 10260 26016 10260 0 S4END[5]
rlabel metal3 26208 10722 26208 10722 0 S4END[6]
rlabel metal3 26400 10764 26400 10764 0 S4END[7]
rlabel metal2 21984 8526 21984 8526 0 S4END[8]
rlabel metal3 2496 9870 2496 9870 0 S4END[9]
rlabel metal3 7008 870 7008 870 0 SLOT_top0
rlabel metal3 8544 870 8544 870 0 SLOT_top1
rlabel metal3 10080 870 10080 870 0 SLOT_top2
rlabel metal3 11616 870 11616 870 0 SLOT_top3
rlabel metal3 28128 10638 28128 10638 0 SS4END[0]
rlabel metal2 40416 8106 40416 8106 0 SS4END[10]
rlabel metal3 42048 6888 42048 6888 0 SS4END[11]
rlabel metal3 43104 6720 43104 6720 0 SS4END[12]
rlabel metal3 43488 6720 43488 6720 0 SS4END[13]
rlabel metal3 42144 6888 42144 6888 0 SS4END[14]
rlabel metal3 38064 6384 38064 6384 0 SS4END[15]
rlabel metal3 28320 10680 28320 10680 0 SS4END[1]
rlabel metal3 28512 10722 28512 10722 0 SS4END[2]
rlabel metal3 28704 10596 28704 10596 0 SS4END[3]
rlabel metal3 28896 10764 28896 10764 0 SS4END[4]
rlabel metal3 29088 10218 29088 10218 0 SS4END[5]
rlabel metal3 29280 10806 29280 10806 0 SS4END[6]
rlabel metal3 29472 10218 29472 10218 0 SS4END[7]
rlabel metal3 41760 10206 41760 10206 0 SS4END[8]
rlabel metal2 43392 8736 43392 8736 0 SS4END[9]
rlabel via2 13152 72 13152 72 0 UserCLK
rlabel metal2 31224 9660 31224 9660 0 UserCLKo
rlabel via1 12773 7224 12773 7224 0 _000_
rlabel via1 12282 7213 12282 7213 0 _001_
rlabel metal2 12072 6636 12072 6636 0 _002_
rlabel via1 11720 7213 11720 7213 0 _003_
rlabel metal2 11136 7056 11136 7056 0 _004_
rlabel via1 11928 8904 11928 8904 0 _005_
rlabel metal3 12432 7224 12432 7224 0 _006_
rlabel metal2 12144 7266 12144 7266 0 _007_
rlabel metal2 11808 6300 11808 6300 0 _008_
rlabel metal3 11808 6132 11808 6132 0 _009_
rlabel metal2 27888 7728 27888 7728 0 _010_
rlabel metal2 27861 8736 27861 8736 0 _011_
rlabel metal2 33744 4284 33744 4284 0 _012_
rlabel metal3 33600 3780 33600 3780 0 _013_
rlabel metal2 21408 3234 21408 3234 0 _014_
rlabel metal2 20760 2688 20760 2688 0 _015_
rlabel metal2 8640 2058 8640 2058 0 net1
rlabel metal2 7872 7056 7872 7056 0 net10
rlabel metal2 42360 8148 42360 8148 0 net100
rlabel metal3 42048 2016 42048 2016 0 net101
rlabel metal2 42264 5124 42264 5124 0 net102
rlabel metal2 43176 3948 43176 3948 0 net103
rlabel metal2 42456 4284 42456 4284 0 net104
rlabel metal2 43296 3906 43296 3906 0 net105
rlabel metal2 41400 3948 41400 3948 0 net106
rlabel metal3 40224 6888 40224 6888 0 net107
rlabel metal2 42792 3528 42792 3528 0 net108
rlabel metal3 41856 3402 41856 3402 0 net109
rlabel metal2 2184 7056 2184 7056 0 net11
rlabel metal2 9672 3612 9672 3612 0 net110
rlabel metal3 10848 7182 10848 7182 0 net111
rlabel metal3 15168 8988 15168 8988 0 net112
rlabel metal2 15672 3444 15672 3444 0 net113
rlabel metal2 4008 7728 4008 7728 0 net114
rlabel metal3 11136 8904 11136 8904 0 net115
rlabel metal2 7752 7728 7752 7728 0 net116
rlabel metal2 3528 7980 3528 7980 0 net117
rlabel metal2 10008 7056 10008 7056 0 net118
rlabel metal2 22848 10122 22848 10122 0 net119
rlabel metal2 1488 7602 1488 7602 0 net12
rlabel metal3 18672 1932 18672 1932 0 net120
rlabel metal2 17304 1680 17304 1680 0 net121
rlabel metal2 13632 8694 13632 8694 0 net122
rlabel metal2 13056 7014 13056 7014 0 net123
rlabel metal2 19968 2814 19968 2814 0 net124
rlabel metal2 18576 3150 18576 3150 0 net125
rlabel metal4 12528 6216 12528 6216 0 net126
rlabel metal2 18624 8190 18624 8190 0 net127
rlabel metal3 19872 2016 19872 2016 0 net128
rlabel metal2 16824 3528 16824 3528 0 net129
rlabel metal2 17856 4200 17856 4200 0 net13
rlabel metal3 14112 8316 14112 8316 0 net130
rlabel metal3 17376 7518 17376 7518 0 net131
rlabel metal2 19992 3948 19992 3948 0 net132
rlabel metal3 10560 8820 10560 8820 0 net133
rlabel metal3 19680 8358 19680 8358 0 net134
rlabel metal2 21888 4326 21888 4326 0 net135
rlabel metal2 17736 3612 17736 3612 0 net136
rlabel metal3 14592 8946 14592 8946 0 net137
rlabel metal3 15552 8274 15552 8274 0 net138
rlabel metal2 42744 8820 42744 8820 0 net139
rlabel metal2 22464 4200 22464 4200 0 net14
rlabel metal2 43512 7812 43512 7812 0 net140
rlabel metal3 15360 8652 15360 8652 0 net141
rlabel metal2 2784 7938 2784 7938 0 net142
rlabel metal2 17880 8148 17880 8148 0 net143
rlabel metal3 16704 8820 16704 8820 0 net144
rlabel metal2 28536 8148 28536 8148 0 net145
rlabel metal3 18240 7686 18240 7686 0 net146
rlabel metal2 21456 2856 21456 2856 0 net147
rlabel metal2 20424 2856 20424 2856 0 net148
rlabel metal2 20256 8610 20256 8610 0 net149
rlabel metal2 1848 8652 1848 8652 0 net15
rlabel metal2 26328 8652 26328 8652 0 net150
rlabel metal3 20928 6888 20928 6888 0 net151
rlabel metal2 19896 4368 19896 4368 0 net152
rlabel metal3 21792 6090 21792 6090 0 net153
rlabel metal3 18624 7266 18624 7266 0 net154
rlabel metal3 18048 8190 18048 8190 0 net155
rlabel metal3 19872 7602 19872 7602 0 net156
rlabel metal3 18432 8568 18432 8568 0 net157
rlabel metal2 22368 9366 22368 9366 0 net158
rlabel metal2 42360 8820 42360 8820 0 net159
rlabel metal2 2232 8652 2232 8652 0 net16
rlabel metal2 11448 7140 11448 7140 0 net160
rlabel metal2 22944 10038 22944 10038 0 net161
rlabel metal3 18624 2562 18624 2562 0 net162
rlabel metal2 13056 1932 13056 1932 0 net163
rlabel metal2 10368 2016 10368 2016 0 net164
rlabel metal2 12048 6552 12048 6552 0 net165
rlabel metal3 38592 6006 38592 6006 0 net166
rlabel metal3 21024 10344 21024 10344 0 net167
rlabel metal2 1608 9240 1608 9240 0 net17
rlabel metal2 1872 9198 1872 9198 0 net18
rlabel metal2 2568 9660 2568 9660 0 net19
rlabel metal2 7584 2604 7584 2604 0 net2
rlabel metal3 18528 8106 18528 8106 0 net20
rlabel metal3 6144 7896 6144 7896 0 net21
rlabel metal3 9024 6048 9024 6048 0 net22
rlabel metal2 9504 2730 9504 2730 0 net23
rlabel metal2 5736 2100 5736 2100 0 net24
rlabel metal2 18336 2730 18336 2730 0 net25
rlabel metal2 22368 8736 22368 8736 0 net26
rlabel via1 26402 7224 26402 7224 0 net27
rlabel metal3 21600 7182 21600 7182 0 net28
rlabel metal4 20400 3192 20400 3192 0 net29
rlabel metal2 2112 5418 2112 5418 0 net3
rlabel metal2 31488 2688 31488 2688 0 net30
rlabel metal2 26640 7140 26640 7140 0 net31
rlabel metal2 13056 6636 13056 6636 0 net32
rlabel metal2 19104 3444 19104 3444 0 net33
rlabel metal2 31776 2646 31776 2646 0 net34
rlabel metal2 27216 7224 27216 7224 0 net35
rlabel metal2 11376 5628 11376 5628 0 net36
rlabel metal2 20016 1932 20016 1932 0 net37
rlabel metal2 22464 9156 22464 9156 0 net38
rlabel metal3 27072 8736 27072 8736 0 net39
rlabel metal2 1728 5334 1728 5334 0 net4
rlabel metal2 17760 6720 17760 6720 0 net40
rlabel metal2 20544 2982 20544 2982 0 net41
rlabel metal3 25824 6132 25824 6132 0 net42
rlabel metal3 26496 8610 26496 8610 0 net43
rlabel metal2 9744 8652 9744 8652 0 net44
rlabel metal2 20352 4158 20352 4158 0 net45
rlabel metal2 33216 3486 33216 3486 0 net46
rlabel metal3 26880 8652 26880 8652 0 net47
rlabel metal2 10128 8652 10128 8652 0 net48
rlabel metal2 19704 4116 19704 4116 0 net49
rlabel metal2 2376 6216 2376 6216 0 net5
rlabel metal2 32400 4116 32400 4116 0 net50
rlabel metal3 26688 8904 26688 8904 0 net51
rlabel metal2 28512 8946 28512 8946 0 net52
rlabel metal2 20496 2604 20496 2604 0 net53
rlabel metal2 33600 3570 33600 3570 0 net54
rlabel metal2 28512 8694 28512 8694 0 net55
rlabel metal3 28896 7980 28896 7980 0 net56
rlabel metal2 6480 1932 6480 1932 0 net57
rlabel metal3 40608 2310 40608 2310 0 net58
rlabel metal2 44256 4074 44256 4074 0 net59
rlabel metal3 14880 6846 14880 6846 0 net6
rlabel metal2 44352 4074 44352 4074 0 net60
rlabel metal2 44544 4998 44544 4998 0 net61
rlabel metal3 43968 4536 43968 4536 0 net62
rlabel metal2 44544 5586 44544 5586 0 net63
rlabel metal2 44928 4872 44928 4872 0 net64
rlabel metal2 14088 2856 14088 2856 0 net65
rlabel metal2 44928 5670 44928 5670 0 net66
rlabel metal3 44256 6636 44256 6636 0 net67
rlabel metal3 43680 5250 43680 5250 0 net68
rlabel metal2 40872 3192 40872 3192 0 net69
rlabel metal2 8976 2688 8976 2688 0 net7
rlabel metal2 16008 3276 16008 3276 0 net70
rlabel metal3 44544 7812 44544 7812 0 net71
rlabel metal3 44928 8694 44928 8694 0 net72
rlabel metal3 43584 9156 43584 9156 0 net73
rlabel metal2 33600 3234 33600 3234 0 net74
rlabel metal3 39072 6720 39072 6720 0 net75
rlabel metal3 44928 9408 44928 9408 0 net76
rlabel metal2 44544 9408 44544 9408 0 net77
rlabel metal3 44160 9240 44160 9240 0 net78
rlabel metal2 44016 9492 44016 9492 0 net79
rlabel metal2 21696 4158 21696 4158 0 net8
rlabel metal2 40632 3276 40632 3276 0 net80
rlabel metal2 43632 9492 43632 9492 0 net81
rlabel metal2 9672 2100 9672 2100 0 net82
rlabel metal2 38664 3276 38664 3276 0 net83
rlabel metal2 41592 2520 41592 2520 0 net84
rlabel metal2 41664 1932 41664 1932 0 net85
rlabel metal2 39072 3108 39072 3108 0 net86
rlabel metal2 41952 2394 41952 2394 0 net87
rlabel metal2 37992 2436 37992 2436 0 net88
rlabel metal3 38688 7728 38688 7728 0 net89
rlabel metal2 17208 7728 17208 7728 0 net9
rlabel metal2 29352 3948 29352 3948 0 net90
rlabel metal2 43560 3612 43560 3612 0 net91
rlabel metal2 42120 3528 42120 3528 0 net92
rlabel metal2 38496 8820 38496 8820 0 net93
rlabel metal2 43584 8148 43584 8148 0 net94
rlabel metal2 34368 8736 34368 8736 0 net95
rlabel metal2 34536 8148 34536 8148 0 net96
rlabel metal2 34872 8148 34872 8148 0 net97
rlabel metal2 35304 8064 35304 8064 0 net98
rlabel metal3 33792 8316 33792 8316 0 net99
<< properties >>
string FIXED_BBOX 0 0 46368 11844
<< end >>
