magic
tech ihp-sg13g2
magscale 1 2
timestamp 1743693518
<< metal1 >>
rect 1152 46892 12576 46916
rect 1152 46852 4928 46892
rect 4968 46852 5010 46892
rect 5050 46852 5092 46892
rect 5132 46852 5174 46892
rect 5214 46852 5256 46892
rect 5296 46852 12576 46892
rect 1152 46828 12576 46852
rect 1659 46724 1701 46733
rect 1659 46684 1660 46724
rect 1700 46684 1701 46724
rect 1659 46675 1701 46684
rect 2235 46724 2277 46733
rect 2235 46684 2236 46724
rect 2276 46684 2277 46724
rect 2235 46675 2277 46684
rect 2811 46724 2853 46733
rect 2811 46684 2812 46724
rect 2852 46684 2853 46724
rect 2811 46675 2853 46684
rect 3387 46724 3429 46733
rect 3387 46684 3388 46724
rect 3428 46684 3429 46724
rect 3387 46675 3429 46684
rect 3963 46724 4005 46733
rect 3963 46684 3964 46724
rect 4004 46684 4005 46724
rect 3963 46675 4005 46684
rect 4539 46724 4581 46733
rect 4539 46684 4540 46724
rect 4580 46684 4581 46724
rect 4539 46675 4581 46684
rect 5115 46724 5157 46733
rect 5115 46684 5116 46724
rect 5156 46684 5157 46724
rect 5115 46675 5157 46684
rect 5691 46724 5733 46733
rect 5691 46684 5692 46724
rect 5732 46684 5733 46724
rect 5691 46675 5733 46684
rect 6267 46724 6309 46733
rect 6267 46684 6268 46724
rect 6308 46684 6309 46724
rect 6267 46675 6309 46684
rect 6843 46724 6885 46733
rect 6843 46684 6844 46724
rect 6884 46684 6885 46724
rect 6843 46675 6885 46684
rect 7419 46724 7461 46733
rect 7419 46684 7420 46724
rect 7460 46684 7461 46724
rect 7419 46675 7461 46684
rect 7995 46724 8037 46733
rect 7995 46684 7996 46724
rect 8036 46684 8037 46724
rect 7995 46675 8037 46684
rect 8571 46724 8613 46733
rect 8571 46684 8572 46724
rect 8612 46684 8613 46724
rect 8571 46675 8613 46684
rect 9147 46724 9189 46733
rect 9147 46684 9148 46724
rect 9188 46684 9189 46724
rect 9147 46675 9189 46684
rect 9723 46724 9765 46733
rect 9723 46684 9724 46724
rect 9764 46684 9765 46724
rect 9723 46675 9765 46684
rect 10299 46724 10341 46733
rect 10299 46684 10300 46724
rect 10340 46684 10341 46724
rect 10299 46675 10341 46684
rect 10875 46724 10917 46733
rect 10875 46684 10876 46724
rect 10916 46684 10917 46724
rect 10875 46675 10917 46684
rect 11451 46724 11493 46733
rect 11451 46684 11452 46724
rect 11492 46684 11493 46724
rect 11451 46675 11493 46684
rect 1227 46472 1269 46481
rect 1227 46432 1228 46472
rect 1268 46432 1269 46472
rect 1227 46423 1269 46432
rect 1899 46472 1941 46481
rect 1899 46432 1900 46472
rect 1940 46432 1941 46472
rect 1899 46423 1941 46432
rect 2475 46472 2517 46481
rect 2475 46432 2476 46472
rect 2516 46432 2517 46472
rect 2475 46423 2517 46432
rect 3051 46472 3093 46481
rect 3051 46432 3052 46472
rect 3092 46432 3093 46472
rect 3051 46423 3093 46432
rect 3627 46472 3669 46481
rect 3627 46432 3628 46472
rect 3668 46432 3669 46472
rect 3627 46423 3669 46432
rect 4203 46472 4245 46481
rect 4203 46432 4204 46472
rect 4244 46432 4245 46472
rect 4203 46423 4245 46432
rect 4779 46472 4821 46481
rect 4779 46432 4780 46472
rect 4820 46432 4821 46472
rect 4779 46423 4821 46432
rect 5355 46472 5397 46481
rect 5355 46432 5356 46472
rect 5396 46432 5397 46472
rect 5355 46423 5397 46432
rect 5931 46472 5973 46481
rect 5931 46432 5932 46472
rect 5972 46432 5973 46472
rect 5931 46423 5973 46432
rect 6507 46472 6549 46481
rect 6507 46432 6508 46472
rect 6548 46432 6549 46472
rect 6507 46423 6549 46432
rect 7083 46472 7125 46481
rect 7083 46432 7084 46472
rect 7124 46432 7125 46472
rect 7083 46423 7125 46432
rect 7659 46472 7701 46481
rect 7659 46432 7660 46472
rect 7700 46432 7701 46472
rect 7659 46423 7701 46432
rect 8235 46472 8277 46481
rect 8235 46432 8236 46472
rect 8276 46432 8277 46472
rect 8235 46423 8277 46432
rect 8811 46472 8853 46481
rect 8811 46432 8812 46472
rect 8852 46432 8853 46472
rect 8811 46423 8853 46432
rect 9387 46472 9429 46481
rect 9387 46432 9388 46472
rect 9428 46432 9429 46472
rect 9387 46423 9429 46432
rect 9963 46472 10005 46481
rect 9963 46432 9964 46472
rect 10004 46432 10005 46472
rect 9963 46423 10005 46432
rect 10539 46472 10581 46481
rect 10539 46432 10540 46472
rect 10580 46432 10581 46472
rect 10539 46423 10581 46432
rect 11115 46472 11157 46481
rect 11115 46432 11116 46472
rect 11156 46432 11157 46472
rect 11115 46423 11157 46432
rect 11691 46472 11733 46481
rect 11691 46432 11692 46472
rect 11732 46432 11733 46472
rect 11691 46423 11733 46432
rect 11883 46472 11925 46481
rect 11883 46432 11884 46472
rect 11924 46432 11925 46472
rect 11883 46423 11925 46432
rect 12267 46472 12309 46481
rect 12267 46432 12268 46472
rect 12308 46432 12309 46472
rect 12267 46423 12309 46432
rect 1467 46304 1509 46313
rect 1467 46264 1468 46304
rect 1508 46264 1509 46304
rect 1467 46255 1509 46264
rect 12123 46304 12165 46313
rect 12123 46264 12124 46304
rect 12164 46264 12165 46304
rect 12123 46255 12165 46264
rect 12507 46304 12549 46313
rect 12507 46264 12508 46304
rect 12548 46264 12549 46304
rect 12507 46255 12549 46264
rect 1152 46136 12576 46160
rect 1152 46096 3688 46136
rect 3728 46096 3770 46136
rect 3810 46096 3852 46136
rect 3892 46096 3934 46136
rect 3974 46096 4016 46136
rect 4056 46096 12576 46136
rect 1152 46072 12576 46096
rect 1563 45968 1605 45977
rect 1563 45928 1564 45968
rect 1604 45928 1605 45968
rect 1563 45919 1605 45928
rect 10395 45968 10437 45977
rect 10395 45928 10396 45968
rect 10436 45928 10437 45968
rect 10395 45919 10437 45928
rect 11259 45968 11301 45977
rect 11259 45928 11260 45968
rect 11300 45928 11301 45968
rect 11259 45919 11301 45928
rect 10779 45884 10821 45893
rect 10779 45844 10780 45884
rect 10820 45844 10821 45884
rect 10779 45835 10821 45844
rect 1227 45800 1269 45809
rect 1227 45760 1228 45800
rect 1268 45760 1269 45800
rect 1227 45751 1269 45760
rect 1803 45800 1845 45809
rect 1803 45760 1804 45800
rect 1844 45760 1845 45800
rect 1803 45751 1845 45760
rect 10155 45800 10197 45809
rect 10155 45760 10156 45800
rect 10196 45760 10197 45800
rect 10155 45751 10197 45760
rect 10539 45800 10581 45809
rect 10539 45760 10540 45800
rect 10580 45760 10581 45800
rect 10539 45751 10581 45760
rect 10923 45800 10965 45809
rect 10923 45760 10924 45800
rect 10964 45760 10965 45800
rect 10923 45751 10965 45760
rect 11499 45800 11541 45809
rect 11499 45760 11500 45800
rect 11540 45760 11541 45800
rect 11499 45751 11541 45760
rect 11883 45800 11925 45809
rect 11883 45760 11884 45800
rect 11924 45760 11925 45800
rect 11883 45751 11925 45760
rect 12267 45800 12309 45809
rect 12267 45760 12268 45800
rect 12308 45760 12309 45800
rect 12267 45751 12309 45760
rect 1467 45548 1509 45557
rect 1467 45508 1468 45548
rect 1508 45508 1509 45548
rect 1467 45499 1509 45508
rect 11163 45548 11205 45557
rect 11163 45508 11164 45548
rect 11204 45508 11205 45548
rect 11163 45499 11205 45508
rect 12123 45548 12165 45557
rect 12123 45508 12124 45548
rect 12164 45508 12165 45548
rect 12123 45499 12165 45508
rect 12507 45548 12549 45557
rect 12507 45508 12508 45548
rect 12548 45508 12549 45548
rect 12507 45499 12549 45508
rect 1152 45380 12576 45404
rect 1152 45340 4928 45380
rect 4968 45340 5010 45380
rect 5050 45340 5092 45380
rect 5132 45340 5174 45380
rect 5214 45340 5256 45380
rect 5296 45340 12576 45380
rect 1152 45316 12576 45340
rect 5691 45212 5733 45221
rect 5691 45172 5692 45212
rect 5732 45172 5733 45212
rect 5691 45163 5733 45172
rect 8667 45212 8709 45221
rect 8667 45172 8668 45212
rect 8708 45172 8709 45212
rect 8667 45163 8709 45172
rect 10683 45212 10725 45221
rect 10683 45172 10684 45212
rect 10724 45172 10725 45212
rect 10683 45163 10725 45172
rect 12027 45212 12069 45221
rect 12027 45172 12028 45212
rect 12068 45172 12069 45212
rect 12027 45163 12069 45172
rect 4635 45128 4677 45137
rect 4635 45088 4636 45128
rect 4676 45088 4677 45128
rect 4635 45079 4677 45088
rect 11643 45128 11685 45137
rect 11643 45088 11644 45128
rect 11684 45088 11685 45128
rect 11643 45079 11685 45088
rect 1227 44960 1269 44969
rect 1227 44920 1228 44960
rect 1268 44920 1269 44960
rect 1227 44911 1269 44920
rect 4395 44960 4437 44969
rect 4395 44920 4396 44960
rect 4436 44920 4437 44960
rect 4395 44911 4437 44920
rect 5451 44960 5493 44969
rect 5451 44920 5452 44960
rect 5492 44920 5493 44960
rect 5451 44911 5493 44920
rect 8907 44960 8949 44969
rect 8907 44920 8908 44960
rect 8948 44920 8949 44960
rect 8907 44911 8949 44920
rect 10347 44960 10389 44969
rect 10347 44920 10348 44960
rect 10388 44920 10389 44960
rect 10347 44911 10389 44920
rect 10923 44960 10965 44969
rect 10923 44920 10924 44960
rect 10964 44920 10965 44960
rect 10923 44911 10965 44920
rect 11259 44960 11301 44969
rect 11259 44920 11260 44960
rect 11300 44920 11301 44960
rect 11259 44911 11301 44920
rect 11499 44960 11541 44969
rect 11499 44920 11500 44960
rect 11540 44920 11541 44960
rect 11499 44911 11541 44920
rect 11883 44960 11925 44969
rect 11883 44920 11884 44960
rect 11924 44920 11925 44960
rect 11883 44911 11925 44920
rect 12267 44960 12309 44969
rect 12267 44920 12268 44960
rect 12308 44920 12309 44960
rect 12267 44911 12309 44920
rect 10587 44876 10629 44885
rect 10587 44836 10588 44876
rect 10628 44836 10629 44876
rect 10587 44827 10629 44836
rect 1467 44792 1509 44801
rect 1467 44752 1468 44792
rect 1508 44752 1509 44792
rect 1467 44743 1509 44752
rect 1152 44624 12576 44648
rect 1152 44584 3688 44624
rect 3728 44584 3770 44624
rect 3810 44584 3852 44624
rect 3892 44584 3934 44624
rect 3974 44584 4016 44624
rect 4056 44584 12576 44624
rect 1152 44560 12576 44584
rect 10491 44456 10533 44465
rect 10491 44416 10492 44456
rect 10532 44416 10533 44456
rect 10491 44407 10533 44416
rect 10875 44456 10917 44465
rect 10875 44416 10876 44456
rect 10916 44416 10917 44456
rect 10875 44407 10917 44416
rect 11643 44456 11685 44465
rect 11643 44416 11644 44456
rect 11684 44416 11685 44456
rect 11643 44407 11685 44416
rect 11259 44372 11301 44381
rect 11259 44332 11260 44372
rect 11300 44332 11301 44372
rect 11259 44323 11301 44332
rect 1227 44288 1269 44297
rect 1227 44248 1228 44288
rect 1268 44248 1269 44288
rect 1227 44239 1269 44248
rect 10731 44288 10773 44297
rect 10731 44248 10732 44288
rect 10772 44248 10773 44288
rect 10731 44239 10773 44248
rect 11115 44288 11157 44297
rect 11115 44248 11116 44288
rect 11156 44248 11157 44288
rect 11115 44239 11157 44248
rect 11499 44288 11541 44297
rect 11499 44248 11500 44288
rect 11540 44248 11541 44288
rect 11499 44239 11541 44248
rect 11883 44288 11925 44297
rect 11883 44248 11884 44288
rect 11924 44248 11925 44288
rect 11883 44239 11925 44248
rect 12267 44288 12309 44297
rect 12267 44248 12268 44288
rect 12308 44248 12309 44288
rect 12267 44239 12309 44248
rect 1467 44036 1509 44045
rect 1467 43996 1468 44036
rect 1508 43996 1509 44036
rect 1467 43987 1509 43996
rect 12507 44036 12549 44045
rect 12507 43996 12508 44036
rect 12548 43996 12549 44036
rect 12507 43987 12549 43996
rect 1152 43868 12576 43892
rect 1152 43828 4928 43868
rect 4968 43828 5010 43868
rect 5050 43828 5092 43868
rect 5132 43828 5174 43868
rect 5214 43828 5256 43868
rect 5296 43828 12576 43868
rect 1152 43804 12576 43828
rect 8379 43700 8421 43709
rect 8379 43660 8380 43700
rect 8420 43660 8421 43700
rect 8379 43651 8421 43660
rect 11355 43616 11397 43625
rect 11355 43576 11356 43616
rect 11396 43576 11397 43616
rect 11355 43567 11397 43576
rect 1227 43448 1269 43457
rect 1227 43408 1228 43448
rect 1268 43408 1269 43448
rect 1227 43399 1269 43408
rect 8619 43448 8661 43457
rect 8619 43408 8620 43448
rect 8660 43408 8661 43448
rect 8619 43399 8661 43408
rect 11115 43448 11157 43457
rect 11115 43408 11116 43448
rect 11156 43408 11157 43448
rect 11115 43399 11157 43408
rect 11499 43448 11541 43457
rect 11499 43408 11500 43448
rect 11540 43408 11541 43448
rect 11499 43399 11541 43408
rect 11883 43448 11925 43457
rect 11883 43408 11884 43448
rect 11924 43408 11925 43448
rect 11883 43399 11925 43408
rect 12267 43448 12309 43457
rect 12267 43408 12268 43448
rect 12308 43408 12309 43448
rect 12267 43399 12309 43408
rect 1467 43280 1509 43289
rect 1467 43240 1468 43280
rect 1508 43240 1509 43280
rect 1467 43231 1509 43240
rect 11739 43280 11781 43289
rect 11739 43240 11740 43280
rect 11780 43240 11781 43280
rect 11739 43231 11781 43240
rect 12123 43280 12165 43289
rect 12123 43240 12124 43280
rect 12164 43240 12165 43280
rect 12123 43231 12165 43240
rect 12507 43280 12549 43289
rect 12507 43240 12508 43280
rect 12548 43240 12549 43280
rect 12507 43231 12549 43240
rect 1152 43112 12576 43136
rect 1152 43072 3688 43112
rect 3728 43072 3770 43112
rect 3810 43072 3852 43112
rect 3892 43072 3934 43112
rect 3974 43072 4016 43112
rect 4056 43072 12576 43112
rect 1152 43048 12576 43072
rect 11259 42944 11301 42953
rect 11259 42904 11260 42944
rect 11300 42904 11301 42944
rect 11259 42895 11301 42904
rect 11739 42944 11781 42953
rect 11739 42904 11740 42944
rect 11780 42904 11781 42944
rect 11739 42895 11781 42904
rect 11355 42860 11397 42869
rect 11355 42820 11356 42860
rect 11396 42820 11397 42860
rect 11355 42811 11397 42820
rect 11019 42776 11061 42785
rect 11019 42736 11020 42776
rect 11060 42736 11061 42776
rect 11019 42727 11061 42736
rect 11595 42776 11637 42785
rect 11595 42736 11596 42776
rect 11636 42736 11637 42776
rect 11595 42727 11637 42736
rect 11979 42776 12021 42785
rect 11979 42736 11980 42776
rect 12020 42736 12021 42776
rect 11979 42727 12021 42736
rect 12267 42776 12309 42785
rect 12267 42736 12268 42776
rect 12308 42736 12309 42776
rect 12267 42727 12309 42736
rect 12507 42524 12549 42533
rect 12507 42484 12508 42524
rect 12548 42484 12549 42524
rect 12507 42475 12549 42484
rect 1152 42356 12576 42380
rect 1152 42316 4928 42356
rect 4968 42316 5010 42356
rect 5050 42316 5092 42356
rect 5132 42316 5174 42356
rect 5214 42316 5256 42356
rect 5296 42316 12576 42356
rect 1152 42292 12576 42316
rect 1227 41936 1269 41945
rect 1227 41896 1228 41936
rect 1268 41896 1269 41936
rect 1227 41887 1269 41896
rect 11883 41936 11925 41945
rect 11883 41896 11884 41936
rect 11924 41896 11925 41936
rect 11883 41887 11925 41896
rect 12267 41936 12309 41945
rect 12267 41896 12268 41936
rect 12308 41896 12309 41936
rect 12267 41887 12309 41896
rect 1467 41852 1509 41861
rect 1467 41812 1468 41852
rect 1508 41812 1509 41852
rect 1467 41803 1509 41812
rect 12123 41768 12165 41777
rect 12123 41728 12124 41768
rect 12164 41728 12165 41768
rect 12123 41719 12165 41728
rect 12507 41768 12549 41777
rect 12507 41728 12508 41768
rect 12548 41728 12549 41768
rect 12507 41719 12549 41728
rect 1152 41600 12576 41624
rect 1152 41560 3688 41600
rect 3728 41560 3770 41600
rect 3810 41560 3852 41600
rect 3892 41560 3934 41600
rect 3974 41560 4016 41600
rect 4056 41560 12576 41600
rect 1152 41536 12576 41560
rect 1227 41264 1269 41273
rect 1227 41224 1228 41264
rect 1268 41224 1269 41264
rect 1227 41215 1269 41224
rect 11499 41264 11541 41273
rect 11499 41224 11500 41264
rect 11540 41224 11541 41264
rect 11499 41215 11541 41224
rect 11883 41264 11925 41273
rect 11883 41224 11884 41264
rect 11924 41224 11925 41264
rect 11883 41215 11925 41224
rect 12267 41264 12309 41273
rect 12267 41224 12268 41264
rect 12308 41224 12309 41264
rect 12267 41215 12309 41224
rect 11739 41096 11781 41105
rect 11739 41056 11740 41096
rect 11780 41056 11781 41096
rect 11739 41047 11781 41056
rect 1467 41012 1509 41021
rect 1467 40972 1468 41012
rect 1508 40972 1509 41012
rect 1467 40963 1509 40972
rect 12123 41012 12165 41021
rect 12123 40972 12124 41012
rect 12164 40972 12165 41012
rect 12123 40963 12165 40972
rect 12507 41012 12549 41021
rect 12507 40972 12508 41012
rect 12548 40972 12549 41012
rect 12507 40963 12549 40972
rect 1152 40844 12576 40868
rect 1152 40804 4928 40844
rect 4968 40804 5010 40844
rect 5050 40804 5092 40844
rect 5132 40804 5174 40844
rect 5214 40804 5256 40844
rect 5296 40804 12576 40844
rect 1152 40780 12576 40804
rect 1227 40424 1269 40433
rect 1227 40384 1228 40424
rect 1268 40384 1269 40424
rect 1227 40375 1269 40384
rect 11499 40424 11541 40433
rect 11499 40384 11500 40424
rect 11540 40384 11541 40424
rect 11499 40375 11541 40384
rect 11883 40424 11925 40433
rect 11883 40384 11884 40424
rect 11924 40384 11925 40424
rect 11883 40375 11925 40384
rect 12267 40424 12309 40433
rect 12267 40384 12268 40424
rect 12308 40384 12309 40424
rect 12267 40375 12309 40384
rect 1467 40340 1509 40349
rect 1467 40300 1468 40340
rect 1508 40300 1509 40340
rect 1467 40291 1509 40300
rect 12507 40340 12549 40349
rect 12507 40300 12508 40340
rect 12548 40300 12549 40340
rect 12507 40291 12549 40300
rect 11739 40256 11781 40265
rect 11739 40216 11740 40256
rect 11780 40216 11781 40256
rect 11739 40207 11781 40216
rect 12123 40256 12165 40265
rect 12123 40216 12124 40256
rect 12164 40216 12165 40256
rect 12123 40207 12165 40216
rect 1152 40088 12576 40112
rect 1152 40048 3688 40088
rect 3728 40048 3770 40088
rect 3810 40048 3852 40088
rect 3892 40048 3934 40088
rect 3974 40048 4016 40088
rect 4056 40048 12576 40088
rect 1152 40024 12576 40048
rect 11115 39752 11157 39761
rect 11115 39712 11116 39752
rect 11156 39712 11157 39752
rect 11115 39703 11157 39712
rect 11499 39752 11541 39761
rect 11499 39712 11500 39752
rect 11540 39712 11541 39752
rect 11499 39703 11541 39712
rect 11883 39752 11925 39761
rect 11883 39712 11884 39752
rect 11924 39712 11925 39752
rect 11883 39703 11925 39712
rect 12267 39752 12309 39761
rect 12267 39712 12268 39752
rect 12308 39712 12309 39752
rect 12267 39703 12309 39712
rect 5931 39668 5973 39677
rect 5931 39628 5932 39668
rect 5972 39628 5973 39668
rect 5931 39619 5973 39628
rect 7171 39668 7229 39669
rect 7171 39628 7180 39668
rect 7220 39628 7229 39668
rect 7171 39627 7229 39628
rect 7563 39668 7605 39677
rect 7563 39628 7564 39668
rect 7604 39628 7605 39668
rect 7563 39619 7605 39628
rect 8803 39668 8861 39669
rect 8803 39628 8812 39668
rect 8852 39628 8861 39668
rect 8803 39627 8861 39628
rect 12123 39584 12165 39593
rect 12123 39544 12124 39584
rect 12164 39544 12165 39584
rect 12123 39535 12165 39544
rect 7371 39500 7413 39509
rect 7371 39460 7372 39500
rect 7412 39460 7413 39500
rect 7371 39451 7413 39460
rect 9003 39500 9045 39509
rect 9003 39460 9004 39500
rect 9044 39460 9045 39500
rect 9003 39451 9045 39460
rect 11355 39500 11397 39509
rect 11355 39460 11356 39500
rect 11396 39460 11397 39500
rect 11355 39451 11397 39460
rect 11739 39500 11781 39509
rect 11739 39460 11740 39500
rect 11780 39460 11781 39500
rect 11739 39451 11781 39460
rect 12507 39500 12549 39509
rect 12507 39460 12508 39500
rect 12548 39460 12549 39500
rect 12507 39451 12549 39460
rect 1152 39332 12576 39356
rect 1152 39292 4928 39332
rect 4968 39292 5010 39332
rect 5050 39292 5092 39332
rect 5132 39292 5174 39332
rect 5214 39292 5256 39332
rect 5296 39292 12576 39332
rect 1152 39268 12576 39292
rect 4827 39164 4869 39173
rect 4827 39124 4828 39164
rect 4868 39124 4869 39164
rect 4827 39115 4869 39124
rect 11355 39164 11397 39173
rect 11355 39124 11356 39164
rect 11396 39124 11397 39164
rect 11355 39115 11397 39124
rect 4443 39080 4485 39089
rect 4443 39040 4444 39080
rect 4484 39040 4485 39080
rect 4443 39031 4485 39040
rect 6411 39080 6453 39089
rect 6411 39040 6412 39080
rect 6452 39040 6453 39080
rect 6411 39031 6453 39040
rect 8859 39080 8901 39089
rect 8859 39040 8860 39080
rect 8900 39040 8901 39080
rect 8859 39031 8901 39040
rect 9243 39080 9285 39089
rect 9243 39040 9244 39080
rect 9284 39040 9285 39080
rect 9243 39031 9285 39040
rect 10971 39080 11013 39089
rect 10971 39040 10972 39080
rect 11012 39040 11013 39080
rect 10971 39031 11013 39040
rect 4971 38996 5013 39005
rect 6682 38996 6740 38997
rect 4971 38956 4972 38996
rect 5012 38956 5013 38996
rect 4971 38947 5013 38956
rect 6219 38987 6261 38996
rect 6219 38947 6220 38987
rect 6260 38947 6261 38987
rect 6682 38956 6691 38996
rect 6731 38956 6740 38996
rect 6682 38955 6740 38956
rect 6795 38996 6837 39005
rect 6795 38956 6796 38996
rect 6836 38956 6837 38996
rect 6795 38947 6837 38956
rect 7179 38996 7221 39005
rect 7179 38956 7180 38996
rect 7220 38956 7221 38996
rect 7179 38947 7221 38956
rect 7755 38987 7797 38996
rect 7755 38947 7756 38987
rect 7796 38947 7797 38987
rect 6219 38938 6261 38947
rect 7755 38938 7797 38947
rect 8235 38987 8277 38996
rect 8235 38947 8236 38987
rect 8276 38947 8277 38987
rect 8235 38938 8277 38947
rect 1227 38912 1269 38921
rect 1227 38872 1228 38912
rect 1268 38872 1269 38912
rect 1227 38863 1269 38872
rect 1467 38912 1509 38921
rect 1467 38872 1468 38912
rect 1508 38872 1509 38912
rect 1467 38863 1509 38872
rect 4203 38912 4245 38921
rect 4203 38872 4204 38912
rect 4244 38872 4245 38912
rect 4203 38863 4245 38872
rect 4587 38912 4629 38921
rect 4587 38872 4588 38912
rect 4628 38872 4629 38912
rect 4587 38863 4629 38872
rect 7275 38912 7317 38921
rect 7275 38872 7276 38912
rect 7316 38872 7317 38912
rect 7275 38863 7317 38872
rect 8458 38912 8516 38913
rect 8458 38872 8467 38912
rect 8507 38872 8516 38912
rect 8458 38871 8516 38872
rect 8619 38912 8661 38921
rect 8619 38872 8620 38912
rect 8660 38872 8661 38912
rect 8619 38863 8661 38872
rect 9003 38912 9045 38921
rect 9003 38872 9004 38912
rect 9044 38872 9045 38912
rect 9003 38863 9045 38872
rect 9387 38912 9429 38921
rect 9387 38872 9388 38912
rect 9428 38872 9429 38912
rect 9387 38863 9429 38872
rect 9627 38912 9669 38921
rect 9627 38872 9628 38912
rect 9668 38872 9669 38912
rect 9627 38863 9669 38872
rect 10731 38912 10773 38921
rect 10731 38872 10732 38912
rect 10772 38872 10773 38912
rect 10731 38863 10773 38872
rect 11115 38912 11157 38921
rect 11115 38872 11116 38912
rect 11156 38872 11157 38912
rect 11115 38863 11157 38872
rect 11499 38912 11541 38921
rect 11499 38872 11500 38912
rect 11540 38872 11541 38912
rect 11499 38863 11541 38872
rect 11883 38912 11925 38921
rect 11883 38872 11884 38912
rect 11924 38872 11925 38912
rect 11883 38863 11925 38872
rect 12123 38912 12165 38921
rect 12123 38872 12124 38912
rect 12164 38872 12165 38912
rect 12123 38863 12165 38872
rect 12267 38912 12309 38921
rect 12267 38872 12268 38912
rect 12308 38872 12309 38912
rect 12267 38863 12309 38872
rect 12507 38912 12549 38921
rect 12507 38872 12508 38912
rect 12548 38872 12549 38912
rect 12507 38863 12549 38872
rect 11739 38744 11781 38753
rect 11739 38704 11740 38744
rect 11780 38704 11781 38744
rect 11739 38695 11781 38704
rect 1152 38576 12576 38600
rect 1152 38536 3688 38576
rect 3728 38536 3770 38576
rect 3810 38536 3852 38576
rect 3892 38536 3934 38576
rect 3974 38536 4016 38576
rect 4056 38536 12576 38576
rect 1152 38512 12576 38536
rect 5259 38408 5301 38417
rect 5259 38368 5260 38408
rect 5300 38368 5301 38408
rect 5259 38359 5301 38368
rect 6891 38324 6933 38333
rect 6891 38284 6892 38324
rect 6932 38284 6933 38324
rect 6891 38275 6933 38284
rect 1227 38240 1269 38249
rect 1227 38200 1228 38240
rect 1268 38200 1269 38240
rect 1227 38191 1269 38200
rect 7659 38240 7701 38249
rect 7659 38200 7660 38240
rect 7700 38200 7701 38240
rect 7659 38191 7701 38200
rect 11019 38240 11061 38249
rect 11019 38200 11020 38240
rect 11060 38200 11061 38240
rect 8715 38189 8757 38198
rect 11019 38191 11061 38200
rect 11499 38240 11541 38249
rect 11499 38200 11500 38240
rect 11540 38200 11541 38240
rect 11499 38191 11541 38200
rect 11883 38240 11925 38249
rect 11883 38200 11884 38240
rect 11924 38200 11925 38240
rect 11883 38191 11925 38200
rect 12267 38240 12309 38249
rect 12267 38200 12268 38240
rect 12308 38200 12309 38240
rect 12267 38191 12309 38200
rect 3819 38156 3861 38165
rect 3819 38116 3820 38156
rect 3860 38116 3861 38156
rect 3819 38107 3861 38116
rect 5059 38156 5117 38157
rect 5059 38116 5068 38156
rect 5108 38116 5117 38156
rect 5059 38115 5117 38116
rect 5451 38156 5493 38165
rect 5451 38116 5452 38156
rect 5492 38116 5493 38156
rect 5451 38107 5493 38116
rect 6691 38156 6749 38157
rect 6691 38116 6700 38156
rect 6740 38116 6749 38156
rect 6691 38115 6749 38116
rect 7162 38156 7220 38157
rect 7162 38116 7171 38156
rect 7211 38116 7220 38156
rect 7162 38115 7220 38116
rect 7275 38156 7317 38165
rect 7275 38116 7276 38156
rect 7316 38116 7317 38156
rect 7275 38107 7317 38116
rect 7755 38156 7797 38165
rect 7755 38116 7756 38156
rect 7796 38116 7797 38156
rect 7755 38107 7797 38116
rect 8227 38156 8285 38157
rect 8227 38116 8236 38156
rect 8276 38116 8285 38156
rect 8715 38149 8716 38189
rect 8756 38149 8757 38189
rect 8715 38140 8757 38149
rect 9099 38156 9141 38165
rect 8227 38115 8285 38116
rect 9099 38116 9100 38156
rect 9140 38116 9141 38156
rect 9099 38107 9141 38116
rect 10339 38156 10397 38157
rect 10339 38116 10348 38156
rect 10388 38116 10397 38156
rect 10339 38115 10397 38116
rect 12123 38072 12165 38081
rect 12123 38032 12124 38072
rect 12164 38032 12165 38072
rect 12123 38023 12165 38032
rect 1467 37988 1509 37997
rect 1467 37948 1468 37988
rect 1508 37948 1509 37988
rect 1467 37939 1509 37948
rect 8907 37988 8949 37997
rect 8907 37948 8908 37988
rect 8948 37948 8949 37988
rect 8907 37939 8949 37948
rect 10539 37988 10581 37997
rect 10539 37948 10540 37988
rect 10580 37948 10581 37988
rect 10539 37939 10581 37948
rect 11259 37988 11301 37997
rect 11259 37948 11260 37988
rect 11300 37948 11301 37988
rect 11259 37939 11301 37948
rect 11739 37988 11781 37997
rect 11739 37948 11740 37988
rect 11780 37948 11781 37988
rect 11739 37939 11781 37948
rect 12507 37988 12549 37997
rect 12507 37948 12508 37988
rect 12548 37948 12549 37988
rect 12507 37939 12549 37948
rect 1152 37820 12576 37844
rect 1152 37780 4928 37820
rect 4968 37780 5010 37820
rect 5050 37780 5092 37820
rect 5132 37780 5174 37820
rect 5214 37780 5256 37820
rect 5296 37780 12576 37820
rect 1152 37756 12576 37780
rect 8811 37652 8853 37661
rect 8811 37612 8812 37652
rect 8852 37612 8853 37652
rect 8811 37603 8853 37612
rect 10923 37652 10965 37661
rect 10923 37612 10924 37652
rect 10964 37612 10965 37652
rect 10923 37603 10965 37612
rect 3723 37484 3765 37493
rect 5355 37484 5397 37493
rect 7053 37484 7095 37493
rect 3723 37444 3724 37484
rect 3764 37444 3765 37484
rect 3723 37435 3765 37444
rect 4971 37475 5013 37484
rect 4971 37435 4972 37475
rect 5012 37435 5013 37475
rect 5355 37444 5356 37484
rect 5396 37444 5397 37484
rect 5355 37435 5397 37444
rect 6603 37475 6645 37484
rect 6603 37435 6604 37475
rect 6644 37435 6645 37475
rect 7053 37444 7054 37484
rect 7094 37444 7095 37484
rect 7053 37435 7095 37444
rect 7179 37484 7221 37493
rect 7179 37444 7180 37484
rect 7220 37444 7221 37484
rect 7179 37435 7221 37444
rect 7563 37484 7605 37493
rect 9178 37484 9236 37485
rect 7563 37444 7564 37484
rect 7604 37444 7605 37484
rect 7563 37435 7605 37444
rect 8139 37475 8181 37484
rect 8139 37435 8140 37475
rect 8180 37435 8181 37475
rect 4971 37426 5013 37435
rect 6603 37426 6645 37435
rect 8139 37426 8181 37435
rect 8619 37475 8661 37484
rect 8619 37435 8620 37475
rect 8660 37435 8661 37475
rect 9178 37444 9187 37484
rect 9227 37444 9236 37484
rect 9178 37443 9236 37444
rect 9291 37484 9333 37493
rect 9291 37444 9292 37484
rect 9332 37444 9333 37484
rect 9291 37435 9333 37444
rect 9675 37484 9717 37493
rect 9675 37444 9676 37484
rect 9716 37444 9717 37484
rect 9675 37435 9717 37444
rect 10251 37475 10293 37484
rect 10251 37435 10252 37475
rect 10292 37435 10293 37475
rect 8619 37426 8661 37435
rect 10251 37426 10293 37435
rect 10731 37475 10773 37484
rect 10731 37435 10732 37475
rect 10772 37435 10773 37475
rect 10731 37426 10773 37435
rect 1227 37400 1269 37409
rect 1227 37360 1228 37400
rect 1268 37360 1269 37400
rect 1227 37351 1269 37360
rect 7659 37400 7701 37409
rect 7659 37360 7660 37400
rect 7700 37360 7701 37400
rect 7659 37351 7701 37360
rect 9771 37400 9813 37409
rect 9771 37360 9772 37400
rect 9812 37360 9813 37400
rect 9771 37351 9813 37360
rect 11307 37400 11349 37409
rect 11307 37360 11308 37400
rect 11348 37360 11349 37400
rect 11307 37351 11349 37360
rect 11499 37400 11541 37409
rect 11499 37360 11500 37400
rect 11540 37360 11541 37400
rect 11499 37351 11541 37360
rect 11883 37400 11925 37409
rect 11883 37360 11884 37400
rect 11924 37360 11925 37400
rect 11883 37351 11925 37360
rect 12267 37400 12309 37409
rect 12267 37360 12268 37400
rect 12308 37360 12309 37400
rect 12267 37351 12309 37360
rect 6795 37316 6837 37325
rect 6795 37276 6796 37316
rect 6836 37276 6837 37316
rect 6795 37267 6837 37276
rect 12123 37316 12165 37325
rect 12123 37276 12124 37316
rect 12164 37276 12165 37316
rect 12123 37267 12165 37276
rect 1467 37232 1509 37241
rect 1467 37192 1468 37232
rect 1508 37192 1509 37232
rect 1467 37183 1509 37192
rect 5163 37232 5205 37241
rect 5163 37192 5164 37232
rect 5204 37192 5205 37232
rect 5163 37183 5205 37192
rect 11067 37232 11109 37241
rect 11067 37192 11068 37232
rect 11108 37192 11109 37232
rect 11067 37183 11109 37192
rect 11739 37232 11781 37241
rect 11739 37192 11740 37232
rect 11780 37192 11781 37232
rect 11739 37183 11781 37192
rect 12507 37232 12549 37241
rect 12507 37192 12508 37232
rect 12548 37192 12549 37232
rect 12507 37183 12549 37192
rect 1152 37064 12576 37088
rect 1152 37024 3688 37064
rect 3728 37024 3770 37064
rect 3810 37024 3852 37064
rect 3892 37024 3934 37064
rect 3974 37024 4016 37064
rect 4056 37024 12576 37064
rect 1152 37000 12576 37024
rect 10491 36896 10533 36905
rect 10491 36856 10492 36896
rect 10532 36856 10533 36896
rect 10491 36847 10533 36856
rect 9483 36728 9525 36737
rect 9483 36688 9484 36728
rect 9524 36688 9525 36728
rect 9483 36679 9525 36688
rect 9867 36728 9909 36737
rect 9867 36688 9868 36728
rect 9908 36688 9909 36728
rect 9867 36679 9909 36688
rect 10251 36728 10293 36737
rect 10251 36688 10252 36728
rect 10292 36688 10293 36728
rect 10251 36679 10293 36688
rect 12267 36728 12309 36737
rect 12267 36688 12268 36728
rect 12308 36688 12309 36728
rect 12267 36679 12309 36688
rect 3147 36644 3189 36653
rect 3147 36604 3148 36644
rect 3188 36604 3189 36644
rect 3147 36595 3189 36604
rect 4387 36644 4445 36645
rect 4387 36604 4396 36644
rect 4436 36604 4445 36644
rect 4387 36603 4445 36604
rect 4779 36644 4821 36653
rect 4779 36604 4780 36644
rect 4820 36604 4821 36644
rect 4779 36595 4821 36604
rect 6019 36644 6077 36645
rect 6019 36604 6028 36644
rect 6068 36604 6077 36644
rect 6019 36603 6077 36604
rect 6411 36644 6453 36653
rect 6411 36604 6412 36644
rect 6452 36604 6453 36644
rect 6411 36595 6453 36604
rect 7651 36644 7709 36645
rect 7651 36604 7660 36644
rect 7700 36604 7709 36644
rect 7651 36603 7709 36604
rect 10819 36644 10877 36645
rect 10819 36604 10828 36644
rect 10868 36604 10877 36644
rect 10819 36603 10877 36604
rect 12075 36644 12117 36653
rect 12075 36604 12076 36644
rect 12116 36604 12117 36644
rect 12075 36595 12117 36604
rect 10635 36560 10677 36569
rect 10635 36520 10636 36560
rect 10676 36520 10677 36560
rect 10635 36511 10677 36520
rect 4587 36476 4629 36485
rect 4587 36436 4588 36476
rect 4628 36436 4629 36476
rect 4587 36427 4629 36436
rect 6219 36476 6261 36485
rect 6219 36436 6220 36476
rect 6260 36436 6261 36476
rect 6219 36427 6261 36436
rect 7851 36476 7893 36485
rect 7851 36436 7852 36476
rect 7892 36436 7893 36476
rect 7851 36427 7893 36436
rect 9723 36476 9765 36485
rect 9723 36436 9724 36476
rect 9764 36436 9765 36476
rect 9723 36427 9765 36436
rect 10107 36476 10149 36485
rect 10107 36436 10108 36476
rect 10148 36436 10149 36476
rect 10107 36427 10149 36436
rect 12507 36476 12549 36485
rect 12507 36436 12508 36476
rect 12548 36436 12549 36476
rect 12507 36427 12549 36436
rect 1152 36308 12576 36332
rect 1152 36268 4928 36308
rect 4968 36268 5010 36308
rect 5050 36268 5092 36308
rect 5132 36268 5174 36308
rect 5214 36268 5256 36308
rect 5296 36268 12576 36308
rect 1152 36244 12576 36268
rect 6315 36140 6357 36149
rect 6315 36100 6316 36140
rect 6356 36100 6357 36140
rect 6315 36091 6357 36100
rect 9963 36140 10005 36149
rect 9963 36100 9964 36140
rect 10004 36100 10005 36140
rect 9963 36091 10005 36100
rect 4875 35972 4917 35981
rect 10138 35972 10196 35973
rect 11115 35972 11157 35981
rect 4875 35932 4876 35972
rect 4916 35932 4917 35972
rect 4875 35923 4917 35932
rect 6123 35963 6165 35972
rect 6123 35923 6124 35963
rect 6164 35923 6165 35963
rect 10138 35932 10147 35972
rect 10187 35932 10196 35972
rect 10138 35931 10196 35932
rect 10635 35963 10677 35972
rect 6123 35914 6165 35923
rect 10635 35923 10636 35963
rect 10676 35923 10677 35963
rect 11115 35932 11116 35972
rect 11156 35932 11157 35972
rect 11115 35923 11157 35932
rect 11595 35972 11637 35981
rect 11595 35932 11596 35972
rect 11636 35932 11637 35972
rect 11595 35923 11637 35932
rect 11705 35972 11763 35973
rect 11705 35932 11714 35972
rect 11754 35932 11763 35972
rect 11705 35931 11763 35932
rect 10635 35914 10677 35923
rect 1227 35888 1269 35897
rect 1227 35848 1228 35888
rect 1268 35848 1269 35888
rect 1227 35839 1269 35848
rect 4059 35888 4101 35897
rect 4059 35848 4060 35888
rect 4100 35848 4101 35888
rect 4059 35839 4101 35848
rect 4299 35888 4341 35897
rect 4299 35848 4300 35888
rect 4340 35848 4341 35888
rect 4299 35839 4341 35848
rect 4491 35888 4533 35897
rect 4491 35848 4492 35888
rect 4532 35848 4533 35888
rect 4491 35839 4533 35848
rect 6507 35888 6549 35897
rect 6507 35848 6508 35888
rect 6548 35848 6549 35888
rect 6507 35839 6549 35848
rect 9195 35888 9237 35897
rect 9195 35848 9196 35888
rect 9236 35848 9237 35888
rect 9195 35839 9237 35848
rect 9579 35888 9621 35897
rect 9579 35848 9580 35888
rect 9620 35848 9621 35888
rect 9579 35839 9621 35848
rect 11211 35888 11253 35897
rect 11211 35848 11212 35888
rect 11252 35848 11253 35888
rect 11211 35839 11253 35848
rect 12267 35888 12309 35897
rect 12267 35848 12268 35888
rect 12308 35848 12309 35888
rect 12267 35839 12309 35848
rect 4731 35804 4773 35813
rect 4731 35764 4732 35804
rect 4772 35764 4773 35804
rect 4731 35755 4773 35764
rect 1467 35720 1509 35729
rect 1467 35680 1468 35720
rect 1508 35680 1509 35720
rect 1467 35671 1509 35680
rect 6747 35720 6789 35729
rect 6747 35680 6748 35720
rect 6788 35680 6789 35720
rect 6747 35671 6789 35680
rect 9435 35720 9477 35729
rect 9435 35680 9436 35720
rect 9476 35680 9477 35720
rect 9435 35671 9477 35680
rect 9819 35720 9861 35729
rect 9819 35680 9820 35720
rect 9860 35680 9861 35720
rect 9819 35671 9861 35680
rect 12507 35720 12549 35729
rect 12507 35680 12508 35720
rect 12548 35680 12549 35720
rect 12507 35671 12549 35680
rect 1152 35552 12576 35576
rect 1152 35512 3688 35552
rect 3728 35512 3770 35552
rect 3810 35512 3852 35552
rect 3892 35512 3934 35552
rect 3974 35512 4016 35552
rect 4056 35512 12576 35552
rect 1152 35488 12576 35512
rect 4155 35384 4197 35393
rect 4155 35344 4156 35384
rect 4196 35344 4197 35384
rect 4155 35335 4197 35344
rect 12459 35384 12501 35393
rect 12459 35344 12460 35384
rect 12500 35344 12501 35384
rect 12459 35335 12501 35344
rect 1227 35216 1269 35225
rect 1227 35176 1228 35216
rect 1268 35176 1269 35216
rect 1227 35167 1269 35176
rect 3915 35216 3957 35225
rect 3915 35176 3916 35216
rect 3956 35176 3957 35216
rect 3915 35167 3957 35176
rect 7563 35216 7605 35225
rect 7563 35176 7564 35216
rect 7604 35176 7605 35216
rect 7563 35167 7605 35176
rect 8842 35216 8900 35217
rect 8842 35176 8851 35216
rect 8891 35176 8900 35216
rect 8842 35175 8900 35176
rect 9003 35216 9045 35225
rect 9003 35176 9004 35216
rect 9044 35176 9045 35216
rect 9003 35167 9045 35176
rect 4299 35132 4341 35141
rect 4299 35092 4300 35132
rect 4340 35092 4341 35132
rect 4299 35083 4341 35092
rect 5539 35132 5597 35133
rect 5539 35092 5548 35132
rect 5588 35092 5597 35132
rect 5539 35091 5597 35092
rect 7066 35132 7124 35133
rect 7066 35092 7075 35132
rect 7115 35092 7124 35132
rect 7066 35091 7124 35092
rect 7179 35132 7221 35141
rect 7179 35092 7180 35132
rect 7220 35092 7221 35132
rect 7179 35083 7221 35092
rect 7659 35132 7701 35141
rect 7659 35092 7660 35132
rect 7700 35092 7701 35132
rect 7659 35083 7701 35092
rect 8131 35132 8189 35133
rect 8131 35092 8140 35132
rect 8180 35092 8189 35132
rect 8131 35091 8189 35092
rect 8619 35132 8677 35133
rect 8619 35092 8628 35132
rect 8668 35092 8677 35132
rect 8619 35091 8677 35092
rect 9571 35132 9629 35133
rect 9571 35092 9580 35132
rect 9620 35092 9629 35132
rect 9571 35091 9629 35092
rect 10827 35132 10869 35141
rect 10827 35092 10828 35132
rect 10868 35092 10869 35132
rect 10827 35083 10869 35092
rect 11019 35132 11061 35141
rect 11019 35092 11020 35132
rect 11060 35092 11061 35132
rect 11019 35083 11061 35092
rect 12259 35132 12317 35133
rect 12259 35092 12268 35132
rect 12308 35092 12317 35132
rect 12259 35091 12317 35092
rect 1467 34964 1509 34973
rect 1467 34924 1468 34964
rect 1508 34924 1509 34964
rect 1467 34915 1509 34924
rect 5739 34964 5781 34973
rect 5739 34924 5740 34964
rect 5780 34924 5781 34964
rect 5739 34915 5781 34924
rect 9243 34964 9285 34973
rect 9243 34924 9244 34964
rect 9284 34924 9285 34964
rect 9243 34915 9285 34924
rect 9387 34964 9429 34973
rect 9387 34924 9388 34964
rect 9428 34924 9429 34964
rect 9387 34915 9429 34924
rect 1152 34796 12576 34820
rect 1152 34756 4928 34796
rect 4968 34756 5010 34796
rect 5050 34756 5092 34796
rect 5132 34756 5174 34796
rect 5214 34756 5256 34796
rect 5296 34756 12576 34796
rect 1152 34732 12576 34756
rect 9771 34544 9813 34553
rect 9771 34504 9772 34544
rect 9812 34504 9813 34544
rect 9771 34495 9813 34504
rect 4491 34460 4533 34469
rect 6123 34460 6165 34469
rect 7834 34460 7892 34461
rect 4491 34420 4492 34460
rect 4532 34420 4533 34460
rect 4491 34411 4533 34420
rect 5739 34451 5781 34460
rect 5739 34411 5740 34451
rect 5780 34411 5781 34451
rect 6123 34420 6124 34460
rect 6164 34420 6165 34460
rect 6123 34411 6165 34420
rect 7371 34451 7413 34460
rect 7371 34411 7372 34451
rect 7412 34411 7413 34451
rect 7834 34420 7843 34460
rect 7883 34420 7892 34460
rect 7834 34419 7892 34420
rect 7947 34460 7989 34469
rect 7947 34420 7948 34460
rect 7988 34420 7989 34460
rect 7947 34411 7989 34420
rect 8331 34460 8373 34469
rect 11211 34460 11253 34469
rect 8331 34420 8332 34460
rect 8372 34420 8373 34460
rect 8331 34411 8373 34420
rect 8907 34451 8949 34460
rect 8907 34411 8908 34451
rect 8948 34411 8949 34451
rect 5739 34402 5781 34411
rect 7371 34402 7413 34411
rect 8907 34402 8949 34411
rect 9387 34451 9429 34460
rect 9387 34411 9388 34451
rect 9428 34411 9429 34451
rect 9387 34402 9429 34411
rect 9963 34451 10005 34460
rect 9963 34411 9964 34451
rect 10004 34411 10005 34451
rect 11211 34420 11212 34460
rect 11252 34420 11253 34460
rect 11211 34411 11253 34420
rect 9963 34402 10005 34411
rect 1227 34376 1269 34385
rect 1227 34336 1228 34376
rect 1268 34336 1269 34376
rect 1227 34327 1269 34336
rect 8427 34376 8469 34385
rect 8427 34336 8428 34376
rect 8468 34336 8469 34376
rect 8427 34327 8469 34336
rect 11595 34376 11637 34385
rect 11595 34336 11596 34376
rect 11636 34336 11637 34376
rect 11595 34327 11637 34336
rect 11883 34376 11925 34385
rect 11883 34336 11884 34376
rect 11924 34336 11925 34376
rect 11883 34327 11925 34336
rect 12267 34376 12309 34385
rect 12267 34336 12268 34376
rect 12308 34336 12309 34376
rect 12267 34327 12309 34336
rect 9627 34292 9669 34301
rect 9627 34252 9628 34292
rect 9668 34252 9669 34292
rect 9627 34243 9669 34252
rect 12123 34292 12165 34301
rect 12123 34252 12124 34292
rect 12164 34252 12165 34292
rect 12123 34243 12165 34252
rect 1467 34208 1509 34217
rect 1467 34168 1468 34208
rect 1508 34168 1509 34208
rect 1467 34159 1509 34168
rect 5931 34208 5973 34217
rect 5931 34168 5932 34208
rect 5972 34168 5973 34208
rect 5931 34159 5973 34168
rect 7563 34208 7605 34217
rect 7563 34168 7564 34208
rect 7604 34168 7605 34208
rect 7563 34159 7605 34168
rect 11355 34208 11397 34217
rect 11355 34168 11356 34208
rect 11396 34168 11397 34208
rect 11355 34159 11397 34168
rect 12507 34208 12549 34217
rect 12507 34168 12508 34208
rect 12548 34168 12549 34208
rect 12507 34159 12549 34168
rect 1152 34040 12576 34064
rect 1152 34000 3688 34040
rect 3728 34000 3770 34040
rect 3810 34000 3852 34040
rect 3892 34000 3934 34040
rect 3974 34000 4016 34040
rect 4056 34000 12576 34040
rect 1152 33976 12576 34000
rect 6555 33872 6597 33881
rect 6555 33832 6556 33872
rect 6596 33832 6597 33872
rect 6555 33823 6597 33832
rect 11211 33788 11253 33797
rect 11211 33748 11212 33788
rect 11252 33748 11253 33788
rect 11211 33739 11253 33748
rect 6315 33704 6357 33713
rect 6315 33664 6316 33704
rect 6356 33664 6357 33704
rect 6315 33655 6357 33664
rect 7275 33704 7317 33713
rect 7275 33664 7276 33704
rect 7316 33664 7317 33704
rect 7275 33655 7317 33664
rect 8554 33704 8612 33705
rect 8554 33664 8563 33704
rect 8603 33664 8612 33704
rect 8554 33663 8612 33664
rect 8715 33704 8757 33713
rect 8715 33664 8716 33704
rect 8756 33664 8757 33704
rect 8715 33655 8757 33664
rect 9195 33704 9237 33713
rect 9195 33664 9196 33704
rect 9236 33664 9237 33704
rect 9195 33655 9237 33664
rect 11883 33704 11925 33713
rect 11883 33664 11884 33704
rect 11924 33664 11925 33704
rect 11883 33655 11925 33664
rect 12267 33704 12309 33713
rect 12267 33664 12268 33704
rect 12308 33664 12309 33704
rect 12267 33655 12309 33664
rect 3339 33620 3381 33629
rect 3339 33580 3340 33620
rect 3380 33580 3381 33620
rect 3339 33571 3381 33580
rect 4579 33620 4637 33621
rect 4579 33580 4588 33620
rect 4628 33580 4637 33620
rect 4579 33579 4637 33580
rect 6778 33620 6836 33621
rect 6778 33580 6787 33620
rect 6827 33580 6836 33620
rect 6778 33579 6836 33580
rect 6891 33620 6933 33629
rect 6891 33580 6892 33620
rect 6932 33580 6933 33620
rect 6891 33571 6933 33580
rect 7371 33620 7413 33629
rect 7371 33580 7372 33620
rect 7412 33580 7413 33620
rect 7371 33571 7413 33580
rect 7843 33620 7901 33621
rect 7843 33580 7852 33620
rect 7892 33580 7901 33620
rect 7843 33579 7901 33580
rect 8331 33620 8389 33621
rect 8331 33580 8340 33620
rect 8380 33580 8389 33620
rect 8331 33579 8389 33580
rect 9579 33620 9621 33629
rect 9579 33580 9580 33620
rect 9620 33580 9621 33620
rect 9579 33571 9621 33580
rect 10819 33620 10877 33621
rect 10819 33580 10828 33620
rect 10868 33580 10877 33620
rect 10819 33579 10877 33580
rect 4779 33452 4821 33461
rect 4779 33412 4780 33452
rect 4820 33412 4821 33452
rect 4779 33403 4821 33412
rect 8955 33452 8997 33461
rect 8955 33412 8956 33452
rect 8996 33412 8997 33452
rect 8955 33403 8997 33412
rect 9435 33452 9477 33461
rect 9435 33412 9436 33452
rect 9476 33412 9477 33452
rect 9435 33403 9477 33412
rect 11019 33452 11061 33461
rect 11019 33412 11020 33452
rect 11060 33412 11061 33452
rect 11019 33403 11061 33412
rect 12123 33452 12165 33461
rect 12123 33412 12124 33452
rect 12164 33412 12165 33452
rect 12123 33403 12165 33412
rect 12507 33452 12549 33461
rect 12507 33412 12508 33452
rect 12548 33412 12549 33452
rect 12507 33403 12549 33412
rect 1152 33284 12576 33308
rect 1152 33244 4928 33284
rect 4968 33244 5010 33284
rect 5050 33244 5092 33284
rect 5132 33244 5174 33284
rect 5214 33244 5256 33284
rect 5296 33244 12576 33284
rect 1152 33220 12576 33244
rect 6315 33116 6357 33125
rect 6315 33076 6316 33116
rect 6356 33076 6357 33116
rect 6315 33067 6357 33076
rect 11403 33116 11445 33125
rect 11403 33076 11404 33116
rect 11444 33076 11445 33116
rect 11403 33067 11445 33076
rect 6747 33032 6789 33041
rect 6747 32992 6748 33032
rect 6788 32992 6789 33032
rect 6747 32983 6789 32992
rect 9387 33032 9429 33041
rect 9387 32992 9388 33032
rect 9428 32992 9429 33032
rect 9387 32983 9429 32992
rect 4570 32948 4628 32949
rect 4570 32908 4579 32948
rect 4619 32908 4628 32948
rect 4570 32907 4628 32908
rect 4683 32948 4725 32957
rect 4683 32908 4684 32948
rect 4724 32908 4725 32948
rect 4683 32899 4725 32908
rect 5067 32948 5109 32957
rect 7947 32948 7989 32957
rect 5067 32908 5068 32948
rect 5108 32908 5109 32948
rect 5067 32899 5109 32908
rect 5643 32939 5685 32948
rect 5643 32899 5644 32939
rect 5684 32899 5685 32939
rect 5643 32890 5685 32899
rect 6123 32939 6165 32948
rect 6123 32899 6124 32939
rect 6164 32899 6165 32939
rect 7947 32908 7948 32948
rect 7988 32908 7989 32948
rect 7947 32899 7989 32908
rect 9658 32948 9716 32949
rect 9658 32908 9667 32948
rect 9707 32908 9716 32948
rect 9658 32907 9716 32908
rect 9771 32948 9813 32957
rect 9771 32908 9772 32948
rect 9812 32908 9813 32948
rect 9191 32906 9249 32907
rect 6123 32890 6165 32899
rect 1227 32864 1269 32873
rect 1227 32824 1228 32864
rect 1268 32824 1269 32864
rect 1227 32815 1269 32824
rect 3723 32864 3765 32873
rect 3723 32824 3724 32864
rect 3764 32824 3765 32864
rect 3723 32815 3765 32824
rect 4107 32864 4149 32873
rect 4107 32824 4108 32864
rect 4148 32824 4149 32864
rect 4107 32815 4149 32824
rect 5163 32864 5205 32873
rect 5163 32824 5164 32864
rect 5204 32824 5205 32864
rect 5163 32815 5205 32824
rect 6538 32864 6596 32865
rect 6538 32824 6547 32864
rect 6587 32824 6596 32864
rect 6538 32823 6596 32824
rect 6891 32864 6933 32873
rect 6891 32824 6892 32864
rect 6932 32824 6933 32864
rect 6891 32815 6933 32824
rect 7563 32864 7605 32873
rect 9191 32866 9200 32906
rect 9240 32866 9249 32906
rect 9771 32899 9813 32908
rect 10251 32948 10293 32957
rect 10251 32908 10252 32948
rect 10292 32908 10293 32948
rect 10251 32899 10293 32908
rect 10731 32939 10773 32948
rect 10731 32899 10732 32939
rect 10772 32899 10773 32939
rect 10731 32890 10773 32899
rect 11211 32939 11253 32948
rect 11211 32899 11212 32939
rect 11252 32899 11253 32939
rect 11211 32890 11253 32899
rect 9191 32865 9249 32866
rect 7563 32824 7564 32864
rect 7604 32824 7605 32864
rect 7563 32815 7605 32824
rect 10155 32864 10197 32873
rect 10155 32824 10156 32864
rect 10196 32824 10197 32864
rect 10155 32815 10197 32824
rect 11883 32864 11925 32873
rect 11883 32824 11884 32864
rect 11924 32824 11925 32864
rect 11883 32815 11925 32824
rect 12267 32864 12309 32873
rect 12267 32824 12268 32864
rect 12308 32824 12309 32864
rect 12267 32815 12309 32824
rect 3963 32780 4005 32789
rect 3963 32740 3964 32780
rect 4004 32740 4005 32780
rect 3963 32731 4005 32740
rect 7803 32780 7845 32789
rect 7803 32740 7804 32780
rect 7844 32740 7845 32780
rect 7803 32731 7845 32740
rect 1467 32696 1509 32705
rect 1467 32656 1468 32696
rect 1508 32656 1509 32696
rect 1467 32647 1509 32656
rect 4347 32696 4389 32705
rect 4347 32656 4348 32696
rect 4388 32656 4389 32696
rect 4347 32647 4389 32656
rect 7131 32696 7173 32705
rect 7131 32656 7132 32696
rect 7172 32656 7173 32696
rect 7131 32647 7173 32656
rect 12123 32696 12165 32705
rect 12123 32656 12124 32696
rect 12164 32656 12165 32696
rect 12123 32647 12165 32656
rect 12507 32696 12549 32705
rect 12507 32656 12508 32696
rect 12548 32656 12549 32696
rect 12507 32647 12549 32656
rect 1152 32528 12576 32552
rect 1152 32488 3688 32528
rect 3728 32488 3770 32528
rect 3810 32488 3852 32528
rect 3892 32488 3934 32528
rect 3974 32488 4016 32528
rect 4056 32488 12576 32528
rect 1152 32464 12576 32488
rect 9819 32360 9861 32369
rect 9819 32320 9820 32360
rect 9860 32320 9861 32360
rect 9819 32311 9861 32320
rect 12459 32360 12501 32369
rect 12459 32320 12460 32360
rect 12500 32320 12501 32360
rect 12459 32311 12501 32320
rect 1227 32192 1269 32201
rect 1227 32152 1228 32192
rect 1268 32152 1269 32192
rect 1227 32143 1269 32152
rect 4875 32192 4917 32201
rect 4875 32152 4876 32192
rect 4916 32152 4917 32192
rect 4875 32143 4917 32152
rect 6315 32192 6357 32201
rect 6315 32152 6316 32192
rect 6356 32152 6357 32192
rect 6315 32143 6357 32152
rect 9579 32192 9621 32201
rect 9579 32152 9580 32192
rect 9620 32152 9621 32192
rect 9579 32143 9621 32152
rect 2667 32108 2709 32117
rect 2667 32068 2668 32108
rect 2708 32068 2709 32108
rect 2667 32059 2709 32068
rect 3907 32108 3965 32109
rect 3907 32068 3916 32108
rect 3956 32068 3965 32108
rect 3907 32067 3965 32068
rect 4365 32108 4407 32117
rect 4365 32068 4366 32108
rect 4406 32068 4407 32108
rect 4365 32059 4407 32068
rect 4491 32108 4533 32117
rect 4491 32068 4492 32108
rect 4532 32068 4533 32108
rect 4491 32059 4533 32068
rect 4971 32108 5013 32117
rect 4971 32068 4972 32108
rect 5012 32068 5013 32108
rect 4971 32059 5013 32068
rect 5443 32108 5501 32109
rect 5443 32068 5452 32108
rect 5492 32068 5501 32108
rect 5443 32067 5501 32068
rect 5931 32108 5989 32109
rect 5931 32068 5940 32108
rect 5980 32068 5989 32108
rect 5931 32067 5989 32068
rect 7947 32108 7989 32117
rect 7947 32068 7948 32108
rect 7988 32068 7989 32108
rect 7947 32059 7989 32068
rect 9187 32108 9245 32109
rect 9187 32068 9196 32108
rect 9236 32068 9245 32108
rect 9187 32067 9245 32068
rect 10522 32108 10580 32109
rect 10522 32068 10531 32108
rect 10571 32068 10580 32108
rect 10522 32067 10580 32068
rect 10138 32024 10196 32025
rect 10138 31984 10147 32024
rect 10187 31984 10196 32024
rect 10138 31983 10196 31984
rect 1467 31940 1509 31949
rect 1467 31900 1468 31940
rect 1508 31900 1509 31940
rect 1467 31891 1509 31900
rect 4107 31940 4149 31949
rect 4107 31900 4108 31940
rect 4148 31900 4149 31940
rect 4107 31891 4149 31900
rect 6123 31940 6165 31949
rect 6123 31900 6124 31940
rect 6164 31900 6165 31940
rect 6123 31891 6165 31900
rect 6555 31940 6597 31949
rect 6555 31900 6556 31940
rect 6596 31900 6597 31940
rect 6555 31891 6597 31900
rect 9387 31940 9429 31949
rect 9387 31900 9388 31940
rect 9428 31900 9429 31940
rect 9387 31891 9429 31900
rect 12459 31940 12501 31949
rect 12459 31900 12460 31940
rect 12500 31900 12501 31940
rect 12459 31891 12501 31900
rect 1152 31772 12576 31796
rect 1152 31732 4928 31772
rect 4968 31732 5010 31772
rect 5050 31732 5092 31772
rect 5132 31732 5174 31772
rect 5214 31732 5256 31772
rect 5296 31732 12576 31772
rect 1152 31708 12576 31732
rect 4299 31604 4341 31613
rect 4299 31564 4300 31604
rect 4340 31564 4341 31604
rect 4299 31555 4341 31564
rect 6315 31604 6357 31613
rect 6315 31564 6316 31604
rect 6356 31564 6357 31604
rect 6315 31555 6357 31564
rect 6843 31604 6885 31613
rect 6843 31564 6844 31604
rect 6884 31564 6885 31604
rect 6843 31555 6885 31564
rect 9243 31604 9285 31613
rect 9243 31564 9244 31604
rect 9284 31564 9285 31604
rect 9243 31555 9285 31564
rect 2859 31436 2901 31445
rect 4570 31436 4628 31437
rect 2859 31396 2860 31436
rect 2900 31396 2901 31436
rect 2859 31387 2901 31396
rect 4107 31427 4149 31436
rect 4107 31387 4108 31427
rect 4148 31387 4149 31427
rect 4570 31396 4579 31436
rect 4619 31396 4628 31436
rect 4570 31395 4628 31396
rect 4683 31436 4725 31445
rect 4683 31396 4684 31436
rect 4724 31396 4725 31436
rect 4683 31387 4725 31396
rect 5067 31436 5109 31445
rect 8811 31436 8853 31445
rect 5067 31396 5068 31436
rect 5108 31396 5109 31436
rect 5067 31387 5109 31396
rect 5643 31427 5685 31436
rect 5643 31387 5644 31427
rect 5684 31387 5685 31427
rect 4107 31378 4149 31387
rect 5643 31378 5685 31387
rect 6123 31427 6165 31436
rect 6123 31387 6124 31427
rect 6164 31387 6165 31427
rect 6123 31378 6165 31387
rect 7563 31427 7605 31436
rect 7563 31387 7564 31427
rect 7604 31387 7605 31427
rect 8811 31396 8812 31436
rect 8852 31396 8853 31436
rect 8811 31387 8853 31396
rect 9579 31436 9621 31445
rect 9579 31396 9580 31436
rect 9620 31396 9621 31436
rect 9579 31387 9621 31396
rect 10827 31427 10869 31436
rect 10827 31387 10828 31427
rect 10868 31387 10869 31427
rect 7563 31378 7605 31387
rect 10827 31378 10869 31387
rect 1227 31352 1269 31361
rect 1227 31312 1228 31352
rect 1268 31312 1269 31352
rect 1227 31303 1269 31312
rect 5163 31352 5205 31361
rect 5163 31312 5164 31352
rect 5204 31312 5205 31352
rect 5163 31303 5205 31312
rect 6699 31352 6741 31361
rect 6699 31312 6700 31352
rect 6740 31312 6741 31352
rect 6699 31303 6741 31312
rect 7083 31352 7125 31361
rect 7083 31312 7084 31352
rect 7124 31312 7125 31352
rect 7083 31303 7125 31312
rect 9003 31352 9045 31361
rect 9003 31312 9004 31352
rect 9044 31312 9045 31352
rect 9003 31303 9045 31312
rect 11499 31352 11541 31361
rect 11499 31312 11500 31352
rect 11540 31312 11541 31352
rect 11499 31303 11541 31312
rect 11883 31352 11925 31361
rect 11883 31312 11884 31352
rect 11924 31312 11925 31352
rect 11883 31303 11925 31312
rect 12267 31352 12309 31361
rect 12267 31312 12268 31352
rect 12308 31312 12309 31352
rect 12267 31303 12309 31312
rect 12123 31268 12165 31277
rect 12123 31228 12124 31268
rect 12164 31228 12165 31268
rect 12123 31219 12165 31228
rect 1467 31184 1509 31193
rect 1467 31144 1468 31184
rect 1508 31144 1509 31184
rect 1467 31135 1509 31144
rect 6459 31184 6501 31193
rect 6459 31144 6460 31184
rect 6500 31144 6501 31184
rect 6459 31135 6501 31144
rect 7371 31184 7413 31193
rect 7371 31144 7372 31184
rect 7412 31144 7413 31184
rect 7371 31135 7413 31144
rect 11019 31184 11061 31193
rect 11019 31144 11020 31184
rect 11060 31144 11061 31184
rect 11019 31135 11061 31144
rect 11739 31184 11781 31193
rect 11739 31144 11740 31184
rect 11780 31144 11781 31184
rect 11739 31135 11781 31144
rect 12507 31184 12549 31193
rect 12507 31144 12508 31184
rect 12548 31144 12549 31184
rect 12507 31135 12549 31144
rect 1152 31016 12576 31040
rect 1152 30976 3688 31016
rect 3728 30976 3770 31016
rect 3810 30976 3852 31016
rect 3892 30976 3934 31016
rect 3974 30976 4016 31016
rect 4056 30976 12576 31016
rect 1152 30952 12576 30976
rect 3675 30848 3717 30857
rect 3675 30808 3676 30848
rect 3716 30808 3717 30848
rect 3675 30799 3717 30808
rect 8091 30848 8133 30857
rect 8091 30808 8092 30848
rect 8132 30808 8133 30848
rect 8091 30799 8133 30808
rect 11643 30848 11685 30857
rect 11643 30808 11644 30848
rect 11684 30808 11685 30848
rect 11643 30799 11685 30808
rect 10827 30764 10869 30773
rect 10827 30724 10828 30764
rect 10868 30724 10869 30764
rect 10827 30715 10869 30724
rect 3435 30680 3477 30689
rect 3435 30640 3436 30680
rect 3476 30640 3477 30680
rect 3435 30631 3477 30640
rect 6027 30680 6069 30689
rect 6027 30640 6028 30680
rect 6068 30640 6069 30680
rect 6027 30631 6069 30640
rect 7306 30680 7364 30681
rect 7306 30640 7315 30680
rect 7355 30640 7364 30680
rect 7306 30639 7364 30640
rect 7467 30680 7509 30689
rect 7467 30640 7468 30680
rect 7508 30640 7509 30680
rect 7467 30631 7509 30640
rect 7851 30680 7893 30689
rect 7851 30640 7852 30680
rect 7892 30640 7893 30680
rect 7851 30631 7893 30640
rect 8187 30680 8229 30689
rect 8187 30640 8188 30680
rect 8228 30640 8229 30680
rect 8187 30631 8229 30640
rect 8427 30680 8469 30689
rect 8427 30640 8428 30680
rect 8468 30640 8469 30680
rect 8427 30631 8469 30640
rect 10443 30680 10485 30689
rect 10443 30640 10444 30680
rect 10484 30640 10485 30680
rect 10443 30631 10485 30640
rect 11019 30680 11061 30689
rect 11019 30640 11020 30680
rect 11060 30640 11061 30680
rect 11019 30631 11061 30640
rect 11403 30680 11445 30689
rect 11403 30640 11404 30680
rect 11444 30640 11445 30680
rect 11403 30631 11445 30640
rect 11883 30680 11925 30689
rect 11883 30640 11884 30680
rect 11924 30640 11925 30680
rect 11883 30631 11925 30640
rect 12267 30680 12309 30689
rect 12267 30640 12268 30680
rect 12308 30640 12309 30680
rect 12267 30631 12309 30640
rect 3819 30596 3861 30605
rect 3819 30556 3820 30596
rect 3860 30556 3861 30596
rect 3819 30547 3861 30556
rect 5059 30596 5117 30597
rect 5059 30556 5068 30596
rect 5108 30556 5117 30596
rect 5059 30555 5117 30556
rect 5530 30596 5588 30597
rect 5530 30556 5539 30596
rect 5579 30556 5588 30596
rect 5530 30555 5588 30556
rect 5643 30596 5685 30605
rect 5643 30556 5644 30596
rect 5684 30556 5685 30596
rect 5643 30547 5685 30556
rect 6123 30596 6165 30605
rect 6123 30556 6124 30596
rect 6164 30556 6165 30596
rect 6123 30547 6165 30556
rect 6595 30596 6653 30597
rect 6595 30556 6604 30596
rect 6644 30556 6653 30596
rect 6595 30555 6653 30556
rect 7114 30596 7172 30597
rect 7114 30556 7123 30596
rect 7163 30556 7172 30596
rect 7114 30555 7172 30556
rect 8619 30596 8661 30605
rect 8619 30556 8620 30596
rect 8660 30556 8661 30596
rect 8619 30547 8661 30556
rect 9859 30596 9917 30597
rect 9859 30556 9868 30596
rect 9908 30556 9917 30596
rect 9859 30555 9917 30556
rect 5259 30512 5301 30521
rect 5259 30472 5260 30512
rect 5300 30472 5301 30512
rect 5259 30463 5301 30472
rect 10059 30512 10101 30521
rect 10059 30472 10060 30512
rect 10100 30472 10101 30512
rect 10059 30463 10101 30472
rect 12123 30512 12165 30521
rect 12123 30472 12124 30512
rect 12164 30472 12165 30512
rect 12123 30463 12165 30472
rect 7707 30428 7749 30437
rect 7707 30388 7708 30428
rect 7748 30388 7749 30428
rect 7707 30379 7749 30388
rect 10203 30428 10245 30437
rect 10203 30388 10204 30428
rect 10244 30388 10245 30428
rect 10203 30379 10245 30388
rect 11259 30428 11301 30437
rect 11259 30388 11260 30428
rect 11300 30388 11301 30428
rect 11259 30379 11301 30388
rect 12507 30428 12549 30437
rect 12507 30388 12508 30428
rect 12548 30388 12549 30428
rect 12507 30379 12549 30388
rect 1152 30260 12576 30284
rect 1152 30220 4928 30260
rect 4968 30220 5010 30260
rect 5050 30220 5092 30260
rect 5132 30220 5174 30260
rect 5214 30220 5256 30260
rect 5296 30220 12576 30260
rect 1152 30196 12576 30220
rect 7467 30092 7509 30101
rect 7467 30052 7468 30092
rect 7508 30052 7509 30092
rect 7467 30043 7509 30052
rect 8283 30092 8325 30101
rect 8283 30052 8284 30092
rect 8324 30052 8325 30092
rect 8283 30043 8325 30052
rect 7899 30008 7941 30017
rect 7899 29968 7900 30008
rect 7940 29968 7941 30008
rect 7899 29959 7941 29968
rect 4077 29924 4119 29933
rect 4077 29884 4078 29924
rect 4118 29884 4119 29924
rect 4077 29875 4119 29884
rect 4203 29924 4245 29933
rect 4203 29884 4204 29924
rect 4244 29884 4245 29924
rect 4203 29875 4245 29884
rect 4587 29924 4629 29933
rect 6027 29924 6069 29933
rect 10155 29924 10197 29933
rect 4587 29884 4588 29924
rect 4628 29884 4629 29924
rect 4587 29875 4629 29884
rect 5163 29915 5205 29924
rect 5163 29875 5164 29915
rect 5204 29875 5205 29915
rect 5163 29866 5205 29875
rect 5643 29915 5685 29924
rect 5643 29875 5644 29915
rect 5684 29875 5685 29915
rect 6027 29884 6028 29924
rect 6068 29884 6069 29924
rect 6027 29875 6069 29884
rect 7275 29915 7317 29924
rect 7275 29875 7276 29915
rect 7316 29875 7317 29915
rect 10155 29884 10156 29924
rect 10196 29884 10197 29924
rect 10155 29875 10197 29884
rect 10522 29924 10580 29925
rect 10522 29884 10531 29924
rect 10571 29884 10580 29924
rect 10522 29883 10580 29884
rect 5643 29866 5685 29875
rect 7275 29866 7317 29875
rect 1227 29840 1269 29849
rect 1227 29800 1228 29840
rect 1268 29800 1269 29840
rect 1227 29791 1269 29800
rect 4683 29840 4725 29849
rect 4683 29800 4684 29840
rect 4724 29800 4725 29840
rect 4683 29791 4725 29800
rect 7659 29840 7701 29849
rect 7659 29800 7660 29840
rect 7700 29800 7701 29840
rect 7659 29791 7701 29800
rect 8043 29840 8085 29849
rect 8043 29800 8044 29840
rect 8084 29800 8085 29840
rect 8043 29791 8085 29800
rect 9387 29840 9429 29849
rect 9387 29800 9388 29840
rect 9428 29800 9429 29840
rect 9387 29791 9429 29800
rect 9771 29840 9813 29849
rect 9771 29800 9772 29840
rect 9812 29800 9813 29840
rect 9771 29791 9813 29800
rect 10011 29840 10053 29849
rect 10011 29800 10012 29840
rect 10052 29800 10053 29840
rect 10011 29791 10053 29800
rect 9627 29756 9669 29765
rect 9627 29716 9628 29756
rect 9668 29716 9669 29756
rect 9627 29707 9669 29716
rect 1467 29672 1509 29681
rect 1467 29632 1468 29672
rect 1508 29632 1509 29672
rect 1467 29623 1509 29632
rect 5866 29672 5924 29673
rect 5866 29632 5875 29672
rect 5915 29632 5924 29672
rect 5866 29631 5924 29632
rect 12459 29672 12501 29681
rect 12459 29632 12460 29672
rect 12500 29632 12501 29672
rect 12459 29623 12501 29632
rect 1152 29504 12576 29528
rect 1152 29464 3688 29504
rect 3728 29464 3770 29504
rect 3810 29464 3852 29504
rect 3892 29464 3934 29504
rect 3974 29464 4016 29504
rect 4056 29464 12576 29504
rect 1152 29440 12576 29464
rect 1467 29336 1509 29345
rect 1467 29296 1468 29336
rect 1508 29296 1509 29336
rect 1467 29287 1509 29296
rect 2619 29336 2661 29345
rect 2619 29296 2620 29336
rect 2660 29296 2661 29336
rect 2619 29287 2661 29296
rect 4587 29336 4629 29345
rect 4587 29296 4588 29336
rect 4628 29296 4629 29336
rect 4587 29287 4629 29296
rect 5979 29336 6021 29345
rect 5979 29296 5980 29336
rect 6020 29296 6021 29336
rect 5979 29287 6021 29296
rect 5595 29252 5637 29261
rect 5595 29212 5596 29252
rect 5636 29212 5637 29252
rect 5595 29203 5637 29212
rect 1227 29168 1269 29177
rect 1227 29128 1228 29168
rect 1268 29128 1269 29168
rect 1227 29119 1269 29128
rect 2379 29168 2421 29177
rect 2379 29128 2380 29168
rect 2420 29128 2421 29168
rect 2379 29119 2421 29128
rect 5355 29168 5397 29177
rect 5355 29128 5356 29168
rect 5396 29128 5397 29168
rect 5355 29119 5397 29128
rect 5739 29168 5781 29177
rect 5739 29128 5740 29168
rect 5780 29128 5781 29168
rect 5739 29119 5781 29128
rect 10347 29168 10389 29177
rect 10347 29128 10348 29168
rect 10388 29128 10389 29168
rect 10347 29119 10389 29128
rect 11883 29168 11925 29177
rect 11883 29128 11884 29168
rect 11924 29128 11925 29168
rect 11883 29119 11925 29128
rect 12267 29168 12309 29177
rect 12267 29128 12268 29168
rect 12308 29128 12309 29168
rect 12267 29119 12309 29128
rect 3147 29084 3189 29093
rect 3147 29044 3148 29084
rect 3188 29044 3189 29084
rect 3147 29035 3189 29044
rect 4387 29084 4445 29085
rect 4387 29044 4396 29084
rect 4436 29044 4445 29084
rect 4387 29043 4445 29044
rect 6411 29084 6453 29093
rect 6411 29044 6412 29084
rect 6452 29044 6453 29084
rect 6411 29035 6453 29044
rect 7651 29084 7709 29085
rect 7651 29044 7660 29084
rect 7700 29044 7709 29084
rect 7651 29043 7709 29044
rect 8043 29084 8085 29093
rect 8043 29044 8044 29084
rect 8084 29044 8085 29084
rect 8043 29035 8085 29044
rect 9283 29084 9341 29085
rect 9283 29044 9292 29084
rect 9332 29044 9341 29084
rect 9283 29043 9341 29044
rect 9850 29084 9908 29085
rect 9850 29044 9859 29084
rect 9899 29044 9908 29084
rect 9850 29043 9908 29044
rect 9963 29084 10005 29093
rect 9963 29044 9964 29084
rect 10004 29044 10005 29084
rect 9963 29035 10005 29044
rect 10443 29084 10485 29093
rect 10443 29044 10444 29084
rect 10484 29044 10485 29084
rect 10443 29035 10485 29044
rect 10914 29084 10972 29085
rect 10914 29044 10923 29084
rect 10963 29044 10972 29084
rect 10914 29043 10972 29044
rect 11403 29084 11461 29085
rect 11403 29044 11412 29084
rect 11452 29044 11461 29084
rect 11403 29043 11461 29044
rect 7851 28916 7893 28925
rect 7851 28876 7852 28916
rect 7892 28876 7893 28916
rect 7851 28867 7893 28876
rect 9483 28916 9525 28925
rect 9483 28876 9484 28916
rect 9524 28876 9525 28916
rect 9483 28867 9525 28876
rect 11595 28916 11637 28925
rect 11595 28876 11596 28916
rect 11636 28876 11637 28916
rect 11595 28867 11637 28876
rect 12123 28916 12165 28925
rect 12123 28876 12124 28916
rect 12164 28876 12165 28916
rect 12123 28867 12165 28876
rect 12507 28916 12549 28925
rect 12507 28876 12508 28916
rect 12548 28876 12549 28916
rect 12507 28867 12549 28876
rect 1152 28748 12576 28772
rect 1152 28708 4928 28748
rect 4968 28708 5010 28748
rect 5050 28708 5092 28748
rect 5132 28708 5174 28748
rect 5214 28708 5256 28748
rect 5296 28708 12576 28748
rect 1152 28684 12576 28708
rect 1467 28580 1509 28589
rect 1467 28540 1468 28580
rect 1508 28540 1509 28580
rect 1467 28531 1509 28540
rect 4011 28580 4053 28589
rect 4011 28540 4012 28580
rect 4052 28540 4053 28580
rect 4011 28531 4053 28540
rect 10347 28580 10389 28589
rect 10347 28540 10348 28580
rect 10388 28540 10389 28580
rect 10347 28531 10389 28540
rect 2571 28412 2613 28421
rect 6891 28412 6933 28421
rect 8602 28412 8660 28413
rect 2571 28372 2572 28412
rect 2612 28372 2613 28412
rect 2571 28363 2613 28372
rect 3819 28403 3861 28412
rect 3819 28363 3820 28403
rect 3860 28363 3861 28403
rect 6891 28372 6892 28412
rect 6932 28372 6933 28412
rect 6891 28363 6933 28372
rect 8139 28403 8181 28412
rect 8139 28363 8140 28403
rect 8180 28363 8181 28403
rect 8602 28372 8611 28412
rect 8651 28372 8660 28412
rect 8602 28371 8660 28372
rect 8715 28412 8757 28421
rect 8715 28372 8716 28412
rect 8756 28372 8757 28412
rect 8715 28363 8757 28372
rect 9099 28412 9141 28421
rect 10539 28412 10581 28421
rect 9099 28372 9100 28412
rect 9140 28372 9141 28412
rect 9099 28363 9141 28372
rect 9675 28403 9717 28412
rect 9675 28363 9676 28403
rect 9716 28363 9717 28403
rect 3819 28354 3861 28363
rect 8139 28354 8181 28363
rect 9675 28354 9717 28363
rect 10155 28403 10197 28412
rect 10155 28363 10156 28403
rect 10196 28363 10197 28403
rect 10539 28372 10540 28412
rect 10580 28372 10581 28412
rect 10539 28363 10581 28372
rect 11787 28403 11829 28412
rect 11787 28363 11788 28403
rect 11828 28363 11829 28403
rect 10155 28354 10197 28363
rect 11787 28354 11829 28363
rect 1227 28328 1269 28337
rect 1227 28288 1228 28328
rect 1268 28288 1269 28328
rect 1227 28279 1269 28288
rect 9195 28328 9237 28337
rect 9195 28288 9196 28328
rect 9236 28288 9237 28328
rect 9195 28279 9237 28288
rect 12363 28328 12405 28337
rect 12363 28288 12364 28328
rect 12404 28288 12405 28328
rect 12363 28279 12405 28288
rect 8331 28160 8373 28169
rect 8331 28120 8332 28160
rect 8372 28120 8373 28160
rect 8331 28111 8373 28120
rect 11979 28160 12021 28169
rect 11979 28120 11980 28160
rect 12020 28120 12021 28160
rect 11979 28111 12021 28120
rect 12123 28160 12165 28169
rect 12123 28120 12124 28160
rect 12164 28120 12165 28160
rect 12123 28111 12165 28120
rect 1152 27992 12576 28016
rect 1152 27952 3688 27992
rect 3728 27952 3770 27992
rect 3810 27952 3852 27992
rect 3892 27952 3934 27992
rect 3974 27952 4016 27992
rect 4056 27952 12576 27992
rect 1152 27928 12576 27952
rect 10570 27824 10628 27825
rect 10570 27784 10579 27824
rect 10619 27784 10628 27824
rect 10570 27783 10628 27784
rect 9291 27656 9333 27665
rect 9291 27616 9292 27656
rect 9332 27616 9333 27656
rect 9291 27607 9333 27616
rect 4299 27572 4341 27581
rect 4299 27532 4300 27572
rect 4340 27532 4341 27572
rect 4299 27523 4341 27532
rect 5539 27572 5597 27573
rect 5539 27532 5548 27572
rect 5588 27532 5597 27572
rect 5539 27531 5597 27532
rect 6795 27572 6837 27581
rect 6795 27532 6796 27572
rect 6836 27532 6837 27572
rect 6795 27523 6837 27532
rect 8035 27572 8093 27573
rect 8035 27532 8044 27572
rect 8084 27532 8093 27572
rect 8035 27531 8093 27532
rect 8794 27572 8852 27573
rect 8794 27532 8803 27572
rect 8843 27532 8852 27572
rect 8794 27531 8852 27532
rect 8907 27572 8949 27581
rect 8907 27532 8908 27572
rect 8948 27532 8949 27572
rect 8907 27523 8949 27532
rect 9387 27572 9429 27581
rect 9387 27532 9388 27572
rect 9428 27532 9429 27572
rect 9387 27523 9429 27532
rect 9859 27572 9917 27573
rect 9859 27532 9868 27572
rect 9908 27532 9917 27572
rect 9859 27531 9917 27532
rect 10347 27572 10405 27573
rect 10347 27532 10356 27572
rect 10396 27532 10405 27572
rect 10347 27531 10405 27532
rect 10915 27572 10973 27573
rect 10915 27532 10924 27572
rect 10964 27532 10973 27572
rect 10915 27531 10973 27532
rect 12171 27572 12213 27581
rect 12171 27532 12172 27572
rect 12212 27532 12213 27572
rect 12171 27523 12213 27532
rect 8235 27488 8277 27497
rect 8235 27448 8236 27488
rect 8276 27448 8277 27488
rect 8235 27439 8277 27448
rect 5739 27404 5781 27413
rect 5739 27364 5740 27404
rect 5780 27364 5781 27404
rect 5739 27355 5781 27364
rect 10731 27404 10773 27413
rect 10731 27364 10732 27404
rect 10772 27364 10773 27404
rect 10731 27355 10773 27364
rect 1152 27236 12576 27260
rect 1152 27196 4928 27236
rect 4968 27196 5010 27236
rect 5050 27196 5092 27236
rect 5132 27196 5174 27236
rect 5214 27196 5256 27236
rect 5296 27196 12576 27236
rect 1152 27172 12576 27196
rect 1467 27068 1509 27077
rect 1467 27028 1468 27068
rect 1508 27028 1509 27068
rect 1467 27019 1509 27028
rect 6555 27068 6597 27077
rect 6555 27028 6556 27068
rect 6596 27028 6597 27068
rect 6555 27019 6597 27028
rect 12027 27068 12069 27077
rect 12027 27028 12028 27068
rect 12068 27028 12069 27068
rect 12027 27019 12069 27028
rect 4107 26984 4149 26993
rect 4107 26944 4108 26984
rect 4148 26944 4149 26984
rect 4107 26935 4149 26944
rect 2667 26900 2709 26909
rect 4378 26900 4436 26901
rect 2667 26860 2668 26900
rect 2708 26860 2709 26900
rect 2667 26851 2709 26860
rect 3915 26891 3957 26900
rect 3915 26851 3916 26891
rect 3956 26851 3957 26891
rect 4378 26860 4387 26900
rect 4427 26860 4436 26900
rect 4378 26859 4436 26860
rect 4491 26900 4533 26909
rect 4491 26860 4492 26900
rect 4532 26860 4533 26900
rect 4491 26851 4533 26860
rect 4875 26900 4917 26909
rect 7222 26900 7264 26909
rect 4875 26860 4876 26900
rect 4916 26860 4917 26900
rect 4875 26851 4917 26860
rect 5451 26891 5493 26900
rect 5451 26851 5452 26891
rect 5492 26851 5493 26891
rect 3915 26842 3957 26851
rect 5451 26842 5493 26851
rect 5931 26891 5973 26900
rect 5931 26851 5932 26891
rect 5972 26851 5973 26891
rect 7222 26860 7223 26900
rect 7263 26860 7264 26900
rect 7222 26851 7264 26860
rect 7467 26900 7509 26909
rect 7467 26860 7468 26900
rect 7508 26860 7509 26900
rect 7467 26851 7509 26860
rect 9754 26900 9812 26901
rect 9754 26860 9763 26900
rect 9803 26860 9812 26900
rect 9754 26859 9812 26860
rect 9867 26900 9909 26909
rect 9867 26860 9868 26900
rect 9908 26860 9909 26900
rect 9867 26851 9909 26860
rect 10251 26900 10293 26909
rect 10251 26860 10252 26900
rect 10292 26860 10293 26900
rect 10251 26851 10293 26860
rect 10827 26891 10869 26900
rect 10827 26851 10828 26891
rect 10868 26851 10869 26891
rect 5931 26842 5973 26851
rect 10827 26842 10869 26851
rect 11307 26891 11349 26900
rect 11307 26851 11308 26891
rect 11348 26851 11349 26891
rect 11307 26842 11349 26851
rect 1227 26816 1269 26825
rect 1227 26776 1228 26816
rect 1268 26776 1269 26816
rect 1227 26767 1269 26776
rect 4971 26816 5013 26825
rect 4971 26776 4972 26816
rect 5012 26776 5013 26816
rect 4971 26767 5013 26776
rect 6154 26816 6212 26817
rect 6154 26776 6163 26816
rect 6203 26776 6212 26816
rect 6154 26775 6212 26776
rect 6315 26816 6357 26825
rect 6315 26776 6316 26816
rect 6356 26776 6357 26816
rect 6315 26767 6357 26776
rect 7354 26816 7412 26817
rect 7354 26776 7363 26816
rect 7403 26776 7412 26816
rect 7354 26775 7412 26776
rect 7563 26816 7605 26825
rect 7563 26776 7564 26816
rect 7604 26776 7605 26816
rect 7563 26767 7605 26776
rect 10347 26816 10389 26825
rect 10347 26776 10348 26816
rect 10388 26776 10389 26816
rect 10347 26767 10389 26776
rect 11691 26816 11733 26825
rect 11691 26776 11692 26816
rect 11732 26776 11733 26816
rect 11691 26767 11733 26776
rect 12267 26816 12309 26825
rect 12267 26776 12268 26816
rect 12308 26776 12309 26816
rect 12267 26767 12309 26776
rect 11530 26648 11588 26649
rect 11530 26608 11539 26648
rect 11579 26608 11588 26648
rect 11530 26607 11588 26608
rect 11931 26648 11973 26657
rect 11931 26608 11932 26648
rect 11972 26608 11973 26648
rect 11931 26599 11973 26608
rect 1152 26480 12576 26504
rect 1152 26440 3688 26480
rect 3728 26440 3770 26480
rect 3810 26440 3852 26480
rect 3892 26440 3934 26480
rect 3974 26440 4016 26480
rect 4056 26440 12576 26480
rect 1152 26416 12576 26440
rect 4731 26312 4773 26321
rect 4731 26272 4732 26312
rect 4772 26272 4773 26312
rect 4731 26263 4773 26272
rect 11722 26312 11780 26313
rect 11722 26272 11731 26312
rect 11771 26272 11780 26312
rect 11722 26271 11780 26272
rect 6699 26228 6741 26237
rect 6699 26188 6700 26228
rect 6740 26188 6741 26228
rect 6699 26179 6741 26188
rect 4491 26144 4533 26153
rect 4491 26104 4492 26144
rect 4532 26104 4533 26144
rect 4491 26095 4533 26104
rect 10443 26144 10485 26153
rect 10443 26104 10444 26144
rect 10484 26104 10485 26144
rect 8662 26093 8704 26102
rect 10443 26095 10485 26104
rect 12075 26144 12117 26153
rect 12075 26104 12076 26144
rect 12116 26104 12117 26144
rect 12075 26095 12117 26104
rect 12267 26144 12309 26153
rect 12267 26104 12268 26144
rect 12308 26104 12309 26144
rect 12267 26095 12309 26104
rect 1411 26060 1469 26061
rect 1411 26020 1420 26060
rect 1460 26020 1469 26060
rect 1411 26019 1469 26020
rect 2667 26060 2709 26069
rect 2667 26020 2668 26060
rect 2708 26020 2709 26060
rect 2667 26011 2709 26020
rect 3043 26060 3101 26061
rect 3043 26020 3052 26060
rect 3092 26020 3101 26060
rect 3043 26019 3101 26020
rect 4299 26060 4341 26069
rect 4299 26020 4300 26060
rect 4340 26020 4341 26060
rect 4299 26011 4341 26020
rect 5259 26060 5301 26069
rect 5259 26020 5260 26060
rect 5300 26020 5301 26060
rect 5259 26011 5301 26020
rect 6499 26060 6557 26061
rect 6499 26020 6508 26060
rect 6548 26020 6557 26060
rect 6499 26019 6557 26020
rect 6891 26060 6933 26069
rect 6891 26020 6892 26060
rect 6932 26020 6933 26060
rect 6891 26011 6933 26020
rect 8131 26060 8189 26061
rect 8131 26020 8140 26060
rect 8180 26020 8189 26060
rect 8131 26019 8189 26020
rect 8523 26060 8565 26069
rect 8523 26020 8524 26060
rect 8564 26020 8565 26060
rect 8662 26053 8663 26093
rect 8703 26053 8704 26093
rect 8662 26044 8704 26053
rect 9946 26060 10004 26061
rect 8523 26011 8565 26020
rect 9946 26020 9955 26060
rect 9995 26020 10004 26060
rect 9946 26019 10004 26020
rect 10059 26060 10101 26069
rect 10059 26020 10060 26060
rect 10100 26020 10101 26060
rect 10059 26011 10101 26020
rect 10539 26060 10581 26069
rect 10539 26020 10540 26060
rect 10580 26020 10581 26060
rect 10539 26011 10581 26020
rect 11006 26060 11064 26061
rect 11006 26020 11015 26060
rect 11055 26020 11064 26060
rect 11006 26019 11064 26020
rect 11530 26060 11588 26061
rect 11530 26020 11539 26060
rect 11579 26020 11588 26060
rect 11530 26019 11588 26020
rect 1227 25976 1269 25985
rect 1227 25936 1228 25976
rect 1268 25936 1269 25976
rect 1227 25927 1269 25936
rect 8331 25976 8373 25985
rect 8331 25936 8332 25976
rect 8372 25936 8373 25976
rect 8331 25927 8373 25936
rect 11835 25976 11877 25985
rect 11835 25936 11836 25976
rect 11876 25936 11877 25976
rect 11835 25927 11877 25936
rect 2859 25892 2901 25901
rect 2859 25852 2860 25892
rect 2900 25852 2901 25892
rect 2859 25843 2901 25852
rect 8811 25892 8853 25901
rect 8811 25852 8812 25892
rect 8852 25852 8853 25892
rect 8811 25843 8853 25852
rect 12507 25892 12549 25901
rect 12507 25852 12508 25892
rect 12548 25852 12549 25892
rect 12507 25843 12549 25852
rect 1152 25724 12576 25748
rect 1152 25684 4928 25724
rect 4968 25684 5010 25724
rect 5050 25684 5092 25724
rect 5132 25684 5174 25724
rect 5214 25684 5256 25724
rect 5296 25684 12576 25724
rect 1152 25660 12576 25684
rect 1467 25556 1509 25565
rect 1467 25516 1468 25556
rect 1508 25516 1509 25556
rect 1467 25507 1509 25516
rect 8026 25556 8084 25557
rect 8026 25516 8035 25556
rect 8075 25516 8084 25556
rect 8026 25515 8084 25516
rect 9771 25556 9813 25565
rect 9771 25516 9772 25556
rect 9812 25516 9813 25556
rect 9771 25507 9813 25516
rect 12507 25556 12549 25565
rect 12507 25516 12508 25556
rect 12548 25516 12549 25556
rect 12507 25507 12549 25516
rect 8794 25472 8852 25473
rect 8794 25432 8803 25472
rect 8843 25432 8852 25472
rect 8794 25431 8852 25432
rect 4203 25388 4245 25397
rect 2955 25379 2997 25388
rect 2955 25339 2956 25379
rect 2996 25339 2997 25379
rect 4203 25348 4204 25388
rect 4244 25348 4245 25388
rect 4203 25339 4245 25348
rect 4683 25388 4725 25397
rect 6315 25388 6357 25397
rect 8187 25388 8229 25397
rect 4683 25348 4684 25388
rect 4724 25348 4725 25388
rect 4683 25339 4725 25348
rect 5931 25379 5973 25388
rect 5931 25339 5932 25379
rect 5972 25339 5973 25379
rect 6315 25348 6316 25388
rect 6356 25348 6357 25388
rect 6315 25339 6357 25348
rect 7563 25379 7605 25388
rect 7563 25339 7564 25379
rect 7604 25339 7605 25379
rect 8187 25348 8188 25388
rect 8228 25348 8229 25388
rect 8187 25339 8229 25348
rect 8331 25388 8373 25397
rect 8331 25348 8332 25388
rect 8372 25348 8373 25388
rect 8715 25388 8757 25397
rect 8331 25339 8373 25348
rect 8475 25346 8517 25355
rect 2955 25330 2997 25339
rect 5931 25330 5973 25339
rect 7563 25330 7605 25339
rect 1227 25304 1269 25313
rect 1227 25264 1228 25304
rect 1268 25264 1269 25304
rect 1227 25255 1269 25264
rect 1611 25304 1653 25313
rect 1611 25264 1612 25304
rect 1652 25264 1653 25304
rect 8475 25306 8476 25346
rect 8516 25306 8517 25346
rect 8715 25348 8716 25388
rect 8756 25348 8757 25388
rect 8715 25339 8757 25348
rect 8950 25388 8992 25397
rect 8950 25348 8951 25388
rect 8991 25348 8992 25388
rect 8950 25339 8992 25348
rect 9195 25388 9237 25397
rect 11211 25388 11253 25397
rect 9195 25348 9196 25388
rect 9236 25348 9237 25388
rect 9195 25339 9237 25348
rect 9963 25379 10005 25388
rect 9963 25339 9964 25379
rect 10004 25339 10005 25379
rect 11211 25348 11212 25388
rect 11252 25348 11253 25388
rect 11211 25339 11253 25348
rect 9963 25330 10005 25339
rect 8475 25297 8517 25306
rect 8602 25304 8660 25305
rect 1611 25255 1653 25264
rect 8602 25264 8611 25304
rect 8651 25264 8660 25304
rect 8602 25263 8660 25264
rect 9082 25304 9140 25305
rect 9082 25264 9091 25304
rect 9131 25264 9140 25304
rect 9082 25263 9140 25264
rect 9291 25304 9333 25313
rect 9291 25264 9292 25304
rect 9332 25264 9333 25304
rect 9291 25255 9333 25264
rect 11499 25304 11541 25313
rect 11499 25264 11500 25304
rect 11540 25264 11541 25304
rect 11499 25255 11541 25264
rect 11883 25304 11925 25313
rect 11883 25264 11884 25304
rect 11924 25264 11925 25304
rect 11883 25255 11925 25264
rect 12267 25304 12309 25313
rect 12267 25264 12268 25304
rect 12308 25264 12309 25304
rect 12267 25255 12309 25264
rect 12123 25220 12165 25229
rect 12123 25180 12124 25220
rect 12164 25180 12165 25220
rect 12123 25171 12165 25180
rect 1851 25136 1893 25145
rect 1851 25096 1852 25136
rect 1892 25096 1893 25136
rect 1851 25087 1893 25096
rect 2763 25136 2805 25145
rect 2763 25096 2764 25136
rect 2804 25096 2805 25136
rect 2763 25087 2805 25096
rect 6123 25136 6165 25145
rect 6123 25096 6124 25136
rect 6164 25096 6165 25136
rect 6123 25087 6165 25096
rect 7755 25136 7797 25145
rect 7755 25096 7756 25136
rect 7796 25096 7797 25136
rect 7755 25087 7797 25096
rect 11739 25136 11781 25145
rect 11739 25096 11740 25136
rect 11780 25096 11781 25136
rect 11739 25087 11781 25096
rect 1152 24968 12576 24992
rect 1152 24928 3688 24968
rect 3728 24928 3770 24968
rect 3810 24928 3852 24968
rect 3892 24928 3934 24968
rect 3974 24928 4016 24968
rect 4056 24928 12576 24968
rect 1152 24904 12576 24928
rect 4731 24800 4773 24809
rect 4731 24760 4732 24800
rect 4772 24760 4773 24800
rect 4731 24751 4773 24760
rect 8650 24800 8708 24801
rect 8650 24760 8659 24800
rect 8699 24760 8708 24800
rect 8650 24759 8708 24760
rect 12075 24800 12117 24809
rect 12075 24760 12076 24800
rect 12116 24760 12117 24800
rect 12075 24751 12117 24760
rect 12507 24800 12549 24809
rect 12507 24760 12508 24800
rect 12548 24760 12549 24800
rect 12507 24751 12549 24760
rect 2170 24632 2228 24633
rect 2170 24592 2179 24632
rect 2219 24592 2228 24632
rect 2170 24591 2228 24592
rect 4491 24632 4533 24641
rect 4491 24592 4492 24632
rect 4532 24592 4533 24632
rect 4491 24583 4533 24592
rect 7371 24632 7413 24641
rect 7371 24592 7372 24632
rect 7412 24592 7413 24632
rect 7371 24583 7413 24592
rect 12267 24632 12309 24641
rect 12267 24592 12268 24632
rect 12308 24592 12309 24632
rect 12267 24583 12309 24592
rect 2371 24548 2429 24549
rect 2371 24508 2380 24548
rect 2420 24508 2429 24548
rect 2371 24507 2429 24508
rect 3627 24548 3669 24557
rect 3627 24508 3628 24548
rect 3668 24508 3669 24548
rect 3627 24499 3669 24508
rect 6874 24548 6932 24549
rect 6874 24508 6883 24548
rect 6923 24508 6932 24548
rect 6874 24507 6932 24508
rect 6987 24548 7029 24557
rect 6987 24508 6988 24548
rect 7028 24508 7029 24548
rect 6987 24499 7029 24508
rect 7467 24548 7509 24557
rect 7467 24508 7468 24548
rect 7508 24508 7509 24548
rect 7467 24499 7509 24508
rect 7939 24548 7997 24549
rect 7939 24508 7948 24548
rect 7988 24508 7997 24548
rect 7939 24507 7997 24508
rect 8427 24548 8485 24549
rect 8427 24508 8436 24548
rect 8476 24508 8485 24548
rect 8427 24507 8485 24508
rect 8811 24548 8853 24557
rect 8811 24508 8812 24548
rect 8852 24508 8853 24548
rect 8811 24499 8853 24508
rect 10051 24548 10109 24549
rect 10051 24508 10060 24548
rect 10100 24508 10109 24548
rect 10051 24507 10109 24508
rect 10635 24548 10677 24557
rect 10635 24508 10636 24548
rect 10676 24508 10677 24548
rect 10635 24499 10677 24508
rect 11875 24548 11933 24549
rect 11875 24508 11884 24548
rect 11924 24508 11933 24548
rect 11875 24507 11933 24508
rect 10251 24380 10293 24389
rect 10251 24340 10252 24380
rect 10292 24340 10293 24380
rect 10251 24331 10293 24340
rect 1152 24212 12576 24236
rect 1152 24172 4928 24212
rect 4968 24172 5010 24212
rect 5050 24172 5092 24212
rect 5132 24172 5174 24212
rect 5214 24172 5256 24212
rect 5296 24172 12576 24212
rect 1152 24148 12576 24172
rect 10011 24044 10053 24053
rect 10011 24004 10012 24044
rect 10052 24004 10053 24044
rect 10011 23995 10053 24004
rect 10683 24044 10725 24053
rect 10683 24004 10684 24044
rect 10724 24004 10725 24044
rect 10683 23995 10725 24004
rect 4107 23876 4149 23885
rect 5739 23876 5781 23885
rect 7834 23876 7892 23877
rect 4107 23836 4108 23876
rect 4148 23836 4149 23876
rect 4107 23827 4149 23836
rect 5355 23867 5397 23876
rect 5355 23827 5356 23867
rect 5396 23827 5397 23867
rect 5739 23836 5740 23876
rect 5780 23836 5781 23876
rect 5739 23827 5781 23836
rect 6987 23867 7029 23876
rect 6987 23827 6988 23867
rect 7028 23827 7029 23867
rect 7834 23836 7843 23876
rect 7883 23836 7892 23876
rect 7834 23835 7892 23836
rect 7947 23876 7989 23885
rect 7947 23836 7948 23876
rect 7988 23836 7989 23876
rect 7947 23827 7989 23836
rect 8331 23876 8373 23885
rect 12267 23876 12309 23885
rect 8331 23836 8332 23876
rect 8372 23836 8373 23876
rect 8331 23827 8373 23836
rect 8907 23867 8949 23876
rect 8907 23827 8908 23867
rect 8948 23827 8949 23867
rect 5355 23818 5397 23827
rect 6987 23818 7029 23827
rect 8907 23818 8949 23827
rect 9387 23867 9429 23876
rect 9387 23827 9388 23867
rect 9428 23827 9429 23867
rect 9387 23818 9429 23827
rect 11019 23867 11061 23876
rect 11019 23827 11020 23867
rect 11060 23827 11061 23867
rect 12267 23836 12268 23876
rect 12308 23836 12309 23876
rect 12267 23827 12309 23836
rect 11019 23818 11061 23827
rect 1227 23792 1269 23801
rect 1227 23752 1228 23792
rect 1268 23752 1269 23792
rect 1227 23743 1269 23752
rect 8427 23792 8469 23801
rect 8427 23752 8428 23792
rect 8468 23752 8469 23792
rect 8427 23743 8469 23752
rect 9610 23792 9668 23793
rect 9610 23752 9619 23792
rect 9659 23752 9668 23792
rect 9610 23751 9668 23752
rect 9771 23792 9813 23801
rect 9771 23752 9772 23792
rect 9812 23752 9813 23792
rect 9771 23743 9813 23752
rect 10443 23792 10485 23801
rect 10443 23752 10444 23792
rect 10484 23752 10485 23792
rect 10443 23743 10485 23752
rect 1467 23624 1509 23633
rect 1467 23584 1468 23624
rect 1508 23584 1509 23624
rect 1467 23575 1509 23584
rect 5547 23624 5589 23633
rect 5547 23584 5548 23624
rect 5588 23584 5589 23624
rect 5547 23575 5589 23584
rect 7179 23624 7221 23633
rect 7179 23584 7180 23624
rect 7220 23584 7221 23624
rect 7179 23575 7221 23584
rect 10827 23624 10869 23633
rect 10827 23584 10828 23624
rect 10868 23584 10869 23624
rect 10827 23575 10869 23584
rect 1152 23456 12576 23480
rect 1152 23416 3688 23456
rect 3728 23416 3770 23456
rect 3810 23416 3852 23456
rect 3892 23416 3934 23456
rect 3974 23416 4016 23456
rect 4056 23416 12576 23456
rect 1152 23392 12576 23416
rect 6363 23288 6405 23297
rect 6363 23248 6364 23288
rect 6404 23248 6405 23288
rect 6363 23239 6405 23248
rect 9819 23288 9861 23297
rect 9819 23248 9820 23288
rect 9860 23248 9861 23288
rect 9819 23239 9861 23248
rect 10203 23288 10245 23297
rect 10203 23248 10204 23288
rect 10244 23248 10245 23288
rect 10203 23239 10245 23248
rect 9435 23204 9477 23213
rect 9435 23164 9436 23204
rect 9476 23164 9477 23204
rect 9435 23155 9477 23164
rect 10827 23204 10869 23213
rect 10827 23164 10828 23204
rect 10868 23164 10869 23204
rect 10827 23155 10869 23164
rect 1227 23120 1269 23129
rect 1227 23080 1228 23120
rect 1268 23080 1269 23120
rect 1227 23071 1269 23080
rect 1467 23120 1509 23129
rect 1467 23080 1468 23120
rect 1508 23080 1509 23120
rect 1467 23071 1509 23080
rect 4683 23120 4725 23129
rect 4683 23080 4684 23120
rect 4724 23080 4725 23120
rect 4683 23071 4725 23080
rect 5962 23120 6020 23121
rect 5962 23080 5971 23120
rect 6011 23080 6020 23120
rect 5962 23079 6020 23080
rect 6123 23120 6165 23129
rect 6123 23080 6124 23120
rect 6164 23080 6165 23120
rect 6123 23071 6165 23080
rect 8139 23120 8181 23129
rect 8139 23080 8140 23120
rect 8180 23080 8181 23120
rect 8139 23071 8181 23080
rect 9579 23120 9621 23129
rect 9579 23080 9580 23120
rect 9620 23080 9621 23120
rect 9579 23071 9621 23080
rect 9963 23120 10005 23129
rect 9963 23080 9964 23120
rect 10004 23080 10005 23120
rect 9963 23071 10005 23080
rect 10347 23120 10389 23129
rect 10347 23080 10348 23120
rect 10388 23080 10389 23120
rect 10347 23071 10389 23080
rect 10587 23120 10629 23129
rect 10587 23080 10588 23120
rect 10628 23080 10629 23120
rect 10587 23071 10629 23080
rect 2475 23036 2517 23045
rect 2475 22996 2476 23036
rect 2516 22996 2517 23036
rect 2475 22987 2517 22996
rect 3715 23036 3773 23037
rect 3715 22996 3724 23036
rect 3764 22996 3773 23036
rect 3715 22995 3773 22996
rect 4173 23036 4215 23045
rect 4173 22996 4174 23036
rect 4214 22996 4215 23036
rect 4173 22987 4215 22996
rect 4297 23036 4339 23045
rect 4297 22996 4298 23036
rect 4338 22996 4339 23036
rect 4297 22987 4339 22996
rect 4779 23036 4821 23045
rect 4779 22996 4780 23036
rect 4820 22996 4821 23036
rect 4779 22987 4821 22996
rect 5251 23036 5309 23037
rect 5251 22996 5260 23036
rect 5300 22996 5309 23036
rect 5251 22995 5309 22996
rect 5739 23036 5797 23037
rect 5739 22996 5748 23036
rect 5788 22996 5797 23036
rect 5739 22995 5797 22996
rect 7642 23036 7700 23037
rect 7642 22996 7651 23036
rect 7691 22996 7700 23036
rect 7642 22995 7700 22996
rect 7755 23036 7797 23045
rect 7755 22996 7756 23036
rect 7796 22996 7797 23036
rect 7755 22987 7797 22996
rect 8235 23036 8277 23045
rect 8235 22996 8236 23036
rect 8276 22996 8277 23036
rect 8235 22987 8277 22996
rect 8707 23036 8765 23037
rect 8707 22996 8716 23036
rect 8756 22996 8765 23036
rect 8707 22995 8765 22996
rect 9195 23036 9253 23037
rect 9195 22996 9204 23036
rect 9244 22996 9253 23036
rect 9195 22995 9253 22996
rect 11011 23036 11069 23037
rect 11011 22996 11020 23036
rect 11060 22996 11069 23036
rect 11011 22995 11069 22996
rect 12267 23036 12309 23045
rect 12267 22996 12268 23036
rect 12308 22996 12309 23036
rect 12267 22987 12309 22996
rect 3915 22868 3957 22877
rect 3915 22828 3916 22868
rect 3956 22828 3957 22868
rect 3915 22819 3957 22828
rect 1152 22700 12576 22724
rect 1152 22660 4928 22700
rect 4968 22660 5010 22700
rect 5050 22660 5092 22700
rect 5132 22660 5174 22700
rect 5214 22660 5256 22700
rect 5296 22660 12576 22700
rect 1152 22636 12576 22660
rect 9099 22532 9141 22541
rect 9099 22492 9100 22532
rect 9140 22492 9141 22532
rect 9099 22483 9141 22492
rect 9915 22532 9957 22541
rect 9915 22492 9916 22532
rect 9956 22492 9957 22532
rect 9915 22483 9957 22492
rect 10299 22532 10341 22541
rect 10299 22492 10300 22532
rect 10340 22492 10341 22532
rect 10299 22483 10341 22492
rect 10683 22532 10725 22541
rect 10683 22492 10684 22532
rect 10724 22492 10725 22532
rect 10683 22483 10725 22492
rect 7131 22448 7173 22457
rect 7131 22408 7132 22448
rect 7172 22408 7173 22448
rect 7131 22399 7173 22408
rect 2859 22364 2901 22373
rect 4570 22364 4628 22365
rect 2859 22324 2860 22364
rect 2900 22324 2901 22364
rect 2859 22315 2901 22324
rect 4107 22355 4149 22364
rect 4107 22315 4108 22355
rect 4148 22315 4149 22355
rect 4570 22324 4579 22364
rect 4619 22324 4628 22364
rect 4570 22323 4628 22324
rect 4683 22364 4725 22373
rect 4683 22324 4684 22364
rect 4724 22324 4725 22364
rect 4683 22315 4725 22324
rect 5067 22364 5109 22373
rect 7354 22364 7412 22365
rect 5067 22324 5068 22364
rect 5108 22324 5109 22364
rect 5067 22315 5109 22324
rect 5643 22355 5685 22364
rect 5643 22315 5644 22355
rect 5684 22315 5685 22355
rect 4107 22306 4149 22315
rect 5643 22306 5685 22315
rect 6123 22355 6165 22364
rect 6123 22315 6124 22355
rect 6164 22315 6165 22355
rect 7354 22324 7363 22364
rect 7403 22324 7412 22364
rect 7354 22323 7412 22324
rect 7467 22364 7509 22373
rect 7467 22324 7468 22364
rect 7508 22324 7509 22364
rect 7467 22315 7509 22324
rect 7851 22364 7893 22373
rect 12267 22364 12309 22373
rect 7851 22324 7852 22364
rect 7892 22324 7893 22364
rect 7851 22315 7893 22324
rect 8427 22355 8469 22364
rect 8427 22315 8428 22355
rect 8468 22315 8469 22355
rect 6123 22306 6165 22315
rect 8427 22306 8469 22315
rect 8907 22355 8949 22364
rect 8907 22315 8908 22355
rect 8948 22315 8949 22355
rect 8907 22306 8949 22315
rect 11019 22355 11061 22364
rect 11019 22315 11020 22355
rect 11060 22315 11061 22355
rect 12267 22324 12268 22364
rect 12308 22324 12309 22364
rect 12267 22315 12309 22324
rect 11019 22306 11061 22315
rect 1227 22280 1269 22289
rect 1227 22240 1228 22280
rect 1268 22240 1269 22280
rect 1227 22231 1269 22240
rect 5163 22280 5205 22289
rect 5163 22240 5164 22280
rect 5204 22240 5205 22280
rect 5163 22231 5205 22240
rect 6346 22280 6404 22281
rect 6346 22240 6355 22280
rect 6395 22240 6404 22280
rect 6346 22239 6404 22240
rect 6507 22280 6549 22289
rect 6507 22240 6508 22280
rect 6548 22240 6549 22280
rect 6507 22231 6549 22240
rect 6891 22280 6933 22289
rect 6891 22240 6892 22280
rect 6932 22240 6933 22280
rect 6891 22231 6933 22240
rect 7947 22280 7989 22289
rect 7947 22240 7948 22280
rect 7988 22240 7989 22280
rect 7947 22231 7989 22240
rect 9291 22280 9333 22289
rect 9291 22240 9292 22280
rect 9332 22240 9333 22280
rect 9291 22231 9333 22240
rect 9675 22280 9717 22289
rect 9675 22240 9676 22280
rect 9716 22240 9717 22280
rect 9675 22231 9717 22240
rect 10059 22280 10101 22289
rect 10059 22240 10060 22280
rect 10100 22240 10101 22280
rect 10059 22231 10101 22240
rect 10443 22280 10485 22289
rect 10443 22240 10444 22280
rect 10484 22240 10485 22280
rect 10443 22231 10485 22240
rect 6747 22196 6789 22205
rect 6747 22156 6748 22196
rect 6788 22156 6789 22196
rect 6747 22147 6789 22156
rect 9531 22196 9573 22205
rect 9531 22156 9532 22196
rect 9572 22156 9573 22196
rect 9531 22147 9573 22156
rect 1467 22112 1509 22121
rect 1467 22072 1468 22112
rect 1508 22072 1509 22112
rect 1467 22063 1509 22072
rect 4299 22112 4341 22121
rect 4299 22072 4300 22112
rect 4340 22072 4341 22112
rect 4299 22063 4341 22072
rect 10827 22112 10869 22121
rect 10827 22072 10828 22112
rect 10868 22072 10869 22112
rect 10827 22063 10869 22072
rect 1152 21944 12576 21968
rect 1152 21904 3688 21944
rect 3728 21904 3770 21944
rect 3810 21904 3852 21944
rect 3892 21904 3934 21944
rect 3974 21904 4016 21944
rect 4056 21904 12576 21944
rect 1152 21880 12576 21904
rect 4107 21776 4149 21785
rect 4107 21736 4108 21776
rect 4148 21736 4149 21776
rect 4107 21727 4149 21736
rect 2283 21608 2325 21617
rect 2283 21568 2284 21608
rect 2324 21568 2325 21608
rect 2283 21559 2325 21568
rect 4395 21608 4437 21617
rect 4395 21568 4396 21608
rect 4436 21568 4437 21608
rect 4395 21559 4437 21568
rect 5355 21608 5397 21617
rect 5355 21568 5356 21608
rect 5396 21568 5397 21608
rect 5355 21559 5397 21568
rect 8907 21608 8949 21617
rect 8907 21568 8908 21608
rect 8948 21568 8949 21608
rect 8907 21559 8949 21568
rect 9291 21608 9333 21617
rect 9291 21568 9292 21608
rect 9332 21568 9333 21608
rect 9291 21559 9333 21568
rect 9675 21608 9717 21617
rect 9675 21568 9676 21608
rect 9716 21568 9717 21608
rect 9675 21559 9717 21568
rect 10251 21608 10293 21617
rect 10251 21568 10252 21608
rect 10292 21568 10293 21608
rect 10251 21559 10293 21568
rect 10443 21608 10485 21617
rect 10443 21568 10444 21608
rect 10484 21568 10485 21608
rect 10443 21559 10485 21568
rect 10683 21608 10725 21617
rect 10683 21568 10684 21608
rect 10724 21568 10725 21608
rect 10683 21559 10725 21568
rect 2667 21524 2709 21533
rect 2667 21484 2668 21524
rect 2708 21484 2709 21524
rect 2667 21475 2709 21484
rect 3907 21524 3965 21525
rect 3907 21484 3916 21524
rect 3956 21484 3965 21524
rect 3907 21483 3965 21484
rect 4858 21524 4916 21525
rect 4858 21484 4867 21524
rect 4907 21484 4916 21524
rect 4858 21483 4916 21484
rect 4971 21524 5013 21533
rect 4971 21484 4972 21524
rect 5012 21484 5013 21524
rect 4971 21475 5013 21484
rect 5451 21524 5493 21533
rect 5451 21484 5452 21524
rect 5492 21484 5493 21524
rect 5451 21475 5493 21484
rect 5923 21524 5981 21525
rect 5923 21484 5932 21524
rect 5972 21484 5981 21524
rect 5923 21483 5981 21484
rect 6442 21524 6500 21525
rect 6442 21484 6451 21524
rect 6491 21484 6500 21524
rect 6442 21483 6500 21484
rect 6795 21524 6837 21533
rect 6795 21484 6796 21524
rect 6836 21484 6837 21524
rect 6795 21475 6837 21484
rect 8035 21524 8093 21525
rect 8035 21484 8044 21524
rect 8084 21484 8093 21524
rect 8035 21483 8093 21484
rect 11011 21524 11069 21525
rect 11011 21484 11020 21524
rect 11060 21484 11069 21524
rect 11011 21483 11069 21484
rect 12267 21524 12309 21533
rect 12267 21484 12268 21524
rect 12308 21484 12309 21524
rect 12267 21475 12309 21484
rect 2523 21440 2565 21449
rect 2523 21400 2524 21440
rect 2564 21400 2565 21440
rect 2523 21391 2565 21400
rect 8235 21440 8277 21449
rect 8235 21400 8236 21440
rect 8276 21400 8277 21440
rect 8235 21391 8277 21400
rect 9915 21440 9957 21449
rect 9915 21400 9916 21440
rect 9956 21400 9957 21440
rect 9915 21391 9957 21400
rect 4635 21356 4677 21365
rect 4635 21316 4636 21356
rect 4676 21316 4677 21356
rect 4635 21307 4677 21316
rect 6603 21356 6645 21365
rect 6603 21316 6604 21356
rect 6644 21316 6645 21356
rect 6603 21307 6645 21316
rect 9147 21356 9189 21365
rect 9147 21316 9148 21356
rect 9188 21316 9189 21356
rect 9147 21307 9189 21316
rect 9531 21356 9573 21365
rect 9531 21316 9532 21356
rect 9572 21316 9573 21356
rect 9531 21307 9573 21316
rect 10011 21356 10053 21365
rect 10011 21316 10012 21356
rect 10052 21316 10053 21356
rect 10011 21307 10053 21316
rect 10827 21356 10869 21365
rect 10827 21316 10828 21356
rect 10868 21316 10869 21356
rect 10827 21307 10869 21316
rect 1152 21188 12576 21212
rect 1152 21148 4928 21188
rect 4968 21148 5010 21188
rect 5050 21148 5092 21188
rect 5132 21148 5174 21188
rect 5214 21148 5256 21188
rect 5296 21148 12576 21188
rect 1152 21124 12576 21148
rect 3819 21020 3861 21029
rect 3819 20980 3820 21020
rect 3860 20980 3861 21020
rect 3819 20971 3861 20980
rect 7275 21020 7317 21029
rect 7275 20980 7276 21020
rect 7316 20980 7317 21020
rect 7275 20971 7317 20980
rect 8379 21020 8421 21029
rect 8379 20980 8380 21020
rect 8420 20980 8421 21020
rect 8379 20971 8421 20980
rect 12123 21020 12165 21029
rect 12123 20980 12124 21020
rect 12164 20980 12165 21020
rect 12123 20971 12165 20980
rect 12507 21020 12549 21029
rect 12507 20980 12508 21020
rect 12548 20980 12549 21020
rect 12507 20971 12549 20980
rect 3627 20936 3669 20945
rect 3627 20896 3628 20936
rect 3668 20896 3669 20936
rect 3627 20887 3669 20896
rect 9675 20936 9717 20945
rect 9675 20896 9676 20936
rect 9716 20896 9717 20936
rect 9675 20887 9717 20896
rect 2187 20852 2229 20861
rect 3994 20852 4052 20853
rect 4971 20852 5013 20861
rect 2187 20812 2188 20852
rect 2228 20812 2229 20852
rect 2187 20803 2229 20812
rect 3435 20843 3477 20852
rect 3435 20803 3436 20843
rect 3476 20803 3477 20843
rect 3994 20812 4003 20852
rect 4043 20812 4052 20852
rect 3994 20811 4052 20812
rect 4491 20843 4533 20852
rect 3435 20794 3477 20803
rect 4491 20803 4492 20843
rect 4532 20803 4533 20843
rect 4971 20812 4972 20852
rect 5012 20812 5013 20852
rect 4971 20803 5013 20812
rect 5451 20852 5493 20861
rect 5451 20812 5452 20852
rect 5492 20812 5493 20852
rect 5451 20803 5493 20812
rect 5561 20852 5619 20853
rect 5561 20812 5570 20852
rect 5610 20812 5619 20852
rect 5561 20811 5619 20812
rect 5835 20852 5877 20861
rect 9291 20852 9333 20861
rect 5835 20812 5836 20852
rect 5876 20812 5877 20852
rect 5835 20803 5877 20812
rect 7083 20843 7125 20852
rect 7083 20803 7084 20843
rect 7124 20803 7125 20843
rect 9291 20812 9292 20852
rect 9332 20812 9333 20852
rect 9291 20803 9333 20812
rect 9562 20852 9620 20853
rect 11595 20852 11637 20861
rect 9562 20812 9571 20852
rect 9611 20812 9620 20852
rect 9562 20811 9620 20812
rect 10347 20843 10389 20852
rect 10347 20803 10348 20843
rect 10388 20803 10389 20843
rect 11595 20812 11596 20852
rect 11636 20812 11637 20852
rect 11595 20803 11637 20812
rect 4491 20794 4533 20803
rect 7083 20794 7125 20803
rect 10347 20794 10389 20803
rect 1227 20768 1269 20777
rect 1227 20728 1228 20768
rect 1268 20728 1269 20768
rect 1227 20719 1269 20728
rect 5067 20768 5109 20777
rect 5067 20728 5068 20768
rect 5108 20728 5109 20768
rect 5067 20719 5109 20728
rect 7947 20768 7989 20777
rect 7947 20728 7948 20768
rect 7988 20728 7989 20768
rect 7947 20719 7989 20728
rect 8379 20768 8421 20777
rect 8379 20728 8380 20768
rect 8420 20728 8421 20768
rect 8379 20719 8421 20728
rect 8619 20768 8661 20777
rect 8619 20728 8620 20768
rect 8660 20728 8661 20768
rect 8619 20719 8661 20728
rect 11883 20768 11925 20777
rect 11883 20728 11884 20768
rect 11924 20728 11925 20768
rect 11883 20719 11925 20728
rect 12267 20768 12309 20777
rect 12267 20728 12268 20768
rect 12308 20728 12309 20768
rect 12267 20719 12309 20728
rect 9963 20684 10005 20693
rect 9963 20644 9964 20684
rect 10004 20644 10005 20684
rect 9963 20635 10005 20644
rect 1467 20600 1509 20609
rect 1467 20560 1468 20600
rect 1508 20560 1509 20600
rect 1467 20551 1509 20560
rect 7707 20600 7749 20609
rect 7707 20560 7708 20600
rect 7748 20560 7749 20600
rect 7707 20551 7749 20560
rect 10155 20600 10197 20609
rect 10155 20560 10156 20600
rect 10196 20560 10197 20600
rect 10155 20551 10197 20560
rect 1152 20432 12576 20456
rect 1152 20392 3688 20432
rect 3728 20392 3770 20432
rect 3810 20392 3852 20432
rect 3892 20392 3934 20432
rect 3974 20392 4016 20432
rect 4056 20392 12576 20432
rect 1152 20368 12576 20392
rect 4107 20264 4149 20273
rect 4107 20224 4108 20264
rect 4148 20224 4149 20264
rect 4107 20215 4149 20224
rect 9387 20264 9429 20273
rect 9387 20224 9388 20264
rect 9428 20224 9429 20264
rect 9387 20215 9429 20224
rect 9819 20180 9861 20189
rect 9819 20140 9820 20180
rect 9860 20140 9861 20180
rect 9819 20131 9861 20140
rect 1227 20096 1269 20105
rect 1227 20056 1228 20096
rect 1268 20056 1269 20096
rect 1227 20047 1269 20056
rect 4587 20096 4629 20105
rect 4587 20056 4588 20096
rect 4628 20056 4629 20096
rect 4587 20047 4629 20056
rect 5547 20096 5589 20105
rect 5547 20056 5548 20096
rect 5588 20056 5589 20096
rect 5547 20047 5589 20056
rect 6987 20096 7029 20105
rect 6987 20056 6988 20096
rect 7028 20056 7029 20096
rect 6987 20047 7029 20056
rect 7227 20096 7269 20105
rect 7227 20056 7228 20096
rect 7268 20056 7269 20096
rect 7227 20047 7269 20056
rect 9579 20096 9621 20105
rect 9579 20056 9580 20096
rect 9620 20056 9621 20096
rect 9579 20047 9621 20056
rect 9915 20096 9957 20105
rect 9915 20056 9916 20096
rect 9956 20056 9957 20096
rect 9915 20047 9957 20056
rect 10155 20096 10197 20105
rect 10155 20056 10156 20096
rect 10196 20056 10197 20096
rect 10155 20047 10197 20056
rect 10923 20096 10965 20105
rect 10923 20056 10924 20096
rect 10964 20056 10965 20096
rect 10923 20047 10965 20056
rect 2667 20012 2709 20021
rect 2667 19972 2668 20012
rect 2708 19972 2709 20012
rect 2667 19963 2709 19972
rect 3907 20012 3965 20013
rect 3907 19972 3916 20012
rect 3956 19972 3965 20012
rect 3907 19971 3965 19972
rect 7947 20012 7989 20021
rect 7947 19972 7948 20012
rect 7988 19972 7989 20012
rect 7947 19963 7989 19972
rect 9187 20012 9245 20013
rect 9187 19972 9196 20012
rect 9236 19972 9245 20012
rect 9187 19971 9245 19972
rect 10426 20012 10484 20013
rect 10426 19972 10435 20012
rect 10475 19972 10484 20012
rect 10426 19971 10484 19972
rect 10539 20012 10581 20021
rect 10539 19972 10540 20012
rect 10580 19972 10581 20012
rect 10539 19963 10581 19972
rect 11019 20012 11061 20021
rect 11019 19972 11020 20012
rect 11060 19972 11061 20012
rect 11019 19963 11061 19972
rect 11491 20012 11549 20013
rect 11491 19972 11500 20012
rect 11540 19972 11549 20012
rect 11491 19971 11549 19972
rect 12010 20012 12068 20013
rect 12010 19972 12019 20012
rect 12059 19972 12068 20012
rect 12010 19971 12068 19972
rect 5307 19928 5349 19937
rect 5307 19888 5308 19928
rect 5348 19888 5349 19928
rect 5307 19879 5349 19888
rect 1467 19844 1509 19853
rect 1467 19804 1468 19844
rect 1508 19804 1509 19844
rect 1467 19795 1509 19804
rect 4827 19844 4869 19853
rect 4827 19804 4828 19844
rect 4868 19804 4869 19844
rect 4827 19795 4869 19804
rect 12171 19844 12213 19853
rect 12171 19804 12172 19844
rect 12212 19804 12213 19844
rect 12171 19795 12213 19804
rect 1152 19676 12576 19700
rect 1152 19636 4928 19676
rect 4968 19636 5010 19676
rect 5050 19636 5092 19676
rect 5132 19636 5174 19676
rect 5214 19636 5256 19676
rect 5296 19636 12576 19676
rect 1152 19612 12576 19636
rect 1467 19508 1509 19517
rect 1467 19468 1468 19508
rect 1508 19468 1509 19508
rect 1467 19459 1509 19468
rect 3627 19508 3669 19517
rect 3627 19468 3628 19508
rect 3668 19468 3669 19508
rect 3627 19459 3669 19468
rect 10587 19508 10629 19517
rect 10587 19468 10588 19508
rect 10628 19468 10629 19508
rect 10587 19459 10629 19468
rect 12171 19508 12213 19517
rect 12171 19468 12172 19508
rect 12212 19468 12213 19508
rect 12171 19459 12213 19468
rect 2187 19340 2229 19349
rect 6603 19340 6645 19349
rect 8235 19340 8277 19349
rect 10731 19340 10773 19349
rect 2187 19300 2188 19340
rect 2228 19300 2229 19340
rect 2187 19291 2229 19300
rect 3435 19331 3477 19340
rect 3435 19291 3436 19331
rect 3476 19291 3477 19331
rect 6603 19300 6604 19340
rect 6644 19300 6645 19340
rect 6603 19291 6645 19300
rect 7851 19331 7893 19340
rect 7851 19291 7852 19331
rect 7892 19291 7893 19331
rect 8235 19300 8236 19340
rect 8276 19300 8277 19340
rect 8235 19291 8277 19300
rect 9483 19331 9525 19340
rect 9483 19291 9484 19331
rect 9524 19291 9525 19331
rect 10731 19300 10732 19340
rect 10772 19300 10773 19340
rect 10731 19291 10773 19300
rect 11979 19331 12021 19340
rect 11979 19291 11980 19331
rect 12020 19291 12021 19331
rect 3435 19282 3477 19291
rect 7851 19282 7893 19291
rect 9483 19282 9525 19291
rect 11979 19282 12021 19291
rect 1227 19256 1269 19265
rect 1227 19216 1228 19256
rect 1268 19216 1269 19256
rect 1227 19207 1269 19216
rect 9963 19256 10005 19265
rect 9963 19216 9964 19256
rect 10004 19216 10005 19256
rect 9963 19207 10005 19216
rect 10347 19256 10389 19265
rect 10347 19216 10348 19256
rect 10388 19216 10389 19256
rect 10347 19207 10389 19216
rect 10203 19172 10245 19181
rect 10203 19132 10204 19172
rect 10244 19132 10245 19172
rect 10203 19123 10245 19132
rect 8043 19088 8085 19097
rect 8043 19048 8044 19088
rect 8084 19048 8085 19088
rect 8043 19039 8085 19048
rect 9675 19088 9717 19097
rect 9675 19048 9676 19088
rect 9716 19048 9717 19088
rect 9675 19039 9717 19048
rect 1152 18920 12576 18944
rect 1152 18880 3688 18920
rect 3728 18880 3770 18920
rect 3810 18880 3852 18920
rect 3892 18880 3934 18920
rect 3974 18880 4016 18920
rect 4056 18880 12576 18920
rect 1152 18856 12576 18880
rect 3387 18668 3429 18677
rect 3387 18628 3388 18668
rect 3428 18628 3429 18668
rect 3387 18619 3429 18628
rect 8859 18668 8901 18677
rect 8859 18628 8860 18668
rect 8900 18628 8901 18668
rect 8859 18619 8901 18628
rect 12507 18668 12549 18677
rect 12507 18628 12508 18668
rect 12548 18628 12549 18668
rect 12507 18619 12549 18628
rect 3147 18584 3189 18593
rect 3147 18544 3148 18584
rect 3188 18544 3189 18584
rect 3147 18535 3189 18544
rect 7179 18584 7221 18593
rect 7179 18544 7180 18584
rect 7220 18544 7221 18584
rect 7179 18535 7221 18544
rect 8458 18584 8516 18585
rect 8458 18544 8467 18584
rect 8507 18544 8516 18584
rect 8458 18543 8516 18544
rect 8619 18584 8661 18593
rect 8619 18544 8620 18584
rect 8660 18544 8661 18584
rect 8619 18535 8661 18544
rect 9771 18584 9813 18593
rect 9771 18544 9772 18584
rect 9812 18544 9813 18584
rect 9771 18535 9813 18544
rect 11403 18584 11445 18593
rect 11403 18544 11404 18584
rect 11444 18544 11445 18584
rect 11403 18535 11445 18544
rect 11883 18584 11925 18593
rect 11883 18544 11884 18584
rect 11924 18544 11925 18584
rect 11883 18535 11925 18544
rect 12123 18584 12165 18593
rect 12123 18544 12124 18584
rect 12164 18544 12165 18584
rect 12123 18535 12165 18544
rect 12267 18584 12309 18593
rect 12267 18544 12268 18584
rect 12308 18544 12309 18584
rect 12267 18535 12309 18544
rect 4011 18500 4053 18509
rect 4011 18460 4012 18500
rect 4052 18460 4053 18500
rect 4011 18451 4053 18460
rect 5251 18500 5309 18501
rect 5251 18460 5260 18500
rect 5300 18460 5309 18500
rect 5251 18459 5309 18460
rect 6682 18500 6740 18501
rect 6682 18460 6691 18500
rect 6731 18460 6740 18500
rect 6682 18459 6740 18460
rect 6795 18500 6837 18509
rect 6795 18460 6796 18500
rect 6836 18460 6837 18500
rect 6795 18451 6837 18460
rect 7275 18500 7317 18509
rect 7275 18460 7276 18500
rect 7316 18460 7317 18500
rect 7275 18451 7317 18460
rect 7747 18500 7805 18501
rect 7747 18460 7756 18500
rect 7796 18460 7805 18500
rect 7747 18459 7805 18460
rect 8235 18500 8293 18501
rect 8235 18460 8244 18500
rect 8284 18460 8293 18500
rect 8235 18459 8293 18460
rect 9274 18500 9332 18501
rect 9274 18460 9283 18500
rect 9323 18460 9332 18500
rect 9274 18459 9332 18460
rect 9387 18500 9429 18509
rect 9387 18460 9388 18500
rect 9428 18460 9429 18500
rect 9387 18451 9429 18460
rect 9867 18500 9909 18509
rect 9867 18460 9868 18500
rect 9908 18460 9909 18500
rect 9867 18451 9909 18460
rect 10339 18500 10397 18501
rect 10339 18460 10348 18500
rect 10388 18460 10397 18500
rect 10339 18459 10397 18460
rect 10858 18500 10916 18501
rect 10858 18460 10867 18500
rect 10907 18460 10916 18500
rect 10858 18459 10916 18460
rect 5451 18416 5493 18425
rect 5451 18376 5452 18416
rect 5492 18376 5493 18416
rect 5451 18367 5493 18376
rect 11019 18332 11061 18341
rect 11019 18292 11020 18332
rect 11060 18292 11061 18332
rect 11019 18283 11061 18292
rect 11643 18332 11685 18341
rect 11643 18292 11644 18332
rect 11684 18292 11685 18332
rect 11643 18283 11685 18292
rect 1152 18164 12576 18188
rect 1152 18124 4928 18164
rect 4968 18124 5010 18164
rect 5050 18124 5092 18164
rect 5132 18124 5174 18164
rect 5214 18124 5256 18164
rect 5296 18124 12576 18164
rect 1152 18100 12576 18124
rect 1467 17996 1509 18005
rect 1467 17956 1468 17996
rect 1508 17956 1509 17996
rect 1467 17947 1509 17956
rect 6027 17996 6069 18005
rect 6027 17956 6028 17996
rect 6068 17956 6069 17996
rect 6027 17947 6069 17956
rect 6795 17996 6837 18005
rect 6795 17956 6796 17996
rect 6836 17956 6837 17996
rect 6795 17947 6837 17956
rect 9099 17996 9141 18005
rect 9099 17956 9100 17996
rect 9140 17956 9141 17996
rect 9099 17947 9141 17956
rect 9915 17996 9957 18005
rect 9915 17956 9916 17996
rect 9956 17956 9957 17996
rect 9915 17947 9957 17956
rect 10299 17996 10341 18005
rect 10299 17956 10300 17996
rect 10340 17956 10341 17996
rect 10299 17947 10341 17956
rect 12267 17996 12309 18005
rect 12267 17956 12268 17996
rect 12308 17956 12309 17996
rect 12267 17947 12309 17956
rect 2331 17912 2373 17921
rect 2331 17872 2332 17912
rect 2372 17872 2373 17912
rect 2331 17863 2373 17872
rect 9243 17912 9285 17921
rect 9243 17872 9244 17912
rect 9284 17872 9285 17912
rect 9243 17863 9285 17872
rect 2475 17828 2517 17837
rect 5530 17828 5588 17829
rect 2475 17788 2476 17828
rect 2516 17788 2517 17828
rect 2475 17779 2517 17788
rect 3723 17819 3765 17828
rect 3723 17779 3724 17819
rect 3764 17779 3765 17819
rect 5530 17788 5539 17828
rect 5579 17788 5588 17828
rect 5530 17787 5588 17788
rect 6132 17828 6174 17837
rect 6132 17788 6133 17828
rect 6173 17788 6174 17828
rect 6507 17828 6549 17837
rect 6132 17779 6174 17788
rect 6363 17786 6405 17795
rect 3723 17770 3765 17779
rect 1227 17744 1269 17753
rect 1227 17704 1228 17744
rect 1268 17704 1269 17744
rect 1227 17695 1269 17704
rect 2091 17744 2133 17753
rect 2091 17704 2092 17744
rect 2132 17704 2133 17744
rect 2091 17695 2133 17704
rect 4107 17744 4149 17753
rect 4107 17704 4108 17744
rect 4148 17704 4149 17744
rect 4107 17695 4149 17704
rect 4779 17744 4821 17753
rect 4779 17704 4780 17744
rect 4820 17704 4821 17744
rect 4779 17695 4821 17704
rect 5019 17744 5061 17753
rect 5019 17704 5020 17744
rect 5060 17704 5061 17744
rect 5019 17695 5061 17704
rect 6242 17744 6284 17753
rect 6242 17704 6243 17744
rect 6283 17704 6284 17744
rect 6363 17746 6364 17786
rect 6404 17746 6405 17786
rect 6507 17788 6508 17828
rect 6548 17788 6549 17828
rect 6507 17779 6549 17788
rect 6641 17828 6699 17829
rect 6641 17788 6650 17828
rect 6690 17788 6699 17828
rect 6641 17787 6699 17788
rect 7659 17828 7701 17837
rect 10522 17828 10580 17829
rect 7659 17788 7660 17828
rect 7700 17788 7701 17828
rect 7659 17779 7701 17788
rect 8907 17819 8949 17828
rect 8907 17779 8908 17819
rect 8948 17779 8949 17819
rect 10522 17788 10531 17828
rect 10571 17788 10580 17828
rect 10522 17787 10580 17788
rect 10635 17828 10677 17837
rect 10635 17788 10636 17828
rect 10676 17788 10677 17828
rect 10635 17779 10677 17788
rect 11019 17828 11061 17837
rect 11019 17788 11020 17828
rect 11060 17788 11061 17828
rect 11019 17779 11061 17788
rect 11595 17819 11637 17828
rect 11595 17779 11596 17819
rect 11636 17779 11637 17819
rect 8907 17770 8949 17779
rect 11595 17770 11637 17779
rect 12075 17819 12117 17828
rect 12075 17779 12076 17819
rect 12116 17779 12117 17819
rect 12075 17770 12117 17779
rect 6363 17737 6405 17746
rect 9483 17744 9525 17753
rect 6242 17695 6284 17704
rect 9483 17704 9484 17744
rect 9524 17704 9525 17744
rect 9483 17695 9525 17704
rect 9675 17744 9717 17753
rect 9675 17704 9676 17744
rect 9716 17704 9717 17744
rect 9675 17695 9717 17704
rect 10059 17744 10101 17753
rect 10059 17704 10060 17744
rect 10100 17704 10101 17744
rect 10059 17695 10101 17704
rect 11115 17744 11157 17753
rect 11115 17704 11116 17744
rect 11156 17704 11157 17744
rect 11115 17695 11157 17704
rect 4347 17660 4389 17669
rect 4347 17620 4348 17660
rect 4388 17620 4389 17660
rect 4347 17611 4389 17620
rect 5510 17660 5552 17669
rect 5510 17620 5511 17660
rect 5551 17620 5552 17660
rect 5510 17611 5552 17620
rect 3915 17576 3957 17585
rect 3915 17536 3916 17576
rect 3956 17536 3957 17576
rect 3915 17527 3957 17536
rect 5722 17576 5780 17577
rect 5722 17536 5731 17576
rect 5771 17536 5780 17576
rect 5722 17535 5780 17536
rect 1152 17408 12576 17432
rect 1152 17368 3688 17408
rect 3728 17368 3770 17408
rect 3810 17368 3852 17408
rect 3892 17368 3934 17408
rect 3974 17368 4016 17408
rect 4056 17368 12576 17408
rect 1152 17344 12576 17368
rect 7467 17240 7509 17249
rect 7467 17200 7468 17240
rect 7508 17200 7509 17240
rect 7467 17191 7509 17200
rect 11835 17240 11877 17249
rect 11835 17200 11836 17240
rect 11876 17200 11877 17240
rect 11835 17191 11877 17200
rect 12507 17240 12549 17249
rect 12507 17200 12508 17240
rect 12548 17200 12549 17240
rect 12507 17191 12549 17200
rect 1467 17156 1509 17165
rect 1467 17116 1468 17156
rect 1508 17116 1509 17156
rect 1467 17107 1509 17116
rect 4587 17156 4629 17165
rect 4587 17116 4588 17156
rect 4628 17116 4629 17156
rect 4587 17107 4629 17116
rect 1227 17072 1269 17081
rect 1227 17032 1228 17072
rect 1268 17032 1269 17072
rect 1227 17023 1269 17032
rect 10443 17072 10485 17081
rect 10443 17032 10444 17072
rect 10484 17032 10485 17072
rect 6843 17021 6885 17030
rect 10443 17023 10485 17032
rect 12075 17072 12117 17081
rect 12075 17032 12076 17072
rect 12116 17032 12117 17072
rect 12075 17023 12117 17032
rect 12267 17072 12309 17081
rect 12267 17032 12268 17072
rect 12308 17032 12309 17072
rect 12267 17023 12309 17032
rect 5856 16999 5898 17008
rect 3147 16988 3189 16997
rect 3147 16948 3148 16988
rect 3188 16948 3189 16988
rect 3147 16939 3189 16948
rect 4387 16988 4445 16989
rect 4387 16948 4396 16988
rect 4436 16948 4445 16988
rect 4387 16947 4445 16948
rect 4858 16988 4916 16989
rect 4858 16948 4867 16988
rect 4907 16948 4916 16988
rect 4858 16947 4916 16948
rect 5164 16988 5206 16997
rect 5164 16948 5165 16988
rect 5205 16948 5206 16988
rect 5164 16939 5206 16948
rect 5331 16988 5389 16989
rect 5331 16948 5340 16988
rect 5380 16948 5389 16988
rect 5331 16947 5389 16948
rect 5493 16988 5551 16989
rect 5730 16988 5788 16989
rect 5493 16948 5502 16988
rect 5542 16948 5551 16988
rect 5493 16947 5551 16948
rect 5634 16979 5680 16988
rect 5634 16939 5635 16979
rect 5675 16939 5680 16979
rect 5730 16948 5739 16988
rect 5779 16948 5788 16988
rect 5856 16959 5857 16999
rect 5897 16959 5898 16999
rect 5856 16950 5898 16959
rect 6219 16988 6261 16997
rect 5730 16947 5788 16948
rect 6219 16948 6220 16988
rect 6260 16948 6261 16988
rect 6219 16939 6261 16948
rect 6338 16988 6380 16997
rect 6338 16948 6339 16988
rect 6379 16948 6380 16988
rect 6338 16939 6380 16948
rect 6448 16988 6506 16989
rect 6448 16948 6457 16988
rect 6497 16948 6506 16988
rect 6448 16947 6506 16948
rect 6699 16988 6741 16997
rect 6699 16948 6700 16988
rect 6740 16948 6741 16988
rect 6843 16981 6844 17021
rect 6884 16981 6885 17021
rect 6843 16972 6885 16981
rect 7162 16988 7220 16989
rect 6699 16939 6741 16948
rect 7162 16948 7171 16988
rect 7211 16948 7220 16988
rect 7162 16947 7220 16948
rect 7478 16988 7520 16997
rect 7478 16948 7479 16988
rect 7519 16948 7520 16988
rect 7478 16939 7520 16948
rect 7648 16988 7690 16997
rect 7648 16948 7649 16988
rect 7689 16948 7690 16988
rect 7648 16939 7690 16948
rect 7939 16988 7997 16989
rect 7939 16948 7948 16988
rect 7988 16948 7997 16988
rect 7939 16947 7997 16948
rect 8235 16988 8277 16997
rect 8235 16948 8236 16988
rect 8276 16948 8277 16988
rect 8235 16939 8277 16948
rect 9475 16988 9533 16989
rect 9475 16948 9484 16988
rect 9524 16948 9533 16988
rect 9475 16947 9533 16948
rect 9946 16988 10004 16989
rect 9946 16948 9955 16988
rect 9995 16948 10004 16988
rect 9946 16947 10004 16948
rect 10059 16988 10101 16997
rect 10059 16948 10060 16988
rect 10100 16948 10101 16988
rect 10059 16939 10101 16948
rect 10539 16988 10581 16997
rect 10539 16948 10540 16988
rect 10580 16948 10581 16988
rect 10539 16939 10581 16948
rect 11011 16988 11069 16989
rect 11011 16948 11020 16988
rect 11060 16948 11069 16988
rect 11011 16947 11069 16948
rect 11530 16988 11588 16989
rect 11530 16948 11539 16988
rect 11579 16948 11588 16988
rect 11530 16947 11588 16948
rect 5634 16930 5680 16939
rect 7851 16904 7893 16913
rect 7851 16864 7852 16904
rect 7892 16864 7893 16904
rect 7851 16855 7893 16864
rect 9675 16904 9717 16913
rect 9675 16864 9676 16904
rect 9716 16864 9717 16904
rect 9675 16855 9717 16864
rect 4587 16820 4629 16829
rect 4587 16780 4588 16820
rect 4628 16780 4629 16820
rect 4587 16771 4629 16780
rect 5067 16820 5109 16829
rect 5067 16780 5068 16820
rect 5108 16780 5109 16820
rect 5067 16771 5109 16780
rect 5818 16820 5876 16821
rect 5818 16780 5827 16820
rect 5867 16780 5876 16820
rect 5818 16779 5876 16780
rect 6123 16820 6165 16829
rect 6123 16780 6124 16820
rect 6164 16780 6165 16820
rect 6123 16771 6165 16780
rect 6987 16820 7029 16829
rect 6987 16780 6988 16820
rect 7028 16780 7029 16820
rect 6987 16771 7029 16780
rect 7258 16820 7316 16821
rect 7258 16780 7267 16820
rect 7307 16780 7316 16820
rect 7258 16779 7316 16780
rect 7738 16820 7796 16821
rect 7738 16780 7747 16820
rect 7787 16780 7796 16820
rect 7738 16779 7796 16780
rect 11691 16820 11733 16829
rect 11691 16780 11692 16820
rect 11732 16780 11733 16820
rect 11691 16771 11733 16780
rect 1152 16652 12576 16676
rect 1152 16612 4928 16652
rect 4968 16612 5010 16652
rect 5050 16612 5092 16652
rect 5132 16612 5174 16652
rect 5214 16612 5256 16652
rect 5296 16612 12576 16652
rect 1152 16588 12576 16612
rect 3339 16484 3381 16493
rect 3339 16444 3340 16484
rect 3380 16444 3381 16484
rect 3339 16435 3381 16444
rect 4971 16484 5013 16493
rect 4971 16444 4972 16484
rect 5012 16444 5013 16484
rect 4971 16435 5013 16444
rect 7275 16484 7317 16493
rect 7275 16444 7276 16484
rect 7316 16444 7317 16484
rect 7275 16435 7317 16444
rect 9723 16484 9765 16493
rect 9723 16444 9724 16484
rect 9764 16444 9765 16484
rect 9723 16435 9765 16444
rect 11403 16484 11445 16493
rect 11403 16444 11404 16484
rect 11444 16444 11445 16484
rect 11403 16435 11445 16444
rect 11835 16484 11877 16493
rect 11835 16444 11836 16484
rect 11876 16444 11877 16484
rect 11835 16435 11877 16444
rect 12507 16484 12549 16493
rect 12507 16444 12508 16484
rect 12548 16444 12549 16484
rect 12507 16435 12549 16444
rect 1467 16400 1509 16409
rect 1467 16360 1468 16400
rect 1508 16360 1509 16400
rect 1467 16351 1509 16360
rect 1899 16316 1941 16325
rect 3531 16316 3573 16325
rect 5530 16316 5588 16317
rect 1899 16276 1900 16316
rect 1940 16276 1941 16316
rect 1899 16267 1941 16276
rect 3147 16307 3189 16316
rect 3147 16267 3148 16307
rect 3188 16267 3189 16307
rect 3531 16276 3532 16316
rect 3572 16276 3573 16316
rect 3531 16267 3573 16276
rect 4779 16307 4821 16316
rect 4779 16267 4780 16307
rect 4820 16267 4821 16307
rect 5530 16276 5539 16316
rect 5579 16276 5588 16316
rect 5530 16275 5588 16276
rect 5643 16316 5685 16325
rect 5643 16276 5644 16316
rect 5684 16276 5685 16316
rect 5643 16267 5685 16276
rect 6027 16316 6069 16325
rect 7546 16316 7604 16317
rect 6027 16276 6028 16316
rect 6068 16276 6069 16316
rect 6027 16267 6069 16276
rect 6603 16307 6645 16316
rect 6603 16267 6604 16307
rect 6644 16267 6645 16307
rect 3147 16258 3189 16267
rect 4779 16258 4821 16267
rect 6603 16258 6645 16267
rect 7083 16307 7125 16316
rect 7083 16267 7084 16307
rect 7124 16267 7125 16307
rect 7546 16276 7555 16316
rect 7595 16276 7604 16316
rect 7546 16275 7604 16276
rect 7659 16316 7701 16325
rect 7659 16276 7660 16316
rect 7700 16276 7701 16316
rect 7659 16267 7701 16276
rect 8043 16316 8085 16325
rect 9963 16316 10005 16325
rect 8043 16276 8044 16316
rect 8084 16276 8085 16316
rect 8043 16267 8085 16276
rect 8619 16307 8661 16316
rect 8619 16267 8620 16307
rect 8660 16267 8661 16307
rect 7083 16258 7125 16267
rect 8619 16258 8661 16267
rect 9099 16307 9141 16316
rect 9099 16267 9100 16307
rect 9140 16267 9141 16307
rect 9963 16276 9964 16316
rect 10004 16276 10005 16316
rect 9963 16267 10005 16276
rect 11211 16307 11253 16316
rect 11211 16267 11212 16307
rect 11252 16267 11253 16307
rect 9099 16258 9141 16267
rect 11211 16258 11253 16267
rect 1227 16232 1269 16241
rect 1227 16192 1228 16232
rect 1268 16192 1269 16232
rect 1227 16183 1269 16192
rect 6123 16232 6165 16241
rect 6123 16192 6124 16232
rect 6164 16192 6165 16232
rect 6123 16183 6165 16192
rect 8139 16232 8181 16241
rect 8139 16192 8140 16232
rect 8180 16192 8181 16232
rect 8139 16183 8181 16192
rect 9322 16232 9380 16233
rect 9322 16192 9331 16232
rect 9371 16192 9380 16232
rect 9322 16191 9380 16192
rect 9483 16232 9525 16241
rect 9483 16192 9484 16232
rect 9524 16192 9525 16232
rect 9483 16183 9525 16192
rect 11595 16232 11637 16241
rect 11595 16192 11596 16232
rect 11636 16192 11637 16232
rect 11595 16183 11637 16192
rect 12267 16232 12309 16241
rect 12267 16192 12268 16232
rect 12308 16192 12309 16232
rect 12267 16183 12309 16192
rect 4971 16064 5013 16073
rect 4971 16024 4972 16064
rect 5012 16024 5013 16064
rect 4971 16015 5013 16024
rect 1152 15896 12576 15920
rect 1152 15856 3688 15896
rect 3728 15856 3770 15896
rect 3810 15856 3852 15896
rect 3892 15856 3934 15896
rect 3974 15856 4016 15896
rect 4056 15856 12576 15896
rect 1152 15832 12576 15856
rect 6154 15728 6212 15729
rect 6154 15688 6163 15728
rect 6203 15688 6212 15728
rect 6154 15687 6212 15688
rect 9003 15728 9045 15737
rect 9003 15688 9004 15728
rect 9044 15688 9045 15728
rect 9003 15679 9045 15688
rect 12267 15728 12309 15737
rect 12267 15688 12268 15728
rect 12308 15688 12309 15728
rect 12267 15679 12309 15688
rect 3915 15644 3957 15653
rect 3915 15604 3916 15644
rect 3956 15604 3957 15644
rect 3915 15595 3957 15604
rect 2091 15560 2133 15569
rect 2091 15520 2092 15560
rect 2132 15520 2133 15560
rect 2091 15511 2133 15520
rect 4875 15560 4917 15569
rect 4875 15520 4876 15560
rect 4916 15520 4917 15560
rect 4875 15511 4917 15520
rect 6891 15560 6933 15569
rect 6891 15520 6892 15560
rect 6932 15520 6933 15560
rect 6891 15511 6933 15520
rect 8410 15560 8468 15561
rect 8410 15520 8419 15560
rect 8459 15520 8468 15560
rect 8410 15519 8468 15520
rect 2475 15476 2517 15485
rect 2475 15436 2476 15476
rect 2516 15436 2517 15476
rect 2475 15427 2517 15436
rect 3715 15476 3773 15477
rect 3715 15436 3724 15476
rect 3764 15436 3773 15476
rect 3715 15435 3773 15436
rect 4378 15476 4436 15477
rect 4378 15436 4387 15476
rect 4427 15436 4436 15476
rect 4378 15435 4436 15436
rect 4491 15476 4533 15485
rect 4491 15436 4492 15476
rect 4532 15436 4533 15476
rect 4491 15427 4533 15436
rect 4971 15476 5013 15485
rect 4971 15436 4972 15476
rect 5012 15436 5013 15476
rect 4971 15427 5013 15436
rect 5443 15476 5501 15477
rect 5443 15436 5452 15476
rect 5492 15436 5501 15476
rect 5443 15435 5501 15436
rect 5931 15476 5989 15477
rect 5931 15436 5940 15476
rect 5980 15436 5989 15476
rect 5931 15435 5989 15436
rect 6394 15476 6452 15477
rect 6394 15436 6403 15476
rect 6443 15436 6452 15476
rect 6394 15435 6452 15436
rect 6507 15476 6549 15485
rect 6507 15436 6508 15476
rect 6548 15436 6549 15476
rect 6507 15427 6549 15436
rect 6987 15476 7029 15485
rect 6987 15436 6988 15476
rect 7028 15436 7029 15476
rect 6987 15427 7029 15436
rect 7459 15476 7517 15477
rect 7459 15436 7468 15476
rect 7508 15436 7517 15476
rect 7459 15435 7517 15436
rect 7947 15476 8005 15477
rect 7947 15436 7956 15476
rect 7996 15436 8005 15476
rect 7947 15435 8005 15436
rect 8278 15476 8320 15485
rect 8278 15436 8279 15476
rect 8319 15436 8320 15476
rect 8278 15427 8320 15436
rect 8523 15476 8565 15485
rect 8523 15436 8524 15476
rect 8564 15436 8565 15476
rect 8523 15427 8565 15436
rect 9187 15476 9245 15477
rect 9187 15436 9196 15476
rect 9236 15436 9245 15476
rect 9187 15435 9245 15436
rect 10443 15476 10485 15485
rect 10443 15436 10444 15476
rect 10484 15436 10485 15476
rect 10443 15427 10485 15436
rect 10827 15476 10869 15485
rect 10827 15436 10828 15476
rect 10868 15436 10869 15476
rect 10827 15427 10869 15436
rect 12067 15476 12125 15477
rect 12067 15436 12076 15476
rect 12116 15436 12125 15476
rect 12067 15435 12125 15436
rect 8602 15392 8660 15393
rect 8602 15352 8611 15392
rect 8651 15352 8660 15392
rect 8602 15351 8660 15352
rect 2331 15308 2373 15317
rect 2331 15268 2332 15308
rect 2372 15268 2373 15308
rect 2331 15259 2373 15268
rect 8139 15308 8181 15317
rect 8139 15268 8140 15308
rect 8180 15268 8181 15308
rect 8139 15259 8181 15268
rect 1152 15140 12576 15164
rect 1152 15100 4928 15140
rect 4968 15100 5010 15140
rect 5050 15100 5092 15140
rect 5132 15100 5174 15140
rect 5214 15100 5256 15140
rect 5296 15100 12576 15140
rect 1152 15076 12576 15100
rect 3610 14972 3668 14973
rect 3610 14932 3619 14972
rect 3659 14932 3668 14972
rect 3610 14931 3668 14932
rect 3723 14972 3765 14981
rect 3723 14932 3724 14972
rect 3764 14932 3765 14972
rect 3723 14923 3765 14932
rect 7947 14972 7989 14981
rect 7947 14932 7948 14972
rect 7988 14932 7989 14972
rect 7947 14923 7989 14932
rect 9483 14972 9525 14981
rect 9483 14932 9484 14972
rect 9524 14932 9525 14972
rect 9483 14923 9525 14932
rect 11355 14972 11397 14981
rect 11355 14932 11356 14972
rect 11396 14932 11397 14972
rect 11355 14923 11397 14932
rect 3833 14888 3875 14897
rect 3833 14848 3834 14888
rect 3874 14848 3875 14888
rect 3833 14839 3875 14848
rect 5259 14888 5301 14897
rect 5259 14848 5260 14888
rect 5300 14848 5301 14888
rect 5259 14839 5301 14848
rect 8427 14888 8469 14897
rect 8427 14848 8428 14888
rect 8468 14848 8469 14888
rect 8427 14839 8469 14848
rect 3130 14804 3188 14805
rect 3130 14764 3139 14804
rect 3179 14764 3188 14804
rect 3130 14763 3188 14764
rect 3514 14804 3572 14805
rect 3514 14764 3523 14804
rect 3563 14764 3572 14804
rect 3514 14763 3572 14764
rect 4027 14804 4085 14805
rect 4027 14764 4036 14804
rect 4076 14764 4085 14804
rect 4027 14763 4085 14764
rect 4186 14804 4244 14805
rect 4186 14764 4195 14804
rect 4235 14764 4244 14804
rect 4186 14763 4244 14764
rect 4330 14804 4388 14805
rect 4330 14764 4339 14804
rect 4379 14764 4388 14804
rect 4330 14763 4388 14764
rect 4474 14804 4532 14805
rect 4474 14764 4483 14804
rect 4523 14764 4532 14804
rect 4474 14763 4532 14764
rect 4576 14804 4634 14805
rect 4576 14764 4585 14804
rect 4625 14764 4634 14804
rect 4576 14763 4634 14764
rect 4875 14804 4917 14813
rect 4875 14764 4876 14804
rect 4916 14764 4917 14804
rect 4875 14755 4917 14764
rect 5146 14804 5204 14805
rect 5146 14764 5155 14804
rect 5195 14764 5204 14804
rect 5146 14763 5204 14764
rect 5739 14804 5781 14813
rect 5739 14764 5740 14804
rect 5780 14764 5781 14804
rect 5739 14755 5781 14764
rect 5931 14804 5973 14813
rect 5931 14764 5932 14804
rect 5972 14764 5973 14804
rect 5931 14755 5973 14764
rect 6202 14804 6260 14805
rect 6202 14764 6211 14804
rect 6251 14764 6260 14804
rect 6202 14763 6260 14764
rect 6315 14804 6357 14813
rect 6315 14764 6316 14804
rect 6356 14764 6357 14804
rect 6315 14755 6357 14764
rect 6699 14804 6741 14813
rect 8528 14804 8586 14805
rect 6699 14764 6700 14804
rect 6740 14764 6741 14804
rect 6699 14755 6741 14764
rect 7275 14795 7317 14804
rect 7275 14755 7276 14795
rect 7316 14755 7317 14795
rect 7275 14746 7317 14755
rect 7755 14795 7797 14804
rect 7755 14755 7756 14795
rect 7796 14755 7797 14795
rect 8528 14764 8537 14804
rect 8577 14764 8586 14804
rect 8528 14763 8586 14764
rect 8811 14804 8853 14813
rect 10923 14804 10965 14813
rect 8811 14764 8812 14804
rect 8852 14764 8853 14804
rect 8811 14755 8853 14764
rect 9675 14795 9717 14804
rect 9675 14755 9676 14795
rect 9716 14755 9717 14795
rect 10923 14764 10924 14804
rect 10964 14764 10965 14804
rect 10923 14755 10965 14764
rect 7755 14746 7797 14755
rect 9675 14746 9717 14755
rect 1419 14720 1461 14729
rect 1419 14680 1420 14720
rect 1460 14680 1461 14720
rect 1419 14671 1461 14680
rect 5835 14720 5877 14729
rect 5835 14680 5836 14720
rect 5876 14680 5877 14720
rect 5835 14671 5877 14680
rect 6795 14720 6837 14729
rect 6795 14680 6796 14720
rect 6836 14680 6837 14720
rect 6795 14671 6837 14680
rect 9291 14720 9333 14729
rect 9291 14680 9292 14720
rect 9332 14680 9333 14720
rect 9291 14671 9333 14680
rect 11115 14720 11157 14729
rect 11115 14680 11116 14720
rect 11156 14680 11157 14720
rect 11115 14671 11157 14680
rect 11691 14720 11733 14729
rect 11691 14680 11692 14720
rect 11732 14680 11733 14720
rect 11691 14671 11733 14680
rect 12075 14720 12117 14729
rect 12075 14680 12076 14720
rect 12116 14680 12117 14720
rect 12075 14671 12117 14680
rect 12459 14720 12501 14729
rect 12459 14680 12460 14720
rect 12500 14680 12501 14720
rect 12459 14671 12501 14680
rect 3110 14636 3152 14645
rect 3110 14596 3111 14636
rect 3151 14596 3152 14636
rect 3110 14587 3152 14596
rect 3322 14636 3380 14637
rect 3322 14596 3331 14636
rect 3371 14596 3380 14636
rect 3322 14595 3380 14596
rect 5547 14636 5589 14645
rect 5547 14596 5548 14636
rect 5588 14596 5589 14636
rect 5547 14587 5589 14596
rect 8139 14636 8181 14645
rect 8139 14596 8140 14636
rect 8180 14596 8181 14636
rect 8139 14587 8181 14596
rect 11451 14636 11493 14645
rect 11451 14596 11452 14636
rect 11492 14596 11493 14636
rect 11451 14587 11493 14596
rect 12219 14636 12261 14645
rect 12219 14596 12220 14636
rect 12260 14596 12261 14636
rect 12219 14587 12261 14596
rect 1179 14552 1221 14561
rect 1179 14512 1180 14552
rect 1220 14512 1221 14552
rect 1179 14503 1221 14512
rect 4587 14552 4629 14561
rect 4587 14512 4588 14552
rect 4628 14512 4629 14552
rect 4587 14503 4629 14512
rect 9051 14552 9093 14561
rect 9051 14512 9052 14552
rect 9092 14512 9093 14552
rect 9051 14503 9093 14512
rect 11835 14552 11877 14561
rect 11835 14512 11836 14552
rect 11876 14512 11877 14552
rect 11835 14503 11877 14512
rect 1152 14384 12576 14408
rect 1152 14344 3688 14384
rect 3728 14344 3770 14384
rect 3810 14344 3852 14384
rect 3892 14344 3934 14384
rect 3974 14344 4016 14384
rect 4056 14344 12576 14384
rect 1152 14320 12576 14344
rect 4875 14216 4917 14225
rect 4875 14176 4876 14216
rect 4916 14176 4917 14216
rect 4875 14167 4917 14176
rect 8667 14216 8709 14225
rect 8667 14176 8668 14216
rect 8708 14176 8709 14216
rect 8667 14167 8709 14176
rect 9051 14216 9093 14225
rect 9051 14176 9052 14216
rect 9092 14176 9093 14216
rect 9051 14167 9093 14176
rect 10491 14216 10533 14225
rect 10491 14176 10492 14216
rect 10532 14176 10533 14216
rect 10491 14167 10533 14176
rect 12075 14216 12117 14225
rect 12075 14176 12076 14216
rect 12116 14176 12117 14216
rect 12075 14167 12117 14176
rect 12219 14216 12261 14225
rect 12219 14176 12220 14216
rect 12260 14176 12261 14216
rect 12219 14167 12261 14176
rect 7563 14132 7605 14141
rect 7563 14092 7564 14132
rect 7604 14092 7605 14132
rect 7563 14083 7605 14092
rect 1419 14048 1461 14057
rect 1419 14008 1420 14048
rect 1460 14008 1461 14048
rect 1419 13999 1461 14008
rect 8907 14048 8949 14057
rect 8907 14008 8908 14048
rect 8948 14008 8949 14048
rect 7894 13997 7936 14006
rect 8907 13999 8949 14008
rect 9291 14048 9333 14057
rect 9291 14008 9292 14048
rect 9332 14008 9333 14048
rect 9291 13999 9333 14008
rect 9675 14048 9717 14057
rect 9675 14008 9676 14048
rect 9716 14008 9717 14048
rect 9675 13999 9717 14008
rect 10059 14048 10101 14057
rect 10059 14008 10060 14048
rect 10100 14008 10101 14048
rect 10059 13999 10101 14008
rect 10251 14048 10293 14057
rect 10251 14008 10252 14048
rect 10292 14008 10293 14048
rect 10251 13999 10293 14008
rect 12459 14048 12501 14057
rect 12459 14008 12460 14048
rect 12500 14008 12501 14048
rect 12459 13999 12501 14008
rect 3147 13964 3189 13973
rect 3147 13924 3148 13964
rect 3188 13924 3189 13964
rect 3147 13915 3189 13924
rect 4387 13964 4445 13965
rect 4387 13924 4396 13964
rect 4436 13924 4445 13964
rect 4387 13923 4445 13924
rect 5163 13964 5205 13973
rect 5547 13964 5589 13973
rect 5163 13924 5164 13964
rect 5204 13924 5205 13964
rect 5163 13915 5205 13924
rect 5259 13955 5301 13964
rect 5259 13915 5260 13955
rect 5300 13915 5301 13955
rect 5547 13924 5548 13964
rect 5588 13924 5589 13964
rect 5547 13915 5589 13924
rect 6070 13964 6112 13973
rect 6070 13924 6071 13964
rect 6111 13924 6112 13964
rect 6070 13915 6112 13924
rect 6202 13964 6260 13965
rect 6202 13924 6211 13964
rect 6251 13924 6260 13964
rect 6202 13923 6260 13924
rect 6315 13964 6357 13973
rect 6315 13924 6316 13964
rect 6356 13924 6357 13964
rect 6315 13915 6357 13924
rect 6891 13964 6933 13973
rect 6891 13924 6892 13964
rect 6932 13924 6933 13964
rect 6891 13915 6933 13924
rect 7138 13964 7196 13965
rect 7138 13924 7147 13964
rect 7187 13924 7196 13964
rect 7138 13923 7196 13924
rect 7258 13964 7316 13965
rect 7258 13924 7267 13964
rect 7307 13924 7316 13964
rect 7258 13923 7316 13924
rect 7755 13964 7797 13973
rect 7755 13924 7756 13964
rect 7796 13924 7797 13964
rect 7894 13957 7895 13997
rect 7935 13957 7936 13997
rect 7894 13948 7936 13957
rect 10635 13964 10677 13973
rect 7755 13915 7797 13924
rect 10635 13924 10636 13964
rect 10676 13924 10677 13964
rect 10635 13915 10677 13924
rect 11875 13964 11933 13965
rect 11875 13924 11884 13964
rect 11924 13924 11933 13964
rect 11875 13923 11933 13924
rect 5259 13906 5301 13915
rect 9435 13880 9477 13889
rect 9435 13840 9436 13880
rect 9476 13840 9477 13880
rect 9435 13831 9477 13840
rect 1179 13796 1221 13805
rect 1179 13756 1180 13796
rect 1220 13756 1221 13796
rect 1179 13747 1221 13756
rect 4587 13796 4629 13805
rect 4587 13756 4588 13796
rect 4628 13756 4629 13796
rect 4587 13747 4629 13756
rect 6394 13796 6452 13797
rect 6394 13756 6403 13796
rect 6443 13756 6452 13796
rect 6394 13755 6452 13756
rect 8043 13796 8085 13805
rect 8043 13756 8044 13796
rect 8084 13756 8085 13796
rect 8043 13747 8085 13756
rect 9819 13796 9861 13805
rect 9819 13756 9820 13796
rect 9860 13756 9861 13796
rect 9819 13747 9861 13756
rect 1152 13628 12576 13652
rect 1152 13588 4928 13628
rect 4968 13588 5010 13628
rect 5050 13588 5092 13628
rect 5132 13588 5174 13628
rect 5214 13588 5256 13628
rect 5296 13588 12576 13628
rect 1152 13564 12576 13588
rect 4395 13460 4437 13469
rect 4395 13420 4396 13460
rect 4436 13420 4437 13460
rect 4395 13411 4437 13420
rect 4666 13460 4724 13461
rect 4666 13420 4675 13460
rect 4715 13420 4724 13460
rect 4666 13419 4724 13420
rect 5259 13460 5301 13469
rect 5259 13420 5260 13460
rect 5300 13420 5301 13460
rect 5259 13411 5301 13420
rect 5547 13460 5589 13469
rect 5547 13420 5548 13460
rect 5588 13420 5589 13460
rect 5547 13411 5589 13420
rect 6394 13460 6452 13461
rect 6394 13420 6403 13460
rect 6443 13420 6452 13460
rect 6394 13419 6452 13420
rect 9723 13460 9765 13469
rect 9723 13420 9724 13460
rect 9764 13420 9765 13460
rect 9723 13411 9765 13420
rect 10107 13460 10149 13469
rect 10107 13420 10108 13460
rect 10148 13420 10149 13460
rect 10107 13411 10149 13420
rect 12219 13460 12261 13469
rect 12219 13420 12220 13460
rect 12260 13420 12261 13460
rect 12219 13411 12261 13420
rect 4573 13376 4615 13385
rect 4573 13336 4574 13376
rect 4614 13336 4615 13376
rect 4573 13327 4615 13336
rect 2955 13292 2997 13301
rect 4779 13292 4821 13301
rect 5050 13292 5108 13293
rect 2955 13252 2956 13292
rect 2996 13252 2997 13292
rect 2955 13243 2997 13252
rect 4203 13283 4245 13292
rect 4203 13243 4204 13283
rect 4244 13243 4245 13283
rect 4779 13252 4780 13292
rect 4820 13252 4821 13292
rect 4779 13243 4821 13252
rect 4875 13283 4917 13292
rect 4875 13243 4876 13283
rect 4916 13243 4917 13283
rect 5050 13252 5059 13292
rect 5099 13252 5108 13292
rect 5050 13251 5108 13252
rect 5355 13292 5397 13301
rect 5355 13252 5356 13292
rect 5396 13252 5397 13292
rect 5762 13292 5804 13301
rect 5355 13243 5397 13252
rect 5643 13250 5685 13259
rect 4203 13234 4245 13243
rect 4875 13234 4917 13243
rect 1419 13208 1461 13217
rect 1419 13168 1420 13208
rect 1460 13168 1461 13208
rect 5643 13210 5644 13250
rect 5684 13210 5685 13250
rect 5762 13252 5763 13292
rect 5803 13252 5804 13292
rect 5762 13243 5804 13252
rect 5872 13292 5930 13293
rect 5872 13252 5881 13292
rect 5921 13252 5930 13292
rect 5872 13251 5930 13252
rect 6070 13292 6112 13301
rect 6070 13252 6071 13292
rect 6111 13252 6112 13292
rect 6070 13243 6112 13252
rect 6315 13292 6357 13301
rect 6315 13252 6316 13292
rect 6356 13252 6357 13292
rect 6315 13243 6357 13252
rect 6742 13292 6784 13301
rect 6742 13252 6743 13292
rect 6783 13252 6784 13292
rect 6742 13243 6784 13252
rect 6987 13292 7029 13301
rect 9291 13292 9333 13301
rect 6987 13252 6988 13292
rect 7028 13252 7029 13292
rect 6987 13243 7029 13252
rect 8043 13283 8085 13292
rect 8043 13243 8044 13283
rect 8084 13243 8085 13283
rect 9291 13252 9292 13292
rect 9332 13252 9333 13292
rect 9291 13243 9333 13252
rect 10539 13292 10581 13301
rect 10539 13252 10540 13292
rect 10580 13252 10581 13292
rect 10539 13243 10581 13252
rect 11787 13283 11829 13292
rect 11787 13243 11788 13283
rect 11828 13243 11829 13283
rect 8043 13234 8085 13243
rect 11787 13234 11829 13243
rect 5643 13201 5685 13210
rect 6202 13208 6260 13209
rect 1419 13159 1461 13168
rect 6202 13168 6211 13208
rect 6251 13168 6260 13208
rect 6202 13167 6260 13168
rect 6874 13208 6932 13209
rect 6874 13168 6883 13208
rect 6923 13168 6932 13208
rect 6874 13167 6932 13168
rect 7083 13208 7125 13217
rect 7083 13168 7084 13208
rect 7124 13168 7125 13208
rect 7083 13159 7125 13168
rect 9483 13208 9525 13217
rect 9483 13168 9484 13208
rect 9524 13168 9525 13208
rect 9483 13159 9525 13168
rect 10347 13208 10389 13217
rect 10347 13168 10348 13208
rect 10388 13168 10389 13208
rect 10347 13159 10389 13168
rect 12459 13208 12501 13217
rect 12459 13168 12460 13208
rect 12500 13168 12501 13208
rect 12459 13159 12501 13168
rect 1179 13040 1221 13049
rect 1179 13000 1180 13040
rect 1220 13000 1221 13040
rect 1179 12991 1221 13000
rect 7851 13040 7893 13049
rect 7851 13000 7852 13040
rect 7892 13000 7893 13040
rect 7851 12991 7893 13000
rect 11979 13040 12021 13049
rect 11979 13000 11980 13040
rect 12020 13000 12021 13040
rect 11979 12991 12021 13000
rect 1152 12872 12576 12896
rect 1152 12832 3688 12872
rect 3728 12832 3770 12872
rect 3810 12832 3852 12872
rect 3892 12832 3934 12872
rect 3974 12832 4016 12872
rect 4056 12832 12576 12872
rect 1152 12808 12576 12832
rect 6027 12704 6069 12713
rect 6027 12664 6028 12704
rect 6068 12664 6069 12704
rect 6027 12655 6069 12664
rect 8859 12704 8901 12713
rect 8859 12664 8860 12704
rect 8900 12664 8901 12704
rect 8859 12655 8901 12664
rect 9531 12704 9573 12713
rect 9531 12664 9532 12704
rect 9572 12664 9573 12704
rect 9531 12655 9573 12664
rect 11835 12704 11877 12713
rect 11835 12664 11836 12704
rect 11876 12664 11877 12704
rect 11835 12655 11877 12664
rect 12219 12704 12261 12713
rect 12219 12664 12220 12704
rect 12260 12664 12261 12704
rect 12219 12655 12261 12664
rect 3819 12536 3861 12545
rect 3819 12496 3820 12536
rect 3860 12496 3861 12536
rect 3819 12487 3861 12496
rect 4971 12536 5013 12545
rect 4971 12496 4972 12536
rect 5012 12496 5013 12536
rect 7467 12536 7509 12545
rect 4971 12487 5013 12496
rect 5307 12494 5349 12503
rect 4107 12452 4149 12461
rect 4107 12412 4108 12452
rect 4148 12412 4149 12452
rect 4107 12403 4149 12412
rect 4354 12452 4412 12453
rect 4354 12412 4363 12452
rect 4403 12412 4412 12452
rect 4354 12411 4412 12412
rect 4474 12452 4532 12453
rect 4474 12412 4483 12452
rect 4523 12412 4532 12452
rect 4474 12411 4532 12412
rect 5067 12452 5109 12461
rect 5067 12412 5068 12452
rect 5108 12412 5109 12452
rect 5067 12403 5109 12412
rect 5186 12452 5228 12461
rect 5186 12412 5187 12452
rect 5227 12412 5228 12452
rect 5307 12454 5308 12494
rect 5348 12454 5349 12494
rect 7467 12496 7468 12536
rect 7508 12496 7509 12536
rect 7467 12487 7509 12496
rect 9099 12536 9141 12545
rect 9099 12496 9100 12536
rect 9140 12496 9141 12536
rect 9099 12487 9141 12496
rect 9291 12536 9333 12545
rect 9291 12496 9292 12536
rect 9332 12496 9333 12536
rect 9291 12487 9333 12496
rect 10251 12536 10293 12545
rect 10251 12496 10252 12536
rect 10292 12496 10293 12536
rect 10251 12487 10293 12496
rect 12075 12536 12117 12545
rect 12075 12496 12076 12536
rect 12116 12496 12117 12536
rect 12075 12487 12117 12496
rect 12459 12536 12501 12545
rect 12459 12496 12460 12536
rect 12500 12496 12501 12536
rect 12459 12487 12501 12496
rect 5307 12445 5349 12454
rect 5451 12452 5493 12461
rect 5186 12403 5228 12412
rect 5451 12412 5452 12452
rect 5492 12412 5493 12452
rect 5451 12403 5493 12412
rect 5585 12452 5643 12453
rect 5585 12412 5594 12452
rect 5634 12412 5643 12452
rect 5585 12411 5643 12412
rect 5931 12452 5973 12461
rect 5931 12412 5932 12452
rect 5972 12412 5973 12452
rect 5931 12403 5973 12412
rect 6123 12452 6165 12461
rect 6123 12412 6124 12452
rect 6164 12412 6165 12452
rect 6123 12403 6165 12412
rect 6970 12452 7028 12453
rect 6970 12412 6979 12452
rect 7019 12412 7028 12452
rect 6970 12411 7028 12412
rect 7083 12452 7125 12461
rect 7083 12412 7084 12452
rect 7124 12412 7125 12452
rect 7083 12403 7125 12412
rect 7563 12452 7605 12461
rect 7563 12412 7564 12452
rect 7604 12412 7605 12452
rect 7563 12403 7605 12412
rect 8035 12452 8093 12453
rect 8035 12412 8044 12452
rect 8084 12412 8093 12452
rect 8035 12411 8093 12412
rect 8523 12452 8581 12453
rect 8523 12412 8532 12452
rect 8572 12412 8581 12452
rect 8523 12411 8581 12412
rect 9754 12452 9812 12453
rect 9754 12412 9763 12452
rect 9803 12412 9812 12452
rect 9754 12411 9812 12412
rect 9867 12452 9909 12461
rect 9867 12412 9868 12452
rect 9908 12412 9909 12452
rect 9867 12403 9909 12412
rect 10347 12452 10389 12461
rect 10347 12412 10348 12452
rect 10388 12412 10389 12452
rect 10347 12403 10389 12412
rect 10819 12452 10877 12453
rect 10819 12412 10828 12452
rect 10868 12412 10877 12452
rect 10819 12411 10877 12412
rect 11338 12452 11396 12453
rect 11338 12412 11347 12452
rect 11387 12412 11396 12452
rect 11338 12411 11396 12412
rect 3579 12284 3621 12293
rect 3579 12244 3580 12284
rect 3620 12244 3621 12284
rect 3579 12235 3621 12244
rect 4827 12284 4869 12293
rect 4827 12244 4828 12284
rect 4868 12244 4869 12284
rect 4827 12235 4869 12244
rect 5739 12284 5781 12293
rect 5739 12244 5740 12284
rect 5780 12244 5781 12284
rect 5739 12235 5781 12244
rect 8715 12284 8757 12293
rect 8715 12244 8716 12284
rect 8756 12244 8757 12284
rect 8715 12235 8757 12244
rect 11499 12284 11541 12293
rect 11499 12244 11500 12284
rect 11540 12244 11541 12284
rect 11499 12235 11541 12244
rect 1152 12116 12576 12140
rect 1152 12076 4928 12116
rect 4968 12076 5010 12116
rect 5050 12076 5092 12116
rect 5132 12076 5174 12116
rect 5214 12076 5256 12116
rect 5296 12076 12576 12116
rect 1152 12052 12576 12076
rect 3195 11948 3237 11957
rect 3195 11908 3196 11948
rect 3236 11908 3237 11948
rect 3195 11899 3237 11908
rect 3867 11948 3909 11957
rect 3867 11908 3868 11948
rect 3908 11908 3909 11948
rect 3867 11899 3909 11908
rect 7995 11948 8037 11957
rect 7995 11908 7996 11948
rect 8036 11908 8037 11948
rect 7995 11899 8037 11908
rect 9099 11948 9141 11957
rect 9099 11908 9100 11948
rect 9140 11908 9141 11948
rect 9099 11899 9141 11908
rect 11355 11948 11397 11957
rect 11355 11908 11356 11948
rect 11396 11908 11397 11948
rect 11355 11899 11397 11908
rect 11835 11948 11877 11957
rect 11835 11908 11836 11948
rect 11876 11908 11877 11948
rect 11835 11899 11877 11908
rect 12219 11948 12261 11957
rect 12219 11908 12220 11948
rect 12260 11908 12261 11948
rect 12219 11899 12261 11908
rect 8091 11864 8133 11873
rect 8091 11824 8092 11864
rect 8132 11824 8133 11864
rect 8091 11815 8133 11824
rect 5818 11780 5876 11781
rect 5818 11740 5827 11780
rect 5867 11740 5876 11780
rect 5818 11739 5876 11740
rect 5931 11780 5973 11789
rect 5931 11740 5932 11780
rect 5972 11740 5973 11780
rect 5931 11731 5973 11740
rect 6315 11780 6357 11789
rect 9274 11780 9332 11781
rect 10251 11780 10293 11789
rect 6315 11740 6316 11780
rect 6356 11740 6357 11780
rect 6315 11731 6357 11740
rect 6891 11771 6933 11780
rect 6891 11731 6892 11771
rect 6932 11731 6933 11771
rect 6891 11722 6933 11731
rect 7371 11771 7413 11780
rect 7371 11731 7372 11771
rect 7412 11731 7413 11771
rect 9274 11740 9283 11780
rect 9323 11740 9332 11780
rect 9274 11739 9332 11740
rect 9771 11771 9813 11780
rect 7371 11722 7413 11731
rect 9771 11731 9772 11771
rect 9812 11731 9813 11771
rect 10251 11740 10252 11780
rect 10292 11740 10293 11780
rect 10251 11731 10293 11740
rect 10731 11780 10773 11789
rect 10731 11740 10732 11780
rect 10772 11740 10773 11780
rect 10731 11731 10773 11740
rect 10841 11780 10899 11781
rect 10841 11740 10850 11780
rect 10890 11740 10899 11780
rect 10841 11739 10899 11740
rect 9771 11722 9813 11731
rect 1419 11696 1461 11705
rect 1419 11656 1420 11696
rect 1460 11656 1461 11696
rect 1419 11647 1461 11656
rect 2955 11696 2997 11705
rect 2955 11656 2956 11696
rect 2996 11656 2997 11696
rect 2955 11647 2997 11656
rect 4107 11696 4149 11705
rect 4107 11656 4108 11696
rect 4148 11656 4149 11696
rect 4107 11647 4149 11656
rect 4299 11696 4341 11705
rect 4299 11656 4300 11696
rect 4340 11656 4341 11696
rect 4299 11647 4341 11656
rect 4683 11696 4725 11705
rect 4683 11656 4684 11696
rect 4724 11656 4725 11696
rect 4683 11647 4725 11656
rect 6411 11696 6453 11705
rect 6411 11656 6412 11696
rect 6452 11656 6453 11696
rect 6411 11647 6453 11656
rect 7594 11696 7652 11697
rect 7594 11656 7603 11696
rect 7643 11656 7652 11696
rect 7594 11655 7652 11656
rect 7755 11696 7797 11705
rect 7755 11656 7756 11696
rect 7796 11656 7797 11696
rect 7755 11647 7797 11656
rect 8331 11696 8373 11705
rect 8331 11656 8332 11696
rect 8372 11656 8373 11696
rect 8331 11647 8373 11656
rect 8715 11696 8757 11705
rect 8715 11656 8716 11696
rect 8756 11656 8757 11696
rect 8715 11647 8757 11656
rect 8955 11696 8997 11705
rect 8955 11656 8956 11696
rect 8996 11656 8997 11696
rect 8955 11647 8997 11656
rect 10347 11696 10389 11705
rect 10347 11656 10348 11696
rect 10388 11656 10389 11696
rect 10347 11647 10389 11656
rect 11115 11696 11157 11705
rect 11115 11656 11116 11696
rect 11156 11656 11157 11696
rect 11115 11647 11157 11656
rect 11691 11696 11733 11705
rect 11691 11656 11692 11696
rect 11732 11656 11733 11696
rect 11691 11647 11733 11656
rect 12075 11696 12117 11705
rect 12075 11656 12076 11696
rect 12116 11656 12117 11696
rect 12075 11647 12117 11656
rect 12459 11696 12501 11705
rect 12459 11656 12460 11696
rect 12500 11656 12501 11696
rect 12459 11647 12501 11656
rect 11451 11612 11493 11621
rect 11451 11572 11452 11612
rect 11492 11572 11493 11612
rect 11451 11563 11493 11572
rect 1179 11528 1221 11537
rect 1179 11488 1180 11528
rect 1220 11488 1221 11528
rect 1179 11479 1221 11488
rect 4539 11528 4581 11537
rect 4539 11488 4540 11528
rect 4580 11488 4581 11528
rect 4539 11479 4581 11488
rect 4923 11528 4965 11537
rect 4923 11488 4924 11528
rect 4964 11488 4965 11528
rect 4923 11479 4965 11488
rect 1152 11360 12576 11384
rect 1152 11320 3688 11360
rect 3728 11320 3770 11360
rect 3810 11320 3852 11360
rect 3892 11320 3934 11360
rect 3974 11320 4016 11360
rect 4056 11320 12576 11360
rect 1152 11296 12576 11320
rect 3915 11192 3957 11201
rect 3915 11152 3916 11192
rect 3956 11152 3957 11192
rect 3915 11143 3957 11152
rect 5115 11192 5157 11201
rect 5115 11152 5116 11192
rect 5156 11152 5157 11192
rect 5115 11143 5157 11152
rect 7611 11192 7653 11201
rect 7611 11152 7612 11192
rect 7652 11152 7653 11192
rect 7611 11143 7653 11152
rect 11595 11192 11637 11201
rect 11595 11152 11596 11192
rect 11636 11152 11637 11192
rect 11595 11143 11637 11152
rect 11835 11108 11877 11117
rect 11835 11068 11836 11108
rect 11876 11068 11877 11108
rect 11835 11059 11877 11068
rect 1419 11024 1461 11033
rect 1419 10984 1420 11024
rect 1460 10984 1461 11024
rect 5530 11024 5588 11025
rect 1419 10975 1461 10984
rect 5403 10982 5445 10991
rect 5530 10984 5539 11024
rect 5579 10984 5588 11024
rect 5530 10983 5588 10984
rect 6027 11024 6069 11033
rect 7371 11024 7413 11033
rect 6027 10984 6028 11024
rect 6068 10984 6069 11024
rect 2475 10940 2517 10949
rect 2475 10900 2476 10940
rect 2516 10900 2517 10940
rect 2475 10891 2517 10900
rect 3715 10940 3773 10941
rect 3715 10900 3724 10940
rect 3764 10900 3773 10940
rect 3715 10899 3773 10900
rect 5259 10940 5301 10949
rect 5259 10900 5260 10940
rect 5300 10900 5301 10940
rect 5403 10942 5404 10982
rect 5444 10942 5445 10982
rect 6027 10975 6069 10984
rect 6258 11015 6304 11024
rect 6258 10975 6259 11015
rect 6299 10975 6304 11015
rect 7371 10984 7372 11024
rect 7412 10984 7413 11024
rect 7371 10975 7413 10984
rect 7755 11024 7797 11033
rect 7755 10984 7756 11024
rect 7796 10984 7797 11024
rect 7755 10975 7797 10984
rect 8715 11024 8757 11033
rect 8715 10984 8716 11024
rect 8756 10984 8757 11024
rect 8715 10975 8757 10984
rect 12075 11024 12117 11033
rect 12075 10984 12076 11024
rect 12116 10984 12117 11024
rect 12075 10975 12117 10984
rect 12459 11024 12501 11033
rect 12459 10984 12460 11024
rect 12500 10984 12501 11024
rect 12459 10975 12501 10984
rect 6258 10966 6304 10975
rect 5403 10933 5445 10942
rect 5643 10940 5685 10949
rect 5259 10891 5301 10900
rect 5643 10900 5644 10940
rect 5684 10900 5685 10940
rect 5643 10891 5685 10900
rect 6123 10940 6165 10949
rect 6123 10900 6124 10940
rect 6164 10900 6165 10940
rect 6123 10891 6165 10900
rect 6352 10940 6410 10941
rect 6352 10900 6361 10940
rect 6401 10900 6410 10940
rect 6352 10899 6410 10900
rect 8218 10940 8276 10941
rect 8218 10900 8227 10940
rect 8267 10900 8276 10940
rect 8218 10899 8276 10900
rect 8331 10940 8373 10949
rect 8331 10900 8332 10940
rect 8372 10900 8373 10940
rect 8331 10891 8373 10900
rect 8811 10940 8853 10949
rect 8811 10900 8812 10940
rect 8852 10900 8853 10940
rect 8811 10891 8853 10900
rect 9283 10940 9341 10941
rect 9283 10900 9292 10940
rect 9332 10900 9341 10940
rect 9283 10899 9341 10900
rect 9771 10940 9829 10941
rect 9771 10900 9780 10940
rect 9820 10900 9829 10940
rect 9771 10899 9829 10900
rect 10155 10940 10197 10949
rect 10155 10900 10156 10940
rect 10196 10900 10197 10940
rect 10155 10891 10197 10900
rect 11395 10940 11453 10941
rect 11395 10900 11404 10940
rect 11444 10900 11453 10940
rect 11395 10899 11453 10900
rect 7995 10856 8037 10865
rect 7995 10816 7996 10856
rect 8036 10816 8037 10856
rect 7995 10807 8037 10816
rect 1179 10772 1221 10781
rect 1179 10732 1180 10772
rect 1220 10732 1221 10772
rect 1179 10723 1221 10732
rect 5722 10772 5780 10773
rect 5722 10732 5731 10772
rect 5771 10732 5780 10772
rect 5722 10731 5780 10732
rect 9963 10772 10005 10781
rect 9963 10732 9964 10772
rect 10004 10732 10005 10772
rect 9963 10723 10005 10732
rect 12219 10772 12261 10781
rect 12219 10732 12220 10772
rect 12260 10732 12261 10772
rect 12219 10723 12261 10732
rect 1152 10604 12576 10628
rect 1152 10564 4928 10604
rect 4968 10564 5010 10604
rect 5050 10564 5092 10604
rect 5132 10564 5174 10604
rect 5214 10564 5256 10604
rect 5296 10564 12576 10604
rect 1152 10540 12576 10564
rect 4107 10436 4149 10445
rect 4107 10396 4108 10436
rect 4148 10396 4149 10436
rect 4107 10387 4149 10396
rect 5739 10436 5781 10445
rect 5739 10396 5740 10436
rect 5780 10396 5781 10436
rect 5739 10387 5781 10396
rect 7755 10436 7797 10445
rect 7755 10396 7756 10436
rect 7796 10396 7797 10436
rect 7755 10387 7797 10396
rect 9867 10436 9909 10445
rect 9867 10396 9868 10436
rect 9908 10396 9909 10436
rect 9867 10387 9909 10396
rect 11835 10436 11877 10445
rect 11835 10396 11836 10436
rect 11876 10396 11877 10436
rect 11835 10387 11877 10396
rect 8043 10352 8085 10361
rect 8043 10312 8044 10352
rect 8084 10312 8085 10352
rect 8043 10303 8085 10312
rect 11451 10352 11493 10361
rect 11451 10312 11452 10352
rect 11492 10312 11493 10352
rect 11451 10303 11493 10312
rect 2667 10268 2709 10277
rect 4299 10268 4341 10277
rect 6010 10268 6068 10269
rect 2667 10228 2668 10268
rect 2708 10228 2709 10268
rect 2667 10219 2709 10228
rect 3915 10259 3957 10268
rect 3915 10219 3916 10259
rect 3956 10219 3957 10259
rect 4299 10228 4300 10268
rect 4340 10228 4341 10268
rect 4299 10219 4341 10228
rect 5547 10259 5589 10268
rect 5547 10219 5548 10259
rect 5588 10219 5589 10259
rect 6010 10228 6019 10268
rect 6059 10228 6068 10268
rect 6010 10227 6068 10228
rect 6128 10268 6170 10277
rect 6128 10228 6129 10268
rect 6169 10228 6170 10268
rect 6128 10219 6170 10228
rect 6507 10268 6549 10277
rect 9483 10268 9525 10277
rect 11307 10268 11349 10277
rect 6507 10228 6508 10268
rect 6548 10228 6549 10268
rect 6507 10219 6549 10228
rect 7083 10259 7125 10268
rect 7083 10219 7084 10259
rect 7124 10219 7125 10259
rect 3915 10210 3957 10219
rect 5547 10210 5589 10219
rect 7083 10210 7125 10219
rect 7563 10259 7605 10268
rect 7563 10219 7564 10259
rect 7604 10219 7605 10259
rect 7563 10210 7605 10219
rect 8235 10259 8277 10268
rect 8235 10219 8236 10259
rect 8276 10219 8277 10259
rect 9483 10228 9484 10268
rect 9524 10228 9525 10268
rect 9483 10219 9525 10228
rect 10059 10259 10101 10268
rect 10059 10219 10060 10259
rect 10100 10219 10101 10259
rect 11307 10228 11308 10268
rect 11348 10228 11349 10268
rect 11307 10219 11349 10228
rect 8235 10210 8277 10219
rect 10059 10210 10101 10219
rect 1419 10184 1461 10193
rect 1419 10144 1420 10184
rect 1460 10144 1461 10184
rect 1419 10135 1461 10144
rect 6603 10184 6645 10193
rect 6603 10144 6604 10184
rect 6644 10144 6645 10184
rect 6603 10135 6645 10144
rect 11691 10184 11733 10193
rect 11691 10144 11692 10184
rect 11732 10144 11733 10184
rect 11691 10135 11733 10144
rect 12075 10184 12117 10193
rect 12075 10144 12076 10184
rect 12116 10144 12117 10184
rect 12075 10135 12117 10144
rect 12459 10184 12501 10193
rect 12459 10144 12460 10184
rect 12500 10144 12501 10184
rect 12459 10135 12501 10144
rect 12219 10100 12261 10109
rect 12219 10060 12220 10100
rect 12260 10060 12261 10100
rect 12219 10051 12261 10060
rect 1179 10016 1221 10025
rect 1179 9976 1180 10016
rect 1220 9976 1221 10016
rect 1179 9967 1221 9976
rect 1152 9848 12576 9872
rect 1152 9808 3688 9848
rect 3728 9808 3770 9848
rect 3810 9808 3852 9848
rect 3892 9808 3934 9848
rect 3974 9808 4016 9848
rect 4056 9808 12576 9848
rect 1152 9784 12576 9808
rect 3003 9680 3045 9689
rect 3003 9640 3004 9680
rect 3044 9640 3045 9680
rect 3003 9631 3045 9640
rect 4971 9680 5013 9689
rect 4971 9640 4972 9680
rect 5012 9640 5013 9680
rect 4971 9631 5013 9640
rect 8091 9680 8133 9689
rect 8091 9640 8092 9680
rect 8132 9640 8133 9680
rect 8091 9631 8133 9640
rect 9771 9680 9813 9689
rect 9771 9640 9772 9680
rect 9812 9640 9813 9680
rect 9771 9631 9813 9640
rect 11835 9680 11877 9689
rect 11835 9640 11836 9680
rect 11876 9640 11877 9680
rect 11835 9631 11877 9640
rect 9963 9596 10005 9605
rect 9963 9556 9964 9596
rect 10004 9556 10005 9596
rect 9963 9547 10005 9556
rect 12219 9596 12261 9605
rect 12219 9556 12220 9596
rect 12260 9556 12261 9596
rect 12219 9547 12261 9556
rect 2763 9512 2805 9521
rect 2763 9472 2764 9512
rect 2804 9472 2805 9512
rect 2763 9463 2805 9472
rect 6123 9512 6165 9521
rect 6123 9472 6124 9512
rect 6164 9472 6165 9512
rect 6123 9463 6165 9472
rect 7851 9512 7893 9521
rect 7851 9472 7852 9512
rect 7892 9472 7893 9512
rect 7851 9463 7893 9472
rect 11595 9512 11637 9521
rect 11595 9472 11596 9512
rect 11636 9472 11637 9512
rect 11595 9463 11637 9472
rect 12459 9512 12501 9521
rect 12459 9472 12460 9512
rect 12500 9472 12501 9512
rect 12459 9463 12501 9472
rect 3531 9428 3573 9437
rect 3531 9388 3532 9428
rect 3572 9388 3573 9428
rect 3531 9379 3573 9388
rect 4771 9428 4829 9429
rect 4771 9388 4780 9428
rect 4820 9388 4829 9428
rect 4771 9387 4829 9388
rect 5163 9428 5205 9437
rect 5163 9388 5164 9428
rect 5204 9388 5205 9428
rect 5163 9379 5205 9388
rect 5355 9428 5397 9437
rect 5355 9388 5356 9428
rect 5396 9388 5397 9428
rect 5355 9379 5397 9388
rect 5626 9428 5684 9429
rect 5626 9388 5635 9428
rect 5675 9388 5684 9428
rect 5626 9387 5684 9388
rect 5739 9428 5781 9437
rect 5739 9388 5740 9428
rect 5780 9388 5781 9428
rect 5739 9379 5781 9388
rect 6219 9428 6261 9437
rect 6219 9388 6220 9428
rect 6260 9388 6261 9428
rect 6219 9379 6261 9388
rect 6691 9428 6749 9429
rect 6691 9388 6700 9428
rect 6740 9388 6749 9428
rect 6691 9387 6749 9388
rect 7210 9428 7268 9429
rect 7210 9388 7219 9428
rect 7259 9388 7268 9428
rect 7210 9387 7268 9388
rect 8331 9428 8373 9437
rect 8331 9388 8332 9428
rect 8372 9388 8373 9428
rect 8331 9379 8373 9388
rect 9571 9428 9629 9429
rect 9571 9388 9580 9428
rect 9620 9388 9629 9428
rect 9571 9387 9629 9388
rect 10147 9428 10205 9429
rect 10147 9388 10156 9428
rect 10196 9388 10205 9428
rect 10147 9387 10205 9388
rect 11403 9428 11445 9437
rect 11403 9388 11404 9428
rect 11444 9388 11445 9428
rect 11403 9379 11445 9388
rect 5338 9260 5396 9261
rect 5338 9220 5347 9260
rect 5387 9220 5396 9260
rect 5338 9219 5396 9220
rect 7371 9260 7413 9269
rect 7371 9220 7372 9260
rect 7412 9220 7413 9260
rect 7371 9211 7413 9220
rect 1152 9092 12576 9116
rect 1152 9052 4928 9092
rect 4968 9052 5010 9092
rect 5050 9052 5092 9092
rect 5132 9052 5174 9092
rect 5214 9052 5256 9092
rect 5296 9052 12576 9092
rect 1152 9028 12576 9052
rect 4491 8924 4533 8933
rect 4491 8884 4492 8924
rect 4532 8884 4533 8924
rect 4491 8875 4533 8884
rect 5547 8924 5589 8933
rect 5547 8884 5548 8924
rect 5588 8884 5589 8924
rect 5547 8875 5589 8884
rect 6298 8924 6356 8925
rect 6298 8884 6307 8924
rect 6347 8884 6356 8924
rect 6298 8883 6356 8884
rect 7066 8924 7124 8925
rect 7066 8884 7075 8924
rect 7115 8884 7124 8924
rect 7066 8883 7124 8884
rect 8907 8924 8949 8933
rect 8907 8884 8908 8924
rect 8948 8884 8949 8924
rect 8907 8875 8949 8884
rect 10299 8924 10341 8933
rect 10299 8884 10300 8924
rect 10340 8884 10341 8924
rect 10299 8875 10341 8884
rect 11067 8924 11109 8933
rect 11067 8884 11068 8924
rect 11108 8884 11109 8924
rect 11067 8875 11109 8884
rect 11451 8924 11493 8933
rect 11451 8884 11452 8924
rect 11492 8884 11493 8924
rect 11451 8875 11493 8884
rect 11835 8924 11877 8933
rect 11835 8884 11836 8924
rect 11876 8884 11877 8924
rect 11835 8875 11877 8884
rect 9339 8840 9381 8849
rect 9339 8800 9340 8840
rect 9380 8800 9381 8840
rect 9339 8791 9381 8800
rect 10683 8840 10725 8849
rect 10683 8800 10684 8840
rect 10724 8800 10725 8840
rect 10683 8791 10725 8800
rect 3051 8756 3093 8765
rect 4779 8756 4821 8765
rect 3051 8716 3052 8756
rect 3092 8716 3093 8756
rect 3051 8707 3093 8716
rect 4299 8747 4341 8756
rect 4299 8707 4300 8747
rect 4340 8707 4341 8747
rect 4779 8716 4780 8756
rect 4820 8716 4821 8756
rect 4779 8707 4821 8716
rect 4923 8756 4965 8765
rect 5739 8756 5781 8765
rect 4923 8716 4924 8756
rect 4964 8716 4965 8756
rect 4923 8707 4965 8716
rect 5163 8747 5205 8756
rect 5163 8707 5164 8747
rect 5204 8707 5205 8747
rect 5394 8747 5440 8756
rect 4299 8698 4341 8707
rect 5163 8698 5205 8707
rect 5262 8736 5304 8745
rect 5262 8696 5263 8736
rect 5303 8696 5304 8736
rect 5394 8707 5395 8747
rect 5435 8707 5440 8747
rect 5739 8716 5740 8756
rect 5780 8716 5781 8756
rect 5739 8707 5781 8716
rect 5979 8756 6021 8765
rect 6651 8756 6693 8765
rect 5979 8716 5980 8756
rect 6020 8716 6021 8756
rect 5866 8714 5924 8715
rect 5394 8698 5440 8707
rect 5262 8687 5304 8696
rect 1419 8672 1461 8681
rect 5866 8674 5875 8714
rect 5915 8674 5924 8714
rect 5979 8707 6021 8716
rect 6078 8747 6120 8756
rect 6078 8707 6079 8747
rect 6119 8707 6120 8747
rect 6078 8698 6120 8707
rect 6453 8742 6495 8751
rect 6453 8702 6454 8742
rect 6494 8702 6495 8742
rect 6651 8716 6652 8756
rect 6692 8716 6693 8756
rect 6651 8707 6693 8716
rect 6754 8756 6812 8757
rect 6754 8716 6763 8756
rect 6803 8716 6812 8756
rect 6754 8715 6812 8716
rect 6987 8756 7029 8765
rect 6987 8716 6988 8756
rect 7028 8716 7029 8756
rect 6987 8707 7029 8716
rect 7467 8756 7509 8765
rect 7467 8716 7468 8756
rect 7508 8716 7509 8756
rect 7467 8707 7509 8716
rect 8715 8747 8757 8756
rect 8715 8707 8716 8747
rect 8756 8707 8757 8747
rect 6453 8693 6495 8702
rect 8715 8698 8757 8707
rect 5866 8673 5924 8674
rect 1419 8632 1420 8672
rect 1460 8632 1461 8672
rect 1419 8623 1461 8632
rect 6874 8672 6932 8673
rect 6874 8632 6883 8672
rect 6923 8632 6932 8672
rect 6874 8631 6932 8632
rect 9099 8672 9141 8681
rect 9099 8632 9100 8672
rect 9140 8632 9141 8672
rect 9099 8623 9141 8632
rect 10539 8672 10581 8681
rect 10539 8632 10540 8672
rect 10580 8632 10581 8672
rect 10539 8623 10581 8632
rect 10923 8672 10965 8681
rect 10923 8632 10924 8672
rect 10964 8632 10965 8672
rect 10923 8623 10965 8632
rect 11307 8672 11349 8681
rect 11307 8632 11308 8672
rect 11348 8632 11349 8672
rect 11307 8623 11349 8632
rect 11691 8672 11733 8681
rect 11691 8632 11692 8672
rect 11732 8632 11733 8672
rect 11691 8623 11733 8632
rect 12075 8672 12117 8681
rect 12075 8632 12076 8672
rect 12116 8632 12117 8672
rect 12075 8623 12117 8632
rect 12459 8672 12501 8681
rect 12459 8632 12460 8672
rect 12500 8632 12501 8672
rect 12459 8623 12501 8632
rect 1179 8504 1221 8513
rect 1179 8464 1180 8504
rect 1220 8464 1221 8504
rect 1179 8455 1221 8464
rect 6027 8504 6069 8513
rect 6027 8464 6028 8504
rect 6068 8464 6069 8504
rect 6027 8455 6069 8464
rect 12219 8504 12261 8513
rect 12219 8464 12220 8504
rect 12260 8464 12261 8504
rect 12219 8455 12261 8464
rect 1152 8336 12576 8360
rect 1152 8296 3688 8336
rect 3728 8296 3770 8336
rect 3810 8296 3852 8336
rect 3892 8296 3934 8336
rect 3974 8296 4016 8336
rect 4056 8296 12576 8336
rect 1152 8272 12576 8296
rect 5547 8168 5589 8177
rect 5547 8128 5548 8168
rect 5588 8128 5589 8168
rect 5547 8119 5589 8128
rect 5835 8168 5877 8177
rect 5835 8128 5836 8168
rect 5876 8128 5877 8168
rect 5835 8119 5877 8128
rect 8571 8168 8613 8177
rect 8571 8128 8572 8168
rect 8612 8128 8613 8168
rect 8571 8119 8613 8128
rect 11067 8168 11109 8177
rect 11067 8128 11068 8168
rect 11108 8128 11109 8168
rect 11067 8119 11109 8128
rect 11451 8168 11493 8177
rect 11451 8128 11452 8168
rect 11492 8128 11493 8168
rect 11451 8119 11493 8128
rect 9675 8084 9717 8093
rect 9675 8044 9676 8084
rect 9716 8044 9717 8084
rect 9675 8035 9717 8044
rect 10107 8084 10149 8093
rect 10107 8044 10108 8084
rect 10148 8044 10149 8084
rect 10107 8035 10149 8044
rect 1419 8000 1461 8009
rect 1419 7960 1420 8000
rect 1460 7960 1461 8000
rect 1419 7951 1461 7960
rect 8331 8000 8373 8009
rect 8331 7960 8332 8000
rect 8372 7960 8373 8000
rect 5871 7958 5929 7959
rect 4107 7916 4149 7925
rect 4107 7876 4108 7916
rect 4148 7876 4149 7916
rect 4107 7867 4149 7876
rect 5347 7916 5405 7917
rect 5347 7876 5356 7916
rect 5396 7876 5405 7916
rect 5347 7875 5405 7876
rect 5739 7916 5781 7925
rect 5871 7918 5880 7958
rect 5920 7918 5929 7958
rect 8331 7951 8373 7960
rect 9867 8000 9909 8009
rect 9867 7960 9868 8000
rect 9908 7960 9909 8000
rect 9867 7951 9909 7960
rect 11307 8000 11349 8009
rect 11307 7960 11308 8000
rect 11348 7960 11349 8000
rect 11307 7951 11349 7960
rect 11691 8000 11733 8009
rect 11691 7960 11692 8000
rect 11732 7960 11733 8000
rect 11691 7951 11733 7960
rect 12075 8000 12117 8009
rect 12075 7960 12076 8000
rect 12116 7960 12117 8000
rect 12075 7951 12117 7960
rect 12219 8000 12261 8009
rect 12219 7960 12220 8000
rect 12260 7960 12261 8000
rect 12219 7951 12261 7960
rect 12459 8000 12501 8009
rect 12459 7960 12460 8000
rect 12500 7960 12501 8000
rect 12459 7951 12501 7960
rect 5871 7917 5929 7918
rect 5739 7876 5740 7916
rect 5780 7876 5781 7916
rect 5739 7867 5781 7876
rect 5980 7916 6038 7917
rect 5980 7876 5989 7916
rect 6029 7876 6038 7916
rect 5980 7875 6038 7876
rect 6699 7916 6741 7925
rect 6699 7876 6700 7916
rect 6740 7876 6741 7916
rect 6699 7867 6741 7876
rect 7939 7916 7997 7917
rect 7939 7876 7948 7916
rect 7988 7876 7997 7916
rect 7939 7875 7997 7876
rect 9003 7916 9045 7925
rect 9003 7876 9004 7916
rect 9044 7876 9045 7916
rect 9003 7867 9045 7876
rect 9274 7916 9332 7917
rect 9274 7876 9283 7916
rect 9323 7876 9332 7916
rect 9274 7875 9332 7876
rect 9387 7832 9429 7841
rect 9387 7792 9388 7832
rect 9428 7792 9429 7832
rect 9387 7783 9429 7792
rect 1179 7748 1221 7757
rect 1179 7708 1180 7748
rect 1220 7708 1221 7748
rect 1179 7699 1221 7708
rect 8139 7748 8181 7757
rect 8139 7708 8140 7748
rect 8180 7708 8181 7748
rect 8139 7699 8181 7708
rect 11835 7748 11877 7757
rect 11835 7708 11836 7748
rect 11876 7708 11877 7748
rect 11835 7699 11877 7708
rect 1152 7580 12576 7604
rect 1152 7540 4928 7580
rect 4968 7540 5010 7580
rect 5050 7540 5092 7580
rect 5132 7540 5174 7580
rect 5214 7540 5256 7580
rect 5296 7540 12576 7580
rect 1152 7516 12576 7540
rect 5434 7328 5492 7329
rect 5434 7288 5443 7328
rect 5483 7288 5492 7328
rect 5434 7287 5492 7288
rect 5110 7244 5152 7253
rect 5110 7204 5111 7244
rect 5151 7204 5152 7244
rect 5110 7195 5152 7204
rect 5242 7244 5300 7245
rect 5242 7204 5251 7244
rect 5291 7204 5300 7244
rect 5242 7203 5300 7204
rect 5355 7244 5397 7253
rect 5355 7204 5356 7244
rect 5396 7204 5397 7244
rect 5355 7195 5397 7204
rect 6795 7244 6837 7253
rect 6795 7204 6796 7244
rect 6836 7204 6837 7244
rect 6795 7195 6837 7204
rect 8043 7235 8085 7244
rect 8043 7195 8044 7235
rect 8084 7195 8085 7235
rect 8043 7186 8085 7195
rect 1419 7160 1461 7169
rect 1419 7120 1420 7160
rect 1460 7120 1461 7160
rect 1419 7111 1461 7120
rect 4683 7160 4725 7169
rect 4683 7120 4684 7160
rect 4724 7120 4725 7160
rect 4683 7111 4725 7120
rect 4923 7160 4965 7169
rect 4923 7120 4924 7160
rect 4964 7120 4965 7160
rect 4923 7111 4965 7120
rect 11307 7160 11349 7169
rect 11307 7120 11308 7160
rect 11348 7120 11349 7160
rect 11307 7111 11349 7120
rect 11691 7160 11733 7169
rect 11691 7120 11692 7160
rect 11732 7120 11733 7160
rect 11691 7111 11733 7120
rect 12075 7160 12117 7169
rect 12075 7120 12076 7160
rect 12116 7120 12117 7160
rect 12075 7111 12117 7120
rect 12219 7160 12261 7169
rect 12219 7120 12220 7160
rect 12260 7120 12261 7160
rect 12219 7111 12261 7120
rect 12459 7160 12501 7169
rect 12459 7120 12460 7160
rect 12500 7120 12501 7160
rect 12459 7111 12501 7120
rect 8235 7076 8277 7085
rect 8235 7036 8236 7076
rect 8276 7036 8277 7076
rect 8235 7027 8277 7036
rect 11451 7076 11493 7085
rect 11451 7036 11452 7076
rect 11492 7036 11493 7076
rect 11451 7027 11493 7036
rect 1179 6992 1221 7001
rect 1179 6952 1180 6992
rect 1220 6952 1221 6992
rect 1179 6943 1221 6952
rect 11067 6992 11109 7001
rect 11067 6952 11068 6992
rect 11108 6952 11109 6992
rect 11067 6943 11109 6952
rect 11835 6992 11877 7001
rect 11835 6952 11836 6992
rect 11876 6952 11877 6992
rect 11835 6943 11877 6952
rect 1152 6824 12576 6848
rect 1152 6784 3688 6824
rect 3728 6784 3770 6824
rect 3810 6784 3852 6824
rect 3892 6784 3934 6824
rect 3974 6784 4016 6824
rect 4056 6784 12576 6824
rect 1152 6760 12576 6784
rect 5163 6656 5205 6665
rect 5163 6616 5164 6656
rect 5204 6616 5205 6656
rect 5163 6607 5205 6616
rect 11835 6656 11877 6665
rect 11835 6616 11836 6656
rect 11876 6616 11877 6656
rect 11835 6607 11877 6616
rect 7371 6572 7413 6581
rect 7371 6532 7372 6572
rect 7412 6532 7413 6572
rect 7371 6523 7413 6532
rect 11691 6488 11733 6497
rect 11691 6448 11692 6488
rect 11732 6448 11733 6488
rect 11691 6439 11733 6448
rect 12075 6488 12117 6497
rect 12075 6448 12076 6488
rect 12116 6448 12117 6488
rect 12075 6439 12117 6448
rect 12459 6488 12501 6497
rect 12459 6448 12460 6488
rect 12500 6448 12501 6488
rect 12459 6439 12501 6448
rect 3723 6404 3765 6413
rect 3723 6364 3724 6404
rect 3764 6364 3765 6404
rect 3723 6355 3765 6364
rect 4963 6404 5021 6405
rect 4963 6364 4972 6404
rect 5012 6364 5021 6404
rect 4963 6363 5021 6364
rect 6699 6404 6741 6413
rect 6699 6364 6700 6404
rect 6740 6364 6741 6404
rect 6699 6355 6741 6364
rect 6970 6404 7028 6405
rect 6970 6364 6979 6404
rect 7019 6364 7028 6404
rect 6970 6363 7028 6364
rect 7563 6404 7605 6413
rect 7563 6364 7564 6404
rect 7604 6364 7605 6404
rect 7563 6355 7605 6364
rect 8803 6404 8861 6405
rect 8803 6364 8812 6404
rect 8852 6364 8861 6404
rect 8803 6363 8861 6364
rect 7083 6320 7125 6329
rect 7083 6280 7084 6320
rect 7124 6280 7125 6320
rect 7083 6271 7125 6280
rect 11451 6320 11493 6329
rect 11451 6280 11452 6320
rect 11492 6280 11493 6320
rect 11451 6271 11493 6280
rect 9003 6236 9045 6245
rect 9003 6196 9004 6236
rect 9044 6196 9045 6236
rect 9003 6187 9045 6196
rect 12219 6236 12261 6245
rect 12219 6196 12220 6236
rect 12260 6196 12261 6236
rect 12219 6187 12261 6196
rect 1152 6068 12576 6092
rect 1152 6028 4928 6068
rect 4968 6028 5010 6068
rect 5050 6028 5092 6068
rect 5132 6028 5174 6068
rect 5214 6028 5256 6068
rect 5296 6028 12576 6068
rect 1152 6004 12576 6028
rect 3051 5732 3093 5741
rect 4683 5732 4725 5741
rect 6315 5732 6357 5741
rect 8026 5732 8084 5733
rect 3051 5692 3052 5732
rect 3092 5692 3093 5732
rect 3051 5683 3093 5692
rect 4299 5723 4341 5732
rect 4299 5683 4300 5723
rect 4340 5683 4341 5723
rect 4683 5692 4684 5732
rect 4724 5692 4725 5732
rect 4683 5683 4725 5692
rect 5931 5723 5973 5732
rect 5931 5683 5932 5723
rect 5972 5683 5973 5723
rect 6315 5692 6316 5732
rect 6356 5692 6357 5732
rect 6315 5683 6357 5692
rect 7563 5723 7605 5732
rect 7563 5683 7564 5723
rect 7604 5683 7605 5723
rect 8026 5692 8035 5732
rect 8075 5692 8084 5732
rect 8026 5691 8084 5692
rect 8144 5732 8186 5741
rect 8144 5692 8145 5732
rect 8185 5692 8186 5732
rect 8144 5683 8186 5692
rect 8523 5732 8565 5741
rect 8523 5692 8524 5732
rect 8564 5692 8565 5732
rect 8523 5683 8565 5692
rect 9099 5723 9141 5732
rect 9099 5683 9100 5723
rect 9140 5683 9141 5723
rect 4299 5674 4341 5683
rect 5931 5674 5973 5683
rect 7563 5674 7605 5683
rect 9099 5674 9141 5683
rect 9579 5723 9621 5732
rect 9579 5683 9580 5723
rect 9620 5683 9621 5723
rect 9579 5674 9621 5683
rect 1419 5648 1461 5657
rect 1419 5608 1420 5648
rect 1460 5608 1461 5648
rect 1419 5599 1461 5608
rect 8619 5648 8661 5657
rect 8619 5608 8620 5648
rect 8660 5608 8661 5648
rect 8619 5599 8661 5608
rect 9802 5648 9860 5649
rect 9802 5608 9811 5648
rect 9851 5608 9860 5648
rect 9802 5607 9860 5608
rect 9963 5648 10005 5657
rect 9963 5608 9964 5648
rect 10004 5608 10005 5648
rect 9963 5599 10005 5608
rect 10203 5648 10245 5657
rect 10203 5608 10204 5648
rect 10244 5608 10245 5648
rect 10203 5599 10245 5608
rect 12075 5648 12117 5657
rect 12075 5608 12076 5648
rect 12116 5608 12117 5648
rect 12075 5599 12117 5608
rect 12219 5648 12261 5657
rect 12219 5608 12220 5648
rect 12260 5608 12261 5648
rect 12219 5599 12261 5608
rect 12459 5648 12501 5657
rect 12459 5608 12460 5648
rect 12500 5608 12501 5648
rect 12459 5599 12501 5608
rect 4491 5564 4533 5573
rect 4491 5524 4492 5564
rect 4532 5524 4533 5564
rect 4491 5515 4533 5524
rect 6123 5564 6165 5573
rect 6123 5524 6124 5564
rect 6164 5524 6165 5564
rect 6123 5515 6165 5524
rect 7755 5564 7797 5573
rect 7755 5524 7756 5564
rect 7796 5524 7797 5564
rect 7755 5515 7797 5524
rect 1179 5480 1221 5489
rect 1179 5440 1180 5480
rect 1220 5440 1221 5480
rect 1179 5431 1221 5440
rect 11835 5480 11877 5489
rect 11835 5440 11836 5480
rect 11876 5440 11877 5480
rect 11835 5431 11877 5440
rect 1152 5312 12576 5336
rect 1152 5272 3688 5312
rect 3728 5272 3770 5312
rect 3810 5272 3852 5312
rect 3892 5272 3934 5312
rect 3974 5272 4016 5312
rect 4056 5272 12576 5312
rect 1152 5248 12576 5272
rect 5355 5144 5397 5153
rect 5355 5104 5356 5144
rect 5396 5104 5397 5144
rect 5355 5095 5397 5104
rect 9819 5144 9861 5153
rect 9819 5104 9820 5144
rect 9860 5104 9861 5144
rect 9819 5095 9861 5104
rect 12219 5060 12261 5069
rect 12219 5020 12220 5060
rect 12260 5020 12261 5060
rect 12219 5011 12261 5020
rect 1227 4976 1269 4985
rect 1227 4936 1228 4976
rect 1268 4936 1269 4976
rect 1227 4927 1269 4936
rect 6123 4976 6165 4985
rect 6123 4936 6124 4976
rect 6164 4936 6165 4976
rect 6123 4927 6165 4936
rect 8139 4976 8181 4985
rect 8139 4936 8140 4976
rect 8180 4936 8181 4976
rect 8139 4927 8181 4936
rect 9579 4976 9621 4985
rect 9579 4936 9580 4976
rect 9620 4936 9621 4976
rect 9579 4927 9621 4936
rect 9915 4976 9957 4985
rect 9915 4936 9916 4976
rect 9956 4936 9957 4976
rect 9915 4927 9957 4936
rect 10155 4976 10197 4985
rect 10155 4936 10156 4976
rect 10196 4936 10197 4976
rect 10155 4927 10197 4936
rect 12075 4976 12117 4985
rect 12075 4936 12076 4976
rect 12116 4936 12117 4976
rect 12075 4927 12117 4936
rect 12459 4976 12501 4985
rect 12459 4936 12460 4976
rect 12500 4936 12501 4976
rect 12459 4927 12501 4936
rect 2283 4892 2325 4901
rect 2283 4852 2284 4892
rect 2324 4852 2325 4892
rect 2283 4843 2325 4852
rect 3523 4892 3581 4893
rect 3523 4852 3532 4892
rect 3572 4852 3581 4892
rect 3523 4851 3581 4852
rect 3915 4892 3957 4901
rect 3915 4852 3916 4892
rect 3956 4852 3957 4892
rect 3915 4843 3957 4852
rect 5155 4892 5213 4893
rect 5155 4852 5164 4892
rect 5204 4852 5213 4892
rect 5155 4851 5213 4852
rect 5626 4892 5684 4893
rect 5626 4852 5635 4892
rect 5675 4852 5684 4892
rect 5626 4851 5684 4852
rect 5739 4892 5781 4901
rect 5739 4852 5740 4892
rect 5780 4852 5781 4892
rect 5739 4843 5781 4852
rect 6219 4892 6261 4901
rect 6219 4852 6220 4892
rect 6260 4852 6261 4892
rect 6219 4843 6261 4852
rect 6691 4892 6749 4893
rect 6691 4852 6700 4892
rect 6740 4852 6749 4892
rect 6691 4851 6749 4852
rect 7179 4892 7237 4893
rect 7179 4852 7188 4892
rect 7228 4852 7237 4892
rect 7179 4851 7237 4852
rect 7642 4892 7700 4893
rect 7642 4852 7651 4892
rect 7691 4852 7700 4892
rect 7642 4851 7700 4852
rect 7755 4892 7797 4901
rect 7755 4852 7756 4892
rect 7796 4852 7797 4892
rect 7755 4843 7797 4852
rect 8235 4892 8277 4901
rect 8235 4852 8236 4892
rect 8276 4852 8277 4892
rect 8235 4843 8277 4852
rect 8707 4892 8765 4893
rect 8707 4852 8716 4892
rect 8756 4852 8765 4892
rect 8707 4851 8765 4852
rect 9195 4892 9253 4893
rect 9195 4852 9204 4892
rect 9244 4852 9253 4892
rect 9195 4851 9253 4852
rect 1467 4724 1509 4733
rect 1467 4684 1468 4724
rect 1508 4684 1509 4724
rect 1467 4675 1509 4684
rect 3723 4724 3765 4733
rect 3723 4684 3724 4724
rect 3764 4684 3765 4724
rect 3723 4675 3765 4684
rect 7371 4724 7413 4733
rect 7371 4684 7372 4724
rect 7412 4684 7413 4724
rect 7371 4675 7413 4684
rect 9387 4724 9429 4733
rect 9387 4684 9388 4724
rect 9428 4684 9429 4724
rect 9387 4675 9429 4684
rect 11835 4724 11877 4733
rect 11835 4684 11836 4724
rect 11876 4684 11877 4724
rect 11835 4675 11877 4684
rect 1152 4556 12576 4580
rect 1152 4516 4928 4556
rect 4968 4516 5010 4556
rect 5050 4516 5092 4556
rect 5132 4516 5174 4556
rect 5214 4516 5256 4556
rect 5296 4516 12576 4556
rect 1152 4492 12576 4516
rect 3387 4304 3429 4313
rect 3387 4264 3388 4304
rect 3428 4264 3429 4304
rect 3387 4255 3429 4264
rect 5355 4304 5397 4313
rect 5355 4264 5356 4304
rect 5396 4264 5397 4304
rect 5355 4255 5397 4264
rect 6987 4304 7029 4313
rect 6987 4264 6988 4304
rect 7028 4264 7029 4304
rect 6987 4255 7029 4264
rect 9195 4304 9237 4313
rect 9195 4264 9196 4304
rect 9236 4264 9237 4304
rect 9195 4255 9237 4264
rect 12219 4304 12261 4313
rect 12219 4264 12220 4304
rect 12260 4264 12261 4304
rect 12219 4255 12261 4264
rect 3915 4220 3957 4229
rect 5547 4220 5589 4229
rect 7258 4220 7316 4221
rect 3915 4180 3916 4220
rect 3956 4180 3957 4220
rect 3915 4171 3957 4180
rect 5163 4211 5205 4220
rect 5163 4171 5164 4211
rect 5204 4171 5205 4211
rect 5547 4180 5548 4220
rect 5588 4180 5589 4220
rect 5547 4171 5589 4180
rect 6795 4211 6837 4220
rect 6795 4171 6796 4211
rect 6836 4171 6837 4211
rect 7258 4180 7267 4220
rect 7307 4180 7316 4220
rect 7258 4179 7316 4180
rect 7371 4220 7413 4229
rect 7371 4180 7372 4220
rect 7412 4180 7413 4220
rect 7371 4171 7413 4180
rect 7755 4220 7797 4229
rect 10635 4220 10677 4229
rect 7755 4180 7756 4220
rect 7796 4180 7797 4220
rect 7755 4171 7797 4180
rect 8331 4211 8373 4220
rect 8331 4171 8332 4211
rect 8372 4171 8373 4211
rect 5163 4162 5205 4171
rect 6795 4162 6837 4171
rect 8331 4162 8373 4171
rect 8811 4211 8853 4220
rect 8811 4171 8812 4211
rect 8852 4171 8853 4211
rect 8811 4162 8853 4171
rect 9387 4211 9429 4220
rect 9387 4171 9388 4211
rect 9428 4171 9429 4211
rect 10635 4180 10636 4220
rect 10676 4180 10677 4220
rect 10635 4171 10677 4180
rect 9387 4162 9429 4171
rect 1419 4136 1461 4145
rect 1419 4096 1420 4136
rect 1460 4096 1461 4136
rect 1419 4087 1461 4096
rect 3147 4136 3189 4145
rect 3147 4096 3148 4136
rect 3188 4096 3189 4136
rect 3147 4087 3189 4096
rect 3531 4136 3573 4145
rect 3531 4096 3532 4136
rect 3572 4096 3573 4136
rect 3531 4087 3573 4096
rect 7851 4136 7893 4145
rect 7851 4096 7852 4136
rect 7892 4096 7893 4136
rect 7851 4087 7893 4096
rect 11691 4136 11733 4145
rect 11691 4096 11692 4136
rect 11732 4096 11733 4136
rect 11691 4087 11733 4096
rect 12075 4136 12117 4145
rect 12075 4096 12076 4136
rect 12116 4096 12117 4136
rect 12075 4087 12117 4096
rect 12459 4136 12501 4145
rect 12459 4096 12460 4136
rect 12500 4096 12501 4136
rect 12459 4087 12501 4096
rect 3771 4052 3813 4061
rect 3771 4012 3772 4052
rect 3812 4012 3813 4052
rect 3771 4003 3813 4012
rect 1179 3968 1221 3977
rect 1179 3928 1180 3968
rect 1220 3928 1221 3968
rect 1179 3919 1221 3928
rect 9034 3968 9092 3969
rect 9034 3928 9043 3968
rect 9083 3928 9092 3968
rect 9034 3927 9092 3928
rect 11451 3968 11493 3977
rect 11451 3928 11452 3968
rect 11492 3928 11493 3968
rect 11451 3919 11493 3928
rect 11835 3968 11877 3977
rect 11835 3928 11836 3968
rect 11876 3928 11877 3968
rect 11835 3919 11877 3928
rect 1152 3800 12576 3824
rect 1152 3760 3688 3800
rect 3728 3760 3770 3800
rect 3810 3760 3852 3800
rect 3892 3760 3934 3800
rect 3974 3760 4016 3800
rect 4056 3760 12576 3800
rect 1152 3736 12576 3760
rect 5547 3632 5589 3641
rect 5547 3592 5548 3632
rect 5588 3592 5589 3632
rect 5547 3583 5589 3592
rect 7179 3632 7221 3641
rect 7179 3592 7180 3632
rect 7220 3592 7221 3632
rect 7179 3583 7221 3592
rect 9099 3632 9141 3641
rect 9099 3592 9100 3632
rect 9140 3592 9141 3632
rect 9099 3583 9141 3592
rect 11835 3632 11877 3641
rect 11835 3592 11836 3632
rect 11876 3592 11877 3632
rect 11835 3583 11877 3592
rect 12219 3632 12261 3641
rect 12219 3592 12220 3632
rect 12260 3592 12261 3632
rect 12219 3583 12261 3592
rect 9627 3548 9669 3557
rect 9627 3508 9628 3548
rect 9668 3508 9669 3548
rect 9627 3499 9669 3508
rect 9243 3464 9285 3473
rect 9243 3424 9244 3464
rect 9284 3424 9285 3464
rect 9243 3415 9285 3424
rect 9483 3464 9525 3473
rect 9483 3424 9484 3464
rect 9524 3424 9525 3464
rect 9483 3415 9525 3424
rect 9867 3464 9909 3473
rect 9867 3424 9868 3464
rect 9908 3424 9909 3464
rect 9867 3415 9909 3424
rect 12075 3464 12117 3473
rect 12075 3424 12076 3464
rect 12116 3424 12117 3464
rect 12075 3415 12117 3424
rect 12459 3464 12501 3473
rect 12459 3424 12460 3464
rect 12500 3424 12501 3464
rect 12459 3415 12501 3424
rect 4107 3380 4149 3389
rect 4107 3340 4108 3380
rect 4148 3340 4149 3380
rect 4107 3331 4149 3340
rect 5347 3380 5405 3381
rect 5347 3340 5356 3380
rect 5396 3340 5405 3380
rect 5347 3339 5405 3340
rect 5739 3380 5781 3389
rect 5739 3340 5740 3380
rect 5780 3340 5781 3380
rect 5739 3331 5781 3340
rect 6979 3380 7037 3381
rect 6979 3340 6988 3380
rect 7028 3340 7037 3380
rect 6979 3339 7037 3340
rect 7659 3380 7701 3389
rect 7659 3340 7660 3380
rect 7700 3340 7701 3380
rect 7659 3331 7701 3340
rect 8899 3380 8957 3381
rect 8899 3340 8908 3380
rect 8948 3340 8957 3380
rect 8899 3339 8957 3340
rect 1152 3044 12576 3068
rect 1152 3004 4928 3044
rect 4968 3004 5010 3044
rect 5050 3004 5092 3044
rect 5132 3004 5174 3044
rect 5214 3004 5256 3044
rect 5296 3004 12576 3044
rect 1152 2980 12576 3004
rect 8187 2876 8229 2885
rect 8187 2836 8188 2876
rect 8228 2836 8229 2876
rect 8187 2827 8229 2836
rect 12219 2876 12261 2885
rect 12219 2836 12220 2876
rect 12260 2836 12261 2876
rect 12219 2827 12261 2836
rect 7227 2792 7269 2801
rect 7227 2752 7228 2792
rect 7268 2752 7269 2792
rect 7227 2743 7269 2752
rect 1419 2624 1461 2633
rect 1419 2584 1420 2624
rect 1460 2584 1461 2624
rect 1419 2575 1461 2584
rect 5163 2624 5205 2633
rect 5163 2584 5164 2624
rect 5204 2584 5205 2624
rect 5163 2575 5205 2584
rect 6987 2624 7029 2633
rect 6987 2584 6988 2624
rect 7028 2584 7029 2624
rect 6987 2575 7029 2584
rect 7947 2624 7989 2633
rect 7947 2584 7948 2624
rect 7988 2584 7989 2624
rect 7947 2575 7989 2584
rect 12459 2624 12501 2633
rect 12459 2584 12460 2624
rect 12500 2584 12501 2624
rect 12459 2575 12501 2584
rect 1179 2456 1221 2465
rect 1179 2416 1180 2456
rect 1220 2416 1221 2456
rect 1179 2407 1221 2416
rect 5403 2456 5445 2465
rect 5403 2416 5404 2456
rect 5444 2416 5445 2456
rect 5403 2407 5445 2416
rect 1152 2288 12576 2312
rect 1152 2248 3688 2288
rect 3728 2248 3770 2288
rect 3810 2248 3852 2288
rect 3892 2248 3934 2288
rect 3974 2248 4016 2288
rect 4056 2248 12576 2288
rect 1152 2224 12576 2248
rect 1467 2120 1509 2129
rect 1467 2080 1468 2120
rect 1508 2080 1509 2120
rect 1467 2071 1509 2080
rect 1227 1952 1269 1961
rect 1227 1912 1228 1952
rect 1268 1912 1269 1952
rect 1227 1903 1269 1912
rect 1152 1532 12576 1556
rect 1152 1492 4928 1532
rect 4968 1492 5010 1532
rect 5050 1492 5092 1532
rect 5132 1492 5174 1532
rect 5214 1492 5256 1532
rect 5296 1492 12576 1532
rect 1152 1468 12576 1492
<< via1 >>
rect 4928 46852 4968 46892
rect 5010 46852 5050 46892
rect 5092 46852 5132 46892
rect 5174 46852 5214 46892
rect 5256 46852 5296 46892
rect 1660 46684 1700 46724
rect 2236 46684 2276 46724
rect 2812 46684 2852 46724
rect 3388 46684 3428 46724
rect 3964 46684 4004 46724
rect 4540 46684 4580 46724
rect 5116 46684 5156 46724
rect 5692 46684 5732 46724
rect 6268 46684 6308 46724
rect 6844 46684 6884 46724
rect 7420 46684 7460 46724
rect 7996 46684 8036 46724
rect 8572 46684 8612 46724
rect 9148 46684 9188 46724
rect 9724 46684 9764 46724
rect 10300 46684 10340 46724
rect 10876 46684 10916 46724
rect 11452 46684 11492 46724
rect 1228 46432 1268 46472
rect 1900 46432 1940 46472
rect 2476 46432 2516 46472
rect 3052 46432 3092 46472
rect 3628 46432 3668 46472
rect 4204 46432 4244 46472
rect 4780 46432 4820 46472
rect 5356 46432 5396 46472
rect 5932 46432 5972 46472
rect 6508 46432 6548 46472
rect 7084 46432 7124 46472
rect 7660 46432 7700 46472
rect 8236 46432 8276 46472
rect 8812 46432 8852 46472
rect 9388 46432 9428 46472
rect 9964 46432 10004 46472
rect 10540 46432 10580 46472
rect 11116 46432 11156 46472
rect 11692 46432 11732 46472
rect 11884 46432 11924 46472
rect 12268 46432 12308 46472
rect 1468 46264 1508 46304
rect 12124 46264 12164 46304
rect 12508 46264 12548 46304
rect 3688 46096 3728 46136
rect 3770 46096 3810 46136
rect 3852 46096 3892 46136
rect 3934 46096 3974 46136
rect 4016 46096 4056 46136
rect 1564 45928 1604 45968
rect 10396 45928 10436 45968
rect 11260 45928 11300 45968
rect 10780 45844 10820 45884
rect 1228 45760 1268 45800
rect 1804 45760 1844 45800
rect 10156 45760 10196 45800
rect 10540 45760 10580 45800
rect 10924 45760 10964 45800
rect 11500 45760 11540 45800
rect 11884 45760 11924 45800
rect 12268 45760 12308 45800
rect 1468 45508 1508 45548
rect 11164 45508 11204 45548
rect 12124 45508 12164 45548
rect 12508 45508 12548 45548
rect 4928 45340 4968 45380
rect 5010 45340 5050 45380
rect 5092 45340 5132 45380
rect 5174 45340 5214 45380
rect 5256 45340 5296 45380
rect 5692 45172 5732 45212
rect 8668 45172 8708 45212
rect 10684 45172 10724 45212
rect 12028 45172 12068 45212
rect 4636 45088 4676 45128
rect 11644 45088 11684 45128
rect 1228 44920 1268 44960
rect 4396 44920 4436 44960
rect 5452 44920 5492 44960
rect 8908 44920 8948 44960
rect 10348 44920 10388 44960
rect 10924 44920 10964 44960
rect 11260 44920 11300 44960
rect 11500 44920 11540 44960
rect 11884 44920 11924 44960
rect 12268 44920 12308 44960
rect 10588 44836 10628 44876
rect 1468 44752 1508 44792
rect 3688 44584 3728 44624
rect 3770 44584 3810 44624
rect 3852 44584 3892 44624
rect 3934 44584 3974 44624
rect 4016 44584 4056 44624
rect 10492 44416 10532 44456
rect 10876 44416 10916 44456
rect 11644 44416 11684 44456
rect 11260 44332 11300 44372
rect 1228 44248 1268 44288
rect 10732 44248 10772 44288
rect 11116 44248 11156 44288
rect 11500 44248 11540 44288
rect 11884 44248 11924 44288
rect 12268 44248 12308 44288
rect 1468 43996 1508 44036
rect 12508 43996 12548 44036
rect 4928 43828 4968 43868
rect 5010 43828 5050 43868
rect 5092 43828 5132 43868
rect 5174 43828 5214 43868
rect 5256 43828 5296 43868
rect 8380 43660 8420 43700
rect 11356 43576 11396 43616
rect 1228 43408 1268 43448
rect 8620 43408 8660 43448
rect 11116 43408 11156 43448
rect 11500 43408 11540 43448
rect 11884 43408 11924 43448
rect 12268 43408 12308 43448
rect 1468 43240 1508 43280
rect 11740 43240 11780 43280
rect 12124 43240 12164 43280
rect 12508 43240 12548 43280
rect 3688 43072 3728 43112
rect 3770 43072 3810 43112
rect 3852 43072 3892 43112
rect 3934 43072 3974 43112
rect 4016 43072 4056 43112
rect 11260 42904 11300 42944
rect 11740 42904 11780 42944
rect 11356 42820 11396 42860
rect 11020 42736 11060 42776
rect 11596 42736 11636 42776
rect 11980 42736 12020 42776
rect 12268 42736 12308 42776
rect 12508 42484 12548 42524
rect 4928 42316 4968 42356
rect 5010 42316 5050 42356
rect 5092 42316 5132 42356
rect 5174 42316 5214 42356
rect 5256 42316 5296 42356
rect 1228 41896 1268 41936
rect 11884 41896 11924 41936
rect 12268 41896 12308 41936
rect 1468 41812 1508 41852
rect 12124 41728 12164 41768
rect 12508 41728 12548 41768
rect 3688 41560 3728 41600
rect 3770 41560 3810 41600
rect 3852 41560 3892 41600
rect 3934 41560 3974 41600
rect 4016 41560 4056 41600
rect 1228 41224 1268 41264
rect 11500 41224 11540 41264
rect 11884 41224 11924 41264
rect 12268 41224 12308 41264
rect 11740 41056 11780 41096
rect 1468 40972 1508 41012
rect 12124 40972 12164 41012
rect 12508 40972 12548 41012
rect 4928 40804 4968 40844
rect 5010 40804 5050 40844
rect 5092 40804 5132 40844
rect 5174 40804 5214 40844
rect 5256 40804 5296 40844
rect 1228 40384 1268 40424
rect 11500 40384 11540 40424
rect 11884 40384 11924 40424
rect 12268 40384 12308 40424
rect 1468 40300 1508 40340
rect 12508 40300 12548 40340
rect 11740 40216 11780 40256
rect 12124 40216 12164 40256
rect 3688 40048 3728 40088
rect 3770 40048 3810 40088
rect 3852 40048 3892 40088
rect 3934 40048 3974 40088
rect 4016 40048 4056 40088
rect 11116 39712 11156 39752
rect 11500 39712 11540 39752
rect 11884 39712 11924 39752
rect 12268 39712 12308 39752
rect 5932 39628 5972 39668
rect 7180 39628 7220 39668
rect 7564 39628 7604 39668
rect 8812 39628 8852 39668
rect 12124 39544 12164 39584
rect 7372 39460 7412 39500
rect 9004 39460 9044 39500
rect 11356 39460 11396 39500
rect 11740 39460 11780 39500
rect 12508 39460 12548 39500
rect 4928 39292 4968 39332
rect 5010 39292 5050 39332
rect 5092 39292 5132 39332
rect 5174 39292 5214 39332
rect 5256 39292 5296 39332
rect 4828 39124 4868 39164
rect 11356 39124 11396 39164
rect 4444 39040 4484 39080
rect 6412 39040 6452 39080
rect 8860 39040 8900 39080
rect 9244 39040 9284 39080
rect 10972 39040 11012 39080
rect 4972 38956 5012 38996
rect 6220 38947 6260 38987
rect 6691 38956 6731 38996
rect 6796 38956 6836 38996
rect 7180 38956 7220 38996
rect 7756 38947 7796 38987
rect 8236 38947 8276 38987
rect 1228 38872 1268 38912
rect 1468 38872 1508 38912
rect 4204 38872 4244 38912
rect 4588 38872 4628 38912
rect 7276 38872 7316 38912
rect 8467 38872 8507 38912
rect 8620 38872 8660 38912
rect 9004 38872 9044 38912
rect 9388 38872 9428 38912
rect 9628 38872 9668 38912
rect 10732 38872 10772 38912
rect 11116 38872 11156 38912
rect 11500 38872 11540 38912
rect 11884 38872 11924 38912
rect 12124 38872 12164 38912
rect 12268 38872 12308 38912
rect 12508 38872 12548 38912
rect 11740 38704 11780 38744
rect 3688 38536 3728 38576
rect 3770 38536 3810 38576
rect 3852 38536 3892 38576
rect 3934 38536 3974 38576
rect 4016 38536 4056 38576
rect 5260 38368 5300 38408
rect 6892 38284 6932 38324
rect 1228 38200 1268 38240
rect 7660 38200 7700 38240
rect 11020 38200 11060 38240
rect 11500 38200 11540 38240
rect 11884 38200 11924 38240
rect 12268 38200 12308 38240
rect 3820 38116 3860 38156
rect 5068 38116 5108 38156
rect 5452 38116 5492 38156
rect 6700 38116 6740 38156
rect 7171 38116 7211 38156
rect 7276 38116 7316 38156
rect 7756 38116 7796 38156
rect 8236 38116 8276 38156
rect 8716 38149 8756 38189
rect 9100 38116 9140 38156
rect 10348 38116 10388 38156
rect 12124 38032 12164 38072
rect 1468 37948 1508 37988
rect 8908 37948 8948 37988
rect 10540 37948 10580 37988
rect 11260 37948 11300 37988
rect 11740 37948 11780 37988
rect 12508 37948 12548 37988
rect 4928 37780 4968 37820
rect 5010 37780 5050 37820
rect 5092 37780 5132 37820
rect 5174 37780 5214 37820
rect 5256 37780 5296 37820
rect 8812 37612 8852 37652
rect 10924 37612 10964 37652
rect 3724 37444 3764 37484
rect 4972 37435 5012 37475
rect 5356 37444 5396 37484
rect 6604 37435 6644 37475
rect 7054 37444 7094 37484
rect 7180 37444 7220 37484
rect 7564 37444 7604 37484
rect 8140 37435 8180 37475
rect 8620 37435 8660 37475
rect 9187 37444 9227 37484
rect 9292 37444 9332 37484
rect 9676 37444 9716 37484
rect 10252 37435 10292 37475
rect 10732 37435 10772 37475
rect 1228 37360 1268 37400
rect 7660 37360 7700 37400
rect 9772 37360 9812 37400
rect 11308 37360 11348 37400
rect 11500 37360 11540 37400
rect 11884 37360 11924 37400
rect 12268 37360 12308 37400
rect 6796 37276 6836 37316
rect 12124 37276 12164 37316
rect 1468 37192 1508 37232
rect 5164 37192 5204 37232
rect 11068 37192 11108 37232
rect 11740 37192 11780 37232
rect 12508 37192 12548 37232
rect 3688 37024 3728 37064
rect 3770 37024 3810 37064
rect 3852 37024 3892 37064
rect 3934 37024 3974 37064
rect 4016 37024 4056 37064
rect 10492 36856 10532 36896
rect 9484 36688 9524 36728
rect 9868 36688 9908 36728
rect 10252 36688 10292 36728
rect 12268 36688 12308 36728
rect 3148 36604 3188 36644
rect 4396 36604 4436 36644
rect 4780 36604 4820 36644
rect 6028 36604 6068 36644
rect 6412 36604 6452 36644
rect 7660 36604 7700 36644
rect 10828 36604 10868 36644
rect 12076 36604 12116 36644
rect 10636 36520 10676 36560
rect 4588 36436 4628 36476
rect 6220 36436 6260 36476
rect 7852 36436 7892 36476
rect 9724 36436 9764 36476
rect 10108 36436 10148 36476
rect 12508 36436 12548 36476
rect 4928 36268 4968 36308
rect 5010 36268 5050 36308
rect 5092 36268 5132 36308
rect 5174 36268 5214 36308
rect 5256 36268 5296 36308
rect 6316 36100 6356 36140
rect 9964 36100 10004 36140
rect 4876 35932 4916 35972
rect 6124 35923 6164 35963
rect 10147 35932 10187 35972
rect 10636 35923 10676 35963
rect 11116 35932 11156 35972
rect 11596 35932 11636 35972
rect 11714 35932 11754 35972
rect 1228 35848 1268 35888
rect 4060 35848 4100 35888
rect 4300 35848 4340 35888
rect 4492 35848 4532 35888
rect 6508 35848 6548 35888
rect 9196 35848 9236 35888
rect 9580 35848 9620 35888
rect 11212 35848 11252 35888
rect 12268 35848 12308 35888
rect 4732 35764 4772 35804
rect 1468 35680 1508 35720
rect 6748 35680 6788 35720
rect 9436 35680 9476 35720
rect 9820 35680 9860 35720
rect 12508 35680 12548 35720
rect 3688 35512 3728 35552
rect 3770 35512 3810 35552
rect 3852 35512 3892 35552
rect 3934 35512 3974 35552
rect 4016 35512 4056 35552
rect 4156 35344 4196 35384
rect 12460 35344 12500 35384
rect 1228 35176 1268 35216
rect 3916 35176 3956 35216
rect 7564 35176 7604 35216
rect 8851 35176 8891 35216
rect 9004 35176 9044 35216
rect 4300 35092 4340 35132
rect 5548 35092 5588 35132
rect 7075 35092 7115 35132
rect 7180 35092 7220 35132
rect 7660 35092 7700 35132
rect 8140 35092 8180 35132
rect 8628 35092 8668 35132
rect 9580 35092 9620 35132
rect 10828 35092 10868 35132
rect 11020 35092 11060 35132
rect 12268 35092 12308 35132
rect 1468 34924 1508 34964
rect 5740 34924 5780 34964
rect 9244 34924 9284 34964
rect 9388 34924 9428 34964
rect 4928 34756 4968 34796
rect 5010 34756 5050 34796
rect 5092 34756 5132 34796
rect 5174 34756 5214 34796
rect 5256 34756 5296 34796
rect 9772 34504 9812 34544
rect 4492 34420 4532 34460
rect 5740 34411 5780 34451
rect 6124 34420 6164 34460
rect 7372 34411 7412 34451
rect 7843 34420 7883 34460
rect 7948 34420 7988 34460
rect 8332 34420 8372 34460
rect 8908 34411 8948 34451
rect 9388 34411 9428 34451
rect 9964 34411 10004 34451
rect 11212 34420 11252 34460
rect 1228 34336 1268 34376
rect 8428 34336 8468 34376
rect 11596 34336 11636 34376
rect 11884 34336 11924 34376
rect 12268 34336 12308 34376
rect 9628 34252 9668 34292
rect 12124 34252 12164 34292
rect 1468 34168 1508 34208
rect 5932 34168 5972 34208
rect 7564 34168 7604 34208
rect 11356 34168 11396 34208
rect 12508 34168 12548 34208
rect 3688 34000 3728 34040
rect 3770 34000 3810 34040
rect 3852 34000 3892 34040
rect 3934 34000 3974 34040
rect 4016 34000 4056 34040
rect 6556 33832 6596 33872
rect 11212 33748 11252 33788
rect 6316 33664 6356 33704
rect 7276 33664 7316 33704
rect 8563 33664 8603 33704
rect 8716 33664 8756 33704
rect 9196 33664 9236 33704
rect 11884 33664 11924 33704
rect 12268 33664 12308 33704
rect 3340 33580 3380 33620
rect 4588 33580 4628 33620
rect 6787 33580 6827 33620
rect 6892 33580 6932 33620
rect 7372 33580 7412 33620
rect 7852 33580 7892 33620
rect 8340 33580 8380 33620
rect 9580 33580 9620 33620
rect 10828 33580 10868 33620
rect 4780 33412 4820 33452
rect 8956 33412 8996 33452
rect 9436 33412 9476 33452
rect 11020 33412 11060 33452
rect 12124 33412 12164 33452
rect 12508 33412 12548 33452
rect 4928 33244 4968 33284
rect 5010 33244 5050 33284
rect 5092 33244 5132 33284
rect 5174 33244 5214 33284
rect 5256 33244 5296 33284
rect 6316 33076 6356 33116
rect 11404 33076 11444 33116
rect 6748 32992 6788 33032
rect 9388 32992 9428 33032
rect 4579 32908 4619 32948
rect 4684 32908 4724 32948
rect 5068 32908 5108 32948
rect 5644 32899 5684 32939
rect 6124 32899 6164 32939
rect 7948 32908 7988 32948
rect 9667 32908 9707 32948
rect 9772 32908 9812 32948
rect 1228 32824 1268 32864
rect 3724 32824 3764 32864
rect 4108 32824 4148 32864
rect 5164 32824 5204 32864
rect 6547 32824 6587 32864
rect 6892 32824 6932 32864
rect 9200 32866 9240 32906
rect 10252 32908 10292 32948
rect 10732 32899 10772 32939
rect 11212 32899 11252 32939
rect 7564 32824 7604 32864
rect 10156 32824 10196 32864
rect 11884 32824 11924 32864
rect 12268 32824 12308 32864
rect 3964 32740 4004 32780
rect 7804 32740 7844 32780
rect 1468 32656 1508 32696
rect 4348 32656 4388 32696
rect 7132 32656 7172 32696
rect 12124 32656 12164 32696
rect 12508 32656 12548 32696
rect 3688 32488 3728 32528
rect 3770 32488 3810 32528
rect 3852 32488 3892 32528
rect 3934 32488 3974 32528
rect 4016 32488 4056 32528
rect 9820 32320 9860 32360
rect 12460 32320 12500 32360
rect 1228 32152 1268 32192
rect 4876 32152 4916 32192
rect 6316 32152 6356 32192
rect 9580 32152 9620 32192
rect 2668 32068 2708 32108
rect 3916 32068 3956 32108
rect 4366 32068 4406 32108
rect 4492 32068 4532 32108
rect 4972 32068 5012 32108
rect 5452 32068 5492 32108
rect 5940 32068 5980 32108
rect 7948 32068 7988 32108
rect 9196 32068 9236 32108
rect 10531 32068 10571 32108
rect 10147 31984 10187 32024
rect 1468 31900 1508 31940
rect 4108 31900 4148 31940
rect 6124 31900 6164 31940
rect 6556 31900 6596 31940
rect 9388 31900 9428 31940
rect 12460 31900 12500 31940
rect 4928 31732 4968 31772
rect 5010 31732 5050 31772
rect 5092 31732 5132 31772
rect 5174 31732 5214 31772
rect 5256 31732 5296 31772
rect 4300 31564 4340 31604
rect 6316 31564 6356 31604
rect 6844 31564 6884 31604
rect 9244 31564 9284 31604
rect 2860 31396 2900 31436
rect 4108 31387 4148 31427
rect 4579 31396 4619 31436
rect 4684 31396 4724 31436
rect 5068 31396 5108 31436
rect 5644 31387 5684 31427
rect 6124 31387 6164 31427
rect 7564 31387 7604 31427
rect 8812 31396 8852 31436
rect 9580 31396 9620 31436
rect 10828 31387 10868 31427
rect 1228 31312 1268 31352
rect 5164 31312 5204 31352
rect 6700 31312 6740 31352
rect 7084 31312 7124 31352
rect 9004 31312 9044 31352
rect 11500 31312 11540 31352
rect 11884 31312 11924 31352
rect 12268 31312 12308 31352
rect 12124 31228 12164 31268
rect 1468 31144 1508 31184
rect 6460 31144 6500 31184
rect 7372 31144 7412 31184
rect 11020 31144 11060 31184
rect 11740 31144 11780 31184
rect 12508 31144 12548 31184
rect 3688 30976 3728 31016
rect 3770 30976 3810 31016
rect 3852 30976 3892 31016
rect 3934 30976 3974 31016
rect 4016 30976 4056 31016
rect 3676 30808 3716 30848
rect 8092 30808 8132 30848
rect 11644 30808 11684 30848
rect 10828 30724 10868 30764
rect 3436 30640 3476 30680
rect 6028 30640 6068 30680
rect 7315 30640 7355 30680
rect 7468 30640 7508 30680
rect 7852 30640 7892 30680
rect 8188 30640 8228 30680
rect 8428 30640 8468 30680
rect 10444 30640 10484 30680
rect 11020 30640 11060 30680
rect 11404 30640 11444 30680
rect 11884 30640 11924 30680
rect 12268 30640 12308 30680
rect 3820 30556 3860 30596
rect 5068 30556 5108 30596
rect 5539 30556 5579 30596
rect 5644 30556 5684 30596
rect 6124 30556 6164 30596
rect 6604 30556 6644 30596
rect 7123 30556 7163 30596
rect 8620 30556 8660 30596
rect 9868 30556 9908 30596
rect 5260 30472 5300 30512
rect 10060 30472 10100 30512
rect 12124 30472 12164 30512
rect 7708 30388 7748 30428
rect 10204 30388 10244 30428
rect 11260 30388 11300 30428
rect 12508 30388 12548 30428
rect 4928 30220 4968 30260
rect 5010 30220 5050 30260
rect 5092 30220 5132 30260
rect 5174 30220 5214 30260
rect 5256 30220 5296 30260
rect 7468 30052 7508 30092
rect 8284 30052 8324 30092
rect 7900 29968 7940 30008
rect 4078 29884 4118 29924
rect 4204 29884 4244 29924
rect 4588 29884 4628 29924
rect 5164 29875 5204 29915
rect 5644 29875 5684 29915
rect 6028 29884 6068 29924
rect 7276 29875 7316 29915
rect 10156 29884 10196 29924
rect 10531 29884 10571 29924
rect 1228 29800 1268 29840
rect 4684 29800 4724 29840
rect 7660 29800 7700 29840
rect 8044 29800 8084 29840
rect 9388 29800 9428 29840
rect 9772 29800 9812 29840
rect 10012 29800 10052 29840
rect 9628 29716 9668 29756
rect 1468 29632 1508 29672
rect 5875 29632 5915 29672
rect 12460 29632 12500 29672
rect 3688 29464 3728 29504
rect 3770 29464 3810 29504
rect 3852 29464 3892 29504
rect 3934 29464 3974 29504
rect 4016 29464 4056 29504
rect 1468 29296 1508 29336
rect 2620 29296 2660 29336
rect 4588 29296 4628 29336
rect 5980 29296 6020 29336
rect 5596 29212 5636 29252
rect 1228 29128 1268 29168
rect 2380 29128 2420 29168
rect 5356 29128 5396 29168
rect 5740 29128 5780 29168
rect 10348 29128 10388 29168
rect 11884 29128 11924 29168
rect 12268 29128 12308 29168
rect 3148 29044 3188 29084
rect 4396 29044 4436 29084
rect 6412 29044 6452 29084
rect 7660 29044 7700 29084
rect 8044 29044 8084 29084
rect 9292 29044 9332 29084
rect 9859 29044 9899 29084
rect 9964 29044 10004 29084
rect 10444 29044 10484 29084
rect 10923 29044 10963 29084
rect 11412 29044 11452 29084
rect 7852 28876 7892 28916
rect 9484 28876 9524 28916
rect 11596 28876 11636 28916
rect 12124 28876 12164 28916
rect 12508 28876 12548 28916
rect 4928 28708 4968 28748
rect 5010 28708 5050 28748
rect 5092 28708 5132 28748
rect 5174 28708 5214 28748
rect 5256 28708 5296 28748
rect 1468 28540 1508 28580
rect 4012 28540 4052 28580
rect 10348 28540 10388 28580
rect 2572 28372 2612 28412
rect 3820 28363 3860 28403
rect 6892 28372 6932 28412
rect 8140 28363 8180 28403
rect 8611 28372 8651 28412
rect 8716 28372 8756 28412
rect 9100 28372 9140 28412
rect 9676 28363 9716 28403
rect 10156 28363 10196 28403
rect 10540 28372 10580 28412
rect 11788 28363 11828 28403
rect 1228 28288 1268 28328
rect 9196 28288 9236 28328
rect 12364 28288 12404 28328
rect 8332 28120 8372 28160
rect 11980 28120 12020 28160
rect 12124 28120 12164 28160
rect 3688 27952 3728 27992
rect 3770 27952 3810 27992
rect 3852 27952 3892 27992
rect 3934 27952 3974 27992
rect 4016 27952 4056 27992
rect 10579 27784 10619 27824
rect 9292 27616 9332 27656
rect 4300 27532 4340 27572
rect 5548 27532 5588 27572
rect 6796 27532 6836 27572
rect 8044 27532 8084 27572
rect 8803 27532 8843 27572
rect 8908 27532 8948 27572
rect 9388 27532 9428 27572
rect 9868 27532 9908 27572
rect 10356 27532 10396 27572
rect 10924 27532 10964 27572
rect 12172 27532 12212 27572
rect 8236 27448 8276 27488
rect 5740 27364 5780 27404
rect 10732 27364 10772 27404
rect 4928 27196 4968 27236
rect 5010 27196 5050 27236
rect 5092 27196 5132 27236
rect 5174 27196 5214 27236
rect 5256 27196 5296 27236
rect 1468 27028 1508 27068
rect 6556 27028 6596 27068
rect 12028 27028 12068 27068
rect 4108 26944 4148 26984
rect 2668 26860 2708 26900
rect 3916 26851 3956 26891
rect 4387 26860 4427 26900
rect 4492 26860 4532 26900
rect 4876 26860 4916 26900
rect 5452 26851 5492 26891
rect 5932 26851 5972 26891
rect 7223 26860 7263 26900
rect 7468 26860 7508 26900
rect 9763 26860 9803 26900
rect 9868 26860 9908 26900
rect 10252 26860 10292 26900
rect 10828 26851 10868 26891
rect 11308 26851 11348 26891
rect 1228 26776 1268 26816
rect 4972 26776 5012 26816
rect 6163 26776 6203 26816
rect 6316 26776 6356 26816
rect 7363 26776 7403 26816
rect 7564 26776 7604 26816
rect 10348 26776 10388 26816
rect 11692 26776 11732 26816
rect 12268 26776 12308 26816
rect 11539 26608 11579 26648
rect 11932 26608 11972 26648
rect 3688 26440 3728 26480
rect 3770 26440 3810 26480
rect 3852 26440 3892 26480
rect 3934 26440 3974 26480
rect 4016 26440 4056 26480
rect 4732 26272 4772 26312
rect 11731 26272 11771 26312
rect 6700 26188 6740 26228
rect 4492 26104 4532 26144
rect 10444 26104 10484 26144
rect 12076 26104 12116 26144
rect 12268 26104 12308 26144
rect 1420 26020 1460 26060
rect 2668 26020 2708 26060
rect 3052 26020 3092 26060
rect 4300 26020 4340 26060
rect 5260 26020 5300 26060
rect 6508 26020 6548 26060
rect 6892 26020 6932 26060
rect 8140 26020 8180 26060
rect 8524 26020 8564 26060
rect 8663 26053 8703 26093
rect 9955 26020 9995 26060
rect 10060 26020 10100 26060
rect 10540 26020 10580 26060
rect 11015 26020 11055 26060
rect 11539 26020 11579 26060
rect 1228 25936 1268 25976
rect 8332 25936 8372 25976
rect 11836 25936 11876 25976
rect 2860 25852 2900 25892
rect 8812 25852 8852 25892
rect 12508 25852 12548 25892
rect 4928 25684 4968 25724
rect 5010 25684 5050 25724
rect 5092 25684 5132 25724
rect 5174 25684 5214 25724
rect 5256 25684 5296 25724
rect 1468 25516 1508 25556
rect 8035 25516 8075 25556
rect 9772 25516 9812 25556
rect 12508 25516 12548 25556
rect 8803 25432 8843 25472
rect 2956 25339 2996 25379
rect 4204 25348 4244 25388
rect 4684 25348 4724 25388
rect 5932 25339 5972 25379
rect 6316 25348 6356 25388
rect 7564 25339 7604 25379
rect 8188 25348 8228 25388
rect 8332 25348 8372 25388
rect 1228 25264 1268 25304
rect 1612 25264 1652 25304
rect 8476 25306 8516 25346
rect 8716 25348 8756 25388
rect 8951 25348 8991 25388
rect 9196 25348 9236 25388
rect 9964 25339 10004 25379
rect 11212 25348 11252 25388
rect 8611 25264 8651 25304
rect 9091 25264 9131 25304
rect 9292 25264 9332 25304
rect 11500 25264 11540 25304
rect 11884 25264 11924 25304
rect 12268 25264 12308 25304
rect 12124 25180 12164 25220
rect 1852 25096 1892 25136
rect 2764 25096 2804 25136
rect 6124 25096 6164 25136
rect 7756 25096 7796 25136
rect 11740 25096 11780 25136
rect 3688 24928 3728 24968
rect 3770 24928 3810 24968
rect 3852 24928 3892 24968
rect 3934 24928 3974 24968
rect 4016 24928 4056 24968
rect 4732 24760 4772 24800
rect 8659 24760 8699 24800
rect 12076 24760 12116 24800
rect 12508 24760 12548 24800
rect 2179 24592 2219 24632
rect 4492 24592 4532 24632
rect 7372 24592 7412 24632
rect 12268 24592 12308 24632
rect 2380 24508 2420 24548
rect 3628 24508 3668 24548
rect 6883 24508 6923 24548
rect 6988 24508 7028 24548
rect 7468 24508 7508 24548
rect 7948 24508 7988 24548
rect 8436 24508 8476 24548
rect 8812 24508 8852 24548
rect 10060 24508 10100 24548
rect 10636 24508 10676 24548
rect 11884 24508 11924 24548
rect 10252 24340 10292 24380
rect 4928 24172 4968 24212
rect 5010 24172 5050 24212
rect 5092 24172 5132 24212
rect 5174 24172 5214 24212
rect 5256 24172 5296 24212
rect 10012 24004 10052 24044
rect 10684 24004 10724 24044
rect 4108 23836 4148 23876
rect 5356 23827 5396 23867
rect 5740 23836 5780 23876
rect 6988 23827 7028 23867
rect 7843 23836 7883 23876
rect 7948 23836 7988 23876
rect 8332 23836 8372 23876
rect 8908 23827 8948 23867
rect 9388 23827 9428 23867
rect 11020 23827 11060 23867
rect 12268 23836 12308 23876
rect 1228 23752 1268 23792
rect 8428 23752 8468 23792
rect 9619 23752 9659 23792
rect 9772 23752 9812 23792
rect 10444 23752 10484 23792
rect 1468 23584 1508 23624
rect 5548 23584 5588 23624
rect 7180 23584 7220 23624
rect 10828 23584 10868 23624
rect 3688 23416 3728 23456
rect 3770 23416 3810 23456
rect 3852 23416 3892 23456
rect 3934 23416 3974 23456
rect 4016 23416 4056 23456
rect 6364 23248 6404 23288
rect 9820 23248 9860 23288
rect 10204 23248 10244 23288
rect 9436 23164 9476 23204
rect 10828 23164 10868 23204
rect 1228 23080 1268 23120
rect 1468 23080 1508 23120
rect 4684 23080 4724 23120
rect 5971 23080 6011 23120
rect 6124 23080 6164 23120
rect 8140 23080 8180 23120
rect 9580 23080 9620 23120
rect 9964 23080 10004 23120
rect 10348 23080 10388 23120
rect 10588 23080 10628 23120
rect 2476 22996 2516 23036
rect 3724 22996 3764 23036
rect 4174 22996 4214 23036
rect 4298 22996 4338 23036
rect 4780 22996 4820 23036
rect 5260 22996 5300 23036
rect 5748 22996 5788 23036
rect 7651 22996 7691 23036
rect 7756 22996 7796 23036
rect 8236 22996 8276 23036
rect 8716 22996 8756 23036
rect 9204 22996 9244 23036
rect 11020 22996 11060 23036
rect 12268 22996 12308 23036
rect 3916 22828 3956 22868
rect 4928 22660 4968 22700
rect 5010 22660 5050 22700
rect 5092 22660 5132 22700
rect 5174 22660 5214 22700
rect 5256 22660 5296 22700
rect 9100 22492 9140 22532
rect 9916 22492 9956 22532
rect 10300 22492 10340 22532
rect 10684 22492 10724 22532
rect 7132 22408 7172 22448
rect 2860 22324 2900 22364
rect 4108 22315 4148 22355
rect 4579 22324 4619 22364
rect 4684 22324 4724 22364
rect 5068 22324 5108 22364
rect 5644 22315 5684 22355
rect 6124 22315 6164 22355
rect 7363 22324 7403 22364
rect 7468 22324 7508 22364
rect 7852 22324 7892 22364
rect 8428 22315 8468 22355
rect 8908 22315 8948 22355
rect 11020 22315 11060 22355
rect 12268 22324 12308 22364
rect 1228 22240 1268 22280
rect 5164 22240 5204 22280
rect 6355 22240 6395 22280
rect 6508 22240 6548 22280
rect 6892 22240 6932 22280
rect 7948 22240 7988 22280
rect 9292 22240 9332 22280
rect 9676 22240 9716 22280
rect 10060 22240 10100 22280
rect 10444 22240 10484 22280
rect 6748 22156 6788 22196
rect 9532 22156 9572 22196
rect 1468 22072 1508 22112
rect 4300 22072 4340 22112
rect 10828 22072 10868 22112
rect 3688 21904 3728 21944
rect 3770 21904 3810 21944
rect 3852 21904 3892 21944
rect 3934 21904 3974 21944
rect 4016 21904 4056 21944
rect 4108 21736 4148 21776
rect 2284 21568 2324 21608
rect 4396 21568 4436 21608
rect 5356 21568 5396 21608
rect 8908 21568 8948 21608
rect 9292 21568 9332 21608
rect 9676 21568 9716 21608
rect 10252 21568 10292 21608
rect 10444 21568 10484 21608
rect 10684 21568 10724 21608
rect 2668 21484 2708 21524
rect 3916 21484 3956 21524
rect 4867 21484 4907 21524
rect 4972 21484 5012 21524
rect 5452 21484 5492 21524
rect 5932 21484 5972 21524
rect 6451 21484 6491 21524
rect 6796 21484 6836 21524
rect 8044 21484 8084 21524
rect 11020 21484 11060 21524
rect 12268 21484 12308 21524
rect 2524 21400 2564 21440
rect 8236 21400 8276 21440
rect 9916 21400 9956 21440
rect 4636 21316 4676 21356
rect 6604 21316 6644 21356
rect 9148 21316 9188 21356
rect 9532 21316 9572 21356
rect 10012 21316 10052 21356
rect 10828 21316 10868 21356
rect 4928 21148 4968 21188
rect 5010 21148 5050 21188
rect 5092 21148 5132 21188
rect 5174 21148 5214 21188
rect 5256 21148 5296 21188
rect 3820 20980 3860 21020
rect 7276 20980 7316 21020
rect 8380 20980 8420 21020
rect 12124 20980 12164 21020
rect 12508 20980 12548 21020
rect 3628 20896 3668 20936
rect 9676 20896 9716 20936
rect 2188 20812 2228 20852
rect 3436 20803 3476 20843
rect 4003 20812 4043 20852
rect 4492 20803 4532 20843
rect 4972 20812 5012 20852
rect 5452 20812 5492 20852
rect 5570 20812 5610 20852
rect 5836 20812 5876 20852
rect 7084 20803 7124 20843
rect 9292 20812 9332 20852
rect 9571 20812 9611 20852
rect 10348 20803 10388 20843
rect 11596 20812 11636 20852
rect 1228 20728 1268 20768
rect 5068 20728 5108 20768
rect 7948 20728 7988 20768
rect 8380 20728 8420 20768
rect 8620 20728 8660 20768
rect 11884 20728 11924 20768
rect 12268 20728 12308 20768
rect 9964 20644 10004 20684
rect 1468 20560 1508 20600
rect 7708 20560 7748 20600
rect 10156 20560 10196 20600
rect 3688 20392 3728 20432
rect 3770 20392 3810 20432
rect 3852 20392 3892 20432
rect 3934 20392 3974 20432
rect 4016 20392 4056 20432
rect 4108 20224 4148 20264
rect 9388 20224 9428 20264
rect 9820 20140 9860 20180
rect 1228 20056 1268 20096
rect 4588 20056 4628 20096
rect 5548 20056 5588 20096
rect 6988 20056 7028 20096
rect 7228 20056 7268 20096
rect 9580 20056 9620 20096
rect 9916 20056 9956 20096
rect 10156 20056 10196 20096
rect 10924 20056 10964 20096
rect 2668 19972 2708 20012
rect 3916 19972 3956 20012
rect 7948 19972 7988 20012
rect 9196 19972 9236 20012
rect 10435 19972 10475 20012
rect 10540 19972 10580 20012
rect 11020 19972 11060 20012
rect 11500 19972 11540 20012
rect 12019 19972 12059 20012
rect 5308 19888 5348 19928
rect 1468 19804 1508 19844
rect 4828 19804 4868 19844
rect 12172 19804 12212 19844
rect 4928 19636 4968 19676
rect 5010 19636 5050 19676
rect 5092 19636 5132 19676
rect 5174 19636 5214 19676
rect 5256 19636 5296 19676
rect 1468 19468 1508 19508
rect 3628 19468 3668 19508
rect 10588 19468 10628 19508
rect 12172 19468 12212 19508
rect 2188 19300 2228 19340
rect 3436 19291 3476 19331
rect 6604 19300 6644 19340
rect 7852 19291 7892 19331
rect 8236 19300 8276 19340
rect 9484 19291 9524 19331
rect 10732 19300 10772 19340
rect 11980 19291 12020 19331
rect 1228 19216 1268 19256
rect 9964 19216 10004 19256
rect 10348 19216 10388 19256
rect 10204 19132 10244 19172
rect 8044 19048 8084 19088
rect 9676 19048 9716 19088
rect 3688 18880 3728 18920
rect 3770 18880 3810 18920
rect 3852 18880 3892 18920
rect 3934 18880 3974 18920
rect 4016 18880 4056 18920
rect 3388 18628 3428 18668
rect 8860 18628 8900 18668
rect 12508 18628 12548 18668
rect 3148 18544 3188 18584
rect 7180 18544 7220 18584
rect 8467 18544 8507 18584
rect 8620 18544 8660 18584
rect 9772 18544 9812 18584
rect 11404 18544 11444 18584
rect 11884 18544 11924 18584
rect 12124 18544 12164 18584
rect 12268 18544 12308 18584
rect 4012 18460 4052 18500
rect 5260 18460 5300 18500
rect 6691 18460 6731 18500
rect 6796 18460 6836 18500
rect 7276 18460 7316 18500
rect 7756 18460 7796 18500
rect 8244 18460 8284 18500
rect 9283 18460 9323 18500
rect 9388 18460 9428 18500
rect 9868 18460 9908 18500
rect 10348 18460 10388 18500
rect 10867 18460 10907 18500
rect 5452 18376 5492 18416
rect 11020 18292 11060 18332
rect 11644 18292 11684 18332
rect 4928 18124 4968 18164
rect 5010 18124 5050 18164
rect 5092 18124 5132 18164
rect 5174 18124 5214 18164
rect 5256 18124 5296 18164
rect 1468 17956 1508 17996
rect 6028 17956 6068 17996
rect 6796 17956 6836 17996
rect 9100 17956 9140 17996
rect 9916 17956 9956 17996
rect 10300 17956 10340 17996
rect 12268 17956 12308 17996
rect 2332 17872 2372 17912
rect 9244 17872 9284 17912
rect 2476 17788 2516 17828
rect 3724 17779 3764 17819
rect 5539 17788 5579 17828
rect 6133 17788 6173 17828
rect 1228 17704 1268 17744
rect 2092 17704 2132 17744
rect 4108 17704 4148 17744
rect 4780 17704 4820 17744
rect 5020 17704 5060 17744
rect 6243 17704 6283 17744
rect 6364 17746 6404 17786
rect 6508 17788 6548 17828
rect 6650 17788 6690 17828
rect 7660 17788 7700 17828
rect 8908 17779 8948 17819
rect 10531 17788 10571 17828
rect 10636 17788 10676 17828
rect 11020 17788 11060 17828
rect 11596 17779 11636 17819
rect 12076 17779 12116 17819
rect 9484 17704 9524 17744
rect 9676 17704 9716 17744
rect 10060 17704 10100 17744
rect 11116 17704 11156 17744
rect 4348 17620 4388 17660
rect 5511 17620 5551 17660
rect 3916 17536 3956 17576
rect 5731 17536 5771 17576
rect 3688 17368 3728 17408
rect 3770 17368 3810 17408
rect 3852 17368 3892 17408
rect 3934 17368 3974 17408
rect 4016 17368 4056 17408
rect 7468 17200 7508 17240
rect 11836 17200 11876 17240
rect 12508 17200 12548 17240
rect 1468 17116 1508 17156
rect 4588 17116 4628 17156
rect 1228 17032 1268 17072
rect 10444 17032 10484 17072
rect 12076 17032 12116 17072
rect 12268 17032 12308 17072
rect 3148 16948 3188 16988
rect 4396 16948 4436 16988
rect 4867 16948 4907 16988
rect 5165 16948 5205 16988
rect 5340 16948 5380 16988
rect 5502 16948 5542 16988
rect 5635 16939 5675 16979
rect 5739 16948 5779 16988
rect 5857 16959 5897 16999
rect 6220 16948 6260 16988
rect 6339 16948 6379 16988
rect 6457 16948 6497 16988
rect 6700 16948 6740 16988
rect 6844 16981 6884 17021
rect 7171 16948 7211 16988
rect 7479 16948 7519 16988
rect 7649 16948 7689 16988
rect 7948 16948 7988 16988
rect 8236 16948 8276 16988
rect 9484 16948 9524 16988
rect 9955 16948 9995 16988
rect 10060 16948 10100 16988
rect 10540 16948 10580 16988
rect 11020 16948 11060 16988
rect 11539 16948 11579 16988
rect 7852 16864 7892 16904
rect 9676 16864 9716 16904
rect 4588 16780 4628 16820
rect 5068 16780 5108 16820
rect 5827 16780 5867 16820
rect 6124 16780 6164 16820
rect 6988 16780 7028 16820
rect 7267 16780 7307 16820
rect 7747 16780 7787 16820
rect 11692 16780 11732 16820
rect 4928 16612 4968 16652
rect 5010 16612 5050 16652
rect 5092 16612 5132 16652
rect 5174 16612 5214 16652
rect 5256 16612 5296 16652
rect 3340 16444 3380 16484
rect 4972 16444 5012 16484
rect 7276 16444 7316 16484
rect 9724 16444 9764 16484
rect 11404 16444 11444 16484
rect 11836 16444 11876 16484
rect 12508 16444 12548 16484
rect 1468 16360 1508 16400
rect 1900 16276 1940 16316
rect 3148 16267 3188 16307
rect 3532 16276 3572 16316
rect 4780 16267 4820 16307
rect 5539 16276 5579 16316
rect 5644 16276 5684 16316
rect 6028 16276 6068 16316
rect 6604 16267 6644 16307
rect 7084 16267 7124 16307
rect 7555 16276 7595 16316
rect 7660 16276 7700 16316
rect 8044 16276 8084 16316
rect 8620 16267 8660 16307
rect 9100 16267 9140 16307
rect 9964 16276 10004 16316
rect 11212 16267 11252 16307
rect 1228 16192 1268 16232
rect 6124 16192 6164 16232
rect 8140 16192 8180 16232
rect 9331 16192 9371 16232
rect 9484 16192 9524 16232
rect 11596 16192 11636 16232
rect 12268 16192 12308 16232
rect 4972 16024 5012 16064
rect 3688 15856 3728 15896
rect 3770 15856 3810 15896
rect 3852 15856 3892 15896
rect 3934 15856 3974 15896
rect 4016 15856 4056 15896
rect 6163 15688 6203 15728
rect 9004 15688 9044 15728
rect 12268 15688 12308 15728
rect 3916 15604 3956 15644
rect 2092 15520 2132 15560
rect 4876 15520 4916 15560
rect 6892 15520 6932 15560
rect 8419 15520 8459 15560
rect 2476 15436 2516 15476
rect 3724 15436 3764 15476
rect 4387 15436 4427 15476
rect 4492 15436 4532 15476
rect 4972 15436 5012 15476
rect 5452 15436 5492 15476
rect 5940 15436 5980 15476
rect 6403 15436 6443 15476
rect 6508 15436 6548 15476
rect 6988 15436 7028 15476
rect 7468 15436 7508 15476
rect 7956 15436 7996 15476
rect 8279 15436 8319 15476
rect 8524 15436 8564 15476
rect 9196 15436 9236 15476
rect 10444 15436 10484 15476
rect 10828 15436 10868 15476
rect 12076 15436 12116 15476
rect 8611 15352 8651 15392
rect 2332 15268 2372 15308
rect 8140 15268 8180 15308
rect 4928 15100 4968 15140
rect 5010 15100 5050 15140
rect 5092 15100 5132 15140
rect 5174 15100 5214 15140
rect 5256 15100 5296 15140
rect 3619 14932 3659 14972
rect 3724 14932 3764 14972
rect 7948 14932 7988 14972
rect 9484 14932 9524 14972
rect 11356 14932 11396 14972
rect 3834 14848 3874 14888
rect 5260 14848 5300 14888
rect 8428 14848 8468 14888
rect 3139 14764 3179 14804
rect 3523 14764 3563 14804
rect 4036 14764 4076 14804
rect 4195 14764 4235 14804
rect 4339 14764 4379 14804
rect 4483 14764 4523 14804
rect 4585 14764 4625 14804
rect 4876 14764 4916 14804
rect 5155 14764 5195 14804
rect 5740 14764 5780 14804
rect 5932 14764 5972 14804
rect 6211 14764 6251 14804
rect 6316 14764 6356 14804
rect 6700 14764 6740 14804
rect 7276 14755 7316 14795
rect 7756 14755 7796 14795
rect 8537 14764 8577 14804
rect 8812 14764 8852 14804
rect 9676 14755 9716 14795
rect 10924 14764 10964 14804
rect 1420 14680 1460 14720
rect 5836 14680 5876 14720
rect 6796 14680 6836 14720
rect 9292 14680 9332 14720
rect 11116 14680 11156 14720
rect 11692 14680 11732 14720
rect 12076 14680 12116 14720
rect 12460 14680 12500 14720
rect 3111 14596 3151 14636
rect 3331 14596 3371 14636
rect 5548 14596 5588 14636
rect 8140 14596 8180 14636
rect 11452 14596 11492 14636
rect 12220 14596 12260 14636
rect 1180 14512 1220 14552
rect 4588 14512 4628 14552
rect 9052 14512 9092 14552
rect 11836 14512 11876 14552
rect 3688 14344 3728 14384
rect 3770 14344 3810 14384
rect 3852 14344 3892 14384
rect 3934 14344 3974 14384
rect 4016 14344 4056 14384
rect 4876 14176 4916 14216
rect 8668 14176 8708 14216
rect 9052 14176 9092 14216
rect 10492 14176 10532 14216
rect 12076 14176 12116 14216
rect 12220 14176 12260 14216
rect 7564 14092 7604 14132
rect 1420 14008 1460 14048
rect 8908 14008 8948 14048
rect 9292 14008 9332 14048
rect 9676 14008 9716 14048
rect 10060 14008 10100 14048
rect 10252 14008 10292 14048
rect 12460 14008 12500 14048
rect 3148 13924 3188 13964
rect 4396 13924 4436 13964
rect 5164 13924 5204 13964
rect 5260 13915 5300 13955
rect 5548 13924 5588 13964
rect 6071 13924 6111 13964
rect 6211 13924 6251 13964
rect 6316 13924 6356 13964
rect 6892 13924 6932 13964
rect 7147 13924 7187 13964
rect 7267 13924 7307 13964
rect 7756 13924 7796 13964
rect 7895 13957 7935 13997
rect 10636 13924 10676 13964
rect 11884 13924 11924 13964
rect 9436 13840 9476 13880
rect 1180 13756 1220 13796
rect 4588 13756 4628 13796
rect 6403 13756 6443 13796
rect 8044 13756 8084 13796
rect 9820 13756 9860 13796
rect 4928 13588 4968 13628
rect 5010 13588 5050 13628
rect 5092 13588 5132 13628
rect 5174 13588 5214 13628
rect 5256 13588 5296 13628
rect 4396 13420 4436 13460
rect 4675 13420 4715 13460
rect 5260 13420 5300 13460
rect 5548 13420 5588 13460
rect 6403 13420 6443 13460
rect 9724 13420 9764 13460
rect 10108 13420 10148 13460
rect 12220 13420 12260 13460
rect 4574 13336 4614 13376
rect 2956 13252 2996 13292
rect 4204 13243 4244 13283
rect 4780 13252 4820 13292
rect 4876 13243 4916 13283
rect 5059 13252 5099 13292
rect 5356 13252 5396 13292
rect 1420 13168 1460 13208
rect 5644 13210 5684 13250
rect 5763 13252 5803 13292
rect 5881 13252 5921 13292
rect 6071 13252 6111 13292
rect 6316 13252 6356 13292
rect 6743 13252 6783 13292
rect 6988 13252 7028 13292
rect 8044 13243 8084 13283
rect 9292 13252 9332 13292
rect 10540 13252 10580 13292
rect 11788 13243 11828 13283
rect 6211 13168 6251 13208
rect 6883 13168 6923 13208
rect 7084 13168 7124 13208
rect 9484 13168 9524 13208
rect 10348 13168 10388 13208
rect 12460 13168 12500 13208
rect 1180 13000 1220 13040
rect 7852 13000 7892 13040
rect 11980 13000 12020 13040
rect 3688 12832 3728 12872
rect 3770 12832 3810 12872
rect 3852 12832 3892 12872
rect 3934 12832 3974 12872
rect 4016 12832 4056 12872
rect 6028 12664 6068 12704
rect 8860 12664 8900 12704
rect 9532 12664 9572 12704
rect 11836 12664 11876 12704
rect 12220 12664 12260 12704
rect 3820 12496 3860 12536
rect 4972 12496 5012 12536
rect 4108 12412 4148 12452
rect 4363 12412 4403 12452
rect 4483 12412 4523 12452
rect 5068 12412 5108 12452
rect 5187 12412 5227 12452
rect 5308 12454 5348 12494
rect 7468 12496 7508 12536
rect 9100 12496 9140 12536
rect 9292 12496 9332 12536
rect 10252 12496 10292 12536
rect 12076 12496 12116 12536
rect 12460 12496 12500 12536
rect 5452 12412 5492 12452
rect 5594 12412 5634 12452
rect 5932 12412 5972 12452
rect 6124 12412 6164 12452
rect 6979 12412 7019 12452
rect 7084 12412 7124 12452
rect 7564 12412 7604 12452
rect 8044 12412 8084 12452
rect 8532 12412 8572 12452
rect 9763 12412 9803 12452
rect 9868 12412 9908 12452
rect 10348 12412 10388 12452
rect 10828 12412 10868 12452
rect 11347 12412 11387 12452
rect 3580 12244 3620 12284
rect 4828 12244 4868 12284
rect 5740 12244 5780 12284
rect 8716 12244 8756 12284
rect 11500 12244 11540 12284
rect 4928 12076 4968 12116
rect 5010 12076 5050 12116
rect 5092 12076 5132 12116
rect 5174 12076 5214 12116
rect 5256 12076 5296 12116
rect 3196 11908 3236 11948
rect 3868 11908 3908 11948
rect 7996 11908 8036 11948
rect 9100 11908 9140 11948
rect 11356 11908 11396 11948
rect 11836 11908 11876 11948
rect 12220 11908 12260 11948
rect 8092 11824 8132 11864
rect 5827 11740 5867 11780
rect 5932 11740 5972 11780
rect 6316 11740 6356 11780
rect 6892 11731 6932 11771
rect 7372 11731 7412 11771
rect 9283 11740 9323 11780
rect 9772 11731 9812 11771
rect 10252 11740 10292 11780
rect 10732 11740 10772 11780
rect 10850 11740 10890 11780
rect 1420 11656 1460 11696
rect 2956 11656 2996 11696
rect 4108 11656 4148 11696
rect 4300 11656 4340 11696
rect 4684 11656 4724 11696
rect 6412 11656 6452 11696
rect 7603 11656 7643 11696
rect 7756 11656 7796 11696
rect 8332 11656 8372 11696
rect 8716 11656 8756 11696
rect 8956 11656 8996 11696
rect 10348 11656 10388 11696
rect 11116 11656 11156 11696
rect 11692 11656 11732 11696
rect 12076 11656 12116 11696
rect 12460 11656 12500 11696
rect 11452 11572 11492 11612
rect 1180 11488 1220 11528
rect 4540 11488 4580 11528
rect 4924 11488 4964 11528
rect 3688 11320 3728 11360
rect 3770 11320 3810 11360
rect 3852 11320 3892 11360
rect 3934 11320 3974 11360
rect 4016 11320 4056 11360
rect 3916 11152 3956 11192
rect 5116 11152 5156 11192
rect 7612 11152 7652 11192
rect 11596 11152 11636 11192
rect 11836 11068 11876 11108
rect 1420 10984 1460 11024
rect 5539 10984 5579 11024
rect 6028 10984 6068 11024
rect 2476 10900 2516 10940
rect 3724 10900 3764 10940
rect 5260 10900 5300 10940
rect 5404 10942 5444 10982
rect 6259 10975 6299 11015
rect 7372 10984 7412 11024
rect 7756 10984 7796 11024
rect 8716 10984 8756 11024
rect 12076 10984 12116 11024
rect 12460 10984 12500 11024
rect 5644 10900 5684 10940
rect 6124 10900 6164 10940
rect 6361 10900 6401 10940
rect 8227 10900 8267 10940
rect 8332 10900 8372 10940
rect 8812 10900 8852 10940
rect 9292 10900 9332 10940
rect 9780 10900 9820 10940
rect 10156 10900 10196 10940
rect 11404 10900 11444 10940
rect 7996 10816 8036 10856
rect 1180 10732 1220 10772
rect 5731 10732 5771 10772
rect 9964 10732 10004 10772
rect 12220 10732 12260 10772
rect 4928 10564 4968 10604
rect 5010 10564 5050 10604
rect 5092 10564 5132 10604
rect 5174 10564 5214 10604
rect 5256 10564 5296 10604
rect 4108 10396 4148 10436
rect 5740 10396 5780 10436
rect 7756 10396 7796 10436
rect 9868 10396 9908 10436
rect 11836 10396 11876 10436
rect 8044 10312 8084 10352
rect 11452 10312 11492 10352
rect 2668 10228 2708 10268
rect 3916 10219 3956 10259
rect 4300 10228 4340 10268
rect 5548 10219 5588 10259
rect 6019 10228 6059 10268
rect 6129 10228 6169 10268
rect 6508 10228 6548 10268
rect 7084 10219 7124 10259
rect 7564 10219 7604 10259
rect 8236 10219 8276 10259
rect 9484 10228 9524 10268
rect 10060 10219 10100 10259
rect 11308 10228 11348 10268
rect 1420 10144 1460 10184
rect 6604 10144 6644 10184
rect 11692 10144 11732 10184
rect 12076 10144 12116 10184
rect 12460 10144 12500 10184
rect 12220 10060 12260 10100
rect 1180 9976 1220 10016
rect 3688 9808 3728 9848
rect 3770 9808 3810 9848
rect 3852 9808 3892 9848
rect 3934 9808 3974 9848
rect 4016 9808 4056 9848
rect 3004 9640 3044 9680
rect 4972 9640 5012 9680
rect 8092 9640 8132 9680
rect 9772 9640 9812 9680
rect 11836 9640 11876 9680
rect 9964 9556 10004 9596
rect 12220 9556 12260 9596
rect 2764 9472 2804 9512
rect 6124 9472 6164 9512
rect 7852 9472 7892 9512
rect 11596 9472 11636 9512
rect 12460 9472 12500 9512
rect 3532 9388 3572 9428
rect 4780 9388 4820 9428
rect 5164 9388 5204 9428
rect 5356 9388 5396 9428
rect 5635 9388 5675 9428
rect 5740 9388 5780 9428
rect 6220 9388 6260 9428
rect 6700 9388 6740 9428
rect 7219 9388 7259 9428
rect 8332 9388 8372 9428
rect 9580 9388 9620 9428
rect 10156 9388 10196 9428
rect 11404 9388 11444 9428
rect 5347 9220 5387 9260
rect 7372 9220 7412 9260
rect 4928 9052 4968 9092
rect 5010 9052 5050 9092
rect 5092 9052 5132 9092
rect 5174 9052 5214 9092
rect 5256 9052 5296 9092
rect 4492 8884 4532 8924
rect 5548 8884 5588 8924
rect 6307 8884 6347 8924
rect 7075 8884 7115 8924
rect 8908 8884 8948 8924
rect 10300 8884 10340 8924
rect 11068 8884 11108 8924
rect 11452 8884 11492 8924
rect 11836 8884 11876 8924
rect 9340 8800 9380 8840
rect 10684 8800 10724 8840
rect 3052 8716 3092 8756
rect 4300 8707 4340 8747
rect 4780 8716 4820 8756
rect 4924 8716 4964 8756
rect 5164 8707 5204 8747
rect 5263 8696 5303 8736
rect 5395 8707 5435 8747
rect 5740 8716 5780 8756
rect 5980 8716 6020 8756
rect 5875 8674 5915 8714
rect 6079 8707 6119 8747
rect 6454 8702 6494 8742
rect 6652 8716 6692 8756
rect 6763 8716 6803 8756
rect 6988 8716 7028 8756
rect 7468 8716 7508 8756
rect 8716 8707 8756 8747
rect 1420 8632 1460 8672
rect 6883 8632 6923 8672
rect 9100 8632 9140 8672
rect 10540 8632 10580 8672
rect 10924 8632 10964 8672
rect 11308 8632 11348 8672
rect 11692 8632 11732 8672
rect 12076 8632 12116 8672
rect 12460 8632 12500 8672
rect 1180 8464 1220 8504
rect 6028 8464 6068 8504
rect 12220 8464 12260 8504
rect 3688 8296 3728 8336
rect 3770 8296 3810 8336
rect 3852 8296 3892 8336
rect 3934 8296 3974 8336
rect 4016 8296 4056 8336
rect 5548 8128 5588 8168
rect 5836 8128 5876 8168
rect 8572 8128 8612 8168
rect 11068 8128 11108 8168
rect 11452 8128 11492 8168
rect 9676 8044 9716 8084
rect 10108 8044 10148 8084
rect 1420 7960 1460 8000
rect 8332 7960 8372 8000
rect 4108 7876 4148 7916
rect 5356 7876 5396 7916
rect 5880 7918 5920 7958
rect 9868 7960 9908 8000
rect 11308 7960 11348 8000
rect 11692 7960 11732 8000
rect 12076 7960 12116 8000
rect 12220 7960 12260 8000
rect 12460 7960 12500 8000
rect 5740 7876 5780 7916
rect 5989 7876 6029 7916
rect 6700 7876 6740 7916
rect 7948 7876 7988 7916
rect 9004 7876 9044 7916
rect 9283 7876 9323 7916
rect 9388 7792 9428 7832
rect 1180 7708 1220 7748
rect 8140 7708 8180 7748
rect 11836 7708 11876 7748
rect 4928 7540 4968 7580
rect 5010 7540 5050 7580
rect 5092 7540 5132 7580
rect 5174 7540 5214 7580
rect 5256 7540 5296 7580
rect 5443 7288 5483 7328
rect 5111 7204 5151 7244
rect 5251 7204 5291 7244
rect 5356 7204 5396 7244
rect 6796 7204 6836 7244
rect 8044 7195 8084 7235
rect 1420 7120 1460 7160
rect 4684 7120 4724 7160
rect 4924 7120 4964 7160
rect 11308 7120 11348 7160
rect 11692 7120 11732 7160
rect 12076 7120 12116 7160
rect 12220 7120 12260 7160
rect 12460 7120 12500 7160
rect 8236 7036 8276 7076
rect 11452 7036 11492 7076
rect 1180 6952 1220 6992
rect 11068 6952 11108 6992
rect 11836 6952 11876 6992
rect 3688 6784 3728 6824
rect 3770 6784 3810 6824
rect 3852 6784 3892 6824
rect 3934 6784 3974 6824
rect 4016 6784 4056 6824
rect 5164 6616 5204 6656
rect 11836 6616 11876 6656
rect 7372 6532 7412 6572
rect 11692 6448 11732 6488
rect 12076 6448 12116 6488
rect 12460 6448 12500 6488
rect 3724 6364 3764 6404
rect 4972 6364 5012 6404
rect 6700 6364 6740 6404
rect 6979 6364 7019 6404
rect 7564 6364 7604 6404
rect 8812 6364 8852 6404
rect 7084 6280 7124 6320
rect 11452 6280 11492 6320
rect 9004 6196 9044 6236
rect 12220 6196 12260 6236
rect 4928 6028 4968 6068
rect 5010 6028 5050 6068
rect 5092 6028 5132 6068
rect 5174 6028 5214 6068
rect 5256 6028 5296 6068
rect 3052 5692 3092 5732
rect 4300 5683 4340 5723
rect 4684 5692 4724 5732
rect 5932 5683 5972 5723
rect 6316 5692 6356 5732
rect 7564 5683 7604 5723
rect 8035 5692 8075 5732
rect 8145 5692 8185 5732
rect 8524 5692 8564 5732
rect 9100 5683 9140 5723
rect 9580 5683 9620 5723
rect 1420 5608 1460 5648
rect 8620 5608 8660 5648
rect 9811 5608 9851 5648
rect 9964 5608 10004 5648
rect 10204 5608 10244 5648
rect 12076 5608 12116 5648
rect 12220 5608 12260 5648
rect 12460 5608 12500 5648
rect 4492 5524 4532 5564
rect 6124 5524 6164 5564
rect 7756 5524 7796 5564
rect 1180 5440 1220 5480
rect 11836 5440 11876 5480
rect 3688 5272 3728 5312
rect 3770 5272 3810 5312
rect 3852 5272 3892 5312
rect 3934 5272 3974 5312
rect 4016 5272 4056 5312
rect 5356 5104 5396 5144
rect 9820 5104 9860 5144
rect 12220 5020 12260 5060
rect 1228 4936 1268 4976
rect 6124 4936 6164 4976
rect 8140 4936 8180 4976
rect 9580 4936 9620 4976
rect 9916 4936 9956 4976
rect 10156 4936 10196 4976
rect 12076 4936 12116 4976
rect 12460 4936 12500 4976
rect 2284 4852 2324 4892
rect 3532 4852 3572 4892
rect 3916 4852 3956 4892
rect 5164 4852 5204 4892
rect 5635 4852 5675 4892
rect 5740 4852 5780 4892
rect 6220 4852 6260 4892
rect 6700 4852 6740 4892
rect 7188 4852 7228 4892
rect 7651 4852 7691 4892
rect 7756 4852 7796 4892
rect 8236 4852 8276 4892
rect 8716 4852 8756 4892
rect 9204 4852 9244 4892
rect 1468 4684 1508 4724
rect 3724 4684 3764 4724
rect 7372 4684 7412 4724
rect 9388 4684 9428 4724
rect 11836 4684 11876 4724
rect 4928 4516 4968 4556
rect 5010 4516 5050 4556
rect 5092 4516 5132 4556
rect 5174 4516 5214 4556
rect 5256 4516 5296 4556
rect 3388 4264 3428 4304
rect 5356 4264 5396 4304
rect 6988 4264 7028 4304
rect 9196 4264 9236 4304
rect 12220 4264 12260 4304
rect 3916 4180 3956 4220
rect 5164 4171 5204 4211
rect 5548 4180 5588 4220
rect 6796 4171 6836 4211
rect 7267 4180 7307 4220
rect 7372 4180 7412 4220
rect 7756 4180 7796 4220
rect 8332 4171 8372 4211
rect 8812 4171 8852 4211
rect 9388 4171 9428 4211
rect 10636 4180 10676 4220
rect 1420 4096 1460 4136
rect 3148 4096 3188 4136
rect 3532 4096 3572 4136
rect 7852 4096 7892 4136
rect 11692 4096 11732 4136
rect 12076 4096 12116 4136
rect 12460 4096 12500 4136
rect 3772 4012 3812 4052
rect 1180 3928 1220 3968
rect 9043 3928 9083 3968
rect 11452 3928 11492 3968
rect 11836 3928 11876 3968
rect 3688 3760 3728 3800
rect 3770 3760 3810 3800
rect 3852 3760 3892 3800
rect 3934 3760 3974 3800
rect 4016 3760 4056 3800
rect 5548 3592 5588 3632
rect 7180 3592 7220 3632
rect 9100 3592 9140 3632
rect 11836 3592 11876 3632
rect 12220 3592 12260 3632
rect 9628 3508 9668 3548
rect 9244 3424 9284 3464
rect 9484 3424 9524 3464
rect 9868 3424 9908 3464
rect 12076 3424 12116 3464
rect 12460 3424 12500 3464
rect 4108 3340 4148 3380
rect 5356 3340 5396 3380
rect 5740 3340 5780 3380
rect 6988 3340 7028 3380
rect 7660 3340 7700 3380
rect 8908 3340 8948 3380
rect 4928 3004 4968 3044
rect 5010 3004 5050 3044
rect 5092 3004 5132 3044
rect 5174 3004 5214 3044
rect 5256 3004 5296 3044
rect 8188 2836 8228 2876
rect 12220 2836 12260 2876
rect 7228 2752 7268 2792
rect 1420 2584 1460 2624
rect 5164 2584 5204 2624
rect 6988 2584 7028 2624
rect 7948 2584 7988 2624
rect 12460 2584 12500 2624
rect 1180 2416 1220 2456
rect 5404 2416 5444 2456
rect 3688 2248 3728 2288
rect 3770 2248 3810 2288
rect 3852 2248 3892 2288
rect 3934 2248 3974 2288
rect 4016 2248 4056 2288
rect 1468 2080 1508 2120
rect 1228 1912 1268 1952
rect 4928 1492 4968 1532
rect 5010 1492 5050 1532
rect 5092 1492 5132 1532
rect 5174 1492 5214 1532
rect 5256 1492 5296 1532
<< metal2 >>
rect 4919 46852 4928 46892
rect 4968 46852 5010 46892
rect 5050 46852 5092 46892
rect 5132 46852 5174 46892
rect 5214 46852 5256 46892
rect 5296 46852 5305 46892
rect 0 46808 90 46828
rect 0 46768 1228 46808
rect 1268 46768 1277 46808
rect 3052 46768 6892 46808
rect 6932 46768 6941 46808
rect 0 46748 90 46768
rect 1603 46684 1612 46724
rect 1652 46684 1660 46724
rect 1700 46684 1783 46724
rect 2179 46684 2188 46724
rect 2228 46684 2236 46724
rect 2276 46684 2359 46724
rect 2755 46684 2764 46724
rect 2804 46684 2812 46724
rect 2852 46684 2935 46724
rect 3052 46472 3092 46768
rect 3331 46684 3340 46724
rect 3380 46684 3388 46724
rect 3428 46684 3511 46724
rect 3907 46684 3916 46724
rect 3956 46684 3964 46724
rect 4004 46684 4087 46724
rect 4483 46684 4492 46724
rect 4532 46684 4540 46724
rect 4580 46684 4663 46724
rect 5107 46684 5116 46724
rect 5156 46684 5356 46724
rect 5396 46684 5405 46724
rect 5635 46684 5644 46724
rect 5684 46684 5692 46724
rect 5732 46684 5815 46724
rect 6211 46684 6220 46724
rect 6260 46684 6268 46724
rect 6308 46684 6391 46724
rect 6787 46684 6796 46724
rect 6836 46684 6844 46724
rect 6884 46684 6967 46724
rect 7363 46684 7372 46724
rect 7412 46684 7420 46724
rect 7460 46684 7543 46724
rect 7939 46684 7948 46724
rect 7988 46684 7996 46724
rect 8036 46684 8119 46724
rect 8515 46684 8524 46724
rect 8564 46684 8572 46724
rect 8612 46684 8695 46724
rect 9091 46684 9100 46724
rect 9140 46684 9148 46724
rect 9188 46684 9271 46724
rect 9667 46684 9676 46724
rect 9716 46684 9724 46724
rect 9764 46684 9847 46724
rect 10243 46684 10252 46724
rect 10292 46684 10300 46724
rect 10340 46684 10423 46724
rect 10819 46684 10828 46724
rect 10868 46684 10876 46724
rect 10916 46684 10999 46724
rect 11395 46684 11404 46724
rect 11444 46684 11452 46724
rect 11492 46684 11575 46724
rect 4204 46600 11020 46640
rect 11060 46600 11069 46640
rect 4204 46472 4244 46600
rect 8236 46516 10732 46556
rect 10772 46516 10781 46556
rect 8236 46472 8276 46516
rect 643 46432 652 46472
rect 692 46432 1228 46472
rect 1268 46432 1277 46472
rect 1769 46432 1900 46472
rect 1940 46432 1949 46472
rect 2345 46432 2476 46472
rect 2516 46432 2525 46472
rect 3043 46432 3052 46472
rect 3092 46432 3101 46472
rect 3619 46432 3628 46472
rect 3668 46432 3677 46472
rect 4195 46432 4204 46472
rect 4244 46432 4253 46472
rect 4771 46432 4780 46472
rect 4820 46432 4829 46472
rect 5347 46432 5356 46472
rect 5396 46432 5405 46472
rect 5801 46432 5932 46472
rect 5972 46432 5981 46472
rect 6377 46432 6508 46472
rect 6548 46432 6557 46472
rect 7075 46432 7084 46472
rect 7124 46432 7133 46472
rect 7529 46432 7660 46472
rect 7700 46432 7709 46472
rect 8227 46432 8236 46472
rect 8276 46432 8285 46472
rect 8803 46432 8812 46472
rect 8852 46432 8861 46472
rect 9257 46432 9388 46472
rect 9428 46432 9437 46472
rect 9955 46432 9964 46472
rect 10004 46432 10348 46472
rect 10388 46432 10397 46472
rect 10531 46432 10540 46472
rect 10580 46432 10828 46472
rect 10868 46432 10877 46472
rect 10985 46432 11116 46472
rect 11156 46432 11165 46472
rect 11299 46432 11308 46472
rect 11348 46432 11692 46472
rect 11732 46432 11741 46472
rect 11875 46432 11884 46472
rect 11924 46432 11933 46472
rect 12259 46432 12268 46472
rect 12308 46432 12748 46472
rect 12788 46432 12797 46472
rect 3628 46388 3668 46432
rect 3628 46348 4204 46388
rect 4244 46348 4253 46388
rect 1459 46264 1468 46304
rect 1508 46264 4684 46304
rect 4724 46264 4733 46304
rect 4780 46220 4820 46432
rect 5356 46304 5396 46432
rect 7084 46388 7124 46432
rect 8812 46388 8852 46432
rect 7084 46348 8620 46388
rect 8660 46348 8669 46388
rect 8812 46348 11212 46388
rect 11252 46348 11261 46388
rect 5356 46264 10060 46304
rect 10100 46264 10109 46304
rect 4780 46180 9964 46220
rect 10004 46180 10013 46220
rect 11884 46136 11924 46432
rect 12115 46264 12124 46304
rect 12164 46264 12364 46304
rect 12404 46264 12413 46304
rect 12499 46264 12508 46304
rect 12548 46264 13132 46304
rect 13172 46264 13181 46304
rect 3679 46096 3688 46136
rect 3728 46096 3770 46136
rect 3810 46096 3852 46136
rect 3892 46096 3934 46136
rect 3974 46096 4016 46136
rect 4056 46096 4065 46136
rect 6691 46096 6700 46136
rect 6740 46096 11924 46136
rect 11020 46012 12556 46052
rect 12596 46012 12605 46052
rect 11020 45968 11060 46012
rect 1027 45928 1036 45968
rect 1076 45928 1564 45968
rect 1604 45928 1613 45968
rect 10387 45928 10396 45968
rect 10436 45928 11060 45968
rect 11107 45928 11116 45968
rect 11156 45928 11260 45968
rect 11300 45928 11309 45968
rect 10771 45844 10780 45884
rect 10820 45844 11980 45884
rect 12020 45844 12029 45884
rect 0 45800 90 45820
rect 0 45760 652 45800
rect 692 45760 701 45800
rect 1097 45760 1228 45800
rect 1268 45760 1277 45800
rect 1673 45760 1804 45800
rect 1844 45760 1853 45800
rect 10147 45760 10156 45800
rect 10196 45760 10205 45800
rect 10409 45760 10540 45800
rect 10580 45760 10589 45800
rect 10915 45760 10924 45800
rect 10964 45760 10973 45800
rect 11369 45760 11500 45800
rect 11540 45760 11549 45800
rect 11753 45760 11788 45800
rect 11828 45760 11884 45800
rect 11924 45760 11933 45800
rect 12137 45760 12172 45800
rect 12212 45760 12268 45800
rect 12308 45760 12317 45800
rect 0 45740 90 45760
rect 10156 45632 10196 45760
rect 10924 45716 10964 45760
rect 10243 45676 10252 45716
rect 10292 45676 10964 45716
rect 10156 45592 11692 45632
rect 11732 45592 11741 45632
rect 1459 45508 1468 45548
rect 1508 45508 3436 45548
rect 3476 45508 3485 45548
rect 11155 45508 11164 45548
rect 11204 45508 12020 45548
rect 12115 45508 12124 45548
rect 12164 45508 12268 45548
rect 12308 45508 12317 45548
rect 12499 45508 12508 45548
rect 12548 45508 13036 45548
rect 13076 45508 13085 45548
rect 11980 45464 12020 45508
rect 13638 45464 13728 45484
rect 11980 45424 13728 45464
rect 13638 45404 13728 45424
rect 4919 45340 4928 45380
rect 4968 45340 5010 45380
rect 5050 45340 5092 45380
rect 5132 45340 5174 45380
rect 5214 45340 5256 45380
rect 5296 45340 5305 45380
rect 5683 45172 5692 45212
rect 5732 45172 5932 45212
rect 5972 45172 5981 45212
rect 8611 45172 8620 45212
rect 8660 45172 8668 45212
rect 8708 45172 8791 45212
rect 10051 45172 10060 45212
rect 10100 45172 10684 45212
rect 10724 45172 10733 45212
rect 10819 45172 10828 45212
rect 10868 45172 12028 45212
rect 12068 45172 12077 45212
rect 13638 45128 13728 45148
rect 4627 45088 4636 45128
rect 4676 45088 6508 45128
rect 6548 45088 6557 45128
rect 10339 45088 10348 45128
rect 10388 45088 11644 45128
rect 11684 45088 11693 45128
rect 12355 45088 12364 45128
rect 12404 45088 13728 45128
rect 13638 45068 13728 45088
rect 10348 45004 10924 45044
rect 10964 45004 10973 45044
rect 10348 44960 10388 45004
rect 67 44920 76 44960
rect 116 44920 1228 44960
rect 1268 44920 1277 44960
rect 4387 44920 4396 44960
rect 4436 44920 4445 44960
rect 5321 44920 5452 44960
rect 5492 44920 5501 44960
rect 8777 44920 8908 44960
rect 8948 44920 8957 44960
rect 10339 44920 10348 44960
rect 10388 44920 10397 44960
rect 10627 44920 10636 44960
rect 10676 44920 10924 44960
rect 10964 44920 10973 44960
rect 11203 44920 11212 44960
rect 11252 44920 11260 44960
rect 11300 44920 11383 44960
rect 11491 44920 11500 44960
rect 11540 44920 11671 44960
rect 11875 44920 11884 44960
rect 11924 44920 12055 44960
rect 12259 44920 12268 44960
rect 12308 44920 12364 44960
rect 12404 44920 12439 44960
rect 4396 44876 4436 44920
rect 4396 44836 5548 44876
rect 5588 44836 5597 44876
rect 10579 44836 10588 44876
rect 10628 44836 12212 44876
rect 0 44792 90 44812
rect 12172 44792 12212 44836
rect 13638 44792 13728 44812
rect 0 44752 76 44792
rect 116 44752 125 44792
rect 1459 44752 1468 44792
rect 1508 44752 2668 44792
rect 2708 44752 2717 44792
rect 12172 44752 13728 44792
rect 0 44732 90 44752
rect 13638 44732 13728 44752
rect 3679 44584 3688 44624
rect 3728 44584 3770 44624
rect 3810 44584 3852 44624
rect 3892 44584 3934 44624
rect 3974 44584 4016 44624
rect 4056 44584 4065 44624
rect 13638 44456 13728 44476
rect 9379 44416 9388 44456
rect 9428 44416 10492 44456
rect 10532 44416 10541 44456
rect 10723 44416 10732 44456
rect 10772 44416 10876 44456
rect 10916 44416 10925 44456
rect 11011 44416 11020 44456
rect 11060 44416 11644 44456
rect 11684 44416 11693 44456
rect 13123 44416 13132 44456
rect 13172 44416 13728 44456
rect 13638 44396 13728 44416
rect 9955 44332 9964 44372
rect 10004 44332 11260 44372
rect 11300 44332 11309 44372
rect 67 44248 76 44288
rect 116 44248 1228 44288
rect 1268 44248 1277 44288
rect 10601 44248 10732 44288
rect 10772 44248 10781 44288
rect 10985 44248 11116 44288
rect 11156 44248 11165 44288
rect 11369 44248 11500 44288
rect 11540 44248 11549 44288
rect 11753 44248 11884 44288
rect 11924 44248 11933 44288
rect 12259 44248 12268 44288
rect 12308 44248 12317 44288
rect 12268 44204 12308 44248
rect 5347 44164 5356 44204
rect 5396 44164 12308 44204
rect 13638 44120 13728 44140
rect 12259 44080 12268 44120
rect 12308 44080 13728 44120
rect 13638 44060 13728 44080
rect 1459 43996 1468 44036
rect 1508 43996 6124 44036
rect 6164 43996 6173 44036
rect 12499 43996 12508 44036
rect 12548 43996 13132 44036
rect 13172 43996 13181 44036
rect 4919 43828 4928 43868
rect 4968 43828 5010 43868
rect 5050 43828 5092 43868
rect 5132 43828 5174 43868
rect 5214 43828 5256 43868
rect 5296 43828 5305 43868
rect 0 43784 90 43804
rect 13638 43784 13728 43804
rect 0 43744 76 43784
rect 116 43744 125 43784
rect 13027 43744 13036 43784
rect 13076 43744 13728 43784
rect 0 43724 90 43744
rect 13638 43724 13728 43744
rect 7651 43660 7660 43700
rect 7700 43660 8380 43700
rect 8420 43660 8429 43700
rect 11347 43576 11356 43616
rect 11396 43576 13556 43616
rect 8035 43492 8044 43532
rect 8084 43492 12308 43532
rect 12268 43448 12308 43492
rect 13516 43448 13556 43576
rect 13638 43448 13728 43468
rect 1097 43408 1228 43448
rect 1268 43408 1277 43448
rect 8489 43408 8620 43448
rect 8660 43408 8669 43448
rect 11107 43408 11116 43448
rect 11156 43408 11165 43448
rect 11369 43408 11500 43448
rect 11540 43408 11549 43448
rect 11596 43408 11884 43448
rect 11924 43408 11933 43448
rect 12259 43408 12268 43448
rect 12308 43408 12317 43448
rect 13516 43408 13728 43448
rect 11116 43364 11156 43408
rect 7843 43324 7852 43364
rect 7892 43324 11156 43364
rect 11596 43280 11636 43408
rect 13638 43388 13728 43408
rect 1459 43240 1468 43280
rect 1508 43240 4588 43280
rect 4628 43240 4637 43280
rect 6499 43240 6508 43280
rect 6548 43240 11636 43280
rect 11731 43240 11740 43280
rect 11780 43240 11789 43280
rect 12115 43240 12124 43280
rect 12164 43240 12364 43280
rect 12404 43240 12413 43280
rect 12499 43240 12508 43280
rect 12548 43240 13036 43280
rect 13076 43240 13085 43280
rect 11740 43112 11780 43240
rect 13638 43112 13728 43132
rect 3679 43072 3688 43112
rect 3728 43072 3770 43112
rect 3810 43072 3852 43112
rect 3892 43072 3934 43112
rect 3974 43072 4016 43112
rect 4056 43072 4065 43112
rect 11740 43072 13728 43112
rect 13638 43052 13728 43072
rect 11177 42904 11260 42944
rect 11300 42904 11308 42944
rect 11348 42904 11357 42944
rect 11683 42904 11692 42944
rect 11732 42904 11740 42944
rect 11780 42904 11863 42944
rect 10531 42820 10540 42860
rect 10580 42820 11356 42860
rect 11396 42820 11405 42860
rect 0 42776 90 42796
rect 13638 42776 13728 42796
rect 0 42736 1228 42776
rect 1268 42736 1277 42776
rect 10889 42736 11020 42776
rect 11060 42736 11069 42776
rect 11465 42736 11596 42776
rect 11636 42736 11645 42776
rect 11849 42736 11980 42776
rect 12020 42736 12029 42776
rect 12259 42736 12268 42776
rect 12308 42736 12317 42776
rect 13123 42736 13132 42776
rect 13172 42736 13728 42776
rect 0 42716 90 42736
rect 12268 42692 12308 42736
rect 13638 42716 13728 42736
rect 7075 42652 7084 42692
rect 7124 42652 12308 42692
rect 12499 42484 12508 42524
rect 12548 42484 13132 42524
rect 13172 42484 13181 42524
rect 13638 42440 13728 42460
rect 12355 42400 12364 42440
rect 12404 42400 13728 42440
rect 13638 42380 13728 42400
rect 4919 42316 4928 42356
rect 4968 42316 5010 42356
rect 5050 42316 5092 42356
rect 5132 42316 5174 42356
rect 5214 42316 5256 42356
rect 5296 42316 5305 42356
rect 13638 42104 13728 42124
rect 13027 42064 13036 42104
rect 13076 42064 13728 42104
rect 13638 42044 13728 42064
rect 67 41896 76 41936
rect 116 41896 1228 41936
rect 1268 41896 1277 41936
rect 5827 41896 5836 41936
rect 5876 41896 11884 41936
rect 11924 41896 11933 41936
rect 12259 41896 12268 41936
rect 12308 41896 12317 41936
rect 12268 41852 12308 41896
rect 1459 41812 1468 41852
rect 1508 41812 2284 41852
rect 2324 41812 2333 41852
rect 10051 41812 10060 41852
rect 10100 41812 12308 41852
rect 0 41768 90 41788
rect 13638 41768 13728 41788
rect 0 41728 76 41768
rect 116 41728 125 41768
rect 12115 41728 12124 41768
rect 12164 41728 12173 41768
rect 12499 41728 12508 41768
rect 12548 41728 12940 41768
rect 12980 41728 12989 41768
rect 13123 41728 13132 41768
rect 13172 41728 13728 41768
rect 0 41708 90 41728
rect 12124 41600 12164 41728
rect 13638 41708 13728 41728
rect 3679 41560 3688 41600
rect 3728 41560 3770 41600
rect 3810 41560 3852 41600
rect 3892 41560 3934 41600
rect 3974 41560 4016 41600
rect 4056 41560 4065 41600
rect 12124 41560 13612 41600
rect 13652 41560 13661 41600
rect 13638 41432 13728 41452
rect 13603 41392 13612 41432
rect 13652 41392 13728 41432
rect 13638 41372 13728 41392
rect 67 41224 76 41264
rect 116 41224 1228 41264
rect 1268 41224 1277 41264
rect 2860 41224 11500 41264
rect 11540 41224 11549 41264
rect 11875 41224 11884 41264
rect 11924 41224 11933 41264
rect 12259 41224 12268 41264
rect 12308 41224 12460 41264
rect 12500 41224 12509 41264
rect 2860 41180 2900 41224
rect 11884 41180 11924 41224
rect 2563 41140 2572 41180
rect 2612 41140 2900 41180
rect 10819 41140 10828 41180
rect 10868 41140 11924 41180
rect 13638 41096 13728 41116
rect 11731 41056 11740 41096
rect 11780 41056 13728 41096
rect 13638 41036 13728 41056
rect 1459 40972 1468 41012
rect 1508 40972 2956 41012
rect 2996 40972 3005 41012
rect 12115 40972 12124 41012
rect 12164 40972 12173 41012
rect 12499 40972 12508 41012
rect 12548 40972 13132 41012
rect 13172 40972 13181 41012
rect 12124 40928 12164 40972
rect 12124 40888 12844 40928
rect 12884 40888 12893 40928
rect 4919 40804 4928 40844
rect 4968 40804 5010 40844
rect 5050 40804 5092 40844
rect 5132 40804 5174 40844
rect 5214 40804 5256 40844
rect 5296 40804 5305 40844
rect 0 40760 90 40780
rect 13638 40760 13728 40780
rect 0 40720 76 40760
rect 116 40720 125 40760
rect 12931 40720 12940 40760
rect 12980 40720 13728 40760
rect 0 40700 90 40720
rect 13638 40700 13728 40720
rect 11500 40468 13228 40508
rect 13268 40468 13277 40508
rect 11500 40424 11540 40468
rect 13638 40424 13728 40444
rect 1097 40384 1228 40424
rect 1268 40384 1277 40424
rect 2860 40384 6220 40424
rect 6260 40384 6269 40424
rect 11491 40384 11500 40424
rect 11540 40384 11549 40424
rect 11875 40384 11884 40424
rect 11924 40384 11933 40424
rect 12259 40384 12268 40424
rect 12308 40384 12556 40424
rect 12596 40384 12605 40424
rect 12835 40384 12844 40424
rect 12884 40384 13728 40424
rect 2860 40340 2900 40384
rect 11884 40340 11924 40384
rect 13638 40364 13728 40384
rect 1459 40300 1468 40340
rect 1508 40300 2900 40340
rect 5731 40300 5740 40340
rect 5780 40300 11924 40340
rect 12499 40300 12508 40340
rect 12548 40300 13420 40340
rect 13460 40300 13469 40340
rect 11731 40216 11740 40256
rect 11780 40216 11789 40256
rect 12115 40216 12124 40256
rect 12164 40216 12364 40256
rect 12404 40216 12413 40256
rect 11740 40088 11780 40216
rect 13638 40088 13728 40108
rect 3679 40048 3688 40088
rect 3728 40048 3770 40088
rect 3810 40048 3852 40088
rect 3892 40048 3934 40088
rect 3974 40048 4016 40088
rect 4056 40048 4065 40088
rect 11740 40048 13728 40088
rect 13638 40028 13728 40048
rect 9475 39796 9484 39836
rect 9524 39796 11540 39836
rect 0 39752 90 39772
rect 11500 39752 11540 39796
rect 13638 39752 13728 39772
rect 0 39712 1228 39752
rect 1268 39712 1277 39752
rect 11107 39712 11116 39752
rect 11156 39712 11165 39752
rect 11491 39712 11500 39752
rect 11540 39712 11549 39752
rect 11875 39712 11884 39752
rect 11924 39712 11933 39752
rect 12259 39712 12268 39752
rect 12308 39712 12317 39752
rect 13123 39712 13132 39752
rect 13172 39712 13728 39752
rect 0 39692 90 39712
rect 7180 39668 7220 39677
rect 8812 39668 8852 39677
rect 5923 39628 5932 39668
rect 5972 39628 6124 39668
rect 6164 39628 6604 39668
rect 6644 39628 6653 39668
rect 7145 39628 7180 39668
rect 7220 39628 7276 39668
rect 7316 39628 7325 39668
rect 7555 39628 7564 39668
rect 7604 39628 8332 39668
rect 8372 39628 8381 39668
rect 8777 39628 8812 39668
rect 8852 39628 8908 39668
rect 8948 39628 8957 39668
rect 7180 39619 7220 39628
rect 8812 39619 8852 39628
rect 7241 39460 7372 39500
rect 7412 39460 7421 39500
rect 8873 39460 9004 39500
rect 9044 39460 9053 39500
rect 4919 39292 4928 39332
rect 4968 39292 5010 39332
rect 5050 39292 5092 39332
rect 5132 39292 5174 39332
rect 5214 39292 5256 39332
rect 5296 39292 5305 39332
rect 11116 39164 11156 39712
rect 11884 39668 11924 39712
rect 11491 39628 11500 39668
rect 11540 39628 11924 39668
rect 12268 39668 12308 39712
rect 13638 39692 13728 39712
rect 12268 39628 13516 39668
rect 13556 39628 13565 39668
rect 12115 39544 12124 39584
rect 12164 39544 13324 39584
rect 13364 39544 13373 39584
rect 11347 39460 11356 39500
rect 11396 39460 11405 39500
rect 11731 39460 11740 39500
rect 11780 39460 11980 39500
rect 12020 39460 12029 39500
rect 12499 39460 12508 39500
rect 12548 39460 13132 39500
rect 13172 39460 13181 39500
rect 11356 39416 11396 39460
rect 13638 39416 13728 39436
rect 11356 39376 13728 39416
rect 13638 39356 13728 39376
rect 4819 39124 4828 39164
rect 4868 39124 11156 39164
rect 11347 39124 11356 39164
rect 11396 39124 12076 39164
rect 12116 39124 12125 39164
rect 12355 39124 12364 39164
rect 12404 39124 13652 39164
rect 13612 39100 13652 39124
rect 4435 39040 4444 39080
rect 4484 39040 5740 39080
rect 5780 39040 5789 39080
rect 6403 39040 6412 39080
rect 6452 39040 8276 39080
rect 8851 39040 8860 39080
rect 8900 39040 9140 39080
rect 9235 39040 9244 39080
rect 9284 39040 9676 39080
rect 9716 39040 9725 39080
rect 10963 39040 10972 39080
rect 11012 39040 13172 39080
rect 13612 39040 13728 39100
rect 4588 38956 4972 38996
rect 5012 38956 5021 38996
rect 6220 38987 6260 38996
rect 4588 38912 4628 38956
rect 6307 38956 6316 38996
rect 6356 38956 6691 38996
rect 6731 38956 6740 38996
rect 6787 38956 6796 38996
rect 6836 38956 6967 38996
rect 7171 38956 7180 38996
rect 7220 38956 7660 38996
rect 7700 38956 7709 38996
rect 7756 38987 8140 38996
rect 67 38872 76 38912
rect 116 38872 1228 38912
rect 1268 38872 1277 38912
rect 1459 38872 1468 38912
rect 1508 38872 2764 38912
rect 2804 38872 2813 38912
rect 4099 38872 4108 38912
rect 4148 38872 4204 38912
rect 4244 38872 4279 38912
rect 4387 38872 4396 38912
rect 4436 38872 4588 38912
rect 4628 38872 4637 38912
rect 6220 38828 6260 38947
rect 7796 38956 8140 38987
rect 8180 38956 8189 38996
rect 8236 38987 8276 39040
rect 7756 38938 7796 38947
rect 9100 38996 9140 39040
rect 9100 38956 10348 38996
rect 10388 38956 10397 38996
rect 12124 38956 12940 38996
rect 12980 38956 12989 38996
rect 8236 38938 8276 38947
rect 12124 38912 12164 38956
rect 13132 38912 13172 39040
rect 13638 39020 13728 39040
rect 7267 38872 7276 38912
rect 7316 38872 7468 38912
rect 7508 38872 7517 38912
rect 8458 38872 8467 38912
rect 8507 38872 8620 38912
rect 8660 38872 8669 38912
rect 8803 38872 8812 38912
rect 8852 38872 9004 38912
rect 9044 38872 9053 38912
rect 9257 38872 9388 38912
rect 9428 38872 9437 38912
rect 9619 38872 9628 38912
rect 9668 38872 9772 38912
rect 9812 38872 9821 38912
rect 9955 38872 9964 38912
rect 10004 38872 10732 38912
rect 10772 38872 10781 38912
rect 10985 38872 11116 38912
rect 11156 38872 11165 38912
rect 11491 38872 11500 38912
rect 11540 38872 11596 38912
rect 11636 38872 11671 38912
rect 11753 38872 11884 38912
rect 11924 38872 11933 38912
rect 12115 38872 12124 38912
rect 12164 38872 12173 38912
rect 12259 38872 12268 38912
rect 12308 38872 12364 38912
rect 12404 38872 12439 38912
rect 12499 38872 12508 38912
rect 12548 38872 13036 38912
rect 13076 38872 13085 38912
rect 13132 38872 13612 38912
rect 13652 38872 13661 38912
rect 6220 38788 8908 38828
rect 8948 38788 8957 38828
rect 0 38744 90 38764
rect 0 38704 76 38744
rect 116 38704 125 38744
rect 0 38684 90 38704
rect 3679 38536 3688 38576
rect 3728 38536 3770 38576
rect 3810 38536 3852 38576
rect 3892 38536 3934 38576
rect 3974 38536 4016 38576
rect 4056 38536 4065 38576
rect 6220 38492 6260 38788
rect 13638 38744 13728 38764
rect 11731 38704 11740 38744
rect 11780 38704 11788 38744
rect 11828 38704 11911 38744
rect 13603 38704 13612 38744
rect 13652 38704 13728 38744
rect 13638 38684 13728 38704
rect 5164 38452 6260 38492
rect 67 38200 76 38240
rect 116 38200 1228 38240
rect 1268 38200 1277 38240
rect 5068 38156 5108 38165
rect 5164 38156 5204 38452
rect 13638 38408 13728 38428
rect 5251 38368 5260 38408
rect 5300 38368 6316 38408
rect 6356 38368 6365 38408
rect 6412 38368 8332 38408
rect 8372 38368 8381 38408
rect 11971 38368 11980 38408
rect 12020 38368 13728 38408
rect 6412 38156 6452 38368
rect 13638 38348 13728 38368
rect 6883 38284 6892 38324
rect 6932 38284 8756 38324
rect 7180 38200 7372 38240
rect 7412 38200 7421 38240
rect 7529 38200 7660 38240
rect 7700 38200 7709 38240
rect 3689 38116 3820 38156
rect 3860 38116 4108 38156
rect 4148 38116 4157 38156
rect 5108 38116 5204 38156
rect 5443 38116 5452 38156
rect 5492 38116 6452 38156
rect 6700 38156 6740 38165
rect 7180 38156 7220 38200
rect 8716 38189 8756 38284
rect 8899 38200 8908 38240
rect 8948 38200 10388 38240
rect 10889 38200 11020 38240
rect 11060 38200 11069 38240
rect 11491 38200 11500 38240
rect 11540 38200 11549 38240
rect 11753 38200 11884 38240
rect 11924 38200 11933 38240
rect 12259 38200 12268 38240
rect 12308 38200 12317 38240
rect 8236 38156 8276 38165
rect 6740 38116 7028 38156
rect 7162 38116 7171 38156
rect 7211 38116 7220 38156
rect 7267 38116 7276 38156
rect 7316 38116 7325 38156
rect 7459 38116 7468 38156
rect 7508 38116 7756 38156
rect 7796 38116 7805 38156
rect 8105 38116 8236 38156
rect 8276 38116 8285 38156
rect 10348 38156 10388 38200
rect 8716 38140 8756 38149
rect 8812 38116 9100 38156
rect 9140 38116 9149 38156
rect 5068 38107 5108 38116
rect 5452 37988 5492 38116
rect 6700 38107 6740 38116
rect 1459 37948 1468 37988
rect 1508 37948 1516 37988
rect 1556 37948 1639 37988
rect 2659 37948 2668 37988
rect 2708 37948 5492 37988
rect 6988 37988 7028 38116
rect 7276 38072 7316 38116
rect 8236 38107 8276 38116
rect 7171 38032 7180 38072
rect 7220 38032 7316 38072
rect 6988 37948 7276 37988
rect 7316 37948 8140 37988
rect 8180 37948 8189 37988
rect 8812 37904 8852 38116
rect 10348 38107 10388 38116
rect 11500 38072 11540 38200
rect 12268 38156 12308 38200
rect 11683 38116 11692 38156
rect 11732 38116 12308 38156
rect 13638 38072 13728 38092
rect 11500 38032 11980 38072
rect 12020 38032 12029 38072
rect 12115 38032 12124 38072
rect 12164 38032 12652 38072
rect 12692 38032 12701 38072
rect 13411 38032 13420 38072
rect 13460 38032 13728 38072
rect 13638 38012 13728 38032
rect 8899 37948 8908 37988
rect 8948 37948 9388 37988
rect 9428 37948 9437 37988
rect 10531 37948 10540 37988
rect 10580 37948 10589 37988
rect 11107 37948 11116 37988
rect 11156 37948 11260 37988
rect 11300 37948 11309 37988
rect 11731 37948 11740 37988
rect 11780 37948 12364 37988
rect 12404 37948 12413 37988
rect 12499 37948 12508 37988
rect 12548 37948 12844 37988
rect 12884 37948 12893 37988
rect 6595 37864 6604 37904
rect 6644 37864 8852 37904
rect 4919 37780 4928 37820
rect 4968 37780 5010 37820
rect 5050 37780 5092 37820
rect 5132 37780 5174 37820
rect 5214 37780 5256 37820
rect 5296 37780 5305 37820
rect 0 37736 90 37756
rect 0 37696 76 37736
rect 116 37696 125 37736
rect 0 37676 90 37696
rect 8681 37612 8812 37652
rect 8852 37612 8861 37652
rect 4099 37528 4108 37568
rect 4148 37528 5396 37568
rect 5356 37484 5396 37528
rect 8140 37528 10292 37568
rect 3331 37444 3340 37484
rect 3380 37444 3724 37484
rect 3764 37444 3820 37484
rect 3860 37444 3924 37484
rect 4387 37444 4396 37484
rect 4436 37475 5012 37484
rect 4436 37444 4972 37475
rect 5347 37444 5356 37484
rect 5396 37444 5405 37484
rect 6019 37444 6028 37484
rect 6068 37475 6644 37484
rect 6068 37444 6604 37475
rect 4972 37426 5012 37435
rect 6923 37444 6988 37484
rect 7028 37444 7054 37484
rect 7094 37444 7103 37484
rect 7171 37444 7180 37484
rect 7220 37444 7276 37484
rect 7316 37444 7351 37484
rect 7459 37444 7468 37484
rect 7508 37444 7564 37484
rect 7604 37444 7639 37484
rect 8140 37475 8180 37528
rect 10252 37484 10292 37528
rect 10540 37484 10580 37948
rect 13638 37736 13728 37756
rect 12067 37696 12076 37736
rect 12116 37696 13728 37736
rect 13638 37676 13728 37696
rect 10915 37612 10924 37652
rect 10964 37612 11020 37652
rect 11060 37612 11095 37652
rect 6604 37426 6644 37435
rect 8140 37426 8180 37435
rect 8620 37475 8660 37484
rect 8995 37444 9004 37484
rect 9044 37444 9187 37484
rect 9227 37444 9236 37484
rect 9283 37444 9292 37484
rect 9332 37444 9463 37484
rect 9580 37444 9676 37484
rect 9716 37444 9725 37484
rect 10252 37475 10444 37484
rect 1097 37360 1228 37400
rect 1268 37360 1277 37400
rect 7625 37360 7660 37400
rect 7700 37360 7756 37400
rect 7796 37360 7805 37400
rect 8620 37316 8660 37435
rect 6787 37276 6796 37316
rect 6836 37276 8660 37316
rect 1459 37192 1468 37232
rect 1508 37192 3148 37232
rect 3188 37192 3197 37232
rect 5155 37192 5164 37232
rect 5204 37192 5740 37232
rect 5780 37192 5789 37232
rect 7747 37192 7756 37232
rect 7796 37192 8236 37232
rect 8276 37192 9292 37232
rect 9332 37192 9341 37232
rect 9580 37064 9620 37444
rect 10292 37444 10444 37475
rect 10484 37444 10493 37484
rect 10540 37475 10772 37484
rect 10540 37444 10732 37475
rect 10252 37426 10292 37435
rect 10732 37426 10772 37435
rect 13638 37400 13728 37420
rect 9676 37360 9772 37400
rect 9812 37360 9821 37400
rect 11177 37360 11308 37400
rect 11348 37360 11357 37400
rect 11491 37360 11500 37400
rect 11540 37360 11549 37400
rect 11753 37360 11884 37400
rect 11924 37360 11933 37400
rect 11980 37360 12268 37400
rect 12308 37360 12317 37400
rect 13315 37360 13324 37400
rect 13364 37360 13728 37400
rect 9676 37148 9716 37360
rect 11500 37316 11540 37360
rect 11980 37316 12020 37360
rect 13638 37340 13728 37360
rect 10051 37276 10060 37316
rect 10100 37276 11540 37316
rect 11596 37276 12020 37316
rect 12115 37276 12124 37316
rect 12164 37276 13420 37316
rect 13460 37276 13469 37316
rect 11596 37232 11636 37276
rect 9763 37192 9772 37232
rect 9812 37192 11068 37232
rect 11108 37192 11117 37232
rect 11395 37192 11404 37232
rect 11444 37192 11636 37232
rect 11731 37192 11740 37232
rect 11780 37192 11980 37232
rect 12020 37192 12029 37232
rect 12499 37192 12508 37232
rect 12548 37192 13612 37232
rect 13652 37192 13661 37232
rect 9676 37108 11020 37148
rect 11060 37108 11069 37148
rect 13638 37064 13728 37084
rect 3679 37024 3688 37064
rect 3728 37024 3770 37064
rect 3810 37024 3852 37064
rect 3892 37024 3934 37064
rect 3974 37024 4016 37064
rect 4056 37024 4065 37064
rect 9580 37024 11212 37064
rect 11252 37024 11261 37064
rect 11779 37024 11788 37064
rect 11828 37024 13728 37064
rect 13638 37004 13728 37024
rect 2179 36940 2188 36980
rect 2228 36940 6356 36980
rect 6316 36812 6356 36940
rect 9964 36940 12308 36980
rect 9964 36896 10004 36940
rect 6403 36856 6412 36896
rect 6452 36856 10004 36896
rect 10483 36856 10492 36896
rect 10532 36856 10828 36896
rect 10868 36856 10877 36896
rect 3331 36772 3340 36812
rect 3380 36772 4820 36812
rect 6316 36772 9908 36812
rect 0 36728 90 36748
rect 0 36688 1228 36728
rect 1268 36688 1277 36728
rect 0 36668 90 36688
rect 4396 36644 4436 36653
rect 4780 36644 4820 36772
rect 9868 36728 9908 36772
rect 10636 36772 12116 36812
rect 10636 36728 10676 36772
rect 6028 36688 7700 36728
rect 9475 36688 9484 36728
rect 9524 36688 9580 36728
rect 9620 36688 9655 36728
rect 9859 36688 9868 36728
rect 9908 36688 9917 36728
rect 10243 36688 10252 36728
rect 10292 36688 10636 36728
rect 10676 36688 10685 36728
rect 6028 36644 6068 36688
rect 7660 36644 7700 36688
rect 10828 36644 10868 36653
rect 12076 36644 12116 36772
rect 12268 36728 12308 36940
rect 13638 36728 13728 36748
rect 12259 36688 12268 36728
rect 12308 36688 12317 36728
rect 13123 36688 13132 36728
rect 13172 36688 13728 36728
rect 13638 36668 13728 36688
rect 3139 36604 3148 36644
rect 3188 36604 3197 36644
rect 4265 36604 4396 36644
rect 4436 36604 4445 36644
rect 4771 36604 4780 36644
rect 4820 36604 4829 36644
rect 5897 36604 6028 36644
rect 6068 36604 6077 36644
rect 6403 36604 6412 36644
rect 6452 36604 6461 36644
rect 10723 36604 10732 36644
rect 10772 36604 10828 36644
rect 10868 36604 10903 36644
rect 12067 36604 12076 36644
rect 12116 36604 12125 36644
rect 3148 36560 3188 36604
rect 4396 36595 4436 36604
rect 6028 36595 6068 36604
rect 3148 36520 4300 36560
rect 4340 36520 4349 36560
rect 4457 36436 4588 36476
rect 4628 36436 4637 36476
rect 6089 36436 6220 36476
rect 6260 36436 6269 36476
rect 6412 36392 6452 36604
rect 7660 36595 7700 36604
rect 10828 36595 10868 36604
rect 9283 36520 9292 36560
rect 9332 36520 10484 36560
rect 10531 36520 10540 36560
rect 10580 36520 10636 36560
rect 10676 36520 10711 36560
rect 10444 36476 10484 36520
rect 7843 36436 7852 36476
rect 7892 36436 8620 36476
rect 8660 36436 8669 36476
rect 9715 36436 9724 36476
rect 9764 36436 10004 36476
rect 10099 36436 10108 36476
rect 10148 36436 10388 36476
rect 10444 36436 11404 36476
rect 11444 36436 11453 36476
rect 12499 36436 12508 36476
rect 12548 36436 13324 36476
rect 13364 36436 13373 36476
rect 4291 36352 4300 36392
rect 4340 36352 6452 36392
rect 4919 36268 4928 36308
rect 4968 36268 5010 36308
rect 5050 36268 5092 36308
rect 5132 36268 5174 36308
rect 5214 36268 5256 36308
rect 5296 36268 5305 36308
rect 9964 36224 10004 36436
rect 10348 36392 10388 36436
rect 13638 36392 13728 36412
rect 10348 36352 12748 36392
rect 12788 36352 12797 36392
rect 12931 36352 12940 36392
rect 12980 36352 13728 36392
rect 13638 36332 13728 36352
rect 10147 36268 10156 36308
rect 10196 36268 10540 36308
rect 10580 36268 10589 36308
rect 9964 36184 13556 36224
rect 6307 36100 6316 36140
rect 6356 36100 6988 36140
rect 7028 36100 7037 36140
rect 9955 36100 9964 36140
rect 10004 36100 11308 36140
rect 11348 36100 11357 36140
rect 13516 36056 13556 36184
rect 13638 36056 13728 36076
rect 9868 36016 12076 36056
rect 12116 36016 12125 36056
rect 13516 36016 13728 36056
rect 9868 35972 9908 36016
rect 13638 35996 13728 36016
rect 4684 35932 4876 35972
rect 4916 35932 4925 35972
rect 6019 35932 6028 35972
rect 6068 35963 6199 35972
rect 6068 35932 6124 35963
rect 4684 35888 4724 35932
rect 6164 35932 6199 35963
rect 6412 35932 9908 35972
rect 10025 35932 10147 35972
rect 10196 35932 10205 35972
rect 10435 35932 10444 35972
rect 10484 35963 10676 35972
rect 10484 35932 10636 35963
rect 6124 35914 6164 35923
rect 6412 35888 6452 35932
rect 11011 35932 11020 35972
rect 11060 35932 11116 35972
rect 11156 35932 11191 35972
rect 11395 35932 11404 35972
rect 11444 35932 11596 35972
rect 11636 35932 11645 35972
rect 11705 35932 11714 35972
rect 11754 35932 12404 35972
rect 10636 35914 10676 35923
rect 11596 35888 11636 35932
rect 67 35848 76 35888
rect 116 35848 1228 35888
rect 1268 35848 1277 35888
rect 2467 35848 2476 35888
rect 2516 35848 4060 35888
rect 4100 35848 4109 35888
rect 4291 35848 4300 35888
rect 4340 35848 4349 35888
rect 4483 35848 4492 35888
rect 4532 35848 4684 35888
rect 4724 35848 4733 35888
rect 6220 35848 6452 35888
rect 6499 35848 6508 35888
rect 6548 35848 6604 35888
rect 6644 35848 6679 35888
rect 9065 35848 9196 35888
rect 9236 35848 9245 35888
rect 9571 35848 9580 35888
rect 9620 35848 10540 35888
rect 10580 35848 10589 35888
rect 10819 35848 10828 35888
rect 10868 35848 11212 35888
rect 11252 35848 11261 35888
rect 11596 35848 12076 35888
rect 12116 35848 12125 35888
rect 12259 35848 12268 35888
rect 12308 35848 12317 35888
rect 4300 35804 4340 35848
rect 6220 35804 6260 35848
rect 12268 35804 12308 35848
rect 4300 35764 4396 35804
rect 4436 35764 4445 35804
rect 4723 35764 4732 35804
rect 4772 35764 6260 35804
rect 9667 35764 9676 35804
rect 9716 35764 12308 35804
rect 0 35720 90 35740
rect 0 35680 76 35720
rect 116 35680 125 35720
rect 1459 35680 1468 35720
rect 1508 35680 2668 35720
rect 2708 35680 2717 35720
rect 6739 35680 6748 35720
rect 6788 35680 9292 35720
rect 9332 35680 9341 35720
rect 9427 35680 9436 35720
rect 9476 35680 9485 35720
rect 9811 35680 9820 35720
rect 9860 35680 9964 35720
rect 10004 35680 10013 35720
rect 0 35660 90 35680
rect 3679 35512 3688 35552
rect 3728 35512 3770 35552
rect 3810 35512 3852 35552
rect 3892 35512 3934 35552
rect 3974 35512 4016 35552
rect 4056 35512 4065 35552
rect 4147 35344 4156 35384
rect 4196 35344 9196 35384
rect 9236 35344 9245 35384
rect 9436 35300 9476 35680
rect 9955 35428 9964 35468
rect 10004 35428 11884 35468
rect 11924 35428 11933 35468
rect 12364 35384 12404 35932
rect 13638 35720 13728 35740
rect 12499 35680 12508 35720
rect 12548 35680 12556 35720
rect 12596 35680 12679 35720
rect 12739 35680 12748 35720
rect 12788 35680 13728 35720
rect 13638 35660 13728 35680
rect 13638 35384 13728 35404
rect 12364 35344 12460 35384
rect 12500 35344 12509 35384
rect 12556 35344 13728 35384
rect 12556 35300 12596 35344
rect 13638 35324 13728 35344
rect 7564 35260 8524 35300
rect 8564 35260 8573 35300
rect 9436 35260 12596 35300
rect 7564 35216 7604 35260
rect 67 35176 76 35216
rect 116 35176 1228 35216
rect 1268 35176 1277 35216
rect 3907 35176 3916 35216
rect 3956 35176 4108 35216
rect 4148 35176 4157 35216
rect 4387 35176 4396 35216
rect 4436 35176 5588 35216
rect 7555 35176 7564 35216
rect 7604 35176 7613 35216
rect 8842 35176 8851 35216
rect 8891 35176 9004 35216
rect 9044 35176 9053 35216
rect 5548 35132 5588 35176
rect 8140 35132 8180 35141
rect 9580 35132 9620 35141
rect 12268 35132 12308 35141
rect 4291 35092 4300 35132
rect 4340 35092 4684 35132
rect 4724 35092 4733 35132
rect 6211 35092 6220 35132
rect 6260 35092 7075 35132
rect 7115 35092 7124 35132
rect 7171 35092 7180 35132
rect 7220 35092 7276 35132
rect 7316 35092 7351 35132
rect 7529 35092 7660 35132
rect 7700 35092 7709 35132
rect 8180 35092 8236 35132
rect 8276 35092 8311 35132
rect 8611 35092 8620 35132
rect 8668 35092 8791 35132
rect 9475 35092 9484 35132
rect 9524 35092 9580 35132
rect 9620 35092 9655 35132
rect 10531 35092 10540 35132
rect 10580 35092 10828 35132
rect 10868 35092 11020 35132
rect 11060 35092 11404 35132
rect 11444 35092 11453 35132
rect 5548 35083 5588 35092
rect 8140 35083 8180 35092
rect 9580 35083 9620 35092
rect 12268 35048 12308 35092
rect 13638 35048 13728 35068
rect 5923 35008 5932 35048
rect 5972 35008 6604 35048
rect 6644 35008 6653 35048
rect 10723 35008 10732 35048
rect 10772 35008 11212 35048
rect 11252 35008 12308 35048
rect 12355 35008 12364 35048
rect 12404 35008 13728 35048
rect 13638 34988 13728 35008
rect 1459 34924 1468 34964
rect 1508 34924 2284 34964
rect 2324 34924 2333 34964
rect 5731 34924 5740 34964
rect 5780 34924 6124 34964
rect 6164 34924 6173 34964
rect 9235 34924 9244 34964
rect 9284 34924 9332 34964
rect 9379 34924 9388 34964
rect 9428 34924 9559 34964
rect 9292 34880 9332 34924
rect 9292 34840 10060 34880
rect 10100 34840 10109 34880
rect 4919 34756 4928 34796
rect 4968 34756 5010 34796
rect 5050 34756 5092 34796
rect 5132 34756 5174 34796
rect 5214 34756 5256 34796
rect 5296 34756 5305 34796
rect 0 34712 90 34732
rect 13638 34712 13728 34732
rect 0 34672 76 34712
rect 116 34672 125 34712
rect 13027 34672 13036 34712
rect 13076 34672 13728 34712
rect 0 34652 90 34672
rect 13638 34652 13728 34672
rect 7756 34588 9484 34628
rect 9524 34588 10004 34628
rect 7756 34544 7796 34588
rect 4099 34504 4108 34544
rect 4148 34504 6164 34544
rect 6124 34460 6164 34504
rect 7372 34504 7796 34544
rect 7852 34504 9772 34544
rect 9812 34504 9821 34544
rect 7372 34460 7412 34504
rect 7852 34460 7892 34504
rect 9964 34460 10004 34588
rect 4483 34420 4492 34460
rect 4532 34420 4684 34460
rect 4724 34420 4733 34460
rect 5740 34451 5780 34460
rect 6115 34420 6124 34460
rect 6164 34420 6173 34460
rect 7180 34451 7412 34460
rect 7180 34420 7372 34451
rect 5740 34376 5780 34411
rect 1097 34336 1228 34376
rect 1268 34336 1277 34376
rect 5740 34336 6604 34376
rect 6644 34336 6653 34376
rect 1459 34168 1468 34208
rect 1508 34168 3052 34208
rect 3092 34168 3101 34208
rect 5923 34168 5932 34208
rect 5972 34168 5981 34208
rect 3679 34000 3688 34040
rect 3728 34000 3770 34040
rect 3810 34000 3852 34040
rect 3892 34000 3934 34040
rect 3974 34000 4016 34040
rect 4056 34000 4065 34040
rect 4099 33748 4108 33788
rect 4148 33748 4157 33788
rect 0 33704 90 33724
rect 4108 33704 4148 33748
rect 0 33664 1228 33704
rect 1268 33664 1277 33704
rect 3340 33664 4148 33704
rect 0 33644 90 33664
rect 3340 33620 3380 33664
rect 4588 33620 4628 33629
rect 3180 33580 3244 33620
rect 3284 33580 3340 33620
rect 3380 33580 3389 33620
rect 4099 33580 4108 33620
rect 4148 33580 4588 33620
rect 5932 33620 5972 34168
rect 7180 33872 7220 34420
rect 7834 34420 7843 34460
rect 7883 34420 7892 34460
rect 7939 34420 7948 34460
rect 7988 34420 8119 34460
rect 8323 34420 8332 34460
rect 8372 34420 8381 34460
rect 8908 34451 8948 34460
rect 7372 34402 7412 34411
rect 8332 34292 8372 34420
rect 9257 34420 9388 34460
rect 9428 34420 9437 34460
rect 9964 34451 10060 34460
rect 8908 34376 8948 34411
rect 9388 34402 9428 34411
rect 10004 34420 10060 34451
rect 10100 34420 10164 34460
rect 10627 34420 10636 34460
rect 10676 34420 11212 34460
rect 11252 34420 11261 34460
rect 9964 34402 10004 34411
rect 13638 34376 13728 34396
rect 8419 34336 8428 34376
rect 8468 34336 8524 34376
rect 8564 34336 8599 34376
rect 8908 34336 9292 34376
rect 9332 34336 9341 34376
rect 11587 34336 11596 34376
rect 11636 34336 11645 34376
rect 11875 34336 11884 34376
rect 11924 34336 11933 34376
rect 12137 34336 12268 34376
rect 12308 34336 12317 34376
rect 12643 34336 12652 34376
rect 12692 34336 13728 34376
rect 11596 34292 11636 34336
rect 7267 34252 7276 34292
rect 7316 34252 8372 34292
rect 9619 34252 9628 34292
rect 9668 34252 11636 34292
rect 7555 34168 7564 34208
rect 7604 34168 7613 34208
rect 10723 34168 10732 34208
rect 10772 34168 11356 34208
rect 11396 34168 11405 34208
rect 6547 33832 6556 33872
rect 6596 33832 7220 33872
rect 7564 33788 7604 34168
rect 11884 34124 11924 34336
rect 13638 34316 13728 34336
rect 12115 34252 12124 34292
rect 12164 34252 12748 34292
rect 12788 34252 12797 34292
rect 12499 34168 12508 34208
rect 12548 34168 13228 34208
rect 13268 34168 13277 34208
rect 9955 34084 9964 34124
rect 10004 34084 11924 34124
rect 13638 34040 13728 34060
rect 11971 34000 11980 34040
rect 12020 34000 13728 34040
rect 13638 33980 13728 34000
rect 7564 33748 7988 33788
rect 11203 33748 11212 33788
rect 11252 33748 11308 33788
rect 11348 33748 11383 33788
rect 6307 33664 6316 33704
rect 6356 33664 6604 33704
rect 6644 33664 6653 33704
rect 7145 33664 7276 33704
rect 7316 33664 7325 33704
rect 7852 33620 7892 33629
rect 5932 33580 6787 33620
rect 6827 33580 6836 33620
rect 6883 33580 6892 33620
rect 6932 33580 6941 33620
rect 7363 33580 7372 33620
rect 7412 33580 7421 33620
rect 7651 33580 7660 33620
rect 7700 33580 7852 33620
rect 7948 33620 7988 33748
rect 13638 33704 13728 33724
rect 8554 33664 8563 33704
rect 8603 33664 8716 33704
rect 8756 33664 8765 33704
rect 9187 33664 9196 33704
rect 9236 33664 10156 33704
rect 10196 33664 10205 33704
rect 11875 33664 11884 33704
rect 11924 33664 11933 33704
rect 12137 33664 12268 33704
rect 12308 33664 12317 33704
rect 12835 33664 12844 33704
rect 12884 33664 13728 33704
rect 10828 33620 10868 33629
rect 7948 33580 8340 33620
rect 8380 33580 8389 33620
rect 9091 33580 9100 33620
rect 9140 33580 9580 33620
rect 9620 33580 9629 33620
rect 10435 33580 10444 33620
rect 10484 33580 10828 33620
rect 10868 33580 11212 33620
rect 11252 33580 11261 33620
rect 4588 33571 4628 33580
rect 6892 33536 6932 33580
rect 6403 33496 6412 33536
rect 6452 33496 6932 33536
rect 7372 33452 7412 33580
rect 7852 33536 7892 33580
rect 10828 33571 10868 33580
rect 7852 33496 9292 33536
rect 9332 33496 9341 33536
rect 10924 33496 11788 33536
rect 11828 33496 11837 33536
rect 10924 33452 10964 33496
rect 4771 33412 4780 33452
rect 4820 33412 4829 33452
rect 7372 33412 8524 33452
rect 8564 33412 8573 33452
rect 8947 33412 8956 33452
rect 8996 33412 9004 33452
rect 9044 33412 9127 33452
rect 9427 33412 9436 33452
rect 9476 33412 10964 33452
rect 11011 33412 11020 33452
rect 11060 33412 11212 33452
rect 11252 33412 11261 33452
rect 4780 33032 4820 33412
rect 11884 33368 11924 33664
rect 13638 33644 13728 33664
rect 12115 33412 12124 33452
rect 12164 33412 12268 33452
rect 12308 33412 12317 33452
rect 12499 33412 12508 33452
rect 12548 33412 13036 33452
rect 13076 33412 13085 33452
rect 13638 33368 13728 33388
rect 6979 33328 6988 33368
rect 7028 33328 11924 33368
rect 13411 33328 13420 33368
rect 13460 33328 13728 33368
rect 13638 33308 13728 33328
rect 4919 33244 4928 33284
rect 4968 33244 5010 33284
rect 5050 33244 5092 33284
rect 5132 33244 5174 33284
rect 5214 33244 5256 33284
rect 5296 33244 5305 33284
rect 9187 33244 9196 33284
rect 9236 33244 10444 33284
rect 10484 33244 10493 33284
rect 6220 33160 6644 33200
rect 6220 33032 6260 33160
rect 6604 33116 6644 33160
rect 6307 33076 6316 33116
rect 6356 33076 6365 33116
rect 6604 33076 8236 33116
rect 8276 33076 8285 33116
rect 8428 33076 11156 33116
rect 11395 33076 11404 33116
rect 11444 33076 11692 33116
rect 11732 33076 11741 33116
rect 4588 32992 4820 33032
rect 5644 32992 6260 33032
rect 4588 32948 4628 32992
rect 5644 32948 5684 32992
rect 6316 32948 6356 33076
rect 8428 33032 8468 33076
rect 11116 33032 11156 33076
rect 13638 33032 13728 33052
rect 6739 32992 6748 33032
rect 6788 32992 8468 33032
rect 9379 32992 9388 33032
rect 9428 32992 9524 33032
rect 9571 32992 9580 33032
rect 9620 32992 9812 33032
rect 11116 32992 12308 33032
rect 13603 32992 13612 33032
rect 13652 32992 13728 33032
rect 9484 32948 9524 32992
rect 9772 32948 9812 32992
rect 4570 32908 4579 32948
rect 4619 32908 4628 32948
rect 4675 32908 4684 32948
rect 4724 32908 4733 32948
rect 4780 32908 5068 32948
rect 5108 32908 5117 32948
rect 5443 32908 5452 32948
rect 5492 32939 5684 32948
rect 5492 32908 5644 32939
rect 67 32824 76 32864
rect 116 32824 1228 32864
rect 1268 32824 1277 32864
rect 3523 32824 3532 32864
rect 3572 32824 3724 32864
rect 3764 32824 3773 32864
rect 3977 32824 4108 32864
rect 4148 32824 4157 32864
rect 4108 32780 4148 32824
rect 3139 32740 3148 32780
rect 3188 32740 3964 32780
rect 4004 32740 4148 32780
rect 4684 32780 4724 32908
rect 4780 32864 4820 32908
rect 5993 32908 6124 32948
rect 6164 32908 6173 32948
rect 6316 32908 6932 32948
rect 7939 32908 7948 32948
rect 7988 32908 8716 32948
rect 8756 32908 8765 32948
rect 5644 32890 5684 32899
rect 6124 32890 6164 32899
rect 6892 32864 6932 32908
rect 9200 32906 9240 32915
rect 9484 32908 9667 32948
rect 9707 32908 9716 32948
rect 9763 32908 9772 32948
rect 9812 32908 9821 32948
rect 10243 32908 10252 32948
rect 10292 32908 10580 32948
rect 10697 32939 10828 32948
rect 10697 32908 10732 32939
rect 9196 32866 9200 32906
rect 9196 32864 9240 32866
rect 10540 32864 10580 32908
rect 10772 32908 10828 32939
rect 10868 32908 10877 32948
rect 11081 32908 11212 32948
rect 11252 32908 11261 32948
rect 10732 32890 10772 32899
rect 11212 32890 11252 32899
rect 12268 32864 12308 32992
rect 13638 32972 13728 32992
rect 4771 32824 4780 32864
rect 4820 32824 4829 32864
rect 5155 32824 5164 32864
rect 5204 32824 5356 32864
rect 5396 32824 5405 32864
rect 6538 32824 6547 32864
rect 6587 32824 6596 32864
rect 6883 32824 6892 32864
rect 6932 32824 6941 32864
rect 7433 32824 7564 32864
rect 7604 32824 7613 32864
rect 7747 32824 7756 32864
rect 7796 32824 9196 32864
rect 9236 32824 9245 32864
rect 10147 32824 10156 32864
rect 10196 32824 10327 32864
rect 10540 32824 10636 32864
rect 10676 32824 10685 32864
rect 11395 32824 11404 32864
rect 11444 32824 11884 32864
rect 11924 32824 11933 32864
rect 12259 32824 12268 32864
rect 12308 32824 12317 32864
rect 6556 32780 6596 32824
rect 4684 32740 4876 32780
rect 4916 32740 4925 32780
rect 6556 32740 7276 32780
rect 7316 32740 7325 32780
rect 7795 32740 7804 32780
rect 7844 32740 12692 32780
rect 0 32696 90 32716
rect 12652 32696 12692 32740
rect 13638 32696 13728 32716
rect 0 32656 76 32696
rect 116 32656 125 32696
rect 1459 32656 1468 32696
rect 1508 32656 2860 32696
rect 2900 32656 2909 32696
rect 4339 32656 4348 32696
rect 4388 32656 5644 32696
rect 5684 32656 5693 32696
rect 7123 32656 7132 32696
rect 7172 32656 9580 32696
rect 9620 32656 9629 32696
rect 10627 32656 10636 32696
rect 10676 32656 11692 32696
rect 11732 32656 11980 32696
rect 12020 32656 12029 32696
rect 12115 32656 12124 32696
rect 12164 32656 12268 32696
rect 12308 32656 12317 32696
rect 12425 32656 12508 32696
rect 12548 32656 12556 32696
rect 12596 32656 12605 32696
rect 12652 32656 13728 32696
rect 0 32636 90 32656
rect 13638 32636 13728 32656
rect 7075 32572 7084 32612
rect 7124 32572 10196 32612
rect 10156 32528 10196 32572
rect 3679 32488 3688 32528
rect 3728 32488 3770 32528
rect 3810 32488 3852 32528
rect 3892 32488 3934 32528
rect 3974 32488 4016 32528
rect 4056 32488 4065 32528
rect 6604 32488 10100 32528
rect 10147 32488 10156 32528
rect 10196 32488 10205 32528
rect 10252 32488 11404 32528
rect 11444 32488 11453 32528
rect 3715 32320 3724 32360
rect 3764 32320 5588 32360
rect 5548 32276 5588 32320
rect 6604 32276 6644 32488
rect 10060 32444 10100 32488
rect 10252 32444 10292 32488
rect 8227 32404 8236 32444
rect 8276 32404 10004 32444
rect 10060 32404 10292 32444
rect 9964 32360 10004 32404
rect 13638 32360 13728 32380
rect 9737 32320 9820 32360
rect 9860 32320 9868 32360
rect 9908 32320 9917 32360
rect 9964 32320 12460 32360
rect 12500 32320 12509 32360
rect 13315 32320 13324 32360
rect 13364 32320 13728 32360
rect 13638 32300 13728 32320
rect 5443 32236 5452 32276
rect 5492 32236 5501 32276
rect 5548 32236 6644 32276
rect 8707 32236 8716 32276
rect 8756 32236 9620 32276
rect 67 32152 76 32192
rect 116 32152 1228 32192
rect 1268 32152 1277 32192
rect 3916 32152 4108 32192
rect 4148 32152 4396 32192
rect 4436 32152 4445 32192
rect 4771 32152 4780 32192
rect 4820 32152 4876 32192
rect 4916 32152 4951 32192
rect 3916 32108 3956 32152
rect 5452 32108 5492 32236
rect 9580 32192 9620 32236
rect 6185 32152 6316 32192
rect 6356 32152 6365 32192
rect 9571 32152 9580 32192
rect 9620 32152 9629 32192
rect 11299 32152 11308 32192
rect 11348 32152 11357 32192
rect 9196 32108 9236 32117
rect 2537 32068 2668 32108
rect 2708 32068 2717 32108
rect 4235 32068 4300 32108
rect 4340 32068 4366 32108
rect 4406 32068 4415 32108
rect 4483 32068 4492 32108
rect 4532 32068 4916 32108
rect 4963 32068 4972 32108
rect 5012 32068 5356 32108
rect 5396 32068 5405 32108
rect 5931 32068 5940 32108
rect 5980 32068 5989 32108
rect 7939 32068 7948 32108
rect 7988 32068 8716 32108
rect 8756 32068 8765 32108
rect 8899 32068 8908 32108
rect 8948 32068 9196 32108
rect 10522 32068 10531 32108
rect 10580 32068 10711 32108
rect 3916 32059 3956 32068
rect 4876 32024 4916 32068
rect 5452 32059 5492 32068
rect 2860 31984 3724 32024
rect 3764 31984 3773 32024
rect 4745 31984 4876 32024
rect 4916 31984 4925 32024
rect 1459 31900 1468 31940
rect 1508 31900 1517 31940
rect 1468 31856 1508 31900
rect 2860 31856 2900 31984
rect 3427 31900 3436 31940
rect 3476 31900 3485 31940
rect 3977 31900 4012 31940
rect 4052 31900 4108 31940
rect 4148 31900 4157 31940
rect 1468 31816 2900 31856
rect 0 31688 90 31708
rect 3436 31688 3476 31900
rect 4876 31856 4916 31984
rect 5949 31940 5989 32068
rect 9196 32059 9236 32068
rect 13638 32024 13728 32044
rect 6124 31984 7276 32024
rect 7316 31984 7325 32024
rect 10138 31984 10147 32024
rect 10187 31984 10444 32024
rect 10484 31984 10493 32024
rect 12451 31984 12460 32024
rect 12500 31984 13728 32024
rect 6124 31940 6164 31984
rect 13638 31964 13728 31984
rect 5155 31900 5164 31940
rect 5204 31900 5989 31940
rect 6115 31900 6124 31940
rect 6164 31900 6173 31940
rect 6547 31900 6556 31940
rect 6596 31900 9140 31940
rect 9187 31900 9196 31940
rect 9236 31900 9388 31940
rect 9428 31900 9437 31940
rect 12451 31900 12460 31940
rect 12500 31900 13132 31940
rect 13172 31900 13181 31940
rect 9100 31856 9140 31900
rect 4876 31816 5684 31856
rect 9100 31816 10924 31856
rect 10964 31816 10973 31856
rect 4919 31732 4928 31772
rect 4968 31732 5010 31772
rect 5050 31732 5092 31772
rect 5132 31732 5174 31772
rect 5214 31732 5256 31772
rect 5296 31732 5305 31772
rect 0 31648 76 31688
rect 116 31648 125 31688
rect 3244 31648 3476 31688
rect 0 31628 90 31648
rect 3244 31436 3284 31648
rect 4169 31564 4300 31604
rect 4340 31564 4349 31604
rect 5644 31520 5684 31816
rect 13638 31688 13728 31708
rect 12739 31648 12748 31688
rect 12788 31648 13728 31688
rect 13638 31628 13728 31648
rect 6185 31564 6316 31604
rect 6356 31564 6365 31604
rect 6761 31564 6844 31604
rect 6884 31564 6892 31604
rect 6932 31564 6941 31604
rect 6988 31564 8236 31604
rect 8276 31564 8285 31604
rect 9235 31564 9244 31604
rect 9284 31564 9676 31604
rect 9716 31564 9725 31604
rect 6988 31520 7028 31564
rect 4579 31480 4588 31520
rect 4628 31480 4675 31520
rect 5644 31480 7028 31520
rect 7564 31480 8908 31520
rect 8948 31480 8957 31520
rect 4588 31436 4628 31480
rect 2851 31396 2860 31436
rect 2900 31396 3244 31436
rect 3284 31396 3293 31436
rect 3977 31396 4108 31436
rect 4148 31396 4157 31436
rect 4570 31396 4579 31436
rect 4619 31396 4628 31436
rect 4675 31396 4684 31436
rect 4724 31396 4876 31436
rect 4916 31396 4925 31436
rect 5059 31396 5068 31436
rect 5108 31396 5260 31436
rect 5300 31396 5309 31436
rect 5644 31427 5684 31480
rect 4108 31378 4148 31387
rect 5731 31396 5740 31436
rect 5780 31427 6164 31436
rect 5780 31396 6124 31427
rect 5644 31378 5684 31387
rect 6124 31378 6164 31387
rect 7564 31427 7604 31480
rect 8611 31396 8620 31436
rect 8660 31396 8812 31436
rect 8852 31396 8861 31436
rect 8908 31396 9580 31436
rect 9620 31396 9629 31436
rect 9859 31396 9868 31436
rect 9908 31427 10868 31436
rect 9908 31396 10828 31427
rect 7564 31378 7604 31387
rect 8908 31352 8948 31396
rect 10828 31378 10868 31387
rect 13638 31352 13728 31372
rect 1097 31312 1228 31352
rect 1268 31312 1277 31352
rect 4579 31312 4588 31352
rect 4628 31312 5164 31352
rect 5204 31312 5213 31352
rect 6691 31312 6700 31352
rect 6740 31312 7084 31352
rect 7124 31312 7133 31352
rect 8707 31312 8716 31352
rect 8756 31312 8948 31352
rect 8995 31312 9004 31352
rect 9044 31312 9100 31352
rect 9140 31312 9292 31352
rect 9332 31312 9341 31352
rect 11369 31312 11500 31352
rect 11540 31312 11549 31352
rect 11753 31312 11788 31352
rect 11828 31312 11884 31352
rect 11924 31312 11933 31352
rect 11980 31312 12268 31352
rect 12308 31312 12317 31352
rect 13219 31312 13228 31352
rect 13268 31312 13728 31352
rect 6700 31268 6740 31312
rect 2860 31228 5012 31268
rect 5059 31228 5068 31268
rect 5108 31228 6740 31268
rect 7084 31268 7124 31312
rect 11980 31268 12020 31312
rect 13638 31292 13728 31312
rect 7084 31228 7756 31268
rect 7796 31228 7805 31268
rect 8803 31228 8812 31268
rect 8852 31228 12020 31268
rect 12115 31228 12124 31268
rect 12164 31228 13324 31268
rect 13364 31228 13373 31268
rect 1459 31144 1468 31184
rect 1508 31144 1517 31184
rect 1468 31100 1508 31144
rect 2860 31100 2900 31228
rect 1468 31060 2900 31100
rect 4972 31016 5012 31228
rect 5251 31144 5260 31184
rect 5300 31144 6316 31184
rect 6356 31144 6365 31184
rect 6451 31144 6460 31184
rect 6500 31144 6604 31184
rect 6644 31144 6892 31184
rect 6932 31144 6941 31184
rect 7241 31144 7372 31184
rect 7412 31144 7421 31184
rect 10889 31144 11020 31184
rect 11060 31144 11069 31184
rect 11731 31144 11740 31184
rect 11780 31144 11980 31184
rect 12020 31144 12029 31184
rect 12499 31144 12508 31184
rect 12548 31144 13228 31184
rect 13268 31144 13277 31184
rect 13638 31016 13728 31036
rect 3679 30976 3688 31016
rect 3728 30976 3770 31016
rect 3810 30976 3852 31016
rect 3892 30976 3934 31016
rect 3974 30976 4016 31016
rect 4056 30976 4065 31016
rect 4972 30976 7276 31016
rect 7316 30976 7325 31016
rect 12355 30976 12364 31016
rect 12404 30976 13728 31016
rect 13638 30956 13728 30976
rect 7843 30892 7852 30932
rect 7892 30892 7901 30932
rect 7852 30848 7892 30892
rect 3148 30808 3244 30848
rect 3284 30808 3293 30848
rect 3667 30808 3676 30848
rect 3716 30808 4108 30848
rect 4148 30808 4300 30848
rect 4340 30808 4349 30848
rect 4396 30808 7892 30848
rect 8083 30808 8092 30848
rect 8132 30808 8908 30848
rect 8948 30808 8957 30848
rect 9859 30808 9868 30848
rect 9908 30808 9917 30848
rect 11587 30808 11596 30848
rect 11636 30808 11644 30848
rect 11684 30808 11767 30848
rect 0 30680 90 30700
rect 0 30640 1228 30680
rect 1268 30640 1277 30680
rect 0 30620 90 30640
rect 3148 30512 3188 30808
rect 4396 30764 4436 30808
rect 3715 30724 3724 30764
rect 3764 30724 4436 30764
rect 4867 30724 4876 30764
rect 4916 30724 7084 30764
rect 7124 30724 7133 30764
rect 3235 30640 3244 30680
rect 3284 30640 3436 30680
rect 3476 30640 3485 30680
rect 5068 30596 5108 30605
rect 5644 30596 5684 30724
rect 6019 30640 6028 30680
rect 6068 30640 6316 30680
rect 6356 30640 6365 30680
rect 7306 30640 7315 30680
rect 7355 30640 7468 30680
rect 7508 30640 7517 30680
rect 7747 30640 7756 30680
rect 7796 30640 7852 30680
rect 7892 30640 8188 30680
rect 8228 30640 8237 30680
rect 8297 30640 8428 30680
rect 8468 30640 8477 30680
rect 6604 30596 6644 30605
rect 9868 30596 9908 30808
rect 10697 30724 10828 30764
rect 10868 30724 10877 30764
rect 13638 30680 13728 30700
rect 10409 30640 10444 30680
rect 10484 30640 10540 30680
rect 10580 30640 10589 30680
rect 10915 30640 10924 30680
rect 10964 30640 11020 30680
rect 11060 30640 11095 30680
rect 11395 30640 11404 30680
rect 11444 30640 11596 30680
rect 11636 30640 11645 30680
rect 11875 30640 11884 30680
rect 11924 30640 11933 30680
rect 12259 30640 12268 30680
rect 12308 30640 12364 30680
rect 12404 30640 12439 30680
rect 13027 30640 13036 30680
rect 13076 30640 13728 30680
rect 11884 30596 11924 30640
rect 13638 30620 13728 30640
rect 3811 30556 3820 30596
rect 3860 30556 4012 30596
rect 4052 30556 4061 30596
rect 4937 30556 5068 30596
rect 5108 30556 5117 30596
rect 5260 30556 5539 30596
rect 5579 30556 5588 30596
rect 5635 30556 5644 30596
rect 5684 30556 5693 30596
rect 6115 30556 6124 30596
rect 6164 30556 6173 30596
rect 6473 30556 6604 30596
rect 6644 30556 6653 30596
rect 7114 30556 7123 30596
rect 7163 30556 7468 30596
rect 7508 30556 7517 30596
rect 8489 30556 8620 30596
rect 8660 30556 9292 30596
rect 9332 30556 9341 30596
rect 11299 30556 11308 30596
rect 11348 30556 11924 30596
rect 5068 30547 5108 30556
rect 5260 30512 5300 30556
rect 3139 30472 3148 30512
rect 3188 30472 3197 30512
rect 4444 30472 4876 30512
rect 4916 30472 4925 30512
rect 5251 30472 5260 30512
rect 5300 30472 5309 30512
rect 4444 30428 4484 30472
rect 6124 30428 6164 30556
rect 6604 30547 6644 30556
rect 9868 30512 9908 30556
rect 7564 30472 9908 30512
rect 10051 30472 10060 30512
rect 10100 30472 10156 30512
rect 10196 30472 10231 30512
rect 12115 30472 12124 30512
rect 12164 30472 12748 30512
rect 12788 30472 12797 30512
rect 7564 30428 7604 30472
rect 4099 30388 4108 30428
rect 4148 30388 4157 30428
rect 4396 30388 4484 30428
rect 4579 30388 4588 30428
rect 4628 30388 6164 30428
rect 6403 30388 6412 30428
rect 6452 30388 7604 30428
rect 7699 30388 7708 30428
rect 7748 30388 8044 30428
rect 8084 30388 8093 30428
rect 10156 30388 10204 30428
rect 10244 30388 10253 30428
rect 11251 30388 11260 30428
rect 11300 30388 11884 30428
rect 11924 30388 11933 30428
rect 12499 30388 12508 30428
rect 12548 30388 13036 30428
rect 13076 30388 13085 30428
rect 1795 30304 1804 30344
rect 1844 30304 2900 30344
rect 2860 30176 2900 30304
rect 4108 30176 4148 30388
rect 2860 30136 4148 30176
rect 4396 30176 4436 30388
rect 10156 30344 10196 30388
rect 13638 30344 13728 30364
rect 5731 30304 5740 30344
rect 5780 30304 10196 30344
rect 12259 30304 12268 30344
rect 12308 30304 13728 30344
rect 13638 30284 13728 30304
rect 4771 30220 4780 30260
rect 4820 30220 4868 30260
rect 4919 30220 4928 30260
rect 4968 30220 5010 30260
rect 5050 30220 5092 30260
rect 5132 30220 5174 30260
rect 5214 30220 5256 30260
rect 5296 30220 5305 30260
rect 5356 30220 6644 30260
rect 10819 30220 10828 30260
rect 10868 30220 10877 30260
rect 4828 30176 4868 30220
rect 5356 30176 5396 30220
rect 6604 30176 6644 30220
rect 10828 30176 10868 30220
rect 4396 30136 4532 30176
rect 4828 30136 4916 30176
rect 4492 30008 4532 30136
rect 4876 30092 4916 30136
rect 5164 30136 5396 30176
rect 6595 30136 6604 30176
rect 6644 30136 9100 30176
rect 9140 30136 9149 30176
rect 10723 30136 10732 30176
rect 10772 30136 10781 30176
rect 10828 30136 10924 30176
rect 10964 30136 10973 30176
rect 4867 30052 4876 30092
rect 4916 30052 4925 30092
rect 4300 29968 4532 30008
rect 4300 29924 4340 29968
rect 4012 29884 4078 29924
rect 4118 29884 4127 29924
rect 4195 29884 4204 29924
rect 4244 29884 4340 29924
rect 4579 29884 4588 29924
rect 4628 29884 4972 29924
rect 5012 29884 5021 29924
rect 5164 29915 5204 30136
rect 7337 30052 7468 30092
rect 7508 30052 7517 30092
rect 8275 30052 8284 30092
rect 8324 30052 9524 30092
rect 9484 30008 9524 30052
rect 10108 30052 10252 30092
rect 10292 30052 10301 30092
rect 10108 30008 10148 30052
rect 10732 30008 10772 30136
rect 13638 30008 13728 30028
rect 5347 29968 5356 30008
rect 5396 29968 5740 30008
rect 5780 29968 6068 30008
rect 7891 29968 7900 30008
rect 7940 29968 9388 30008
rect 9428 29968 9437 30008
rect 9484 29968 10148 30008
rect 10204 29968 10444 30008
rect 10484 29968 10493 30008
rect 10723 29968 10732 30008
rect 10772 29968 10781 30008
rect 12547 29968 12556 30008
rect 12596 29968 13728 30008
rect 6028 29924 6068 29968
rect 10204 29924 10244 29968
rect 13638 29948 13728 29968
rect 4012 29840 4052 29884
rect 5513 29884 5644 29924
rect 5684 29884 5693 29924
rect 6019 29884 6028 29924
rect 6068 29884 6077 29924
rect 7276 29915 7756 29924
rect 5164 29866 5204 29875
rect 5644 29866 5684 29875
rect 7316 29884 7756 29915
rect 7796 29884 7805 29924
rect 7852 29884 8332 29924
rect 8372 29884 8381 29924
rect 10147 29884 10156 29924
rect 10196 29884 10244 29924
rect 10522 29884 10531 29924
rect 10571 29884 10924 29924
rect 10964 29884 10973 29924
rect 7276 29866 7316 29875
rect 7852 29840 7892 29884
rect 67 29800 76 29840
rect 116 29800 1228 29840
rect 1268 29800 1277 29840
rect 4012 29800 4108 29840
rect 4148 29800 4157 29840
rect 4483 29800 4492 29840
rect 4532 29800 4684 29840
rect 4724 29800 4733 29840
rect 7459 29800 7468 29840
rect 7508 29800 7660 29840
rect 7700 29800 7892 29840
rect 8035 29800 8044 29840
rect 8084 29800 8093 29840
rect 9257 29800 9388 29840
rect 9428 29800 9437 29840
rect 9641 29800 9772 29840
rect 9812 29800 9821 29840
rect 10003 29800 10012 29840
rect 10052 29800 10060 29840
rect 10100 29800 10183 29840
rect 10819 29800 10828 29840
rect 10868 29800 10877 29840
rect 8044 29756 8084 29800
rect 1027 29716 1036 29756
rect 1076 29716 1652 29756
rect 4003 29716 4012 29756
rect 4052 29716 7756 29756
rect 7796 29716 8084 29756
rect 9619 29716 9628 29756
rect 9668 29716 10292 29756
rect 0 29672 90 29692
rect 0 29632 76 29672
rect 116 29632 125 29672
rect 1459 29632 1468 29672
rect 1508 29632 1517 29672
rect 0 29612 90 29632
rect 1468 29420 1508 29632
rect 1612 29588 1652 29716
rect 10252 29672 10292 29716
rect 13638 29672 13728 29692
rect 5347 29632 5356 29672
rect 5396 29632 5875 29672
rect 5915 29632 5924 29672
rect 10252 29632 10484 29672
rect 10627 29632 10636 29672
rect 10676 29632 12460 29672
rect 12500 29632 12509 29672
rect 12556 29632 13728 29672
rect 10444 29588 10484 29632
rect 12556 29588 12596 29632
rect 13638 29612 13728 29632
rect 1612 29548 10100 29588
rect 10444 29548 12596 29588
rect 10060 29504 10100 29548
rect 2851 29464 2860 29504
rect 2900 29464 3052 29504
rect 3092 29464 3101 29504
rect 3679 29464 3688 29504
rect 3728 29464 3770 29504
rect 3810 29464 3852 29504
rect 3892 29464 3934 29504
rect 3974 29464 4016 29504
rect 4056 29464 4065 29504
rect 4963 29464 4972 29504
rect 5012 29464 6316 29504
rect 6356 29464 6365 29504
rect 10060 29464 10292 29504
rect 10252 29420 10292 29464
rect 1468 29380 10100 29420
rect 10147 29380 10156 29420
rect 10196 29380 10205 29420
rect 10252 29380 10924 29420
rect 10964 29380 10973 29420
rect 10060 29336 10100 29380
rect 10156 29336 10196 29380
rect 13638 29336 13728 29356
rect 1459 29296 1468 29336
rect 1508 29296 1996 29336
rect 2036 29296 2045 29336
rect 2563 29296 2572 29336
rect 2612 29296 2620 29336
rect 2660 29296 2743 29336
rect 4579 29296 4588 29336
rect 4628 29296 5644 29336
rect 5684 29296 5693 29336
rect 5971 29296 5980 29336
rect 6020 29296 6700 29336
rect 6740 29296 6749 29336
rect 10051 29296 10060 29336
rect 10100 29296 10109 29336
rect 10156 29296 13728 29336
rect 13638 29276 13728 29296
rect 5587 29212 5596 29252
rect 5636 29212 9388 29252
rect 9428 29212 9437 29252
rect 9571 29212 9580 29252
rect 9620 29212 12308 29252
rect 12268 29168 12308 29212
rect 67 29128 76 29168
rect 116 29128 1228 29168
rect 1268 29128 1277 29168
rect 2371 29128 2380 29168
rect 2420 29128 2860 29168
rect 2900 29128 2909 29168
rect 5225 29128 5356 29168
rect 5396 29128 5405 29168
rect 5609 29128 5740 29168
rect 5780 29128 6452 29168
rect 2860 29084 2900 29128
rect 4396 29084 4436 29093
rect 6412 29084 6452 29128
rect 7660 29128 8140 29168
rect 8180 29128 9100 29168
rect 9140 29128 9332 29168
rect 7660 29084 7700 29128
rect 9292 29084 9332 29128
rect 9868 29128 10156 29168
rect 10196 29128 10205 29168
rect 10339 29128 10348 29168
rect 10388 29128 10828 29168
rect 10868 29128 10877 29168
rect 11875 29128 11884 29168
rect 11924 29128 12212 29168
rect 12259 29128 12268 29168
rect 12308 29128 12317 29168
rect 9868 29084 9908 29128
rect 10923 29084 10963 29093
rect 12172 29084 12212 29128
rect 2860 29044 3148 29084
rect 3188 29044 3197 29084
rect 4265 29044 4396 29084
rect 4436 29044 4445 29084
rect 6403 29044 6412 29084
rect 6452 29044 6461 29084
rect 7747 29044 7756 29084
rect 7796 29044 8044 29084
rect 8084 29044 8093 29084
rect 9850 29044 9859 29084
rect 9899 29044 9908 29084
rect 9955 29044 9964 29084
rect 10004 29044 10013 29084
rect 10435 29044 10444 29084
rect 10484 29044 10580 29084
rect 10627 29044 10636 29084
rect 10676 29044 10923 29084
rect 11011 29044 11020 29084
rect 11060 29044 11412 29084
rect 11452 29044 11461 29084
rect 12163 29044 12172 29084
rect 12212 29044 12221 29084
rect 4396 29035 4436 29044
rect 7660 29035 7700 29044
rect 9292 29035 9332 29044
rect 9964 29000 10004 29044
rect 10540 29000 10580 29044
rect 10923 29035 10963 29044
rect 13638 29000 13728 29020
rect 9667 28960 9676 29000
rect 9716 28960 10004 29000
rect 10051 28960 10060 29000
rect 10100 28960 10580 29000
rect 11971 28960 11980 29000
rect 12020 28960 13728 29000
rect 10540 28916 10580 28960
rect 13638 28940 13728 28960
rect 7843 28876 7852 28916
rect 7892 28876 8620 28916
rect 8660 28876 8669 28916
rect 9475 28876 9484 28916
rect 9524 28876 10156 28916
rect 10196 28876 10205 28916
rect 10540 28876 11020 28916
rect 11060 28876 11069 28916
rect 11465 28876 11596 28916
rect 11636 28876 11645 28916
rect 12115 28876 12124 28916
rect 12164 28876 12364 28916
rect 12404 28876 12413 28916
rect 12499 28876 12508 28916
rect 12548 28876 13132 28916
rect 13172 28876 13181 28916
rect 6307 28792 6316 28832
rect 6356 28792 10060 28832
rect 10100 28792 10109 28832
rect 4919 28708 4928 28748
rect 4968 28708 5010 28748
rect 5050 28708 5092 28748
rect 5132 28708 5174 28748
rect 5214 28708 5256 28748
rect 5296 28708 5305 28748
rect 0 28664 90 28684
rect 13638 28664 13728 28684
rect 0 28624 76 28664
rect 116 28624 125 28664
rect 7267 28624 7276 28664
rect 7316 28624 10540 28664
rect 10580 28624 10589 28664
rect 11875 28624 11884 28664
rect 11924 28624 13728 28664
rect 0 28604 90 28624
rect 13638 28604 13728 28624
rect 1459 28540 1468 28580
rect 1508 28540 3436 28580
rect 3476 28540 3485 28580
rect 3977 28540 4012 28580
rect 4052 28540 4108 28580
rect 4148 28540 4157 28580
rect 8332 28540 8908 28580
rect 8948 28540 8957 28580
rect 10339 28540 10348 28580
rect 10388 28540 10397 28580
rect 2659 28456 2668 28496
rect 2708 28456 6932 28496
rect 6892 28412 6932 28456
rect 8332 28412 8372 28540
rect 10348 28496 10388 28540
rect 8573 28456 8620 28496
rect 8660 28456 8669 28496
rect 9379 28456 9388 28496
rect 9428 28456 9868 28496
rect 9908 28456 10292 28496
rect 10348 28456 11924 28496
rect 8620 28412 8660 28456
rect 2275 28372 2284 28412
rect 2324 28372 2476 28412
rect 2516 28372 2572 28412
rect 2612 28372 2621 28412
rect 3820 28403 4396 28412
rect 3860 28372 4396 28403
rect 4436 28372 4445 28412
rect 6883 28372 6892 28412
rect 6932 28372 6941 28412
rect 8140 28403 8372 28412
rect 3820 28354 3860 28363
rect 8180 28372 8372 28403
rect 8602 28372 8611 28412
rect 8651 28372 8660 28412
rect 8707 28372 8716 28412
rect 8756 28372 8765 28412
rect 9091 28372 9100 28412
rect 9140 28372 9580 28412
rect 9620 28372 9629 28412
rect 9676 28403 9716 28412
rect 8140 28354 8180 28363
rect 8716 28328 8756 28372
rect 10025 28372 10156 28412
rect 10196 28372 10205 28412
rect 9676 28328 9716 28363
rect 10156 28354 10196 28363
rect 10252 28328 10292 28456
rect 10409 28372 10540 28412
rect 10580 28372 11596 28412
rect 11636 28372 11645 28412
rect 11788 28403 11828 28412
rect 11788 28328 11828 28363
rect 1097 28288 1228 28328
rect 1268 28288 1277 28328
rect 8419 28288 8428 28328
rect 8468 28288 8756 28328
rect 9187 28288 9196 28328
rect 9236 28288 9245 28328
rect 9676 28288 10060 28328
rect 10100 28288 10109 28328
rect 10252 28288 11828 28328
rect 11884 28328 11924 28456
rect 13638 28328 13728 28348
rect 11884 28288 12364 28328
rect 12404 28288 12413 28328
rect 13315 28288 13324 28328
rect 13364 28288 13728 28328
rect 9196 28244 9236 28288
rect 13638 28268 13728 28288
rect 9196 28204 10924 28244
rect 10964 28204 10973 28244
rect 8323 28120 8332 28160
rect 8372 28120 8381 28160
rect 11849 28120 11980 28160
rect 12020 28120 12029 28160
rect 12115 28120 12124 28160
rect 12164 28120 12173 28160
rect 3679 27952 3688 27992
rect 3728 27952 3770 27992
rect 3810 27952 3852 27992
rect 3892 27952 3934 27992
rect 3974 27952 4016 27992
rect 4056 27952 4065 27992
rect 8332 27908 8372 28120
rect 12124 28076 12164 28120
rect 9475 28036 9484 28076
rect 9524 28036 12164 28076
rect 13638 27992 13728 28012
rect 13219 27952 13228 27992
rect 13268 27952 13728 27992
rect 13638 27932 13728 27952
rect 8332 27868 10004 27908
rect 9292 27700 9772 27740
rect 9812 27700 9821 27740
rect 0 27656 90 27676
rect 9292 27656 9332 27700
rect 0 27616 1228 27656
rect 1268 27616 1277 27656
rect 8044 27616 8908 27656
rect 8948 27616 8957 27656
rect 9283 27616 9292 27656
rect 9332 27616 9341 27656
rect 0 27596 90 27616
rect 5548 27572 5588 27581
rect 8044 27572 8084 27616
rect 4291 27532 4300 27572
rect 4340 27532 4588 27572
rect 4628 27532 4637 27572
rect 5417 27532 5548 27572
rect 5588 27532 5597 27572
rect 6691 27532 6700 27572
rect 6740 27532 6796 27572
rect 6836 27532 6871 27572
rect 5548 27523 5588 27532
rect 8044 27523 8084 27532
rect 8236 27532 8803 27572
rect 8843 27532 8852 27572
rect 8899 27532 8908 27572
rect 8948 27532 8957 27572
rect 8236 27488 8276 27532
rect 8227 27448 8236 27488
rect 8276 27448 8285 27488
rect 8908 27404 8948 27532
rect 9292 27488 9332 27616
rect 9868 27572 9908 27581
rect 9379 27532 9388 27572
rect 9428 27532 9772 27572
rect 9812 27532 9821 27572
rect 9964 27572 10004 27868
rect 10570 27784 10579 27824
rect 10619 27784 11884 27824
rect 11924 27784 11933 27824
rect 11587 27700 11596 27740
rect 11636 27700 11645 27740
rect 11596 27656 11636 27700
rect 13638 27656 13728 27676
rect 11596 27616 12212 27656
rect 12739 27616 12748 27656
rect 12788 27616 13728 27656
rect 10924 27572 10964 27581
rect 12172 27572 12212 27616
rect 13638 27596 13728 27616
rect 9964 27532 10356 27572
rect 10396 27532 10405 27572
rect 10964 27532 11596 27572
rect 11636 27532 11645 27572
rect 12163 27532 12172 27572
rect 12212 27532 12268 27572
rect 12308 27532 12372 27572
rect 9868 27488 9908 27532
rect 10924 27523 10964 27532
rect 9292 27448 9428 27488
rect 9868 27448 10252 27488
rect 10292 27448 10301 27488
rect 5731 27364 5740 27404
rect 5780 27364 5932 27404
rect 5972 27364 5981 27404
rect 8908 27364 9332 27404
rect 9292 27236 9332 27364
rect 9388 27320 9428 27448
rect 10601 27364 10732 27404
rect 10772 27364 10781 27404
rect 13638 27320 13728 27340
rect 9388 27280 10348 27320
rect 10388 27280 10397 27320
rect 13027 27280 13036 27320
rect 13076 27280 13728 27320
rect 13638 27260 13728 27280
rect 4919 27196 4928 27236
rect 4968 27196 5010 27236
rect 5050 27196 5092 27236
rect 5132 27196 5174 27236
rect 5214 27196 5256 27236
rect 5296 27196 5305 27236
rect 9292 27196 10060 27236
rect 10100 27196 10109 27236
rect 11683 27196 11692 27236
rect 11732 27196 11884 27236
rect 11924 27196 11933 27236
rect 1468 27112 8716 27152
rect 8756 27112 8765 27152
rect 8812 27112 13324 27152
rect 13364 27112 13373 27152
rect 1468 27068 1508 27112
rect 1459 27028 1468 27068
rect 1508 27028 1517 27068
rect 3916 27028 5548 27068
rect 5588 27028 5597 27068
rect 6547 27028 6556 27068
rect 6596 27028 6988 27068
rect 7028 27028 7037 27068
rect 2537 26860 2668 26900
rect 2708 26860 3436 26900
rect 3476 26860 3485 26900
rect 3916 26891 3956 27028
rect 8812 26984 8852 27112
rect 11491 27028 11500 27068
rect 11540 27028 12028 27068
rect 12068 27028 12077 27068
rect 13638 26984 13728 27004
rect 4099 26944 4108 26984
rect 4148 26944 4436 26984
rect 4396 26900 4436 26944
rect 6028 26944 8852 26984
rect 9667 26944 9676 26984
rect 9716 26944 12116 26984
rect 12355 26944 12364 26984
rect 12404 26944 13728 26984
rect 4378 26860 4387 26900
rect 4427 26860 4436 26900
rect 4483 26860 4492 26900
rect 4532 26860 4541 26900
rect 4675 26860 4684 26900
rect 4724 26860 4876 26900
rect 4916 26860 4925 26900
rect 5452 26891 5548 26900
rect 3916 26842 3956 26851
rect 4492 26816 4532 26860
rect 5492 26860 5548 26891
rect 5588 26860 5623 26900
rect 5801 26860 5932 26900
rect 5972 26860 5981 26900
rect 5452 26842 5492 26851
rect 5932 26842 5972 26851
rect 1219 26776 1228 26816
rect 1268 26776 1277 26816
rect 4291 26776 4300 26816
rect 4340 26776 4532 26816
rect 4841 26776 4972 26816
rect 5012 26776 5021 26816
rect 0 26648 90 26668
rect 1228 26648 1268 26776
rect 0 26608 1268 26648
rect 0 26588 90 26608
rect 3679 26440 3688 26480
rect 3728 26440 3770 26480
rect 3810 26440 3852 26480
rect 3892 26440 3934 26480
rect 3974 26440 4016 26480
rect 4056 26440 4065 26480
rect 6028 26312 6068 26944
rect 10252 26900 10292 26944
rect 12076 26900 12116 26944
rect 13638 26924 13728 26944
rect 6403 26860 6412 26900
rect 6452 26860 6796 26900
rect 6836 26860 7223 26900
rect 7263 26860 7272 26900
rect 7459 26860 7468 26900
rect 7508 26860 7756 26900
rect 7796 26860 7805 26900
rect 9754 26860 9763 26900
rect 9803 26860 9812 26900
rect 9859 26860 9868 26900
rect 9908 26860 10004 26900
rect 10243 26860 10252 26900
rect 10292 26860 10301 26900
rect 10828 26891 11020 26900
rect 9772 26816 9812 26860
rect 6154 26776 6163 26816
rect 6203 26776 6316 26816
rect 6356 26776 6365 26816
rect 7267 26776 7276 26816
rect 7316 26776 7363 26816
rect 7403 26776 7447 26816
rect 7555 26776 7564 26816
rect 7604 26776 8140 26816
rect 8180 26776 8189 26816
rect 9763 26776 9772 26816
rect 9812 26776 9859 26816
rect 9964 26732 10004 26860
rect 10868 26860 11020 26891
rect 11060 26860 11069 26900
rect 11308 26891 11980 26900
rect 10828 26842 10868 26851
rect 10339 26776 10348 26816
rect 10388 26776 10397 26816
rect 8620 26692 10004 26732
rect 10348 26732 10388 26776
rect 11020 26732 11060 26860
rect 11348 26860 11980 26891
rect 12020 26860 12029 26900
rect 12076 26860 13324 26900
rect 13364 26860 13373 26900
rect 11308 26842 11348 26851
rect 11561 26776 11692 26816
rect 11732 26776 11741 26816
rect 11875 26776 11884 26816
rect 11924 26776 12268 26816
rect 12308 26776 12317 26816
rect 10348 26692 10924 26732
rect 10964 26692 10973 26732
rect 11020 26692 13228 26732
rect 13268 26692 13277 26732
rect 6979 26356 6988 26396
rect 7028 26356 7660 26396
rect 7700 26356 8524 26396
rect 8564 26356 8573 26396
rect 8620 26312 8660 26692
rect 13638 26648 13728 26668
rect 11530 26608 11539 26648
rect 11579 26608 11828 26648
rect 11923 26608 11932 26648
rect 11972 26608 12308 26648
rect 13123 26608 13132 26648
rect 13172 26608 13728 26648
rect 11788 26564 11828 26608
rect 11788 26524 12116 26564
rect 10339 26356 10348 26396
rect 10388 26356 10484 26396
rect 4723 26272 4732 26312
rect 4772 26272 6068 26312
rect 6307 26272 6316 26312
rect 6356 26272 8660 26312
rect 4457 26188 4588 26228
rect 4628 26188 6644 26228
rect 6691 26188 6700 26228
rect 6740 26188 7276 26228
rect 7316 26188 8372 26228
rect 4492 26144 4532 26188
rect 6604 26144 6644 26188
rect 4483 26104 4492 26144
rect 4532 26104 4541 26144
rect 6604 26104 6700 26144
rect 6740 26104 6749 26144
rect 1420 26060 1460 26069
rect 3052 26060 3092 26069
rect 6508 26060 6548 26069
rect 8140 26060 8180 26069
rect 8332 26060 8372 26188
rect 8620 26102 8660 26272
rect 10444 26228 10484 26356
rect 11722 26272 11731 26312
rect 11771 26272 11884 26312
rect 11924 26272 11933 26312
rect 10051 26188 10060 26228
rect 10100 26188 10340 26228
rect 8620 26093 8703 26102
rect 8620 26062 8663 26093
rect 2467 26020 2476 26060
rect 2516 26020 2668 26060
rect 2708 26020 2717 26060
rect 2860 26020 3052 26060
rect 4099 26020 4108 26060
rect 4148 26020 4300 26060
rect 4340 26020 4349 26060
rect 5251 26020 5260 26060
rect 5300 26020 5644 26060
rect 5684 26020 5693 26060
rect 6857 26020 6892 26060
rect 6932 26020 6988 26060
rect 7028 26020 7037 26060
rect 7651 26020 7660 26060
rect 7700 26020 8140 26060
rect 8323 26020 8332 26060
rect 8372 26020 8524 26060
rect 8564 26020 8573 26060
rect 10300 26060 10340 26188
rect 10444 26188 11404 26228
rect 11444 26188 11453 26228
rect 10444 26144 10484 26188
rect 12076 26144 12116 26524
rect 12268 26144 12308 26608
rect 13638 26588 13728 26608
rect 13638 26312 13728 26332
rect 13027 26272 13036 26312
rect 13076 26272 13728 26312
rect 13638 26252 13728 26272
rect 10435 26104 10444 26144
rect 10484 26104 10493 26144
rect 12067 26104 12076 26144
rect 12116 26104 12125 26144
rect 12259 26104 12268 26144
rect 12308 26104 12317 26144
rect 8663 26044 8703 26053
rect 9946 26020 9955 26060
rect 9995 26020 10004 26060
rect 10051 26020 10060 26060
rect 10100 26020 10231 26060
rect 10300 26020 10540 26060
rect 10580 26020 10589 26060
rect 11006 26020 11015 26060
rect 11055 26020 11064 26060
rect 11530 26020 11539 26060
rect 11579 26020 12076 26060
rect 12116 26020 12125 26060
rect 1420 25976 1460 26020
rect 2860 25976 2900 26020
rect 3052 26011 3092 26020
rect 1097 25936 1228 25976
rect 1268 25936 1277 25976
rect 1420 25936 2668 25976
rect 2708 25936 2900 25976
rect 6508 25976 6548 26020
rect 7660 25976 7700 26020
rect 8140 26011 8180 26020
rect 9964 25976 10004 26020
rect 6508 25936 7700 25976
rect 8323 25936 8332 25976
rect 8372 25936 8716 25976
rect 8756 25936 8765 25976
rect 9964 25936 10732 25976
rect 10772 25936 10781 25976
rect 11020 25892 11060 26020
rect 13638 25976 13728 25996
rect 11827 25936 11836 25976
rect 11876 25936 11884 25976
rect 11924 25936 12007 25976
rect 13123 25936 13132 25976
rect 13172 25936 13728 25976
rect 13638 25916 13728 25936
rect 2851 25852 2860 25892
rect 2900 25852 2956 25892
rect 2996 25852 3031 25892
rect 8611 25852 8620 25892
rect 8660 25852 8812 25892
rect 8852 25852 8861 25892
rect 10243 25852 10252 25892
rect 10292 25852 11060 25892
rect 12499 25852 12508 25892
rect 12548 25852 12557 25892
rect 4919 25684 4928 25724
rect 4968 25684 5010 25724
rect 5050 25684 5092 25724
rect 5132 25684 5174 25724
rect 5214 25684 5256 25724
rect 5296 25684 5305 25724
rect 0 25640 90 25660
rect 12508 25640 12548 25852
rect 13638 25640 13728 25660
rect 0 25580 116 25640
rect 76 25472 116 25580
rect 2860 25600 9292 25640
rect 9332 25600 9341 25640
rect 12508 25600 13728 25640
rect 2860 25556 2900 25600
rect 13638 25580 13728 25600
rect 1459 25516 1468 25556
rect 1508 25516 2900 25556
rect 8026 25516 8035 25556
rect 8075 25516 9236 25556
rect 9641 25516 9772 25556
rect 9812 25516 9821 25556
rect 12499 25516 12508 25556
rect 12548 25516 13132 25556
rect 13172 25516 13181 25556
rect 25 25432 116 25472
rect 6316 25432 7468 25472
rect 7508 25432 7517 25472
rect 8332 25432 8803 25472
rect 8843 25432 8852 25472
rect 25 25304 65 25432
rect 6316 25388 6356 25432
rect 8332 25388 8372 25432
rect 9196 25388 9236 25516
rect 2659 25348 2668 25388
rect 2708 25379 2996 25388
rect 2708 25348 2956 25379
rect 4099 25348 4108 25388
rect 4148 25348 4204 25388
rect 4244 25348 4279 25388
rect 4675 25348 4684 25388
rect 4724 25348 5644 25388
rect 5684 25348 5693 25388
rect 5932 25379 5972 25388
rect 2956 25330 2996 25339
rect 6307 25348 6316 25388
rect 6356 25348 6365 25388
rect 7529 25379 7660 25388
rect 7529 25348 7564 25379
rect 25 25264 1228 25304
rect 1268 25264 1277 25304
rect 1603 25264 1612 25304
rect 1652 25264 1661 25304
rect 1612 25136 1652 25264
rect 25 25096 1652 25136
rect 1843 25096 1852 25136
rect 1892 25096 2284 25136
rect 2324 25096 2333 25136
rect 2563 25096 2572 25136
rect 2612 25096 2764 25136
rect 2804 25096 2813 25136
rect 25 24800 65 25096
rect 5932 25052 5972 25339
rect 7604 25348 7660 25379
rect 7700 25348 7709 25388
rect 8057 25348 8140 25388
rect 8180 25348 8188 25388
rect 8228 25348 8237 25388
rect 8323 25348 8332 25388
rect 8372 25348 8381 25388
rect 8707 25348 8716 25388
rect 8756 25348 8951 25388
rect 8991 25348 9000 25388
rect 9187 25348 9196 25388
rect 9236 25348 9245 25388
rect 9379 25348 9388 25388
rect 9428 25348 9580 25388
rect 9620 25379 10004 25388
rect 9620 25348 9964 25379
rect 7564 25330 7604 25339
rect 8428 25306 8476 25346
rect 8516 25306 8525 25346
rect 11177 25348 11212 25388
rect 11252 25348 11308 25388
rect 11348 25348 11357 25388
rect 11884 25348 12364 25388
rect 12404 25348 12413 25388
rect 9964 25330 10004 25339
rect 8428 25304 8468 25306
rect 11884 25304 11924 25348
rect 13638 25304 13728 25324
rect 7756 25264 8468 25304
rect 8602 25264 8611 25304
rect 8651 25264 8660 25304
rect 8969 25264 9091 25304
rect 9140 25264 9149 25304
rect 9283 25264 9292 25304
rect 9332 25264 9463 25304
rect 11491 25264 11500 25304
rect 11540 25264 11549 25304
rect 11875 25264 11884 25304
rect 11924 25264 11933 25304
rect 11980 25264 12268 25304
rect 12308 25264 12317 25304
rect 12940 25264 13728 25304
rect 7756 25136 7796 25264
rect 8620 25220 8660 25264
rect 11500 25220 11540 25264
rect 11980 25220 12020 25264
rect 12940 25220 12980 25264
rect 13638 25244 13728 25264
rect 8573 25180 8620 25220
rect 8660 25180 8669 25220
rect 9763 25180 9772 25220
rect 9812 25180 11540 25220
rect 11596 25180 12020 25220
rect 12115 25180 12124 25220
rect 12164 25180 12980 25220
rect 11596 25136 11636 25180
rect 6115 25096 6124 25136
rect 6164 25096 7468 25136
rect 7508 25096 7517 25136
rect 7625 25096 7756 25136
rect 7796 25096 7805 25136
rect 11107 25096 11116 25136
rect 11156 25096 11636 25136
rect 11731 25096 11740 25136
rect 11780 25096 12404 25136
rect 5932 25012 8236 25052
rect 8276 25012 8285 25052
rect 12364 24968 12404 25096
rect 13638 24968 13728 24988
rect 3679 24928 3688 24968
rect 3728 24928 3770 24968
rect 3810 24928 3852 24968
rect 3892 24928 3934 24968
rect 3974 24928 4016 24968
rect 4056 24928 4065 24968
rect 12364 24928 13728 24968
rect 13638 24908 13728 24928
rect 7180 24844 9676 24884
rect 9716 24844 9725 24884
rect 7180 24800 7220 24844
rect 25 24760 116 24800
rect 4723 24760 4732 24800
rect 4772 24760 7220 24800
rect 8650 24760 8659 24800
rect 8699 24760 9100 24800
rect 9140 24760 9149 24800
rect 11945 24760 12076 24800
rect 12116 24760 12125 24800
rect 12499 24760 12508 24800
rect 12548 24760 13036 24800
rect 13076 24760 13085 24800
rect 76 24652 116 24760
rect 0 24592 116 24652
rect 6892 24676 7756 24716
rect 7796 24676 7805 24716
rect 8035 24676 8044 24716
rect 8084 24676 12308 24716
rect 2057 24592 2092 24632
rect 2132 24592 2179 24632
rect 2219 24592 2237 24632
rect 4099 24592 4108 24632
rect 4148 24592 4492 24632
rect 4532 24592 4541 24632
rect 0 24572 90 24592
rect 2380 24548 2420 24557
rect 6892 24548 6932 24676
rect 12268 24632 12308 24676
rect 13638 24632 13728 24652
rect 7241 24592 7276 24632
rect 7316 24592 7372 24632
rect 7412 24592 7421 24632
rect 8227 24592 8236 24632
rect 8276 24592 10100 24632
rect 12259 24592 12268 24632
rect 12308 24592 12317 24632
rect 12451 24592 12460 24632
rect 12500 24592 13728 24632
rect 7948 24548 7988 24557
rect 10060 24548 10100 24592
rect 13638 24572 13728 24592
rect 11884 24548 11924 24557
rect 2420 24508 2668 24548
rect 2708 24508 2717 24548
rect 3139 24508 3148 24548
rect 3188 24508 3628 24548
rect 3668 24508 3677 24548
rect 6874 24508 6883 24548
rect 6923 24508 6932 24548
rect 6979 24508 6988 24548
rect 7028 24508 7180 24548
rect 7220 24508 7229 24548
rect 7459 24508 7468 24548
rect 7508 24508 7517 24548
rect 7817 24508 7948 24548
rect 7988 24508 7997 24548
rect 8314 24508 8332 24548
rect 8372 24508 8436 24548
rect 8476 24508 8494 24548
rect 8611 24508 8620 24548
rect 8660 24508 8812 24548
rect 8852 24508 8861 24548
rect 10627 24508 10636 24548
rect 10676 24508 11308 24548
rect 11348 24508 11357 24548
rect 11587 24508 11596 24548
rect 11636 24508 11884 24548
rect 2380 24499 2420 24508
rect 7468 24464 7508 24508
rect 7948 24499 7988 24508
rect 10060 24499 10100 24508
rect 11884 24499 11924 24508
rect 6595 24424 6604 24464
rect 6644 24424 7508 24464
rect 10121 24340 10252 24380
rect 10292 24340 10301 24380
rect 13638 24296 13728 24316
rect 12835 24256 12844 24296
rect 12884 24256 13728 24296
rect 13638 24236 13728 24256
rect 4919 24172 4928 24212
rect 4968 24172 5010 24212
rect 5050 24172 5092 24212
rect 5132 24172 5174 24212
rect 5214 24172 5256 24212
rect 5296 24172 5305 24212
rect 5539 24004 5548 24044
rect 5588 24004 8948 24044
rect 9955 24004 9964 24044
rect 10004 24004 10012 24044
rect 10052 24004 10135 24044
rect 10675 24004 10684 24044
rect 10724 24004 12460 24044
rect 12500 24004 12509 24044
rect 8908 23960 8948 24004
rect 13638 23960 13728 23980
rect 4003 23920 4012 23960
rect 4052 23920 5780 23960
rect 5740 23876 5780 23920
rect 8908 23920 10348 23960
rect 10388 23920 10397 23960
rect 11491 23920 11500 23960
rect 11540 23920 13728 23960
rect 3977 23836 4108 23876
rect 4148 23836 4157 23876
rect 4963 23836 4972 23876
rect 5012 23867 5396 23876
rect 5012 23836 5356 23867
rect 5731 23836 5740 23876
rect 5780 23836 5789 23876
rect 6988 23867 7028 23876
rect 5356 23792 5396 23827
rect 7459 23836 7468 23876
rect 7508 23836 7843 23876
rect 7883 23836 7892 23876
rect 7939 23836 7948 23876
rect 7988 23836 7997 23876
rect 8201 23836 8332 23876
rect 8372 23836 8381 23876
rect 8908 23867 8948 23920
rect 13638 23900 13728 23920
rect 1219 23752 1228 23792
rect 1268 23752 1277 23792
rect 5356 23752 5740 23792
rect 5780 23752 5789 23792
rect 0 23624 90 23644
rect 1228 23624 1268 23752
rect 6988 23708 7028 23827
rect 7948 23792 7988 23836
rect 8908 23818 8948 23827
rect 9388 23867 10252 23876
rect 9428 23836 10252 23867
rect 10292 23836 10301 23876
rect 10889 23836 11020 23876
rect 11060 23836 11069 23876
rect 11299 23836 11308 23876
rect 11348 23836 12268 23876
rect 12308 23836 12317 23876
rect 9388 23818 9428 23827
rect 11020 23818 11060 23827
rect 7747 23752 7756 23792
rect 7796 23752 7988 23792
rect 8131 23752 8140 23792
rect 8180 23752 8428 23792
rect 8468 23752 8524 23792
rect 8564 23752 8573 23792
rect 9610 23752 9619 23792
rect 9659 23752 9772 23792
rect 9812 23752 9821 23792
rect 10051 23752 10060 23792
rect 10100 23752 10444 23792
rect 10484 23752 10493 23792
rect 2860 23668 4244 23708
rect 6988 23668 9100 23708
rect 9140 23668 9149 23708
rect 0 23584 1268 23624
rect 1459 23584 1468 23624
rect 1508 23584 1517 23624
rect 0 23564 90 23584
rect 1468 23540 1508 23584
rect 2860 23540 2900 23668
rect 4003 23584 4012 23624
rect 4052 23584 4061 23624
rect 1468 23500 2900 23540
rect 4012 23540 4052 23584
rect 4204 23540 4244 23668
rect 13638 23624 13728 23644
rect 5539 23584 5548 23624
rect 5588 23584 5740 23624
rect 5780 23584 5789 23624
rect 7049 23584 7180 23624
rect 7220 23584 7229 23624
rect 10819 23584 10828 23624
rect 10868 23584 10999 23624
rect 12163 23584 12172 23624
rect 12212 23584 13728 23624
rect 13638 23564 13728 23584
rect 4012 23500 4148 23540
rect 4204 23500 9388 23540
rect 9428 23500 9437 23540
rect 3679 23416 3688 23456
rect 3728 23416 3770 23456
rect 3810 23416 3852 23456
rect 3892 23416 3934 23456
rect 3974 23416 4016 23456
rect 4056 23416 4065 23456
rect 2659 23332 2668 23372
rect 2708 23332 2900 23372
rect 2860 23288 2900 23332
rect 4108 23288 4148 23500
rect 13315 23416 13324 23456
rect 13364 23416 13556 23456
rect 13516 23372 13556 23416
rect 2860 23248 3860 23288
rect 3907 23248 3916 23288
rect 3956 23248 4148 23288
rect 4300 23332 7604 23372
rect 13507 23332 13516 23372
rect 13556 23332 13565 23372
rect 3820 23204 3860 23248
rect 4300 23204 4340 23332
rect 7564 23288 7604 23332
rect 13638 23288 13728 23308
rect 6211 23248 6220 23288
rect 6260 23248 6364 23288
rect 6404 23248 6413 23288
rect 7564 23248 9820 23288
rect 9860 23248 10060 23288
rect 10100 23248 10109 23288
rect 10195 23248 10204 23288
rect 10244 23248 10348 23288
rect 10388 23248 10397 23288
rect 10444 23248 13728 23288
rect 10444 23204 10484 23248
rect 13638 23228 13728 23248
rect 3820 23164 4340 23204
rect 4483 23164 4492 23204
rect 4532 23164 5644 23204
rect 5684 23164 5693 23204
rect 8236 23164 8332 23204
rect 8372 23164 8381 23204
rect 9427 23164 9436 23204
rect 9476 23164 10388 23204
rect 10435 23164 10444 23204
rect 10484 23164 10493 23204
rect 10697 23164 10828 23204
rect 10868 23164 10877 23204
rect 25 23080 1228 23120
rect 1268 23080 1277 23120
rect 1459 23080 1468 23120
rect 1508 23080 1804 23120
rect 1844 23080 1853 23120
rect 4553 23080 4684 23120
rect 4724 23080 4733 23120
rect 25 22868 65 23080
rect 3724 23036 3764 23045
rect 4780 23036 4820 23164
rect 5962 23080 5971 23120
rect 6011 23080 6124 23120
rect 6164 23080 6173 23120
rect 7747 23080 7756 23120
rect 7796 23080 8140 23120
rect 8180 23080 8189 23120
rect 5260 23036 5300 23045
rect 8236 23036 8276 23164
rect 10348 23120 10388 23164
rect 8995 23080 9004 23120
rect 9044 23080 9580 23120
rect 9620 23080 9629 23120
rect 9955 23080 9964 23120
rect 10004 23080 10135 23120
rect 10339 23080 10348 23120
rect 10388 23080 10397 23120
rect 10531 23080 10540 23120
rect 10580 23080 10588 23120
rect 10628 23080 10711 23120
rect 8716 23036 8756 23045
rect 11020 23036 11060 23045
rect 2179 22996 2188 23036
rect 2228 22996 2476 23036
rect 2516 22996 2525 23036
rect 4043 22996 4108 23036
rect 4148 22996 4174 23036
rect 4214 22996 4223 23036
rect 4289 22996 4298 23036
rect 4340 22996 4469 23036
rect 4771 22996 4780 23036
rect 4820 22996 4829 23036
rect 5129 22996 5260 23036
rect 5300 22996 5309 23036
rect 5731 22996 5740 23036
rect 5788 22996 5911 23036
rect 7363 22996 7372 23036
rect 7412 22996 7651 23036
rect 7691 22996 7700 23036
rect 7747 22996 7756 23036
rect 7796 22996 7805 23036
rect 8035 22996 8044 23036
rect 8084 22996 8236 23036
rect 8276 22996 8285 23036
rect 9187 22996 9196 23036
rect 9244 22996 9367 23036
rect 10051 22996 10060 23036
rect 10100 22996 11020 23036
rect 11060 22996 11069 23036
rect 11203 22996 11212 23036
rect 11252 22996 12268 23036
rect 12308 22996 12317 23036
rect 3724 22952 3764 22996
rect 5260 22987 5300 22996
rect 7756 22952 7796 22996
rect 8716 22952 8756 22996
rect 11020 22987 11060 22996
rect 13638 22952 13728 22972
rect 3724 22912 5204 22952
rect 5443 22912 5452 22952
rect 5492 22912 7796 22952
rect 8611 22912 8620 22952
rect 8660 22912 8756 22952
rect 11587 22912 11596 22952
rect 11636 22912 13728 22952
rect 5164 22868 5204 22912
rect 13638 22892 13728 22912
rect 25 22828 76 22868
rect 116 22828 125 22868
rect 3907 22828 3916 22868
rect 3956 22828 3965 22868
rect 5164 22828 5740 22868
rect 5780 22828 6892 22868
rect 6932 22828 6941 22868
rect 0 22616 90 22636
rect 0 22576 76 22616
rect 116 22576 125 22616
rect 0 22556 90 22576
rect 3916 22448 3956 22828
rect 4919 22660 4928 22700
rect 4968 22660 5010 22700
rect 5050 22660 5092 22700
rect 5132 22660 5174 22700
rect 5214 22660 5256 22700
rect 5296 22660 5305 22700
rect 13638 22616 13728 22636
rect 9100 22576 9964 22616
rect 10004 22576 10013 22616
rect 10204 22576 13728 22616
rect 9100 22532 9140 22576
rect 10204 22532 10244 22576
rect 13638 22556 13728 22576
rect 9091 22492 9100 22532
rect 9140 22492 9149 22532
rect 9907 22492 9916 22532
rect 9956 22492 10244 22532
rect 10291 22492 10300 22532
rect 10340 22492 10444 22532
rect 10484 22492 10493 22532
rect 10675 22492 10684 22532
rect 10724 22492 11500 22532
rect 11540 22492 11549 22532
rect 3916 22408 4340 22448
rect 7123 22408 7132 22448
rect 7172 22408 12076 22448
rect 12116 22408 12125 22448
rect 4300 22364 4340 22408
rect 2851 22324 2860 22364
rect 2900 22324 4012 22364
rect 4052 22324 4061 22364
rect 4108 22355 4244 22364
rect 1097 22240 1228 22280
rect 1268 22240 1277 22280
rect 3148 22112 3188 22324
rect 4148 22324 4244 22355
rect 4300 22324 4579 22364
rect 4619 22324 4628 22364
rect 4675 22324 4684 22364
rect 4724 22324 4876 22364
rect 4916 22324 4925 22364
rect 5059 22324 5068 22364
rect 5108 22324 5117 22364
rect 5513 22324 5644 22364
rect 5684 22324 5693 22364
rect 5740 22355 6164 22364
rect 5740 22324 6124 22355
rect 4108 22306 4148 22315
rect 1459 22072 1468 22112
rect 1508 22072 2860 22112
rect 2900 22072 2909 22112
rect 3139 22072 3148 22112
rect 3188 22072 3197 22112
rect 4204 22028 4244 22324
rect 5068 22280 5108 22324
rect 5644 22306 5684 22315
rect 4579 22240 4588 22280
rect 4628 22240 5108 22280
rect 5155 22240 5164 22280
rect 5204 22240 5335 22280
rect 5740 22112 5780 22324
rect 7171 22324 7180 22364
rect 7220 22324 7363 22364
rect 7403 22324 7412 22364
rect 7459 22324 7468 22364
rect 7508 22324 7517 22364
rect 7843 22324 7852 22364
rect 7892 22324 8140 22364
rect 8180 22324 8189 22364
rect 8428 22355 8620 22364
rect 6124 22306 6164 22315
rect 7468 22280 7508 22324
rect 8468 22324 8620 22355
rect 8660 22324 8669 22364
rect 8777 22324 8908 22364
rect 8948 22324 8957 22364
rect 10889 22324 11020 22364
rect 11060 22324 11069 22364
rect 11299 22324 11308 22364
rect 11348 22324 12268 22364
rect 12308 22324 12317 22364
rect 8428 22306 8468 22315
rect 8908 22306 8948 22315
rect 11020 22306 11060 22315
rect 13638 22280 13728 22300
rect 6346 22240 6355 22280
rect 6395 22240 6508 22280
rect 6548 22240 6557 22280
rect 6761 22240 6892 22280
rect 6932 22240 6941 22280
rect 7267 22240 7276 22280
rect 7316 22240 7756 22280
rect 7796 22240 7805 22280
rect 7913 22240 7948 22280
rect 7988 22240 8044 22280
rect 8084 22240 8093 22280
rect 9161 22240 9196 22280
rect 9236 22240 9292 22280
rect 9332 22240 9341 22280
rect 9667 22240 9676 22280
rect 9716 22240 9868 22280
rect 9908 22240 9917 22280
rect 10051 22240 10060 22280
rect 10100 22240 10156 22280
rect 10196 22240 10231 22280
rect 10435 22240 10444 22280
rect 10484 22240 10636 22280
rect 10676 22240 10685 22280
rect 11596 22240 13728 22280
rect 11596 22196 11636 22240
rect 13638 22220 13728 22240
rect 6739 22156 6748 22196
rect 6788 22156 9292 22196
rect 9332 22156 9341 22196
rect 9523 22156 9532 22196
rect 9572 22156 11636 22196
rect 4291 22072 4300 22112
rect 4340 22072 5780 22112
rect 8035 22072 8044 22112
rect 8084 22072 10444 22112
rect 10484 22072 10493 22112
rect 10819 22072 10828 22112
rect 10868 22072 10877 22112
rect 4204 21988 9580 22028
rect 9620 21988 9629 22028
rect 3679 21904 3688 21944
rect 3728 21904 3770 21944
rect 3810 21904 3852 21944
rect 3892 21904 3934 21944
rect 3974 21904 4016 21944
rect 4056 21904 4065 21944
rect 10828 21860 10868 22072
rect 13638 21944 13728 21964
rect 11491 21904 11500 21944
rect 11540 21904 13728 21944
rect 13638 21884 13728 21904
rect 1603 21820 1612 21860
rect 1652 21820 10868 21860
rect 3977 21736 4108 21776
rect 4148 21736 4157 21776
rect 4867 21652 4876 21692
rect 4916 21652 7180 21692
rect 7220 21652 7229 21692
rect 8812 21652 9100 21692
rect 9140 21652 9149 21692
rect 10924 21652 11596 21692
rect 11636 21652 11645 21692
rect 0 21608 90 21628
rect 8812 21608 8852 21652
rect 10924 21608 10964 21652
rect 13638 21608 13728 21628
rect 0 21568 1228 21608
rect 1268 21568 1277 21608
rect 2179 21568 2188 21608
rect 2228 21568 2284 21608
rect 2324 21568 2708 21608
rect 4099 21568 4108 21608
rect 4148 21568 4396 21608
rect 4436 21568 4445 21608
rect 5347 21568 5356 21608
rect 5396 21568 5548 21608
rect 5588 21568 5597 21608
rect 5932 21568 6412 21608
rect 6452 21568 6461 21608
rect 8716 21568 8852 21608
rect 8899 21568 8908 21608
rect 8948 21568 8957 21608
rect 9161 21568 9292 21608
rect 9332 21568 9341 21608
rect 9667 21568 9676 21608
rect 9716 21568 9725 21608
rect 10243 21568 10252 21608
rect 10292 21568 10388 21608
rect 10435 21568 10444 21608
rect 10484 21568 10540 21608
rect 10580 21568 10615 21608
rect 10675 21568 10684 21608
rect 10724 21568 10964 21608
rect 11884 21568 13728 21608
rect 0 21548 90 21568
rect 2668 21524 2708 21568
rect 3916 21524 3956 21533
rect 5932 21524 5972 21568
rect 8044 21524 8084 21533
rect 8716 21524 8756 21568
rect 8908 21524 8948 21568
rect 2659 21484 2668 21524
rect 2708 21484 2717 21524
rect 3956 21484 4396 21524
rect 4436 21484 4445 21524
rect 4858 21484 4867 21524
rect 4907 21484 4916 21524
rect 4963 21484 4972 21524
rect 5012 21484 5143 21524
rect 5443 21484 5452 21524
rect 5492 21484 5876 21524
rect 3916 21475 3956 21484
rect 4876 21440 4916 21484
rect 2371 21400 2380 21440
rect 2420 21400 2524 21440
rect 2564 21400 2573 21440
rect 4204 21400 4916 21440
rect 3811 20980 3820 21020
rect 3860 20980 4108 21020
rect 4148 20980 4157 21020
rect 4204 20936 4244 21400
rect 5836 21356 5876 21484
rect 6442 21484 6451 21524
rect 6491 21484 6548 21524
rect 6665 21484 6796 21524
rect 6836 21484 6845 21524
rect 8084 21484 8716 21524
rect 8756 21484 8765 21524
rect 8908 21484 9484 21524
rect 9524 21484 9533 21524
rect 5932 21475 5972 21484
rect 4627 21316 4636 21356
rect 4676 21316 5396 21356
rect 5836 21316 6412 21356
rect 6452 21316 6461 21356
rect 4919 21148 4928 21188
rect 4968 21148 5010 21188
rect 5050 21148 5092 21188
rect 5132 21148 5174 21188
rect 5214 21148 5256 21188
rect 5296 21148 5305 21188
rect 5356 21104 5396 21316
rect 5356 21064 6404 21104
rect 3619 20896 3628 20936
rect 3668 20896 4244 20936
rect 6364 20936 6404 21064
rect 6508 21020 6548 21484
rect 8044 21475 8084 21484
rect 9676 21440 9716 21568
rect 10348 21524 10388 21568
rect 11020 21524 11060 21533
rect 10348 21484 10636 21524
rect 10676 21484 10685 21524
rect 10889 21484 11020 21524
rect 11060 21484 11069 21524
rect 11020 21475 11060 21484
rect 8227 21400 8236 21440
rect 8276 21400 8908 21440
rect 8948 21400 8957 21440
rect 9091 21400 9100 21440
rect 9140 21400 9716 21440
rect 9907 21400 9916 21440
rect 9956 21400 10964 21440
rect 10924 21356 10964 21400
rect 6595 21316 6604 21356
rect 6644 21316 6892 21356
rect 6932 21316 6941 21356
rect 9139 21316 9148 21356
rect 9188 21316 9476 21356
rect 9523 21316 9532 21356
rect 9572 21316 9581 21356
rect 10003 21316 10012 21356
rect 10052 21316 10060 21356
rect 10100 21316 10183 21356
rect 10697 21316 10828 21356
rect 10868 21316 10877 21356
rect 10924 21316 11500 21356
rect 11540 21316 11549 21356
rect 9436 21104 9476 21316
rect 9532 21272 9572 21316
rect 11884 21272 11924 21568
rect 13638 21548 13728 21568
rect 11971 21484 11980 21524
rect 12020 21484 12268 21524
rect 12308 21484 12317 21524
rect 13638 21272 13728 21292
rect 9532 21232 11924 21272
rect 13612 21212 13728 21272
rect 13612 21188 13652 21212
rect 12547 21148 12556 21188
rect 12596 21148 13652 21188
rect 6691 21064 6700 21104
rect 6740 21064 7948 21104
rect 7988 21064 7997 21104
rect 9436 21064 12308 21104
rect 6508 20980 7276 21020
rect 7316 20980 7325 21020
rect 8371 20980 8380 21020
rect 8420 20980 9004 21020
rect 9044 20980 9053 21020
rect 9580 20980 11924 21020
rect 12041 20980 12124 21020
rect 12164 20980 12172 21020
rect 12212 20980 12221 21020
rect 9580 20936 9620 20980
rect 6364 20896 9620 20936
rect 9667 20896 9676 20936
rect 9716 20896 11500 20936
rect 11540 20896 11549 20936
rect 11884 20852 11924 20980
rect 12268 20936 12308 21064
rect 12499 20980 12508 21020
rect 12548 20980 12844 21020
rect 12884 20980 12893 21020
rect 13638 20936 13728 20956
rect 12268 20896 13728 20936
rect 13638 20876 13728 20896
rect 2057 20812 2188 20852
rect 2228 20812 2237 20852
rect 3235 20812 3244 20852
rect 3284 20843 3476 20852
rect 3284 20812 3436 20843
rect 3994 20812 4003 20852
rect 4043 20812 4108 20852
rect 4148 20812 4183 20852
rect 4361 20812 4492 20852
rect 4532 20812 4541 20852
rect 4963 20812 4972 20852
rect 5012 20812 5143 20852
rect 5321 20812 5452 20852
rect 5492 20812 5501 20852
rect 5561 20812 5570 20852
rect 5610 20812 5644 20852
rect 5684 20812 5750 20852
rect 5827 20812 5836 20852
rect 5876 20812 5885 20852
rect 6403 20812 6412 20852
rect 6452 20812 6700 20852
rect 6740 20812 6749 20852
rect 7084 20843 8236 20852
rect 3436 20794 3476 20803
rect 4492 20794 4532 20803
rect 5836 20768 5876 20812
rect 7124 20812 8236 20843
rect 8276 20812 8285 20852
rect 8620 20812 9004 20852
rect 9044 20812 9053 20852
rect 9161 20812 9292 20852
rect 9332 20812 9341 20852
rect 9449 20812 9571 20852
rect 9620 20812 9629 20852
rect 10051 20812 10060 20852
rect 10100 20812 10109 20852
rect 10348 20843 10540 20852
rect 7084 20794 7124 20803
rect 8620 20768 8660 20812
rect 10060 20768 10100 20812
rect 10388 20812 10540 20843
rect 10580 20812 10589 20852
rect 11299 20812 11308 20852
rect 11348 20812 11596 20852
rect 11636 20812 11645 20852
rect 11884 20812 12308 20852
rect 10348 20794 10388 20803
rect 12268 20768 12308 20812
rect 67 20728 76 20768
rect 116 20728 1228 20768
rect 1268 20728 1277 20768
rect 4579 20728 4588 20768
rect 4628 20728 5068 20768
rect 5108 20728 5117 20768
rect 5740 20728 5876 20768
rect 7939 20728 7948 20768
rect 7988 20728 8380 20768
rect 8420 20728 8429 20768
rect 8611 20728 8620 20768
rect 8660 20728 8669 20768
rect 8716 20728 10100 20768
rect 11753 20728 11884 20768
rect 11924 20728 11933 20768
rect 12259 20728 12268 20768
rect 12308 20728 12317 20768
rect 5740 20684 5780 20728
rect 8716 20684 8756 20728
rect 3139 20644 3148 20684
rect 3188 20644 5780 20684
rect 5836 20644 8756 20684
rect 9955 20644 9964 20684
rect 10004 20644 10060 20684
rect 10100 20644 10135 20684
rect 0 20600 90 20620
rect 5836 20600 5876 20644
rect 13638 20600 13728 20620
rect 0 20560 76 20600
rect 116 20560 125 20600
rect 1459 20560 1468 20600
rect 1508 20560 1708 20600
rect 1748 20560 1757 20600
rect 4387 20560 4396 20600
rect 4436 20560 5876 20600
rect 7699 20560 7708 20600
rect 7748 20560 8716 20600
rect 8756 20560 8765 20600
rect 10025 20560 10156 20600
rect 10196 20560 10205 20600
rect 12067 20560 12076 20600
rect 12116 20560 13728 20600
rect 0 20540 90 20560
rect 13638 20540 13728 20560
rect 1987 20476 1996 20516
rect 2036 20476 10828 20516
rect 10868 20476 10877 20516
rect 3139 20392 3148 20432
rect 3188 20392 3197 20432
rect 3679 20392 3688 20432
rect 3728 20392 3770 20432
rect 3810 20392 3852 20432
rect 3892 20392 3934 20432
rect 3974 20392 4016 20432
rect 4056 20392 4065 20432
rect 4963 20392 4972 20432
rect 5012 20392 11308 20432
rect 11348 20392 11357 20432
rect 3148 20096 3188 20392
rect 9571 20308 9580 20348
rect 9620 20308 10828 20348
rect 10868 20308 10877 20348
rect 13638 20264 13728 20284
rect 3977 20224 4108 20264
rect 4148 20224 4157 20264
rect 9283 20224 9292 20264
rect 9332 20224 9388 20264
rect 9428 20224 9463 20264
rect 11587 20224 11596 20264
rect 11636 20224 13728 20264
rect 13638 20204 13728 20224
rect 3235 20140 3244 20180
rect 3284 20140 4628 20180
rect 9811 20140 9820 20180
rect 9860 20140 10340 20180
rect 4588 20096 4628 20140
rect 10300 20096 10340 20140
rect 10828 20140 11060 20180
rect 10828 20096 10868 20140
rect 11020 20096 11060 20140
rect 67 20056 76 20096
rect 116 20056 1228 20096
rect 1268 20056 1277 20096
rect 3148 20056 3284 20096
rect 4579 20056 4588 20096
rect 4628 20056 4637 20096
rect 5539 20056 5548 20096
rect 5588 20056 5740 20096
rect 5780 20056 6988 20096
rect 7028 20056 7037 20096
rect 7219 20056 7228 20096
rect 7268 20056 8908 20096
rect 8948 20056 8957 20096
rect 9571 20056 9580 20096
rect 9620 20056 9916 20096
rect 9956 20056 9965 20096
rect 10051 20056 10060 20096
rect 10100 20056 10156 20096
rect 10196 20056 10231 20096
rect 10300 20056 10868 20096
rect 10915 20056 10924 20096
rect 10964 20056 10973 20096
rect 11020 20056 11156 20096
rect 11369 20056 11500 20096
rect 11540 20056 13324 20096
rect 13364 20056 13373 20096
rect 3244 20012 3284 20056
rect 3916 20012 3956 20021
rect 9196 20012 9236 20021
rect 2467 19972 2476 20012
rect 2516 19972 2668 20012
rect 2708 19972 2717 20012
rect 3235 19972 3244 20012
rect 3284 19972 3293 20012
rect 3956 19972 4588 20012
rect 4628 19972 4637 20012
rect 7939 19972 7948 20012
rect 7988 19972 7997 20012
rect 8995 19972 9004 20012
rect 9044 19972 9196 20012
rect 9236 19972 9292 20012
rect 9332 19972 9341 20012
rect 10147 19972 10156 20012
rect 10196 19972 10435 20012
rect 10475 19972 10484 20012
rect 10531 19972 10540 20012
rect 10580 19972 10828 20012
rect 10868 19972 10877 20012
rect 3916 19963 3956 19972
rect 4588 19928 4628 19972
rect 4588 19888 5308 19928
rect 5348 19888 5357 19928
rect 1459 19804 1468 19844
rect 1508 19804 2284 19844
rect 2324 19804 2333 19844
rect 4387 19804 4396 19844
rect 4436 19804 4828 19844
rect 4868 19804 4877 19844
rect 4919 19636 4928 19676
rect 4968 19636 5010 19676
rect 5050 19636 5092 19676
rect 5132 19636 5174 19676
rect 5214 19636 5256 19676
rect 5296 19636 5305 19676
rect 0 19592 90 19612
rect 0 19552 76 19592
rect 116 19552 125 19592
rect 0 19532 90 19552
rect 1459 19468 1468 19508
rect 1508 19468 3244 19508
rect 3284 19468 3293 19508
rect 3619 19468 3628 19508
rect 3668 19468 5644 19508
rect 5684 19468 5693 19508
rect 7948 19424 7988 19972
rect 9196 19963 9236 19972
rect 10924 19928 10964 20056
rect 11011 19972 11020 20012
rect 11060 19972 11069 20012
rect 10051 19888 10060 19928
rect 10100 19888 10964 19928
rect 11020 19844 11060 19972
rect 10147 19804 10156 19844
rect 10196 19804 10924 19844
rect 10964 19804 11060 19844
rect 11116 19844 11156 20056
rect 11500 20012 11540 20056
rect 12010 19972 12019 20012
rect 12059 19972 12116 20012
rect 11500 19963 11540 19972
rect 11116 19804 11884 19844
rect 11924 19804 11933 19844
rect 12076 19508 12116 19972
rect 13638 19928 13728 19948
rect 12451 19888 12460 19928
rect 12500 19888 13728 19928
rect 13638 19868 13728 19888
rect 12163 19804 12172 19844
rect 12212 19804 12343 19844
rect 13638 19592 13728 19612
rect 12835 19552 12844 19592
rect 12884 19552 13728 19592
rect 13638 19532 13728 19552
rect 10579 19468 10588 19508
rect 10628 19468 11596 19508
rect 11636 19468 11645 19508
rect 12076 19468 12172 19508
rect 12212 19468 12221 19508
rect 4099 19384 4108 19424
rect 4148 19384 7988 19424
rect 7948 19340 7988 19384
rect 2179 19300 2188 19340
rect 2228 19300 2572 19340
rect 2612 19300 2621 19340
rect 3436 19331 4588 19340
rect 3476 19300 4588 19331
rect 4628 19300 4637 19340
rect 6115 19300 6124 19340
rect 6164 19300 6604 19340
rect 6644 19300 7084 19340
rect 7124 19300 7133 19340
rect 7852 19331 7892 19340
rect 3436 19282 3476 19291
rect 7948 19300 8236 19340
rect 8276 19300 8285 19340
rect 9004 19331 9524 19340
rect 9004 19300 9484 19331
rect 7852 19256 7892 19291
rect 67 19216 76 19256
rect 116 19216 1228 19256
rect 1268 19216 1277 19256
rect 4387 19216 4396 19256
rect 4436 19216 7892 19256
rect 9004 19172 9044 19300
rect 10723 19300 10732 19340
rect 10772 19300 11212 19340
rect 11252 19300 11261 19340
rect 11980 19331 12020 19340
rect 9484 19282 9524 19291
rect 11980 19256 12020 19291
rect 13638 19256 13728 19276
rect 9955 19216 9964 19256
rect 10004 19216 10013 19256
rect 10217 19216 10348 19256
rect 10388 19216 10397 19256
rect 10531 19216 10540 19256
rect 10580 19216 12020 19256
rect 12844 19216 13728 19256
rect 9964 19172 10004 19216
rect 12844 19172 12884 19216
rect 13638 19196 13728 19216
rect 4579 19132 4588 19172
rect 4628 19132 8524 19172
rect 8564 19132 9044 19172
rect 9091 19132 9100 19172
rect 9140 19132 10004 19172
rect 10195 19132 10204 19172
rect 10244 19132 12884 19172
rect 7913 19048 8044 19088
rect 8084 19048 8093 19088
rect 9667 19048 9676 19088
rect 9716 19048 10924 19088
rect 10964 19048 10973 19088
rect 4579 18964 4588 19004
rect 4628 18964 9292 19004
rect 9332 18964 9341 19004
rect 13638 18920 13728 18940
rect 3679 18880 3688 18920
rect 3728 18880 3770 18920
rect 3810 18880 3852 18920
rect 3892 18880 3934 18920
rect 3974 18880 4016 18920
rect 4056 18880 4065 18920
rect 12739 18880 12748 18920
rect 12788 18880 13728 18920
rect 13638 18860 13728 18880
rect 10060 18796 11692 18836
rect 11732 18796 11741 18836
rect 10060 18668 10100 18796
rect 3305 18628 3388 18668
rect 3428 18628 3436 18668
rect 3476 18628 3485 18668
rect 7180 18628 8332 18668
rect 8372 18628 8381 18668
rect 8851 18628 8860 18668
rect 8900 18628 10100 18668
rect 10252 18712 12308 18752
rect 0 18584 90 18604
rect 7180 18584 7220 18628
rect 0 18544 76 18584
rect 116 18544 125 18584
rect 3017 18544 3148 18584
rect 3188 18544 4052 18584
rect 7171 18544 7180 18584
rect 7220 18544 7229 18584
rect 8458 18544 8467 18584
rect 8507 18544 8620 18584
rect 8660 18544 8669 18584
rect 9763 18544 9772 18584
rect 9812 18544 10060 18584
rect 10100 18544 10109 18584
rect 0 18524 90 18544
rect 4012 18500 4052 18544
rect 5260 18500 5300 18509
rect 7756 18500 7796 18509
rect 3977 18460 4012 18500
rect 4052 18460 4108 18500
rect 4148 18460 4157 18500
rect 4387 18460 4396 18500
rect 4436 18460 5260 18500
rect 5260 18451 5300 18460
rect 5452 18460 6691 18500
rect 6731 18460 6740 18500
rect 6787 18460 6796 18500
rect 6836 18460 6892 18500
rect 6932 18460 6967 18500
rect 7145 18460 7276 18500
rect 7316 18460 7325 18500
rect 7625 18460 7756 18500
rect 7796 18460 7805 18500
rect 8035 18460 8044 18500
rect 8084 18460 8244 18500
rect 8284 18460 8293 18500
rect 9274 18460 9283 18500
rect 9323 18460 9332 18500
rect 9379 18460 9388 18500
rect 9428 18460 9484 18500
rect 9524 18460 9559 18500
rect 9859 18460 9868 18500
rect 9908 18460 9917 18500
rect 5452 18416 5492 18460
rect 7756 18451 7796 18460
rect 5443 18376 5452 18416
rect 5492 18376 5501 18416
rect 4919 18124 4928 18164
rect 4968 18124 5010 18164
rect 5050 18124 5092 18164
rect 5132 18124 5174 18164
rect 5214 18124 5256 18164
rect 5296 18124 5305 18164
rect 4675 18040 4684 18080
rect 4724 18040 9044 18080
rect 1459 17956 1468 17996
rect 1508 17956 2188 17996
rect 2228 17956 2237 17996
rect 6019 17956 6028 17996
rect 6068 17956 6124 17996
rect 6164 17956 6199 17996
rect 6787 17956 6796 17996
rect 6836 17956 7180 17996
rect 7220 17956 7229 17996
rect 8515 17956 8524 17996
rect 8564 17956 8660 17996
rect 2323 17872 2332 17912
rect 2372 17872 5836 17912
rect 5876 17872 5885 17912
rect 8620 17828 8660 17956
rect 9004 17912 9044 18040
rect 9292 17996 9332 18460
rect 9868 18332 9908 18460
rect 10252 18416 10292 18712
rect 11404 18628 12172 18668
rect 12212 18628 12221 18668
rect 11404 18584 11444 18628
rect 12268 18584 12308 18712
rect 12425 18628 12508 18668
rect 12548 18628 12556 18668
rect 12596 18628 12605 18668
rect 13638 18584 13728 18604
rect 11395 18544 11404 18584
rect 11444 18544 11453 18584
rect 11875 18544 11884 18584
rect 11924 18544 12055 18584
rect 12115 18544 12124 18584
rect 12164 18544 12212 18584
rect 12259 18544 12268 18584
rect 12308 18544 12317 18584
rect 12460 18544 13728 18584
rect 10348 18500 10388 18509
rect 12172 18500 12212 18544
rect 10388 18460 10435 18500
rect 10793 18460 10867 18500
rect 10907 18460 10924 18500
rect 10964 18460 10973 18500
rect 12067 18460 12076 18500
rect 12116 18460 12212 18500
rect 10348 18416 10388 18460
rect 9955 18376 9964 18416
rect 10004 18376 10292 18416
rect 10339 18376 10348 18416
rect 10388 18376 10397 18416
rect 9868 18292 10964 18332
rect 11011 18292 11020 18332
rect 11060 18292 11069 18332
rect 11635 18292 11644 18332
rect 11684 18292 11732 18332
rect 10924 18248 10964 18292
rect 11020 18248 11060 18292
rect 11692 18248 11732 18292
rect 10339 18208 10348 18248
rect 10388 18208 10636 18248
rect 10676 18208 10685 18248
rect 10915 18208 10924 18248
rect 10964 18208 10973 18248
rect 11020 18208 11500 18248
rect 11540 18208 11549 18248
rect 11692 18208 12076 18248
rect 12116 18208 12125 18248
rect 12460 18164 12500 18544
rect 13638 18524 13728 18544
rect 13638 18248 13728 18268
rect 13123 18208 13132 18248
rect 13172 18208 13728 18248
rect 13638 18188 13728 18208
rect 9091 17956 9100 17996
rect 9140 17956 9332 17996
rect 9484 18124 12500 18164
rect 9004 17872 9244 17912
rect 9284 17872 9293 17912
rect 2092 17788 2476 17828
rect 2516 17788 2525 17828
rect 3593 17788 3724 17828
rect 3764 17788 3773 17828
rect 5020 17788 5539 17828
rect 5579 17788 5740 17828
rect 5780 17788 5789 17828
rect 6124 17788 6133 17828
rect 6173 17788 6211 17828
rect 6499 17788 6508 17828
rect 6548 17788 6595 17828
rect 6641 17788 6650 17828
rect 6690 17788 6700 17828
rect 6740 17788 6830 17828
rect 6979 17788 6988 17828
rect 7028 17788 7660 17828
rect 7700 17788 7709 17828
rect 8620 17819 8948 17828
rect 8620 17788 8908 17819
rect 2092 17744 2132 17788
rect 3724 17770 3764 17779
rect 5020 17744 5060 17788
rect 6129 17744 6169 17788
rect 6339 17746 6364 17786
rect 6404 17746 6413 17786
rect 67 17704 76 17744
rect 116 17704 1228 17744
rect 1268 17704 1277 17744
rect 2083 17704 2092 17744
rect 2132 17704 2141 17744
rect 4099 17704 4108 17744
rect 4148 17704 4300 17744
rect 4340 17704 4349 17744
rect 4649 17704 4780 17744
rect 4820 17704 4829 17744
rect 5011 17704 5020 17744
rect 5060 17704 5069 17744
rect 6115 17704 6124 17744
rect 6164 17704 6173 17744
rect 6220 17704 6243 17744
rect 6283 17704 6292 17744
rect 4339 17620 4348 17660
rect 4388 17620 4972 17660
rect 5012 17620 5021 17660
rect 5251 17620 5260 17660
rect 5300 17620 5511 17660
rect 5551 17620 5560 17660
rect 0 17576 90 17596
rect 0 17536 76 17576
rect 116 17536 125 17576
rect 3907 17536 3916 17576
rect 3956 17536 4204 17576
rect 4244 17536 4253 17576
rect 5059 17536 5068 17576
rect 5108 17536 5731 17576
rect 5771 17536 5780 17576
rect 0 17516 90 17536
rect 3679 17368 3688 17408
rect 3728 17368 3770 17408
rect 3810 17368 3852 17408
rect 3892 17368 3934 17408
rect 3974 17368 4016 17408
rect 4056 17368 4065 17408
rect 6220 17324 6260 17704
rect 6339 17660 6379 17746
rect 6508 17744 6548 17788
rect 9283 17788 9292 17828
rect 9332 17788 9341 17828
rect 8908 17770 8948 17779
rect 6499 17704 6508 17744
rect 6548 17704 6557 17744
rect 6883 17704 6892 17744
rect 6932 17704 7124 17744
rect 7084 17660 7124 17704
rect 9292 17660 9332 17788
rect 9484 17744 9524 18124
rect 9833 17956 9916 17996
rect 9956 17956 9964 17996
rect 10004 17956 10013 17996
rect 10291 17956 10300 17996
rect 10340 17956 10540 17996
rect 10580 17956 10589 17996
rect 11587 17956 11596 17996
rect 11636 17956 12268 17996
rect 12308 17956 12317 17996
rect 13638 17912 13728 17932
rect 12259 17872 12268 17912
rect 12308 17872 13728 17912
rect 13638 17852 13728 17872
rect 10522 17788 10531 17828
rect 10571 17788 10580 17828
rect 10627 17788 10636 17828
rect 10676 17788 10868 17828
rect 10915 17788 10924 17828
rect 10964 17788 11020 17828
rect 11060 17788 11095 17828
rect 11561 17819 11692 17828
rect 11561 17788 11596 17819
rect 10540 17744 10580 17788
rect 10828 17744 10868 17788
rect 11636 17788 11692 17819
rect 11732 17788 11741 17828
rect 11945 17788 12076 17828
rect 12116 17788 12125 17828
rect 11596 17770 11636 17779
rect 12076 17770 12116 17779
rect 9475 17704 9484 17744
rect 9524 17704 9533 17744
rect 9667 17704 9676 17744
rect 9716 17704 9725 17744
rect 10051 17704 10060 17744
rect 10100 17704 10348 17744
rect 10388 17704 10397 17744
rect 10531 17704 10540 17744
rect 10580 17704 10627 17744
rect 10697 17704 10828 17744
rect 10868 17704 10877 17744
rect 10985 17704 11116 17744
rect 11156 17704 11165 17744
rect 9676 17660 9716 17704
rect 10828 17660 10868 17704
rect 6339 17620 7028 17660
rect 7075 17620 7084 17660
rect 7124 17620 7133 17660
rect 8611 17620 8620 17660
rect 8660 17620 9964 17660
rect 10004 17620 10013 17660
rect 10828 17620 13036 17660
rect 13076 17620 13085 17660
rect 6988 17576 7028 17620
rect 13638 17576 13728 17596
rect 6988 17536 7468 17576
rect 7508 17536 7517 17576
rect 12451 17536 12460 17576
rect 12500 17536 13728 17576
rect 13638 17516 13728 17536
rect 7267 17452 7276 17492
rect 7316 17452 11692 17492
rect 11732 17452 11741 17492
rect 3436 17284 6028 17324
rect 6068 17284 6077 17324
rect 6220 17284 6412 17324
rect 6452 17284 6461 17324
rect 1891 17200 1900 17240
rect 1940 17200 3244 17240
rect 3284 17200 3293 17240
rect 1459 17116 1468 17156
rect 1508 17116 3340 17156
rect 3380 17116 3389 17156
rect 3436 17072 3476 17284
rect 13638 17240 13728 17260
rect 3619 17200 3628 17240
rect 3668 17200 6220 17240
rect 6260 17200 6269 17240
rect 7337 17200 7468 17240
rect 7508 17200 7517 17240
rect 7747 17200 7756 17240
rect 7796 17200 7805 17240
rect 11827 17200 11836 17240
rect 11876 17200 12172 17240
rect 12212 17200 12221 17240
rect 12499 17200 12508 17240
rect 12548 17200 12844 17240
rect 12884 17200 12893 17240
rect 13315 17200 13324 17240
rect 13364 17200 13728 17240
rect 7756 17156 7796 17200
rect 13638 17180 13728 17200
rect 4579 17116 4588 17156
rect 4628 17116 7276 17156
rect 7316 17116 7325 17156
rect 7756 17116 7948 17156
rect 7988 17116 7997 17156
rect 5740 17072 5780 17116
rect 67 17032 76 17072
rect 116 17032 1228 17072
rect 1268 17032 1277 17072
rect 3235 17032 3244 17072
rect 3284 17032 3476 17072
rect 4396 17032 4876 17072
rect 4916 17032 4925 17072
rect 5059 17032 5068 17072
rect 5108 17032 5643 17072
rect 5740 17032 5803 17072
rect 4396 16988 4436 17032
rect 5603 16989 5643 17032
rect 3139 16948 3148 16988
rect 3188 16948 4300 16988
rect 4340 16948 4349 16988
rect 4396 16939 4436 16948
rect 4828 16948 4867 16988
rect 4907 16948 4916 16988
rect 5034 16948 5164 16988
rect 5205 16948 5214 16988
rect 5331 16948 5340 16988
rect 5380 16948 5396 16988
rect 5493 16948 5502 16988
rect 5542 16948 5551 16988
rect 5603 16979 5684 16989
rect 5763 16988 5803 17032
rect 5949 17032 6028 17072
rect 6068 17032 6077 17072
rect 5949 17030 5989 17032
rect 5871 16999 5989 17030
rect 5603 16948 5635 16979
rect 3331 16864 3340 16904
rect 3380 16864 3628 16904
rect 3668 16864 3677 16904
rect 4457 16780 4588 16820
rect 4628 16780 4637 16820
rect 0 16568 90 16588
rect 4828 16568 4868 16948
rect 4963 16780 4972 16820
rect 5012 16780 5068 16820
rect 5108 16780 5143 16820
rect 4919 16612 4928 16652
rect 4968 16612 5010 16652
rect 5050 16612 5092 16652
rect 5132 16612 5174 16652
rect 5214 16612 5256 16652
rect 5296 16612 5305 16652
rect 5356 16568 5396 16948
rect 5511 16904 5551 16948
rect 5626 16939 5635 16948
rect 5675 16939 5684 16979
rect 5730 16948 5739 16988
rect 5779 16948 5803 16988
rect 5848 16959 5857 16999
rect 5897 16990 5989 16999
rect 5897 16959 5911 16990
rect 6129 16988 6169 17116
rect 6211 17032 6220 17072
rect 6260 17032 6740 17072
rect 6700 16988 6740 17032
rect 6892 17032 7660 17072
rect 7700 17032 7709 17072
rect 6892 17030 6932 17032
rect 6844 17021 6932 17030
rect 6129 16948 6220 16988
rect 6260 16948 6269 16988
rect 6316 16948 6339 16988
rect 6379 16948 6388 16988
rect 6448 16948 6457 16988
rect 6497 16948 6506 16988
rect 6691 16948 6700 16988
rect 6740 16948 6749 16988
rect 6884 16990 6932 17021
rect 7756 16988 7796 17116
rect 7843 17032 7852 17072
rect 7892 17032 7988 17072
rect 10051 17032 10060 17072
rect 10100 17032 10444 17072
rect 10484 17032 10828 17072
rect 10868 17032 10877 17072
rect 11491 17032 11500 17072
rect 11540 17032 12076 17072
rect 12116 17032 12125 17072
rect 12259 17032 12268 17072
rect 12308 17032 12317 17072
rect 6844 16972 6884 16981
rect 7049 16948 7171 16988
rect 7220 16948 7229 16988
rect 7363 16948 7372 16988
rect 7412 16948 7479 16988
rect 7519 16948 7543 16988
rect 7640 16948 7649 16988
rect 7689 16948 7796 16988
rect 7948 16988 7988 17032
rect 9484 16988 9524 16997
rect 11020 16988 11060 16997
rect 8227 16948 8236 16988
rect 8276 16948 8620 16988
rect 8660 16948 8669 16988
rect 9449 16948 9484 16988
rect 9524 16948 9580 16988
rect 9620 16948 9629 16988
rect 9676 16948 9955 16988
rect 9995 16948 10004 16988
rect 10051 16948 10060 16988
rect 10100 16948 10109 16988
rect 10435 16948 10444 16988
rect 10484 16948 10540 16988
rect 10580 16948 10924 16988
rect 10964 16948 10973 16988
rect 11530 16948 11539 16988
rect 11579 16948 11884 16988
rect 11924 16948 11933 16988
rect 5626 16938 5684 16939
rect 6316 16904 6356 16948
rect 6466 16904 6506 16948
rect 7948 16939 7988 16948
rect 9484 16939 9524 16948
rect 9676 16904 9716 16948
rect 5452 16864 5551 16904
rect 6019 16864 6028 16904
rect 6068 16864 6316 16904
rect 6356 16864 6365 16904
rect 6412 16864 6508 16904
rect 6548 16864 6666 16904
rect 7468 16864 7852 16904
rect 7892 16864 7901 16904
rect 9667 16864 9676 16904
rect 9716 16864 9725 16904
rect 5452 16820 5492 16864
rect 5443 16780 5452 16820
rect 5492 16780 5501 16820
rect 5818 16780 5827 16820
rect 5867 16780 5876 16820
rect 6115 16780 6124 16820
rect 6164 16780 6220 16820
rect 6260 16780 6295 16820
rect 5836 16736 5876 16780
rect 5836 16696 6316 16736
rect 6356 16696 6365 16736
rect 6412 16652 6452 16864
rect 6857 16780 6988 16820
rect 7028 16780 7037 16820
rect 7241 16780 7267 16820
rect 7307 16780 7372 16820
rect 7412 16780 7421 16820
rect 7468 16736 7508 16864
rect 7738 16780 7747 16820
rect 7787 16780 7796 16820
rect 7756 16736 7796 16780
rect 6691 16696 6700 16736
rect 6740 16696 7508 16736
rect 7747 16696 7756 16736
rect 7796 16696 7843 16736
rect 10060 16652 10100 16948
rect 11020 16904 11060 16948
rect 12268 16904 12308 17032
rect 13638 16904 13728 16924
rect 10147 16864 10156 16904
rect 10196 16864 11060 16904
rect 11779 16864 11788 16904
rect 11828 16864 12308 16904
rect 12931 16864 12940 16904
rect 12980 16864 13728 16904
rect 13638 16844 13728 16864
rect 11561 16780 11692 16820
rect 11732 16780 11741 16820
rect 5731 16612 5740 16652
rect 5780 16612 6452 16652
rect 6499 16612 6508 16652
rect 6548 16612 10100 16652
rect 13638 16568 13728 16588
rect 0 16528 76 16568
rect 116 16528 125 16568
rect 4828 16528 4916 16568
rect 0 16508 90 16528
rect 3331 16444 3340 16484
rect 3380 16444 4780 16484
rect 4820 16444 4829 16484
rect 1459 16360 1468 16400
rect 1508 16360 4684 16400
rect 4724 16360 4733 16400
rect 4876 16316 4916 16528
rect 4972 16528 5396 16568
rect 12547 16528 12556 16568
rect 12596 16528 13728 16568
rect 4972 16484 5012 16528
rect 13638 16508 13728 16528
rect 4963 16444 4972 16484
rect 5012 16444 5021 16484
rect 5836 16444 6508 16484
rect 6548 16444 6557 16484
rect 7267 16444 7276 16484
rect 7316 16444 7852 16484
rect 7892 16444 7901 16484
rect 8803 16444 8812 16484
rect 8852 16444 9724 16484
rect 9764 16444 9773 16484
rect 10531 16444 10540 16484
rect 10580 16444 11404 16484
rect 11444 16444 11453 16484
rect 11827 16444 11836 16484
rect 11876 16444 11980 16484
rect 12020 16444 12029 16484
rect 12499 16444 12508 16484
rect 12548 16444 12748 16484
rect 12788 16444 12797 16484
rect 5836 16400 5876 16444
rect 4963 16360 4972 16400
rect 5012 16360 5876 16400
rect 5836 16316 5876 16360
rect 1769 16276 1900 16316
rect 1940 16276 1949 16316
rect 3148 16307 3476 16316
rect 3188 16276 3476 16307
rect 3523 16276 3532 16316
rect 3572 16276 3581 16316
rect 4195 16276 4204 16316
rect 4244 16307 4820 16316
rect 4244 16276 4780 16307
rect 3148 16258 3188 16267
rect 1097 16192 1228 16232
rect 1268 16192 1277 16232
rect 3436 16064 3476 16276
rect 3532 16148 3572 16276
rect 4876 16276 5539 16316
rect 5579 16276 5588 16316
rect 5635 16276 5644 16316
rect 5684 16276 5876 16316
rect 5932 16360 6796 16400
rect 6836 16360 6845 16400
rect 6988 16360 7180 16400
rect 7220 16360 7229 16400
rect 7555 16360 7564 16400
rect 7604 16360 8660 16400
rect 4780 16258 4820 16267
rect 5548 16232 5588 16276
rect 5548 16192 5740 16232
rect 5780 16192 5789 16232
rect 5932 16148 5972 16360
rect 6988 16316 7028 16360
rect 6019 16276 6028 16316
rect 6068 16276 6077 16316
rect 6604 16307 7028 16316
rect 3532 16108 5972 16148
rect 6028 16064 6068 16276
rect 6644 16276 7028 16307
rect 7084 16307 7276 16316
rect 6604 16258 6644 16267
rect 7124 16276 7276 16307
rect 7316 16276 7325 16316
rect 7546 16276 7555 16316
rect 7595 16276 7604 16316
rect 7651 16276 7660 16316
rect 7700 16276 7748 16316
rect 8035 16276 8044 16316
rect 8084 16276 8332 16316
rect 8372 16276 8381 16316
rect 8620 16307 8660 16360
rect 7084 16258 7124 16267
rect 6115 16192 6124 16232
rect 6164 16192 6173 16232
rect 6124 16148 6164 16192
rect 6124 16108 6796 16148
rect 6836 16108 6845 16148
rect 3436 16024 4204 16064
rect 4244 16024 4253 16064
rect 4963 16024 4972 16064
rect 5012 16024 5021 16064
rect 5155 16024 5164 16064
rect 5204 16024 7084 16064
rect 7124 16024 7133 16064
rect 4972 15980 5012 16024
rect 4972 15940 5644 15980
rect 5684 15940 5693 15980
rect 7564 15896 7604 16276
rect 7708 16148 7748 16276
rect 8969 16276 9100 16316
rect 9140 16276 9149 16316
rect 9833 16276 9964 16316
rect 10004 16276 10013 16316
rect 10627 16276 10636 16316
rect 10676 16276 11212 16316
rect 11252 16276 11261 16316
rect 8620 16258 8660 16267
rect 9100 16258 9140 16267
rect 9964 16232 10004 16276
rect 11212 16258 11252 16267
rect 13638 16232 13728 16252
rect 8009 16192 8140 16232
rect 8180 16192 8189 16232
rect 9322 16192 9331 16232
rect 9371 16192 9484 16232
rect 9524 16192 9533 16232
rect 9964 16192 10540 16232
rect 10580 16192 10589 16232
rect 11465 16192 11596 16232
rect 11636 16192 11645 16232
rect 12259 16192 12268 16232
rect 12308 16192 12317 16232
rect 12835 16192 12844 16232
rect 12884 16192 13728 16232
rect 12268 16148 12308 16192
rect 13638 16172 13728 16192
rect 7708 16108 8180 16148
rect 9859 16108 9868 16148
rect 9908 16108 12308 16148
rect 8140 16064 8180 16108
rect 8131 16024 8140 16064
rect 8180 16024 8189 16064
rect 9571 15940 9580 15980
rect 9620 15940 11404 15980
rect 11444 15940 11453 15980
rect 13638 15896 13728 15916
rect 3679 15856 3688 15896
rect 3728 15856 3770 15896
rect 3810 15856 3852 15896
rect 3892 15856 3934 15896
rect 3974 15856 4016 15896
rect 4056 15856 4065 15896
rect 7564 15856 9484 15896
rect 9524 15856 9533 15896
rect 10051 15856 10060 15896
rect 10100 15856 13728 15896
rect 13638 15836 13728 15856
rect 4780 15772 4972 15812
rect 5012 15772 5021 15812
rect 8515 15772 8524 15812
rect 8564 15772 9908 15812
rect 9955 15772 9964 15812
rect 10004 15772 10252 15812
rect 10292 15772 10301 15812
rect 2860 15604 3916 15644
rect 3956 15604 3965 15644
rect 0 15560 90 15580
rect 2860 15560 2900 15604
rect 0 15520 1228 15560
rect 1268 15520 1277 15560
rect 2083 15520 2092 15560
rect 2132 15520 2900 15560
rect 0 15500 90 15520
rect 3724 15476 3764 15485
rect 2345 15436 2476 15476
rect 2516 15436 2525 15476
rect 3916 15476 3956 15604
rect 4780 15476 4820 15772
rect 4876 15688 5164 15728
rect 5204 15688 5213 15728
rect 6154 15688 6163 15728
rect 6203 15688 7084 15728
rect 7124 15688 7133 15728
rect 7180 15688 7564 15728
rect 7604 15688 7613 15728
rect 8969 15688 9004 15728
rect 9044 15688 9100 15728
rect 9140 15688 9149 15728
rect 4876 15560 4916 15688
rect 4972 15604 6796 15644
rect 6836 15604 6845 15644
rect 4867 15520 4876 15560
rect 4916 15520 4925 15560
rect 4972 15476 5012 15604
rect 7180 15560 7220 15688
rect 7267 15604 7276 15644
rect 7316 15604 7604 15644
rect 8227 15604 8236 15644
rect 8276 15604 8620 15644
rect 8660 15604 9236 15644
rect 6883 15520 6892 15560
rect 6932 15520 6941 15560
rect 7180 15520 7508 15560
rect 5452 15476 5492 15485
rect 3916 15436 4387 15476
rect 4427 15436 4436 15476
rect 4483 15436 4492 15476
rect 4532 15436 4820 15476
rect 4963 15436 4972 15476
rect 5012 15436 5021 15476
rect 5251 15436 5260 15476
rect 5300 15436 5452 15476
rect 3724 15392 3764 15436
rect 5452 15427 5492 15436
rect 5644 15436 5940 15476
rect 5980 15436 5989 15476
rect 6394 15436 6403 15476
rect 6443 15436 6452 15476
rect 6499 15436 6508 15476
rect 6548 15436 6644 15476
rect 3724 15352 4204 15392
rect 4244 15352 4253 15392
rect 5644 15308 5684 15436
rect 6412 15392 6452 15436
rect 5731 15352 5740 15392
rect 5780 15352 6452 15392
rect 2323 15268 2332 15308
rect 2372 15268 2476 15308
rect 2516 15268 2525 15308
rect 4291 15268 4300 15308
rect 4340 15268 5684 15308
rect 4919 15100 4928 15140
rect 4968 15100 5010 15140
rect 5050 15100 5092 15140
rect 5132 15100 5174 15140
rect 5214 15100 5256 15140
rect 5296 15100 5305 15140
rect 5736 15056 5776 15352
rect 6604 15224 6644 15436
rect 6892 15392 6932 15520
rect 7468 15476 7508 15520
rect 6979 15436 6988 15476
rect 7028 15436 7084 15476
rect 7124 15436 7159 15476
rect 7564 15476 7604 15604
rect 8297 15520 8419 15560
rect 8468 15520 8477 15560
rect 9196 15476 9236 15604
rect 9868 15560 9908 15772
rect 12067 15688 12076 15728
rect 12116 15688 12268 15728
rect 12308 15688 12317 15728
rect 13638 15560 13728 15580
rect 9868 15520 10868 15560
rect 10828 15476 10868 15520
rect 12172 15520 13728 15560
rect 12076 15476 12116 15485
rect 7564 15436 7956 15476
rect 7996 15436 8005 15476
rect 8227 15436 8236 15476
rect 8276 15436 8279 15476
rect 8319 15436 8407 15476
rect 8515 15436 8524 15476
rect 8564 15436 8695 15476
rect 9236 15436 9580 15476
rect 9620 15436 9629 15476
rect 10409 15436 10444 15476
rect 10484 15436 10540 15476
rect 10580 15436 10589 15476
rect 10819 15436 10828 15476
rect 10868 15436 10924 15476
rect 10964 15436 11028 15476
rect 11203 15436 11212 15476
rect 11252 15436 12076 15476
rect 7468 15427 7508 15436
rect 9196 15427 9236 15436
rect 12076 15427 12116 15436
rect 6892 15352 7316 15392
rect 7276 15224 7316 15352
rect 2572 15016 2860 15056
rect 2900 15016 2909 15056
rect 3628 15016 5776 15056
rect 2572 14720 2612 15016
rect 3628 14972 3668 15016
rect 3610 14932 3619 14972
rect 3659 14932 3668 14972
rect 3715 14932 3724 14972
rect 3764 14932 5452 14972
rect 5492 14932 5501 14972
rect 3148 14848 3628 14888
rect 3668 14848 3677 14888
rect 3825 14848 3834 14888
rect 3874 14848 4012 14888
rect 4052 14848 4061 14888
rect 4204 14848 4300 14888
rect 4340 14848 4349 14888
rect 5225 14848 5260 14888
rect 5300 14848 5356 14888
rect 5396 14848 5405 14888
rect 3148 14804 3188 14848
rect 4204 14804 4244 14848
rect 5736 14804 5776 15016
rect 6466 15184 6644 15224
rect 7180 15184 7316 15224
rect 7564 15352 8611 15392
rect 8651 15352 8660 15392
rect 6466 14804 6506 15184
rect 7180 14888 7220 15184
rect 7564 15140 7604 15352
rect 12172 15308 12212 15520
rect 13638 15500 13728 15520
rect 8131 15268 8140 15308
rect 8180 15268 8189 15308
rect 9292 15268 12212 15308
rect 7267 15100 7276 15140
rect 7316 15100 7604 15140
rect 7939 15016 7948 15056
rect 7988 15016 8084 15056
rect 7267 14932 7276 14972
rect 7316 14932 7948 14972
rect 7988 14932 7997 14972
rect 8044 14888 8084 15016
rect 6700 14848 7700 14888
rect 6700 14804 6740 14848
rect 3130 14764 3139 14804
rect 3179 14764 3188 14804
rect 3514 14764 3523 14804
rect 3563 14764 3724 14804
rect 3764 14764 3773 14804
rect 4027 14764 4036 14804
rect 4076 14764 4099 14804
rect 4186 14764 4195 14804
rect 4235 14764 4244 14804
rect 4330 14764 4339 14804
rect 4379 14764 4388 14804
rect 4474 14764 4483 14804
rect 4523 14764 4532 14804
rect 4576 14764 4585 14804
rect 4628 14764 4759 14804
rect 4867 14764 4876 14804
rect 4916 14764 5047 14804
rect 5146 14764 5155 14804
rect 5204 14764 5548 14804
rect 5588 14764 5597 14804
rect 5731 14764 5740 14804
rect 5780 14764 5789 14804
rect 5923 14764 5932 14804
rect 5972 14764 6103 14804
rect 6202 14764 6211 14804
rect 6251 14764 6260 14804
rect 6307 14764 6316 14804
rect 6356 14764 6506 14804
rect 6691 14764 6700 14804
rect 6740 14764 6749 14804
rect 7276 14795 7564 14804
rect 4045 14720 4085 14764
rect 1411 14680 1420 14720
rect 1460 14680 2612 14720
rect 4003 14680 4012 14720
rect 4052 14680 4085 14720
rect 4348 14636 4388 14764
rect 4492 14720 4532 14764
rect 6220 14720 6260 14764
rect 7316 14764 7564 14795
rect 7604 14764 7613 14804
rect 7276 14746 7316 14755
rect 7660 14720 7700 14848
rect 7756 14848 8084 14888
rect 8140 14888 8180 15268
rect 8140 14848 8428 14888
rect 8468 14848 8477 14888
rect 7756 14795 7796 14848
rect 7843 14764 7852 14804
rect 7892 14764 8537 14804
rect 8577 14764 8586 14804
rect 8803 14764 8812 14804
rect 8852 14764 8861 14804
rect 7756 14746 7796 14755
rect 8812 14720 8852 14764
rect 9292 14720 9332 15268
rect 13638 15224 13728 15244
rect 13612 15164 13728 15224
rect 13612 15140 13652 15164
rect 12163 15100 12172 15140
rect 12212 15100 13652 15140
rect 12172 15016 13612 15056
rect 13652 15016 13661 15056
rect 12172 14972 12212 15016
rect 9475 14932 9484 14972
rect 9524 14932 9655 14972
rect 11347 14932 11356 14972
rect 11396 14932 12212 14972
rect 13638 14888 13728 14908
rect 10339 14848 10348 14888
rect 10388 14848 13728 14888
rect 13638 14828 13728 14848
rect 9571 14764 9580 14804
rect 9620 14795 9751 14804
rect 9620 14764 9676 14795
rect 9716 14764 9751 14795
rect 10793 14764 10924 14804
rect 10964 14764 10973 14804
rect 9676 14746 9716 14755
rect 10924 14720 10964 14764
rect 4492 14680 4684 14720
rect 4724 14680 4733 14720
rect 5731 14680 5740 14720
rect 5780 14680 5836 14720
rect 5876 14680 5911 14720
rect 6129 14680 6260 14720
rect 6787 14680 6796 14720
rect 6836 14680 7084 14720
rect 7124 14680 7133 14720
rect 7564 14680 7700 14720
rect 7939 14680 7948 14720
rect 7988 14680 8852 14720
rect 9283 14680 9292 14720
rect 9332 14680 9341 14720
rect 10924 14680 11116 14720
rect 11156 14680 11165 14720
rect 11561 14680 11692 14720
rect 11732 14680 11741 14720
rect 12067 14680 12076 14720
rect 12116 14680 12268 14720
rect 12308 14680 12317 14720
rect 12451 14680 12460 14720
rect 12500 14680 13132 14720
rect 13172 14680 13181 14720
rect 2467 14596 2476 14636
rect 2516 14596 3111 14636
rect 3151 14596 3236 14636
rect 3322 14596 3331 14636
rect 3371 14596 4388 14636
rect 5539 14596 5548 14636
rect 5588 14596 5836 14636
rect 5876 14596 5885 14636
rect 0 14552 90 14572
rect 0 14512 1180 14552
rect 1220 14512 1229 14552
rect 0 14492 90 14512
rect 3196 14468 3236 14596
rect 4579 14512 4588 14552
rect 4628 14512 5068 14552
rect 5108 14512 5117 14552
rect 6129 14468 6169 14680
rect 3196 14428 5836 14468
rect 5876 14428 6169 14468
rect 7564 14552 7604 14680
rect 7651 14596 7660 14636
rect 7700 14596 8140 14636
rect 8180 14596 8189 14636
rect 9091 14596 9100 14636
rect 9140 14596 9484 14636
rect 9524 14596 9533 14636
rect 9763 14596 9772 14636
rect 9812 14596 11452 14636
rect 11492 14596 11501 14636
rect 11596 14596 12220 14636
rect 12260 14596 12269 14636
rect 11596 14552 11636 14596
rect 13638 14552 13728 14572
rect 7564 14512 8332 14552
rect 8372 14512 8381 14552
rect 8524 14512 9052 14552
rect 9092 14512 9676 14552
rect 9716 14512 9725 14552
rect 10723 14512 10732 14552
rect 10772 14512 11636 14552
rect 11827 14512 11836 14552
rect 11876 14512 11885 14552
rect 13123 14512 13132 14552
rect 13172 14512 13728 14552
rect 7564 14384 7604 14512
rect 8524 14384 8564 14512
rect 11836 14468 11876 14512
rect 13638 14492 13728 14512
rect 9475 14428 9484 14468
rect 9524 14428 11876 14468
rect 3679 14344 3688 14384
rect 3728 14344 3770 14384
rect 3810 14344 3852 14384
rect 3892 14344 3934 14384
rect 3974 14344 4016 14384
rect 4056 14344 4065 14384
rect 7555 14344 7564 14384
rect 7604 14344 7613 14384
rect 8227 14344 8236 14384
rect 8276 14344 8564 14384
rect 8707 14344 8716 14384
rect 8756 14344 9100 14384
rect 9140 14344 9149 14384
rect 9667 14344 9676 14384
rect 9716 14344 10252 14384
rect 10292 14344 10301 14384
rect 11011 14344 11020 14384
rect 11060 14344 11069 14384
rect 11020 14300 11060 14344
rect 3139 14260 3148 14300
rect 3188 14260 7372 14300
rect 7412 14260 7421 14300
rect 9964 14260 11060 14300
rect 11107 14260 11116 14300
rect 11156 14260 12260 14300
rect 9964 14216 10004 14260
rect 12220 14216 12260 14260
rect 13638 14216 13728 14236
rect 4291 14176 4300 14216
rect 4340 14176 4876 14216
rect 4916 14176 4925 14216
rect 5059 14176 5068 14216
rect 5108 14176 7028 14216
rect 8585 14176 8668 14216
rect 8708 14176 8716 14216
rect 8756 14176 8765 14216
rect 9043 14176 9052 14216
rect 9092 14176 10004 14216
rect 10409 14176 10492 14216
rect 10532 14176 10540 14216
rect 10580 14176 10589 14216
rect 11875 14176 11884 14216
rect 11924 14176 12076 14216
rect 12116 14176 12125 14216
rect 12211 14176 12220 14216
rect 12260 14176 12269 14216
rect 12739 14176 12748 14216
rect 12788 14176 13728 14216
rect 4579 14092 4588 14132
rect 4628 14092 6356 14132
rect 1411 14008 1420 14048
rect 1460 14008 2380 14048
rect 2420 14008 2429 14048
rect 5164 14008 5356 14048
rect 5396 14008 5405 14048
rect 5548 14008 5836 14048
rect 5876 14008 5885 14048
rect 4396 13964 4436 13973
rect 5164 13964 5204 14008
rect 5548 13964 5588 14008
rect 6316 13964 6356 14092
rect 3043 13924 3052 13964
rect 3092 13924 3148 13964
rect 3188 13924 3223 13964
rect 4195 13924 4204 13964
rect 4244 13924 4396 13964
rect 5155 13924 5164 13964
rect 5204 13924 5213 13964
rect 5260 13955 5300 13964
rect 4396 13915 4436 13924
rect 5539 13924 5548 13964
rect 5588 13924 5597 13964
rect 5644 13924 6071 13964
rect 6111 13924 6120 13964
rect 6202 13924 6211 13964
rect 6251 13924 6260 13964
rect 6307 13924 6316 13964
rect 6356 13924 6892 13964
rect 6932 13924 6941 13964
rect 5260 13880 5300 13915
rect 5155 13840 5164 13880
rect 5204 13840 5300 13880
rect 67 13756 76 13796
rect 116 13756 1180 13796
rect 1220 13756 1229 13796
rect 4579 13756 4588 13796
rect 4628 13756 5068 13796
rect 5108 13756 5117 13796
rect 0 13544 90 13564
rect 0 13504 76 13544
rect 116 13504 125 13544
rect 4396 13504 4588 13544
rect 4628 13504 4637 13544
rect 0 13484 90 13504
rect 4396 13460 4436 13504
rect 4780 13460 4820 13756
rect 4919 13588 4928 13628
rect 4968 13588 5010 13628
rect 5050 13588 5092 13628
rect 5132 13588 5174 13628
rect 5214 13588 5256 13628
rect 5296 13588 5305 13628
rect 5644 13544 5684 13924
rect 6220 13880 6260 13924
rect 5260 13504 5684 13544
rect 5932 13840 6260 13880
rect 6988 13880 7028 14176
rect 13638 14156 13728 14176
rect 7555 14092 7564 14132
rect 7604 14092 7613 14132
rect 9292 14092 12020 14132
rect 7564 14048 7604 14092
rect 9292 14048 9332 14092
rect 7156 14008 7180 14048
rect 7220 14008 7229 14048
rect 7564 14008 7892 14048
rect 8323 14008 8332 14048
rect 8372 14008 8620 14048
rect 8660 14008 8669 14048
rect 8899 14008 8908 14048
rect 8948 14008 8957 14048
rect 9283 14008 9292 14048
rect 9332 14008 9341 14048
rect 9545 14008 9676 14048
rect 9716 14008 9725 14048
rect 9929 14008 10060 14048
rect 10100 14008 10109 14048
rect 10243 14008 10252 14048
rect 10292 14008 11596 14048
rect 11636 14008 11645 14048
rect 7156 13964 7196 14008
rect 7852 14006 7892 14008
rect 7852 13997 7935 14006
rect 7852 13966 7895 13997
rect 7133 13924 7147 13964
rect 7187 13924 7196 13964
rect 7258 13924 7267 13964
rect 7316 13924 7447 13964
rect 7747 13924 7756 13964
rect 7796 13924 7805 13964
rect 7895 13948 7935 13957
rect 8908 13964 8948 14008
rect 11884 13964 11924 13973
rect 8908 13924 10100 13964
rect 10627 13924 10636 13964
rect 10676 13924 10924 13964
rect 10964 13924 10973 13964
rect 11395 13924 11404 13964
rect 11444 13924 11884 13964
rect 7756 13880 7796 13924
rect 6988 13840 7796 13880
rect 8611 13840 8620 13880
rect 8660 13840 9436 13880
rect 9476 13840 9485 13880
rect 5260 13460 5300 13504
rect 5932 13460 5972 13840
rect 10060 13796 10100 13924
rect 11884 13915 11924 13924
rect 11980 13880 12020 14092
rect 12329 14008 12460 14048
rect 12500 14008 12509 14048
rect 13638 13880 13728 13900
rect 11980 13840 13728 13880
rect 13638 13820 13728 13840
rect 6281 13756 6316 13796
rect 6356 13756 6403 13796
rect 6443 13756 6461 13796
rect 8035 13756 8044 13796
rect 8084 13756 8524 13796
rect 8564 13756 8573 13796
rect 9811 13756 9820 13796
rect 9860 13756 9869 13796
rect 10060 13756 12404 13796
rect 9820 13712 9860 13756
rect 8419 13672 8428 13712
rect 8468 13672 9860 13712
rect 12364 13544 12404 13756
rect 13638 13544 13728 13564
rect 6403 13504 6412 13544
rect 6452 13504 6461 13544
rect 9091 13504 9100 13544
rect 9140 13504 12260 13544
rect 12364 13504 13728 13544
rect 6412 13460 6452 13504
rect 12220 13460 12260 13504
rect 13638 13484 13728 13504
rect 4387 13420 4396 13460
rect 4436 13420 4445 13460
rect 4553 13420 4675 13460
rect 4724 13420 4733 13460
rect 4780 13420 4876 13460
rect 4916 13420 4925 13460
rect 5251 13420 5260 13460
rect 5300 13420 5309 13460
rect 5539 13420 5548 13460
rect 5588 13420 5972 13460
rect 6394 13420 6403 13460
rect 6443 13420 6499 13460
rect 9641 13420 9724 13460
rect 9764 13420 9772 13460
rect 9812 13420 9821 13460
rect 10099 13420 10108 13460
rect 10148 13420 10156 13460
rect 10196 13420 10279 13460
rect 12211 13420 12220 13460
rect 12260 13420 12269 13460
rect 4291 13336 4300 13376
rect 4340 13336 4574 13376
rect 4614 13336 5551 13376
rect 5511 13292 5551 13336
rect 5740 13336 5836 13376
rect 5876 13336 5885 13376
rect 6019 13336 6028 13376
rect 6068 13336 6111 13376
rect 5740 13292 5780 13336
rect 6071 13292 6111 13336
rect 6316 13336 7948 13376
rect 7988 13336 7997 13376
rect 10243 13336 10252 13376
rect 10292 13336 11828 13376
rect 6316 13292 6356 13336
rect 2947 13252 2956 13292
rect 2996 13252 3127 13292
rect 4003 13252 4012 13292
rect 4052 13283 4244 13292
rect 4052 13252 4204 13283
rect 4649 13252 4684 13292
rect 4724 13252 4780 13292
rect 4820 13252 4829 13292
rect 4876 13283 4972 13292
rect 4204 13234 4244 13243
rect 4916 13252 4972 13283
rect 5012 13252 5059 13292
rect 5099 13252 5108 13292
rect 5251 13252 5260 13292
rect 5300 13252 5356 13292
rect 5396 13252 5431 13292
rect 5511 13252 5588 13292
rect 5740 13252 5763 13292
rect 5803 13252 5812 13292
rect 5872 13252 5881 13292
rect 5921 13271 5957 13292
rect 5921 13252 5972 13271
rect 6062 13252 6071 13292
rect 6111 13252 6120 13292
rect 6307 13252 6316 13292
rect 6356 13252 6365 13292
rect 6412 13252 6743 13292
rect 6783 13252 6792 13292
rect 6979 13252 6988 13292
rect 7028 13252 7159 13292
rect 8009 13283 8140 13292
rect 8009 13252 8044 13283
rect 4876 13234 4916 13243
rect 5548 13250 5588 13252
rect 5548 13210 5644 13250
rect 5684 13210 5693 13250
rect 5917 13231 5972 13252
rect 5932 13208 5972 13231
rect 6412 13208 6452 13252
rect 8084 13252 8140 13283
rect 8180 13252 8332 13292
rect 8372 13252 8381 13292
rect 8428 13252 9292 13292
rect 9332 13252 9341 13292
rect 10531 13252 10540 13292
rect 10580 13252 11596 13292
rect 11636 13252 11645 13292
rect 11788 13283 11828 13336
rect 8044 13234 8084 13243
rect 1289 13168 1324 13208
rect 1364 13168 1420 13208
rect 1460 13168 1469 13208
rect 5932 13168 5989 13208
rect 6202 13168 6211 13208
rect 6251 13168 6308 13208
rect 6403 13168 6412 13208
rect 6452 13168 6461 13208
rect 6761 13168 6883 13208
rect 6932 13168 6941 13208
rect 7075 13168 7084 13208
rect 7124 13168 7133 13208
rect 5949 13124 5989 13168
rect 6268 13124 6308 13168
rect 5836 13084 5989 13124
rect 6211 13084 6220 13124
rect 6260 13084 6308 13124
rect 25 13000 1180 13040
rect 1220 13000 1229 13040
rect 25 12704 65 13000
rect 5836 12956 5876 13084
rect 7084 13040 7124 13168
rect 8428 13124 8468 13252
rect 11788 13234 11828 13243
rect 12460 13252 13324 13292
rect 13364 13252 13373 13292
rect 12460 13208 12500 13252
rect 13638 13208 13728 13228
rect 8707 13168 8716 13208
rect 8756 13168 9484 13208
rect 9524 13168 9533 13208
rect 10217 13168 10348 13208
rect 10388 13168 10397 13208
rect 12451 13168 12460 13208
rect 12500 13168 12509 13208
rect 12556 13168 13728 13208
rect 12556 13124 12596 13168
rect 13638 13148 13728 13168
rect 7363 13084 7372 13124
rect 7412 13084 7948 13124
rect 7988 13084 8468 13124
rect 12067 13084 12076 13124
rect 12116 13084 12596 13124
rect 6883 13000 6892 13040
rect 6932 13000 7124 13040
rect 7843 13000 7852 13040
rect 7892 13000 8332 13040
rect 8372 13000 8381 13040
rect 11395 13000 11404 13040
rect 11444 13000 11980 13040
rect 12020 13000 12029 13040
rect 5836 12916 6124 12956
rect 6164 12916 7084 12956
rect 7124 12916 7133 12956
rect 13638 12872 13728 12892
rect 3679 12832 3688 12872
rect 3728 12832 3770 12872
rect 3810 12832 3852 12872
rect 3892 12832 3934 12872
rect 3974 12832 4016 12872
rect 4056 12832 4065 12872
rect 4684 12832 9772 12872
rect 9812 12832 9821 12872
rect 12451 12832 12460 12872
rect 12500 12832 13728 12872
rect 25 12664 116 12704
rect 76 12556 116 12664
rect 0 12496 116 12556
rect 3689 12496 3820 12536
rect 3860 12496 3869 12536
rect 0 12476 90 12496
rect 4684 12452 4724 12832
rect 13638 12812 13728 12832
rect 5356 12748 7756 12788
rect 7796 12748 7805 12788
rect 7948 12748 11692 12788
rect 11732 12748 11741 12788
rect 4841 12496 4972 12536
rect 5012 12496 5021 12536
rect 5356 12494 5396 12748
rect 6019 12664 6028 12704
rect 6068 12664 6700 12704
rect 6740 12664 6749 12704
rect 7948 12620 7988 12748
rect 8035 12664 8044 12704
rect 8084 12664 8860 12704
rect 8900 12664 8909 12704
rect 9449 12664 9532 12704
rect 9572 12664 9580 12704
rect 9620 12664 9629 12704
rect 11827 12664 11836 12704
rect 11876 12664 11980 12704
rect 12020 12664 12029 12704
rect 12163 12664 12172 12704
rect 12212 12664 12220 12704
rect 12260 12664 12343 12704
rect 6883 12580 6892 12620
rect 6932 12580 7180 12620
rect 7220 12580 7988 12620
rect 8803 12580 8812 12620
rect 8852 12580 9196 12620
rect 9236 12580 9245 12620
rect 9763 12580 9772 12620
rect 9812 12580 11500 12620
rect 11540 12580 11549 12620
rect 12076 12580 12556 12620
rect 12596 12580 12605 12620
rect 5299 12454 5308 12494
rect 5348 12454 5396 12494
rect 5452 12496 5836 12536
rect 5876 12496 5972 12536
rect 6979 12496 6988 12536
rect 7028 12496 7316 12536
rect 7459 12496 7468 12536
rect 7508 12496 7639 12536
rect 5452 12452 5492 12496
rect 5932 12452 5972 12496
rect 7276 12452 7316 12496
rect 7948 12452 7988 12580
rect 9091 12496 9100 12536
rect 9140 12496 9149 12536
rect 9283 12496 9292 12536
rect 9332 12496 9428 12536
rect 10243 12496 10252 12536
rect 10292 12496 10540 12536
rect 10580 12496 10589 12536
rect 8044 12452 8084 12461
rect 9100 12452 9140 12496
rect 3977 12412 4108 12452
rect 4148 12412 4157 12452
rect 4300 12412 4363 12452
rect 4403 12412 4412 12452
rect 4474 12412 4483 12452
rect 4523 12412 4724 12452
rect 4771 12412 4780 12452
rect 4820 12412 5068 12452
rect 5108 12412 5117 12452
rect 5164 12412 5187 12452
rect 5227 12412 5236 12452
rect 5443 12412 5452 12452
rect 5492 12412 5501 12452
rect 5585 12412 5594 12452
rect 5634 12412 5740 12452
rect 5780 12412 5789 12452
rect 5923 12412 5932 12452
rect 5972 12412 5981 12452
rect 6115 12412 6124 12452
rect 6164 12412 6508 12452
rect 6548 12412 6796 12452
rect 6836 12412 6845 12452
rect 6970 12412 6979 12452
rect 7019 12412 7028 12452
rect 7075 12412 7084 12452
rect 7124 12412 7220 12452
rect 7276 12412 7564 12452
rect 7604 12412 7892 12452
rect 7948 12412 8044 12452
rect 8323 12412 8332 12452
rect 8372 12412 8532 12452
rect 8572 12412 8581 12452
rect 9100 12412 9196 12452
rect 9236 12412 9245 12452
rect 4300 12368 4340 12412
rect 5164 12368 5204 12412
rect 6988 12368 7028 12412
rect 7180 12368 7220 12412
rect 4300 12328 4396 12368
rect 4436 12328 4445 12368
rect 5164 12328 6316 12368
rect 6356 12328 6365 12368
rect 6979 12328 6988 12368
rect 7028 12328 7075 12368
rect 7171 12328 7180 12368
rect 7220 12328 7229 12368
rect 3571 12244 3580 12284
rect 3620 12244 4204 12284
rect 4244 12244 4253 12284
rect 4819 12244 4828 12284
rect 4868 12244 4877 12284
rect 5731 12244 5740 12284
rect 5780 12244 7276 12284
rect 7316 12244 7325 12284
rect 3043 11908 3052 11948
rect 3092 11908 3196 11948
rect 3236 11908 3245 11948
rect 3859 11908 3868 11948
rect 3908 11908 4012 11948
rect 4052 11908 4061 11948
rect 4828 11780 4868 12244
rect 7852 12200 7892 12412
rect 8044 12403 8084 12412
rect 9388 12368 9428 12496
rect 10828 12452 10868 12580
rect 12076 12536 12116 12580
rect 13638 12536 13728 12556
rect 12067 12496 12076 12536
rect 12116 12496 12125 12536
rect 12451 12496 12460 12536
rect 12500 12496 12940 12536
rect 12980 12496 12989 12536
rect 13315 12496 13324 12536
rect 13364 12496 13728 12536
rect 13638 12476 13728 12496
rect 9754 12412 9763 12452
rect 9803 12412 9812 12452
rect 9859 12412 9868 12452
rect 9908 12412 10060 12452
rect 10100 12412 10109 12452
rect 10339 12412 10348 12452
rect 10388 12412 10397 12452
rect 11338 12412 11347 12452
rect 11387 12412 11404 12452
rect 11444 12412 11527 12452
rect 9100 12328 9428 12368
rect 9772 12368 9812 12412
rect 10348 12368 10388 12412
rect 10828 12403 10868 12412
rect 9772 12328 9868 12368
rect 9908 12328 9917 12368
rect 10147 12328 10156 12368
rect 10196 12328 10388 12368
rect 8585 12244 8716 12284
rect 8756 12244 8765 12284
rect 6403 12160 6412 12200
rect 6452 12160 8524 12200
rect 8564 12160 8573 12200
rect 4919 12076 4928 12116
rect 4968 12076 5010 12116
rect 5050 12076 5092 12116
rect 5132 12076 5174 12116
rect 5214 12076 5256 12116
rect 5296 12076 5305 12116
rect 6211 12076 6220 12116
rect 6260 12076 7180 12116
rect 7220 12076 7229 12116
rect 9100 11948 9140 12328
rect 11491 12244 11500 12284
rect 11540 12244 11596 12284
rect 11636 12244 11671 12284
rect 13638 12200 13728 12220
rect 13027 12160 13036 12200
rect 13076 12160 13728 12200
rect 13638 12140 13728 12160
rect 9187 12076 9196 12116
rect 9236 12076 13556 12116
rect 10147 11992 10156 12032
rect 10196 11992 11636 12032
rect 11596 11948 11636 11992
rect 7913 11908 7996 11948
rect 8036 11908 8044 11948
rect 8084 11908 8093 11948
rect 9091 11908 9100 11948
rect 9140 11908 9149 11948
rect 9484 11908 10252 11948
rect 10292 11908 10301 11948
rect 11347 11908 11356 11948
rect 11396 11908 11500 11948
rect 11540 11908 11549 11948
rect 11596 11908 11836 11948
rect 11876 11908 11885 11948
rect 12211 11908 12220 11948
rect 12260 11908 12364 11948
rect 12404 11908 12413 11948
rect 6115 11824 6124 11864
rect 6164 11824 8092 11864
rect 8132 11824 8141 11864
rect 4108 11740 4300 11780
rect 4340 11740 4349 11780
rect 4684 11740 4868 11780
rect 5347 11740 5356 11780
rect 5396 11740 5827 11780
rect 5867 11740 5876 11780
rect 5923 11740 5932 11780
rect 5972 11740 5981 11780
rect 6185 11740 6316 11780
rect 6356 11740 6365 11780
rect 6761 11740 6892 11780
rect 6932 11740 6941 11780
rect 7075 11740 7084 11780
rect 7124 11771 7412 11780
rect 7124 11740 7372 11771
rect 4108 11696 4148 11740
rect 4684 11696 4724 11740
rect 5932 11696 5972 11740
rect 6892 11722 6932 11731
rect 9161 11740 9283 11780
rect 9332 11740 9341 11780
rect 7372 11722 7412 11731
rect 9484 11696 9524 11908
rect 13516 11864 13556 12076
rect 13638 11864 13728 11884
rect 13516 11824 13728 11864
rect 13638 11804 13728 11824
rect 9641 11740 9772 11780
rect 9812 11740 9821 11780
rect 10243 11740 10252 11780
rect 10292 11740 10301 11780
rect 10723 11740 10732 11780
rect 10772 11740 10781 11780
rect 10841 11740 10850 11780
rect 10890 11740 11500 11780
rect 11540 11740 11549 11780
rect 11692 11740 12748 11780
rect 12788 11740 12797 11780
rect 9772 11722 9812 11731
rect 1411 11656 1420 11696
rect 1460 11656 2092 11696
rect 2132 11656 2141 11696
rect 2947 11656 2956 11696
rect 2996 11656 3127 11696
rect 4099 11656 4108 11696
rect 4148 11656 4157 11696
rect 4291 11656 4300 11696
rect 4340 11656 4349 11696
rect 4675 11656 4684 11696
rect 4724 11656 4733 11696
rect 5932 11656 6124 11696
rect 6164 11656 6173 11696
rect 6281 11656 6412 11696
rect 6452 11656 6461 11696
rect 7594 11656 7603 11696
rect 7643 11656 7756 11696
rect 7796 11656 7805 11696
rect 8323 11656 8332 11696
rect 8372 11656 8620 11696
rect 8660 11656 8716 11696
rect 8756 11656 8765 11696
rect 8947 11656 8956 11696
rect 8996 11656 9524 11696
rect 4300 11612 4340 11656
rect 10252 11612 10292 11740
rect 10339 11656 10348 11696
rect 10388 11656 10519 11696
rect 10732 11612 10772 11740
rect 11692 11696 11732 11740
rect 11107 11656 11116 11696
rect 11156 11656 11308 11696
rect 11348 11656 11357 11696
rect 11683 11656 11692 11696
rect 11732 11656 11741 11696
rect 12067 11656 12076 11696
rect 12116 11656 12268 11696
rect 12308 11656 12317 11696
rect 12451 11656 12460 11696
rect 12500 11656 12844 11696
rect 12884 11656 12893 11696
rect 13411 11656 13420 11696
rect 13460 11656 13469 11696
rect 13420 11612 13460 11656
rect 3331 11572 3340 11612
rect 3380 11572 4340 11612
rect 4972 11572 8812 11612
rect 8852 11572 8861 11612
rect 9091 11572 9100 11612
rect 9140 11572 10292 11612
rect 10348 11572 10772 11612
rect 11395 11572 11404 11612
rect 11444 11572 11452 11612
rect 11492 11572 11575 11612
rect 13324 11572 13460 11612
rect 0 11528 90 11548
rect 4972 11528 5012 11572
rect 10348 11528 10388 11572
rect 0 11488 1180 11528
rect 1220 11488 1229 11528
rect 4291 11488 4300 11528
rect 4340 11488 4540 11528
rect 4580 11488 4589 11528
rect 4915 11488 4924 11528
rect 4964 11488 5012 11528
rect 10051 11488 10060 11528
rect 10100 11488 10388 11528
rect 0 11468 90 11488
rect 13324 11444 13364 11572
rect 13638 11528 13728 11548
rect 13411 11488 13420 11528
rect 13460 11488 13728 11528
rect 13638 11468 13728 11488
rect 8035 11404 8044 11444
rect 8084 11404 13364 11444
rect 3679 11320 3688 11360
rect 3728 11320 3770 11360
rect 3810 11320 3852 11360
rect 3892 11320 3934 11360
rect 3974 11320 4016 11360
rect 4056 11320 4065 11360
rect 6595 11320 6604 11360
rect 6644 11320 9100 11360
rect 9140 11320 10156 11360
rect 10196 11320 10205 11360
rect 7276 11236 7852 11276
rect 7892 11236 7901 11276
rect 8620 11236 11788 11276
rect 11828 11236 11837 11276
rect 7276 11192 7316 11236
rect 8620 11192 8660 11236
rect 13638 11192 13728 11212
rect 3907 11152 3916 11192
rect 3956 11152 4108 11192
rect 4148 11152 4157 11192
rect 4675 11152 4684 11192
rect 4724 11152 5116 11192
rect 5156 11152 5165 11192
rect 6307 11152 6316 11192
rect 6356 11152 7276 11192
rect 7316 11152 7325 11192
rect 7603 11152 7612 11192
rect 7652 11152 8660 11192
rect 8716 11152 10540 11192
rect 10580 11152 10589 11192
rect 11491 11152 11500 11192
rect 11540 11152 11596 11192
rect 11636 11152 11671 11192
rect 12259 11152 12268 11192
rect 12308 11152 13728 11192
rect 1795 11068 1804 11108
rect 1844 11068 8332 11108
rect 8372 11068 8381 11108
rect 7372 11024 7412 11068
rect 8716 11024 8756 11152
rect 13638 11132 13728 11152
rect 9004 11068 10348 11108
rect 10388 11068 10397 11108
rect 10723 11068 10732 11108
rect 10772 11068 11836 11108
rect 11876 11068 11885 11108
rect 1289 10984 1420 11024
rect 1460 10984 1469 11024
rect 4675 10984 4684 11024
rect 4724 10984 5396 11024
rect 5530 10984 5539 11024
rect 5579 10984 6028 11024
rect 6068 10984 6077 11024
rect 6250 11015 6412 11024
rect 5356 10982 5396 10984
rect 3724 10940 3764 10949
rect 5356 10942 5404 10982
rect 5444 10942 5453 10982
rect 6250 10975 6259 11015
rect 6299 10984 6412 11015
rect 6452 10984 6461 11024
rect 7363 10984 7372 11024
rect 7412 10984 7421 11024
rect 7555 10984 7564 11024
rect 7604 10984 7756 11024
rect 7796 10984 7805 11024
rect 7852 10984 8716 11024
rect 8756 10984 8765 11024
rect 6299 10975 6308 10984
rect 6250 10974 6308 10975
rect 7852 10940 7892 10984
rect 9004 10940 9044 11068
rect 10243 10984 10252 11024
rect 10292 10984 11444 11024
rect 11945 10984 12076 11024
rect 12116 10984 12125 11024
rect 12451 10984 12460 11024
rect 12500 10984 13132 11024
rect 13172 10984 13181 11024
rect 9292 10940 9332 10949
rect 11404 10940 11444 10984
rect 2345 10900 2476 10940
rect 2516 10900 2525 10940
rect 3764 10900 4300 10940
rect 4340 10900 4349 10940
rect 5251 10900 5260 10940
rect 5300 10900 5309 10940
rect 5635 10900 5644 10940
rect 5684 10900 5836 10940
rect 5876 10900 5885 10940
rect 5993 10900 6124 10940
rect 6164 10900 6173 10940
rect 6352 10900 6361 10940
rect 6401 10900 6452 10940
rect 6499 10900 6508 10940
rect 6548 10900 7892 10940
rect 8218 10900 8227 10940
rect 8267 10900 8276 10940
rect 8323 10900 8332 10940
rect 8372 10900 8428 10940
rect 8468 10900 8503 10940
rect 8803 10900 8812 10940
rect 8852 10900 9044 10940
rect 9091 10900 9100 10940
rect 9140 10900 9292 10940
rect 9658 10900 9772 10940
rect 9820 10900 9838 10940
rect 10147 10900 10156 10940
rect 10196 10900 10205 10940
rect 3724 10891 3764 10900
rect 5260 10856 5300 10900
rect 6412 10856 6452 10900
rect 8236 10856 8276 10900
rect 5260 10816 5740 10856
rect 5780 10816 5789 10856
rect 6307 10816 6316 10856
rect 6356 10816 6452 10856
rect 7913 10816 7996 10856
rect 8036 10816 8044 10856
rect 8084 10816 8093 10856
rect 8236 10816 8908 10856
rect 8948 10816 8957 10856
rect 9004 10772 9044 10900
rect 9292 10891 9332 10900
rect 10156 10856 10196 10900
rect 11404 10891 11444 10900
rect 13638 10856 13728 10876
rect 1171 10732 1180 10772
rect 1220 10732 1229 10772
rect 5722 10732 5731 10772
rect 5771 10732 6892 10772
rect 6932 10732 6941 10772
rect 8908 10732 9044 10772
rect 9868 10816 10196 10856
rect 13123 10816 13132 10856
rect 13172 10816 13728 10856
rect 0 10520 90 10540
rect 1180 10520 1220 10732
rect 8908 10688 8948 10732
rect 6604 10648 8948 10688
rect 4919 10564 4928 10604
rect 4968 10564 5010 10604
rect 5050 10564 5092 10604
rect 5132 10564 5174 10604
rect 5214 10564 5256 10604
rect 5296 10564 5305 10604
rect 0 10480 1220 10520
rect 0 10460 90 10480
rect 4099 10396 4108 10436
rect 4148 10396 4684 10436
rect 4724 10396 5452 10436
rect 5492 10396 5501 10436
rect 5731 10396 5740 10436
rect 5780 10396 6028 10436
rect 6068 10396 6077 10436
rect 4300 10312 6220 10352
rect 6260 10312 6269 10352
rect 4300 10268 4340 10312
rect 2467 10228 2476 10268
rect 2516 10228 2668 10268
rect 2708 10228 2717 10268
rect 3916 10259 3956 10268
rect 4291 10228 4300 10268
rect 4340 10228 4349 10268
rect 4675 10228 4684 10268
rect 4724 10259 5588 10268
rect 4724 10228 5548 10259
rect 3916 10184 3956 10219
rect 4684 10184 4724 10228
rect 5731 10228 5740 10268
rect 5780 10228 5789 10268
rect 5897 10228 5932 10268
rect 5972 10228 6019 10268
rect 6059 10228 6077 10268
rect 6120 10228 6129 10268
rect 6169 10228 6178 10268
rect 6377 10228 6508 10268
rect 6548 10228 6557 10268
rect 5548 10210 5588 10219
rect 1411 10144 1420 10184
rect 1460 10144 1996 10184
rect 2036 10144 2045 10184
rect 3916 10144 4204 10184
rect 4244 10144 4724 10184
rect 5740 10184 5780 10228
rect 6124 10184 6164 10228
rect 6604 10184 6644 10648
rect 9868 10604 9908 10816
rect 13638 10796 13728 10816
rect 9955 10732 9964 10772
rect 10004 10732 10013 10772
rect 10627 10732 10636 10772
rect 10676 10732 12220 10772
rect 12260 10732 12269 10772
rect 7555 10564 7564 10604
rect 7604 10564 9908 10604
rect 9964 10436 10004 10732
rect 13638 10520 13728 10540
rect 10339 10480 10348 10520
rect 10388 10480 11828 10520
rect 11875 10480 11884 10520
rect 11924 10480 13728 10520
rect 11788 10436 11828 10480
rect 13638 10460 13728 10480
rect 7625 10396 7756 10436
rect 7796 10396 7805 10436
rect 9737 10396 9868 10436
rect 9908 10396 9917 10436
rect 9964 10396 11732 10436
rect 11788 10396 11836 10436
rect 11876 10396 11885 10436
rect 6979 10312 6988 10352
rect 7028 10312 8044 10352
rect 8084 10312 8093 10352
rect 9187 10312 9196 10352
rect 9236 10312 11452 10352
rect 11492 10312 11501 10352
rect 6691 10228 6700 10268
rect 6740 10259 7124 10268
rect 6740 10228 7084 10259
rect 7084 10210 7124 10219
rect 7564 10259 7604 10268
rect 8131 10228 8140 10268
rect 8180 10259 8311 10268
rect 8180 10228 8236 10259
rect 5740 10144 6028 10184
rect 6068 10144 6164 10184
rect 6595 10144 6604 10184
rect 6644 10144 6653 10184
rect 7564 10100 7604 10219
rect 8276 10228 8311 10259
rect 8419 10228 8428 10268
rect 8468 10228 9484 10268
rect 9524 10228 9533 10268
rect 10060 10259 10252 10268
rect 8236 10210 8276 10219
rect 10100 10228 10252 10259
rect 10292 10228 10301 10268
rect 11177 10228 11308 10268
rect 11348 10228 11357 10268
rect 10060 10210 10100 10219
rect 11692 10184 11732 10396
rect 12076 10228 13324 10268
rect 13364 10228 13373 10268
rect 12076 10184 12116 10228
rect 13638 10184 13728 10204
rect 11683 10144 11692 10184
rect 11732 10144 11741 10184
rect 12067 10144 12076 10184
rect 12116 10144 12125 10184
rect 12329 10144 12460 10184
rect 12500 10144 12509 10184
rect 12835 10144 12844 10184
rect 12884 10144 13728 10184
rect 13638 10124 13728 10144
rect 5731 10060 5740 10100
rect 5780 10060 7604 10100
rect 8419 10060 8428 10100
rect 8468 10060 12220 10100
rect 12260 10060 12269 10100
rect 67 9976 76 10016
rect 116 9976 1180 10016
rect 1220 9976 1229 10016
rect 13638 9848 13728 9868
rect 3679 9808 3688 9848
rect 3728 9808 3770 9848
rect 3810 9808 3852 9848
rect 3892 9808 3934 9848
rect 3974 9808 4016 9848
rect 4056 9808 4065 9848
rect 11299 9808 11308 9848
rect 11348 9808 13728 9848
rect 13638 9788 13728 9808
rect 4387 9724 4396 9764
rect 4436 9724 5260 9764
rect 5300 9724 5309 9764
rect 5539 9724 5548 9764
rect 5588 9724 11404 9764
rect 11444 9724 11453 9764
rect 2995 9640 3004 9680
rect 3044 9640 3436 9680
rect 3476 9640 3485 9680
rect 4963 9640 4972 9680
rect 5012 9640 5356 9680
rect 5396 9640 5405 9680
rect 8083 9640 8092 9680
rect 8132 9640 9388 9680
rect 9428 9640 9437 9680
rect 9641 9640 9772 9680
rect 9812 9640 9821 9680
rect 11779 9640 11788 9680
rect 11828 9640 11836 9680
rect 11876 9640 11959 9680
rect 4771 9556 4780 9596
rect 4820 9556 4829 9596
rect 5164 9556 6412 9596
rect 6452 9556 6461 9596
rect 6604 9556 6796 9596
rect 6836 9556 9100 9596
rect 9140 9556 9149 9596
rect 9283 9556 9292 9596
rect 9332 9556 9964 9596
rect 10004 9556 10013 9596
rect 10435 9556 10444 9596
rect 10484 9556 12220 9596
rect 12260 9556 12269 9596
rect 12460 9556 13036 9596
rect 13076 9556 13085 9596
rect 0 9512 90 9532
rect 0 9472 76 9512
rect 116 9472 125 9512
rect 2467 9472 2476 9512
rect 2516 9472 2764 9512
rect 2804 9472 2900 9512
rect 0 9452 90 9472
rect 2860 9428 2900 9472
rect 4780 9428 4820 9556
rect 5164 9428 5204 9556
rect 5539 9472 5548 9512
rect 5588 9472 6124 9512
rect 6164 9472 6173 9512
rect 6604 9428 6644 9556
rect 12460 9512 12500 9556
rect 13638 9512 13728 9532
rect 7721 9472 7756 9512
rect 7796 9472 7852 9512
rect 7892 9472 7901 9512
rect 10156 9472 10252 9512
rect 10292 9472 10301 9512
rect 11465 9472 11596 9512
rect 11636 9472 11645 9512
rect 12451 9472 12460 9512
rect 12500 9472 12509 9512
rect 12556 9472 13728 9512
rect 2860 9388 3532 9428
rect 3572 9388 3581 9428
rect 4579 9388 4588 9428
rect 4628 9388 4780 9428
rect 4867 9388 4876 9428
rect 4916 9388 5164 9428
rect 5204 9388 5213 9428
rect 5347 9388 5356 9428
rect 5396 9388 5527 9428
rect 5626 9388 5635 9428
rect 5675 9388 5684 9428
rect 5731 9388 5740 9428
rect 5780 9388 6028 9428
rect 6068 9388 6077 9428
rect 6211 9388 6220 9428
rect 6260 9388 6644 9428
rect 6700 9428 6740 9437
rect 9580 9428 9620 9437
rect 10156 9428 10196 9472
rect 12556 9428 12596 9472
rect 13638 9452 13728 9472
rect 6740 9388 6988 9428
rect 7028 9388 7037 9428
rect 7210 9388 7219 9428
rect 7259 9388 7660 9428
rect 7700 9388 7709 9428
rect 8201 9388 8332 9428
rect 8372 9388 8381 9428
rect 9449 9388 9580 9428
rect 9620 9388 9629 9428
rect 4780 9379 4820 9388
rect 4876 9304 5492 9344
rect 4876 9176 4916 9304
rect 5338 9220 5347 9260
rect 5387 9220 5396 9260
rect 4492 9136 4916 9176
rect 4492 8924 4532 9136
rect 4919 9052 4928 9092
rect 4968 9052 5010 9092
rect 5050 9052 5092 9092
rect 5132 9052 5174 9092
rect 5214 9052 5256 9092
rect 5296 9052 5305 9092
rect 4483 8884 4492 8924
rect 4532 8884 4541 8924
rect 5356 8840 5396 9220
rect 5452 9176 5492 9304
rect 5644 9260 5684 9388
rect 6700 9379 6740 9388
rect 8332 9260 8372 9388
rect 9580 9379 9620 9388
rect 10156 9379 10196 9388
rect 10252 9388 11404 9428
rect 11444 9388 11453 9428
rect 12547 9388 12556 9428
rect 12596 9388 12605 9428
rect 10252 9260 10292 9388
rect 5539 9220 5548 9260
rect 5588 9220 5684 9260
rect 7363 9220 7372 9260
rect 7412 9220 7421 9260
rect 8332 9220 10292 9260
rect 7372 9176 7412 9220
rect 13638 9176 13728 9196
rect 5452 9136 5740 9176
rect 5780 9136 5789 9176
rect 7372 9136 8332 9176
rect 8372 9136 8381 9176
rect 8908 9136 10484 9176
rect 11683 9136 11692 9176
rect 11732 9136 13728 9176
rect 8908 9008 8948 9136
rect 5731 8968 5740 9008
rect 5780 8968 7124 9008
rect 7171 8968 7180 9008
rect 7220 8968 8948 9008
rect 7084 8924 7124 8968
rect 5539 8884 5548 8924
rect 5588 8884 6020 8924
rect 6115 8884 6124 8924
rect 6164 8884 6307 8924
rect 6347 8884 6356 8924
rect 7066 8884 7075 8924
rect 7115 8884 7124 8924
rect 8777 8884 8908 8924
rect 8948 8884 8957 8924
rect 9091 8884 9100 8924
rect 9140 8884 10300 8924
rect 10340 8884 10349 8924
rect 5164 8800 5260 8840
rect 5300 8800 5309 8840
rect 5356 8800 5684 8840
rect 2467 8716 2476 8756
rect 2516 8716 3052 8756
rect 3092 8716 3101 8756
rect 4300 8747 4492 8756
rect 4340 8716 4492 8747
rect 4532 8716 4541 8756
rect 4649 8716 4780 8756
rect 4820 8716 4829 8756
rect 4915 8716 4924 8756
rect 4964 8716 5068 8756
rect 5108 8716 5117 8756
rect 5164 8747 5204 8800
rect 5644 8756 5684 8800
rect 5980 8756 6020 8884
rect 10444 8840 10484 9136
rect 13638 9116 13728 9136
rect 10531 8884 10540 8924
rect 10580 8884 11068 8924
rect 11108 8884 11117 8924
rect 11395 8884 11404 8924
rect 11444 8884 11452 8924
rect 11492 8884 11575 8924
rect 11827 8884 11836 8924
rect 11876 8884 13516 8924
rect 13556 8884 13565 8924
rect 13638 8840 13728 8860
rect 6370 8800 6412 8840
rect 6452 8800 6461 8840
rect 6787 8800 6796 8840
rect 6836 8800 6845 8840
rect 8131 8800 8140 8840
rect 8180 8800 9340 8840
rect 9380 8800 9389 8840
rect 10444 8800 10684 8840
rect 10724 8800 10733 8840
rect 10924 8800 13728 8840
rect 4300 8698 4340 8707
rect 5386 8747 5452 8756
rect 5164 8698 5204 8707
rect 5254 8696 5263 8736
rect 5303 8696 5315 8736
rect 5386 8707 5395 8747
rect 5435 8716 5452 8747
rect 5492 8716 5575 8756
rect 5644 8716 5740 8756
rect 5780 8716 5789 8756
rect 5971 8716 5980 8756
rect 6020 8716 6029 8756
rect 6079 8747 6220 8756
rect 5435 8707 5444 8716
rect 5386 8706 5444 8707
rect 1411 8632 1420 8672
rect 1460 8632 1900 8672
rect 1940 8632 1949 8672
rect 0 8504 90 8524
rect 5275 8504 5315 8696
rect 5866 8674 5875 8714
rect 5915 8674 5929 8714
rect 6119 8716 6220 8747
rect 6260 8716 6269 8756
rect 6370 8742 6410 8800
rect 6796 8756 6836 8800
rect 6079 8698 6119 8707
rect 6370 8702 6454 8742
rect 6494 8702 6503 8742
rect 6604 8716 6652 8756
rect 6692 8716 6701 8756
rect 6749 8716 6763 8756
rect 6803 8716 6836 8756
rect 6979 8716 6988 8756
rect 7028 8716 7037 8756
rect 7459 8716 7468 8756
rect 7508 8716 7564 8756
rect 7604 8716 7639 8756
rect 8716 8747 8908 8756
rect 5889 8588 5929 8674
rect 6604 8672 6644 8716
rect 6595 8632 6604 8672
rect 6644 8632 6653 8672
rect 6761 8632 6883 8672
rect 6932 8632 6941 8672
rect 5889 8548 6028 8588
rect 6068 8548 6077 8588
rect 6988 8504 7028 8716
rect 8756 8716 8908 8747
rect 8948 8716 9580 8756
rect 9620 8716 9629 8756
rect 8716 8698 8756 8707
rect 10924 8672 10964 8800
rect 13638 8780 13728 8800
rect 9091 8632 9100 8672
rect 9140 8632 9292 8672
rect 9332 8632 9341 8672
rect 10531 8632 10540 8672
rect 10580 8632 10589 8672
rect 10915 8632 10924 8672
rect 10964 8632 10973 8672
rect 11177 8632 11308 8672
rect 11348 8632 11357 8672
rect 11683 8632 11692 8672
rect 11732 8632 11884 8672
rect 11924 8632 11933 8672
rect 12067 8632 12076 8672
rect 12116 8632 12268 8672
rect 12308 8632 12317 8672
rect 12451 8632 12460 8672
rect 12500 8632 13420 8672
rect 13460 8632 13469 8672
rect 10540 8588 10580 8632
rect 10540 8548 12500 8588
rect 12460 8504 12500 8548
rect 13638 8504 13728 8524
rect 0 8464 1180 8504
rect 1220 8464 1229 8504
rect 5275 8464 5644 8504
rect 5684 8464 5693 8504
rect 6019 8464 6028 8504
rect 6068 8464 7028 8504
rect 12163 8464 12172 8504
rect 12212 8464 12220 8504
rect 12260 8464 12343 8504
rect 12460 8464 13728 8504
rect 0 8444 90 8464
rect 13638 8444 13728 8464
rect 3679 8296 3688 8336
rect 3728 8296 3770 8336
rect 3810 8296 3852 8336
rect 3892 8296 3934 8336
rect 3974 8296 4016 8336
rect 4056 8296 4065 8336
rect 6979 8212 6988 8252
rect 7028 8212 11252 8252
rect 11212 8168 11252 8212
rect 13638 8168 13728 8188
rect 4771 8128 4780 8168
rect 4820 8128 5548 8168
rect 5588 8128 5597 8168
rect 5705 8128 5836 8168
rect 5876 8128 5885 8168
rect 8515 8128 8524 8168
rect 8564 8128 8572 8168
rect 8612 8128 8695 8168
rect 9379 8128 9388 8168
rect 9428 8128 11068 8168
rect 11108 8128 11117 8168
rect 11212 8128 11452 8168
rect 11492 8128 11501 8168
rect 12067 8128 12076 8168
rect 12116 8128 13728 8168
rect 13638 8108 13728 8128
rect 5347 8044 5356 8084
rect 5396 8044 5930 8084
rect 7939 8044 7948 8084
rect 7988 8044 8468 8084
rect 9667 8044 9676 8084
rect 9716 8044 9908 8084
rect 10099 8044 10108 8084
rect 10148 8044 11980 8084
rect 12020 8044 12029 8084
rect 12076 8044 12844 8084
rect 12884 8044 12893 8084
rect 1289 7960 1420 8000
rect 1460 7960 1469 8000
rect 5890 7958 5930 8044
rect 8201 7960 8332 8000
rect 8372 7960 8381 8000
rect 5356 7916 5396 7925
rect 5871 7918 5880 7958
rect 5920 7918 5930 7958
rect 7948 7916 7988 7925
rect 4099 7876 4108 7916
rect 4148 7876 4157 7916
rect 4675 7876 4684 7916
rect 4724 7876 5356 7916
rect 5609 7876 5740 7916
rect 5780 7876 5789 7916
rect 5980 7876 5989 7916
rect 6029 7876 6124 7916
rect 6164 7876 6173 7916
rect 6569 7876 6700 7916
rect 6740 7876 6749 7916
rect 7988 7876 8140 7916
rect 8180 7876 8189 7916
rect 4108 7832 4148 7876
rect 5356 7867 5396 7876
rect 7948 7867 7988 7876
rect 8428 7832 8468 8044
rect 9868 8000 9908 8044
rect 12076 8000 12116 8044
rect 9859 7960 9868 8000
rect 9908 7960 9917 8000
rect 11299 7960 11308 8000
rect 11348 7960 11357 8000
rect 11561 7960 11692 8000
rect 11732 7960 11741 8000
rect 12067 7960 12076 8000
rect 12116 7960 12125 8000
rect 12211 7960 12220 8000
rect 12260 7960 12268 8000
rect 12308 7960 12391 8000
rect 12451 7960 12460 8000
rect 12500 7960 13132 8000
rect 13172 7960 13181 8000
rect 8873 7876 9004 7916
rect 9044 7876 9053 7916
rect 9274 7876 9283 7916
rect 9323 7876 10060 7916
rect 10100 7876 10109 7916
rect 11308 7832 11348 7960
rect 13638 7832 13728 7852
rect 4108 7792 4724 7832
rect 8323 7792 8332 7832
rect 8372 7792 8468 7832
rect 9091 7792 9100 7832
rect 9140 7792 9388 7832
rect 9428 7792 9484 7832
rect 9524 7792 9533 7832
rect 11308 7792 13728 7832
rect 1171 7708 1180 7748
rect 1220 7708 1229 7748
rect 0 7496 90 7516
rect 1180 7496 1220 7708
rect 0 7456 1220 7496
rect 0 7436 90 7456
rect 4684 7160 4724 7792
rect 13638 7772 13728 7792
rect 7939 7708 7948 7748
rect 7988 7708 8140 7748
rect 8180 7708 8189 7748
rect 8236 7708 11836 7748
rect 11876 7708 11885 7748
rect 8236 7664 8276 7708
rect 8131 7624 8140 7664
rect 8180 7624 8276 7664
rect 4919 7540 4928 7580
rect 4968 7540 5010 7580
rect 5050 7540 5092 7580
rect 5132 7540 5174 7580
rect 5214 7540 5256 7580
rect 5296 7540 5305 7580
rect 13638 7496 13728 7516
rect 12451 7456 12460 7496
rect 12500 7456 13728 7496
rect 13638 7436 13728 7456
rect 5251 7372 5260 7412
rect 5300 7372 8084 7412
rect 4771 7288 4780 7328
rect 4820 7288 5300 7328
rect 5434 7288 5443 7328
rect 5483 7288 6028 7328
rect 6068 7288 6077 7328
rect 5260 7244 5300 7288
rect 8044 7244 8084 7372
rect 4867 7204 4876 7244
rect 4916 7204 5111 7244
rect 5151 7204 5160 7244
rect 5242 7204 5251 7244
rect 5291 7204 5300 7244
rect 5347 7204 5356 7244
rect 5396 7204 5527 7244
rect 6665 7204 6796 7244
rect 6836 7204 6845 7244
rect 8044 7235 8716 7244
rect 1289 7120 1420 7160
rect 1460 7120 1469 7160
rect 4675 7120 4684 7160
rect 4724 7120 4733 7160
rect 4841 7120 4924 7160
rect 4964 7120 4972 7160
rect 5012 7120 5021 7160
rect 4684 7076 4724 7120
rect 6796 7076 6836 7204
rect 8084 7204 8716 7235
rect 8756 7204 8765 7244
rect 11212 7204 12212 7244
rect 8044 7186 8084 7195
rect 11212 7160 11252 7204
rect 12172 7160 12212 7204
rect 13638 7160 13728 7180
rect 10819 7120 10828 7160
rect 10868 7120 11252 7160
rect 11299 7120 11308 7160
rect 11348 7120 11479 7160
rect 11683 7120 11692 7160
rect 11732 7120 11741 7160
rect 11945 7120 12076 7160
rect 12116 7120 12125 7160
rect 12172 7120 12220 7160
rect 12260 7120 12269 7160
rect 12451 7120 12460 7160
rect 12500 7120 12556 7160
rect 12596 7120 12631 7160
rect 12748 7120 13728 7160
rect 11692 7076 11732 7120
rect 12748 7076 12788 7120
rect 13638 7100 13728 7120
rect 4684 7036 6836 7076
rect 8227 7036 8236 7076
rect 8276 7036 9004 7076
rect 9044 7036 9053 7076
rect 9100 7036 11452 7076
rect 11492 7036 11501 7076
rect 11692 7036 12788 7076
rect 9100 6992 9140 7036
rect 547 6952 556 6992
rect 596 6952 1180 6992
rect 1220 6952 1229 6992
rect 6115 6952 6124 6992
rect 6164 6952 9140 6992
rect 9196 6952 11068 6992
rect 11108 6952 11117 6992
rect 11212 6952 11836 6992
rect 11876 6952 11885 6992
rect 9196 6908 9236 6952
rect 7267 6868 7276 6908
rect 7316 6868 9236 6908
rect 11212 6824 11252 6952
rect 13638 6824 13728 6844
rect 3679 6784 3688 6824
rect 3728 6784 3770 6824
rect 3810 6784 3852 6824
rect 3892 6784 3934 6824
rect 3974 6784 4016 6824
rect 4056 6784 4065 6824
rect 4387 6784 4396 6824
rect 4436 6784 11252 6824
rect 12076 6784 13728 6824
rect 5164 6700 6220 6740
rect 6260 6700 6269 6740
rect 5164 6656 5204 6700
rect 5155 6616 5164 6656
rect 5204 6616 5213 6656
rect 5635 6616 5644 6656
rect 5684 6616 11836 6656
rect 11876 6616 11885 6656
rect 4867 6532 4876 6572
rect 4916 6532 5684 6572
rect 7363 6532 7372 6572
rect 7412 6532 9484 6572
rect 9524 6532 9533 6572
rect 0 6488 90 6508
rect 5644 6488 5684 6532
rect 12076 6488 12116 6784
rect 13638 6764 13728 6784
rect 13638 6488 13728 6508
rect 0 6448 556 6488
rect 596 6448 605 6488
rect 5635 6448 5644 6488
rect 5684 6448 5693 6488
rect 11561 6448 11692 6488
rect 11732 6448 11741 6488
rect 12067 6448 12076 6488
rect 12116 6448 12125 6488
rect 12329 6448 12460 6488
rect 12500 6448 12509 6488
rect 12556 6448 13728 6488
rect 0 6428 90 6448
rect 4972 6404 5012 6413
rect 8812 6404 8852 6413
rect 12556 6404 12596 6448
rect 13638 6428 13728 6448
rect 1507 6364 1516 6404
rect 1556 6364 3724 6404
rect 3764 6364 3773 6404
rect 4675 6364 4684 6404
rect 4724 6364 4972 6404
rect 6569 6364 6700 6404
rect 6740 6364 6749 6404
rect 6970 6364 6979 6404
rect 7019 6364 7316 6404
rect 7433 6364 7564 6404
rect 7604 6364 7613 6404
rect 8681 6364 8812 6404
rect 8852 6364 9292 6404
rect 9332 6364 9341 6404
rect 11299 6364 11308 6404
rect 11348 6364 12596 6404
rect 4972 6355 5012 6364
rect 7276 6320 7316 6364
rect 8812 6355 8852 6364
rect 5731 6280 5740 6320
rect 5780 6280 7084 6320
rect 7124 6280 7133 6320
rect 7276 6280 7756 6320
rect 7796 6280 7805 6320
rect 8908 6280 11452 6320
rect 11492 6280 11501 6320
rect 5740 6236 5780 6280
rect 8908 6236 8948 6280
rect 4771 6196 4780 6236
rect 4820 6196 5780 6236
rect 7459 6196 7468 6236
rect 7508 6196 8948 6236
rect 8995 6196 9004 6236
rect 9044 6196 9580 6236
rect 9620 6196 9629 6236
rect 12211 6196 12220 6236
rect 12260 6196 12269 6236
rect 12220 6152 12260 6196
rect 13638 6152 13728 6172
rect 5635 6112 5644 6152
rect 5684 6112 12260 6152
rect 12451 6112 12460 6152
rect 12500 6112 13728 6152
rect 13638 6092 13728 6112
rect 4919 6028 4928 6068
rect 4968 6028 5010 6068
rect 5050 6028 5092 6068
rect 5132 6028 5174 6068
rect 5214 6028 5256 6068
rect 5296 6028 5305 6068
rect 13638 5816 13728 5836
rect 3715 5776 3724 5816
rect 3764 5776 4108 5816
rect 4148 5776 4436 5816
rect 4396 5732 4436 5776
rect 7756 5776 8812 5816
rect 8852 5776 8861 5816
rect 11683 5776 11692 5816
rect 11732 5776 13728 5816
rect 7756 5732 7796 5776
rect 13638 5756 13728 5776
rect 3017 5692 3052 5732
rect 3092 5692 3148 5732
rect 3188 5692 3197 5732
rect 4300 5723 4340 5732
rect 4396 5692 4684 5732
rect 4724 5692 4733 5732
rect 5932 5723 5972 5732
rect 4300 5648 4340 5683
rect 6211 5692 6220 5732
rect 6260 5692 6316 5732
rect 6356 5692 6391 5732
rect 7564 5723 7796 5732
rect 5932 5648 5972 5683
rect 7604 5692 7796 5723
rect 7913 5692 7948 5732
rect 7988 5692 8035 5732
rect 8075 5692 8093 5732
rect 8136 5692 8145 5732
rect 8185 5692 8194 5732
rect 8419 5692 8428 5732
rect 8468 5692 8524 5732
rect 8564 5692 8599 5732
rect 8969 5692 9100 5732
rect 9140 5692 9149 5732
rect 9449 5692 9580 5732
rect 9620 5692 9629 5732
rect 11779 5692 11788 5732
rect 11828 5692 12260 5732
rect 7564 5648 7604 5683
rect 8140 5648 8180 5692
rect 9100 5674 9140 5683
rect 9580 5674 9620 5683
rect 12220 5648 12260 5692
rect 1411 5608 1420 5648
rect 1460 5608 4244 5648
rect 4300 5608 4492 5648
rect 4532 5608 4541 5648
rect 4675 5608 4684 5648
rect 4724 5608 5452 5648
rect 5492 5608 7604 5648
rect 7747 5608 7756 5648
rect 7796 5608 8180 5648
rect 8611 5608 8620 5648
rect 8660 5608 8669 5648
rect 9802 5608 9811 5648
rect 9851 5608 9964 5648
rect 10004 5608 10013 5648
rect 10195 5608 10204 5648
rect 10244 5608 10348 5648
rect 10388 5608 10397 5648
rect 12067 5608 12076 5648
rect 12116 5608 12125 5648
rect 12211 5608 12220 5648
rect 12260 5608 12269 5648
rect 12329 5608 12460 5648
rect 12500 5608 12509 5648
rect 0 5480 90 5500
rect 4204 5480 4244 5608
rect 8620 5564 8660 5608
rect 12076 5564 12116 5608
rect 4483 5524 4492 5564
rect 4532 5524 5836 5564
rect 5876 5524 5885 5564
rect 6115 5524 6124 5564
rect 6164 5524 7084 5564
rect 7124 5524 7133 5564
rect 7651 5524 7660 5564
rect 7700 5524 7756 5564
rect 7796 5524 7831 5564
rect 8620 5524 9676 5564
rect 9716 5524 9725 5564
rect 12076 5524 12884 5564
rect 12844 5480 12884 5524
rect 13638 5480 13728 5500
rect 0 5440 1180 5480
rect 1220 5440 1229 5480
rect 1699 5440 1708 5480
rect 1748 5440 2900 5480
rect 4204 5440 6316 5480
rect 6356 5440 6365 5480
rect 8323 5440 8332 5480
rect 8372 5440 11836 5480
rect 11876 5440 11885 5480
rect 12844 5440 13728 5480
rect 0 5420 90 5440
rect 2860 5396 2900 5440
rect 13638 5420 13728 5440
rect 2860 5356 6220 5396
rect 6260 5356 6988 5396
rect 7028 5356 7037 5396
rect 3679 5272 3688 5312
rect 3728 5272 3770 5312
rect 3810 5272 3852 5312
rect 3892 5272 3934 5312
rect 3974 5272 4016 5312
rect 4056 5272 4065 5312
rect 4588 5188 9004 5228
rect 9044 5188 9053 5228
rect 1097 4936 1228 4976
rect 1268 4936 1277 4976
rect 3532 4936 4492 4976
rect 4532 4936 4541 4976
rect 3532 4892 3572 4936
rect 2275 4852 2284 4892
rect 2324 4852 2956 4892
rect 2996 4852 3005 4892
rect 3907 4852 3916 4892
rect 3956 4852 4108 4892
rect 4148 4852 4157 4892
rect 3532 4843 3572 4852
rect 4588 4808 4628 5188
rect 13638 5144 13728 5164
rect 5347 5104 5356 5144
rect 5396 5104 6700 5144
rect 6740 5104 6749 5144
rect 9811 5104 9820 5144
rect 9860 5104 9964 5144
rect 10004 5104 10013 5144
rect 12460 5104 13728 5144
rect 5827 5020 5836 5060
rect 5876 5020 6836 5060
rect 7363 5020 7372 5060
rect 7412 5020 12220 5060
rect 12260 5020 12269 5060
rect 5164 4936 5356 4976
rect 5396 4936 5405 4976
rect 5635 4936 5644 4976
rect 5684 4936 5780 4976
rect 6115 4936 6124 4976
rect 6164 4936 6644 4976
rect 5164 4892 5204 4936
rect 5740 4892 5780 4936
rect 5164 4843 5204 4852
rect 5260 4852 5635 4892
rect 5675 4852 5684 4892
rect 5731 4852 5740 4892
rect 5780 4852 5789 4892
rect 6211 4852 6220 4892
rect 6260 4852 6269 4892
rect 3628 4768 4628 4808
rect 3628 4724 3668 4768
rect 5260 4724 5300 4852
rect 1459 4684 1468 4724
rect 1508 4684 3668 4724
rect 3715 4684 3724 4724
rect 3764 4684 5300 4724
rect 6220 4556 6260 4852
rect 6604 4640 6644 4936
rect 6700 4892 6740 4901
rect 6796 4892 6836 5020
rect 12460 4976 12500 5104
rect 13638 5084 13728 5104
rect 8009 4936 8140 4976
rect 8180 4936 8189 4976
rect 8716 4936 9004 4976
rect 9044 4936 9053 4976
rect 9475 4936 9484 4976
rect 9524 4936 9580 4976
rect 9620 4936 9655 4976
rect 9833 4936 9916 4976
rect 9956 4936 9964 4976
rect 10004 4936 10013 4976
rect 10147 4936 10156 4976
rect 10196 4936 10205 4976
rect 12067 4936 12076 4976
rect 12116 4936 12125 4976
rect 12451 4936 12460 4976
rect 12500 4936 12509 4976
rect 8716 4892 8756 4936
rect 10156 4892 10196 4936
rect 6796 4852 7188 4892
rect 7228 4852 7237 4892
rect 7459 4852 7468 4892
rect 7508 4852 7651 4892
rect 7691 4852 7700 4892
rect 7747 4852 7756 4892
rect 7796 4852 7927 4892
rect 8105 4852 8236 4892
rect 8276 4852 8285 4892
rect 9091 4852 9100 4892
rect 9140 4852 9204 4892
rect 9244 4852 9271 4892
rect 9388 4852 10196 4892
rect 6700 4808 6740 4852
rect 8236 4808 8276 4852
rect 8716 4843 8756 4852
rect 6700 4768 8276 4808
rect 9388 4724 9428 4852
rect 12076 4808 12116 4936
rect 13638 4808 13728 4828
rect 12076 4768 13728 4808
rect 13638 4748 13728 4768
rect 7241 4684 7372 4724
rect 7412 4684 7421 4724
rect 9379 4684 9388 4724
rect 9428 4684 9437 4724
rect 9484 4684 11836 4724
rect 11876 4684 11885 4724
rect 6604 4600 8140 4640
rect 8180 4600 8189 4640
rect 4919 4516 4928 4556
rect 4968 4516 5010 4556
rect 5050 4516 5092 4556
rect 5132 4516 5174 4556
rect 5214 4516 5256 4556
rect 5296 4516 5305 4556
rect 6220 4516 8428 4556
rect 8468 4516 8477 4556
rect 0 4472 90 4492
rect 9484 4472 9524 4684
rect 13638 4472 13728 4492
rect 0 4432 1228 4472
rect 1268 4432 1277 4472
rect 7171 4432 7180 4472
rect 7220 4432 9524 4472
rect 12451 4432 12460 4472
rect 12500 4432 13728 4472
rect 0 4412 90 4432
rect 3305 4264 3388 4304
rect 3428 4264 3436 4304
rect 3476 4264 3485 4304
rect 5347 4264 5356 4304
rect 5396 4264 5932 4304
rect 5972 4264 5981 4304
rect 6979 4264 6988 4304
rect 7028 4264 7468 4304
rect 7508 4264 7517 4304
rect 7660 4220 7700 4432
rect 13638 4412 13728 4432
rect 7843 4348 7852 4388
rect 7892 4348 9332 4388
rect 9292 4304 9332 4348
rect 8227 4264 8236 4304
rect 8276 4264 8372 4304
rect 3532 4180 3916 4220
rect 3956 4180 4108 4220
rect 4148 4180 4157 4220
rect 4483 4180 4492 4220
rect 4532 4211 5204 4220
rect 4532 4180 5164 4211
rect 3532 4136 3572 4180
rect 5513 4180 5548 4220
rect 5588 4180 5644 4220
rect 5684 4180 5693 4220
rect 6796 4211 7124 4220
rect 5164 4162 5204 4171
rect 6836 4180 7124 4211
rect 7258 4180 7267 4220
rect 7307 4180 7316 4220
rect 7363 4180 7372 4220
rect 7412 4180 7700 4220
rect 7747 4180 7756 4220
rect 7796 4180 8140 4220
rect 8180 4180 8189 4220
rect 8332 4211 8372 4264
rect 6796 4162 6836 4171
rect 1411 4096 1420 4136
rect 1460 4096 1612 4136
rect 1652 4096 1661 4136
rect 3017 4096 3148 4136
rect 3188 4096 3197 4136
rect 3523 4096 3532 4136
rect 3572 4096 3581 4136
rect 7084 4052 7124 4180
rect 7276 4136 7316 4180
rect 8332 4162 8372 4171
rect 8812 4264 9196 4304
rect 9236 4264 9245 4304
rect 9292 4264 12220 4304
rect 12260 4264 12269 4304
rect 8812 4211 8852 4264
rect 8995 4180 9004 4220
rect 9044 4211 9428 4220
rect 9044 4180 9388 4211
rect 8812 4162 8852 4171
rect 9388 4162 9428 4171
rect 9484 4180 10636 4220
rect 10676 4180 10685 4220
rect 12076 4180 12884 4220
rect 7276 4096 7468 4136
rect 7508 4096 7517 4136
rect 7843 4096 7852 4136
rect 7892 4096 8236 4136
rect 8276 4096 8285 4136
rect 9484 4052 9524 4180
rect 12076 4136 12116 4180
rect 12844 4136 12884 4180
rect 13638 4136 13728 4156
rect 11683 4096 11692 4136
rect 11732 4096 11741 4136
rect 12067 4096 12076 4136
rect 12116 4096 12125 4136
rect 12329 4096 12460 4136
rect 12500 4096 12509 4136
rect 12844 4096 13728 4136
rect 3235 4012 3244 4052
rect 3284 4012 3772 4052
rect 3812 4012 3821 4052
rect 7084 4012 8620 4052
rect 8660 4012 8669 4052
rect 8908 4012 9524 4052
rect 11692 4052 11732 4096
rect 13638 4076 13728 4096
rect 11692 4012 12652 4052
rect 12692 4012 12701 4052
rect 8908 3968 8948 4012
rect 67 3928 76 3968
rect 116 3928 1180 3968
rect 1220 3928 1229 3968
rect 6979 3928 6988 3968
rect 7028 3928 8948 3968
rect 9034 3928 9043 3968
rect 9083 3928 9676 3968
rect 9716 3928 9725 3968
rect 9955 3928 9964 3968
rect 10004 3928 11452 3968
rect 11492 3928 11501 3968
rect 11596 3928 11836 3968
rect 11876 3928 11885 3968
rect 11596 3884 11636 3928
rect 6499 3844 6508 3884
rect 6548 3844 11636 3884
rect 13638 3800 13728 3820
rect 3679 3760 3688 3800
rect 3728 3760 3770 3800
rect 3810 3760 3852 3800
rect 3892 3760 3934 3800
rect 3974 3760 4016 3800
rect 4056 3760 4065 3800
rect 4387 3760 4396 3800
rect 4436 3760 9772 3800
rect 9812 3760 9821 3800
rect 12460 3760 13728 3800
rect 7747 3676 7756 3716
rect 7796 3676 12260 3716
rect 12220 3632 12260 3676
rect 5417 3592 5548 3632
rect 5588 3592 5597 3632
rect 7171 3592 7180 3632
rect 7220 3592 7468 3632
rect 7508 3592 7517 3632
rect 8969 3592 9100 3632
rect 9140 3592 9149 3632
rect 10051 3592 10060 3632
rect 10100 3592 11836 3632
rect 11876 3592 11885 3632
rect 12211 3592 12220 3632
rect 12260 3592 12269 3632
rect 4108 3508 5356 3548
rect 5396 3508 5644 3548
rect 5684 3508 5780 3548
rect 0 3464 90 3484
rect 0 3424 76 3464
rect 116 3424 125 3464
rect 0 3404 90 3424
rect 4108 3380 4148 3508
rect 5356 3380 5396 3389
rect 5740 3380 5780 3508
rect 6988 3508 9004 3548
rect 9044 3508 9053 3548
rect 9187 3508 9196 3548
rect 9236 3508 9628 3548
rect 9668 3508 9677 3548
rect 6988 3380 7028 3508
rect 12460 3464 12500 3760
rect 13638 3740 13728 3760
rect 13638 3464 13728 3484
rect 8908 3424 9244 3464
rect 9284 3424 9293 3464
rect 9475 3424 9484 3464
rect 9524 3424 9533 3464
rect 9667 3424 9676 3464
rect 9716 3424 9868 3464
rect 9908 3424 9917 3464
rect 12067 3424 12076 3464
rect 12116 3424 12125 3464
rect 12451 3424 12460 3464
rect 12500 3424 12509 3464
rect 12643 3424 12652 3464
rect 12692 3424 13728 3464
rect 8908 3380 8948 3424
rect 2275 3340 2284 3380
rect 2324 3340 4108 3380
rect 4148 3340 4157 3380
rect 5321 3340 5356 3380
rect 5396 3340 5452 3380
rect 5492 3340 5501 3380
rect 5731 3340 5740 3380
rect 5780 3340 5789 3380
rect 7075 3340 7084 3380
rect 7124 3340 7660 3380
rect 7700 3340 7709 3380
rect 8611 3340 8620 3380
rect 8660 3340 8908 3380
rect 5356 3331 5396 3340
rect 6988 3331 7028 3340
rect 8908 3331 8948 3340
rect 9484 3296 9524 3424
rect 9004 3256 9524 3296
rect 12076 3296 12116 3424
rect 13638 3404 13728 3424
rect 12076 3256 12884 3296
rect 9004 3212 9044 3256
rect 1603 3172 1612 3212
rect 1652 3172 9044 3212
rect 12844 3128 12884 3256
rect 13638 3128 13728 3148
rect 12844 3088 13728 3128
rect 13638 3068 13728 3088
rect 4919 3004 4928 3044
rect 4968 3004 5010 3044
rect 5050 3004 5092 3044
rect 5132 3004 5174 3044
rect 5214 3004 5256 3044
rect 5296 3004 5305 3044
rect 8105 2836 8188 2876
rect 8228 2836 8236 2876
rect 8276 2836 8285 2876
rect 12211 2836 12220 2876
rect 12260 2836 13516 2876
rect 13556 2836 13565 2876
rect 13638 2792 13728 2812
rect 7219 2752 7228 2792
rect 7268 2752 13228 2792
rect 13268 2752 13277 2792
rect 13516 2752 13728 2792
rect 13516 2624 13556 2752
rect 13638 2732 13728 2752
rect 1411 2584 1420 2624
rect 1460 2584 2572 2624
rect 2612 2584 2621 2624
rect 5155 2584 5164 2624
rect 5204 2584 5356 2624
rect 5396 2584 5405 2624
rect 6857 2584 6988 2624
rect 7028 2584 7037 2624
rect 7363 2584 7372 2624
rect 7412 2584 7948 2624
rect 7988 2584 7997 2624
rect 12451 2584 12460 2624
rect 12500 2584 13556 2624
rect 0 2456 90 2476
rect 0 2416 1180 2456
rect 1220 2416 1229 2456
rect 5395 2416 5404 2456
rect 5444 2416 5740 2456
rect 5780 2416 5789 2456
rect 0 2396 90 2416
rect 3679 2248 3688 2288
rect 3728 2248 3770 2288
rect 3810 2248 3852 2288
rect 3892 2248 3934 2288
rect 3974 2248 4016 2288
rect 4056 2248 4065 2288
rect 1459 2080 1468 2120
rect 1508 2080 4780 2120
rect 4820 2080 4829 2120
rect 67 1912 76 1952
rect 116 1912 1228 1952
rect 1268 1912 1277 1952
rect 4919 1492 4928 1532
rect 4968 1492 5010 1532
rect 5050 1492 5092 1532
rect 5132 1492 5174 1532
rect 5214 1492 5256 1532
rect 5296 1492 5305 1532
rect 0 1448 90 1468
rect 0 1408 76 1448
rect 116 1408 125 1448
rect 2179 1408 2188 1448
rect 2228 1408 4108 1448
rect 4148 1408 4157 1448
rect 0 1388 90 1408
<< via2 >>
rect 4928 46852 4968 46892
rect 5010 46852 5050 46892
rect 5092 46852 5132 46892
rect 5174 46852 5214 46892
rect 5256 46852 5296 46892
rect 1228 46768 1268 46808
rect 6892 46768 6932 46808
rect 1612 46684 1652 46724
rect 2188 46684 2228 46724
rect 2764 46684 2804 46724
rect 3340 46684 3380 46724
rect 3916 46684 3956 46724
rect 4492 46684 4532 46724
rect 5356 46684 5396 46724
rect 5644 46684 5684 46724
rect 6220 46684 6260 46724
rect 6796 46684 6836 46724
rect 7372 46684 7412 46724
rect 7948 46684 7988 46724
rect 8524 46684 8564 46724
rect 9100 46684 9140 46724
rect 9676 46684 9716 46724
rect 10252 46684 10292 46724
rect 10828 46684 10868 46724
rect 11404 46684 11444 46724
rect 11020 46600 11060 46640
rect 10732 46516 10772 46556
rect 652 46432 692 46472
rect 1900 46432 1940 46472
rect 2476 46432 2516 46472
rect 5932 46432 5972 46472
rect 6508 46432 6548 46472
rect 7660 46432 7700 46472
rect 9388 46432 9428 46472
rect 10348 46432 10388 46472
rect 10828 46432 10868 46472
rect 11116 46432 11156 46472
rect 11308 46432 11348 46472
rect 12748 46432 12788 46472
rect 4204 46348 4244 46388
rect 4684 46264 4724 46304
rect 8620 46348 8660 46388
rect 11212 46348 11252 46388
rect 10060 46264 10100 46304
rect 9964 46180 10004 46220
rect 12364 46264 12404 46304
rect 13132 46264 13172 46304
rect 3688 46096 3728 46136
rect 3770 46096 3810 46136
rect 3852 46096 3892 46136
rect 3934 46096 3974 46136
rect 4016 46096 4056 46136
rect 6700 46096 6740 46136
rect 12556 46012 12596 46052
rect 1036 45928 1076 45968
rect 11116 45928 11156 45968
rect 11980 45844 12020 45884
rect 652 45760 692 45800
rect 1228 45760 1268 45800
rect 1804 45760 1844 45800
rect 10540 45760 10580 45800
rect 11500 45760 11540 45800
rect 11788 45760 11828 45800
rect 12172 45760 12212 45800
rect 10252 45676 10292 45716
rect 11692 45592 11732 45632
rect 3436 45508 3476 45548
rect 12268 45508 12308 45548
rect 13036 45508 13076 45548
rect 4928 45340 4968 45380
rect 5010 45340 5050 45380
rect 5092 45340 5132 45380
rect 5174 45340 5214 45380
rect 5256 45340 5296 45380
rect 5932 45172 5972 45212
rect 8620 45172 8660 45212
rect 10060 45172 10100 45212
rect 10828 45172 10868 45212
rect 6508 45088 6548 45128
rect 10348 45088 10388 45128
rect 12364 45088 12404 45128
rect 10924 45004 10964 45044
rect 76 44920 116 44960
rect 5452 44920 5492 44960
rect 8908 44920 8948 44960
rect 10636 44920 10676 44960
rect 11212 44920 11252 44960
rect 11500 44920 11540 44960
rect 11884 44920 11924 44960
rect 12364 44920 12404 44960
rect 5548 44836 5588 44876
rect 76 44752 116 44792
rect 2668 44752 2708 44792
rect 3688 44584 3728 44624
rect 3770 44584 3810 44624
rect 3852 44584 3892 44624
rect 3934 44584 3974 44624
rect 4016 44584 4056 44624
rect 9388 44416 9428 44456
rect 10732 44416 10772 44456
rect 11020 44416 11060 44456
rect 13132 44416 13172 44456
rect 9964 44332 10004 44372
rect 76 44248 116 44288
rect 10732 44248 10772 44288
rect 11116 44248 11156 44288
rect 11500 44248 11540 44288
rect 11884 44248 11924 44288
rect 5356 44164 5396 44204
rect 12268 44080 12308 44120
rect 6124 43996 6164 44036
rect 13132 43996 13172 44036
rect 4928 43828 4968 43868
rect 5010 43828 5050 43868
rect 5092 43828 5132 43868
rect 5174 43828 5214 43868
rect 5256 43828 5296 43868
rect 76 43744 116 43784
rect 13036 43744 13076 43784
rect 7660 43660 7700 43700
rect 8044 43492 8084 43532
rect 1228 43408 1268 43448
rect 8620 43408 8660 43448
rect 11500 43408 11540 43448
rect 7852 43324 7892 43364
rect 4588 43240 4628 43280
rect 6508 43240 6548 43280
rect 12364 43240 12404 43280
rect 13036 43240 13076 43280
rect 3688 43072 3728 43112
rect 3770 43072 3810 43112
rect 3852 43072 3892 43112
rect 3934 43072 3974 43112
rect 4016 43072 4056 43112
rect 11308 42904 11348 42944
rect 11692 42904 11732 42944
rect 10540 42820 10580 42860
rect 1228 42736 1268 42776
rect 11020 42736 11060 42776
rect 11596 42736 11636 42776
rect 11980 42736 12020 42776
rect 13132 42736 13172 42776
rect 7084 42652 7124 42692
rect 13132 42484 13172 42524
rect 12364 42400 12404 42440
rect 4928 42316 4968 42356
rect 5010 42316 5050 42356
rect 5092 42316 5132 42356
rect 5174 42316 5214 42356
rect 5256 42316 5296 42356
rect 13036 42064 13076 42104
rect 76 41896 116 41936
rect 5836 41896 5876 41936
rect 2284 41812 2324 41852
rect 10060 41812 10100 41852
rect 76 41728 116 41768
rect 12940 41728 12980 41768
rect 13132 41728 13172 41768
rect 3688 41560 3728 41600
rect 3770 41560 3810 41600
rect 3852 41560 3892 41600
rect 3934 41560 3974 41600
rect 4016 41560 4056 41600
rect 13612 41560 13652 41600
rect 13612 41392 13652 41432
rect 76 41224 116 41264
rect 12460 41224 12500 41264
rect 2572 41140 2612 41180
rect 10828 41140 10868 41180
rect 2956 40972 2996 41012
rect 13132 40972 13172 41012
rect 12844 40888 12884 40928
rect 4928 40804 4968 40844
rect 5010 40804 5050 40844
rect 5092 40804 5132 40844
rect 5174 40804 5214 40844
rect 5256 40804 5296 40844
rect 76 40720 116 40760
rect 12940 40720 12980 40760
rect 13228 40468 13268 40508
rect 1228 40384 1268 40424
rect 6220 40384 6260 40424
rect 12556 40384 12596 40424
rect 12844 40384 12884 40424
rect 5740 40300 5780 40340
rect 13420 40300 13460 40340
rect 12364 40216 12404 40256
rect 3688 40048 3728 40088
rect 3770 40048 3810 40088
rect 3852 40048 3892 40088
rect 3934 40048 3974 40088
rect 4016 40048 4056 40088
rect 9484 39796 9524 39836
rect 1228 39712 1268 39752
rect 13132 39712 13172 39752
rect 6124 39628 6164 39668
rect 6604 39628 6644 39668
rect 7276 39628 7316 39668
rect 8332 39628 8372 39668
rect 8908 39628 8948 39668
rect 7372 39460 7412 39500
rect 9004 39460 9044 39500
rect 4928 39292 4968 39332
rect 5010 39292 5050 39332
rect 5092 39292 5132 39332
rect 5174 39292 5214 39332
rect 5256 39292 5296 39332
rect 11500 39628 11540 39668
rect 13516 39628 13556 39668
rect 13324 39544 13364 39584
rect 11980 39460 12020 39500
rect 13132 39460 13172 39500
rect 12076 39124 12116 39164
rect 12364 39124 12404 39164
rect 5740 39040 5780 39080
rect 9676 39040 9716 39080
rect 6316 38956 6356 38996
rect 6796 38956 6836 38996
rect 7660 38956 7700 38996
rect 76 38872 116 38912
rect 2764 38872 2804 38912
rect 4108 38872 4148 38912
rect 4396 38872 4436 38912
rect 8140 38956 8180 38996
rect 10348 38956 10388 38996
rect 12940 38956 12980 38996
rect 7468 38872 7508 38912
rect 8812 38872 8852 38912
rect 9388 38872 9428 38912
rect 9772 38872 9812 38912
rect 9964 38872 10004 38912
rect 11116 38872 11156 38912
rect 11596 38872 11636 38912
rect 11884 38872 11924 38912
rect 12364 38872 12404 38912
rect 13036 38872 13076 38912
rect 13612 38872 13652 38912
rect 8908 38788 8948 38828
rect 76 38704 116 38744
rect 3688 38536 3728 38576
rect 3770 38536 3810 38576
rect 3852 38536 3892 38576
rect 3934 38536 3974 38576
rect 4016 38536 4056 38576
rect 11788 38704 11828 38744
rect 13612 38704 13652 38744
rect 76 38200 116 38240
rect 6316 38368 6356 38408
rect 8332 38368 8372 38408
rect 11980 38368 12020 38408
rect 7372 38200 7412 38240
rect 7660 38200 7700 38240
rect 3820 38116 3860 38156
rect 4108 38116 4148 38156
rect 8908 38200 8948 38240
rect 11020 38200 11060 38240
rect 11884 38200 11924 38240
rect 7468 38116 7508 38156
rect 8236 38116 8276 38156
rect 1516 37948 1556 37988
rect 2668 37948 2708 37988
rect 7180 38032 7220 38072
rect 7276 37948 7316 37988
rect 8140 37948 8180 37988
rect 11692 38116 11732 38156
rect 11980 38032 12020 38072
rect 12652 38032 12692 38072
rect 13420 38032 13460 38072
rect 9388 37948 9428 37988
rect 11116 37948 11156 37988
rect 12364 37948 12404 37988
rect 12844 37948 12884 37988
rect 6604 37864 6644 37904
rect 4928 37780 4968 37820
rect 5010 37780 5050 37820
rect 5092 37780 5132 37820
rect 5174 37780 5214 37820
rect 5256 37780 5296 37820
rect 76 37696 116 37736
rect 8812 37612 8852 37652
rect 4108 37528 4148 37568
rect 3340 37444 3380 37484
rect 3820 37444 3860 37484
rect 4396 37444 4436 37484
rect 6028 37444 6068 37484
rect 6988 37444 7028 37484
rect 7276 37444 7316 37484
rect 7468 37444 7508 37484
rect 12076 37696 12116 37736
rect 11020 37612 11060 37652
rect 9004 37444 9044 37484
rect 9292 37444 9332 37484
rect 1228 37360 1268 37400
rect 7756 37360 7796 37400
rect 3148 37192 3188 37232
rect 5740 37192 5780 37232
rect 7756 37192 7796 37232
rect 8236 37192 8276 37232
rect 9292 37192 9332 37232
rect 10444 37444 10484 37484
rect 11308 37360 11348 37400
rect 11884 37360 11924 37400
rect 13324 37360 13364 37400
rect 10060 37276 10100 37316
rect 13420 37276 13460 37316
rect 9772 37192 9812 37232
rect 11404 37192 11444 37232
rect 11980 37192 12020 37232
rect 13612 37192 13652 37232
rect 11020 37108 11060 37148
rect 3688 37024 3728 37064
rect 3770 37024 3810 37064
rect 3852 37024 3892 37064
rect 3934 37024 3974 37064
rect 4016 37024 4056 37064
rect 11212 37024 11252 37064
rect 11788 37024 11828 37064
rect 2188 36940 2228 36980
rect 6412 36856 6452 36896
rect 10828 36856 10868 36896
rect 3340 36772 3380 36812
rect 1228 36688 1268 36728
rect 9580 36688 9620 36728
rect 10636 36688 10676 36728
rect 13132 36688 13172 36728
rect 4396 36604 4436 36644
rect 6028 36604 6068 36644
rect 10732 36604 10772 36644
rect 4300 36520 4340 36560
rect 4588 36436 4628 36476
rect 6220 36436 6260 36476
rect 9292 36520 9332 36560
rect 10540 36520 10580 36560
rect 8620 36436 8660 36476
rect 11404 36436 11444 36476
rect 13324 36436 13364 36476
rect 4300 36352 4340 36392
rect 4928 36268 4968 36308
rect 5010 36268 5050 36308
rect 5092 36268 5132 36308
rect 5174 36268 5214 36308
rect 5256 36268 5296 36308
rect 12748 36352 12788 36392
rect 12940 36352 12980 36392
rect 10156 36268 10196 36308
rect 10540 36268 10580 36308
rect 6988 36100 7028 36140
rect 11308 36100 11348 36140
rect 12076 36016 12116 36056
rect 6028 35932 6068 35972
rect 10156 35932 10187 35972
rect 10187 35932 10196 35972
rect 10444 35932 10484 35972
rect 11020 35932 11060 35972
rect 11404 35932 11444 35972
rect 76 35848 116 35888
rect 2476 35848 2516 35888
rect 4684 35848 4724 35888
rect 6604 35848 6644 35888
rect 9196 35848 9236 35888
rect 10540 35848 10580 35888
rect 10828 35848 10868 35888
rect 11212 35848 11252 35888
rect 12076 35848 12116 35888
rect 4396 35764 4436 35804
rect 9676 35764 9716 35804
rect 76 35680 116 35720
rect 2668 35680 2708 35720
rect 9292 35680 9332 35720
rect 9964 35680 10004 35720
rect 3688 35512 3728 35552
rect 3770 35512 3810 35552
rect 3852 35512 3892 35552
rect 3934 35512 3974 35552
rect 4016 35512 4056 35552
rect 9196 35344 9236 35384
rect 9964 35428 10004 35468
rect 11884 35428 11924 35468
rect 12556 35680 12596 35720
rect 12748 35680 12788 35720
rect 8524 35260 8564 35300
rect 76 35176 116 35216
rect 4108 35176 4148 35216
rect 4396 35176 4436 35216
rect 4684 35092 4724 35132
rect 6220 35092 6260 35132
rect 7276 35092 7316 35132
rect 7660 35092 7700 35132
rect 8236 35092 8276 35132
rect 8620 35092 8628 35132
rect 8628 35092 8660 35132
rect 9484 35092 9524 35132
rect 10540 35092 10580 35132
rect 11404 35092 11444 35132
rect 5932 35008 5972 35048
rect 6604 35008 6644 35048
rect 10732 35008 10772 35048
rect 11212 35008 11252 35048
rect 12364 35008 12404 35048
rect 2284 34924 2324 34964
rect 6124 34924 6164 34964
rect 9388 34924 9428 34964
rect 10060 34840 10100 34880
rect 4928 34756 4968 34796
rect 5010 34756 5050 34796
rect 5092 34756 5132 34796
rect 5174 34756 5214 34796
rect 5256 34756 5296 34796
rect 76 34672 116 34712
rect 13036 34672 13076 34712
rect 9484 34588 9524 34628
rect 4108 34504 4148 34544
rect 4684 34420 4724 34460
rect 1228 34336 1268 34376
rect 6604 34336 6644 34376
rect 3052 34168 3092 34208
rect 3688 34000 3728 34040
rect 3770 34000 3810 34040
rect 3852 34000 3892 34040
rect 3934 34000 3974 34040
rect 4016 34000 4056 34040
rect 4108 33748 4148 33788
rect 1228 33664 1268 33704
rect 3244 33580 3284 33620
rect 4108 33580 4148 33620
rect 7948 34420 7988 34460
rect 9388 34451 9428 34460
rect 9388 34420 9428 34451
rect 10060 34420 10100 34460
rect 10636 34420 10676 34460
rect 8524 34336 8564 34376
rect 9292 34336 9332 34376
rect 12268 34336 12308 34376
rect 12652 34336 12692 34376
rect 7276 34252 7316 34292
rect 10732 34168 10772 34208
rect 12748 34252 12788 34292
rect 13228 34168 13268 34208
rect 9964 34084 10004 34124
rect 11980 34000 12020 34040
rect 11308 33748 11348 33788
rect 6604 33664 6644 33704
rect 7276 33664 7316 33704
rect 7660 33580 7700 33620
rect 10156 33664 10196 33704
rect 12268 33664 12308 33704
rect 12844 33664 12884 33704
rect 9100 33580 9140 33620
rect 10444 33580 10484 33620
rect 11212 33580 11252 33620
rect 6412 33496 6452 33536
rect 9292 33496 9332 33536
rect 11788 33496 11828 33536
rect 8524 33412 8564 33452
rect 9004 33412 9044 33452
rect 11212 33412 11252 33452
rect 12268 33412 12308 33452
rect 13036 33412 13076 33452
rect 6988 33328 7028 33368
rect 13420 33328 13460 33368
rect 4928 33244 4968 33284
rect 5010 33244 5050 33284
rect 5092 33244 5132 33284
rect 5174 33244 5214 33284
rect 5256 33244 5296 33284
rect 9196 33244 9236 33284
rect 10444 33244 10484 33284
rect 8236 33076 8276 33116
rect 11692 33076 11732 33116
rect 9580 32992 9620 33032
rect 13612 32992 13652 33032
rect 5452 32908 5492 32948
rect 76 32824 116 32864
rect 3532 32824 3572 32864
rect 4108 32824 4148 32864
rect 3148 32740 3188 32780
rect 6124 32939 6164 32948
rect 6124 32908 6164 32939
rect 8716 32908 8756 32948
rect 10828 32908 10868 32948
rect 11212 32939 11252 32948
rect 11212 32908 11252 32939
rect 4780 32824 4820 32864
rect 5356 32824 5396 32864
rect 7564 32824 7604 32864
rect 7756 32824 7796 32864
rect 9196 32824 9236 32864
rect 10156 32824 10196 32864
rect 10636 32824 10676 32864
rect 11404 32824 11444 32864
rect 4876 32740 4916 32780
rect 7276 32740 7316 32780
rect 76 32656 116 32696
rect 2860 32656 2900 32696
rect 5644 32656 5684 32696
rect 9580 32656 9620 32696
rect 10636 32656 10676 32696
rect 11692 32656 11732 32696
rect 11980 32656 12020 32696
rect 12268 32656 12308 32696
rect 12556 32656 12596 32696
rect 7084 32572 7124 32612
rect 3688 32488 3728 32528
rect 3770 32488 3810 32528
rect 3852 32488 3892 32528
rect 3934 32488 3974 32528
rect 4016 32488 4056 32528
rect 10156 32488 10196 32528
rect 11404 32488 11444 32528
rect 3724 32320 3764 32360
rect 8236 32404 8276 32444
rect 9868 32320 9908 32360
rect 13324 32320 13364 32360
rect 5452 32236 5492 32276
rect 8716 32236 8756 32276
rect 76 32152 116 32192
rect 4108 32152 4148 32192
rect 4396 32152 4436 32192
rect 4780 32152 4820 32192
rect 6316 32152 6356 32192
rect 11308 32152 11348 32192
rect 2668 32068 2708 32108
rect 4300 32068 4340 32108
rect 5356 32068 5396 32108
rect 8716 32068 8756 32108
rect 8908 32068 8948 32108
rect 10540 32068 10571 32108
rect 10571 32068 10580 32108
rect 3724 31984 3764 32024
rect 4876 31984 4916 32024
rect 3436 31900 3476 31940
rect 4012 31900 4052 31940
rect 7276 31984 7316 32024
rect 10444 31984 10484 32024
rect 12460 31984 12500 32024
rect 5164 31900 5204 31940
rect 9196 31900 9236 31940
rect 13132 31900 13172 31940
rect 10924 31816 10964 31856
rect 4928 31732 4968 31772
rect 5010 31732 5050 31772
rect 5092 31732 5132 31772
rect 5174 31732 5214 31772
rect 5256 31732 5296 31772
rect 76 31648 116 31688
rect 4300 31564 4340 31604
rect 12748 31648 12788 31688
rect 6316 31564 6356 31604
rect 6892 31564 6932 31604
rect 8236 31564 8276 31604
rect 9676 31564 9716 31604
rect 4588 31480 4628 31520
rect 8908 31480 8948 31520
rect 3244 31396 3284 31436
rect 4108 31427 4148 31436
rect 4108 31396 4148 31427
rect 4876 31396 4916 31436
rect 5260 31396 5300 31436
rect 5740 31396 5780 31436
rect 8620 31396 8660 31436
rect 9868 31396 9908 31436
rect 1228 31312 1268 31352
rect 4588 31312 4628 31352
rect 8716 31312 8756 31352
rect 9100 31312 9140 31352
rect 9292 31312 9332 31352
rect 11500 31312 11540 31352
rect 11788 31312 11828 31352
rect 13228 31312 13268 31352
rect 5068 31228 5108 31268
rect 7756 31228 7796 31268
rect 8812 31228 8852 31268
rect 13324 31228 13364 31268
rect 5260 31144 5300 31184
rect 6316 31144 6356 31184
rect 6604 31144 6644 31184
rect 6892 31144 6932 31184
rect 7372 31144 7412 31184
rect 11020 31144 11060 31184
rect 11980 31144 12020 31184
rect 13228 31144 13268 31184
rect 3688 30976 3728 31016
rect 3770 30976 3810 31016
rect 3852 30976 3892 31016
rect 3934 30976 3974 31016
rect 4016 30976 4056 31016
rect 7276 30976 7316 31016
rect 12364 30976 12404 31016
rect 7852 30892 7892 30932
rect 3244 30808 3284 30848
rect 4108 30808 4148 30848
rect 4300 30808 4340 30848
rect 8908 30808 8948 30848
rect 9868 30808 9908 30848
rect 11596 30808 11636 30848
rect 1228 30640 1268 30680
rect 3724 30724 3764 30764
rect 4876 30724 4916 30764
rect 7084 30724 7124 30764
rect 3244 30640 3284 30680
rect 6316 30640 6356 30680
rect 7756 30640 7796 30680
rect 8428 30640 8468 30680
rect 10828 30724 10868 30764
rect 10540 30640 10580 30680
rect 10924 30640 10964 30680
rect 11596 30640 11636 30680
rect 12364 30640 12404 30680
rect 13036 30640 13076 30680
rect 4012 30556 4052 30596
rect 5068 30556 5108 30596
rect 6604 30556 6644 30596
rect 7468 30556 7508 30596
rect 8620 30556 8660 30596
rect 9292 30556 9332 30596
rect 11308 30556 11348 30596
rect 3148 30472 3188 30512
rect 4876 30472 4916 30512
rect 10156 30472 10196 30512
rect 12748 30472 12788 30512
rect 4108 30388 4148 30428
rect 4588 30388 4628 30428
rect 6412 30388 6452 30428
rect 8044 30388 8084 30428
rect 11884 30388 11924 30428
rect 13036 30388 13076 30428
rect 1804 30304 1844 30344
rect 5740 30304 5780 30344
rect 12268 30304 12308 30344
rect 4780 30220 4820 30260
rect 4928 30220 4968 30260
rect 5010 30220 5050 30260
rect 5092 30220 5132 30260
rect 5174 30220 5214 30260
rect 5256 30220 5296 30260
rect 10828 30220 10868 30260
rect 6604 30136 6644 30176
rect 9100 30136 9140 30176
rect 10732 30136 10772 30176
rect 10924 30136 10964 30176
rect 4876 30052 4916 30092
rect 4972 29884 5012 29924
rect 7468 30052 7508 30092
rect 10252 30052 10292 30092
rect 5356 29968 5396 30008
rect 5740 29968 5780 30008
rect 9388 29968 9428 30008
rect 10444 29968 10484 30008
rect 10732 29968 10772 30008
rect 12556 29968 12596 30008
rect 5644 29915 5684 29924
rect 5644 29884 5684 29915
rect 7756 29884 7796 29924
rect 8332 29884 8372 29924
rect 10924 29884 10964 29924
rect 76 29800 116 29840
rect 4108 29800 4148 29840
rect 4492 29800 4532 29840
rect 7468 29800 7508 29840
rect 9388 29800 9428 29840
rect 9772 29800 9812 29840
rect 10060 29800 10100 29840
rect 10828 29800 10868 29840
rect 1036 29716 1076 29756
rect 4012 29716 4052 29756
rect 7756 29716 7796 29756
rect 76 29632 116 29672
rect 5356 29632 5396 29672
rect 10636 29632 10676 29672
rect 2860 29464 2900 29504
rect 3052 29464 3092 29504
rect 3688 29464 3728 29504
rect 3770 29464 3810 29504
rect 3852 29464 3892 29504
rect 3934 29464 3974 29504
rect 4016 29464 4056 29504
rect 4972 29464 5012 29504
rect 6316 29464 6356 29504
rect 10156 29380 10196 29420
rect 10924 29380 10964 29420
rect 1996 29296 2036 29336
rect 2572 29296 2612 29336
rect 5644 29296 5684 29336
rect 6700 29296 6740 29336
rect 10060 29296 10100 29336
rect 9388 29212 9428 29252
rect 9580 29212 9620 29252
rect 76 29128 116 29168
rect 2860 29128 2900 29168
rect 5356 29128 5396 29168
rect 5740 29128 5780 29168
rect 8140 29128 8180 29168
rect 9100 29128 9140 29168
rect 10156 29128 10196 29168
rect 10828 29128 10868 29168
rect 3148 29044 3188 29084
rect 4396 29044 4436 29084
rect 7756 29044 7796 29084
rect 10636 29044 10676 29084
rect 11020 29044 11060 29084
rect 12172 29044 12212 29084
rect 9676 28960 9716 29000
rect 10060 28960 10100 29000
rect 11980 28960 12020 29000
rect 8620 28876 8660 28916
rect 10156 28876 10196 28916
rect 11020 28876 11060 28916
rect 11596 28876 11636 28916
rect 12364 28876 12404 28916
rect 13132 28876 13172 28916
rect 6316 28792 6356 28832
rect 10060 28792 10100 28832
rect 4928 28708 4968 28748
rect 5010 28708 5050 28748
rect 5092 28708 5132 28748
rect 5174 28708 5214 28748
rect 5256 28708 5296 28748
rect 76 28624 116 28664
rect 7276 28624 7316 28664
rect 10540 28624 10580 28664
rect 11884 28624 11924 28664
rect 3436 28540 3476 28580
rect 4108 28540 4148 28580
rect 8908 28540 8948 28580
rect 2668 28456 2708 28496
rect 8620 28456 8660 28496
rect 9388 28456 9428 28496
rect 9868 28456 9908 28496
rect 2284 28372 2324 28412
rect 2476 28372 2516 28412
rect 4396 28372 4436 28412
rect 9580 28372 9620 28412
rect 10156 28403 10196 28412
rect 10156 28372 10196 28403
rect 10540 28372 10580 28412
rect 11596 28372 11636 28412
rect 1228 28288 1268 28328
rect 8428 28288 8468 28328
rect 10060 28288 10100 28328
rect 13324 28288 13364 28328
rect 10924 28204 10964 28244
rect 11980 28120 12020 28160
rect 3688 27952 3728 27992
rect 3770 27952 3810 27992
rect 3852 27952 3892 27992
rect 3934 27952 3974 27992
rect 4016 27952 4056 27992
rect 9484 28036 9524 28076
rect 13228 27952 13268 27992
rect 9772 27700 9812 27740
rect 1228 27616 1268 27656
rect 8908 27616 8948 27656
rect 4588 27532 4628 27572
rect 5548 27532 5588 27572
rect 6700 27532 6740 27572
rect 9772 27532 9812 27572
rect 11884 27784 11924 27824
rect 11596 27700 11636 27740
rect 12748 27616 12788 27656
rect 11596 27532 11636 27572
rect 12268 27532 12308 27572
rect 10252 27448 10292 27488
rect 5932 27364 5972 27404
rect 10732 27364 10772 27404
rect 10348 27280 10388 27320
rect 13036 27280 13076 27320
rect 4928 27196 4968 27236
rect 5010 27196 5050 27236
rect 5092 27196 5132 27236
rect 5174 27196 5214 27236
rect 5256 27196 5296 27236
rect 10060 27196 10100 27236
rect 11692 27196 11732 27236
rect 11884 27196 11924 27236
rect 8716 27112 8756 27152
rect 13324 27112 13364 27152
rect 5548 27028 5588 27068
rect 6988 27028 7028 27068
rect 2668 26860 2708 26900
rect 3436 26860 3476 26900
rect 11500 27028 11540 27068
rect 9676 26944 9716 26984
rect 12364 26944 12404 26984
rect 4684 26860 4724 26900
rect 5548 26860 5588 26900
rect 5932 26891 5972 26900
rect 5932 26860 5972 26891
rect 4300 26776 4340 26816
rect 4972 26776 5012 26816
rect 3688 26440 3728 26480
rect 3770 26440 3810 26480
rect 3852 26440 3892 26480
rect 3934 26440 3974 26480
rect 4016 26440 4056 26480
rect 6412 26860 6452 26900
rect 6796 26860 6836 26900
rect 7756 26860 7796 26900
rect 7276 26776 7316 26816
rect 8140 26776 8180 26816
rect 9772 26776 9812 26816
rect 11020 26860 11060 26900
rect 11980 26860 12020 26900
rect 13324 26860 13364 26900
rect 11692 26776 11732 26816
rect 11884 26776 11924 26816
rect 10924 26692 10964 26732
rect 13228 26692 13268 26732
rect 6988 26356 7028 26396
rect 7660 26356 7700 26396
rect 8524 26356 8564 26396
rect 13132 26608 13172 26648
rect 10348 26356 10388 26396
rect 6316 26272 6356 26312
rect 4588 26188 4628 26228
rect 7276 26188 7316 26228
rect 6700 26104 6740 26144
rect 11884 26272 11924 26312
rect 10060 26188 10100 26228
rect 2476 26020 2516 26060
rect 4108 26020 4148 26060
rect 5644 26020 5684 26060
rect 6988 26020 7028 26060
rect 7660 26020 7700 26060
rect 8332 26020 8372 26060
rect 11404 26188 11444 26228
rect 13036 26272 13076 26312
rect 10060 26020 10100 26060
rect 12076 26020 12116 26060
rect 1228 25936 1268 25976
rect 2668 25936 2708 25976
rect 8716 25936 8756 25976
rect 10732 25936 10772 25976
rect 11884 25936 11924 25976
rect 13132 25936 13172 25976
rect 2956 25852 2996 25892
rect 8620 25852 8660 25892
rect 10252 25852 10292 25892
rect 4928 25684 4968 25724
rect 5010 25684 5050 25724
rect 5092 25684 5132 25724
rect 5174 25684 5214 25724
rect 5256 25684 5296 25724
rect 9292 25600 9332 25640
rect 9772 25516 9812 25556
rect 13132 25516 13172 25556
rect 7468 25432 7508 25472
rect 2668 25348 2708 25388
rect 4108 25348 4148 25388
rect 5644 25348 5684 25388
rect 2284 25096 2324 25136
rect 2572 25096 2612 25136
rect 7660 25348 7700 25388
rect 8140 25348 8180 25388
rect 8716 25348 8756 25388
rect 9388 25348 9428 25388
rect 9580 25348 9620 25388
rect 11308 25348 11348 25388
rect 12364 25348 12404 25388
rect 9100 25264 9131 25304
rect 9131 25264 9140 25304
rect 9292 25264 9332 25304
rect 8620 25180 8660 25220
rect 9772 25180 9812 25220
rect 7468 25096 7508 25136
rect 7756 25096 7796 25136
rect 11116 25096 11156 25136
rect 8236 25012 8276 25052
rect 3688 24928 3728 24968
rect 3770 24928 3810 24968
rect 3852 24928 3892 24968
rect 3934 24928 3974 24968
rect 4016 24928 4056 24968
rect 9676 24844 9716 24884
rect 9100 24760 9140 24800
rect 12076 24760 12116 24800
rect 13036 24760 13076 24800
rect 7756 24676 7796 24716
rect 8044 24676 8084 24716
rect 2092 24592 2132 24632
rect 4108 24592 4148 24632
rect 7276 24592 7316 24632
rect 8236 24592 8276 24632
rect 12460 24592 12500 24632
rect 2668 24508 2708 24548
rect 3148 24508 3188 24548
rect 7180 24508 7220 24548
rect 7948 24508 7988 24548
rect 8332 24508 8372 24548
rect 8620 24508 8660 24548
rect 11308 24508 11348 24548
rect 11596 24508 11636 24548
rect 6604 24424 6644 24464
rect 10252 24340 10292 24380
rect 12844 24256 12884 24296
rect 4928 24172 4968 24212
rect 5010 24172 5050 24212
rect 5092 24172 5132 24212
rect 5174 24172 5214 24212
rect 5256 24172 5296 24212
rect 5548 24004 5588 24044
rect 9964 24004 10004 24044
rect 12460 24004 12500 24044
rect 4012 23920 4052 23960
rect 10348 23920 10388 23960
rect 11500 23920 11540 23960
rect 4108 23836 4148 23876
rect 4972 23836 5012 23876
rect 7468 23836 7508 23876
rect 8332 23836 8372 23876
rect 5740 23752 5780 23792
rect 10252 23836 10292 23876
rect 11020 23867 11060 23876
rect 11020 23836 11060 23867
rect 11308 23836 11348 23876
rect 7756 23752 7796 23792
rect 8140 23752 8180 23792
rect 8524 23752 8564 23792
rect 10060 23752 10100 23792
rect 9100 23668 9140 23708
rect 4012 23584 4052 23624
rect 5740 23584 5780 23624
rect 7180 23584 7220 23624
rect 10828 23584 10868 23624
rect 12172 23584 12212 23624
rect 9388 23500 9428 23540
rect 3688 23416 3728 23456
rect 3770 23416 3810 23456
rect 3852 23416 3892 23456
rect 3934 23416 3974 23456
rect 4016 23416 4056 23456
rect 2668 23332 2708 23372
rect 13324 23416 13364 23456
rect 3916 23248 3956 23288
rect 13516 23332 13556 23372
rect 6220 23248 6260 23288
rect 10060 23248 10100 23288
rect 10348 23248 10388 23288
rect 4492 23164 4532 23204
rect 5644 23164 5684 23204
rect 8332 23164 8372 23204
rect 10444 23164 10484 23204
rect 10828 23164 10868 23204
rect 1804 23080 1844 23120
rect 4684 23080 4724 23120
rect 7756 23080 7796 23120
rect 8140 23080 8180 23120
rect 9004 23080 9044 23120
rect 9964 23080 10004 23120
rect 10540 23080 10580 23120
rect 2188 22996 2228 23036
rect 4108 22996 4148 23036
rect 4300 22996 4338 23036
rect 4338 22996 4340 23036
rect 5260 22996 5300 23036
rect 5740 22996 5748 23036
rect 5748 22996 5780 23036
rect 7372 22996 7412 23036
rect 8044 22996 8084 23036
rect 9196 22996 9204 23036
rect 9204 22996 9236 23036
rect 10060 22996 10100 23036
rect 11020 22996 11060 23036
rect 11212 22996 11252 23036
rect 5452 22912 5492 22952
rect 8620 22912 8660 22952
rect 11596 22912 11636 22952
rect 76 22828 116 22868
rect 5740 22828 5780 22868
rect 6892 22828 6932 22868
rect 76 22576 116 22616
rect 4928 22660 4968 22700
rect 5010 22660 5050 22700
rect 5092 22660 5132 22700
rect 5174 22660 5214 22700
rect 5256 22660 5296 22700
rect 9964 22576 10004 22616
rect 10444 22492 10484 22532
rect 11500 22492 11540 22532
rect 12076 22408 12116 22448
rect 4012 22324 4052 22364
rect 1228 22240 1268 22280
rect 4876 22324 4916 22364
rect 5644 22355 5684 22364
rect 5644 22324 5684 22355
rect 2860 22072 2900 22112
rect 3148 22072 3188 22112
rect 4588 22240 4628 22280
rect 5164 22240 5204 22280
rect 7180 22324 7220 22364
rect 8140 22324 8180 22364
rect 8620 22324 8660 22364
rect 8908 22355 8948 22364
rect 8908 22324 8948 22355
rect 11020 22355 11060 22364
rect 11020 22324 11060 22355
rect 11308 22324 11348 22364
rect 6892 22240 6932 22280
rect 7276 22240 7316 22280
rect 7756 22240 7796 22280
rect 8044 22240 8084 22280
rect 9196 22240 9236 22280
rect 9868 22240 9908 22280
rect 10156 22240 10196 22280
rect 10636 22240 10676 22280
rect 9292 22156 9332 22196
rect 8044 22072 8084 22112
rect 10444 22072 10484 22112
rect 9580 21988 9620 22028
rect 3688 21904 3728 21944
rect 3770 21904 3810 21944
rect 3852 21904 3892 21944
rect 3934 21904 3974 21944
rect 4016 21904 4056 21944
rect 11500 21904 11540 21944
rect 1612 21820 1652 21860
rect 4108 21736 4148 21776
rect 4876 21652 4916 21692
rect 7180 21652 7220 21692
rect 9100 21652 9140 21692
rect 11596 21652 11636 21692
rect 1228 21568 1268 21608
rect 2188 21568 2228 21608
rect 4108 21568 4148 21608
rect 5548 21568 5588 21608
rect 6412 21568 6452 21608
rect 9292 21568 9332 21608
rect 10540 21568 10580 21608
rect 4396 21484 4436 21524
rect 4972 21484 5012 21524
rect 2380 21400 2420 21440
rect 4108 20980 4148 21020
rect 6796 21484 6836 21524
rect 8716 21484 8756 21524
rect 9484 21484 9524 21524
rect 6412 21316 6452 21356
rect 4928 21148 4968 21188
rect 5010 21148 5050 21188
rect 5092 21148 5132 21188
rect 5174 21148 5214 21188
rect 5256 21148 5296 21188
rect 10636 21484 10676 21524
rect 11020 21484 11060 21524
rect 8908 21400 8948 21440
rect 9100 21400 9140 21440
rect 6892 21316 6932 21356
rect 10060 21316 10100 21356
rect 10828 21316 10868 21356
rect 11500 21316 11540 21356
rect 11980 21484 12020 21524
rect 12268 21484 12308 21524
rect 12556 21148 12596 21188
rect 6700 21064 6740 21104
rect 7948 21064 7988 21104
rect 9004 20980 9044 21020
rect 12172 20980 12212 21020
rect 11500 20896 11540 20936
rect 12844 20980 12884 21020
rect 2188 20812 2228 20852
rect 3244 20812 3284 20852
rect 4108 20812 4148 20852
rect 4492 20843 4532 20852
rect 4492 20812 4532 20843
rect 4972 20812 5012 20852
rect 5452 20812 5492 20852
rect 5644 20812 5684 20852
rect 6412 20812 6452 20852
rect 6700 20812 6740 20852
rect 8236 20812 8276 20852
rect 9004 20812 9044 20852
rect 9292 20812 9332 20852
rect 9580 20812 9611 20852
rect 9611 20812 9620 20852
rect 10060 20812 10100 20852
rect 10540 20812 10580 20852
rect 11308 20812 11348 20852
rect 76 20728 116 20768
rect 4588 20728 4628 20768
rect 11884 20728 11924 20768
rect 3148 20644 3188 20684
rect 10060 20644 10100 20684
rect 76 20560 116 20600
rect 1708 20560 1748 20600
rect 4396 20560 4436 20600
rect 8716 20560 8756 20600
rect 10156 20560 10196 20600
rect 12076 20560 12116 20600
rect 1996 20476 2036 20516
rect 10828 20476 10868 20516
rect 3148 20392 3188 20432
rect 3688 20392 3728 20432
rect 3770 20392 3810 20432
rect 3852 20392 3892 20432
rect 3934 20392 3974 20432
rect 4016 20392 4056 20432
rect 4972 20392 5012 20432
rect 11308 20392 11348 20432
rect 9580 20308 9620 20348
rect 10828 20308 10868 20348
rect 4108 20224 4148 20264
rect 9292 20224 9332 20264
rect 11596 20224 11636 20264
rect 3244 20140 3284 20180
rect 76 20056 116 20096
rect 5740 20056 5780 20096
rect 8908 20056 8948 20096
rect 10060 20056 10100 20096
rect 11500 20056 11540 20096
rect 13324 20056 13364 20096
rect 2476 19972 2516 20012
rect 3244 19972 3284 20012
rect 4588 19972 4628 20012
rect 9004 19972 9044 20012
rect 9292 19972 9332 20012
rect 10156 19972 10196 20012
rect 10828 19972 10868 20012
rect 2284 19804 2324 19844
rect 4396 19804 4436 19844
rect 4928 19636 4968 19676
rect 5010 19636 5050 19676
rect 5092 19636 5132 19676
rect 5174 19636 5214 19676
rect 5256 19636 5296 19676
rect 76 19552 116 19592
rect 3244 19468 3284 19508
rect 5644 19468 5684 19508
rect 10060 19888 10100 19928
rect 10156 19804 10196 19844
rect 10924 19804 10964 19844
rect 11884 19804 11924 19844
rect 12460 19888 12500 19928
rect 12172 19804 12212 19844
rect 12844 19552 12884 19592
rect 11596 19468 11636 19508
rect 4108 19384 4148 19424
rect 2572 19300 2612 19340
rect 4588 19300 4628 19340
rect 6124 19300 6164 19340
rect 7084 19300 7124 19340
rect 76 19216 116 19256
rect 4396 19216 4436 19256
rect 11212 19300 11252 19340
rect 10348 19216 10388 19256
rect 10540 19216 10580 19256
rect 4588 19132 4628 19172
rect 8524 19132 8564 19172
rect 9100 19132 9140 19172
rect 8044 19048 8084 19088
rect 10924 19048 10964 19088
rect 4588 18964 4628 19004
rect 9292 18964 9332 19004
rect 3688 18880 3728 18920
rect 3770 18880 3810 18920
rect 3852 18880 3892 18920
rect 3934 18880 3974 18920
rect 4016 18880 4056 18920
rect 12748 18880 12788 18920
rect 11692 18796 11732 18836
rect 3436 18628 3476 18668
rect 8332 18628 8372 18668
rect 76 18544 116 18584
rect 3148 18544 3188 18584
rect 10060 18544 10100 18584
rect 4108 18460 4148 18500
rect 4396 18460 4436 18500
rect 6892 18460 6932 18500
rect 7276 18460 7316 18500
rect 7756 18460 7796 18500
rect 8044 18460 8084 18500
rect 9484 18460 9524 18500
rect 4928 18124 4968 18164
rect 5010 18124 5050 18164
rect 5092 18124 5132 18164
rect 5174 18124 5214 18164
rect 5256 18124 5296 18164
rect 4684 18040 4724 18080
rect 2188 17956 2228 17996
rect 6124 17956 6164 17996
rect 7180 17956 7220 17996
rect 8524 17956 8564 17996
rect 5836 17872 5876 17912
rect 12172 18628 12212 18668
rect 12556 18628 12596 18668
rect 11884 18544 11924 18584
rect 10924 18460 10964 18500
rect 12076 18460 12116 18500
rect 9964 18376 10004 18416
rect 10348 18376 10388 18416
rect 10348 18208 10388 18248
rect 10636 18208 10676 18248
rect 10924 18208 10964 18248
rect 11500 18208 11540 18248
rect 12076 18208 12116 18248
rect 13132 18208 13172 18248
rect 2476 17788 2516 17828
rect 3724 17819 3764 17828
rect 3724 17788 3764 17819
rect 5740 17788 5780 17828
rect 6700 17788 6740 17828
rect 6988 17788 7028 17828
rect 76 17704 116 17744
rect 4300 17704 4340 17744
rect 4780 17704 4820 17744
rect 6124 17704 6164 17744
rect 4972 17620 5012 17660
rect 5260 17620 5300 17660
rect 76 17536 116 17576
rect 4204 17536 4244 17576
rect 5068 17536 5108 17576
rect 3688 17368 3728 17408
rect 3770 17368 3810 17408
rect 3852 17368 3892 17408
rect 3934 17368 3974 17408
rect 4016 17368 4056 17408
rect 9292 17788 9332 17828
rect 6508 17704 6548 17744
rect 6892 17704 6932 17744
rect 9964 17956 10004 17996
rect 10540 17956 10580 17996
rect 11596 17956 11636 17996
rect 12268 17872 12308 17912
rect 10924 17788 10964 17828
rect 11692 17788 11732 17828
rect 12076 17819 12116 17828
rect 12076 17788 12116 17819
rect 10348 17704 10388 17744
rect 10540 17704 10580 17744
rect 10828 17704 10868 17744
rect 11116 17704 11156 17744
rect 7084 17620 7124 17660
rect 8620 17620 8660 17660
rect 9964 17620 10004 17660
rect 13036 17620 13076 17660
rect 7468 17536 7508 17576
rect 12460 17536 12500 17576
rect 7276 17452 7316 17492
rect 11692 17452 11732 17492
rect 6028 17284 6068 17324
rect 6412 17284 6452 17324
rect 1900 17200 1940 17240
rect 3244 17200 3284 17240
rect 3340 17116 3380 17156
rect 3628 17200 3668 17240
rect 6220 17200 6260 17240
rect 7468 17200 7508 17240
rect 7756 17200 7796 17240
rect 12172 17200 12212 17240
rect 12844 17200 12884 17240
rect 13324 17200 13364 17240
rect 7276 17116 7316 17156
rect 7948 17116 7988 17156
rect 76 17032 116 17072
rect 3244 17032 3284 17072
rect 4876 17032 4916 17072
rect 5068 17032 5108 17072
rect 4300 16948 4340 16988
rect 5164 16948 5165 16988
rect 5165 16948 5204 16988
rect 6028 17032 6068 17072
rect 3340 16864 3380 16904
rect 3628 16864 3668 16904
rect 4588 16780 4628 16820
rect 4972 16780 5012 16820
rect 4928 16612 4968 16652
rect 5010 16612 5050 16652
rect 5092 16612 5132 16652
rect 5174 16612 5214 16652
rect 5256 16612 5296 16652
rect 6220 17032 6260 17072
rect 7660 17032 7700 17072
rect 7852 17032 7892 17072
rect 10060 17032 10100 17072
rect 10828 17032 10868 17072
rect 11500 17032 11540 17072
rect 7180 16948 7211 16988
rect 7211 16948 7220 16988
rect 7372 16948 7412 16988
rect 8620 16948 8660 16988
rect 9580 16948 9620 16988
rect 10444 16948 10484 16988
rect 10924 16948 10964 16988
rect 11884 16948 11924 16988
rect 6028 16864 6068 16904
rect 6316 16864 6356 16904
rect 6508 16864 6548 16904
rect 5452 16780 5492 16820
rect 6220 16780 6260 16820
rect 6316 16696 6356 16736
rect 6988 16780 7028 16820
rect 7372 16780 7412 16820
rect 6700 16696 6740 16736
rect 7756 16696 7796 16736
rect 10156 16864 10196 16904
rect 11788 16864 11828 16904
rect 12940 16864 12980 16904
rect 11692 16780 11732 16820
rect 5740 16612 5780 16652
rect 6508 16612 6548 16652
rect 76 16528 116 16568
rect 4780 16444 4820 16484
rect 4684 16360 4724 16400
rect 12556 16528 12596 16568
rect 6508 16444 6548 16484
rect 7852 16444 7892 16484
rect 8812 16444 8852 16484
rect 10540 16444 10580 16484
rect 11980 16444 12020 16484
rect 12748 16444 12788 16484
rect 4972 16360 5012 16400
rect 1900 16276 1940 16316
rect 4204 16276 4244 16316
rect 1228 16192 1268 16232
rect 6796 16360 6836 16400
rect 7180 16360 7220 16400
rect 7564 16360 7604 16400
rect 5740 16192 5780 16232
rect 7276 16276 7316 16316
rect 8332 16276 8372 16316
rect 6796 16108 6836 16148
rect 4204 16024 4244 16064
rect 5164 16024 5204 16064
rect 7084 16024 7124 16064
rect 5644 15940 5684 15980
rect 9100 16307 9140 16316
rect 9100 16276 9140 16307
rect 9964 16276 10004 16316
rect 10636 16276 10676 16316
rect 11212 16307 11252 16316
rect 11212 16276 11252 16307
rect 8140 16192 8180 16232
rect 10540 16192 10580 16232
rect 11596 16192 11636 16232
rect 12844 16192 12884 16232
rect 9868 16108 9908 16148
rect 8140 16024 8180 16064
rect 9580 15940 9620 15980
rect 11404 15940 11444 15980
rect 3688 15856 3728 15896
rect 3770 15856 3810 15896
rect 3852 15856 3892 15896
rect 3934 15856 3974 15896
rect 4016 15856 4056 15896
rect 9484 15856 9524 15896
rect 10060 15856 10100 15896
rect 4972 15772 5012 15812
rect 8524 15772 8564 15812
rect 9964 15772 10004 15812
rect 10252 15772 10292 15812
rect 1228 15520 1268 15560
rect 2476 15436 2516 15476
rect 5164 15688 5204 15728
rect 7084 15688 7124 15728
rect 7564 15688 7604 15728
rect 9100 15688 9140 15728
rect 6796 15604 6836 15644
rect 7276 15604 7316 15644
rect 8236 15604 8276 15644
rect 8620 15604 8660 15644
rect 5260 15436 5300 15476
rect 4204 15352 4244 15392
rect 5740 15352 5780 15392
rect 2476 15268 2516 15308
rect 4300 15268 4340 15308
rect 4928 15100 4968 15140
rect 5010 15100 5050 15140
rect 5092 15100 5132 15140
rect 5174 15100 5214 15140
rect 5256 15100 5296 15140
rect 7084 15436 7124 15476
rect 8428 15520 8459 15560
rect 8459 15520 8468 15560
rect 12076 15688 12116 15728
rect 8236 15436 8276 15476
rect 8524 15436 8564 15476
rect 9580 15436 9620 15476
rect 10540 15436 10580 15476
rect 10924 15436 10964 15476
rect 11212 15436 11252 15476
rect 2860 15016 2900 15056
rect 5452 14932 5492 14972
rect 3628 14848 3668 14888
rect 4012 14848 4052 14888
rect 4300 14848 4340 14888
rect 5356 14848 5396 14888
rect 7276 15100 7316 15140
rect 7948 15016 7988 15056
rect 7276 14932 7316 14972
rect 3724 14764 3764 14804
rect 4588 14764 4625 14804
rect 4625 14764 4628 14804
rect 4876 14764 4916 14804
rect 5164 14764 5195 14804
rect 5195 14764 5204 14804
rect 5548 14764 5588 14804
rect 5932 14764 5972 14804
rect 6316 14764 6356 14804
rect 4012 14680 4052 14720
rect 7564 14764 7604 14804
rect 7852 14764 7892 14804
rect 12172 15100 12212 15140
rect 13612 15016 13652 15056
rect 9484 14932 9524 14972
rect 10348 14848 10388 14888
rect 9580 14764 9620 14804
rect 10924 14764 10964 14804
rect 4684 14680 4724 14720
rect 5740 14680 5780 14720
rect 7084 14680 7124 14720
rect 7948 14680 7988 14720
rect 11692 14680 11732 14720
rect 12268 14680 12308 14720
rect 13132 14680 13172 14720
rect 2476 14596 2516 14636
rect 5836 14596 5876 14636
rect 5068 14512 5108 14552
rect 5836 14428 5876 14468
rect 7660 14596 7700 14636
rect 9100 14596 9140 14636
rect 9484 14596 9524 14636
rect 9772 14596 9812 14636
rect 8332 14512 8372 14552
rect 9676 14512 9716 14552
rect 10732 14512 10772 14552
rect 13132 14512 13172 14552
rect 9484 14428 9524 14468
rect 3688 14344 3728 14384
rect 3770 14344 3810 14384
rect 3852 14344 3892 14384
rect 3934 14344 3974 14384
rect 4016 14344 4056 14384
rect 7564 14344 7604 14384
rect 8236 14344 8276 14384
rect 8716 14344 8756 14384
rect 9100 14344 9140 14384
rect 9676 14344 9716 14384
rect 10252 14344 10292 14384
rect 11020 14344 11060 14384
rect 3148 14260 3188 14300
rect 7372 14260 7412 14300
rect 11116 14260 11156 14300
rect 4300 14176 4340 14216
rect 5068 14176 5108 14216
rect 8716 14176 8756 14216
rect 10540 14176 10580 14216
rect 11884 14176 11924 14216
rect 12748 14176 12788 14216
rect 4588 14092 4628 14132
rect 2380 14008 2420 14048
rect 5356 14008 5396 14048
rect 5836 14008 5876 14048
rect 3052 13924 3092 13964
rect 4204 13924 4244 13964
rect 5164 13840 5204 13880
rect 76 13756 116 13796
rect 5068 13756 5108 13796
rect 76 13504 116 13544
rect 4588 13504 4628 13544
rect 4928 13588 4968 13628
rect 5010 13588 5050 13628
rect 5092 13588 5132 13628
rect 5174 13588 5214 13628
rect 5256 13588 5296 13628
rect 7180 14008 7220 14048
rect 8332 14008 8372 14048
rect 8620 14008 8660 14048
rect 9676 14008 9716 14048
rect 10060 14008 10100 14048
rect 11596 14008 11636 14048
rect 7276 13924 7307 13964
rect 7307 13924 7316 13964
rect 10924 13924 10964 13964
rect 11404 13924 11444 13964
rect 8620 13840 8660 13880
rect 12460 14008 12500 14048
rect 6316 13756 6356 13796
rect 8524 13756 8564 13796
rect 8428 13672 8468 13712
rect 6412 13504 6452 13544
rect 9100 13504 9140 13544
rect 4684 13420 4715 13460
rect 4715 13420 4724 13460
rect 4876 13420 4916 13460
rect 9772 13420 9812 13460
rect 10156 13420 10196 13460
rect 4300 13336 4340 13376
rect 5836 13336 5876 13376
rect 6028 13336 6068 13376
rect 7948 13336 7988 13376
rect 10252 13336 10292 13376
rect 2956 13252 2996 13292
rect 4012 13252 4052 13292
rect 4684 13252 4724 13292
rect 4972 13252 5012 13292
rect 5260 13252 5300 13292
rect 6988 13252 7028 13292
rect 8140 13252 8180 13292
rect 8332 13252 8372 13292
rect 11596 13252 11636 13292
rect 1324 13168 1364 13208
rect 6412 13168 6452 13208
rect 6892 13168 6923 13208
rect 6923 13168 6932 13208
rect 6220 13084 6260 13124
rect 13324 13252 13364 13292
rect 8716 13168 8756 13208
rect 10348 13168 10388 13208
rect 7372 13084 7412 13124
rect 7948 13084 7988 13124
rect 12076 13084 12116 13124
rect 6892 13000 6932 13040
rect 8332 13000 8372 13040
rect 11404 13000 11444 13040
rect 6124 12916 6164 12956
rect 7084 12916 7124 12956
rect 3688 12832 3728 12872
rect 3770 12832 3810 12872
rect 3852 12832 3892 12872
rect 3934 12832 3974 12872
rect 4016 12832 4056 12872
rect 9772 12832 9812 12872
rect 12460 12832 12500 12872
rect 3820 12496 3860 12536
rect 7756 12748 7796 12788
rect 11692 12748 11732 12788
rect 4972 12496 5012 12536
rect 6700 12664 6740 12704
rect 8044 12664 8084 12704
rect 9580 12664 9620 12704
rect 11980 12664 12020 12704
rect 12172 12664 12212 12704
rect 6892 12580 6932 12620
rect 7180 12580 7220 12620
rect 8812 12580 8852 12620
rect 9196 12580 9236 12620
rect 9772 12580 9812 12620
rect 11500 12580 11540 12620
rect 12556 12580 12596 12620
rect 5836 12496 5876 12536
rect 6988 12496 7028 12536
rect 7468 12496 7508 12536
rect 10540 12496 10580 12536
rect 4108 12412 4148 12452
rect 4780 12412 4820 12452
rect 5740 12412 5780 12452
rect 6508 12412 6548 12452
rect 6796 12412 6836 12452
rect 8332 12412 8372 12452
rect 9196 12412 9236 12452
rect 4396 12328 4436 12368
rect 6316 12328 6356 12368
rect 6988 12328 7028 12368
rect 7180 12328 7220 12368
rect 4204 12244 4244 12284
rect 7276 12244 7316 12284
rect 3052 11908 3092 11948
rect 4012 11908 4052 11948
rect 12940 12496 12980 12536
rect 13324 12496 13364 12536
rect 10060 12412 10100 12452
rect 11404 12412 11444 12452
rect 9868 12328 9908 12368
rect 10156 12328 10196 12368
rect 8716 12244 8756 12284
rect 6412 12160 6452 12200
rect 8524 12160 8564 12200
rect 4928 12076 4968 12116
rect 5010 12076 5050 12116
rect 5092 12076 5132 12116
rect 5174 12076 5214 12116
rect 5256 12076 5296 12116
rect 6220 12076 6260 12116
rect 7180 12076 7220 12116
rect 11596 12244 11636 12284
rect 13036 12160 13076 12200
rect 9196 12076 9236 12116
rect 10156 11992 10196 12032
rect 8044 11908 8084 11948
rect 10252 11908 10292 11948
rect 11500 11908 11540 11948
rect 12364 11908 12404 11948
rect 6124 11824 6164 11864
rect 4300 11740 4340 11780
rect 5356 11740 5396 11780
rect 6316 11740 6356 11780
rect 6892 11771 6932 11780
rect 6892 11740 6932 11771
rect 7084 11740 7124 11780
rect 9292 11740 9323 11780
rect 9323 11740 9332 11780
rect 9772 11771 9812 11780
rect 9772 11740 9812 11771
rect 11500 11740 11540 11780
rect 12748 11740 12788 11780
rect 2092 11656 2132 11696
rect 2956 11656 2996 11696
rect 6124 11656 6164 11696
rect 6412 11656 6452 11696
rect 8620 11656 8660 11696
rect 10348 11656 10388 11696
rect 11308 11656 11348 11696
rect 12268 11656 12308 11696
rect 12844 11656 12884 11696
rect 13420 11656 13460 11696
rect 3340 11572 3380 11612
rect 8812 11572 8852 11612
rect 9100 11572 9140 11612
rect 11404 11572 11444 11612
rect 4300 11488 4340 11528
rect 10060 11488 10100 11528
rect 13420 11488 13460 11528
rect 8044 11404 8084 11444
rect 3688 11320 3728 11360
rect 3770 11320 3810 11360
rect 3852 11320 3892 11360
rect 3934 11320 3974 11360
rect 4016 11320 4056 11360
rect 6604 11320 6644 11360
rect 9100 11320 9140 11360
rect 10156 11320 10196 11360
rect 7852 11236 7892 11276
rect 11788 11236 11828 11276
rect 4108 11152 4148 11192
rect 4684 11152 4724 11192
rect 6316 11152 6356 11192
rect 7276 11152 7316 11192
rect 10540 11152 10580 11192
rect 11500 11152 11540 11192
rect 12268 11152 12308 11192
rect 1804 11068 1844 11108
rect 8332 11068 8372 11108
rect 10348 11068 10388 11108
rect 10732 11068 10772 11108
rect 1420 10984 1460 11024
rect 4684 10984 4724 11024
rect 6412 10984 6452 11024
rect 7564 10984 7604 11024
rect 7756 10984 7796 11024
rect 10252 10984 10292 11024
rect 12076 10984 12116 11024
rect 13132 10984 13172 11024
rect 2476 10900 2516 10940
rect 4300 10900 4340 10940
rect 5836 10900 5876 10940
rect 6124 10900 6164 10940
rect 6508 10900 6548 10940
rect 8428 10900 8468 10940
rect 9100 10900 9140 10940
rect 9772 10900 9780 10940
rect 9780 10900 9812 10940
rect 5740 10816 5780 10856
rect 6316 10816 6356 10856
rect 8044 10816 8084 10856
rect 8908 10816 8948 10856
rect 6892 10732 6932 10772
rect 13132 10816 13172 10856
rect 4928 10564 4968 10604
rect 5010 10564 5050 10604
rect 5092 10564 5132 10604
rect 5174 10564 5214 10604
rect 5256 10564 5296 10604
rect 4684 10396 4724 10436
rect 5452 10396 5492 10436
rect 6028 10396 6068 10436
rect 6220 10312 6260 10352
rect 2476 10228 2516 10268
rect 4684 10228 4724 10268
rect 5740 10228 5780 10268
rect 5932 10228 5972 10268
rect 6508 10228 6548 10268
rect 1996 10144 2036 10184
rect 4204 10144 4244 10184
rect 10636 10732 10676 10772
rect 7564 10564 7604 10604
rect 10348 10480 10388 10520
rect 11884 10480 11924 10520
rect 7756 10396 7796 10436
rect 9868 10396 9908 10436
rect 6988 10312 7028 10352
rect 9196 10312 9236 10352
rect 6700 10228 6740 10268
rect 8140 10228 8180 10268
rect 6028 10144 6068 10184
rect 8428 10228 8468 10268
rect 10252 10228 10292 10268
rect 11308 10228 11348 10268
rect 13324 10228 13364 10268
rect 12460 10144 12500 10184
rect 12844 10144 12884 10184
rect 5740 10060 5780 10100
rect 8428 10060 8468 10100
rect 76 9976 116 10016
rect 3688 9808 3728 9848
rect 3770 9808 3810 9848
rect 3852 9808 3892 9848
rect 3934 9808 3974 9848
rect 4016 9808 4056 9848
rect 11308 9808 11348 9848
rect 4396 9724 4436 9764
rect 5260 9724 5300 9764
rect 5548 9724 5588 9764
rect 11404 9724 11444 9764
rect 3436 9640 3476 9680
rect 5356 9640 5396 9680
rect 9388 9640 9428 9680
rect 9772 9640 9812 9680
rect 11788 9640 11828 9680
rect 4780 9556 4820 9596
rect 6412 9556 6452 9596
rect 6796 9556 6836 9596
rect 9100 9556 9140 9596
rect 9292 9556 9332 9596
rect 10444 9556 10484 9596
rect 13036 9556 13076 9596
rect 76 9472 116 9512
rect 2476 9472 2516 9512
rect 5548 9472 5588 9512
rect 7756 9472 7796 9512
rect 10252 9472 10292 9512
rect 11596 9472 11636 9512
rect 4588 9388 4628 9428
rect 4876 9388 4916 9428
rect 5356 9388 5396 9428
rect 6028 9388 6068 9428
rect 6988 9388 7028 9428
rect 7660 9388 7700 9428
rect 8332 9388 8372 9428
rect 9580 9388 9620 9428
rect 4928 9052 4968 9092
rect 5010 9052 5050 9092
rect 5092 9052 5132 9092
rect 5174 9052 5214 9092
rect 5256 9052 5296 9092
rect 12556 9388 12596 9428
rect 5548 9220 5588 9260
rect 5740 9136 5780 9176
rect 8332 9136 8372 9176
rect 11692 9136 11732 9176
rect 5740 8968 5780 9008
rect 7180 8968 7220 9008
rect 6124 8884 6164 8924
rect 8908 8884 8948 8924
rect 9100 8884 9140 8924
rect 5260 8800 5300 8840
rect 2476 8716 2516 8756
rect 4492 8716 4532 8756
rect 4780 8716 4820 8756
rect 5068 8716 5108 8756
rect 10540 8884 10580 8924
rect 11404 8884 11444 8924
rect 13516 8884 13556 8924
rect 6412 8800 6452 8840
rect 6796 8800 6836 8840
rect 8140 8800 8180 8840
rect 5452 8716 5492 8756
rect 1900 8632 1940 8672
rect 6220 8716 6260 8756
rect 7564 8716 7604 8756
rect 6604 8632 6644 8672
rect 6892 8632 6923 8672
rect 6923 8632 6932 8672
rect 6028 8548 6068 8588
rect 8908 8716 8948 8756
rect 9580 8716 9620 8756
rect 9292 8632 9332 8672
rect 11308 8632 11348 8672
rect 11884 8632 11924 8672
rect 12268 8632 12308 8672
rect 13420 8632 13460 8672
rect 5644 8464 5684 8504
rect 12172 8464 12212 8504
rect 3688 8296 3728 8336
rect 3770 8296 3810 8336
rect 3852 8296 3892 8336
rect 3934 8296 3974 8336
rect 4016 8296 4056 8336
rect 6988 8212 7028 8252
rect 4780 8128 4820 8168
rect 5836 8128 5876 8168
rect 8524 8128 8564 8168
rect 9388 8128 9428 8168
rect 12076 8128 12116 8168
rect 5356 8044 5396 8084
rect 7948 8044 7988 8084
rect 11980 8044 12020 8084
rect 12844 8044 12884 8084
rect 1420 7960 1460 8000
rect 8332 7960 8372 8000
rect 4684 7876 4724 7916
rect 5740 7876 5780 7916
rect 6124 7876 6164 7916
rect 6700 7876 6740 7916
rect 8140 7876 8180 7916
rect 11692 7960 11732 8000
rect 12268 7960 12308 8000
rect 13132 7960 13172 8000
rect 9004 7876 9044 7916
rect 10060 7876 10100 7916
rect 8332 7792 8372 7832
rect 9100 7792 9140 7832
rect 9484 7792 9524 7832
rect 7948 7708 7988 7748
rect 8140 7624 8180 7664
rect 4928 7540 4968 7580
rect 5010 7540 5050 7580
rect 5092 7540 5132 7580
rect 5174 7540 5214 7580
rect 5256 7540 5296 7580
rect 12460 7456 12500 7496
rect 5260 7372 5300 7412
rect 4780 7288 4820 7328
rect 6028 7288 6068 7328
rect 4876 7204 4916 7244
rect 5356 7204 5396 7244
rect 6796 7204 6836 7244
rect 1420 7120 1460 7160
rect 4972 7120 5012 7160
rect 8716 7204 8756 7244
rect 10828 7120 10868 7160
rect 11308 7120 11348 7160
rect 12076 7120 12116 7160
rect 12556 7120 12596 7160
rect 9004 7036 9044 7076
rect 556 6952 596 6992
rect 6124 6952 6164 6992
rect 7276 6868 7316 6908
rect 3688 6784 3728 6824
rect 3770 6784 3810 6824
rect 3852 6784 3892 6824
rect 3934 6784 3974 6824
rect 4016 6784 4056 6824
rect 4396 6784 4436 6824
rect 6220 6700 6260 6740
rect 5644 6616 5684 6656
rect 4876 6532 4916 6572
rect 9484 6532 9524 6572
rect 556 6448 596 6488
rect 5644 6448 5684 6488
rect 11692 6448 11732 6488
rect 12460 6448 12500 6488
rect 1516 6364 1556 6404
rect 3724 6364 3764 6404
rect 4684 6364 4724 6404
rect 6700 6364 6740 6404
rect 7564 6364 7604 6404
rect 8812 6364 8852 6404
rect 9292 6364 9332 6404
rect 11308 6364 11348 6404
rect 5740 6280 5780 6320
rect 7756 6280 7796 6320
rect 4780 6196 4820 6236
rect 7468 6196 7508 6236
rect 9580 6196 9620 6236
rect 5644 6112 5684 6152
rect 12460 6112 12500 6152
rect 4928 6028 4968 6068
rect 5010 6028 5050 6068
rect 5092 6028 5132 6068
rect 5174 6028 5214 6068
rect 5256 6028 5296 6068
rect 3724 5776 3764 5816
rect 4108 5776 4148 5816
rect 8812 5776 8852 5816
rect 11692 5776 11732 5816
rect 3148 5692 3188 5732
rect 6220 5692 6260 5732
rect 7948 5692 7988 5732
rect 8428 5692 8468 5732
rect 9100 5723 9140 5732
rect 9100 5692 9140 5723
rect 9580 5723 9620 5732
rect 9580 5692 9620 5723
rect 11788 5692 11828 5732
rect 4492 5608 4532 5648
rect 4684 5608 4724 5648
rect 5452 5608 5492 5648
rect 7756 5608 7796 5648
rect 10348 5608 10388 5648
rect 12460 5608 12500 5648
rect 5836 5524 5876 5564
rect 7084 5524 7124 5564
rect 7660 5524 7700 5564
rect 9676 5524 9716 5564
rect 1708 5440 1748 5480
rect 6316 5440 6356 5480
rect 8332 5440 8372 5480
rect 6220 5356 6260 5396
rect 6988 5356 7028 5396
rect 3688 5272 3728 5312
rect 3770 5272 3810 5312
rect 3852 5272 3892 5312
rect 3934 5272 3974 5312
rect 4016 5272 4056 5312
rect 9004 5188 9044 5228
rect 1228 4936 1268 4976
rect 4492 4936 4532 4976
rect 2956 4852 2996 4892
rect 4108 4852 4148 4892
rect 6700 5104 6740 5144
rect 9964 5104 10004 5144
rect 5836 5020 5876 5060
rect 7372 5020 7412 5060
rect 5356 4936 5396 4976
rect 5644 4936 5684 4976
rect 8140 4936 8180 4976
rect 9004 4936 9044 4976
rect 9484 4936 9524 4976
rect 9964 4936 10004 4976
rect 7468 4852 7508 4892
rect 7756 4852 7796 4892
rect 8236 4852 8276 4892
rect 9100 4852 9140 4892
rect 7372 4684 7412 4724
rect 8140 4600 8180 4640
rect 4928 4516 4968 4556
rect 5010 4516 5050 4556
rect 5092 4516 5132 4556
rect 5174 4516 5214 4556
rect 5256 4516 5296 4556
rect 8428 4516 8468 4556
rect 1228 4432 1268 4472
rect 7180 4432 7220 4472
rect 12460 4432 12500 4472
rect 3436 4264 3476 4304
rect 5932 4264 5972 4304
rect 7468 4264 7508 4304
rect 7852 4348 7892 4388
rect 8236 4264 8276 4304
rect 4108 4180 4148 4220
rect 4492 4180 4532 4220
rect 5644 4180 5684 4220
rect 8140 4180 8180 4220
rect 1612 4096 1652 4136
rect 3148 4096 3188 4136
rect 9004 4180 9044 4220
rect 7468 4096 7508 4136
rect 8236 4096 8276 4136
rect 12460 4096 12500 4136
rect 3244 4012 3284 4052
rect 8620 4012 8660 4052
rect 12652 4012 12692 4052
rect 76 3928 116 3968
rect 6988 3928 7028 3968
rect 9676 3928 9716 3968
rect 9964 3928 10004 3968
rect 6508 3844 6548 3884
rect 3688 3760 3728 3800
rect 3770 3760 3810 3800
rect 3852 3760 3892 3800
rect 3934 3760 3974 3800
rect 4016 3760 4056 3800
rect 4396 3760 4436 3800
rect 9772 3760 9812 3800
rect 7756 3676 7796 3716
rect 5548 3592 5588 3632
rect 7468 3592 7508 3632
rect 9100 3592 9140 3632
rect 10060 3592 10100 3632
rect 5356 3508 5396 3548
rect 5644 3508 5684 3548
rect 76 3424 116 3464
rect 9004 3508 9044 3548
rect 9196 3508 9236 3548
rect 9676 3424 9716 3464
rect 12652 3424 12692 3464
rect 2284 3340 2324 3380
rect 5452 3340 5492 3380
rect 7084 3340 7124 3380
rect 8620 3340 8660 3380
rect 1612 3172 1652 3212
rect 4928 3004 4968 3044
rect 5010 3004 5050 3044
rect 5092 3004 5132 3044
rect 5174 3004 5214 3044
rect 5256 3004 5296 3044
rect 8236 2836 8276 2876
rect 13516 2836 13556 2876
rect 13228 2752 13268 2792
rect 2572 2584 2612 2624
rect 5356 2584 5396 2624
rect 6988 2584 7028 2624
rect 7372 2584 7412 2624
rect 5740 2416 5780 2456
rect 3688 2248 3728 2288
rect 3770 2248 3810 2288
rect 3852 2248 3892 2288
rect 3934 2248 3974 2288
rect 4016 2248 4056 2288
rect 4780 2080 4820 2120
rect 76 1912 116 1952
rect 4928 1492 4968 1532
rect 5010 1492 5050 1532
rect 5092 1492 5132 1532
rect 5174 1492 5214 1532
rect 5256 1492 5296 1532
rect 76 1408 116 1448
rect 2188 1408 2228 1448
rect 4108 1408 4148 1448
<< metal3 >>
rect 1016 48304 1096 48384
rect 1592 48304 1672 48384
rect 2168 48304 2248 48384
rect 2744 48304 2824 48384
rect 3320 48304 3400 48384
rect 3896 48304 3976 48384
rect 4472 48304 4552 48384
rect 5048 48364 5128 48384
rect 5048 48324 5396 48364
rect 5048 48304 5156 48324
rect 652 46472 692 46481
rect 652 45800 692 46432
rect 1036 45968 1076 48304
rect 1036 45919 1076 45928
rect 1228 46808 1268 46817
rect 652 45751 692 45760
rect 1228 45800 1268 46768
rect 1612 46724 1652 48304
rect 1612 46675 1652 46684
rect 2188 46724 2228 48304
rect 2188 46675 2228 46684
rect 2764 46724 2804 48304
rect 2764 46675 2804 46684
rect 3340 46724 3380 48304
rect 3340 46675 3380 46684
rect 3916 46724 3956 48304
rect 3916 46675 3956 46684
rect 4492 46724 4532 48304
rect 5068 48280 5156 48304
rect 4928 46892 5296 46901
rect 4968 46852 5010 46892
rect 5050 46852 5092 46892
rect 5132 46852 5174 46892
rect 5214 46852 5256 46892
rect 4928 46843 5296 46852
rect 4492 46675 4532 46684
rect 5356 46724 5396 48324
rect 5624 48304 5704 48384
rect 6200 48304 6280 48384
rect 6776 48304 6856 48384
rect 7352 48304 7432 48384
rect 7928 48304 8008 48384
rect 8504 48304 8584 48384
rect 9080 48304 9160 48384
rect 9656 48304 9736 48384
rect 10232 48304 10312 48384
rect 10808 48304 10888 48384
rect 11384 48304 11464 48384
rect 11960 48304 12040 48384
rect 12536 48304 12616 48384
rect 5356 46675 5396 46684
rect 5644 46724 5684 48304
rect 5644 46675 5684 46684
rect 6220 46724 6260 48304
rect 6220 46675 6260 46684
rect 6796 46724 6836 48304
rect 6796 46675 6836 46684
rect 6892 46808 6932 46817
rect 1900 46472 1940 46481
rect 1900 46337 1940 46432
rect 2476 46472 2516 46481
rect 1228 45751 1268 45760
rect 1804 45800 1844 45809
rect 76 44960 116 44969
rect 76 44792 116 44920
rect 76 44743 116 44752
rect 76 44288 116 44297
rect 76 43784 116 44248
rect 76 43735 116 43744
rect 1228 43448 1268 43457
rect 1228 42776 1268 43408
rect 1228 42727 1268 42736
rect 76 41936 116 41945
rect 76 41768 116 41896
rect 76 41719 116 41728
rect 76 41264 116 41273
rect 76 40760 116 41224
rect 76 40711 116 40720
rect 1228 40424 1268 40433
rect 1228 39752 1268 40384
rect 1228 39703 1268 39712
rect 76 38912 116 38921
rect 76 38744 116 38872
rect 76 38695 116 38704
rect 76 38240 116 38249
rect 76 37736 116 38200
rect 76 37687 116 37696
rect 1516 37988 1556 37997
rect 1228 37400 1268 37409
rect 1228 36728 1268 37360
rect 1228 36679 1268 36688
rect 76 35888 116 35897
rect 76 35720 116 35848
rect 76 35671 116 35680
rect 76 35216 116 35225
rect 76 34712 116 35176
rect 76 34663 116 34672
rect 1228 34376 1268 34385
rect 1228 33704 1268 34336
rect 1228 33655 1268 33664
rect 76 32864 116 32873
rect 76 32696 116 32824
rect 76 32647 116 32656
rect 76 32192 116 32201
rect 76 31688 116 32152
rect 76 31639 116 31648
rect 1228 31352 1268 31361
rect 1228 30680 1268 31312
rect 1228 30631 1268 30640
rect 76 29840 116 29849
rect 76 29672 116 29800
rect 76 29623 116 29632
rect 1036 29756 1076 29765
rect 76 29168 116 29177
rect 76 28664 116 29128
rect 76 28615 116 28624
rect 76 22868 116 22877
rect 76 22616 116 22828
rect 76 22567 116 22576
rect 76 20768 116 20777
rect 76 20600 116 20728
rect 76 20551 116 20560
rect 76 20096 116 20105
rect 76 19592 116 20056
rect 76 19543 116 19552
rect 76 19256 116 19265
rect 76 18584 116 19216
rect 76 18535 116 18544
rect 76 17744 116 17753
rect 76 17576 116 17704
rect 76 17527 116 17536
rect 76 17072 116 17081
rect 76 16568 116 17032
rect 76 16519 116 16528
rect 76 13796 116 13805
rect 76 13544 116 13756
rect 76 13495 116 13504
rect 76 10016 116 10025
rect 76 9512 116 9976
rect 76 9463 116 9472
rect 556 6992 596 7001
rect 556 6488 596 6952
rect 556 6439 596 6448
rect 76 3968 116 3977
rect 76 3464 116 3928
rect 76 3415 116 3424
rect 76 1952 116 1961
rect 76 1448 116 1912
rect 76 1399 116 1408
rect 1036 80 1076 29716
rect 1228 28328 1268 28337
rect 1228 27656 1268 28288
rect 1228 27607 1268 27616
rect 1228 25976 1268 25985
rect 1268 25936 1364 25976
rect 1228 25927 1268 25936
rect 1228 22280 1268 22289
rect 1228 21608 1268 22240
rect 1228 21559 1268 21568
rect 1228 16232 1268 16241
rect 1228 15560 1268 16192
rect 1228 15511 1268 15520
rect 1324 13208 1364 25936
rect 1324 13159 1364 13168
rect 1420 11024 1460 11033
rect 1420 10889 1460 10984
rect 1420 8000 1460 8009
rect 1420 7865 1460 7960
rect 1420 7160 1460 7169
rect 1420 7025 1460 7120
rect 1516 6404 1556 37948
rect 1804 30344 1844 45760
rect 2284 41852 2324 41861
rect 2284 37460 2324 41812
rect 2284 37420 2420 37460
rect 1804 30295 1844 30304
rect 2188 36980 2228 36989
rect 1996 30176 2036 30185
rect 1996 29336 2036 30136
rect 1996 29287 2036 29296
rect 2188 27380 2228 36940
rect 2284 34964 2324 34973
rect 2284 28412 2324 34924
rect 2380 29084 2420 37420
rect 2476 35888 2516 46432
rect 5932 46472 5972 46481
rect 4204 46388 4244 46397
rect 3688 46136 4056 46145
rect 3728 46096 3770 46136
rect 3810 46096 3852 46136
rect 3892 46096 3934 46136
rect 3974 46096 4016 46136
rect 3688 46087 4056 46096
rect 3436 45548 3476 45557
rect 2668 44792 2708 44801
rect 2476 35839 2516 35848
rect 2572 41180 2612 41189
rect 2572 29336 2612 41140
rect 2668 37988 2708 44752
rect 2956 41012 2996 41021
rect 2668 37939 2708 37948
rect 2764 38912 2804 38921
rect 2668 35720 2708 35729
rect 2668 32108 2708 35680
rect 2668 30848 2708 32068
rect 2668 30799 2708 30808
rect 2572 29287 2612 29296
rect 2380 29044 2708 29084
rect 2668 28496 2708 29044
rect 2284 28363 2324 28372
rect 2476 28412 2516 28421
rect 2188 27340 2420 27380
rect 2284 25136 2324 25145
rect 2284 25001 2324 25096
rect 2092 24632 2132 24641
rect 1804 23120 1844 23129
rect 1612 21860 1652 21869
rect 1612 15980 1652 21820
rect 1612 15931 1652 15940
rect 1708 20600 1748 20609
rect 1516 6355 1556 6364
rect 1612 9008 1652 9017
rect 1228 4976 1268 4985
rect 1228 4472 1268 4936
rect 1228 4423 1268 4432
rect 1612 4136 1652 8968
rect 1708 5480 1748 20560
rect 1804 11108 1844 23080
rect 1996 20516 2036 20525
rect 1900 17240 1940 17249
rect 1900 16316 1940 17200
rect 1900 16267 1940 16276
rect 1996 16148 2036 20476
rect 1804 11059 1844 11068
rect 1900 16108 2036 16148
rect 1900 8672 1940 16108
rect 1996 15980 2036 15989
rect 1996 10184 2036 15940
rect 2092 11696 2132 24592
rect 2188 23036 2228 23045
rect 2188 21608 2228 22996
rect 2188 20852 2228 21568
rect 2284 22448 2324 22457
rect 2284 21272 2324 22408
rect 2380 21440 2420 27340
rect 2380 21391 2420 21400
rect 2476 26060 2516 28372
rect 2668 26900 2708 28456
rect 2668 26851 2708 26860
rect 2284 21232 2420 21272
rect 2188 17996 2228 20812
rect 2188 17947 2228 17956
rect 2284 19844 2324 19853
rect 2092 11647 2132 11656
rect 1996 10135 2036 10144
rect 1900 8623 1940 8632
rect 1708 5431 1748 5440
rect 1612 4087 1652 4096
rect 2284 3380 2324 19804
rect 2380 14048 2420 21232
rect 2476 20012 2516 26020
rect 2668 25976 2708 25985
rect 2668 25388 2708 25936
rect 2572 25136 2612 25145
rect 2572 22448 2612 25096
rect 2668 24548 2708 25348
rect 2668 23372 2708 24508
rect 2668 23323 2708 23332
rect 2572 22399 2612 22408
rect 2668 23036 2708 23045
rect 2476 17828 2516 19972
rect 2476 17779 2516 17788
rect 2572 22280 2612 22289
rect 2572 19340 2612 22240
rect 2668 20264 2708 22996
rect 2668 20215 2708 20224
rect 2572 15560 2612 19300
rect 2476 15520 2612 15560
rect 2668 15980 2708 15989
rect 2476 15476 2516 15520
rect 2476 15427 2516 15436
rect 2476 15308 2516 15317
rect 2476 14636 2516 15268
rect 2476 14587 2516 14596
rect 2572 15224 2612 15233
rect 2380 13999 2420 14008
rect 2476 12956 2516 12965
rect 2476 10940 2516 12916
rect 2476 10268 2516 10900
rect 2476 9512 2516 10228
rect 2476 8756 2516 9472
rect 2476 8707 2516 8716
rect 2284 3331 2324 3340
rect 1612 3212 1652 3221
rect 1612 80 1652 3172
rect 2572 2624 2612 15184
rect 2668 13040 2708 15940
rect 2668 12991 2708 13000
rect 2764 12956 2804 38872
rect 2860 32696 2900 32705
rect 2860 32612 2900 32656
rect 2860 32561 2900 32572
rect 2860 29504 2900 29513
rect 2860 29168 2900 29464
rect 2860 29119 2900 29128
rect 2956 26312 2996 40972
rect 3436 40340 3476 45508
rect 3688 44624 4056 44633
rect 3728 44584 3770 44624
rect 3810 44584 3852 44624
rect 3892 44584 3934 44624
rect 3974 44584 4016 44624
rect 3688 44575 4056 44584
rect 3688 43112 4056 43121
rect 3728 43072 3770 43112
rect 3810 43072 3852 43112
rect 3892 43072 3934 43112
rect 3974 43072 4016 43112
rect 3688 43063 4056 43072
rect 3688 41600 4056 41609
rect 3728 41560 3770 41600
rect 3810 41560 3852 41600
rect 3892 41560 3934 41600
rect 3974 41560 4016 41600
rect 3688 41551 4056 41560
rect 3436 40291 3476 40300
rect 3688 40088 4056 40097
rect 3728 40048 3770 40088
rect 3810 40048 3852 40088
rect 3892 40048 3934 40088
rect 3974 40048 4016 40088
rect 3688 40039 4056 40048
rect 4108 38912 4148 38921
rect 3688 38576 4056 38585
rect 3728 38536 3770 38576
rect 3810 38536 3852 38576
rect 3892 38536 3934 38576
rect 3974 38536 4016 38576
rect 3688 38527 4056 38536
rect 3820 38156 3860 38165
rect 3340 37484 3380 37493
rect 3148 37232 3188 37241
rect 3052 34208 3092 34217
rect 3052 29504 3092 34168
rect 3148 32948 3188 37192
rect 3340 36812 3380 37444
rect 3820 37484 3860 38116
rect 4108 38156 4148 38872
rect 4108 38107 4148 38116
rect 3820 37435 3860 37444
rect 4108 37568 4148 37577
rect 3688 37064 4056 37073
rect 3728 37024 3770 37064
rect 3810 37024 3852 37064
rect 3892 37024 3934 37064
rect 3974 37024 4016 37064
rect 3688 37015 4056 37024
rect 3148 32899 3188 32908
rect 3244 33620 3284 33629
rect 3148 32780 3188 32789
rect 3148 30680 3188 32740
rect 3244 31688 3284 33580
rect 3340 31772 3380 36772
rect 3688 35552 4056 35561
rect 3728 35512 3770 35552
rect 3810 35512 3852 35552
rect 3892 35512 3934 35552
rect 3974 35512 4016 35552
rect 3688 35503 4056 35512
rect 4108 35216 4148 37528
rect 4108 34544 4148 35176
rect 3688 34040 4056 34049
rect 3728 34000 3770 34040
rect 3810 34000 3852 34040
rect 3892 34000 3934 34040
rect 3974 34000 4016 34040
rect 3688 33991 4056 34000
rect 4108 33788 4148 34504
rect 4108 33739 4148 33748
rect 4108 33620 4148 33629
rect 3436 32948 3476 32957
rect 3436 31940 3476 32908
rect 3436 31891 3476 31900
rect 3532 32864 3572 32873
rect 3340 31732 3476 31772
rect 3244 31648 3380 31688
rect 3244 31436 3284 31445
rect 3244 30848 3284 31396
rect 3244 30799 3284 30808
rect 3244 30680 3284 30689
rect 3148 30640 3244 30680
rect 3052 29455 3092 29464
rect 3148 30512 3188 30521
rect 3148 29252 3188 30472
rect 3148 29203 3188 29212
rect 3148 29084 3188 29093
rect 2956 26272 3092 26312
rect 2956 25892 2996 25901
rect 2860 22112 2900 22121
rect 2860 21977 2900 22072
rect 2956 17576 2996 25852
rect 3052 23204 3092 26272
rect 3052 23155 3092 23164
rect 3148 24548 3188 29044
rect 3148 22280 3188 24508
rect 3148 22231 3188 22240
rect 3148 22112 3188 22121
rect 3148 20684 3188 22072
rect 3148 20432 3188 20644
rect 3148 20383 3188 20392
rect 3244 20852 3284 30640
rect 3148 20264 3188 20273
rect 2956 17527 2996 17536
rect 3052 20180 3092 20189
rect 2956 17408 2996 17417
rect 2860 15056 2900 15065
rect 2860 14921 2900 15016
rect 2956 13292 2996 17368
rect 3052 13964 3092 20140
rect 3148 18584 3188 20224
rect 3244 20180 3284 20812
rect 3244 20131 3284 20140
rect 3244 20012 3284 20021
rect 3244 19508 3284 19972
rect 3244 19459 3284 19468
rect 3188 18544 3284 18584
rect 3148 18535 3188 18544
rect 3148 17576 3188 17585
rect 3148 15056 3188 17536
rect 3244 17240 3284 18544
rect 3244 17191 3284 17200
rect 3340 17156 3380 31648
rect 3436 28580 3476 31732
rect 3436 28531 3476 28540
rect 3436 26900 3476 26909
rect 3436 25556 3476 26860
rect 3436 25507 3476 25516
rect 3532 23204 3572 32824
rect 4108 32864 4148 33580
rect 4108 32815 4148 32824
rect 3688 32528 4056 32537
rect 3728 32488 3770 32528
rect 3810 32488 3852 32528
rect 3892 32488 3934 32528
rect 3974 32488 4016 32528
rect 3688 32479 4056 32488
rect 3724 32360 3764 32369
rect 3724 32024 3764 32320
rect 3724 31975 3764 31984
rect 4108 32192 4148 32201
rect 4012 31940 4052 31949
rect 4012 31805 4052 31900
rect 4108 31436 4148 32152
rect 3688 31016 4056 31025
rect 3728 30976 3770 31016
rect 3810 30976 3852 31016
rect 3892 30976 3934 31016
rect 3974 30976 4016 31016
rect 3688 30967 4056 30976
rect 3820 30848 3860 30857
rect 3724 30764 3764 30773
rect 3724 29672 3764 30724
rect 3820 29756 3860 30808
rect 4108 30848 4148 31396
rect 4108 30799 4148 30808
rect 3820 29707 3860 29716
rect 4012 30764 4052 30773
rect 4012 30596 4052 30724
rect 4012 29756 4052 30556
rect 4108 30512 4148 30521
rect 4108 30428 4148 30472
rect 4108 30377 4148 30388
rect 4204 30260 4244 46348
rect 4684 46304 4724 46313
rect 4588 43280 4628 43289
rect 4588 40340 4628 43240
rect 4588 40291 4628 40300
rect 4396 38912 4436 38921
rect 4396 38072 4436 38872
rect 4684 38324 4724 46264
rect 4928 45380 5296 45389
rect 4968 45340 5010 45380
rect 5050 45340 5092 45380
rect 5132 45340 5174 45380
rect 5214 45340 5256 45380
rect 4928 45331 5296 45340
rect 5932 45212 5972 46432
rect 5932 45163 5972 45172
rect 6508 46472 6548 46481
rect 6508 45128 6548 46432
rect 6508 45079 6548 45088
rect 6700 46136 6740 46145
rect 5452 44960 5492 44969
rect 5452 44825 5492 44920
rect 5548 44876 5588 44885
rect 5356 44204 5396 44213
rect 4928 43868 5296 43877
rect 4968 43828 5010 43868
rect 5050 43828 5092 43868
rect 5132 43828 5174 43868
rect 5214 43828 5256 43868
rect 4928 43819 5296 43828
rect 4928 42356 5296 42365
rect 4968 42316 5010 42356
rect 5050 42316 5092 42356
rect 5132 42316 5174 42356
rect 5214 42316 5256 42356
rect 4928 42307 5296 42316
rect 4928 40844 5296 40853
rect 4968 40804 5010 40844
rect 5050 40804 5092 40844
rect 5132 40804 5174 40844
rect 5214 40804 5256 40844
rect 4928 40795 5296 40804
rect 4928 39332 5296 39341
rect 4968 39292 5010 39332
rect 5050 39292 5092 39332
rect 5132 39292 5174 39332
rect 5214 39292 5256 39332
rect 4928 39283 5296 39292
rect 4684 38275 4724 38284
rect 4300 38032 4436 38072
rect 4300 36560 4340 38032
rect 4492 37988 4532 37997
rect 4300 36392 4340 36520
rect 4300 32276 4340 36352
rect 4300 32227 4340 32236
rect 4396 37484 4436 37493
rect 4396 36644 4436 37444
rect 4396 35804 4436 36604
rect 4396 35216 4436 35764
rect 4396 32192 4436 35176
rect 4396 32143 4436 32152
rect 4300 32108 4340 32117
rect 4300 31604 4340 32068
rect 4300 31555 4340 31564
rect 4396 32024 4436 32033
rect 4108 30220 4244 30260
rect 4300 30848 4340 30857
rect 4300 30260 4340 30808
rect 4108 30008 4148 30220
rect 4300 30211 4340 30220
rect 4396 30176 4436 31984
rect 4492 30260 4532 37948
rect 5356 37988 5396 44164
rect 5356 37939 5396 37948
rect 5452 38324 5492 38333
rect 4928 37820 5296 37829
rect 4968 37780 5010 37820
rect 5050 37780 5092 37820
rect 5132 37780 5174 37820
rect 5214 37780 5256 37820
rect 4928 37771 5296 37780
rect 4588 36476 4628 36485
rect 4588 31520 4628 36436
rect 4928 36308 5296 36317
rect 4968 36268 5010 36308
rect 5050 36268 5092 36308
rect 5132 36268 5174 36308
rect 5214 36268 5256 36308
rect 4928 36259 5296 36268
rect 4588 31471 4628 31480
rect 4684 35888 4724 35897
rect 4684 35132 4724 35848
rect 4684 34460 4724 35092
rect 4928 34796 5296 34805
rect 4968 34756 5010 34796
rect 5050 34756 5092 34796
rect 5132 34756 5174 34796
rect 5214 34756 5256 34796
rect 4928 34747 5296 34756
rect 4492 30211 4532 30220
rect 4588 31352 4628 31361
rect 4588 30428 4628 31312
rect 4396 30127 4436 30136
rect 4588 30176 4628 30388
rect 4684 30260 4724 34420
rect 4928 33284 5296 33293
rect 4968 33244 5010 33284
rect 5050 33244 5092 33284
rect 5132 33244 5174 33284
rect 5214 33244 5256 33284
rect 4928 33235 5296 33244
rect 5452 33140 5492 38284
rect 5260 33100 5492 33140
rect 4684 30211 4724 30220
rect 4780 32864 4820 32873
rect 4780 32192 4820 32824
rect 4780 30260 4820 32152
rect 4876 32780 4916 32789
rect 4876 32024 4916 32740
rect 4876 31975 4916 31984
rect 5164 31940 5204 32035
rect 5260 31940 5300 33100
rect 5452 32948 5492 32957
rect 5356 32864 5396 32873
rect 5356 32108 5396 32824
rect 5452 32276 5492 32908
rect 5452 32227 5492 32236
rect 5396 32068 5492 32108
rect 5356 32059 5396 32068
rect 5260 31900 5396 31940
rect 5164 31891 5204 31900
rect 4928 31772 5296 31781
rect 4968 31732 5010 31772
rect 5050 31732 5092 31772
rect 5132 31732 5174 31772
rect 5214 31732 5256 31772
rect 4928 31723 5296 31732
rect 4876 31436 4916 31445
rect 4876 30764 4916 31396
rect 5260 31436 5300 31445
rect 4876 30512 4916 30724
rect 5068 31268 5108 31277
rect 5068 30596 5108 31228
rect 5260 31184 5300 31396
rect 5260 31135 5300 31144
rect 5068 30547 5108 30556
rect 4876 30463 4916 30472
rect 4780 30211 4820 30220
rect 4928 30260 5296 30269
rect 4968 30220 5010 30260
rect 5050 30220 5092 30260
rect 5132 30220 5174 30260
rect 5214 30220 5256 30260
rect 4928 30211 5296 30220
rect 4588 30127 4628 30136
rect 4876 30092 4916 30101
rect 4780 30008 4820 30017
rect 4108 29968 4244 30008
rect 4012 29707 4052 29716
rect 4108 29840 4148 29849
rect 3724 29623 3764 29632
rect 3688 29504 4056 29513
rect 3728 29464 3770 29504
rect 3810 29464 3852 29504
rect 3892 29464 3934 29504
rect 3974 29464 4016 29504
rect 3688 29455 4056 29464
rect 4108 28580 4148 29800
rect 4108 28531 4148 28540
rect 3688 27992 4056 28001
rect 3728 27952 3770 27992
rect 3810 27952 3852 27992
rect 3892 27952 3934 27992
rect 3974 27952 4016 27992
rect 3688 27943 4056 27952
rect 3688 26480 4056 26489
rect 3728 26440 3770 26480
rect 3810 26440 3852 26480
rect 3892 26440 3934 26480
rect 3974 26440 4016 26480
rect 3688 26431 4056 26440
rect 4108 26060 4148 26069
rect 4108 25925 4148 26020
rect 4012 25556 4052 25565
rect 4012 25136 4052 25516
rect 4108 25388 4148 25397
rect 4108 25253 4148 25348
rect 4012 25096 4148 25136
rect 3688 24968 4056 24977
rect 3728 24928 3770 24968
rect 3810 24928 3852 24968
rect 3892 24928 3934 24968
rect 3974 24928 4016 24968
rect 3688 24919 4056 24928
rect 4108 24800 4148 25096
rect 4012 24760 4148 24800
rect 4012 23960 4052 24760
rect 4012 23624 4052 23920
rect 4012 23575 4052 23584
rect 4108 24632 4148 24641
rect 4108 23876 4148 24592
rect 3688 23456 4056 23465
rect 3728 23416 3770 23456
rect 3810 23416 3852 23456
rect 3892 23416 3934 23456
rect 3974 23416 4016 23456
rect 3688 23407 4056 23416
rect 3916 23288 3956 23297
rect 4108 23288 4148 23836
rect 3532 23164 3668 23204
rect 3436 23036 3476 23045
rect 3436 18668 3476 22996
rect 3628 22952 3668 23164
rect 3436 18619 3476 18628
rect 3532 22912 3668 22952
rect 3340 17107 3380 17116
rect 3148 15007 3188 15016
rect 3244 17072 3284 17081
rect 3148 14888 3188 14897
rect 3148 14300 3188 14848
rect 3148 14251 3188 14260
rect 3092 13924 3188 13964
rect 3052 13915 3092 13924
rect 2764 12907 2804 12916
rect 2860 13040 2900 13049
rect 2860 12704 2900 13000
rect 2764 12664 2900 12704
rect 2764 9848 2804 12664
rect 2764 9799 2804 9808
rect 2956 11696 2996 13252
rect 3052 13796 3092 13805
rect 3052 11948 3092 13756
rect 3052 11899 3092 11908
rect 2956 4892 2996 11656
rect 2956 4843 2996 4852
rect 3052 9848 3092 9857
rect 3052 2900 3092 9808
rect 3148 5732 3188 13924
rect 3244 13796 3284 17032
rect 3244 13747 3284 13756
rect 3340 16904 3380 16913
rect 3340 13628 3380 16864
rect 3148 4136 3188 5692
rect 3148 4087 3188 4096
rect 3244 13588 3380 13628
rect 3436 15140 3476 15149
rect 3244 4052 3284 13588
rect 3244 4003 3284 4012
rect 3340 11612 3380 11621
rect 3052 2860 3284 2900
rect 2572 2575 2612 2584
rect 2188 1448 2228 1457
rect 2188 80 2228 1408
rect 2764 1448 2804 1457
rect 2764 80 2804 1408
rect 3244 188 3284 2860
rect 3244 139 3284 148
rect 3340 80 3380 11572
rect 3436 9680 3476 15100
rect 3436 9631 3476 9640
rect 3436 4304 3476 4313
rect 3436 4169 3476 4264
rect 3532 2900 3572 22912
rect 3916 22112 3956 23248
rect 4012 23248 4148 23288
rect 4012 22364 4052 23248
rect 4012 22315 4052 22324
rect 4108 23036 4148 23045
rect 3916 22063 3956 22072
rect 3688 21944 4056 21953
rect 3728 21904 3770 21944
rect 3810 21904 3852 21944
rect 3892 21904 3934 21944
rect 3974 21904 4016 21944
rect 3688 21895 4056 21904
rect 4108 21776 4148 22996
rect 4108 21727 4148 21736
rect 4108 21608 4148 21617
rect 4108 21020 4148 21568
rect 4108 20971 4148 20980
rect 4108 20852 4148 20861
rect 3688 20432 4056 20441
rect 3728 20392 3770 20432
rect 3810 20392 3852 20432
rect 3892 20392 3934 20432
rect 3974 20392 4016 20432
rect 3688 20383 4056 20392
rect 3628 20264 3668 20273
rect 3628 19088 3668 20224
rect 4108 20264 4148 20812
rect 4108 20215 4148 20224
rect 3628 19039 3668 19048
rect 4108 19424 4148 19433
rect 3688 18920 4056 18929
rect 3728 18880 3770 18920
rect 3810 18880 3852 18920
rect 3892 18880 3934 18920
rect 3974 18880 4016 18920
rect 3688 18871 4056 18880
rect 4108 18500 4148 19384
rect 4108 18451 4148 18460
rect 3724 18080 3764 18089
rect 3724 17828 3764 18040
rect 4204 17996 4244 29968
rect 4492 29840 4532 29849
rect 4396 29084 4436 29093
rect 4396 28412 4436 29044
rect 4396 28363 4436 28372
rect 4300 26816 4340 26825
rect 4300 23036 4340 26776
rect 4492 23204 4532 29800
rect 4588 27572 4628 27581
rect 4588 26228 4628 27532
rect 4588 26179 4628 26188
rect 4684 26900 4724 26909
rect 4684 26060 4724 26860
rect 4492 23155 4532 23164
rect 4588 26020 4724 26060
rect 4300 22901 4340 22996
rect 4396 22784 4436 22793
rect 3724 17779 3764 17788
rect 4108 17956 4244 17996
rect 4300 22112 4340 22121
rect 3688 17408 4056 17417
rect 3728 17368 3770 17408
rect 3810 17368 3852 17408
rect 3892 17368 3934 17408
rect 3974 17368 4016 17408
rect 3688 17359 4056 17368
rect 3628 17240 3668 17249
rect 3628 16904 3668 17200
rect 3628 16855 3668 16864
rect 3688 15896 4056 15905
rect 3728 15856 3770 15896
rect 3810 15856 3852 15896
rect 3892 15856 3934 15896
rect 3974 15856 4016 15896
rect 3688 15847 4056 15856
rect 4012 15728 4052 15737
rect 3628 14888 3668 14897
rect 3628 14753 3668 14848
rect 4012 14888 4052 15688
rect 4012 14839 4052 14848
rect 3724 14804 3764 14813
rect 3724 14636 3764 14764
rect 3724 14587 3764 14596
rect 4012 14720 4052 14729
rect 4012 14585 4052 14680
rect 3688 14384 4056 14393
rect 3728 14344 3770 14384
rect 3810 14344 3852 14384
rect 3892 14344 3934 14384
rect 3974 14344 4016 14384
rect 3688 14335 4056 14344
rect 4012 13292 4052 13301
rect 4012 13157 4052 13252
rect 3688 12872 4056 12881
rect 3728 12832 3770 12872
rect 3810 12832 3852 12872
rect 3892 12832 3934 12872
rect 3974 12832 4016 12872
rect 3688 12823 4056 12832
rect 4108 12620 4148 17956
rect 4300 17744 4340 22072
rect 4396 21524 4436 22744
rect 4588 22532 4628 26020
rect 4588 22483 4628 22492
rect 4684 23120 4724 23129
rect 4396 20600 4436 21484
rect 4588 22280 4628 22289
rect 4684 22280 4724 23080
rect 4628 22240 4724 22280
rect 4492 20852 4532 20861
rect 4492 20717 4532 20812
rect 4588 20768 4628 22240
rect 4396 20551 4436 20560
rect 4588 20180 4628 20728
rect 4492 20140 4628 20180
rect 4684 20180 4724 20189
rect 4204 17576 4244 17585
rect 4204 17324 4244 17536
rect 4204 16484 4244 17284
rect 4300 16988 4340 17704
rect 4300 16939 4340 16948
rect 4396 19844 4436 19853
rect 4396 19256 4436 19804
rect 4396 18500 4436 19216
rect 4204 16444 4340 16484
rect 4012 12580 4148 12620
rect 4204 16316 4244 16325
rect 4204 16064 4244 16276
rect 4204 15392 4244 16024
rect 4204 13964 4244 15352
rect 4300 15308 4340 16444
rect 4300 14888 4340 15268
rect 4396 15056 4436 18460
rect 4396 15007 4436 15016
rect 4340 14848 4436 14888
rect 4300 14839 4340 14848
rect 4300 14720 4340 14729
rect 4300 14216 4340 14680
rect 4396 14552 4436 14848
rect 4492 14804 4532 20140
rect 4588 20012 4628 20021
rect 4588 19340 4628 19972
rect 4588 19172 4628 19300
rect 4588 19123 4628 19132
rect 4588 19004 4628 19013
rect 4588 16988 4628 18964
rect 4684 18080 4724 20140
rect 4684 18031 4724 18040
rect 4780 17912 4820 29968
rect 4876 28916 4916 30052
rect 5260 30092 5300 30101
rect 4972 29924 5012 29933
rect 4972 29504 5012 29884
rect 4972 29455 5012 29464
rect 5260 29000 5300 30052
rect 5356 30008 5396 31900
rect 5356 29959 5396 29968
rect 5356 29672 5396 29681
rect 5356 29168 5396 29632
rect 5356 29119 5396 29128
rect 5260 28960 5396 29000
rect 4876 28867 4916 28876
rect 4928 28748 5296 28757
rect 4968 28708 5010 28748
rect 5050 28708 5092 28748
rect 5132 28708 5174 28748
rect 5214 28708 5256 28748
rect 4928 28699 5296 28708
rect 4928 27236 5296 27245
rect 4968 27196 5010 27236
rect 5050 27196 5092 27236
rect 5132 27196 5174 27236
rect 5214 27196 5256 27236
rect 4928 27187 5296 27196
rect 5356 27068 5396 28960
rect 5260 27028 5396 27068
rect 4972 26816 5012 26825
rect 4972 26681 5012 26776
rect 5260 26480 5300 27028
rect 5260 26431 5300 26440
rect 4928 25724 5296 25733
rect 4968 25684 5010 25724
rect 5050 25684 5092 25724
rect 5132 25684 5174 25724
rect 5214 25684 5256 25724
rect 4928 25675 5296 25684
rect 5452 25220 5492 32068
rect 5548 30260 5588 44836
rect 6124 44036 6164 44045
rect 5836 41936 5876 41945
rect 5740 40340 5780 40349
rect 5740 39080 5780 40300
rect 5740 39031 5780 39040
rect 5740 37232 5780 37241
rect 5548 30211 5588 30220
rect 5644 32864 5684 32873
rect 5644 32696 5684 32824
rect 5644 30092 5684 32656
rect 5740 31436 5780 37192
rect 5740 31387 5780 31396
rect 5740 30512 5780 30521
rect 5740 30344 5780 30472
rect 5740 30295 5780 30304
rect 5548 30052 5684 30092
rect 5548 27572 5588 30052
rect 5740 30008 5780 30017
rect 5644 29924 5684 29933
rect 5644 29336 5684 29884
rect 5644 29287 5684 29296
rect 5740 29168 5780 29968
rect 5548 27068 5588 27532
rect 5548 27019 5588 27028
rect 5644 29128 5740 29168
rect 5452 25171 5492 25180
rect 5548 26900 5588 26909
rect 4928 24212 5296 24221
rect 4968 24172 5010 24212
rect 5050 24172 5092 24212
rect 5132 24172 5174 24212
rect 5214 24172 5256 24212
rect 4928 24163 5296 24172
rect 5548 24044 5588 26860
rect 5644 26060 5684 29128
rect 5740 29119 5780 29128
rect 5740 28076 5780 28085
rect 5740 26648 5780 28036
rect 5836 26732 5876 41896
rect 6124 39668 6164 43996
rect 6508 43280 6548 43289
rect 6124 39619 6164 39628
rect 6220 40424 6260 40433
rect 6220 38240 6260 40384
rect 6316 38996 6356 39005
rect 6316 38408 6356 38956
rect 6316 38359 6356 38368
rect 6220 38200 6356 38240
rect 6028 37484 6068 37493
rect 6028 36644 6068 37444
rect 6028 35972 6068 36604
rect 5932 35048 5972 35057
rect 5932 28076 5972 35008
rect 6028 33368 6068 35932
rect 6220 36476 6260 36485
rect 6220 35132 6260 36436
rect 6220 35083 6260 35092
rect 6028 33319 6068 33328
rect 6124 34964 6164 34973
rect 5932 28027 5972 28036
rect 6028 33200 6068 33209
rect 5932 27404 5972 27413
rect 5932 26900 5972 27364
rect 5932 26851 5972 26860
rect 5836 26692 5972 26732
rect 5740 26608 5876 26648
rect 5644 25388 5684 26020
rect 5644 25339 5684 25348
rect 5740 26480 5780 26489
rect 4972 23876 5012 23885
rect 4972 22868 5012 23836
rect 5548 23120 5588 24004
rect 5740 23792 5780 26440
rect 5740 23743 5780 23752
rect 5740 23624 5780 23633
rect 5548 23071 5588 23080
rect 5644 23204 5684 23213
rect 5260 23036 5300 23045
rect 5260 22901 5300 22996
rect 5452 22952 5492 22961
rect 4972 22819 5012 22828
rect 4928 22700 5296 22709
rect 4968 22660 5010 22700
rect 5050 22660 5092 22700
rect 5132 22660 5174 22700
rect 5214 22660 5256 22700
rect 4928 22651 5296 22660
rect 5164 22532 5204 22541
rect 4876 22364 4916 22373
rect 4876 21692 4916 22324
rect 4876 21643 4916 21652
rect 5164 22280 5204 22492
rect 4972 21524 5012 21533
rect 4972 21389 5012 21484
rect 5164 21356 5204 22240
rect 5164 21307 5204 21316
rect 5356 21524 5396 21533
rect 4928 21188 5296 21197
rect 4968 21148 5010 21188
rect 5050 21148 5092 21188
rect 5132 21148 5174 21188
rect 5214 21148 5256 21188
rect 4928 21139 5296 21148
rect 4972 21020 5012 21029
rect 4972 20852 5012 20980
rect 5260 21020 5300 21029
rect 4972 20432 5012 20812
rect 4972 20383 5012 20392
rect 5068 20936 5108 20945
rect 5068 19844 5108 20896
rect 5260 20180 5300 20980
rect 5356 20936 5396 21484
rect 5452 21020 5492 22912
rect 5644 22364 5684 23164
rect 5740 23036 5780 23584
rect 5740 22987 5780 22996
rect 5452 20971 5492 20980
rect 5548 21608 5588 21617
rect 5356 20887 5396 20896
rect 5452 20852 5492 20861
rect 5260 20140 5396 20180
rect 5068 19795 5108 19804
rect 4928 19676 5296 19685
rect 4968 19636 5010 19676
rect 5050 19636 5092 19676
rect 5132 19636 5174 19676
rect 5214 19636 5256 19676
rect 4928 19627 5296 19636
rect 4928 18164 5296 18173
rect 4968 18124 5010 18164
rect 5050 18124 5092 18164
rect 5132 18124 5174 18164
rect 5214 18124 5256 18164
rect 4928 18115 5296 18124
rect 4588 16939 4628 16948
rect 4684 17872 4820 17912
rect 4876 17996 4916 18005
rect 5356 17996 5396 20140
rect 4588 16820 4628 16829
rect 4588 15728 4628 16780
rect 4684 16400 4724 17872
rect 4684 16351 4724 16360
rect 4780 17744 4820 17753
rect 4780 16484 4820 17704
rect 4876 17072 4916 17956
rect 5164 17956 5396 17996
rect 4972 17660 5012 17669
rect 4972 17492 5012 17620
rect 4972 17443 5012 17452
rect 5068 17576 5108 17585
rect 4876 17023 4916 17032
rect 5068 17072 5108 17536
rect 5068 17023 5108 17032
rect 5164 17240 5204 17956
rect 5260 17660 5300 17669
rect 5260 17525 5300 17620
rect 5452 17300 5492 20812
rect 5164 16988 5204 17200
rect 5164 16939 5204 16948
rect 5356 17260 5492 17300
rect 4972 16820 5012 16915
rect 4972 16771 5012 16780
rect 4928 16652 5296 16661
rect 4968 16612 5010 16652
rect 5050 16612 5092 16652
rect 5132 16612 5174 16652
rect 5214 16612 5256 16652
rect 4928 16603 5296 16612
rect 4588 15679 4628 15688
rect 4492 14755 4532 14764
rect 4588 14804 4628 14813
rect 4780 14804 4820 16444
rect 4972 16400 5012 16409
rect 4972 15812 5012 16360
rect 5260 16232 5300 16241
rect 4972 15763 5012 15772
rect 5164 16064 5204 16073
rect 5164 15728 5204 16024
rect 5164 15679 5204 15688
rect 5260 15476 5300 16192
rect 5260 15427 5300 15436
rect 4928 15140 5296 15149
rect 4968 15100 5010 15140
rect 5050 15100 5092 15140
rect 5132 15100 5174 15140
rect 5214 15100 5256 15140
rect 4928 15091 5296 15100
rect 5260 14972 5300 14981
rect 4876 14804 4916 14813
rect 4780 14764 4876 14804
rect 4396 14512 4532 14552
rect 4300 14167 4340 14176
rect 4396 14384 4436 14393
rect 3820 12536 3860 12545
rect 3820 12401 3860 12496
rect 4012 11948 4052 12580
rect 4012 11899 4052 11908
rect 4108 12452 4148 12461
rect 3688 11360 4056 11369
rect 3728 11320 3770 11360
rect 3810 11320 3852 11360
rect 3892 11320 3934 11360
rect 3974 11320 4016 11360
rect 3688 11311 4056 11320
rect 4108 11192 4148 12412
rect 4108 11143 4148 11152
rect 4204 12284 4244 13924
rect 4300 14048 4340 14057
rect 4300 13376 4340 14008
rect 4300 13327 4340 13336
rect 4204 10184 4244 12244
rect 4300 13124 4340 13133
rect 4300 11780 4340 13084
rect 4300 11528 4340 11740
rect 4396 12368 4436 14344
rect 4492 14048 4532 14512
rect 4492 13999 4532 14008
rect 4588 14132 4628 14764
rect 4876 14755 4916 14764
rect 5164 14804 5204 14813
rect 4588 13544 4628 14092
rect 4588 13495 4628 13504
rect 4684 14720 4724 14729
rect 4684 13460 4724 14680
rect 4684 13411 4724 13420
rect 4780 14636 4820 14645
rect 4684 13292 4724 13301
rect 4780 13292 4820 14596
rect 5068 14552 5108 14561
rect 5068 14417 5108 14512
rect 5068 14216 5108 14225
rect 5068 13796 5108 14176
rect 5068 13747 5108 13756
rect 5164 13880 5204 14764
rect 5260 14048 5300 14932
rect 5260 13999 5300 14008
rect 5356 14888 5396 17260
rect 5548 17072 5588 21568
rect 5644 21020 5684 22324
rect 5644 20971 5684 20980
rect 5740 22868 5780 22877
rect 5644 20852 5684 20861
rect 5644 19508 5684 20812
rect 5740 20096 5780 22828
rect 5740 20047 5780 20056
rect 5644 19459 5684 19468
rect 5548 17023 5588 17032
rect 5644 19340 5684 19349
rect 5644 16988 5684 19300
rect 5836 18248 5876 26608
rect 5836 18199 5876 18208
rect 5932 18080 5972 26692
rect 5836 18040 5972 18080
rect 5836 17912 5876 18040
rect 5836 17863 5876 17872
rect 5932 17912 5972 17921
rect 5644 16939 5684 16948
rect 5740 17828 5780 17837
rect 5548 16904 5588 16913
rect 5452 16820 5492 16829
rect 5452 14972 5492 16780
rect 5452 14923 5492 14932
rect 5356 14048 5396 14848
rect 5452 14804 5492 14813
rect 5452 14216 5492 14764
rect 5548 14804 5588 16864
rect 5740 16652 5780 17788
rect 5740 16232 5780 16612
rect 5644 15980 5684 15989
rect 5644 14888 5684 15940
rect 5740 15392 5780 16192
rect 5740 15343 5780 15352
rect 5836 17072 5876 17081
rect 5644 14839 5684 14848
rect 5740 15056 5780 15065
rect 5548 14755 5588 14764
rect 5740 14720 5780 15016
rect 5740 14671 5780 14680
rect 5836 14636 5876 17032
rect 5932 14804 5972 17872
rect 6028 17324 6068 33160
rect 6124 32948 6164 34924
rect 6124 32899 6164 32908
rect 6220 34964 6260 34973
rect 6124 32360 6164 32369
rect 6124 19340 6164 32320
rect 6220 23288 6260 34924
rect 6316 32360 6356 38200
rect 6412 36896 6452 36905
rect 6412 34964 6452 36856
rect 6412 34915 6452 34924
rect 6316 32311 6356 32320
rect 6412 33536 6452 33545
rect 6316 32192 6356 32201
rect 6316 31604 6356 32152
rect 6412 31772 6452 33496
rect 6412 31723 6452 31732
rect 6316 31555 6356 31564
rect 6316 31184 6356 31193
rect 6316 30680 6356 31144
rect 6316 29504 6356 30640
rect 6412 30428 6452 30437
rect 6412 30092 6452 30388
rect 6412 30043 6452 30052
rect 6316 28832 6356 29464
rect 6316 28783 6356 28792
rect 6412 26900 6452 26909
rect 6220 23239 6260 23248
rect 6316 26312 6356 26321
rect 6316 23060 6356 26272
rect 6124 19291 6164 19300
rect 6220 23020 6356 23060
rect 6124 17996 6164 18007
rect 6124 17912 6164 17956
rect 6220 17996 6260 23020
rect 6412 21608 6452 26860
rect 6220 17947 6260 17956
rect 6316 21568 6412 21608
rect 6124 17863 6164 17872
rect 6220 17828 6260 17837
rect 6028 17275 6068 17284
rect 6124 17744 6164 17753
rect 6028 17072 6068 17167
rect 6028 17023 6068 17032
rect 6124 17072 6164 17704
rect 6220 17240 6260 17788
rect 6220 17191 6260 17200
rect 6220 17072 6260 17081
rect 6124 17032 6220 17072
rect 6028 16904 6068 16913
rect 6028 16769 6068 16864
rect 5932 14720 5972 14764
rect 5932 14671 5972 14680
rect 6028 16568 6068 16577
rect 5836 14587 5876 14596
rect 5740 14468 5780 14477
rect 5452 14176 5588 14216
rect 5164 13796 5204 13840
rect 5164 13747 5204 13756
rect 4928 13628 5296 13637
rect 4968 13588 5010 13628
rect 5050 13588 5092 13628
rect 5132 13588 5174 13628
rect 5214 13588 5256 13628
rect 4928 13579 5296 13588
rect 4724 13252 4820 13292
rect 4876 13460 4916 13469
rect 4396 11780 4436 12328
rect 4396 11731 4436 11740
rect 4492 13208 4532 13217
rect 4300 10940 4340 11488
rect 4300 10891 4340 10900
rect 4396 11612 4436 11621
rect 4204 10135 4244 10144
rect 4300 10772 4340 10781
rect 3688 9848 4056 9857
rect 3728 9808 3770 9848
rect 3810 9808 3852 9848
rect 3892 9808 3934 9848
rect 3974 9808 4016 9848
rect 3688 9799 4056 9808
rect 4300 9764 4340 10732
rect 4204 9724 4340 9764
rect 4396 9764 4436 11572
rect 4204 8672 4244 9724
rect 4204 8632 4340 8672
rect 3688 8336 4056 8345
rect 3728 8296 3770 8336
rect 3810 8296 3852 8336
rect 3892 8296 3934 8336
rect 3974 8296 4016 8336
rect 3688 8287 4056 8296
rect 3688 6824 4056 6833
rect 3728 6784 3770 6824
rect 3810 6784 3852 6824
rect 3892 6784 3934 6824
rect 3974 6784 4016 6824
rect 3688 6775 4056 6784
rect 4300 6656 4340 8632
rect 4396 6824 4436 9724
rect 4396 6775 4436 6784
rect 4492 8756 4532 13168
rect 4588 12284 4628 12293
rect 4588 9596 4628 12244
rect 4684 11192 4724 13252
rect 4876 13124 4916 13420
rect 4972 13460 5012 13469
rect 4972 13292 5012 13420
rect 4972 13243 5012 13252
rect 5260 13292 5300 13303
rect 5260 13208 5300 13252
rect 5356 13292 5396 14008
rect 5356 13243 5396 13252
rect 5452 14048 5492 14057
rect 5260 13159 5300 13168
rect 5452 13124 5492 14008
rect 4780 13084 4916 13124
rect 5356 13084 5492 13124
rect 5548 13124 5588 14176
rect 5548 13084 5684 13124
rect 4780 12452 4820 13084
rect 4972 12620 5012 12629
rect 4972 12536 5012 12580
rect 4972 12485 5012 12496
rect 4780 12403 4820 12412
rect 4928 12116 5296 12125
rect 4968 12076 5010 12116
rect 5050 12076 5092 12116
rect 5132 12076 5174 12116
rect 5214 12076 5256 12116
rect 4928 12067 5296 12076
rect 5356 11948 5396 13084
rect 5644 12980 5684 13084
rect 4684 11143 4724 11152
rect 4780 11908 5396 11948
rect 5548 12940 5684 12980
rect 4684 11024 4724 11033
rect 4684 10436 4724 10984
rect 4684 10387 4724 10396
rect 4588 9547 4628 9556
rect 4684 10268 4724 10277
rect 4300 6616 4436 6656
rect 3724 6404 3764 6413
rect 3724 5816 3764 6364
rect 3724 5767 3764 5776
rect 4108 5816 4148 5825
rect 3688 5312 4056 5321
rect 3728 5272 3770 5312
rect 3810 5272 3852 5312
rect 3892 5272 3934 5312
rect 3974 5272 4016 5312
rect 3688 5263 4056 5272
rect 4108 4892 4148 5776
rect 4108 4220 4148 4852
rect 4108 4171 4148 4180
rect 3688 3800 4056 3809
rect 3728 3760 3770 3800
rect 3810 3760 3852 3800
rect 3892 3760 3934 3800
rect 3974 3760 4016 3800
rect 3688 3751 4056 3760
rect 4396 3800 4436 6616
rect 4492 5648 4532 8716
rect 4588 9428 4628 9437
rect 4588 5648 4628 9388
rect 4684 7916 4724 10228
rect 4780 9596 4820 11908
rect 5356 11780 5396 11789
rect 4928 10604 5296 10613
rect 4968 10564 5010 10604
rect 5050 10564 5092 10604
rect 5132 10564 5174 10604
rect 5214 10564 5256 10604
rect 4928 10555 5296 10564
rect 4780 9547 4820 9556
rect 5260 9764 5300 9773
rect 4876 9428 4916 9437
rect 4684 6404 4724 7876
rect 4780 9388 4876 9428
rect 5260 9428 5300 9724
rect 5356 9680 5396 11740
rect 5356 9631 5396 9640
rect 5452 10436 5492 10445
rect 5356 9428 5396 9437
rect 5260 9388 5356 9428
rect 4780 8756 4820 9388
rect 4876 9379 4916 9388
rect 5356 9379 5396 9388
rect 4928 9092 5296 9101
rect 5452 9092 5492 10396
rect 5548 9764 5588 12940
rect 5740 12620 5780 14428
rect 5740 12571 5780 12580
rect 5836 14468 5876 14477
rect 5836 14048 5876 14428
rect 5836 13460 5876 14008
rect 5836 13376 5876 13420
rect 5836 12536 5876 13336
rect 6028 13376 6068 16528
rect 6028 13327 6068 13336
rect 6124 13208 6164 17032
rect 6220 17023 6260 17032
rect 6316 16904 6356 21568
rect 6412 21559 6452 21568
rect 6412 21356 6452 21365
rect 6412 20852 6452 21316
rect 6412 20803 6452 20812
rect 6508 18080 6548 43240
rect 6604 39668 6644 39677
rect 6604 37904 6644 39628
rect 6604 35888 6644 37864
rect 6604 35048 6644 35848
rect 6604 34999 6644 35008
rect 6604 34376 6644 34385
rect 6604 33704 6644 34336
rect 6604 31184 6644 33664
rect 6604 31135 6644 31144
rect 6604 30596 6644 30605
rect 6604 30176 6644 30556
rect 6604 30127 6644 30136
rect 6700 29336 6740 46096
rect 6700 29287 6740 29296
rect 6796 38996 6836 39005
rect 6700 27572 6740 27581
rect 6700 26144 6740 27532
rect 6796 26900 6836 38956
rect 6892 31604 6932 46768
rect 7372 46724 7412 48304
rect 7372 46675 7412 46684
rect 7948 46724 7988 48304
rect 7948 46675 7988 46684
rect 8524 46724 8564 48304
rect 8524 46675 8564 46684
rect 9100 46724 9140 48304
rect 9100 46675 9140 46684
rect 9676 46724 9716 48304
rect 9676 46675 9716 46684
rect 10252 46724 10292 48304
rect 10252 46675 10292 46684
rect 10828 46724 10868 48304
rect 10828 46675 10868 46684
rect 11404 46724 11444 48304
rect 11404 46675 11444 46684
rect 11020 46640 11060 46649
rect 10732 46556 10772 46565
rect 7660 46472 7700 46481
rect 7660 43700 7700 46432
rect 9388 46472 9428 46481
rect 8620 46388 8660 46397
rect 8620 45212 8660 46348
rect 8620 45163 8660 45172
rect 8908 44960 8948 44969
rect 8908 44825 8948 44920
rect 9388 44456 9428 46432
rect 10348 46472 10388 46481
rect 10060 46304 10100 46313
rect 9388 44407 9428 44416
rect 9964 46220 10004 46229
rect 9964 44372 10004 46180
rect 10060 45212 10100 46264
rect 10060 45163 10100 45172
rect 10252 45716 10292 45725
rect 9964 44323 10004 44332
rect 7660 43651 7700 43660
rect 8044 43532 8084 43541
rect 7852 43364 7892 43373
rect 7084 42692 7124 42701
rect 6988 37484 7028 37493
rect 6988 36140 7028 37444
rect 6988 36091 7028 36100
rect 6892 31555 6932 31564
rect 6988 33368 7028 33377
rect 6796 26851 6836 26860
rect 6892 31184 6932 31193
rect 6604 24464 6644 24473
rect 6604 21524 6644 24424
rect 6700 21524 6740 26104
rect 6892 22868 6932 31144
rect 6988 27068 7028 33328
rect 7084 33284 7124 42652
rect 7276 39668 7316 39677
rect 7084 33235 7124 33244
rect 7180 38072 7220 38081
rect 7084 32612 7124 32621
rect 7084 32477 7124 32572
rect 6988 27019 7028 27028
rect 7084 30764 7124 30773
rect 6988 26396 7028 26405
rect 6988 26060 7028 26356
rect 6988 26011 7028 26020
rect 6892 22819 6932 22828
rect 6892 22280 6932 22289
rect 6796 21524 6836 21533
rect 6700 21484 6796 21524
rect 6604 21475 6644 21484
rect 6412 18040 6548 18080
rect 6700 21104 6740 21113
rect 6700 20852 6740 21064
rect 6412 17828 6452 18040
rect 6412 17779 6452 17788
rect 6604 17996 6644 18005
rect 6508 17744 6548 17753
rect 6316 16855 6356 16864
rect 6412 17324 6452 17333
rect 5836 12487 5876 12496
rect 6028 13168 6164 13208
rect 6220 16820 6260 16829
rect 5740 12452 5780 12461
rect 5740 12368 5780 12412
rect 5740 11612 5780 12328
rect 5740 11563 5780 11572
rect 5836 10940 5876 10949
rect 5740 10856 5780 10865
rect 5740 10268 5780 10816
rect 5740 10219 5780 10228
rect 5548 9715 5588 9724
rect 5740 10100 5780 10109
rect 5548 9512 5588 9607
rect 5548 9463 5588 9472
rect 5644 9344 5684 9353
rect 4968 9052 5010 9092
rect 5050 9052 5092 9092
rect 5132 9052 5174 9092
rect 5214 9052 5256 9092
rect 4928 9043 5296 9052
rect 5356 9052 5492 9092
rect 5548 9260 5588 9269
rect 5260 8840 5300 8849
rect 5356 8840 5396 9052
rect 5300 8800 5396 8840
rect 5260 8791 5300 8800
rect 4780 8168 4820 8716
rect 5068 8756 5108 8765
rect 5068 8621 5108 8716
rect 4780 7328 4820 8128
rect 5356 8084 5396 8800
rect 5452 8756 5492 8765
rect 5452 8621 5492 8716
rect 4928 7580 5296 7589
rect 4968 7540 5010 7580
rect 5050 7540 5092 7580
rect 5132 7540 5174 7580
rect 5214 7540 5256 7580
rect 4928 7531 5296 7540
rect 5260 7412 5300 7421
rect 4780 7279 4820 7288
rect 4876 7244 4916 7339
rect 4876 6572 4916 7204
rect 4972 7160 5012 7169
rect 4972 7025 5012 7120
rect 4876 6523 4916 6532
rect 4684 6355 4724 6364
rect 4780 6236 4820 6245
rect 5260 6236 5300 7372
rect 5356 7244 5396 8044
rect 5356 7195 5396 7204
rect 5260 6196 5396 6236
rect 4684 5648 4724 5657
rect 4588 5608 4684 5648
rect 4492 4976 4532 5608
rect 4684 5599 4724 5608
rect 4492 4220 4532 4936
rect 4492 4171 4532 4180
rect 4396 3751 4436 3760
rect 3532 2860 4148 2900
rect 3688 2288 4056 2297
rect 3728 2248 3770 2288
rect 3810 2248 3852 2288
rect 3892 2248 3934 2288
rect 3974 2248 4016 2288
rect 3688 2239 4056 2248
rect 4108 1448 4148 2860
rect 4780 2120 4820 6196
rect 4928 6068 5296 6077
rect 4968 6028 5010 6068
rect 5050 6028 5092 6068
rect 5132 6028 5174 6068
rect 5214 6028 5256 6068
rect 4928 6019 5296 6028
rect 5356 4976 5396 6196
rect 5356 4927 5396 4936
rect 5452 5648 5492 5657
rect 4928 4556 5296 4565
rect 4968 4516 5010 4556
rect 5050 4516 5092 4556
rect 5132 4516 5174 4556
rect 5214 4516 5256 4556
rect 4928 4507 5296 4516
rect 5356 3548 5396 3557
rect 4928 3044 5296 3053
rect 4968 3004 5010 3044
rect 5050 3004 5092 3044
rect 5132 3004 5174 3044
rect 5214 3004 5256 3044
rect 4928 2995 5296 3004
rect 5356 2624 5396 3508
rect 5452 3380 5492 5608
rect 5548 3632 5588 9220
rect 5644 8504 5684 9304
rect 5740 9176 5780 10060
rect 5740 9127 5780 9136
rect 5740 9008 5780 9017
rect 5740 8873 5780 8968
rect 5644 6656 5684 8464
rect 5740 8756 5780 8765
rect 5740 7916 5780 8716
rect 5836 8168 5876 10900
rect 6028 10436 6068 13168
rect 6220 13124 6260 16780
rect 6316 16736 6356 16745
rect 6316 16601 6356 16696
rect 6316 14804 6356 14813
rect 6316 14669 6356 14764
rect 6220 13075 6260 13084
rect 6316 13796 6356 13805
rect 6124 12956 6164 12965
rect 6124 12821 6164 12916
rect 6124 12452 6164 12461
rect 6124 11864 6164 12412
rect 6316 12368 6356 13756
rect 6412 13544 6452 17284
rect 6508 16904 6548 17704
rect 6508 16855 6548 16864
rect 6508 16652 6548 16661
rect 6508 16484 6548 16612
rect 6508 16064 6548 16444
rect 6508 16015 6548 16024
rect 6412 13495 6452 13504
rect 6508 14720 6548 14729
rect 6412 13292 6452 13301
rect 6412 13208 6452 13252
rect 6412 13157 6452 13168
rect 6508 12452 6548 14680
rect 6508 12403 6548 12412
rect 6316 12319 6356 12328
rect 6412 12200 6452 12209
rect 6124 11815 6164 11824
rect 6220 12116 6260 12125
rect 6124 11696 6164 11705
rect 6220 11696 6260 12076
rect 6164 11656 6260 11696
rect 6124 11647 6164 11656
rect 6028 10387 6068 10396
rect 6124 10940 6164 10949
rect 5836 8119 5876 8128
rect 5932 10268 5972 10277
rect 5740 7867 5780 7876
rect 5644 6607 5684 6616
rect 5740 7748 5780 7757
rect 5644 6488 5684 6497
rect 5644 6152 5684 6448
rect 5740 6320 5780 7708
rect 5740 6271 5780 6280
rect 5644 4976 5684 6112
rect 5836 5564 5876 5573
rect 5836 5060 5876 5524
rect 5836 5011 5876 5020
rect 5644 4927 5684 4936
rect 5932 4304 5972 10228
rect 6028 10184 6068 10193
rect 6028 9428 6068 10144
rect 6028 8756 6068 9388
rect 6124 8924 6164 10900
rect 6220 10520 6260 11656
rect 6316 11780 6356 11789
rect 6316 11645 6356 11740
rect 6412 11696 6452 12160
rect 6412 11647 6452 11656
rect 6604 11360 6644 17956
rect 6700 17828 6740 20812
rect 6700 17744 6740 17788
rect 6700 17695 6740 17704
rect 6700 16736 6740 16745
rect 6700 12704 6740 16696
rect 6796 16400 6836 21484
rect 6892 21356 6932 22240
rect 6892 21307 6932 21316
rect 7084 20180 7124 30724
rect 7180 24548 7220 38032
rect 7276 37988 7316 39628
rect 7372 39500 7412 39509
rect 7372 38240 7412 39460
rect 7660 38996 7700 39005
rect 7372 38191 7412 38200
rect 7468 38912 7508 38921
rect 7276 37939 7316 37948
rect 7468 38156 7508 38872
rect 7276 37484 7316 37493
rect 7276 37349 7316 37444
rect 7468 37484 7508 38116
rect 7276 35132 7316 35141
rect 7276 34292 7316 35092
rect 7276 33704 7316 34252
rect 7276 33569 7316 33664
rect 7276 32780 7316 32789
rect 7276 32024 7316 32740
rect 7276 31975 7316 31984
rect 7372 31184 7412 31193
rect 7276 31016 7316 31025
rect 7276 28664 7316 30976
rect 7276 28615 7316 28624
rect 7276 26816 7316 26825
rect 7276 26228 7316 26776
rect 7276 26179 7316 26188
rect 7180 24413 7220 24508
rect 7276 24632 7316 24641
rect 7180 23624 7220 23633
rect 7180 22364 7220 23584
rect 7180 22315 7220 22324
rect 7276 22280 7316 24592
rect 7372 23036 7412 31144
rect 7468 30764 7508 37444
rect 7660 38240 7700 38956
rect 7660 37484 7700 38200
rect 7660 37435 7700 37444
rect 7756 37400 7796 37409
rect 7756 37232 7796 37360
rect 7756 37183 7796 37192
rect 7660 35132 7700 35141
rect 7660 33620 7700 35092
rect 7660 33571 7700 33580
rect 7468 30715 7508 30724
rect 7564 32864 7604 32873
rect 7468 30596 7508 30605
rect 7468 30092 7508 30556
rect 7468 30043 7508 30052
rect 7468 29840 7508 29849
rect 7468 25472 7508 29800
rect 7468 25337 7508 25432
rect 7468 25136 7508 25145
rect 7468 23876 7508 25096
rect 7468 23827 7508 23836
rect 7372 22987 7412 22996
rect 7276 22231 7316 22240
rect 6988 20140 7124 20180
rect 7180 21692 7220 21701
rect 7180 20180 7220 21652
rect 7180 20140 7316 20180
rect 6892 18500 6932 18509
rect 6892 17744 6932 18460
rect 6988 17996 7028 20140
rect 6988 17947 7028 17956
rect 7084 19340 7124 19349
rect 6892 17695 6932 17704
rect 6988 17828 7028 17837
rect 7084 17828 7124 19300
rect 7276 18500 7316 20140
rect 7564 18584 7604 32824
rect 7756 32864 7796 32873
rect 7756 32729 7796 32824
rect 7756 31268 7796 31277
rect 7756 30680 7796 31228
rect 7852 30932 7892 43324
rect 7852 30883 7892 30892
rect 7948 34460 7988 34469
rect 7756 29924 7796 30640
rect 7756 29875 7796 29884
rect 7852 30764 7892 30773
rect 7756 29756 7796 29765
rect 7756 29084 7796 29716
rect 7660 29044 7756 29084
rect 7660 26396 7700 29044
rect 7756 29035 7796 29044
rect 7660 26347 7700 26356
rect 7756 26900 7796 26909
rect 7028 17788 7124 17828
rect 7180 17996 7220 18005
rect 6988 17240 7028 17788
rect 6988 17191 7028 17200
rect 7084 17660 7124 17669
rect 6796 16351 6836 16360
rect 6988 16820 7028 16829
rect 6892 16316 6932 16325
rect 6796 16148 6836 16157
rect 6796 15644 6836 16108
rect 6796 12788 6836 15604
rect 6892 13208 6932 16276
rect 6988 13292 7028 16780
rect 7084 16064 7124 17620
rect 7180 16988 7220 17956
rect 7276 17996 7316 18460
rect 7276 17947 7316 17956
rect 7372 18544 7604 18584
rect 7660 26060 7700 26069
rect 7660 25388 7700 26020
rect 7276 17492 7316 17501
rect 7276 17357 7316 17452
rect 7372 17240 7412 18544
rect 7660 18080 7700 25348
rect 7756 25136 7796 26860
rect 7756 24716 7796 25096
rect 7756 24667 7796 24676
rect 7756 23792 7796 23801
rect 7756 23120 7796 23752
rect 7756 23071 7796 23080
rect 7660 18031 7700 18040
rect 7756 22280 7796 22289
rect 7756 18500 7796 22240
rect 7852 21692 7892 30724
rect 7948 24548 7988 34420
rect 8044 30596 8084 43492
rect 8620 43448 8660 43457
rect 8620 43313 8660 43408
rect 10060 41852 10100 41861
rect 9484 39836 9524 39845
rect 8332 39668 8372 39677
rect 8140 38996 8180 39005
rect 8180 38956 8276 38996
rect 8140 38947 8180 38956
rect 8236 38156 8276 38956
rect 8044 30547 8084 30556
rect 8140 37988 8180 37997
rect 8044 30428 8084 30437
rect 8044 24716 8084 30388
rect 8140 29168 8180 37948
rect 8236 37232 8276 38116
rect 8236 37183 8276 37192
rect 8332 38408 8372 39628
rect 8908 39668 8948 39677
rect 8236 35132 8276 35141
rect 8236 33116 8276 35092
rect 8236 32444 8276 33076
rect 8236 32395 8276 32404
rect 8140 29119 8180 29128
rect 8236 31604 8276 31613
rect 8140 26816 8180 26825
rect 8140 25388 8180 26776
rect 8140 25339 8180 25348
rect 8236 25220 8276 31564
rect 8332 29924 8372 38368
rect 8812 38912 8852 38921
rect 8812 37652 8852 38872
rect 8812 37603 8852 37612
rect 8908 38828 8948 39628
rect 8908 38240 8948 38788
rect 8620 36476 8660 36485
rect 8524 35300 8564 35309
rect 8524 34376 8564 35260
rect 8620 35132 8660 36436
rect 8620 35083 8660 35092
rect 8524 33452 8564 34336
rect 8428 30680 8468 30689
rect 8428 30428 8468 30640
rect 8428 30379 8468 30388
rect 8332 29875 8372 29884
rect 8524 28832 8564 33412
rect 8716 32948 8756 32957
rect 8716 32276 8756 32908
rect 8716 32108 8756 32236
rect 8620 31436 8660 31445
rect 8620 30596 8660 31396
rect 8620 30547 8660 30556
rect 8716 31352 8756 32068
rect 8524 28783 8564 28792
rect 8620 28916 8660 28925
rect 8620 28496 8660 28876
rect 8620 28447 8660 28456
rect 8428 28328 8468 28337
rect 8044 24667 8084 24676
rect 8140 25180 8276 25220
rect 8332 26060 8372 26069
rect 7988 24508 8084 24548
rect 7948 24499 7988 24508
rect 8044 23204 8084 24508
rect 8140 23792 8180 25180
rect 8140 23743 8180 23752
rect 8236 25052 8276 25061
rect 8236 24632 8276 25012
rect 7852 21643 7892 21652
rect 7948 23164 8084 23204
rect 7948 21104 7988 23164
rect 8140 23120 8180 23129
rect 8044 23036 8084 23045
rect 8044 22280 8084 22996
rect 8044 22112 8084 22240
rect 8044 22063 8084 22072
rect 8140 22364 8180 23080
rect 7948 21055 7988 21064
rect 7756 17660 7796 18460
rect 8044 19088 8084 19097
rect 8044 18500 8084 19048
rect 8044 18451 8084 18460
rect 8140 18332 8180 22324
rect 7564 17620 7796 17660
rect 8044 18292 8180 18332
rect 8236 20852 8276 24592
rect 8332 24548 8372 26020
rect 8332 24499 8372 24508
rect 8332 23876 8372 23885
rect 8332 23204 8372 23836
rect 8332 23155 8372 23164
rect 8428 23060 8468 28288
rect 8716 27152 8756 31312
rect 8908 32108 8948 38200
rect 9004 39500 9044 39509
rect 9004 37484 9044 39460
rect 9388 38912 9428 38921
rect 9388 37988 9428 38872
rect 9388 37939 9428 37948
rect 9004 37435 9044 37444
rect 9292 37484 9332 37493
rect 9292 37232 9332 37444
rect 9292 36560 9332 37192
rect 9292 36511 9332 36520
rect 9196 35888 9236 35897
rect 9196 35384 9236 35848
rect 9292 35720 9332 35729
rect 9292 35468 9332 35680
rect 9484 35636 9524 39796
rect 9676 39080 9716 39089
rect 9484 35587 9524 35596
rect 9580 36728 9620 36737
rect 9292 35419 9332 35428
rect 9196 35335 9236 35344
rect 9484 35132 9524 35141
rect 9388 34964 9428 34973
rect 9388 34460 9428 34924
rect 9484 34628 9524 35092
rect 9484 34579 9524 34588
rect 9388 34411 9428 34420
rect 9292 34376 9332 34385
rect 9100 33620 9140 33629
rect 8908 31520 8948 32068
rect 8716 27103 8756 27112
rect 8812 31268 8852 31277
rect 8524 26396 8564 26405
rect 8524 24548 8564 26356
rect 8716 25976 8756 25985
rect 8620 25892 8660 25901
rect 8620 25220 8660 25852
rect 8716 25388 8756 25936
rect 8716 25339 8756 25348
rect 8620 25171 8660 25180
rect 8620 24548 8660 24557
rect 8524 24508 8620 24548
rect 8620 24499 8660 24508
rect 7372 17191 7412 17200
rect 7468 17576 7508 17585
rect 7468 17240 7508 17536
rect 7468 17191 7508 17200
rect 7180 16939 7220 16948
rect 7276 17156 7316 17165
rect 7276 16988 7316 17116
rect 7468 17072 7508 17081
rect 7372 16988 7412 17016
rect 7276 16948 7372 16988
rect 7180 16400 7220 16409
rect 7180 16232 7220 16360
rect 7180 16183 7220 16192
rect 7276 16316 7316 16948
rect 7372 16939 7412 16948
rect 7084 15929 7124 16024
rect 7084 15728 7124 15737
rect 7124 15688 7220 15728
rect 7084 15679 7124 15688
rect 6988 13243 7028 13252
rect 7084 15476 7124 15485
rect 7084 14720 7124 15436
rect 6892 13159 6932 13168
rect 7084 13124 7124 14680
rect 7180 14048 7220 15688
rect 7276 15644 7316 16276
rect 7276 15595 7316 15604
rect 7372 16820 7412 16829
rect 7276 15140 7316 15235
rect 7276 15091 7316 15100
rect 7372 15056 7412 16780
rect 7372 15007 7412 15016
rect 7180 13999 7220 14008
rect 7276 14972 7316 14981
rect 7276 13964 7316 14932
rect 7276 13915 7316 13924
rect 7372 14300 7412 14309
rect 7084 13075 7124 13084
rect 7180 13796 7220 13805
rect 6892 13040 6932 13049
rect 6892 12956 6932 13000
rect 7180 12980 7220 13756
rect 7372 13124 7412 14260
rect 7372 13075 7412 13084
rect 6892 12905 6932 12916
rect 7084 12956 7124 12965
rect 7180 12931 7220 12940
rect 7372 12956 7412 12965
rect 6796 12748 7028 12788
rect 6700 12655 6740 12664
rect 6892 12620 6932 12629
rect 6316 11192 6356 11201
rect 6316 10856 6356 11152
rect 6316 10807 6356 10816
rect 6412 11024 6452 11033
rect 6220 10471 6260 10480
rect 6316 10688 6356 10697
rect 6220 10352 6260 10361
rect 6220 10100 6260 10312
rect 6220 10051 6260 10060
rect 6124 8875 6164 8884
rect 6220 8840 6260 8880
rect 6220 8756 6260 8800
rect 6028 8716 6164 8756
rect 6028 8588 6068 8597
rect 6028 7328 6068 8548
rect 6028 7279 6068 7288
rect 6124 7916 6164 8716
rect 6124 6992 6164 7876
rect 6124 6943 6164 6952
rect 6220 6740 6260 8716
rect 6220 6691 6260 6700
rect 6220 5732 6260 5741
rect 6220 5396 6260 5692
rect 6316 5480 6356 10648
rect 6412 9596 6452 10984
rect 6508 10940 6548 10949
rect 6508 10268 6548 10900
rect 6604 10268 6644 11320
rect 6796 12452 6836 12461
rect 6700 10268 6740 10277
rect 6604 10228 6700 10268
rect 6508 10219 6548 10228
rect 6700 10219 6740 10228
rect 6700 10100 6740 10109
rect 6412 8840 6452 9556
rect 6412 8791 6452 8800
rect 6508 10016 6548 10025
rect 6316 5431 6356 5440
rect 6220 5347 6260 5356
rect 5932 4255 5972 4264
rect 5548 3583 5588 3592
rect 5644 4220 5684 4229
rect 5644 3548 5684 4180
rect 6508 3884 6548 9976
rect 6604 9512 6644 9521
rect 6604 8672 6644 9472
rect 6604 8623 6644 8632
rect 6700 7916 6740 10060
rect 6796 9596 6836 12412
rect 6892 11780 6932 12580
rect 6988 12536 7028 12748
rect 6988 12487 7028 12496
rect 6892 11731 6932 11740
rect 6988 12368 7028 12377
rect 6796 9547 6836 9556
rect 6892 10772 6932 10781
rect 6796 8840 6836 8935
rect 6796 8791 6836 8800
rect 6700 7867 6740 7876
rect 6796 8672 6836 8681
rect 6796 7244 6836 8632
rect 6892 8672 6932 10732
rect 6988 10352 7028 12328
rect 7084 11948 7124 12916
rect 7180 12872 7220 12881
rect 7180 12620 7220 12832
rect 7180 12571 7220 12580
rect 7276 12704 7316 12713
rect 7180 12452 7220 12492
rect 7180 12368 7220 12412
rect 7180 12116 7220 12328
rect 7276 12284 7316 12664
rect 7276 12235 7316 12244
rect 7180 12067 7220 12076
rect 7084 11908 7220 11948
rect 6988 10303 7028 10312
rect 7084 11780 7124 11789
rect 6892 8623 6932 8632
rect 6988 9428 7028 9437
rect 6988 8252 7028 9388
rect 6988 8203 7028 8212
rect 6796 7195 6836 7204
rect 6700 6404 6740 6413
rect 6700 5144 6740 6364
rect 7084 5564 7124 11740
rect 7180 9008 7220 11908
rect 7180 8959 7220 8968
rect 7276 11192 7316 11201
rect 7084 5515 7124 5524
rect 7180 8840 7220 8849
rect 6700 5095 6740 5104
rect 6988 5396 7028 5405
rect 6508 3835 6548 3844
rect 6988 3968 7028 5356
rect 7180 4472 7220 8800
rect 7276 6908 7316 11152
rect 7276 6859 7316 6868
rect 7372 5060 7412 12916
rect 7468 12704 7508 17032
rect 7564 16400 7604 17620
rect 7756 17324 7796 17333
rect 7756 17240 7796 17284
rect 7756 17189 7796 17200
rect 7948 17156 7988 17165
rect 7564 15728 7604 16360
rect 7564 14804 7604 15688
rect 7564 14636 7604 14764
rect 7564 14587 7604 14596
rect 7660 17072 7700 17081
rect 7660 14636 7700 17032
rect 7852 17072 7892 17081
rect 7852 16937 7892 17032
rect 7660 14587 7700 14596
rect 7756 16736 7796 16745
rect 7468 12655 7508 12664
rect 7564 14384 7604 14393
rect 7468 12536 7508 12545
rect 7468 12368 7508 12496
rect 7468 12319 7508 12328
rect 7564 12200 7604 14344
rect 7756 12788 7796 16696
rect 7852 16484 7892 16493
rect 7852 14804 7892 16444
rect 7948 15056 7988 17116
rect 7948 15007 7988 15016
rect 7852 14755 7892 14764
rect 7948 14888 7988 14897
rect 7948 14720 7988 14848
rect 7756 12739 7796 12748
rect 7852 14636 7892 14645
rect 7468 12160 7604 12200
rect 7660 12368 7700 12377
rect 7468 6236 7508 12160
rect 7564 11024 7604 11033
rect 7564 10604 7604 10984
rect 7660 10856 7700 12328
rect 7852 11276 7892 14596
rect 7948 13376 7988 14680
rect 7948 13327 7988 13336
rect 7852 11227 7892 11236
rect 7948 13124 7988 13133
rect 7756 11024 7796 11033
rect 7948 11024 7988 13084
rect 8044 12704 8084 18292
rect 8140 16232 8180 16327
rect 8140 16183 8180 16192
rect 8140 16064 8180 16073
rect 8140 13544 8180 16024
rect 8236 15644 8276 20812
rect 8236 15595 8276 15604
rect 8332 23020 8468 23060
rect 8524 23792 8564 23801
rect 8332 18668 8372 23020
rect 8524 22952 8564 23752
rect 8620 22952 8660 22961
rect 8524 22912 8620 22952
rect 8620 22364 8660 22912
rect 8332 16316 8372 18628
rect 8236 15476 8276 15485
rect 8236 14552 8276 15436
rect 8236 14503 8276 14512
rect 8332 14552 8372 16276
rect 8428 20852 8468 20861
rect 8428 15728 8468 20812
rect 8524 19172 8564 19181
rect 8524 17996 8564 19132
rect 8524 17947 8564 17956
rect 8620 17828 8660 22324
rect 8524 17788 8660 17828
rect 8716 21524 8756 21533
rect 8716 20600 8756 21484
rect 8524 16820 8564 17788
rect 8620 17660 8660 17669
rect 8620 16988 8660 17620
rect 8620 16939 8660 16948
rect 8524 16780 8660 16820
rect 8524 16652 8564 16661
rect 8524 15812 8564 16612
rect 8620 16232 8660 16780
rect 8716 16316 8756 20560
rect 8812 16484 8852 31228
rect 8908 30848 8948 31480
rect 8908 28580 8948 30808
rect 8908 27656 8948 28540
rect 8908 27607 8948 27616
rect 9004 33452 9044 33461
rect 9004 26564 9044 33412
rect 9100 31352 9140 33580
rect 9292 33536 9332 34336
rect 9196 33284 9236 33293
rect 9196 32864 9236 33244
rect 9292 33140 9332 33496
rect 9580 33140 9620 36688
rect 9676 35804 9716 39040
rect 9772 38912 9812 38921
rect 9964 38912 10004 38921
rect 9772 38777 9812 38872
rect 9868 38872 9964 38912
rect 9676 35755 9716 35764
rect 9772 37232 9812 37241
rect 9292 33100 9428 33140
rect 9196 32815 9236 32824
rect 9388 33032 9428 33100
rect 9100 31303 9140 31312
rect 9196 31940 9236 31949
rect 9100 30176 9140 30185
rect 9100 29336 9140 30136
rect 9100 29287 9140 29296
rect 8908 26524 9044 26564
rect 9100 29168 9140 29177
rect 8908 22532 8948 26524
rect 9100 26480 9140 29128
rect 8908 22483 8948 22492
rect 9004 26440 9140 26480
rect 9004 23120 9044 26440
rect 9100 25304 9140 25313
rect 9100 24800 9140 25264
rect 9100 24751 9140 24760
rect 8908 22364 8948 22373
rect 8908 21440 8948 22324
rect 8908 21391 8948 21400
rect 9004 21020 9044 23080
rect 9100 23708 9140 23717
rect 9100 21692 9140 23668
rect 9196 23036 9236 31900
rect 9388 31436 9428 32992
rect 9388 31387 9428 31396
rect 9484 33100 9620 33140
rect 9676 35636 9716 35645
rect 9292 31352 9332 31361
rect 9292 30596 9332 31312
rect 9292 25640 9332 30556
rect 9388 30932 9428 30941
rect 9388 30008 9428 30892
rect 9388 29959 9428 29968
rect 9388 29840 9428 29849
rect 9388 29252 9428 29800
rect 9388 29203 9428 29212
rect 9292 25591 9332 25600
rect 9388 28496 9428 28505
rect 9388 25388 9428 28456
rect 9484 28244 9524 33100
rect 9580 33032 9620 33041
rect 9580 32897 9620 32992
rect 9580 32696 9620 32705
rect 9580 29252 9620 32656
rect 9676 31604 9716 35596
rect 9676 31555 9716 31564
rect 9676 31436 9716 31445
rect 9676 29672 9716 31396
rect 9772 29840 9812 37192
rect 9868 32360 9908 38872
rect 9964 38863 10004 38872
rect 10060 37484 10100 41812
rect 9964 37444 10100 37484
rect 9964 35720 10004 37444
rect 9964 35671 10004 35680
rect 10060 37316 10100 37325
rect 9964 35468 10004 35477
rect 9964 35333 10004 35428
rect 10060 34880 10100 37276
rect 10156 36308 10196 36317
rect 10156 35972 10196 36268
rect 10156 35923 10196 35932
rect 10060 34831 10100 34840
rect 10060 34460 10100 34469
rect 9868 32311 9908 32320
rect 9964 34124 10004 34133
rect 9868 31436 9908 31445
rect 9868 30848 9908 31396
rect 9868 30799 9908 30808
rect 9772 29791 9812 29800
rect 9868 30680 9908 30689
rect 9676 29632 9812 29672
rect 9580 29203 9620 29212
rect 9676 29000 9716 29009
rect 9580 28412 9620 28440
rect 9676 28412 9716 28960
rect 9620 28372 9716 28412
rect 9580 28363 9620 28372
rect 9484 28204 9620 28244
rect 9388 25339 9428 25348
rect 9484 28076 9524 28085
rect 9292 25304 9332 25313
rect 9292 24632 9332 25264
rect 9292 24583 9332 24592
rect 9196 22987 9236 22996
rect 9388 23540 9428 23549
rect 9100 21643 9140 21652
rect 9196 22280 9236 22289
rect 9004 20971 9044 20980
rect 9100 21440 9140 21449
rect 9004 20852 9044 20861
rect 8812 16435 8852 16444
rect 8908 20096 8948 20105
rect 8716 16276 8852 16316
rect 8620 16192 8756 16232
rect 8524 15763 8564 15772
rect 8428 15679 8468 15688
rect 8620 15644 8660 15653
rect 8332 14503 8372 14512
rect 8428 15560 8468 15569
rect 8428 14468 8468 15520
rect 8428 14419 8468 14428
rect 8524 15476 8564 15485
rect 8140 13495 8180 13504
rect 8236 14384 8276 14393
rect 8044 12655 8084 12664
rect 8140 13292 8180 13301
rect 8044 11948 8084 11957
rect 8044 11813 8084 11908
rect 7796 10984 7988 11024
rect 8044 11444 8084 11453
rect 7756 10975 7796 10984
rect 8044 10856 8084 11404
rect 7660 10816 7988 10856
rect 7564 8756 7604 10564
rect 7852 10688 7892 10697
rect 7756 10436 7796 10445
rect 7756 9512 7796 10396
rect 7756 9463 7796 9472
rect 7564 8707 7604 8716
rect 7660 9428 7700 9437
rect 7564 6404 7604 6413
rect 7564 6269 7604 6364
rect 7468 6187 7508 6196
rect 7660 5564 7700 9388
rect 7660 5515 7700 5524
rect 7756 6320 7796 6329
rect 7756 5648 7796 6280
rect 7372 5011 7412 5020
rect 7468 4892 7508 4901
rect 7180 4423 7220 4432
rect 7372 4724 7412 4733
rect 5644 3499 5684 3508
rect 5452 3331 5492 3340
rect 6988 3380 7028 3928
rect 7084 3380 7124 3408
rect 6988 3340 7084 3380
rect 5356 2575 5396 2584
rect 6988 2624 7028 3340
rect 7084 3331 7124 3340
rect 6988 2575 7028 2584
rect 7372 2624 7412 4684
rect 7468 4304 7508 4852
rect 7468 4255 7508 4264
rect 7756 4892 7796 5608
rect 7468 4136 7508 4145
rect 7468 3632 7508 4096
rect 7756 3716 7796 4852
rect 7852 4388 7892 10648
rect 7948 8084 7988 10816
rect 8044 10807 8084 10816
rect 7948 8035 7988 8044
rect 8140 10268 8180 13252
rect 8140 8840 8180 10228
rect 8044 7916 8084 7925
rect 7948 7748 7988 7757
rect 7948 5732 7988 7708
rect 7948 5683 7988 5692
rect 7852 4339 7892 4348
rect 7756 3667 7796 3676
rect 7468 3583 7508 3592
rect 8044 2900 8084 7876
rect 8140 7916 8180 8800
rect 8140 7867 8180 7876
rect 8140 7664 8180 7673
rect 8140 4976 8180 7624
rect 8140 4640 8180 4936
rect 8140 4220 8180 4600
rect 8236 4892 8276 14344
rect 8428 14300 8468 14309
rect 8332 14048 8372 14057
rect 8332 13292 8372 14008
rect 8428 13712 8468 14260
rect 8524 13796 8564 15436
rect 8620 14048 8660 15604
rect 8716 14384 8756 16192
rect 8716 14335 8756 14344
rect 8716 14216 8756 14225
rect 8716 14081 8756 14176
rect 8620 13999 8660 14008
rect 8524 13747 8564 13756
rect 8620 13880 8660 13889
rect 8620 13745 8660 13840
rect 8428 13663 8468 13672
rect 8332 13243 8372 13252
rect 8428 13544 8468 13553
rect 8332 13040 8372 13049
rect 8332 12452 8372 13000
rect 8332 12403 8372 12412
rect 8332 11108 8372 11117
rect 8332 10268 8372 11068
rect 8428 10940 8468 13504
rect 8716 13208 8756 13217
rect 8620 12788 8660 12797
rect 8428 10688 8468 10900
rect 8428 10639 8468 10648
rect 8524 12200 8564 12209
rect 8428 10268 8468 10296
rect 8332 10228 8428 10268
rect 8332 9428 8372 10228
rect 8428 10219 8468 10228
rect 8332 9379 8372 9388
rect 8428 10100 8468 10109
rect 8332 9176 8372 9185
rect 8332 8000 8372 9136
rect 8332 7951 8372 7960
rect 8332 7832 8372 7841
rect 8332 5480 8372 7792
rect 8332 5431 8372 5440
rect 8428 5732 8468 10060
rect 8524 8840 8564 12160
rect 8620 11864 8660 12748
rect 8716 12284 8756 13168
rect 8812 13040 8852 16276
rect 8812 12991 8852 13000
rect 8716 12235 8756 12244
rect 8812 12620 8852 12629
rect 8620 11824 8756 11864
rect 8524 8791 8564 8800
rect 8620 11696 8660 11705
rect 8524 8168 8564 8177
rect 8524 8033 8564 8128
rect 8236 4304 8276 4852
rect 8236 4255 8276 4264
rect 8428 4556 8468 5692
rect 8140 4171 8180 4180
rect 8236 4136 8276 4145
rect 8428 4136 8468 4516
rect 8276 4096 8468 4136
rect 8524 7580 8564 7589
rect 8236 4087 8276 4096
rect 7372 2575 7412 2584
rect 7948 2860 8084 2900
rect 8236 2876 8276 2885
rect 5740 2456 5780 2465
rect 5740 2321 5780 2416
rect 4780 2071 4820 2080
rect 4928 1532 5296 1541
rect 4968 1492 5010 1532
rect 5050 1492 5092 1532
rect 5132 1492 5174 1532
rect 5214 1492 5256 1532
rect 4928 1483 5296 1492
rect 4108 1399 4148 1408
rect 5644 1448 5684 1457
rect 4492 944 4532 953
rect 3916 104 3956 113
rect 1016 0 1096 80
rect 1592 0 1672 80
rect 2168 0 2248 80
rect 2744 0 2824 80
rect 3320 0 3400 80
rect 3896 64 3916 80
rect 4492 80 4532 904
rect 5068 188 5108 197
rect 5068 80 5108 148
rect 5644 80 5684 1408
rect 6220 1448 6260 1457
rect 6220 80 6260 1408
rect 6796 1280 6836 1289
rect 6796 80 6836 1240
rect 7372 272 7412 281
rect 7372 80 7412 232
rect 7948 80 7988 2860
rect 8236 2741 8276 2836
rect 8524 80 8564 7540
rect 8620 4052 8660 11656
rect 8716 7244 8756 11824
rect 8812 11612 8852 12580
rect 8812 11563 8852 11572
rect 8908 11024 8948 20056
rect 9004 20012 9044 20812
rect 9004 19963 9044 19972
rect 9100 19340 9140 21400
rect 8812 10984 8948 11024
rect 9004 19300 9140 19340
rect 8812 8756 8852 10984
rect 8908 10856 8948 10865
rect 8908 8924 8948 10816
rect 8908 8875 8948 8884
rect 8908 8756 8948 8765
rect 8812 8716 8908 8756
rect 8716 7195 8756 7204
rect 8812 6404 8852 6413
rect 8812 5816 8852 6364
rect 8812 5767 8852 5776
rect 8908 4220 8948 8716
rect 9004 8084 9044 19300
rect 9100 19172 9140 19181
rect 9100 16484 9140 19132
rect 9196 17660 9236 22240
rect 9292 22196 9332 22205
rect 9292 21608 9332 22156
rect 9292 21559 9332 21568
rect 9292 20852 9332 20861
rect 9292 20264 9332 20812
rect 9292 20215 9332 20224
rect 9292 20012 9332 20021
rect 9292 19004 9332 19972
rect 9292 18955 9332 18964
rect 9388 18080 9428 23500
rect 9484 21524 9524 28036
rect 9580 25556 9620 28204
rect 9676 26984 9716 28372
rect 9772 27740 9812 29632
rect 9868 28496 9908 30640
rect 9868 28447 9908 28456
rect 9772 27691 9812 27700
rect 9772 27572 9812 27581
rect 9812 27532 9908 27572
rect 9772 27523 9812 27532
rect 9676 26935 9716 26944
rect 9772 26816 9812 26825
rect 9772 25556 9812 26776
rect 9580 25516 9716 25556
rect 9484 21475 9524 21484
rect 9580 25388 9620 25397
rect 9580 22028 9620 25348
rect 9676 24884 9716 25516
rect 9772 25507 9812 25516
rect 9868 26060 9908 27532
rect 9676 24835 9716 24844
rect 9772 25220 9812 25229
rect 9580 21020 9620 21988
rect 9484 20980 9620 21020
rect 9676 22700 9716 22709
rect 9484 20180 9524 20980
rect 9580 20852 9620 20861
rect 9580 20348 9620 20812
rect 9580 20299 9620 20308
rect 9484 20140 9620 20180
rect 9292 18040 9428 18080
rect 9484 18500 9524 18509
rect 9292 17828 9332 18040
rect 9292 17779 9332 17788
rect 9388 17912 9428 17921
rect 9196 17620 9332 17660
rect 9100 16444 9236 16484
rect 9100 16316 9140 16325
rect 9100 15728 9140 16276
rect 9100 15679 9140 15688
rect 9100 15560 9140 15569
rect 9100 14636 9140 15520
rect 9100 14587 9140 14596
rect 9100 14384 9140 14393
rect 9100 13544 9140 14344
rect 9100 13495 9140 13504
rect 9100 13376 9140 13385
rect 9100 11612 9140 13336
rect 9196 12620 9236 16444
rect 9196 12571 9236 12580
rect 9196 12452 9236 12461
rect 9196 12116 9236 12412
rect 9196 12067 9236 12076
rect 9292 11948 9332 17620
rect 9100 11563 9140 11572
rect 9196 11908 9332 11948
rect 9100 11360 9140 11369
rect 9100 10940 9140 11320
rect 9100 10891 9140 10900
rect 9196 10352 9236 11908
rect 9196 10303 9236 10312
rect 9292 11780 9332 11789
rect 9100 9596 9140 9605
rect 9100 8924 9140 9556
rect 9292 9596 9332 11740
rect 9388 9680 9428 17872
rect 9484 17660 9524 18460
rect 9484 17611 9524 17620
rect 9580 16988 9620 20140
rect 9580 15980 9620 16948
rect 9580 15931 9620 15940
rect 9484 15896 9524 15905
rect 9484 14972 9524 15856
rect 9484 14923 9524 14932
rect 9580 15476 9620 15485
rect 9580 14804 9620 15436
rect 9580 14755 9620 14764
rect 9484 14636 9524 14645
rect 9484 14468 9524 14596
rect 9484 13376 9524 14428
rect 9484 13327 9524 13336
rect 9580 14552 9620 14561
rect 9580 12980 9620 14512
rect 9676 14552 9716 22660
rect 9772 17912 9812 25180
rect 9868 22700 9908 26020
rect 9964 24044 10004 34084
rect 10060 30680 10100 34420
rect 10156 33704 10196 33713
rect 10156 33200 10196 33664
rect 10156 33151 10196 33160
rect 10156 32864 10196 32875
rect 10156 32780 10196 32824
rect 10156 32731 10196 32740
rect 10156 32528 10196 32537
rect 10156 32393 10196 32488
rect 10060 30631 10100 30640
rect 10156 30512 10196 30521
rect 10060 29840 10100 29849
rect 10060 29504 10100 29800
rect 10156 29672 10196 30472
rect 10252 30092 10292 45676
rect 10348 45128 10388 46432
rect 10348 45079 10388 45088
rect 10540 45800 10580 45809
rect 10540 42860 10580 45760
rect 10636 44960 10676 44969
rect 10636 44792 10676 44920
rect 10636 44743 10676 44752
rect 10732 44456 10772 46516
rect 10828 46472 10868 46481
rect 10828 45212 10868 46432
rect 10828 45163 10868 45172
rect 10732 44407 10772 44416
rect 10924 45044 10964 45053
rect 10540 42811 10580 42820
rect 10732 44288 10772 44297
rect 10252 30043 10292 30052
rect 10348 38996 10388 39005
rect 10156 29632 10292 29672
rect 10060 29464 10196 29504
rect 10156 29420 10196 29464
rect 10156 29371 10196 29380
rect 10060 29336 10100 29345
rect 10060 29252 10100 29296
rect 10060 29201 10100 29212
rect 10156 29168 10196 29177
rect 10252 29168 10292 29632
rect 10196 29128 10292 29168
rect 10156 29119 10196 29128
rect 10060 29000 10100 29009
rect 10060 28832 10100 28960
rect 10252 29000 10292 29009
rect 10060 28328 10100 28792
rect 10156 28916 10196 28925
rect 10156 28412 10196 28876
rect 10156 28363 10196 28372
rect 10060 28279 10100 28288
rect 10156 27488 10196 27497
rect 10060 27236 10100 27245
rect 10060 27101 10100 27196
rect 10060 26228 10100 26323
rect 10060 26179 10100 26188
rect 10060 26060 10100 26071
rect 10060 25976 10100 26020
rect 10060 25927 10100 25936
rect 9964 23995 10004 24004
rect 10060 23792 10100 23801
rect 10060 23657 10100 23752
rect 10060 23288 10100 23297
rect 9868 22651 9908 22660
rect 9964 23120 10004 23129
rect 9964 22616 10004 23080
rect 10060 23036 10100 23248
rect 10060 22987 10100 22996
rect 9964 22567 10004 22576
rect 9868 22532 9908 22541
rect 9868 22448 9908 22492
rect 9868 22408 10004 22448
rect 9772 17863 9812 17872
rect 9868 22280 9908 22289
rect 9868 16316 9908 22240
rect 9964 18416 10004 22408
rect 10156 22280 10196 27448
rect 10252 27488 10292 28960
rect 10252 25892 10292 27448
rect 10348 27488 10388 38956
rect 10444 37484 10484 37493
rect 10444 35972 10484 37444
rect 10732 37316 10772 44248
rect 10732 37267 10772 37276
rect 10828 41180 10868 41189
rect 10828 36896 10868 41140
rect 10828 36847 10868 36856
rect 10636 36728 10676 36737
rect 10540 36560 10580 36569
rect 10540 36308 10580 36520
rect 10540 36259 10580 36268
rect 10444 34964 10484 35932
rect 10540 35888 10580 35897
rect 10540 35132 10580 35848
rect 10540 35083 10580 35092
rect 10444 34924 10580 34964
rect 10444 33620 10484 33629
rect 10444 33284 10484 33580
rect 10444 32444 10484 33244
rect 10444 32395 10484 32404
rect 10540 32276 10580 34924
rect 10636 34460 10676 36688
rect 10732 36644 10772 36653
rect 10732 35048 10772 36604
rect 10732 34999 10772 35008
rect 10828 35888 10868 35897
rect 10636 33032 10676 34420
rect 10636 32983 10676 32992
rect 10732 34208 10772 34217
rect 10636 32864 10676 32873
rect 10636 32696 10676 32824
rect 10636 32647 10676 32656
rect 10444 32236 10580 32276
rect 10636 32444 10676 32453
rect 10444 32024 10484 32236
rect 10444 30260 10484 31984
rect 10444 30211 10484 30220
rect 10540 32108 10580 32117
rect 10540 30680 10580 32068
rect 10540 30176 10580 30640
rect 10636 30344 10676 32404
rect 10636 30295 10676 30304
rect 10540 30127 10580 30136
rect 10732 30176 10772 34168
rect 10828 32948 10868 35848
rect 10828 32696 10868 32908
rect 10828 32647 10868 32656
rect 10924 32024 10964 45004
rect 11020 44456 11060 46600
rect 11116 46472 11156 46481
rect 11116 45968 11156 46432
rect 11308 46472 11348 46481
rect 11116 45919 11156 45928
rect 11212 46388 11252 46397
rect 11212 44960 11252 46348
rect 11212 44911 11252 44920
rect 11020 44407 11060 44416
rect 11116 44288 11156 44297
rect 11116 44153 11156 44248
rect 11308 42944 11348 46432
rect 11980 45884 12020 48304
rect 11980 45835 12020 45844
rect 12364 46304 12404 46313
rect 11500 45800 11540 45809
rect 11500 45665 11540 45760
rect 11788 45800 11828 45809
rect 11692 45632 11732 45641
rect 11500 44960 11540 44969
rect 11500 44825 11540 44920
rect 11500 44288 11540 44297
rect 11500 43700 11540 44248
rect 11500 43651 11540 43660
rect 11308 42895 11348 42904
rect 11500 43448 11540 43457
rect 11020 42776 11060 42785
rect 11020 41852 11060 42736
rect 11020 41803 11060 41812
rect 11500 40340 11540 43408
rect 11692 42944 11732 45592
rect 11692 42895 11732 42904
rect 11596 42776 11636 42785
rect 11596 42641 11636 42736
rect 11500 40291 11540 40300
rect 11500 39668 11540 39677
rect 11116 38912 11156 38921
rect 11116 38777 11156 38872
rect 11020 38240 11060 38249
rect 11020 37652 11060 38200
rect 11020 37603 11060 37612
rect 11116 37988 11156 37997
rect 11020 37148 11060 37157
rect 11020 35972 11060 37108
rect 11020 32780 11060 35932
rect 11020 32731 11060 32740
rect 10828 31984 10964 32024
rect 10828 30932 10868 31984
rect 10828 30883 10868 30892
rect 10924 31856 10964 31865
rect 10828 30764 10868 30773
rect 10828 30260 10868 30724
rect 10924 30680 10964 31816
rect 10924 30631 10964 30640
rect 11020 31184 11060 31193
rect 10828 30211 10868 30220
rect 10732 30127 10772 30136
rect 10924 30176 10964 30185
rect 10924 30092 10964 30136
rect 10828 30052 10964 30092
rect 10444 30008 10484 30017
rect 10444 29000 10484 29968
rect 10732 30008 10772 30017
rect 10444 28951 10484 28960
rect 10540 29924 10580 29933
rect 10540 28832 10580 29884
rect 10636 29672 10676 29681
rect 10636 29336 10676 29632
rect 10636 29084 10676 29296
rect 10636 29000 10676 29044
rect 10636 28920 10676 28960
rect 10348 27439 10388 27448
rect 10444 28792 10580 28832
rect 10348 27320 10388 27329
rect 10348 26396 10388 27280
rect 10348 26347 10388 26356
rect 10292 25852 10388 25892
rect 10252 25843 10292 25852
rect 10252 24380 10292 24389
rect 10252 23876 10292 24340
rect 10348 23960 10388 25852
rect 10348 23911 10388 23920
rect 10252 23827 10292 23836
rect 10444 23708 10484 28792
rect 10540 28664 10580 28673
rect 10540 28412 10580 28624
rect 10540 28363 10580 28372
rect 10732 27572 10772 29968
rect 10828 29840 10868 30052
rect 10828 29791 10868 29800
rect 10924 29924 10964 29933
rect 10924 29420 10964 29884
rect 10924 29371 10964 29380
rect 10828 29168 10868 29177
rect 10868 29128 10964 29168
rect 10828 29119 10868 29128
rect 10636 27532 10772 27572
rect 10828 29000 10868 29009
rect 10156 22231 10196 22240
rect 10252 23668 10484 23708
rect 10540 27404 10580 27413
rect 10060 21356 10100 21365
rect 10060 20852 10100 21316
rect 10060 20803 10100 20812
rect 10060 20684 10100 20693
rect 10060 20096 10100 20644
rect 10060 20047 10100 20056
rect 10156 20600 10196 20609
rect 10156 20012 10196 20560
rect 10156 19963 10196 19972
rect 9964 18367 10004 18376
rect 10060 19928 10100 19937
rect 10060 18584 10100 19888
rect 9964 17996 10004 18005
rect 9964 17861 10004 17956
rect 9772 16276 9908 16316
rect 9964 17660 10004 17669
rect 9964 16316 10004 17620
rect 10060 17072 10100 18544
rect 10060 17023 10100 17032
rect 10156 19844 10196 19853
rect 10156 18416 10196 19804
rect 9772 14636 9812 16276
rect 9964 16267 10004 16276
rect 10156 16904 10196 18376
rect 9772 14587 9812 14596
rect 9868 16148 9908 16157
rect 9676 14503 9716 14512
rect 9772 14468 9812 14477
rect 9676 14384 9716 14393
rect 9676 14048 9716 14344
rect 9676 13999 9716 14008
rect 9772 13460 9812 14428
rect 9772 13411 9812 13420
rect 9580 12940 9716 12980
rect 9388 9631 9428 9640
rect 9484 12788 9524 12797
rect 9292 9547 9332 9556
rect 9100 8875 9140 8884
rect 9388 9512 9428 9521
rect 9292 8672 9332 8681
rect 9004 8044 9236 8084
rect 9004 7916 9044 7925
rect 9004 7076 9044 7876
rect 9004 7027 9044 7036
rect 9100 7832 9140 7841
rect 9100 5732 9140 7792
rect 9004 5692 9100 5732
rect 9004 5228 9044 5692
rect 9100 5683 9140 5692
rect 9004 4976 9044 5188
rect 9004 4927 9044 4936
rect 9100 4892 9140 4901
rect 9004 4220 9044 4229
rect 8908 4180 9004 4220
rect 8620 3380 8660 4012
rect 9004 3548 9044 4180
rect 9100 3632 9140 4852
rect 9100 3583 9140 3592
rect 9004 3499 9044 3508
rect 9196 3548 9236 8044
rect 9292 6404 9332 8632
rect 9388 8168 9428 9472
rect 9388 8119 9428 8128
rect 9484 7832 9524 12748
rect 9580 12704 9620 12713
rect 9580 12569 9620 12664
rect 9580 9428 9620 9437
rect 9580 8756 9620 9388
rect 9580 8707 9620 8716
rect 9484 7783 9524 7792
rect 9292 6355 9332 6364
rect 9484 6572 9524 6581
rect 9484 4976 9524 6532
rect 9580 6236 9620 6245
rect 9580 5732 9620 6196
rect 9580 5683 9620 5692
rect 9676 5564 9716 12940
rect 9772 12872 9812 12881
rect 9772 12620 9812 12832
rect 9772 11780 9812 12580
rect 9868 12536 9908 16108
rect 10060 15896 10100 15905
rect 9964 15812 10004 15821
rect 9964 12788 10004 15772
rect 10060 14048 10100 15856
rect 10060 13999 10100 14008
rect 10156 13460 10196 16864
rect 10252 15812 10292 23668
rect 10540 23456 10580 27364
rect 10540 23407 10580 23416
rect 10348 23288 10388 23297
rect 10348 19256 10388 23248
rect 10444 23204 10484 23213
rect 10444 22532 10484 23164
rect 10444 22483 10484 22492
rect 10540 23120 10580 23129
rect 10348 19207 10388 19216
rect 10444 22112 10484 22121
rect 10444 19256 10484 22072
rect 10540 21608 10580 23080
rect 10636 22280 10676 27532
rect 10732 27404 10772 27413
rect 10732 25976 10772 27364
rect 10732 25927 10772 25936
rect 10828 25808 10868 28960
rect 10924 28244 10964 29128
rect 11020 29084 11060 31144
rect 11020 29035 11060 29044
rect 10924 26732 10964 28204
rect 11020 28916 11060 28925
rect 11020 26900 11060 28876
rect 11020 26851 11060 26860
rect 10924 26597 10964 26692
rect 10636 22231 10676 22240
rect 10732 25768 10868 25808
rect 10540 21559 10580 21568
rect 10636 21524 10676 21533
rect 10444 19207 10484 19216
rect 10540 20852 10580 20861
rect 10540 19256 10580 20812
rect 10348 18416 10388 18511
rect 10348 18367 10388 18376
rect 10252 15763 10292 15772
rect 10348 18248 10388 18257
rect 10348 17744 10388 18208
rect 10540 17996 10580 19216
rect 10636 18248 10676 21484
rect 10636 18199 10676 18208
rect 10580 17956 10676 17996
rect 10540 17947 10580 17956
rect 10348 15056 10388 17704
rect 10540 17744 10580 17753
rect 10156 13411 10196 13420
rect 10252 15016 10388 15056
rect 10444 16988 10484 16997
rect 10252 14384 10292 15016
rect 9964 12739 10004 12748
rect 10252 13376 10292 14344
rect 9868 12496 10004 12536
rect 9772 11731 9812 11740
rect 9868 12368 9908 12377
rect 9772 10940 9812 10949
rect 9772 9680 9812 10900
rect 9868 10436 9908 12328
rect 9868 10387 9908 10396
rect 9772 9631 9812 9640
rect 9676 5515 9716 5524
rect 9964 5144 10004 12496
rect 9964 5095 10004 5104
rect 10060 12452 10100 12461
rect 10060 11528 10100 12412
rect 10060 7916 10100 11488
rect 10156 12368 10196 12377
rect 10156 12032 10196 12328
rect 10156 11360 10196 11992
rect 10156 11311 10196 11320
rect 10252 11948 10292 13336
rect 10348 14888 10388 14897
rect 10348 13208 10388 14848
rect 10348 13159 10388 13168
rect 10252 11024 10292 11908
rect 10252 10268 10292 10984
rect 10348 11696 10388 11705
rect 10348 11108 10388 11656
rect 10348 10520 10388 11068
rect 10348 10471 10388 10480
rect 10252 9512 10292 10228
rect 10444 9596 10484 16948
rect 10540 16484 10580 17704
rect 10540 16435 10580 16444
rect 10636 16316 10676 17956
rect 10732 16904 10772 25768
rect 11116 25136 11156 37948
rect 11308 37400 11348 37409
rect 11212 37064 11252 37073
rect 11212 35888 11252 37024
rect 11308 36140 11348 37360
rect 11404 37232 11444 37241
rect 11404 37097 11444 37192
rect 11308 36091 11348 36100
rect 11404 36476 11444 36485
rect 11404 35972 11444 36436
rect 11404 35923 11444 35932
rect 11212 35839 11252 35848
rect 11404 35132 11444 35141
rect 11212 35048 11252 35057
rect 11212 33620 11252 35008
rect 11212 33571 11252 33580
rect 11308 33788 11348 33797
rect 11212 33452 11252 33461
rect 11212 32948 11252 33412
rect 11212 32899 11252 32908
rect 11116 25087 11156 25096
rect 11212 32780 11252 32789
rect 11212 24968 11252 32740
rect 11308 32192 11348 33748
rect 11404 33116 11444 35092
rect 11404 33067 11444 33076
rect 11404 32864 11444 32873
rect 11404 32729 11444 32824
rect 11308 32143 11348 32152
rect 11404 32612 11444 32621
rect 11404 32528 11444 32572
rect 11308 30596 11348 30605
rect 11308 30461 11348 30556
rect 11404 30344 11444 32488
rect 11500 31520 11540 39628
rect 11788 39416 11828 45760
rect 12172 45800 12212 45809
rect 11884 44960 11924 44969
rect 11884 44708 11924 44920
rect 11884 44659 11924 44668
rect 11884 44288 11924 44297
rect 11884 43364 11924 44248
rect 11884 43315 11924 43324
rect 11980 42776 12020 42785
rect 11980 41936 12020 42736
rect 11980 41887 12020 41896
rect 11788 39367 11828 39376
rect 11980 39500 12020 39509
rect 11596 38912 11636 38921
rect 11596 33872 11636 38872
rect 11884 38912 11924 38921
rect 11884 38777 11924 38872
rect 11788 38744 11828 38753
rect 11596 33823 11636 33832
rect 11692 38156 11732 38165
rect 11692 33368 11732 38116
rect 11788 37064 11828 38704
rect 11980 38408 12020 39460
rect 11980 38359 12020 38368
rect 12076 39164 12116 39173
rect 11884 38240 11924 38249
rect 11884 38105 11924 38200
rect 11980 38072 12020 38081
rect 11884 37400 11924 37409
rect 11980 37400 12020 38032
rect 12076 37736 12116 39124
rect 12076 37687 12116 37696
rect 11980 37360 12116 37400
rect 11884 37265 11924 37360
rect 11788 37015 11828 37024
rect 11980 37232 12020 37241
rect 11884 36560 11924 36569
rect 11884 35468 11924 36520
rect 11884 35419 11924 35428
rect 11980 34040 12020 37192
rect 12076 36056 12116 37360
rect 12076 36007 12116 36016
rect 11980 33991 12020 34000
rect 12076 35888 12116 35897
rect 11980 33872 12020 33881
rect 11500 31471 11540 31480
rect 11596 33328 11732 33368
rect 11788 33536 11828 33545
rect 11308 30304 11444 30344
rect 11500 31352 11540 31361
rect 11308 29588 11348 30304
rect 11308 29539 11348 29548
rect 11116 24928 11252 24968
rect 11308 29252 11348 29261
rect 11308 25388 11348 29212
rect 11404 28832 11444 28841
rect 11404 26900 11444 28792
rect 11500 27068 11540 31312
rect 11596 30848 11636 33328
rect 11692 33200 11732 33211
rect 11692 33116 11732 33160
rect 11692 33067 11732 33076
rect 11596 30799 11636 30808
rect 11692 32696 11732 32705
rect 11596 30680 11636 30689
rect 11596 28916 11636 30640
rect 11596 28867 11636 28876
rect 11596 28412 11636 28421
rect 11596 27740 11636 28372
rect 11596 27691 11636 27700
rect 11500 27019 11540 27028
rect 11596 27572 11636 27581
rect 11404 26860 11540 26900
rect 11404 26228 11444 26237
rect 11404 26093 11444 26188
rect 11020 23876 11060 23885
rect 10828 23624 10868 23633
rect 10828 23540 10868 23584
rect 10828 23489 10868 23500
rect 10828 23288 10868 23297
rect 10828 23204 10868 23248
rect 10828 23153 10868 23164
rect 11020 23036 11060 23836
rect 10924 22700 10964 22709
rect 10828 21356 10868 21365
rect 10828 20516 10868 21316
rect 10828 20467 10868 20476
rect 10828 20348 10868 20357
rect 10828 20012 10868 20308
rect 10828 17744 10868 19972
rect 10924 19844 10964 22660
rect 11020 22364 11060 22996
rect 11020 21524 11060 22324
rect 11020 21475 11060 21484
rect 10924 19795 10964 19804
rect 11020 21356 11060 21365
rect 10924 19088 10964 19097
rect 10924 18500 10964 19048
rect 10924 18451 10964 18460
rect 10828 17695 10868 17704
rect 10924 18248 10964 18257
rect 10924 17828 10964 18208
rect 10732 16855 10772 16864
rect 10828 17072 10868 17081
rect 10636 16267 10676 16276
rect 10732 16736 10772 16745
rect 10540 16232 10580 16241
rect 10540 15476 10580 16192
rect 10732 16148 10772 16696
rect 10540 15427 10580 15436
rect 10636 16108 10772 16148
rect 10540 14216 10580 14225
rect 10540 14081 10580 14176
rect 10444 9547 10484 9556
rect 10540 12536 10580 12545
rect 10540 11192 10580 12496
rect 10252 9463 10292 9472
rect 10540 8924 10580 11152
rect 10636 10772 10676 16108
rect 10732 15980 10772 15989
rect 10732 14720 10772 15940
rect 10732 14671 10772 14680
rect 10732 14552 10772 14561
rect 10732 14417 10772 14512
rect 10732 14300 10772 14309
rect 10732 11108 10772 14260
rect 10732 11059 10772 11068
rect 10636 10723 10676 10732
rect 10540 8875 10580 8884
rect 9484 4927 9524 4936
rect 9964 4976 10004 4985
rect 9964 4841 10004 4936
rect 9196 3499 9236 3508
rect 9676 3968 9716 3977
rect 9676 3464 9716 3928
rect 9964 3968 10004 3977
rect 9772 3800 9812 3809
rect 9964 3800 10004 3928
rect 9812 3760 10004 3800
rect 9772 3751 9812 3760
rect 10060 3632 10100 7876
rect 10828 7160 10868 17032
rect 10924 16988 10964 17788
rect 10924 16939 10964 16948
rect 10924 16820 10964 16829
rect 10924 15980 10964 16780
rect 10924 15931 10964 15940
rect 10924 15476 10964 15485
rect 10924 14804 10964 15436
rect 10924 13964 10964 14764
rect 11020 14384 11060 21316
rect 11020 14335 11060 14344
rect 11116 17744 11156 24928
rect 11212 24800 11252 24809
rect 11212 23708 11252 24760
rect 11308 24548 11348 25348
rect 11500 24800 11540 26860
rect 11500 24751 11540 24760
rect 11308 23876 11348 24508
rect 11596 24548 11636 27532
rect 11692 27404 11732 32656
rect 11788 31352 11828 33496
rect 11980 33200 12020 33832
rect 11884 33160 12020 33200
rect 11884 31352 11924 33160
rect 11980 32696 12020 32705
rect 12076 32696 12116 35848
rect 12020 32656 12116 32696
rect 11980 32647 12020 32656
rect 11884 31312 12116 31352
rect 11788 31303 11828 31312
rect 11980 31184 12020 31193
rect 11884 30428 11924 30437
rect 11692 27355 11732 27364
rect 11788 28832 11828 28841
rect 11692 27236 11732 27245
rect 11692 26816 11732 27196
rect 11692 26767 11732 26776
rect 11788 26648 11828 28792
rect 11884 28664 11924 30388
rect 11980 29000 12020 31144
rect 11980 28951 12020 28960
rect 11884 28615 11924 28624
rect 11980 28160 12020 28169
rect 11884 27824 11924 27833
rect 11884 27236 11924 27784
rect 11884 27187 11924 27196
rect 11980 26900 12020 28120
rect 11980 26851 12020 26860
rect 11596 24499 11636 24508
rect 11692 26608 11828 26648
rect 11884 26816 11924 26825
rect 11500 23960 11540 23969
rect 11348 23836 11444 23876
rect 11308 23827 11348 23836
rect 11212 23668 11348 23708
rect 11212 23456 11252 23465
rect 11212 23036 11252 23416
rect 11212 19340 11252 22996
rect 11308 22364 11348 23668
rect 11308 20852 11348 22324
rect 11308 20803 11348 20812
rect 11212 19291 11252 19300
rect 11308 20432 11348 20441
rect 11116 14300 11156 17704
rect 11212 19172 11252 19181
rect 11212 16736 11252 19132
rect 11308 16820 11348 20392
rect 11308 16771 11348 16780
rect 11212 16687 11252 16696
rect 11404 16400 11444 23836
rect 11500 22532 11540 23920
rect 11500 22483 11540 22492
rect 11596 22952 11636 22961
rect 11500 21944 11540 21953
rect 11500 21356 11540 21904
rect 11596 21692 11636 22912
rect 11596 21643 11636 21652
rect 11500 21307 11540 21316
rect 11500 20936 11540 20945
rect 11500 20096 11540 20896
rect 11500 18416 11540 20056
rect 11596 20264 11636 20273
rect 11596 19508 11636 20224
rect 11596 19459 11636 19468
rect 11692 18836 11732 26608
rect 11692 18787 11732 18796
rect 11788 26480 11828 26489
rect 11500 18376 11636 18416
rect 11500 18248 11540 18257
rect 11500 17072 11540 18208
rect 11596 18164 11636 18376
rect 11596 18124 11732 18164
rect 11500 17023 11540 17032
rect 11596 17996 11636 18005
rect 11308 16360 11444 16400
rect 11500 16904 11540 16913
rect 11212 16316 11252 16325
rect 11212 15476 11252 16276
rect 11212 15427 11252 15436
rect 11116 14251 11156 14260
rect 10924 13915 10964 13924
rect 11308 11696 11348 16360
rect 11404 15980 11444 15989
rect 11404 13964 11444 15940
rect 11404 13915 11444 13924
rect 11404 13040 11444 13049
rect 11404 12452 11444 13000
rect 11500 12620 11540 16864
rect 11596 16232 11636 17956
rect 11692 17828 11732 18124
rect 11692 17779 11732 17788
rect 11692 17492 11732 17501
rect 11692 17357 11732 17452
rect 11788 17072 11828 26440
rect 11884 26312 11924 26776
rect 12076 26732 12116 31312
rect 12172 29252 12212 45760
rect 12268 45548 12308 45557
rect 12268 44120 12308 45508
rect 12364 45128 12404 46264
rect 12556 46052 12596 48304
rect 12556 46003 12596 46012
rect 12748 46472 12788 46481
rect 12364 45079 12404 45088
rect 12364 44960 12404 44969
rect 12364 44876 12404 44920
rect 12364 44825 12404 44836
rect 12268 44071 12308 44080
rect 12364 43280 12404 43289
rect 12364 42440 12404 43240
rect 12364 42391 12404 42400
rect 12460 41264 12500 41273
rect 12364 40256 12404 40265
rect 12268 39416 12308 39425
rect 12268 34880 12308 39376
rect 12364 39164 12404 40216
rect 12364 39115 12404 39124
rect 12364 38996 12404 39007
rect 12364 38912 12404 38956
rect 12364 38863 12404 38872
rect 12364 37988 12404 37997
rect 12364 35048 12404 37948
rect 12364 34999 12404 35008
rect 12268 34840 12404 34880
rect 12268 34376 12308 34385
rect 12268 34241 12308 34336
rect 12268 33704 12308 33799
rect 12268 33655 12308 33664
rect 12268 33452 12308 33461
rect 12268 32864 12308 33412
rect 12364 33032 12404 34840
rect 12460 34124 12500 41224
rect 12556 40424 12596 40433
rect 12556 36224 12596 40384
rect 12556 36175 12596 36184
rect 12652 38072 12692 38081
rect 12556 35720 12596 35729
rect 12556 34376 12596 35680
rect 12556 34327 12596 34336
rect 12652 34376 12692 38032
rect 12748 36560 12788 46432
rect 13132 46304 13172 46313
rect 13036 45548 13076 45557
rect 13036 43784 13076 45508
rect 13132 44456 13172 46264
rect 13132 44407 13172 44416
rect 13036 43735 13076 43744
rect 13132 44036 13172 44045
rect 13036 43280 13076 43289
rect 13036 42104 13076 43240
rect 13132 42776 13172 43996
rect 13132 42727 13172 42736
rect 13036 42055 13076 42064
rect 13132 42524 13172 42533
rect 12940 41768 12980 41777
rect 12844 40928 12884 40937
rect 12844 40424 12884 40888
rect 12940 40760 12980 41728
rect 13132 41768 13172 42484
rect 13132 41719 13172 41728
rect 13612 41600 13652 41609
rect 13612 41432 13652 41560
rect 13612 41383 13652 41392
rect 12940 40711 12980 40720
rect 13132 41012 13172 41021
rect 12844 40375 12884 40384
rect 13132 39752 13172 40972
rect 13132 39703 13172 39712
rect 13228 40508 13268 40517
rect 13132 39500 13172 39509
rect 12940 38996 12980 39005
rect 12748 36511 12788 36520
rect 12844 37988 12884 37997
rect 12748 36392 12788 36401
rect 12748 35720 12788 36352
rect 12748 35671 12788 35680
rect 12652 34327 12692 34336
rect 12748 34292 12788 34301
rect 12460 34084 12692 34124
rect 12556 33872 12596 33881
rect 12556 33140 12596 33832
rect 12364 32983 12404 32992
rect 12460 33100 12596 33140
rect 12268 32824 12404 32864
rect 12268 32696 12308 32705
rect 12268 30344 12308 32656
rect 12364 31016 12404 32824
rect 12460 32024 12500 33100
rect 12460 31975 12500 31984
rect 12556 32696 12596 32705
rect 12364 30967 12404 30976
rect 12460 31520 12500 31529
rect 12268 30295 12308 30304
rect 12364 30680 12404 30689
rect 12364 29840 12404 30640
rect 12364 29791 12404 29800
rect 12172 29203 12212 29212
rect 11884 26263 11924 26272
rect 11980 26692 12116 26732
rect 12172 29084 12212 29093
rect 11884 25976 11924 25985
rect 11884 20768 11924 25936
rect 11980 24632 12020 26692
rect 12076 26060 12116 26069
rect 12076 24800 12116 26020
rect 12076 24751 12116 24760
rect 12172 24632 12212 29044
rect 12364 28916 12404 28925
rect 11980 24583 12020 24592
rect 12076 24592 12212 24632
rect 12268 27572 12308 27581
rect 12076 22448 12116 24592
rect 12076 22399 12116 22408
rect 12172 23624 12212 23633
rect 11884 20719 11924 20728
rect 11980 21524 12020 21533
rect 11884 19928 11924 19937
rect 11884 19844 11924 19888
rect 11884 19793 11924 19804
rect 11884 18668 11924 18679
rect 11884 18584 11924 18628
rect 11884 18535 11924 18544
rect 11980 17492 12020 21484
rect 12172 21020 12212 23584
rect 12268 21524 12308 27532
rect 12364 26984 12404 28876
rect 12460 27488 12500 31480
rect 12556 30008 12596 32656
rect 12556 29959 12596 29968
rect 12652 28076 12692 34084
rect 12748 31688 12788 34252
rect 12844 33704 12884 37948
rect 12940 36392 12980 38956
rect 12940 36343 12980 36352
rect 13036 38912 13076 38921
rect 12844 33655 12884 33664
rect 12940 36224 12980 36233
rect 12748 31639 12788 31648
rect 12844 33536 12884 33545
rect 12460 27439 12500 27448
rect 12556 28036 12692 28076
rect 12748 30512 12788 30521
rect 12364 26935 12404 26944
rect 12268 21475 12308 21484
rect 12364 25388 12404 25397
rect 12172 20971 12212 20980
rect 12268 21356 12308 21365
rect 12076 20600 12116 20609
rect 12076 18500 12116 20560
rect 12172 19844 12212 19853
rect 12172 18668 12212 19804
rect 12172 18619 12212 18628
rect 12076 18451 12116 18460
rect 12268 18332 12308 21316
rect 12268 18283 12308 18292
rect 12076 18248 12116 18257
rect 12076 18113 12116 18208
rect 12364 18164 12404 25348
rect 12460 24632 12500 24641
rect 12460 24044 12500 24592
rect 12460 23995 12500 24004
rect 12556 21356 12596 28036
rect 12748 27656 12788 30472
rect 12844 28076 12884 33496
rect 12844 28027 12884 28036
rect 12748 27607 12788 27616
rect 12844 27908 12884 27917
rect 12748 27488 12788 27497
rect 12556 21307 12596 21316
rect 12652 26228 12692 26237
rect 12556 21188 12596 21197
rect 12460 19928 12500 19937
rect 12460 19793 12500 19888
rect 12172 18124 12404 18164
rect 12460 19088 12500 19097
rect 11884 17452 12020 17492
rect 12076 17828 12116 17837
rect 11884 17156 11924 17452
rect 11884 17107 11924 17116
rect 11980 17324 12020 17333
rect 11788 17023 11828 17032
rect 11884 16988 11924 16997
rect 11788 16904 11828 16913
rect 11596 16183 11636 16192
rect 11692 16820 11732 16829
rect 11596 16064 11636 16073
rect 11596 14048 11636 16024
rect 11692 14720 11732 16780
rect 11692 14671 11732 14680
rect 11788 14048 11828 16864
rect 11884 14216 11924 16948
rect 11980 16484 12020 17284
rect 11980 16435 12020 16444
rect 11884 14167 11924 14176
rect 11980 16316 12020 16325
rect 11788 14008 11924 14048
rect 11596 13292 11636 14008
rect 11596 13243 11636 13252
rect 11788 13880 11828 13889
rect 11500 12571 11540 12580
rect 11692 12788 11732 12797
rect 11404 12403 11444 12412
rect 11596 12284 11636 12293
rect 11500 11948 11540 12043
rect 11500 11899 11540 11908
rect 11308 10268 11348 11656
rect 11500 11780 11540 11789
rect 11404 11612 11444 11621
rect 11404 11477 11444 11572
rect 11500 11192 11540 11740
rect 11500 11143 11540 11152
rect 11308 10219 11348 10228
rect 11308 9848 11348 9857
rect 11308 8672 11348 9808
rect 11404 9764 11444 9773
rect 11404 8924 11444 9724
rect 11596 9512 11636 12244
rect 11596 9463 11636 9472
rect 11692 9428 11732 12748
rect 11788 11276 11828 13840
rect 11788 11227 11828 11236
rect 11884 10688 11924 14008
rect 11980 12704 12020 16276
rect 12076 15728 12116 17788
rect 12172 17240 12212 18124
rect 12364 17996 12404 18005
rect 12172 17191 12212 17200
rect 12268 17912 12308 17921
rect 12076 15679 12116 15688
rect 12172 17072 12212 17081
rect 12172 15560 12212 17032
rect 12076 15520 12212 15560
rect 12076 14048 12116 15520
rect 12172 15140 12212 15149
rect 12172 14132 12212 15100
rect 12268 14720 12308 17872
rect 12268 14671 12308 14680
rect 12172 14092 12308 14132
rect 12076 14008 12212 14048
rect 11980 12655 12020 12664
rect 12076 13124 12116 13133
rect 12076 11024 12116 13084
rect 12172 12704 12212 14008
rect 12172 12655 12212 12664
rect 12268 11696 12308 14092
rect 12364 11948 12404 17956
rect 12460 17744 12500 19048
rect 12556 18668 12596 21148
rect 12556 18619 12596 18628
rect 12652 17996 12692 26188
rect 12748 19088 12788 27448
rect 12844 25220 12884 27868
rect 12844 25171 12884 25180
rect 12844 24296 12884 24305
rect 12844 21020 12884 24256
rect 12844 20971 12884 20980
rect 12748 19039 12788 19048
rect 12844 19592 12884 19601
rect 12652 17947 12692 17956
rect 12748 18920 12788 18929
rect 12460 17704 12692 17744
rect 12460 17576 12500 17585
rect 12460 14048 12500 17536
rect 12460 13999 12500 14008
rect 12556 16568 12596 16577
rect 12364 11899 12404 11908
rect 12460 12872 12500 12881
rect 12268 11647 12308 11656
rect 12076 10975 12116 10984
rect 12268 11192 12308 11201
rect 11884 10648 12020 10688
rect 11884 10520 11924 10529
rect 11788 9680 11828 9689
rect 11788 9545 11828 9640
rect 11692 9388 11828 9428
rect 11404 8875 11444 8884
rect 11692 9176 11732 9185
rect 11308 8623 11348 8632
rect 11692 8000 11732 9136
rect 11692 7951 11732 7960
rect 10828 7111 10868 7120
rect 11308 7160 11348 7169
rect 11308 6404 11348 7120
rect 11308 6355 11348 6364
rect 11692 6488 11732 6497
rect 11692 5816 11732 6448
rect 11692 5767 11732 5776
rect 11788 5732 11828 9388
rect 11884 8672 11924 10480
rect 11884 8623 11924 8632
rect 11980 8084 12020 10648
rect 12172 8672 12212 8681
rect 12172 8504 12212 8632
rect 12268 8672 12308 11152
rect 12460 10184 12500 12832
rect 12556 12620 12596 16528
rect 12652 13880 12692 17704
rect 12748 16484 12788 18880
rect 12844 17240 12884 19552
rect 12940 18584 12980 36184
rect 13036 34712 13076 38872
rect 13132 36728 13172 39460
rect 13132 36679 13172 36688
rect 13036 34663 13076 34672
rect 13228 34460 13268 40468
rect 13420 40340 13460 40349
rect 13324 39584 13364 39593
rect 13324 37400 13364 39544
rect 13420 38072 13460 40300
rect 13420 38023 13460 38032
rect 13516 39668 13556 39677
rect 13324 37351 13364 37360
rect 13420 37316 13460 37325
rect 13132 34420 13268 34460
rect 13324 36476 13364 36485
rect 13132 33536 13172 34420
rect 13132 33487 13172 33496
rect 13228 34208 13268 34217
rect 13036 33452 13076 33461
rect 13036 30680 13076 33412
rect 13036 30631 13076 30640
rect 13132 31940 13172 31949
rect 13036 30428 13076 30437
rect 13036 27320 13076 30388
rect 13132 29084 13172 31900
rect 13228 31352 13268 34168
rect 13324 32360 13364 36436
rect 13420 33368 13460 37276
rect 13420 33319 13460 33328
rect 13324 32311 13364 32320
rect 13420 33032 13460 33041
rect 13228 31303 13268 31312
rect 13324 31268 13364 31277
rect 13132 29035 13172 29044
rect 13228 31184 13268 31193
rect 13036 27271 13076 27280
rect 13132 28916 13172 28925
rect 13132 26648 13172 28876
rect 13228 27992 13268 31144
rect 13324 28328 13364 31228
rect 13324 28279 13364 28288
rect 13420 28160 13460 32992
rect 13228 27943 13268 27952
rect 13324 28120 13460 28160
rect 13324 27152 13364 28120
rect 13324 27103 13364 27112
rect 13420 27992 13460 28001
rect 13324 26900 13364 26909
rect 13132 26599 13172 26608
rect 13228 26732 13268 26741
rect 13036 26312 13076 26321
rect 13036 24800 13076 26272
rect 13132 25976 13172 25985
rect 13132 25556 13172 25936
rect 13132 25507 13172 25516
rect 13228 25388 13268 26692
rect 13036 24751 13076 24760
rect 13132 25348 13268 25388
rect 13036 24632 13076 24641
rect 13036 18668 13076 24592
rect 13036 18619 13076 18628
rect 12940 18535 12980 18544
rect 13132 18416 13172 25348
rect 13228 25220 13268 25229
rect 13228 23288 13268 25180
rect 13324 23456 13364 26860
rect 13324 23407 13364 23416
rect 13228 23248 13364 23288
rect 12844 17191 12884 17200
rect 12940 18376 13172 18416
rect 13228 23120 13268 23129
rect 12940 17072 12980 18376
rect 13132 18248 13172 18257
rect 12748 16435 12788 16444
rect 12844 17032 12980 17072
rect 13036 17660 13076 17669
rect 12844 16400 12884 17032
rect 12844 16351 12884 16360
rect 12940 16904 12980 16913
rect 12844 16232 12884 16241
rect 12652 13831 12692 13840
rect 12748 14216 12788 14225
rect 12556 12571 12596 12580
rect 12748 11780 12788 14176
rect 12748 11731 12788 11740
rect 12844 11696 12884 16192
rect 12940 12536 12980 16864
rect 13036 14888 13076 17620
rect 13036 14839 13076 14848
rect 13132 14720 13172 18208
rect 13132 14671 13172 14680
rect 12940 12487 12980 12496
rect 13132 14552 13172 14561
rect 12844 11647 12884 11656
rect 13036 12200 13076 12209
rect 12460 10135 12500 10144
rect 12844 10184 12884 10193
rect 12268 8623 12308 8632
rect 12556 9428 12596 9437
rect 12172 8455 12212 8464
rect 11980 8035 12020 8044
rect 12076 8168 12116 8177
rect 12076 7160 12116 8128
rect 12268 8000 12308 8009
rect 12268 7865 12308 7960
rect 12076 7111 12116 7120
rect 12460 7496 12500 7505
rect 12460 6488 12500 7456
rect 12556 7160 12596 9388
rect 12844 8084 12884 10144
rect 13036 9596 13076 12160
rect 13132 11024 13172 14512
rect 13132 10975 13172 10984
rect 13036 9547 13076 9556
rect 13132 10856 13172 10865
rect 12844 8035 12884 8044
rect 13132 8000 13172 10816
rect 13132 7951 13172 7960
rect 12556 7111 12596 7120
rect 12460 6439 12500 6448
rect 11788 5683 11828 5692
rect 12460 6152 12500 6161
rect 10348 5648 10388 5657
rect 10348 5513 10388 5608
rect 12460 5648 12500 6112
rect 12460 5599 12500 5608
rect 12460 4472 12500 4481
rect 12460 4136 12500 4432
rect 12460 4087 12500 4096
rect 12556 4304 12596 4313
rect 10060 3583 10100 3592
rect 9676 3415 9716 3424
rect 8620 3331 8660 3340
rect 9100 1028 9140 1037
rect 9100 80 9140 988
rect 9676 1028 9716 1037
rect 9676 80 9716 988
rect 10252 1028 10292 1037
rect 10252 80 10292 988
rect 10828 1028 10868 1037
rect 10828 80 10868 988
rect 11404 1028 11444 1037
rect 11404 80 11444 988
rect 11980 692 12020 701
rect 11980 80 12020 652
rect 12556 80 12596 4264
rect 12652 4052 12692 4061
rect 12652 3464 12692 4012
rect 12652 3415 12692 3424
rect 13228 2792 13268 23080
rect 13324 20096 13364 23248
rect 13324 20047 13364 20056
rect 13324 18668 13364 18677
rect 13324 18248 13364 18628
rect 13420 18416 13460 27952
rect 13516 23540 13556 39628
rect 13612 38912 13652 38921
rect 13612 38744 13652 38872
rect 13612 38695 13652 38704
rect 13612 37232 13652 37241
rect 13612 33032 13652 37192
rect 13612 32983 13652 32992
rect 13516 23491 13556 23500
rect 13612 29252 13652 29261
rect 13420 18367 13460 18376
rect 13516 23372 13556 23381
rect 13324 18208 13460 18248
rect 13324 17240 13364 17249
rect 13324 13292 13364 17200
rect 13324 13243 13364 13252
rect 13324 12536 13364 12545
rect 13324 10268 13364 12496
rect 13420 11696 13460 18208
rect 13420 11647 13460 11656
rect 13324 10219 13364 10228
rect 13420 11528 13460 11537
rect 13420 8672 13460 11488
rect 13516 8924 13556 23332
rect 13612 20180 13652 29212
rect 13612 20131 13652 20140
rect 13612 18584 13652 18593
rect 13612 15056 13652 18544
rect 13612 15007 13652 15016
rect 13516 8875 13556 8884
rect 13612 14888 13652 14897
rect 13420 8623 13460 8632
rect 13516 2876 13556 2885
rect 13612 2876 13652 14848
rect 13556 2836 13652 2876
rect 13516 2827 13556 2836
rect 13228 2743 13268 2752
rect 3956 64 3976 80
rect 3896 0 3976 64
rect 4472 0 4552 80
rect 5048 0 5128 80
rect 5624 0 5704 80
rect 6200 0 6280 80
rect 6776 0 6856 80
rect 7352 0 7432 80
rect 7928 0 8008 80
rect 8504 0 8584 80
rect 9080 0 9160 80
rect 9656 0 9736 80
rect 10232 0 10312 80
rect 10808 0 10888 80
rect 11384 0 11464 80
rect 11960 0 12040 80
rect 12536 0 12616 80
<< via3 >>
rect 4928 46852 4968 46892
rect 5010 46852 5050 46892
rect 5092 46852 5132 46892
rect 5174 46852 5214 46892
rect 5256 46852 5296 46892
rect 1900 46432 1940 46472
rect 1420 10984 1460 11024
rect 1420 7960 1460 8000
rect 1420 7120 1460 7160
rect 1996 30136 2036 30176
rect 3688 46096 3728 46136
rect 3770 46096 3810 46136
rect 3852 46096 3892 46136
rect 3934 46096 3974 46136
rect 4016 46096 4056 46136
rect 2668 30808 2708 30848
rect 2284 25096 2324 25136
rect 1612 15940 1652 15980
rect 1612 8968 1652 9008
rect 1996 15940 2036 15980
rect 2284 22408 2324 22448
rect 2572 22408 2612 22448
rect 2668 22996 2708 23036
rect 2572 22240 2612 22280
rect 2668 20224 2708 20264
rect 2668 15940 2708 15980
rect 2572 15184 2612 15224
rect 2476 12916 2516 12956
rect 2668 13000 2708 13040
rect 2860 32572 2900 32612
rect 3688 44584 3728 44624
rect 3770 44584 3810 44624
rect 3852 44584 3892 44624
rect 3934 44584 3974 44624
rect 4016 44584 4056 44624
rect 3688 43072 3728 43112
rect 3770 43072 3810 43112
rect 3852 43072 3892 43112
rect 3934 43072 3974 43112
rect 4016 43072 4056 43112
rect 3688 41560 3728 41600
rect 3770 41560 3810 41600
rect 3852 41560 3892 41600
rect 3934 41560 3974 41600
rect 4016 41560 4056 41600
rect 3436 40300 3476 40340
rect 3688 40048 3728 40088
rect 3770 40048 3810 40088
rect 3852 40048 3892 40088
rect 3934 40048 3974 40088
rect 4016 40048 4056 40088
rect 3688 38536 3728 38576
rect 3770 38536 3810 38576
rect 3852 38536 3892 38576
rect 3934 38536 3974 38576
rect 4016 38536 4056 38576
rect 3688 37024 3728 37064
rect 3770 37024 3810 37064
rect 3852 37024 3892 37064
rect 3934 37024 3974 37064
rect 4016 37024 4056 37064
rect 3148 32908 3188 32948
rect 3688 35512 3728 35552
rect 3770 35512 3810 35552
rect 3852 35512 3892 35552
rect 3934 35512 3974 35552
rect 4016 35512 4056 35552
rect 3688 34000 3728 34040
rect 3770 34000 3810 34040
rect 3852 34000 3892 34040
rect 3934 34000 3974 34040
rect 4016 34000 4056 34040
rect 3436 32908 3476 32948
rect 3148 29212 3188 29252
rect 2860 22072 2900 22112
rect 3052 23164 3092 23204
rect 3148 22240 3188 22280
rect 3148 20224 3188 20264
rect 2956 17536 2996 17576
rect 3052 20140 3092 20180
rect 2956 17368 2996 17408
rect 2860 15016 2900 15056
rect 3148 17536 3188 17576
rect 3436 25516 3476 25556
rect 3688 32488 3728 32528
rect 3770 32488 3810 32528
rect 3852 32488 3892 32528
rect 3934 32488 3974 32528
rect 4016 32488 4056 32528
rect 4012 31900 4052 31940
rect 3688 30976 3728 31016
rect 3770 30976 3810 31016
rect 3852 30976 3892 31016
rect 3934 30976 3974 31016
rect 4016 30976 4056 31016
rect 3820 30808 3860 30848
rect 3820 29716 3860 29756
rect 4012 30724 4052 30764
rect 4108 30472 4148 30512
rect 4588 40300 4628 40340
rect 4928 45340 4968 45380
rect 5010 45340 5050 45380
rect 5092 45340 5132 45380
rect 5174 45340 5214 45380
rect 5256 45340 5296 45380
rect 5452 44920 5492 44960
rect 4928 43828 4968 43868
rect 5010 43828 5050 43868
rect 5092 43828 5132 43868
rect 5174 43828 5214 43868
rect 5256 43828 5296 43868
rect 4928 42316 4968 42356
rect 5010 42316 5050 42356
rect 5092 42316 5132 42356
rect 5174 42316 5214 42356
rect 5256 42316 5296 42356
rect 4928 40804 4968 40844
rect 5010 40804 5050 40844
rect 5092 40804 5132 40844
rect 5174 40804 5214 40844
rect 5256 40804 5296 40844
rect 4928 39292 4968 39332
rect 5010 39292 5050 39332
rect 5092 39292 5132 39332
rect 5174 39292 5214 39332
rect 5256 39292 5296 39332
rect 4684 38284 4724 38324
rect 4492 37948 4532 37988
rect 4300 32236 4340 32276
rect 4396 31984 4436 32024
rect 4300 30220 4340 30260
rect 5356 37948 5396 37988
rect 5452 38284 5492 38324
rect 4928 37780 4968 37820
rect 5010 37780 5050 37820
rect 5092 37780 5132 37820
rect 5174 37780 5214 37820
rect 5256 37780 5296 37820
rect 4928 36268 4968 36308
rect 5010 36268 5050 36308
rect 5092 36268 5132 36308
rect 5174 36268 5214 36308
rect 5256 36268 5296 36308
rect 4928 34756 4968 34796
rect 5010 34756 5050 34796
rect 5092 34756 5132 34796
rect 5174 34756 5214 34796
rect 5256 34756 5296 34796
rect 4492 30220 4532 30260
rect 4396 30136 4436 30176
rect 4928 33244 4968 33284
rect 5010 33244 5050 33284
rect 5092 33244 5132 33284
rect 5174 33244 5214 33284
rect 5256 33244 5296 33284
rect 4684 30220 4724 30260
rect 5164 31900 5204 31940
rect 4928 31732 4968 31772
rect 5010 31732 5050 31772
rect 5092 31732 5132 31772
rect 5174 31732 5214 31772
rect 5256 31732 5296 31772
rect 4928 30220 4968 30260
rect 5010 30220 5050 30260
rect 5092 30220 5132 30260
rect 5174 30220 5214 30260
rect 5256 30220 5296 30260
rect 4588 30136 4628 30176
rect 3724 29632 3764 29672
rect 3688 29464 3728 29504
rect 3770 29464 3810 29504
rect 3852 29464 3892 29504
rect 3934 29464 3974 29504
rect 4016 29464 4056 29504
rect 3688 27952 3728 27992
rect 3770 27952 3810 27992
rect 3852 27952 3892 27992
rect 3934 27952 3974 27992
rect 4016 27952 4056 27992
rect 3688 26440 3728 26480
rect 3770 26440 3810 26480
rect 3852 26440 3892 26480
rect 3934 26440 3974 26480
rect 4016 26440 4056 26480
rect 4108 26020 4148 26060
rect 4012 25516 4052 25556
rect 4108 25348 4148 25388
rect 3688 24928 3728 24968
rect 3770 24928 3810 24968
rect 3852 24928 3892 24968
rect 3934 24928 3974 24968
rect 4016 24928 4056 24968
rect 3688 23416 3728 23456
rect 3770 23416 3810 23456
rect 3852 23416 3892 23456
rect 3934 23416 3974 23456
rect 4016 23416 4056 23456
rect 3436 22996 3476 23036
rect 3148 15016 3188 15056
rect 3148 14848 3188 14888
rect 2764 12916 2804 12956
rect 2860 13000 2900 13040
rect 2764 9808 2804 9848
rect 3052 13756 3092 13796
rect 3052 9808 3092 9848
rect 3244 13756 3284 13796
rect 3436 15100 3476 15140
rect 2764 1408 2804 1448
rect 3244 148 3284 188
rect 3436 4264 3476 4304
rect 3916 22072 3956 22112
rect 3688 21904 3728 21944
rect 3770 21904 3810 21944
rect 3852 21904 3892 21944
rect 3934 21904 3974 21944
rect 4016 21904 4056 21944
rect 3688 20392 3728 20432
rect 3770 20392 3810 20432
rect 3852 20392 3892 20432
rect 3934 20392 3974 20432
rect 4016 20392 4056 20432
rect 3628 20224 3668 20264
rect 3628 19048 3668 19088
rect 3688 18880 3728 18920
rect 3770 18880 3810 18920
rect 3852 18880 3892 18920
rect 3934 18880 3974 18920
rect 4016 18880 4056 18920
rect 3724 18040 3764 18080
rect 4780 29968 4820 30008
rect 4492 29800 4532 29840
rect 4396 29044 4436 29084
rect 4588 27532 4628 27572
rect 4300 22996 4340 23036
rect 4396 22744 4436 22784
rect 4300 22072 4340 22112
rect 3688 17368 3728 17408
rect 3770 17368 3810 17408
rect 3852 17368 3892 17408
rect 3934 17368 3974 17408
rect 4016 17368 4056 17408
rect 3688 15856 3728 15896
rect 3770 15856 3810 15896
rect 3852 15856 3892 15896
rect 3934 15856 3974 15896
rect 4016 15856 4056 15896
rect 4012 15688 4052 15728
rect 3628 14848 3668 14888
rect 3724 14596 3764 14636
rect 4012 14680 4052 14720
rect 3688 14344 3728 14384
rect 3770 14344 3810 14384
rect 3852 14344 3892 14384
rect 3934 14344 3974 14384
rect 4016 14344 4056 14384
rect 4012 13252 4052 13292
rect 3688 12832 3728 12872
rect 3770 12832 3810 12872
rect 3852 12832 3892 12872
rect 3934 12832 3974 12872
rect 4016 12832 4056 12872
rect 4588 22492 4628 22532
rect 4492 20812 4532 20852
rect 4684 20140 4724 20180
rect 4204 17284 4244 17324
rect 4396 15016 4436 15056
rect 4300 14680 4340 14720
rect 4588 19132 4628 19172
rect 5260 30052 5300 30092
rect 4876 28876 4916 28916
rect 4928 28708 4968 28748
rect 5010 28708 5050 28748
rect 5092 28708 5132 28748
rect 5174 28708 5214 28748
rect 5256 28708 5296 28748
rect 4928 27196 4968 27236
rect 5010 27196 5050 27236
rect 5092 27196 5132 27236
rect 5174 27196 5214 27236
rect 5256 27196 5296 27236
rect 4972 26776 5012 26816
rect 5260 26440 5300 26480
rect 4928 25684 4968 25724
rect 5010 25684 5050 25724
rect 5092 25684 5132 25724
rect 5174 25684 5214 25724
rect 5256 25684 5296 25724
rect 5548 30220 5588 30260
rect 5644 32824 5684 32864
rect 5740 30472 5780 30512
rect 5452 25180 5492 25220
rect 4928 24172 4968 24212
rect 5010 24172 5050 24212
rect 5092 24172 5132 24212
rect 5174 24172 5214 24212
rect 5256 24172 5296 24212
rect 5740 28036 5780 28076
rect 6028 33328 6068 33368
rect 5932 28036 5972 28076
rect 6028 33160 6068 33200
rect 5740 26440 5780 26480
rect 5548 23080 5588 23120
rect 5260 22996 5300 23036
rect 4972 22828 5012 22868
rect 4928 22660 4968 22700
rect 5010 22660 5050 22700
rect 5092 22660 5132 22700
rect 5174 22660 5214 22700
rect 5256 22660 5296 22700
rect 5164 22492 5204 22532
rect 4972 21484 5012 21524
rect 5164 21316 5204 21356
rect 5356 21484 5396 21524
rect 4928 21148 4968 21188
rect 5010 21148 5050 21188
rect 5092 21148 5132 21188
rect 5174 21148 5214 21188
rect 5256 21148 5296 21188
rect 4972 20980 5012 21020
rect 5260 20980 5300 21020
rect 5068 20896 5108 20936
rect 5452 20980 5492 21020
rect 5356 20896 5396 20936
rect 5068 19804 5108 19844
rect 4928 19636 4968 19676
rect 5010 19636 5050 19676
rect 5092 19636 5132 19676
rect 5174 19636 5214 19676
rect 5256 19636 5296 19676
rect 4928 18124 4968 18164
rect 5010 18124 5050 18164
rect 5092 18124 5132 18164
rect 5174 18124 5214 18164
rect 5256 18124 5296 18164
rect 4588 16948 4628 16988
rect 4876 17956 4916 17996
rect 4972 17452 5012 17492
rect 5260 17620 5300 17660
rect 5164 17200 5204 17240
rect 4972 16780 5012 16820
rect 4928 16612 4968 16652
rect 5010 16612 5050 16652
rect 5092 16612 5132 16652
rect 5174 16612 5214 16652
rect 5256 16612 5296 16652
rect 4588 15688 4628 15728
rect 4492 14764 4532 14804
rect 5260 16192 5300 16232
rect 4928 15100 4968 15140
rect 5010 15100 5050 15140
rect 5092 15100 5132 15140
rect 5174 15100 5214 15140
rect 5256 15100 5296 15140
rect 5260 14932 5300 14972
rect 4396 14344 4436 14384
rect 3820 12496 3860 12536
rect 3688 11320 3728 11360
rect 3770 11320 3810 11360
rect 3852 11320 3892 11360
rect 3934 11320 3974 11360
rect 4016 11320 4056 11360
rect 4300 14008 4340 14048
rect 4300 13084 4340 13124
rect 4492 14008 4532 14048
rect 4780 14596 4820 14636
rect 5068 14512 5108 14552
rect 5260 14008 5300 14048
rect 5644 20980 5684 21020
rect 5548 17032 5588 17072
rect 5644 19300 5684 19340
rect 5836 18208 5876 18248
rect 5932 17872 5972 17912
rect 5644 16948 5684 16988
rect 5548 16864 5588 16904
rect 5452 14764 5492 14804
rect 5836 17032 5876 17072
rect 5644 14848 5684 14888
rect 5740 15016 5780 15056
rect 6220 34924 6260 34964
rect 6124 32320 6164 32360
rect 6412 34924 6452 34964
rect 6316 32320 6356 32360
rect 6412 31732 6452 31772
rect 6412 30052 6452 30092
rect 6220 17956 6260 17996
rect 6124 17872 6164 17912
rect 6220 17788 6260 17828
rect 6028 17032 6068 17072
rect 6028 16864 6068 16904
rect 5932 14680 5972 14720
rect 6028 16528 6068 16568
rect 5740 14428 5780 14468
rect 5164 13756 5204 13796
rect 4928 13588 4968 13628
rect 5010 13588 5050 13628
rect 5092 13588 5132 13628
rect 5174 13588 5214 13628
rect 5256 13588 5296 13628
rect 4396 11740 4436 11780
rect 4492 13168 4532 13208
rect 4396 11572 4436 11612
rect 4300 10732 4340 10772
rect 3688 9808 3728 9848
rect 3770 9808 3810 9848
rect 3852 9808 3892 9848
rect 3934 9808 3974 9848
rect 4016 9808 4056 9848
rect 3688 8296 3728 8336
rect 3770 8296 3810 8336
rect 3852 8296 3892 8336
rect 3934 8296 3974 8336
rect 4016 8296 4056 8336
rect 3688 6784 3728 6824
rect 3770 6784 3810 6824
rect 3852 6784 3892 6824
rect 3934 6784 3974 6824
rect 4016 6784 4056 6824
rect 4588 12244 4628 12284
rect 4972 13420 5012 13460
rect 5356 13252 5396 13292
rect 5452 14008 5492 14048
rect 5260 13168 5300 13208
rect 4972 12580 5012 12620
rect 4928 12076 4968 12116
rect 5010 12076 5050 12116
rect 5092 12076 5132 12116
rect 5174 12076 5214 12116
rect 5256 12076 5296 12116
rect 4588 9556 4628 9596
rect 3688 5272 3728 5312
rect 3770 5272 3810 5312
rect 3852 5272 3892 5312
rect 3934 5272 3974 5312
rect 4016 5272 4056 5312
rect 3688 3760 3728 3800
rect 3770 3760 3810 3800
rect 3852 3760 3892 3800
rect 3934 3760 3974 3800
rect 4016 3760 4056 3800
rect 4928 10564 4968 10604
rect 5010 10564 5050 10604
rect 5092 10564 5132 10604
rect 5174 10564 5214 10604
rect 5256 10564 5296 10604
rect 5740 12580 5780 12620
rect 5836 13420 5876 13460
rect 8908 44920 8948 44960
rect 6604 21484 6644 21524
rect 7084 33244 7124 33284
rect 7084 32572 7124 32612
rect 6412 17788 6452 17828
rect 6604 17956 6644 17996
rect 5740 12328 5780 12368
rect 5740 11572 5780 11612
rect 5548 9472 5588 9512
rect 5644 9304 5684 9344
rect 4928 9052 4968 9092
rect 5010 9052 5050 9092
rect 5092 9052 5132 9092
rect 5174 9052 5214 9092
rect 5256 9052 5296 9092
rect 5068 8716 5108 8756
rect 5452 8716 5492 8756
rect 4928 7540 4968 7580
rect 5010 7540 5050 7580
rect 5092 7540 5132 7580
rect 5174 7540 5214 7580
rect 5256 7540 5296 7580
rect 4876 7204 4916 7244
rect 4972 7120 5012 7160
rect 3688 2248 3728 2288
rect 3770 2248 3810 2288
rect 3852 2248 3892 2288
rect 3934 2248 3974 2288
rect 4016 2248 4056 2288
rect 4928 6028 4968 6068
rect 5010 6028 5050 6068
rect 5092 6028 5132 6068
rect 5174 6028 5214 6068
rect 5256 6028 5296 6068
rect 4928 4516 4968 4556
rect 5010 4516 5050 4556
rect 5092 4516 5132 4556
rect 5174 4516 5214 4556
rect 5256 4516 5296 4556
rect 4928 3004 4968 3044
rect 5010 3004 5050 3044
rect 5092 3004 5132 3044
rect 5174 3004 5214 3044
rect 5256 3004 5296 3044
rect 5740 8968 5780 9008
rect 5740 8716 5780 8756
rect 6316 16696 6356 16736
rect 6316 14764 6356 14804
rect 6124 12916 6164 12956
rect 6124 12412 6164 12452
rect 6508 16024 6548 16064
rect 6508 14680 6548 14720
rect 6412 13252 6452 13292
rect 5740 7708 5780 7748
rect 6316 11740 6356 11780
rect 6700 17704 6740 17744
rect 7276 37444 7316 37484
rect 7276 33664 7316 33704
rect 7180 24508 7220 24548
rect 7660 37444 7700 37484
rect 7468 30724 7508 30764
rect 7468 25432 7508 25472
rect 6988 17956 7028 17996
rect 7756 32824 7796 32864
rect 7852 30724 7892 30764
rect 6988 17200 7028 17240
rect 6892 16276 6932 16316
rect 7276 17956 7316 17996
rect 7276 17452 7316 17492
rect 7660 18040 7700 18080
rect 8620 43408 8660 43448
rect 8044 30556 8084 30596
rect 8428 30388 8468 30428
rect 8524 28792 8564 28832
rect 7852 21652 7892 21692
rect 9484 35596 9524 35636
rect 9292 35428 9332 35468
rect 7372 17200 7412 17240
rect 7468 17032 7508 17072
rect 7180 16192 7220 16232
rect 7084 16024 7124 16064
rect 7084 14680 7124 14720
rect 7276 15100 7316 15140
rect 7372 15016 7412 15056
rect 7084 13084 7124 13124
rect 7180 13756 7220 13796
rect 6892 12916 6932 12956
rect 7180 12940 7220 12980
rect 6220 10480 6260 10520
rect 6316 10648 6356 10688
rect 6220 10060 6260 10100
rect 6220 8800 6260 8840
rect 6700 10060 6740 10100
rect 6508 9976 6548 10016
rect 6604 9472 6644 9512
rect 6796 8800 6836 8840
rect 6796 8632 6836 8672
rect 7372 12916 7412 12956
rect 7180 12832 7220 12872
rect 7276 12664 7316 12704
rect 7180 12412 7220 12452
rect 6988 9388 7028 9428
rect 7180 8800 7220 8840
rect 7756 17284 7796 17324
rect 7564 14596 7604 14636
rect 7852 17032 7892 17072
rect 7468 12664 7508 12704
rect 7468 12328 7508 12368
rect 7948 14848 7988 14888
rect 7852 14596 7892 14636
rect 7660 12328 7700 12368
rect 8140 16192 8180 16232
rect 8140 16024 8180 16064
rect 8236 14512 8276 14552
rect 8428 20812 8468 20852
rect 8524 16612 8564 16652
rect 9772 38872 9812 38912
rect 9388 32992 9428 33032
rect 9100 29296 9140 29336
rect 8908 22492 8948 22532
rect 9388 31396 9428 31436
rect 9676 35596 9716 35636
rect 9388 30892 9428 30932
rect 9580 32992 9620 33032
rect 9676 31396 9716 31436
rect 9964 35428 10004 35468
rect 9868 30640 9908 30680
rect 9292 24592 9332 24632
rect 8428 15688 8468 15728
rect 8428 14428 8468 14468
rect 8140 13504 8180 13544
rect 8044 11908 8084 11948
rect 7852 10648 7892 10688
rect 7564 6364 7604 6404
rect 8044 7876 8084 7916
rect 8428 14260 8468 14300
rect 8716 14176 8756 14216
rect 8620 13840 8660 13880
rect 8428 13504 8468 13544
rect 8620 12748 8660 12788
rect 8428 10648 8468 10688
rect 8812 13000 8852 13040
rect 8524 8800 8564 8840
rect 8524 8128 8564 8168
rect 8524 7540 8564 7580
rect 5740 2416 5780 2456
rect 4928 1492 4968 1532
rect 5010 1492 5050 1532
rect 5092 1492 5132 1532
rect 5174 1492 5214 1532
rect 5256 1492 5296 1532
rect 5644 1408 5684 1448
rect 4492 904 4532 944
rect 3916 64 3956 104
rect 5068 148 5108 188
rect 6220 1408 6260 1448
rect 6796 1240 6836 1280
rect 7372 232 7412 272
rect 8236 2836 8276 2876
rect 9868 26020 9908 26060
rect 9676 22660 9716 22700
rect 9388 17872 9428 17912
rect 9100 15520 9140 15560
rect 9100 13336 9140 13376
rect 9484 17620 9524 17660
rect 9484 13336 9524 13376
rect 9580 14512 9620 14552
rect 10156 33160 10196 33200
rect 10156 32740 10196 32780
rect 10156 32488 10196 32528
rect 10060 30640 10100 30680
rect 10636 44752 10676 44792
rect 10060 29212 10100 29252
rect 10252 28960 10292 29000
rect 10156 27448 10196 27488
rect 10060 27196 10100 27236
rect 10060 26188 10100 26228
rect 10060 25936 10100 25976
rect 10060 23752 10100 23792
rect 9868 22660 9908 22700
rect 9868 22492 9908 22532
rect 9772 17872 9812 17912
rect 10732 37276 10772 37316
rect 10444 32404 10484 32444
rect 10636 32992 10676 33032
rect 10636 32404 10676 32444
rect 10444 30220 10484 30260
rect 10636 30304 10676 30344
rect 10540 30136 10580 30176
rect 10828 32656 10868 32696
rect 11116 44248 11156 44288
rect 11500 45760 11540 45800
rect 11500 44920 11540 44960
rect 11500 43660 11540 43700
rect 11020 41812 11060 41852
rect 11596 42736 11636 42776
rect 11500 40300 11540 40340
rect 11116 38872 11156 38912
rect 11020 32740 11060 32780
rect 10828 30892 10868 30932
rect 10444 28960 10484 29000
rect 10540 29884 10580 29924
rect 10636 29296 10676 29336
rect 10636 28960 10676 29000
rect 10348 27448 10388 27488
rect 10924 29884 10964 29924
rect 10828 28960 10868 29000
rect 10540 27364 10580 27404
rect 9964 17956 10004 17996
rect 10156 18376 10196 18416
rect 9772 14428 9812 14468
rect 9484 12748 9524 12788
rect 9388 9472 9428 9512
rect 9580 12664 9620 12704
rect 10540 23416 10580 23456
rect 10924 26692 10964 26732
rect 10444 19216 10484 19256
rect 10348 18376 10388 18416
rect 9964 12748 10004 12788
rect 11404 37192 11444 37232
rect 11212 32740 11252 32780
rect 11404 33076 11444 33116
rect 11404 32824 11444 32864
rect 11404 32572 11444 32612
rect 11308 30556 11348 30596
rect 11884 44668 11924 44708
rect 11884 43324 11924 43364
rect 11980 41896 12020 41936
rect 11788 39376 11828 39416
rect 11884 38872 11924 38912
rect 11596 33832 11636 33872
rect 11884 38200 11924 38240
rect 11884 37360 11924 37400
rect 11884 36520 11924 36560
rect 11980 33832 12020 33872
rect 11500 31480 11540 31520
rect 11308 29548 11348 29588
rect 11308 29212 11348 29252
rect 11404 28792 11444 28832
rect 11692 33160 11732 33200
rect 11596 27532 11636 27572
rect 11404 26188 11444 26228
rect 10828 23500 10868 23540
rect 10828 23248 10868 23288
rect 10924 22660 10964 22700
rect 11020 21316 11060 21356
rect 10732 16864 10772 16904
rect 10732 16696 10772 16736
rect 10540 14176 10580 14216
rect 10732 15940 10772 15980
rect 10732 14680 10772 14720
rect 10732 14512 10772 14552
rect 10732 14260 10772 14300
rect 9964 4936 10004 4976
rect 10924 16780 10964 16820
rect 10924 15940 10964 15980
rect 11212 24760 11252 24800
rect 11500 24760 11540 24800
rect 11692 27364 11732 27404
rect 11788 28792 11828 28832
rect 11212 23416 11252 23456
rect 11212 19132 11252 19172
rect 11308 16780 11348 16820
rect 11212 16696 11252 16736
rect 11788 26440 11828 26480
rect 11500 16864 11540 16904
rect 11692 17452 11732 17492
rect 12364 44836 12404 44876
rect 12268 39376 12308 39416
rect 12364 38956 12404 38996
rect 12268 34336 12308 34376
rect 12268 33664 12308 33704
rect 12556 36184 12596 36224
rect 12556 34336 12596 34376
rect 12748 36520 12788 36560
rect 12556 33832 12596 33872
rect 12364 32992 12404 33032
rect 12460 31480 12500 31520
rect 12364 29800 12404 29840
rect 12172 29212 12212 29252
rect 11980 24592 12020 24632
rect 11884 19888 11924 19928
rect 11884 18628 11924 18668
rect 12940 36184 12980 36224
rect 12844 33496 12884 33536
rect 12460 27448 12500 27488
rect 12268 21316 12308 21356
rect 12268 18292 12308 18332
rect 12076 18208 12116 18248
rect 12844 28036 12884 28076
rect 12844 27868 12884 27908
rect 12748 27448 12788 27488
rect 12556 21316 12596 21356
rect 12652 26188 12692 26228
rect 12460 19888 12500 19928
rect 12460 19048 12500 19088
rect 11884 17116 11924 17156
rect 11980 17284 12020 17324
rect 11788 17032 11828 17072
rect 11596 16024 11636 16064
rect 11980 16276 12020 16316
rect 11788 13840 11828 13880
rect 11500 11908 11540 11948
rect 11404 11572 11444 11612
rect 12364 17956 12404 17996
rect 12172 17032 12212 17072
rect 12844 25180 12884 25220
rect 12748 19048 12788 19088
rect 12652 17956 12692 17996
rect 11788 9640 11828 9680
rect 12172 8632 12212 8672
rect 13132 33496 13172 33536
rect 13420 32992 13460 33032
rect 13132 29044 13172 29084
rect 13420 27952 13460 27992
rect 13036 24592 13076 24632
rect 13036 18628 13076 18668
rect 12940 18544 12980 18584
rect 13228 25180 13268 25220
rect 13228 23080 13268 23120
rect 12844 16360 12884 16400
rect 12652 13840 12692 13880
rect 13036 14848 13076 14888
rect 12268 7960 12308 8000
rect 10348 5608 10388 5648
rect 12556 4264 12596 4304
rect 9100 988 9140 1028
rect 9676 988 9716 1028
rect 10252 988 10292 1028
rect 10828 988 10868 1028
rect 11404 988 11444 1028
rect 11980 652 12020 692
rect 13324 18628 13364 18668
rect 13516 23500 13556 23540
rect 13612 29212 13652 29252
rect 13420 18376 13460 18416
rect 13612 20140 13652 20180
rect 13612 18544 13652 18584
rect 13612 14848 13652 14888
<< metal4 >>
rect 4919 46852 4928 46892
rect 4968 46852 5010 46892
rect 5050 46852 5092 46892
rect 5132 46852 5174 46892
rect 5214 46852 5256 46892
rect 5296 46852 5305 46892
rect 1805 46432 1900 46472
rect 1940 46432 1949 46472
rect 3679 46096 3688 46136
rect 3728 46096 3770 46136
rect 3810 46096 3852 46136
rect 3892 46096 3934 46136
rect 3974 46096 4016 46136
rect 4056 46096 4065 46136
rect 10819 45760 10828 45800
rect 10868 45760 11500 45800
rect 11540 45760 11549 45800
rect 4919 45340 4928 45380
rect 4968 45340 5010 45380
rect 5050 45340 5092 45380
rect 5132 45340 5174 45380
rect 5214 45340 5256 45380
rect 5296 45340 5305 45380
rect 5443 44920 5452 44960
rect 5492 44920 5644 44960
rect 5684 44920 5693 44960
rect 8813 44920 8908 44960
rect 8948 44920 8957 44960
rect 9283 44920 9292 44960
rect 9332 44920 11500 44960
rect 11540 44920 11549 44960
rect 10243 44836 10252 44876
rect 10292 44836 12364 44876
rect 12404 44836 12413 44876
rect 6403 44752 6412 44792
rect 6452 44752 10636 44792
rect 10676 44752 10685 44792
rect 10627 44668 10636 44708
rect 10676 44668 11884 44708
rect 11924 44668 11933 44708
rect 3679 44584 3688 44624
rect 3728 44584 3770 44624
rect 3810 44584 3852 44624
rect 3892 44584 3934 44624
rect 3974 44584 4016 44624
rect 4056 44584 4065 44624
rect 9475 44248 9484 44288
rect 9524 44248 11116 44288
rect 11156 44248 11165 44288
rect 4919 43828 4928 43868
rect 4968 43828 5010 43868
rect 5050 43828 5092 43868
rect 5132 43828 5174 43868
rect 5214 43828 5256 43868
rect 5296 43828 5305 43868
rect 6595 43660 6604 43700
rect 6644 43660 11500 43700
rect 11540 43660 11549 43700
rect 8525 43408 8620 43448
rect 8660 43408 8669 43448
rect 6787 43324 6796 43364
rect 6836 43324 11884 43364
rect 11924 43324 11933 43364
rect 3679 43072 3688 43112
rect 3728 43072 3770 43112
rect 3810 43072 3852 43112
rect 3892 43072 3934 43112
rect 3974 43072 4016 43112
rect 4056 43072 4065 43112
rect 11203 42736 11212 42776
rect 11252 42736 11596 42776
rect 11636 42736 11645 42776
rect 4919 42316 4928 42356
rect 4968 42316 5010 42356
rect 5050 42316 5092 42356
rect 5132 42316 5174 42356
rect 5214 42316 5256 42356
rect 5296 42316 5305 42356
rect 10435 41896 10444 41936
rect 10484 41896 11980 41936
rect 12020 41896 12029 41936
rect 11011 41812 11020 41852
rect 11060 41812 11404 41852
rect 11444 41812 11453 41852
rect 3679 41560 3688 41600
rect 3728 41560 3770 41600
rect 3810 41560 3852 41600
rect 3892 41560 3934 41600
rect 3974 41560 4016 41600
rect 4056 41560 4065 41600
rect 4919 40804 4928 40844
rect 4968 40804 5010 40844
rect 5050 40804 5092 40844
rect 5132 40804 5174 40844
rect 5214 40804 5256 40844
rect 5296 40804 5305 40844
rect 3341 40300 3436 40340
rect 3476 40300 3485 40340
rect 4493 40300 4588 40340
rect 4628 40300 4637 40340
rect 6499 40300 6508 40340
rect 6548 40300 11500 40340
rect 11540 40300 11549 40340
rect 3679 40048 3688 40088
rect 3728 40048 3770 40088
rect 3810 40048 3852 40088
rect 3892 40048 3934 40088
rect 3974 40048 4016 40088
rect 4056 40048 4065 40088
rect 11779 39376 11788 39416
rect 11828 39376 12268 39416
rect 12308 39376 12317 39416
rect 4919 39292 4928 39332
rect 4968 39292 5010 39332
rect 5050 39292 5092 39332
rect 5132 39292 5174 39332
rect 5214 39292 5256 39332
rect 5296 39292 5305 39332
rect 10915 38956 10924 38996
rect 10964 38956 12364 38996
rect 12404 38956 12413 38996
rect 9677 38872 9772 38912
rect 9812 38872 9821 38912
rect 11021 38872 11116 38912
rect 11156 38872 11165 38912
rect 11789 38872 11884 38912
rect 11924 38872 11933 38912
rect 3679 38536 3688 38576
rect 3728 38536 3770 38576
rect 3810 38536 3852 38576
rect 3892 38536 3934 38576
rect 3974 38536 4016 38576
rect 4056 38536 4065 38576
rect 4675 38284 4684 38324
rect 4724 38284 5452 38324
rect 5492 38284 5501 38324
rect 11011 38200 11020 38240
rect 11060 38200 11884 38240
rect 11924 38200 11933 38240
rect 4483 37948 4492 37988
rect 4532 37948 5356 37988
rect 5396 37948 5405 37988
rect 4919 37780 4928 37820
rect 4968 37780 5010 37820
rect 5050 37780 5092 37820
rect 5132 37780 5174 37820
rect 5214 37780 5256 37820
rect 5296 37780 5305 37820
rect 7171 37444 7180 37484
rect 7220 37444 7276 37484
rect 7316 37444 7660 37484
rect 7700 37444 7709 37484
rect 11875 37360 11884 37400
rect 11924 37360 11980 37400
rect 12020 37360 12029 37400
rect 9091 37276 9100 37316
rect 9140 37276 10732 37316
rect 10772 37276 10781 37316
rect 9571 37192 9580 37232
rect 9620 37192 11404 37232
rect 11444 37192 11453 37232
rect 3679 37024 3688 37064
rect 3728 37024 3770 37064
rect 3810 37024 3852 37064
rect 3892 37024 3934 37064
rect 3974 37024 4016 37064
rect 4056 37024 4065 37064
rect 11875 36520 11884 36560
rect 11924 36520 12748 36560
rect 12788 36520 12797 36560
rect 4919 36268 4928 36308
rect 4968 36268 5010 36308
rect 5050 36268 5092 36308
rect 5132 36268 5174 36308
rect 5214 36268 5256 36308
rect 5296 36268 5305 36308
rect 12547 36184 12556 36224
rect 12596 36184 12940 36224
rect 12980 36184 12989 36224
rect 9475 35596 9484 35636
rect 9524 35596 9676 35636
rect 9716 35596 9725 35636
rect 3679 35512 3688 35552
rect 3728 35512 3770 35552
rect 3810 35512 3852 35552
rect 3892 35512 3934 35552
rect 3974 35512 4016 35552
rect 4056 35512 4065 35552
rect 9283 35428 9292 35468
rect 9332 35428 9964 35468
rect 10004 35428 10013 35468
rect 6211 34924 6220 34964
rect 6260 34924 6412 34964
rect 6452 34924 6461 34964
rect 4919 34756 4928 34796
rect 4968 34756 5010 34796
rect 5050 34756 5092 34796
rect 5132 34756 5174 34796
rect 5214 34756 5256 34796
rect 5296 34756 5305 34796
rect 10339 34336 10348 34376
rect 10388 34336 12268 34376
rect 12308 34336 12317 34376
rect 12547 34336 12556 34376
rect 12596 34336 12605 34376
rect 3679 34000 3688 34040
rect 3728 34000 3770 34040
rect 3810 34000 3852 34040
rect 3892 34000 3934 34040
rect 3974 34000 4016 34040
rect 4056 34000 4065 34040
rect 12556 33872 12596 34336
rect 11587 33832 11596 33872
rect 11636 33832 11980 33872
rect 12020 33832 12029 33872
rect 12547 33832 12556 33872
rect 12596 33832 12605 33872
rect 7181 33664 7276 33704
rect 7316 33664 7325 33704
rect 12067 33664 12076 33704
rect 12116 33664 12268 33704
rect 12308 33664 12317 33704
rect 12835 33496 12844 33536
rect 12884 33496 13132 33536
rect 13172 33496 13181 33536
rect 6019 33328 6028 33368
rect 6068 33328 6124 33368
rect 6164 33328 6173 33368
rect 4919 33244 4928 33284
rect 4968 33244 5010 33284
rect 5050 33244 5092 33284
rect 5132 33244 5174 33284
rect 5214 33244 5256 33284
rect 5296 33244 5305 33284
rect 7075 33244 7084 33284
rect 7124 33244 7133 33284
rect 7084 33200 7124 33244
rect 6019 33160 6028 33200
rect 6068 33160 7124 33200
rect 10147 33160 10156 33200
rect 10196 33160 11692 33200
rect 11732 33160 11741 33200
rect 10531 33076 10540 33116
rect 10580 33076 11404 33116
rect 11444 33076 11453 33116
rect 9379 32992 9388 33032
rect 9428 32992 9580 33032
rect 9620 32992 9629 33032
rect 10627 32992 10636 33032
rect 10676 32992 11540 33032
rect 12355 32992 12364 33032
rect 12404 32992 13420 33032
rect 13460 32992 13469 33032
rect 3139 32908 3148 32948
rect 3188 32908 3436 32948
rect 3476 32908 3485 32948
rect 5635 32824 5644 32864
rect 5684 32824 7756 32864
rect 7796 32824 7805 32864
rect 8035 32824 8044 32864
rect 8084 32824 11404 32864
rect 11444 32824 11453 32864
rect 11500 32780 11540 32992
rect 10147 32740 10156 32780
rect 10196 32740 11020 32780
rect 11060 32740 11212 32780
rect 11252 32740 11261 32780
rect 11404 32740 11540 32780
rect 10723 32656 10732 32696
rect 10772 32656 10828 32696
rect 10868 32656 10877 32696
rect 11404 32612 11444 32740
rect 2851 32572 2860 32612
rect 2900 32572 7084 32612
rect 7124 32572 7133 32612
rect 11395 32572 11404 32612
rect 11444 32572 11453 32612
rect 3679 32488 3688 32528
rect 3728 32488 3770 32528
rect 3810 32488 3852 32528
rect 3892 32488 3934 32528
rect 3974 32488 4016 32528
rect 4056 32488 4065 32528
rect 10147 32488 10156 32528
rect 10196 32488 10540 32528
rect 10580 32488 10589 32528
rect 10435 32404 10444 32444
rect 10484 32404 10636 32444
rect 10676 32404 10685 32444
rect 6115 32320 6124 32360
rect 6164 32320 6316 32360
rect 6356 32320 6365 32360
rect 4291 32236 4300 32276
rect 4340 32236 4349 32276
rect 4300 32024 4340 32236
rect 4300 31984 4396 32024
rect 4436 31984 4445 32024
rect 4003 31900 4012 31940
rect 4052 31900 5164 31940
rect 5204 31900 5213 31940
rect 4919 31732 4928 31772
rect 4968 31732 5010 31772
rect 5050 31732 5092 31772
rect 5132 31732 5174 31772
rect 5214 31732 5256 31772
rect 5296 31732 5305 31772
rect 6307 31732 6316 31772
rect 6356 31732 6412 31772
rect 6452 31732 6461 31772
rect 11491 31480 11500 31520
rect 11540 31480 12460 31520
rect 12500 31480 12509 31520
rect 9379 31396 9388 31436
rect 9428 31396 9676 31436
rect 9716 31396 9725 31436
rect 3679 30976 3688 31016
rect 3728 30976 3770 31016
rect 3810 30976 3852 31016
rect 3892 30976 3934 31016
rect 3974 30976 4016 31016
rect 4056 30976 4065 31016
rect 9379 30892 9388 30932
rect 9428 30892 10828 30932
rect 10868 30892 10877 30932
rect 2659 30808 2668 30848
rect 2708 30808 3820 30848
rect 3860 30808 3869 30848
rect 3427 30724 3436 30764
rect 3476 30724 4012 30764
rect 4052 30724 4061 30764
rect 7459 30724 7468 30764
rect 7508 30724 7852 30764
rect 7892 30724 7901 30764
rect 9859 30640 9868 30680
rect 9908 30640 10060 30680
rect 10100 30640 10109 30680
rect 3427 30556 3436 30596
rect 3476 30556 8044 30596
rect 8084 30556 8093 30596
rect 10147 30556 10156 30596
rect 10196 30556 11308 30596
rect 11348 30556 11357 30596
rect 4099 30472 4108 30512
rect 4148 30472 5740 30512
rect 5780 30472 5789 30512
rect 2755 30388 2764 30428
rect 2804 30388 8428 30428
rect 8468 30388 8477 30428
rect 10627 30304 10636 30344
rect 10676 30304 10868 30344
rect 4205 30220 4300 30260
rect 4340 30220 4349 30260
rect 4397 30220 4492 30260
rect 4532 30220 4541 30260
rect 4589 30220 4684 30260
rect 4724 30220 4733 30260
rect 4919 30220 4928 30260
rect 4968 30220 5010 30260
rect 5050 30220 5092 30260
rect 5132 30220 5174 30260
rect 5214 30220 5256 30260
rect 5296 30220 5305 30260
rect 5539 30220 5548 30260
rect 5588 30220 6220 30260
rect 6260 30220 6269 30260
rect 8515 30220 8524 30260
rect 8564 30220 10100 30260
rect 10435 30220 10444 30260
rect 10484 30220 10493 30260
rect 1987 30136 1996 30176
rect 2036 30136 4396 30176
rect 4436 30136 4445 30176
rect 4492 30136 4588 30176
rect 4628 30136 4637 30176
rect 4492 29840 4532 30136
rect 10060 30092 10100 30220
rect 10444 30092 10484 30220
rect 10828 30176 10868 30304
rect 10531 30136 10540 30176
rect 10580 30136 10772 30176
rect 10828 30136 11596 30176
rect 11636 30136 11645 30176
rect 5251 30052 5260 30092
rect 5300 30052 6124 30092
rect 6164 30052 6412 30092
rect 6452 30052 6461 30092
rect 10060 30052 10292 30092
rect 10444 30052 10676 30092
rect 4675 29968 4684 30008
rect 4724 29968 4780 30008
rect 4820 29968 4829 30008
rect 10252 29840 10292 30052
rect 10636 29924 10676 30052
rect 10531 29884 10540 29924
rect 10580 29884 10676 29924
rect 10732 29924 10772 30136
rect 10732 29884 10924 29924
rect 10964 29884 10973 29924
rect 4483 29800 4492 29840
rect 4532 29800 4541 29840
rect 10252 29800 12364 29840
rect 12404 29800 12413 29840
rect 3523 29716 3532 29756
rect 3572 29716 3820 29756
rect 3860 29716 3869 29756
rect 3331 29632 3340 29672
rect 3380 29632 3724 29672
rect 3764 29632 3773 29672
rect 11299 29548 11308 29588
rect 11348 29548 11444 29588
rect 3679 29464 3688 29504
rect 3728 29464 3770 29504
rect 3810 29464 3852 29504
rect 3892 29464 3934 29504
rect 3974 29464 4016 29504
rect 4056 29464 4065 29504
rect 9091 29296 9100 29336
rect 9140 29296 10636 29336
rect 10676 29296 10685 29336
rect 3043 29212 3052 29252
rect 3092 29212 3148 29252
rect 3188 29212 3197 29252
rect 10051 29212 10060 29252
rect 10100 29212 11308 29252
rect 11348 29212 11357 29252
rect 4291 29044 4300 29084
rect 4340 29044 4396 29084
rect 4436 29044 4445 29084
rect 10243 28960 10252 29000
rect 10292 28960 10444 29000
rect 10484 28960 10493 29000
rect 10627 28960 10636 29000
rect 10676 28960 10828 29000
rect 10868 28960 10877 29000
rect 4675 28876 4684 28916
rect 4724 28876 4876 28916
rect 4916 28876 4925 28916
rect 11404 28832 11444 29548
rect 12163 29212 12172 29252
rect 12212 29212 13612 29252
rect 13652 29212 13661 29252
rect 12835 29044 12844 29084
rect 12884 29044 13132 29084
rect 13172 29044 13181 29084
rect 8515 28792 8524 28832
rect 8564 28792 8716 28832
rect 8756 28792 8765 28832
rect 11395 28792 11404 28832
rect 11444 28792 11453 28832
rect 11779 28792 11788 28832
rect 11828 28792 12076 28832
rect 12116 28792 12125 28832
rect 4919 28708 4928 28748
rect 4968 28708 5010 28748
rect 5050 28708 5092 28748
rect 5132 28708 5174 28748
rect 5214 28708 5256 28748
rect 5296 28708 5305 28748
rect 5731 28036 5740 28076
rect 5780 28036 5932 28076
rect 5972 28036 5981 28076
rect 12835 28036 12844 28076
rect 12884 28036 12893 28076
rect 12844 27992 12884 28036
rect 3679 27952 3688 27992
rect 3728 27952 3770 27992
rect 3810 27952 3852 27992
rect 3892 27952 3934 27992
rect 3974 27952 4016 27992
rect 4056 27952 4065 27992
rect 12844 27952 13420 27992
rect 13460 27952 13469 27992
rect 12749 27868 12844 27908
rect 12884 27868 12893 27908
rect 4579 27532 4588 27572
rect 4628 27532 4780 27572
rect 4820 27532 4829 27572
rect 11501 27532 11596 27572
rect 11636 27532 11645 27572
rect 10147 27448 10156 27488
rect 10196 27448 10348 27488
rect 10388 27448 10397 27488
rect 12451 27448 12460 27488
rect 12500 27448 12748 27488
rect 12788 27448 12797 27488
rect 10445 27364 10540 27404
rect 10580 27364 10589 27404
rect 11597 27364 11692 27404
rect 11732 27364 11741 27404
rect 4919 27196 4928 27236
rect 4968 27196 5010 27236
rect 5050 27196 5092 27236
rect 5132 27196 5174 27236
rect 5214 27196 5256 27236
rect 5296 27196 5305 27236
rect 10051 27196 10060 27236
rect 10100 27196 10540 27236
rect 10580 27196 10589 27236
rect 4675 26776 4684 26816
rect 4724 26776 4972 26816
rect 5012 26776 5021 26816
rect 10915 26692 10924 26732
rect 10964 26692 11308 26732
rect 11348 26692 11357 26732
rect 3679 26440 3688 26480
rect 3728 26440 3770 26480
rect 3810 26440 3852 26480
rect 3892 26440 3934 26480
rect 3974 26440 4016 26480
rect 4056 26440 4065 26480
rect 5251 26440 5260 26480
rect 5300 26440 5740 26480
rect 5780 26440 5789 26480
rect 11683 26440 11692 26480
rect 11732 26440 11788 26480
rect 11828 26440 11837 26480
rect 10051 26188 10060 26228
rect 10100 26188 10109 26228
rect 11395 26188 11404 26228
rect 11444 26188 12652 26228
rect 12692 26188 12701 26228
rect 10060 26060 10100 26188
rect 3043 26020 3052 26060
rect 3092 26020 4108 26060
rect 4148 26020 4157 26060
rect 9859 26020 9868 26060
rect 9908 26020 10100 26060
rect 10051 25936 10060 25976
rect 10100 25936 10540 25976
rect 10580 25936 10589 25976
rect 4919 25684 4928 25724
rect 4968 25684 5010 25724
rect 5050 25684 5092 25724
rect 5132 25684 5174 25724
rect 5214 25684 5256 25724
rect 5296 25684 5305 25724
rect 3427 25516 3436 25556
rect 3476 25516 4012 25556
rect 4052 25516 4061 25556
rect 7459 25432 7468 25472
rect 7508 25432 7564 25472
rect 7604 25432 7613 25472
rect 2659 25348 2668 25388
rect 2708 25348 3532 25388
rect 3572 25348 4108 25388
rect 4148 25348 4157 25388
rect 5443 25180 5452 25220
rect 5492 25180 5740 25220
rect 5780 25180 5789 25220
rect 12835 25180 12844 25220
rect 12884 25180 13228 25220
rect 13268 25180 13277 25220
rect 2275 25096 2284 25136
rect 2324 25096 5548 25136
rect 5588 25096 5597 25136
rect 3679 24928 3688 24968
rect 3728 24928 3770 24968
rect 3810 24928 3852 24968
rect 3892 24928 3934 24968
rect 3974 24928 4016 24968
rect 4056 24928 4065 24968
rect 11203 24760 11212 24800
rect 11252 24760 11500 24800
rect 11540 24760 11549 24800
rect 1411 24592 1420 24632
rect 1460 24592 9292 24632
rect 9332 24592 9341 24632
rect 11971 24592 11980 24632
rect 12020 24592 13036 24632
rect 13076 24592 13085 24632
rect 7171 24508 7180 24548
rect 7220 24508 7468 24548
rect 7508 24508 7517 24548
rect 9667 24340 9676 24380
rect 9716 24340 10636 24380
rect 10676 24340 10685 24380
rect 4919 24172 4928 24212
rect 4968 24172 5010 24212
rect 5050 24172 5092 24212
rect 5132 24172 5174 24212
rect 5214 24172 5256 24212
rect 5296 24172 5305 24212
rect 8227 23752 8236 23792
rect 8276 23752 10060 23792
rect 10100 23752 10109 23792
rect 1507 23500 1516 23540
rect 1556 23500 10828 23540
rect 10868 23500 10877 23540
rect 13507 23500 13516 23540
rect 13556 23500 13565 23540
rect 3679 23416 3688 23456
rect 3728 23416 3770 23456
rect 3810 23416 3852 23456
rect 3892 23416 3934 23456
rect 3974 23416 4016 23456
rect 4056 23416 4065 23456
rect 10531 23416 10540 23456
rect 10580 23416 11212 23456
rect 11252 23416 11261 23456
rect 2860 23248 10828 23288
rect 10868 23248 10877 23288
rect 2860 23120 2900 23248
rect 13516 23204 13556 23500
rect 2947 23164 2956 23204
rect 2996 23164 3052 23204
rect 3092 23164 3101 23204
rect 13228 23164 13556 23204
rect 13228 23120 13268 23164
rect 1699 23080 1708 23120
rect 1748 23080 2900 23120
rect 5539 23080 5548 23120
rect 5588 23080 5597 23120
rect 13219 23080 13228 23120
rect 13268 23080 13277 23120
rect 5548 23036 5588 23080
rect 2659 22996 2668 23036
rect 2708 22996 2860 23036
rect 2900 22996 2909 23036
rect 3331 22996 3340 23036
rect 3380 22996 3436 23036
rect 3476 22996 3485 23036
rect 4205 22996 4300 23036
rect 4340 22996 4349 23036
rect 5251 22996 5260 23036
rect 5300 22996 5452 23036
rect 5492 22996 5588 23036
rect 4963 22828 4972 22868
rect 5012 22828 5021 22868
rect 4972 22784 5012 22828
rect 4387 22744 4396 22784
rect 4436 22744 5012 22784
rect 4919 22660 4928 22700
rect 4968 22660 5010 22700
rect 5050 22660 5092 22700
rect 5132 22660 5174 22700
rect 5214 22660 5256 22700
rect 5296 22660 5305 22700
rect 9667 22660 9676 22700
rect 9716 22660 9868 22700
rect 9908 22660 9917 22700
rect 10531 22660 10540 22700
rect 10580 22660 10924 22700
rect 10964 22660 10973 22700
rect 4579 22492 4588 22532
rect 4628 22492 5164 22532
rect 5204 22492 5213 22532
rect 8899 22492 8908 22532
rect 8948 22492 9868 22532
rect 9908 22492 9917 22532
rect 2275 22408 2284 22448
rect 2324 22408 2572 22448
rect 2612 22408 2621 22448
rect 2563 22240 2572 22280
rect 2612 22240 3148 22280
rect 3188 22240 3197 22280
rect 2851 22072 2860 22112
rect 2900 22072 3148 22112
rect 3188 22072 3197 22112
rect 3907 22072 3916 22112
rect 3956 22072 4300 22112
rect 4340 22072 4349 22112
rect 3679 21904 3688 21944
rect 3728 21904 3770 21944
rect 3810 21904 3852 21944
rect 3892 21904 3934 21944
rect 3974 21904 4016 21944
rect 4056 21904 4065 21944
rect 7843 21652 7852 21692
rect 7892 21652 9388 21692
rect 9428 21652 9437 21692
rect 4963 21484 4972 21524
rect 5012 21484 5356 21524
rect 5396 21484 6604 21524
rect 6644 21484 6653 21524
rect 5155 21316 5164 21356
rect 5204 21316 5396 21356
rect 11011 21316 11020 21356
rect 11060 21316 11308 21356
rect 11348 21316 11357 21356
rect 12259 21316 12268 21356
rect 12308 21316 12556 21356
rect 12596 21316 12605 21356
rect 4919 21148 4928 21188
rect 4968 21148 5010 21188
rect 5050 21148 5092 21188
rect 5132 21148 5174 21188
rect 5214 21148 5256 21188
rect 5296 21148 5305 21188
rect 5356 21104 5396 21316
rect 4972 21064 5396 21104
rect 4972 21020 5012 21064
rect 4963 20980 4972 21020
rect 5012 20980 5021 21020
rect 5251 20980 5260 21020
rect 5300 20980 5452 21020
rect 5492 20980 5501 21020
rect 5635 20980 5644 21020
rect 5684 20980 5693 21020
rect 5059 20896 5068 20936
rect 5108 20896 5356 20936
rect 5396 20896 5405 20936
rect 5644 20852 5684 20980
rect 4483 20812 4492 20852
rect 4532 20812 8428 20852
rect 8468 20812 8477 20852
rect 3679 20392 3688 20432
rect 3728 20392 3770 20432
rect 3810 20392 3852 20432
rect 3892 20392 3934 20432
rect 3974 20392 4016 20432
rect 4056 20392 4065 20432
rect 2659 20224 2668 20264
rect 2708 20224 3148 20264
rect 3188 20224 3197 20264
rect 3619 20224 3628 20264
rect 3668 20224 4492 20264
rect 4532 20224 4541 20264
rect 2957 20140 3052 20180
rect 3092 20140 3101 20180
rect 4589 20140 4684 20180
rect 4724 20140 4733 20180
rect 13517 20140 13612 20180
rect 13652 20140 13661 20180
rect 11875 19888 11884 19928
rect 11924 19888 12460 19928
rect 12500 19888 12509 19928
rect 4387 19804 4396 19844
rect 4436 19804 5068 19844
rect 5108 19804 5117 19844
rect 4919 19636 4928 19676
rect 4968 19636 5010 19676
rect 5050 19636 5092 19676
rect 5132 19636 5174 19676
rect 5214 19636 5256 19676
rect 5296 19636 5305 19676
rect 5539 19300 5548 19340
rect 5588 19300 5644 19340
rect 5684 19300 5693 19340
rect 10435 19216 10444 19256
rect 10484 19216 11252 19256
rect 11212 19172 11252 19216
rect 4483 19132 4492 19172
rect 4532 19132 4588 19172
rect 4628 19132 4637 19172
rect 11203 19132 11212 19172
rect 11252 19132 11261 19172
rect 3523 19048 3532 19088
rect 3572 19048 3628 19088
rect 3668 19048 3677 19088
rect 12451 19048 12460 19088
rect 12500 19048 12748 19088
rect 12788 19048 12797 19088
rect 3679 18880 3688 18920
rect 3728 18880 3770 18920
rect 3810 18880 3852 18920
rect 3892 18880 3934 18920
rect 3974 18880 4016 18920
rect 4056 18880 4065 18920
rect 9763 18628 9772 18668
rect 9812 18628 11884 18668
rect 11924 18628 11933 18668
rect 13027 18628 13036 18668
rect 13076 18628 13324 18668
rect 13364 18628 13373 18668
rect 12931 18544 12940 18584
rect 12980 18544 13612 18584
rect 13652 18544 13661 18584
rect 10147 18376 10156 18416
rect 10196 18376 10348 18416
rect 10388 18376 10397 18416
rect 13325 18376 13420 18416
rect 13460 18376 13469 18416
rect 11491 18292 11500 18332
rect 11540 18292 12268 18332
rect 12308 18292 12317 18332
rect 5827 18208 5836 18248
rect 5876 18208 6796 18248
rect 6836 18208 6845 18248
rect 10915 18208 10924 18248
rect 10964 18208 12076 18248
rect 12116 18208 12125 18248
rect 4919 18124 4928 18164
rect 4968 18124 5010 18164
rect 5050 18124 5092 18164
rect 5132 18124 5174 18164
rect 5214 18124 5256 18164
rect 5296 18124 5305 18164
rect 3715 18040 3724 18080
rect 3764 18040 4204 18080
rect 4244 18040 7660 18080
rect 7700 18040 7709 18080
rect 4876 17996 4916 18040
rect 4867 17956 4876 17996
rect 4916 17956 4956 17996
rect 5932 17956 6220 17996
rect 6260 17956 6269 17996
rect 6595 17956 6604 17996
rect 6644 17956 6988 17996
rect 7028 17956 7037 17996
rect 7181 17956 7276 17996
rect 7316 17956 7325 17996
rect 9955 17956 9964 17996
rect 10004 17956 11116 17996
rect 11156 17956 11165 17996
rect 12355 17956 12364 17996
rect 12404 17956 12652 17996
rect 12692 17956 12701 17996
rect 5932 17912 5972 17956
rect 5923 17872 5932 17912
rect 5972 17872 5981 17912
rect 6115 17872 6124 17912
rect 6164 17872 6892 17912
rect 6932 17872 6941 17912
rect 9379 17872 9388 17912
rect 9428 17872 9772 17912
rect 9812 17872 9821 17912
rect 6211 17788 6220 17828
rect 6260 17788 6412 17828
rect 6452 17788 6461 17828
rect 6115 17704 6124 17744
rect 6164 17704 6700 17744
rect 6740 17704 6749 17744
rect 4387 17620 4396 17660
rect 4436 17620 5260 17660
rect 5300 17620 9484 17660
rect 9524 17620 9533 17660
rect 2947 17536 2956 17576
rect 2996 17536 3148 17576
rect 3188 17536 3197 17576
rect 4963 17452 4972 17492
rect 5012 17452 7276 17492
rect 7316 17452 7325 17492
rect 11683 17452 11692 17492
rect 11732 17452 13612 17492
rect 13652 17452 13661 17492
rect 2659 17368 2668 17408
rect 2708 17368 2956 17408
rect 2996 17368 3005 17408
rect 3679 17368 3688 17408
rect 3728 17368 3770 17408
rect 3810 17368 3852 17408
rect 3892 17368 3934 17408
rect 3974 17368 4016 17408
rect 4056 17368 4065 17408
rect 4195 17284 4204 17324
rect 4244 17284 7756 17324
rect 7796 17284 7805 17324
rect 11885 17284 11980 17324
rect 12020 17284 12029 17324
rect 5155 17200 5164 17240
rect 5204 17200 5836 17240
rect 5876 17200 5885 17240
rect 6893 17200 6988 17240
rect 7028 17200 7037 17240
rect 7363 17200 7372 17240
rect 7412 17200 9964 17240
rect 10004 17200 10013 17240
rect 10531 17200 10540 17240
rect 10580 17200 13420 17240
rect 13460 17200 13469 17240
rect 11587 17116 11596 17156
rect 11636 17116 11884 17156
rect 11924 17116 11933 17156
rect 5539 17032 5548 17072
rect 5588 17032 5597 17072
rect 5827 17032 5836 17072
rect 5876 17032 6028 17072
rect 6068 17032 6077 17072
rect 7459 17032 7468 17072
rect 7508 17032 7852 17072
rect 7892 17032 7901 17072
rect 11779 17032 11788 17072
rect 11828 17032 12172 17072
rect 12212 17032 12221 17072
rect 4493 16948 4588 16988
rect 4628 16948 4637 16988
rect 5548 16904 5588 17032
rect 5635 16948 5644 16988
rect 5684 16948 5693 16988
rect 5539 16864 5548 16904
rect 5588 16864 5597 16904
rect 4963 16780 4972 16820
rect 5012 16780 5021 16820
rect 4972 16736 5012 16780
rect 4972 16696 5588 16736
rect 4919 16612 4928 16652
rect 4968 16612 5010 16652
rect 5050 16612 5092 16652
rect 5132 16612 5174 16652
rect 5214 16612 5256 16652
rect 5296 16612 5305 16652
rect 5548 16568 5588 16696
rect 5644 16652 5684 16948
rect 5933 16864 6028 16904
rect 6068 16864 6077 16904
rect 10723 16864 10732 16904
rect 10772 16864 11500 16904
rect 11540 16864 11549 16904
rect 10915 16780 10924 16820
rect 10964 16780 11308 16820
rect 11348 16780 11357 16820
rect 5923 16696 5932 16736
rect 5972 16696 6316 16736
rect 6356 16696 6365 16736
rect 10723 16696 10732 16736
rect 10772 16696 11212 16736
rect 11252 16696 11261 16736
rect 5644 16612 8524 16652
rect 8564 16612 8573 16652
rect 5548 16528 6028 16568
rect 6068 16528 6077 16568
rect 11980 16360 12844 16400
rect 12884 16360 12893 16400
rect 11980 16316 12020 16360
rect 6797 16276 6892 16316
rect 6932 16276 6941 16316
rect 11971 16276 11980 16316
rect 12020 16276 12029 16316
rect 5251 16192 5260 16232
rect 5300 16192 7180 16232
rect 7220 16192 7276 16232
rect 7316 16192 8140 16232
rect 8180 16192 8189 16232
rect 6499 16024 6508 16064
rect 6548 16024 6892 16064
rect 6932 16024 6941 16064
rect 7075 16024 7084 16064
rect 7124 16024 8140 16064
rect 8180 16024 8189 16064
rect 11501 16024 11596 16064
rect 11636 16024 11645 16064
rect 1603 15940 1612 15980
rect 1652 15940 1996 15980
rect 2036 15940 2045 15980
rect 2659 15940 2668 15980
rect 2708 15940 6700 15980
rect 6740 15940 6749 15980
rect 10723 15940 10732 15980
rect 10772 15940 10924 15980
rect 10964 15940 10973 15980
rect 3679 15856 3688 15896
rect 3728 15856 3770 15896
rect 3810 15856 3852 15896
rect 3892 15856 3934 15896
rect 3974 15856 4016 15896
rect 4056 15856 4065 15896
rect 5731 15856 5740 15896
rect 5780 15856 9140 15896
rect 4003 15688 4012 15728
rect 4052 15688 4588 15728
rect 4628 15688 4637 15728
rect 8333 15688 8428 15728
rect 8468 15688 8477 15728
rect 9100 15560 9140 15856
rect 9091 15520 9100 15560
rect 9140 15520 9149 15560
rect 2563 15184 2572 15224
rect 2612 15184 7316 15224
rect 7276 15140 7316 15184
rect 3427 15100 3436 15140
rect 3476 15100 3532 15140
rect 3572 15100 3581 15140
rect 4919 15100 4928 15140
rect 4968 15100 5010 15140
rect 5050 15100 5092 15140
rect 5132 15100 5174 15140
rect 5214 15100 5256 15140
rect 5296 15100 5305 15140
rect 7267 15100 7276 15140
rect 7316 15100 7325 15140
rect 2851 15016 2860 15056
rect 2900 15016 3148 15056
rect 3188 15016 3197 15056
rect 4387 15016 4396 15056
rect 4436 15016 4445 15056
rect 5731 15016 5740 15056
rect 5780 15016 7372 15056
rect 7412 15016 7421 15056
rect 4396 14972 4436 15016
rect 4396 14932 5260 14972
rect 5300 14932 5309 14972
rect 3053 14848 3148 14888
rect 3188 14848 3197 14888
rect 3619 14848 3628 14888
rect 3668 14848 4396 14888
rect 4436 14848 4445 14888
rect 5635 14848 5644 14888
rect 5684 14848 7948 14888
rect 7988 14848 7997 14888
rect 13027 14848 13036 14888
rect 13076 14848 13612 14888
rect 13652 14848 13661 14888
rect 4483 14764 4492 14804
rect 4532 14764 5452 14804
rect 5492 14764 5501 14804
rect 6221 14764 6316 14804
rect 6356 14764 6365 14804
rect 4003 14680 4012 14720
rect 4052 14680 4300 14720
rect 4340 14680 4349 14720
rect 5923 14680 5932 14720
rect 5972 14680 6508 14720
rect 6548 14680 6557 14720
rect 7075 14680 7084 14720
rect 7124 14680 7468 14720
rect 7508 14680 7517 14720
rect 10723 14680 10732 14720
rect 10772 14680 10868 14720
rect 3715 14596 3724 14636
rect 3764 14596 4780 14636
rect 4820 14596 4829 14636
rect 7555 14596 7564 14636
rect 7604 14596 7852 14636
rect 7892 14596 7901 14636
rect 5059 14512 5068 14552
rect 5108 14512 8236 14552
rect 8276 14512 8285 14552
rect 9571 14512 9580 14552
rect 9620 14512 10732 14552
rect 10772 14512 10781 14552
rect 10828 14468 10868 14680
rect 5731 14428 5740 14468
rect 5780 14428 8428 14468
rect 8468 14428 8477 14468
rect 9763 14428 9772 14468
rect 9812 14428 10156 14468
rect 10196 14428 10205 14468
rect 10732 14428 10868 14468
rect 3679 14344 3688 14384
rect 3728 14344 3770 14384
rect 3810 14344 3852 14384
rect 3892 14344 3934 14384
rect 3974 14344 4016 14384
rect 4056 14344 4065 14384
rect 4291 14344 4300 14384
rect 4340 14344 4396 14384
rect 4436 14344 4445 14384
rect 10732 14300 10772 14428
rect 8333 14260 8428 14300
rect 8468 14260 8477 14300
rect 10723 14260 10732 14300
rect 10772 14260 10781 14300
rect 8621 14176 8716 14216
rect 8756 14176 8765 14216
rect 10445 14176 10540 14216
rect 10580 14176 10589 14216
rect 4291 14008 4300 14048
rect 4340 14008 4492 14048
rect 4532 14008 4541 14048
rect 5251 14008 5260 14048
rect 5300 14008 5452 14048
rect 5492 14008 5501 14048
rect 1891 13840 1900 13880
rect 1940 13840 8620 13880
rect 8660 13840 8669 13880
rect 11779 13840 11788 13880
rect 11828 13840 12652 13880
rect 12692 13840 12701 13880
rect 3043 13756 3052 13796
rect 3092 13756 3244 13796
rect 3284 13756 3293 13796
rect 4771 13756 4780 13796
rect 4820 13756 5164 13796
rect 5204 13756 5213 13796
rect 6883 13756 6892 13796
rect 6932 13756 7180 13796
rect 7220 13756 7229 13796
rect 4919 13588 4928 13628
rect 4968 13588 5010 13628
rect 5050 13588 5092 13628
rect 5132 13588 5174 13628
rect 5214 13588 5256 13628
rect 5296 13588 5305 13628
rect 8131 13504 8140 13544
rect 8180 13504 8428 13544
rect 8468 13504 8477 13544
rect 4963 13420 4972 13460
rect 5012 13420 5836 13460
rect 5876 13420 5885 13460
rect 9091 13336 9100 13376
rect 9140 13336 9484 13376
rect 9524 13336 9533 13376
rect 4003 13252 4012 13292
rect 4052 13252 4204 13292
rect 4244 13252 4253 13292
rect 5347 13252 5356 13292
rect 5396 13252 5548 13292
rect 5588 13252 5597 13292
rect 5923 13252 5932 13292
rect 5972 13252 6412 13292
rect 6452 13252 6461 13292
rect 4397 13168 4492 13208
rect 4532 13168 4541 13208
rect 5251 13168 5260 13208
rect 5300 13168 5836 13208
rect 5876 13168 5885 13208
rect 4291 13084 4300 13124
rect 4340 13084 4588 13124
rect 4628 13084 4637 13124
rect 7075 13084 7084 13124
rect 7124 13084 7276 13124
rect 7316 13084 7325 13124
rect 2659 13000 2668 13040
rect 2708 13000 2860 13040
rect 2900 13000 2909 13040
rect 8717 13000 8812 13040
rect 8852 13000 8861 13040
rect 7171 12956 7180 12980
rect 2467 12916 2476 12956
rect 2516 12916 2764 12956
rect 2804 12916 2813 12956
rect 6019 12916 6028 12956
rect 6068 12916 6124 12956
rect 6164 12916 6173 12956
rect 6797 12916 6892 12956
rect 6932 12916 6941 12956
rect 7084 12940 7180 12956
rect 7220 12940 7229 12980
rect 7084 12916 7220 12940
rect 7363 12916 7372 12956
rect 7412 12916 8140 12956
rect 8180 12916 8189 12956
rect 3679 12832 3688 12872
rect 3728 12832 3770 12872
rect 3810 12832 3852 12872
rect 3892 12832 3934 12872
rect 3974 12832 4016 12872
rect 4056 12832 4065 12872
rect 7084 12788 7124 12916
rect 7171 12832 7180 12872
rect 7220 12832 7276 12872
rect 7316 12832 7325 12872
rect 7084 12748 7220 12788
rect 8611 12748 8620 12788
rect 8660 12748 8812 12788
rect 8852 12748 8861 12788
rect 9475 12748 9484 12788
rect 9524 12748 9964 12788
rect 10004 12748 10013 12788
rect 4963 12580 4972 12620
rect 5012 12580 5740 12620
rect 5780 12580 5789 12620
rect 3811 12496 3820 12536
rect 3860 12496 4204 12536
rect 4244 12496 5108 12536
rect 5068 12452 5108 12496
rect 7180 12452 7220 12748
rect 7267 12664 7276 12704
rect 7316 12664 7468 12704
rect 7508 12664 7517 12704
rect 9485 12664 9580 12704
rect 9620 12664 9629 12704
rect 5068 12412 6124 12452
rect 6164 12412 6173 12452
rect 7171 12412 7180 12452
rect 7220 12412 7229 12452
rect 5731 12328 5740 12368
rect 5780 12328 6124 12368
rect 6164 12328 6173 12368
rect 6307 12328 6316 12368
rect 6356 12328 7468 12368
rect 7508 12328 7660 12368
rect 7700 12328 7709 12368
rect 4387 12244 4396 12284
rect 4436 12244 4588 12284
rect 4628 12244 4637 12284
rect 4919 12076 4928 12116
rect 4968 12076 5010 12116
rect 5050 12076 5092 12116
rect 5132 12076 5174 12116
rect 5214 12076 5256 12116
rect 5296 12076 5305 12116
rect 7949 11908 8044 11948
rect 8084 11908 8093 11948
rect 11405 11908 11500 11948
rect 11540 11908 11549 11948
rect 4301 11740 4396 11780
rect 4436 11740 4445 11780
rect 6221 11740 6316 11780
rect 6356 11740 6365 11780
rect 4387 11572 4396 11612
rect 4436 11572 5740 11612
rect 5780 11572 5789 11612
rect 9379 11572 9388 11612
rect 9428 11572 11404 11612
rect 11444 11572 11453 11612
rect 3679 11320 3688 11360
rect 3728 11320 3770 11360
rect 3810 11320 3852 11360
rect 3892 11320 3934 11360
rect 3974 11320 4016 11360
rect 4056 11320 4065 11360
rect 1411 10984 1420 11024
rect 1460 10984 1708 11024
rect 1748 10984 1757 11024
rect 4291 10732 4300 10772
rect 4340 10732 4396 10772
rect 4436 10732 4445 10772
rect 6307 10648 6316 10688
rect 6356 10648 6892 10688
rect 6932 10648 6941 10688
rect 7843 10648 7852 10688
rect 7892 10648 8428 10688
rect 8468 10648 8477 10688
rect 4919 10564 4928 10604
rect 4968 10564 5010 10604
rect 5050 10564 5092 10604
rect 5132 10564 5174 10604
rect 5214 10564 5256 10604
rect 5296 10564 5305 10604
rect 6211 10480 6220 10520
rect 6260 10480 6316 10520
rect 6356 10480 6365 10520
rect 6211 10060 6220 10100
rect 6260 10060 6700 10100
rect 6740 10060 6796 10100
rect 6836 10060 6845 10100
rect 6307 9976 6316 10016
rect 6356 9976 6508 10016
rect 6548 9976 6557 10016
rect 2755 9808 2764 9848
rect 2804 9808 3052 9848
rect 3092 9808 3101 9848
rect 3679 9808 3688 9848
rect 3728 9808 3770 9848
rect 3810 9808 3852 9848
rect 3892 9808 3934 9848
rect 3974 9808 4016 9848
rect 4056 9808 4065 9848
rect 11011 9640 11020 9680
rect 11060 9640 11788 9680
rect 11828 9640 11837 9680
rect 4579 9556 4588 9596
rect 4628 9556 4637 9596
rect 4588 9344 4628 9556
rect 5453 9472 5548 9512
rect 5588 9472 6604 9512
rect 6644 9472 9388 9512
rect 9428 9472 9437 9512
rect 5827 9388 5836 9428
rect 5876 9388 6988 9428
rect 7028 9388 7037 9428
rect 4588 9304 5644 9344
rect 5684 9304 5693 9344
rect 4919 9052 4928 9092
rect 4968 9052 5010 9092
rect 5050 9052 5092 9092
rect 5132 9052 5174 9092
rect 5214 9052 5256 9092
rect 5296 9052 5305 9092
rect 1603 8968 1612 9008
rect 1652 8968 5740 9008
rect 5780 8968 5789 9008
rect 6211 8800 6220 8840
rect 6260 8800 6796 8840
rect 6836 8800 6845 8840
rect 7171 8800 7180 8840
rect 7220 8800 8524 8840
rect 8564 8800 8573 8840
rect 5059 8716 5068 8756
rect 5108 8716 5452 8756
rect 5492 8716 5740 8756
rect 5780 8716 5789 8756
rect 6787 8632 6796 8672
rect 6836 8632 6988 8672
rect 7028 8632 7037 8672
rect 7171 8632 7180 8672
rect 7220 8632 12172 8672
rect 12212 8632 12221 8672
rect 3679 8296 3688 8336
rect 3728 8296 3770 8336
rect 3810 8296 3852 8336
rect 3892 8296 3934 8336
rect 3974 8296 4016 8336
rect 4056 8296 4065 8336
rect 8429 8128 8524 8168
rect 8564 8128 8573 8168
rect 1411 7960 1420 8000
rect 1460 7960 1516 8000
rect 1556 7960 1565 8000
rect 7363 7960 7372 8000
rect 7412 7960 12268 8000
rect 12308 7960 12317 8000
rect 8035 7876 8044 7916
rect 8084 7876 9484 7916
rect 9524 7876 9533 7916
rect 5443 7708 5452 7748
rect 5492 7708 5740 7748
rect 5780 7708 5789 7748
rect 4919 7540 4928 7580
rect 4968 7540 5010 7580
rect 5050 7540 5092 7580
rect 5132 7540 5174 7580
rect 5214 7540 5256 7580
rect 5296 7540 5305 7580
rect 8515 7540 8524 7580
rect 8564 7540 9292 7580
rect 9332 7540 9341 7580
rect 4771 7204 4780 7244
rect 4820 7204 4876 7244
rect 4916 7204 4925 7244
rect 1325 7120 1420 7160
rect 1460 7120 1469 7160
rect 4963 7120 4972 7160
rect 5012 7120 6508 7160
rect 6548 7120 6557 7160
rect 3679 6784 3688 6824
rect 3728 6784 3770 6824
rect 3810 6784 3852 6824
rect 3892 6784 3934 6824
rect 3974 6784 4016 6824
rect 4056 6784 4065 6824
rect 7469 6364 7564 6404
rect 7604 6364 7613 6404
rect 4919 6028 4928 6068
rect 4968 6028 5010 6068
rect 5050 6028 5092 6068
rect 5132 6028 5174 6068
rect 5214 6028 5256 6068
rect 5296 6028 5305 6068
rect 10253 5608 10348 5648
rect 10388 5608 10397 5648
rect 3679 5272 3688 5312
rect 3728 5272 3770 5312
rect 3810 5272 3852 5312
rect 3892 5272 3934 5312
rect 3974 5272 4016 5312
rect 4056 5272 4065 5312
rect 9869 4936 9964 4976
rect 10004 4936 10013 4976
rect 4919 4516 4928 4556
rect 4968 4516 5010 4556
rect 5050 4516 5092 4556
rect 5132 4516 5174 4556
rect 5214 4516 5256 4556
rect 5296 4516 5305 4556
rect 3341 4264 3436 4304
rect 3476 4264 3485 4304
rect 10435 4264 10444 4304
rect 10484 4264 12556 4304
rect 12596 4264 12605 4304
rect 3679 3760 3688 3800
rect 3728 3760 3770 3800
rect 3810 3760 3852 3800
rect 3892 3760 3934 3800
rect 3974 3760 4016 3800
rect 4056 3760 4065 3800
rect 4919 3004 4928 3044
rect 4968 3004 5010 3044
rect 5050 3004 5092 3044
rect 5132 3004 5174 3044
rect 5214 3004 5256 3044
rect 5296 3004 5305 3044
rect 8141 2836 8236 2876
rect 8276 2836 8285 2876
rect 5731 2416 5740 2456
rect 5780 2416 11884 2456
rect 11924 2416 11933 2456
rect 3679 2248 3688 2288
rect 3728 2248 3770 2288
rect 3810 2248 3852 2288
rect 3892 2248 3934 2288
rect 3974 2248 4016 2288
rect 4056 2248 4065 2288
rect 4919 1492 4928 1532
rect 4968 1492 5010 1532
rect 5050 1492 5092 1532
rect 5132 1492 5174 1532
rect 5214 1492 5256 1532
rect 5296 1492 5305 1532
rect 2669 1408 2764 1448
rect 2804 1408 2813 1448
rect 5549 1408 5644 1448
rect 5684 1408 5693 1448
rect 6125 1408 6220 1448
rect 6260 1408 6269 1448
rect 6787 1240 6796 1280
rect 6836 1240 8908 1280
rect 8948 1240 8957 1280
rect 9005 988 9100 1028
rect 9140 988 9149 1028
rect 9581 988 9676 1028
rect 9716 988 9725 1028
rect 10157 988 10252 1028
rect 10292 988 10301 1028
rect 10733 988 10828 1028
rect 10868 988 10877 1028
rect 11309 988 11404 1028
rect 11444 988 11453 1028
rect 4483 904 4492 944
rect 4532 904 6604 944
rect 6644 904 6653 944
rect 11203 652 11212 692
rect 11252 652 11980 692
rect 12020 652 12029 692
rect 7363 232 7372 272
rect 7412 232 8620 272
rect 8660 232 8669 272
rect 3235 148 3244 188
rect 3284 148 3956 188
rect 5059 148 5068 188
rect 5108 148 6412 188
rect 6452 148 6461 188
rect 3916 104 3956 148
rect 3907 64 3916 104
rect 3956 64 3965 104
<< via4 >>
rect 4928 46852 4968 46892
rect 5010 46852 5050 46892
rect 5092 46852 5132 46892
rect 5174 46852 5214 46892
rect 5256 46852 5296 46892
rect 1900 46432 1940 46472
rect 3688 46096 3728 46136
rect 3770 46096 3810 46136
rect 3852 46096 3892 46136
rect 3934 46096 3974 46136
rect 4016 46096 4056 46136
rect 10828 45760 10868 45800
rect 4928 45340 4968 45380
rect 5010 45340 5050 45380
rect 5092 45340 5132 45380
rect 5174 45340 5214 45380
rect 5256 45340 5296 45380
rect 5644 44920 5684 44960
rect 8908 44920 8948 44960
rect 9292 44920 9332 44960
rect 10252 44836 10292 44876
rect 6412 44752 6452 44792
rect 10636 44668 10676 44708
rect 3688 44584 3728 44624
rect 3770 44584 3810 44624
rect 3852 44584 3892 44624
rect 3934 44584 3974 44624
rect 4016 44584 4056 44624
rect 9484 44248 9524 44288
rect 4928 43828 4968 43868
rect 5010 43828 5050 43868
rect 5092 43828 5132 43868
rect 5174 43828 5214 43868
rect 5256 43828 5296 43868
rect 6604 43660 6644 43700
rect 8620 43408 8660 43448
rect 6796 43324 6836 43364
rect 3688 43072 3728 43112
rect 3770 43072 3810 43112
rect 3852 43072 3892 43112
rect 3934 43072 3974 43112
rect 4016 43072 4056 43112
rect 11212 42736 11252 42776
rect 4928 42316 4968 42356
rect 5010 42316 5050 42356
rect 5092 42316 5132 42356
rect 5174 42316 5214 42356
rect 5256 42316 5296 42356
rect 10444 41896 10484 41936
rect 11404 41812 11444 41852
rect 3688 41560 3728 41600
rect 3770 41560 3810 41600
rect 3852 41560 3892 41600
rect 3934 41560 3974 41600
rect 4016 41560 4056 41600
rect 4928 40804 4968 40844
rect 5010 40804 5050 40844
rect 5092 40804 5132 40844
rect 5174 40804 5214 40844
rect 5256 40804 5296 40844
rect 3436 40300 3476 40340
rect 4588 40300 4628 40340
rect 6508 40300 6548 40340
rect 3688 40048 3728 40088
rect 3770 40048 3810 40088
rect 3852 40048 3892 40088
rect 3934 40048 3974 40088
rect 4016 40048 4056 40088
rect 4928 39292 4968 39332
rect 5010 39292 5050 39332
rect 5092 39292 5132 39332
rect 5174 39292 5214 39332
rect 5256 39292 5296 39332
rect 10924 38956 10964 38996
rect 9772 38872 9812 38912
rect 11116 38872 11156 38912
rect 11884 38872 11924 38912
rect 3688 38536 3728 38576
rect 3770 38536 3810 38576
rect 3852 38536 3892 38576
rect 3934 38536 3974 38576
rect 4016 38536 4056 38576
rect 11020 38200 11060 38240
rect 4928 37780 4968 37820
rect 5010 37780 5050 37820
rect 5092 37780 5132 37820
rect 5174 37780 5214 37820
rect 5256 37780 5296 37820
rect 7180 37444 7220 37484
rect 11980 37360 12020 37400
rect 9100 37276 9140 37316
rect 9580 37192 9620 37232
rect 3688 37024 3728 37064
rect 3770 37024 3810 37064
rect 3852 37024 3892 37064
rect 3934 37024 3974 37064
rect 4016 37024 4056 37064
rect 4928 36268 4968 36308
rect 5010 36268 5050 36308
rect 5092 36268 5132 36308
rect 5174 36268 5214 36308
rect 5256 36268 5296 36308
rect 3688 35512 3728 35552
rect 3770 35512 3810 35552
rect 3852 35512 3892 35552
rect 3934 35512 3974 35552
rect 4016 35512 4056 35552
rect 4928 34756 4968 34796
rect 5010 34756 5050 34796
rect 5092 34756 5132 34796
rect 5174 34756 5214 34796
rect 5256 34756 5296 34796
rect 10348 34336 10388 34376
rect 3688 34000 3728 34040
rect 3770 34000 3810 34040
rect 3852 34000 3892 34040
rect 3934 34000 3974 34040
rect 4016 34000 4056 34040
rect 7276 33664 7316 33704
rect 12076 33664 12116 33704
rect 6124 33328 6164 33368
rect 4928 33244 4968 33284
rect 5010 33244 5050 33284
rect 5092 33244 5132 33284
rect 5174 33244 5214 33284
rect 5256 33244 5296 33284
rect 10540 33076 10580 33116
rect 8044 32824 8084 32864
rect 10732 32656 10772 32696
rect 3688 32488 3728 32528
rect 3770 32488 3810 32528
rect 3852 32488 3892 32528
rect 3934 32488 3974 32528
rect 4016 32488 4056 32528
rect 10540 32488 10580 32528
rect 4928 31732 4968 31772
rect 5010 31732 5050 31772
rect 5092 31732 5132 31772
rect 5174 31732 5214 31772
rect 5256 31732 5296 31772
rect 6316 31732 6356 31772
rect 3688 30976 3728 31016
rect 3770 30976 3810 31016
rect 3852 30976 3892 31016
rect 3934 30976 3974 31016
rect 4016 30976 4056 31016
rect 3436 30724 3476 30764
rect 3436 30556 3476 30596
rect 10156 30556 10196 30596
rect 2764 30388 2804 30428
rect 4300 30220 4340 30260
rect 4492 30220 4532 30260
rect 4684 30220 4724 30260
rect 4928 30220 4968 30260
rect 5010 30220 5050 30260
rect 5092 30220 5132 30260
rect 5174 30220 5214 30260
rect 5256 30220 5296 30260
rect 6220 30220 6260 30260
rect 8524 30220 8564 30260
rect 11596 30136 11636 30176
rect 6124 30052 6164 30092
rect 4684 29968 4724 30008
rect 3532 29716 3572 29756
rect 3340 29632 3380 29672
rect 3688 29464 3728 29504
rect 3770 29464 3810 29504
rect 3852 29464 3892 29504
rect 3934 29464 3974 29504
rect 4016 29464 4056 29504
rect 3052 29212 3092 29252
rect 4300 29044 4340 29084
rect 4684 28876 4724 28916
rect 12844 29044 12884 29084
rect 8716 28792 8756 28832
rect 12076 28792 12116 28832
rect 4928 28708 4968 28748
rect 5010 28708 5050 28748
rect 5092 28708 5132 28748
rect 5174 28708 5214 28748
rect 5256 28708 5296 28748
rect 3688 27952 3728 27992
rect 3770 27952 3810 27992
rect 3852 27952 3892 27992
rect 3934 27952 3974 27992
rect 4016 27952 4056 27992
rect 12844 27868 12884 27908
rect 4780 27532 4820 27572
rect 11596 27532 11636 27572
rect 10540 27364 10580 27404
rect 11692 27364 11732 27404
rect 4928 27196 4968 27236
rect 5010 27196 5050 27236
rect 5092 27196 5132 27236
rect 5174 27196 5214 27236
rect 5256 27196 5296 27236
rect 10540 27196 10580 27236
rect 4684 26776 4724 26816
rect 11308 26692 11348 26732
rect 3688 26440 3728 26480
rect 3770 26440 3810 26480
rect 3852 26440 3892 26480
rect 3934 26440 3974 26480
rect 4016 26440 4056 26480
rect 11692 26440 11732 26480
rect 3052 26020 3092 26060
rect 10540 25936 10580 25976
rect 4928 25684 4968 25724
rect 5010 25684 5050 25724
rect 5092 25684 5132 25724
rect 5174 25684 5214 25724
rect 5256 25684 5296 25724
rect 7564 25432 7604 25472
rect 2668 25348 2708 25388
rect 3532 25348 3572 25388
rect 5740 25180 5780 25220
rect 5548 25096 5588 25136
rect 3688 24928 3728 24968
rect 3770 24928 3810 24968
rect 3852 24928 3892 24968
rect 3934 24928 3974 24968
rect 4016 24928 4056 24968
rect 1420 24592 1460 24632
rect 7468 24508 7508 24548
rect 9676 24340 9716 24380
rect 10636 24340 10676 24380
rect 4928 24172 4968 24212
rect 5010 24172 5050 24212
rect 5092 24172 5132 24212
rect 5174 24172 5214 24212
rect 5256 24172 5296 24212
rect 8236 23752 8276 23792
rect 1516 23500 1556 23540
rect 3688 23416 3728 23456
rect 3770 23416 3810 23456
rect 3852 23416 3892 23456
rect 3934 23416 3974 23456
rect 4016 23416 4056 23456
rect 2956 23164 2996 23204
rect 1708 23080 1748 23120
rect 2860 22996 2900 23036
rect 3340 22996 3380 23036
rect 4300 22996 4340 23036
rect 5452 22996 5492 23036
rect 4928 22660 4968 22700
rect 5010 22660 5050 22700
rect 5092 22660 5132 22700
rect 5174 22660 5214 22700
rect 5256 22660 5296 22700
rect 10540 22660 10580 22700
rect 3148 22072 3188 22112
rect 3688 21904 3728 21944
rect 3770 21904 3810 21944
rect 3852 21904 3892 21944
rect 3934 21904 3974 21944
rect 4016 21904 4056 21944
rect 9388 21652 9428 21692
rect 11308 21316 11348 21356
rect 4928 21148 4968 21188
rect 5010 21148 5050 21188
rect 5092 21148 5132 21188
rect 5174 21148 5214 21188
rect 5256 21148 5296 21188
rect 3688 20392 3728 20432
rect 3770 20392 3810 20432
rect 3852 20392 3892 20432
rect 3934 20392 3974 20432
rect 4016 20392 4056 20432
rect 4492 20224 4532 20264
rect 3052 20140 3092 20180
rect 4684 20140 4724 20180
rect 13612 20140 13652 20180
rect 4396 19804 4436 19844
rect 4928 19636 4968 19676
rect 5010 19636 5050 19676
rect 5092 19636 5132 19676
rect 5174 19636 5214 19676
rect 5256 19636 5296 19676
rect 5548 19300 5588 19340
rect 4492 19132 4532 19172
rect 3532 19048 3572 19088
rect 3688 18880 3728 18920
rect 3770 18880 3810 18920
rect 3852 18880 3892 18920
rect 3934 18880 3974 18920
rect 4016 18880 4056 18920
rect 9772 18628 9812 18668
rect 13420 18376 13460 18416
rect 11500 18292 11540 18332
rect 6796 18208 6836 18248
rect 10924 18208 10964 18248
rect 4928 18124 4968 18164
rect 5010 18124 5050 18164
rect 5092 18124 5132 18164
rect 5174 18124 5214 18164
rect 5256 18124 5296 18164
rect 4204 18040 4244 18080
rect 7276 17956 7316 17996
rect 11116 17956 11156 17996
rect 6892 17872 6932 17912
rect 6124 17704 6164 17744
rect 4396 17620 4436 17660
rect 13612 17452 13652 17492
rect 2668 17368 2708 17408
rect 3688 17368 3728 17408
rect 3770 17368 3810 17408
rect 3852 17368 3892 17408
rect 3934 17368 3974 17408
rect 4016 17368 4056 17408
rect 11980 17284 12020 17324
rect 5836 17200 5876 17240
rect 6988 17200 7028 17240
rect 9964 17200 10004 17240
rect 10540 17200 10580 17240
rect 13420 17200 13460 17240
rect 11596 17116 11636 17156
rect 4588 16948 4628 16988
rect 4928 16612 4968 16652
rect 5010 16612 5050 16652
rect 5092 16612 5132 16652
rect 5174 16612 5214 16652
rect 5256 16612 5296 16652
rect 6028 16864 6068 16904
rect 5932 16696 5972 16736
rect 6892 16276 6932 16316
rect 7276 16192 7316 16232
rect 8140 16192 8180 16232
rect 6892 16024 6932 16064
rect 11596 16024 11636 16064
rect 6700 15940 6740 15980
rect 3688 15856 3728 15896
rect 3770 15856 3810 15896
rect 3852 15856 3892 15896
rect 3934 15856 3974 15896
rect 4016 15856 4056 15896
rect 5740 15856 5780 15896
rect 8428 15688 8468 15728
rect 3532 15100 3572 15140
rect 4928 15100 4968 15140
rect 5010 15100 5050 15140
rect 5092 15100 5132 15140
rect 5174 15100 5214 15140
rect 5256 15100 5296 15140
rect 3148 14848 3188 14888
rect 4396 14848 4436 14888
rect 6316 14764 6356 14804
rect 7468 14680 7508 14720
rect 10732 14512 10772 14552
rect 10156 14428 10196 14468
rect 3688 14344 3728 14384
rect 3770 14344 3810 14384
rect 3852 14344 3892 14384
rect 3934 14344 3974 14384
rect 4016 14344 4056 14384
rect 4300 14344 4340 14384
rect 8428 14260 8468 14300
rect 8716 14176 8756 14216
rect 10540 14176 10580 14216
rect 1900 13840 1940 13880
rect 4780 13756 4820 13796
rect 6892 13756 6932 13796
rect 4928 13588 4968 13628
rect 5010 13588 5050 13628
rect 5092 13588 5132 13628
rect 5174 13588 5214 13628
rect 5256 13588 5296 13628
rect 4204 13252 4244 13292
rect 5548 13252 5588 13292
rect 5932 13252 5972 13292
rect 4492 13168 4532 13208
rect 5836 13168 5876 13208
rect 4588 13084 4628 13124
rect 7276 13084 7316 13124
rect 8812 13000 8852 13040
rect 6028 12916 6068 12956
rect 6892 12916 6932 12956
rect 8140 12916 8180 12956
rect 3688 12832 3728 12872
rect 3770 12832 3810 12872
rect 3852 12832 3892 12872
rect 3934 12832 3974 12872
rect 4016 12832 4056 12872
rect 7276 12832 7316 12872
rect 8812 12748 8852 12788
rect 4204 12496 4244 12536
rect 9580 12664 9620 12704
rect 6124 12328 6164 12368
rect 6316 12328 6356 12368
rect 4396 12244 4436 12284
rect 4928 12076 4968 12116
rect 5010 12076 5050 12116
rect 5092 12076 5132 12116
rect 5174 12076 5214 12116
rect 5256 12076 5296 12116
rect 8044 11908 8084 11948
rect 11500 11908 11540 11948
rect 4396 11740 4436 11780
rect 6316 11740 6356 11780
rect 9388 11572 9428 11612
rect 3688 11320 3728 11360
rect 3770 11320 3810 11360
rect 3852 11320 3892 11360
rect 3934 11320 3974 11360
rect 4016 11320 4056 11360
rect 1708 10984 1748 11024
rect 4396 10732 4436 10772
rect 6892 10648 6932 10688
rect 4928 10564 4968 10604
rect 5010 10564 5050 10604
rect 5092 10564 5132 10604
rect 5174 10564 5214 10604
rect 5256 10564 5296 10604
rect 6316 10480 6356 10520
rect 6796 10060 6836 10100
rect 6316 9976 6356 10016
rect 3688 9808 3728 9848
rect 3770 9808 3810 9848
rect 3852 9808 3892 9848
rect 3934 9808 3974 9848
rect 4016 9808 4056 9848
rect 11020 9640 11060 9680
rect 5548 9472 5588 9512
rect 5836 9388 5876 9428
rect 4928 9052 4968 9092
rect 5010 9052 5050 9092
rect 5092 9052 5132 9092
rect 5174 9052 5214 9092
rect 5256 9052 5296 9092
rect 6988 8632 7028 8672
rect 7180 8632 7220 8672
rect 3688 8296 3728 8336
rect 3770 8296 3810 8336
rect 3852 8296 3892 8336
rect 3934 8296 3974 8336
rect 4016 8296 4056 8336
rect 8524 8128 8564 8168
rect 1516 7960 1556 8000
rect 7372 7960 7412 8000
rect 9484 7876 9524 7916
rect 5452 7708 5492 7748
rect 4928 7540 4968 7580
rect 5010 7540 5050 7580
rect 5092 7540 5132 7580
rect 5174 7540 5214 7580
rect 5256 7540 5296 7580
rect 9292 7540 9332 7580
rect 4780 7204 4820 7244
rect 1420 7120 1460 7160
rect 6508 7120 6548 7160
rect 3688 6784 3728 6824
rect 3770 6784 3810 6824
rect 3852 6784 3892 6824
rect 3934 6784 3974 6824
rect 4016 6784 4056 6824
rect 7564 6364 7604 6404
rect 4928 6028 4968 6068
rect 5010 6028 5050 6068
rect 5092 6028 5132 6068
rect 5174 6028 5214 6068
rect 5256 6028 5296 6068
rect 10348 5608 10388 5648
rect 3688 5272 3728 5312
rect 3770 5272 3810 5312
rect 3852 5272 3892 5312
rect 3934 5272 3974 5312
rect 4016 5272 4056 5312
rect 9964 4936 10004 4976
rect 4928 4516 4968 4556
rect 5010 4516 5050 4556
rect 5092 4516 5132 4556
rect 5174 4516 5214 4556
rect 5256 4516 5296 4556
rect 3436 4264 3476 4304
rect 10444 4264 10484 4304
rect 3688 3760 3728 3800
rect 3770 3760 3810 3800
rect 3852 3760 3892 3800
rect 3934 3760 3974 3800
rect 4016 3760 4056 3800
rect 4928 3004 4968 3044
rect 5010 3004 5050 3044
rect 5092 3004 5132 3044
rect 5174 3004 5214 3044
rect 5256 3004 5296 3044
rect 8236 2836 8276 2876
rect 11884 2416 11924 2456
rect 3688 2248 3728 2288
rect 3770 2248 3810 2288
rect 3852 2248 3892 2288
rect 3934 2248 3974 2288
rect 4016 2248 4056 2288
rect 4928 1492 4968 1532
rect 5010 1492 5050 1532
rect 5092 1492 5132 1532
rect 5174 1492 5214 1532
rect 5256 1492 5296 1532
rect 2764 1408 2804 1448
rect 5644 1408 5684 1448
rect 6220 1408 6260 1448
rect 8908 1240 8948 1280
rect 9100 988 9140 1028
rect 9676 988 9716 1028
rect 10252 988 10292 1028
rect 10828 988 10868 1028
rect 11404 988 11444 1028
rect 6604 904 6644 944
rect 11212 652 11252 692
rect 8620 232 8660 272
rect 6412 148 6452 188
<< metal5 >>
rect 1900 46472 1940 46481
rect 1420 24632 1460 24641
rect 1420 7160 1460 24592
rect 1516 23540 1556 23549
rect 1516 8000 1556 23500
rect 1708 23120 1748 23129
rect 1708 11024 1748 23080
rect 1900 13880 1940 46432
rect 3652 46136 4092 48384
rect 3652 46096 3688 46136
rect 3728 46096 3770 46136
rect 3810 46096 3852 46136
rect 3892 46096 3934 46136
rect 3974 46096 4016 46136
rect 4056 46096 4092 46136
rect 3652 44624 4092 46096
rect 3652 44584 3688 44624
rect 3728 44584 3770 44624
rect 3810 44584 3852 44624
rect 3892 44584 3934 44624
rect 3974 44584 4016 44624
rect 4056 44584 4092 44624
rect 3652 43112 4092 44584
rect 3652 43072 3688 43112
rect 3728 43072 3770 43112
rect 3810 43072 3852 43112
rect 3892 43072 3934 43112
rect 3974 43072 4016 43112
rect 4056 43072 4092 43112
rect 3652 41600 4092 43072
rect 3652 41560 3688 41600
rect 3728 41560 3770 41600
rect 3810 41560 3852 41600
rect 3892 41560 3934 41600
rect 3974 41560 4016 41600
rect 4056 41560 4092 41600
rect 3436 40340 3476 40349
rect 3436 30764 3476 40300
rect 3436 30715 3476 30724
rect 3652 40088 4092 41560
rect 4892 46892 5332 48384
rect 4892 46852 4928 46892
rect 4968 46852 5010 46892
rect 5050 46852 5092 46892
rect 5132 46852 5174 46892
rect 5214 46852 5256 46892
rect 5296 46852 5332 46892
rect 4892 45380 5332 46852
rect 4892 45340 4928 45380
rect 4968 45340 5010 45380
rect 5050 45340 5092 45380
rect 5132 45340 5174 45380
rect 5214 45340 5256 45380
rect 5296 45340 5332 45380
rect 4892 43868 5332 45340
rect 10828 45800 10868 45809
rect 4892 43828 4928 43868
rect 4968 43828 5010 43868
rect 5050 43828 5092 43868
rect 5132 43828 5174 43868
rect 5214 43828 5256 43868
rect 5296 43828 5332 43868
rect 4892 42356 5332 43828
rect 4892 42316 4928 42356
rect 4968 42316 5010 42356
rect 5050 42316 5092 42356
rect 5132 42316 5174 42356
rect 5214 42316 5256 42356
rect 5296 42316 5332 42356
rect 4892 40844 5332 42316
rect 4892 40804 4928 40844
rect 4968 40804 5010 40844
rect 5050 40804 5092 40844
rect 5132 40804 5174 40844
rect 5214 40804 5256 40844
rect 5296 40804 5332 40844
rect 3652 40048 3688 40088
rect 3728 40048 3770 40088
rect 3810 40048 3852 40088
rect 3892 40048 3934 40088
rect 3974 40048 4016 40088
rect 4056 40048 4092 40088
rect 3652 38576 4092 40048
rect 4588 40340 4628 40349
rect 4588 38900 4628 40300
rect 4892 39332 5332 40804
rect 4892 39292 4928 39332
rect 4968 39292 5010 39332
rect 5050 39292 5092 39332
rect 5132 39292 5174 39332
rect 5214 39292 5256 39332
rect 5296 39292 5332 39332
rect 4588 38860 4820 38900
rect 3652 38536 3688 38576
rect 3728 38536 3770 38576
rect 3810 38536 3852 38576
rect 3892 38536 3934 38576
rect 3974 38536 4016 38576
rect 4056 38536 4092 38576
rect 3652 37064 4092 38536
rect 3652 37024 3688 37064
rect 3728 37024 3770 37064
rect 3810 37024 3852 37064
rect 3892 37024 3934 37064
rect 3974 37024 4016 37064
rect 4056 37024 4092 37064
rect 3652 35552 4092 37024
rect 3652 35512 3688 35552
rect 3728 35512 3770 35552
rect 3810 35512 3852 35552
rect 3892 35512 3934 35552
rect 3974 35512 4016 35552
rect 4056 35512 4092 35552
rect 3652 34040 4092 35512
rect 3652 34000 3688 34040
rect 3728 34000 3770 34040
rect 3810 34000 3852 34040
rect 3892 34000 3934 34040
rect 3974 34000 4016 34040
rect 4056 34000 4092 34040
rect 3652 32528 4092 34000
rect 3652 32488 3688 32528
rect 3728 32488 3770 32528
rect 3810 32488 3852 32528
rect 3892 32488 3934 32528
rect 3974 32488 4016 32528
rect 4056 32488 4092 32528
rect 3652 31016 4092 32488
rect 3652 30976 3688 31016
rect 3728 30976 3770 31016
rect 3810 30976 3852 31016
rect 3892 30976 3934 31016
rect 3974 30976 4016 31016
rect 4056 30976 4092 31016
rect 3436 30596 3476 30605
rect 2764 30428 2804 30437
rect 2668 25388 2708 25397
rect 2668 17408 2708 25348
rect 2668 17359 2708 17368
rect 1900 13831 1940 13840
rect 1708 10975 1748 10984
rect 1516 7951 1556 7960
rect 1420 7111 1460 7120
rect 2764 1448 2804 30388
rect 3340 29672 3380 29681
rect 3052 29252 3092 29261
rect 3052 26060 3092 29212
rect 2956 23204 2996 23213
rect 2956 23060 2996 23164
rect 2860 23036 2996 23060
rect 2900 23020 2996 23036
rect 2860 22987 2900 22996
rect 3052 20180 3092 26020
rect 3340 23036 3380 29632
rect 3340 22987 3380 22996
rect 3052 20131 3092 20140
rect 3148 22112 3188 22121
rect 3148 14888 3188 22072
rect 3148 14839 3188 14848
rect 3436 4304 3476 30556
rect 3532 29756 3572 29765
rect 3532 25388 3572 29716
rect 3532 25339 3572 25348
rect 3652 29504 4092 30976
rect 3652 29464 3688 29504
rect 3728 29464 3770 29504
rect 3810 29464 3852 29504
rect 3892 29464 3934 29504
rect 3974 29464 4016 29504
rect 4056 29464 4092 29504
rect 3652 27992 4092 29464
rect 4300 30260 4340 30269
rect 4300 29084 4340 30220
rect 4300 29035 4340 29044
rect 4492 30260 4532 30269
rect 3652 27952 3688 27992
rect 3728 27952 3770 27992
rect 3810 27952 3852 27992
rect 3892 27952 3934 27992
rect 3974 27952 4016 27992
rect 4056 27952 4092 27992
rect 3652 26480 4092 27952
rect 3652 26440 3688 26480
rect 3728 26440 3770 26480
rect 3810 26440 3852 26480
rect 3892 26440 3934 26480
rect 3974 26440 4016 26480
rect 4056 26440 4092 26480
rect 3652 24968 4092 26440
rect 3652 24928 3688 24968
rect 3728 24928 3770 24968
rect 3810 24928 3852 24968
rect 3892 24928 3934 24968
rect 3974 24928 4016 24968
rect 4056 24928 4092 24968
rect 3652 23456 4092 24928
rect 3652 23416 3688 23456
rect 3728 23416 3770 23456
rect 3810 23416 3852 23456
rect 3892 23416 3934 23456
rect 3974 23416 4016 23456
rect 4056 23416 4092 23456
rect 3652 21944 4092 23416
rect 3652 21904 3688 21944
rect 3728 21904 3770 21944
rect 3810 21904 3852 21944
rect 3892 21904 3934 21944
rect 3974 21904 4016 21944
rect 4056 21904 4092 21944
rect 3652 20432 4092 21904
rect 3652 20392 3688 20432
rect 3728 20392 3770 20432
rect 3810 20392 3852 20432
rect 3892 20392 3934 20432
rect 3974 20392 4016 20432
rect 4056 20392 4092 20432
rect 3532 19088 3572 19097
rect 3532 15140 3572 19048
rect 3532 15091 3572 15100
rect 3652 18920 4092 20392
rect 3652 18880 3688 18920
rect 3728 18880 3770 18920
rect 3810 18880 3852 18920
rect 3892 18880 3934 18920
rect 3974 18880 4016 18920
rect 4056 18880 4092 18920
rect 3652 17408 4092 18880
rect 4300 23036 4340 23045
rect 3652 17368 3688 17408
rect 3728 17368 3770 17408
rect 3810 17368 3852 17408
rect 3892 17368 3934 17408
rect 3974 17368 4016 17408
rect 4056 17368 4092 17408
rect 3652 15896 4092 17368
rect 3652 15856 3688 15896
rect 3728 15856 3770 15896
rect 3810 15856 3852 15896
rect 3892 15856 3934 15896
rect 3974 15856 4016 15896
rect 4056 15856 4092 15896
rect 3436 4255 3476 4264
rect 3652 14384 4092 15856
rect 3652 14344 3688 14384
rect 3728 14344 3770 14384
rect 3810 14344 3852 14384
rect 3892 14344 3934 14384
rect 3974 14344 4016 14384
rect 4056 14344 4092 14384
rect 3652 12872 4092 14344
rect 3652 12832 3688 12872
rect 3728 12832 3770 12872
rect 3810 12832 3852 12872
rect 3892 12832 3934 12872
rect 3974 12832 4016 12872
rect 4056 12832 4092 12872
rect 3652 11360 4092 12832
rect 4204 18080 4244 18089
rect 4204 13292 4244 18040
rect 4300 14384 4340 22996
rect 4492 20264 4532 30220
rect 4684 30260 4724 30269
rect 4684 30008 4724 30220
rect 4684 29959 4724 29968
rect 4492 20215 4532 20224
rect 4684 28916 4724 28925
rect 4684 26816 4724 28876
rect 4780 27572 4820 38860
rect 4780 27523 4820 27532
rect 4892 37820 5332 39292
rect 4892 37780 4928 37820
rect 4968 37780 5010 37820
rect 5050 37780 5092 37820
rect 5132 37780 5174 37820
rect 5214 37780 5256 37820
rect 5296 37780 5332 37820
rect 4892 36308 5332 37780
rect 4892 36268 4928 36308
rect 4968 36268 5010 36308
rect 5050 36268 5092 36308
rect 5132 36268 5174 36308
rect 5214 36268 5256 36308
rect 5296 36268 5332 36308
rect 4892 34796 5332 36268
rect 4892 34756 4928 34796
rect 4968 34756 5010 34796
rect 5050 34756 5092 34796
rect 5132 34756 5174 34796
rect 5214 34756 5256 34796
rect 5296 34756 5332 34796
rect 4892 33284 5332 34756
rect 4892 33244 4928 33284
rect 4968 33244 5010 33284
rect 5050 33244 5092 33284
rect 5132 33244 5174 33284
rect 5214 33244 5256 33284
rect 5296 33244 5332 33284
rect 4892 31772 5332 33244
rect 4892 31732 4928 31772
rect 4968 31732 5010 31772
rect 5050 31732 5092 31772
rect 5132 31732 5174 31772
rect 5214 31732 5256 31772
rect 5296 31732 5332 31772
rect 4892 30260 5332 31732
rect 4892 30220 4928 30260
rect 4968 30220 5010 30260
rect 5050 30220 5092 30260
rect 5132 30220 5174 30260
rect 5214 30220 5256 30260
rect 5296 30220 5332 30260
rect 4892 28748 5332 30220
rect 4892 28708 4928 28748
rect 4968 28708 5010 28748
rect 5050 28708 5092 28748
rect 5132 28708 5174 28748
rect 5214 28708 5256 28748
rect 5296 28708 5332 28748
rect 4684 20180 4724 26776
rect 4684 20131 4724 20140
rect 4892 27236 5332 28708
rect 4892 27196 4928 27236
rect 4968 27196 5010 27236
rect 5050 27196 5092 27236
rect 5132 27196 5174 27236
rect 5214 27196 5256 27236
rect 5296 27196 5332 27236
rect 4892 25724 5332 27196
rect 4892 25684 4928 25724
rect 4968 25684 5010 25724
rect 5050 25684 5092 25724
rect 5132 25684 5174 25724
rect 5214 25684 5256 25724
rect 5296 25684 5332 25724
rect 4892 24212 5332 25684
rect 5644 44960 5684 44969
rect 4892 24172 4928 24212
rect 4968 24172 5010 24212
rect 5050 24172 5092 24212
rect 5132 24172 5174 24212
rect 5214 24172 5256 24212
rect 5296 24172 5332 24212
rect 4892 22700 5332 24172
rect 5548 25136 5588 25145
rect 4892 22660 4928 22700
rect 4968 22660 5010 22700
rect 5050 22660 5092 22700
rect 5132 22660 5174 22700
rect 5214 22660 5256 22700
rect 5296 22660 5332 22700
rect 4892 21188 5332 22660
rect 4892 21148 4928 21188
rect 4968 21148 5010 21188
rect 5050 21148 5092 21188
rect 5132 21148 5174 21188
rect 5214 21148 5256 21188
rect 5296 21148 5332 21188
rect 4300 14335 4340 14344
rect 4396 19844 4436 19853
rect 4396 17660 4436 19804
rect 4892 19676 5332 21148
rect 4892 19636 4928 19676
rect 4968 19636 5010 19676
rect 5050 19636 5092 19676
rect 5132 19636 5174 19676
rect 5214 19636 5256 19676
rect 5296 19636 5332 19676
rect 4396 14888 4436 17620
rect 4204 12536 4244 13252
rect 4204 12487 4244 12496
rect 4396 12284 4436 14848
rect 4492 19172 4532 19181
rect 4492 13208 4532 19132
rect 4892 18164 5332 19636
rect 4892 18124 4928 18164
rect 4968 18124 5010 18164
rect 5050 18124 5092 18164
rect 5132 18124 5174 18164
rect 5214 18124 5256 18164
rect 5296 18124 5332 18164
rect 4492 13159 4532 13168
rect 4588 16988 4628 16997
rect 4588 13124 4628 16948
rect 4892 16652 5332 18124
rect 4892 16612 4928 16652
rect 4968 16612 5010 16652
rect 5050 16612 5092 16652
rect 5132 16612 5174 16652
rect 5214 16612 5256 16652
rect 5296 16612 5332 16652
rect 4892 15140 5332 16612
rect 4892 15100 4928 15140
rect 4968 15100 5010 15140
rect 5050 15100 5092 15140
rect 5132 15100 5174 15140
rect 5214 15100 5256 15140
rect 5296 15100 5332 15140
rect 4588 13075 4628 13084
rect 4780 13796 4820 13805
rect 4396 12235 4436 12244
rect 3652 11320 3688 11360
rect 3728 11320 3770 11360
rect 3810 11320 3852 11360
rect 3892 11320 3934 11360
rect 3974 11320 4016 11360
rect 4056 11320 4092 11360
rect 3652 9848 4092 11320
rect 4396 11780 4436 11789
rect 4396 10772 4436 11740
rect 4396 10723 4436 10732
rect 3652 9808 3688 9848
rect 3728 9808 3770 9848
rect 3810 9808 3852 9848
rect 3892 9808 3934 9848
rect 3974 9808 4016 9848
rect 4056 9808 4092 9848
rect 3652 8336 4092 9808
rect 3652 8296 3688 8336
rect 3728 8296 3770 8336
rect 3810 8296 3852 8336
rect 3892 8296 3934 8336
rect 3974 8296 4016 8336
rect 4056 8296 4092 8336
rect 3652 6824 4092 8296
rect 4780 7244 4820 13756
rect 4780 7195 4820 7204
rect 4892 13628 5332 15100
rect 4892 13588 4928 13628
rect 4968 13588 5010 13628
rect 5050 13588 5092 13628
rect 5132 13588 5174 13628
rect 5214 13588 5256 13628
rect 5296 13588 5332 13628
rect 4892 12116 5332 13588
rect 4892 12076 4928 12116
rect 4968 12076 5010 12116
rect 5050 12076 5092 12116
rect 5132 12076 5174 12116
rect 5214 12076 5256 12116
rect 5296 12076 5332 12116
rect 4892 10604 5332 12076
rect 4892 10564 4928 10604
rect 4968 10564 5010 10604
rect 5050 10564 5092 10604
rect 5132 10564 5174 10604
rect 5214 10564 5256 10604
rect 5296 10564 5332 10604
rect 4892 9092 5332 10564
rect 4892 9052 4928 9092
rect 4968 9052 5010 9092
rect 5050 9052 5092 9092
rect 5132 9052 5174 9092
rect 5214 9052 5256 9092
rect 5296 9052 5332 9092
rect 4892 7580 5332 9052
rect 5452 23036 5492 23045
rect 5452 7748 5492 22996
rect 5548 19340 5588 25096
rect 5548 19291 5588 19300
rect 5548 13292 5588 13301
rect 5548 9512 5588 13252
rect 5548 9463 5588 9472
rect 5452 7699 5492 7708
rect 4892 7540 4928 7580
rect 4968 7540 5010 7580
rect 5050 7540 5092 7580
rect 5132 7540 5174 7580
rect 5214 7540 5256 7580
rect 5296 7540 5332 7580
rect 3652 6784 3688 6824
rect 3728 6784 3770 6824
rect 3810 6784 3852 6824
rect 3892 6784 3934 6824
rect 3974 6784 4016 6824
rect 4056 6784 4092 6824
rect 3652 5312 4092 6784
rect 3652 5272 3688 5312
rect 3728 5272 3770 5312
rect 3810 5272 3852 5312
rect 3892 5272 3934 5312
rect 3974 5272 4016 5312
rect 4056 5272 4092 5312
rect 2764 1399 2804 1408
rect 3652 3800 4092 5272
rect 3652 3760 3688 3800
rect 3728 3760 3770 3800
rect 3810 3760 3852 3800
rect 3892 3760 3934 3800
rect 3974 3760 4016 3800
rect 4056 3760 4092 3800
rect 3652 2288 4092 3760
rect 3652 2248 3688 2288
rect 3728 2248 3770 2288
rect 3810 2248 3852 2288
rect 3892 2248 3934 2288
rect 3974 2248 4016 2288
rect 4056 2248 4092 2288
rect 3652 0 4092 2248
rect 4892 6068 5332 7540
rect 4892 6028 4928 6068
rect 4968 6028 5010 6068
rect 5050 6028 5092 6068
rect 5132 6028 5174 6068
rect 5214 6028 5256 6068
rect 5296 6028 5332 6068
rect 4892 4556 5332 6028
rect 4892 4516 4928 4556
rect 4968 4516 5010 4556
rect 5050 4516 5092 4556
rect 5132 4516 5174 4556
rect 5214 4516 5256 4556
rect 5296 4516 5332 4556
rect 4892 3044 5332 4516
rect 4892 3004 4928 3044
rect 4968 3004 5010 3044
rect 5050 3004 5092 3044
rect 5132 3004 5174 3044
rect 5214 3004 5256 3044
rect 5296 3004 5332 3044
rect 4892 1532 5332 3004
rect 4892 1492 4928 1532
rect 4968 1492 5010 1532
rect 5050 1492 5092 1532
rect 5132 1492 5174 1532
rect 5214 1492 5256 1532
rect 5296 1492 5332 1532
rect 4892 0 5332 1492
rect 5644 1448 5684 44920
rect 8908 44960 8948 44969
rect 6412 44792 6452 44801
rect 6124 33368 6164 33377
rect 6124 30092 6164 33328
rect 6316 31772 6356 31781
rect 6124 30043 6164 30052
rect 6220 30260 6260 30269
rect 5740 25220 5780 25229
rect 5740 15896 5780 25180
rect 6124 17744 6164 17753
rect 5740 15847 5780 15856
rect 5836 17240 5876 17249
rect 5836 13208 5876 17200
rect 6028 16904 6068 16913
rect 5932 16736 5972 16745
rect 5932 13292 5972 16696
rect 5932 13243 5972 13252
rect 5836 9428 5876 13168
rect 6028 12956 6068 16864
rect 6028 12907 6068 12916
rect 6124 12368 6164 17704
rect 6124 12319 6164 12328
rect 5836 9379 5876 9388
rect 5644 1399 5684 1408
rect 6220 1448 6260 30220
rect 6316 14804 6356 31732
rect 6316 12368 6356 14764
rect 6316 11780 6356 12328
rect 6316 11731 6356 11740
rect 6316 10520 6356 10529
rect 6316 10016 6356 10480
rect 6316 9967 6356 9976
rect 6220 1399 6260 1408
rect 6412 188 6452 44752
rect 6604 43700 6644 43709
rect 6508 40340 6548 40349
rect 6508 7160 6548 40300
rect 6508 7111 6548 7120
rect 6604 944 6644 43660
rect 8620 43448 8660 43457
rect 6796 43364 6836 43373
rect 6796 23060 6836 43324
rect 6700 23020 6836 23060
rect 7180 37484 7220 37493
rect 6700 15980 6740 23020
rect 6700 15931 6740 15940
rect 6796 18248 6836 18257
rect 6796 10100 6836 18208
rect 6892 17912 6932 17921
rect 6892 16316 6932 17872
rect 6892 16267 6932 16276
rect 6988 17240 7028 17249
rect 6892 16064 6932 16073
rect 6892 13796 6932 16024
rect 6892 13747 6932 13756
rect 6892 12956 6932 12965
rect 6892 10688 6932 12916
rect 6892 10639 6932 10648
rect 6796 10051 6836 10060
rect 6988 8672 7028 17200
rect 6988 8623 7028 8632
rect 7180 8672 7220 37444
rect 7276 33704 7316 33713
rect 7276 18096 7316 33664
rect 8044 32864 8084 32873
rect 7564 25472 7604 25481
rect 7468 24548 7508 24557
rect 7276 18056 7412 18096
rect 7276 17996 7316 18005
rect 7276 16232 7316 17956
rect 7276 16183 7316 16192
rect 7276 13124 7316 13133
rect 7276 12872 7316 13084
rect 7276 12823 7316 12832
rect 7180 8623 7220 8632
rect 7372 8000 7412 18056
rect 7468 14720 7508 24508
rect 7468 14671 7508 14680
rect 7372 7951 7412 7960
rect 7564 6404 7604 25432
rect 8044 11948 8084 32824
rect 8524 30260 8564 30269
rect 8236 23792 8276 23801
rect 8140 16232 8180 16241
rect 8140 12956 8180 16192
rect 8140 12907 8180 12916
rect 8044 11899 8084 11908
rect 7564 6355 7604 6364
rect 8236 2876 8276 23752
rect 8428 15728 8468 15737
rect 8428 14300 8468 15688
rect 8428 14251 8468 14260
rect 8524 8168 8564 30220
rect 8524 8119 8564 8128
rect 8236 2827 8276 2836
rect 6604 895 6644 904
rect 8620 272 8660 43408
rect 8716 28832 8756 28841
rect 8716 14216 8756 28792
rect 8716 14167 8756 14176
rect 8812 13040 8852 13049
rect 8812 12788 8852 13000
rect 8812 12739 8852 12748
rect 8908 1280 8948 44920
rect 9292 44960 9332 44969
rect 8908 1231 8948 1240
rect 9100 37316 9140 37325
rect 9100 1028 9140 37276
rect 9292 7580 9332 44920
rect 10252 44876 10292 44885
rect 9484 44288 9524 44297
rect 9388 21692 9428 21701
rect 9388 11612 9428 21652
rect 9388 11563 9428 11572
rect 9484 7916 9524 44248
rect 9772 38912 9812 38921
rect 9580 37232 9620 37241
rect 9580 12704 9620 37192
rect 9580 12655 9620 12664
rect 9676 24380 9716 24389
rect 9484 7867 9524 7876
rect 9292 7531 9332 7540
rect 9100 979 9140 988
rect 9676 1028 9716 24340
rect 9772 18668 9812 38872
rect 9772 18619 9812 18628
rect 10156 30596 10196 30605
rect 9964 17240 10004 17249
rect 9964 4976 10004 17200
rect 10156 14468 10196 30556
rect 10156 14419 10196 14428
rect 9964 4927 10004 4936
rect 9676 979 9716 988
rect 10252 1028 10292 44836
rect 10636 44708 10676 44717
rect 10444 41936 10484 41945
rect 10348 34376 10388 34385
rect 10348 5648 10388 34336
rect 10348 5599 10388 5608
rect 10444 4304 10484 41896
rect 10540 33116 10580 33125
rect 10540 32528 10580 33076
rect 10540 27404 10580 32488
rect 10540 27355 10580 27364
rect 10540 27236 10580 27245
rect 10540 25976 10580 27196
rect 10540 22700 10580 25936
rect 10636 24380 10676 44668
rect 10636 24331 10676 24340
rect 10732 32696 10772 32705
rect 10540 22651 10580 22660
rect 10540 17240 10580 17249
rect 10540 14216 10580 17200
rect 10732 14552 10772 32656
rect 10732 14503 10772 14512
rect 10540 14167 10580 14176
rect 10444 4255 10484 4264
rect 10252 979 10292 988
rect 10828 1028 10868 45760
rect 11212 42776 11252 42785
rect 10924 38996 10964 39005
rect 10924 18248 10964 38956
rect 11116 38912 11156 38921
rect 10924 18199 10964 18208
rect 11020 38240 11060 38249
rect 11020 9680 11060 38200
rect 11116 17996 11156 38872
rect 11116 17947 11156 17956
rect 11020 9631 11060 9640
rect 10828 979 10868 988
rect 11212 692 11252 42736
rect 11404 41852 11444 41861
rect 11308 26732 11348 26741
rect 11308 21356 11348 26692
rect 11308 21307 11348 21316
rect 11404 1028 11444 41812
rect 11884 38912 11924 38921
rect 11596 30176 11636 30185
rect 11596 27572 11636 30136
rect 11596 27523 11636 27532
rect 11692 27404 11732 27413
rect 11692 26480 11732 27364
rect 11692 26431 11732 26440
rect 11500 18332 11540 18341
rect 11500 11948 11540 18292
rect 11596 17156 11636 17165
rect 11596 16064 11636 17116
rect 11596 16015 11636 16024
rect 11500 11899 11540 11908
rect 11884 2456 11924 38872
rect 11980 37400 12020 37409
rect 11980 17324 12020 37360
rect 12076 33704 12116 33713
rect 12076 28832 12116 33664
rect 12076 28783 12116 28792
rect 12844 29084 12884 29093
rect 12844 27908 12884 29044
rect 12844 27859 12884 27868
rect 13612 20180 13652 20189
rect 11980 17275 12020 17284
rect 13420 18416 13460 18425
rect 13420 17240 13460 18376
rect 13612 17492 13652 20140
rect 13612 17443 13652 17452
rect 13420 17191 13460 17200
rect 11884 2407 11924 2416
rect 11404 979 11444 988
rect 11212 643 11252 652
rect 8620 223 8660 232
rect 6412 139 6452 148
use sg13g2_inv_1  _049_
timestamp 1676382929
transform -1 0 5376 0 1 10584
box -48 -56 336 834
use sg13g2_inv_1  _050_
timestamp 1676382929
transform 1 0 4704 0 -1 9072
box -48 -56 336 834
use sg13g2_mux2_1  _051_
timestamp 1677247768
transform 1 0 4704 0 -1 15120
box -48 -56 1008 834
use sg13g2_or2_1  _052_
timestamp 1684236171
transform 1 0 5376 0 -1 18144
box -48 -56 528 834
use sg13g2_a21oi_1  _053_
timestamp 1683973020
transform -1 0 3936 0 -1 15120
box -48 -56 528 834
use sg13g2_a221oi_1  _054_
timestamp 1685197497
transform 1 0 5280 0 1 16632
box -48 -56 816 834
use sg13g2_nand2_1  _055_
timestamp 1676557249
transform -1 0 6048 0 -1 15120
box -48 -56 432 834
use sg13g2_nand2b_1  _056_
timestamp 1676567195
transform 1 0 6432 0 -1 18144
box -48 -56 528 834
use sg13g2_a21oi_1  _057_
timestamp 1683973020
transform -1 0 7584 0 1 16632
box -48 -56 528 834
use sg13g2_nor2b_1  _058_
timestamp 1685181386
transform 1 0 4800 0 1 16632
box -54 -56 528 834
use sg13g2_o21ai_1  _059_
timestamp 1685175443
transform -1 0 6528 0 1 16632
box -48 -56 538 834
use sg13g2_o21ai_1  _060_
timestamp 1685175443
transform 1 0 6048 0 -1 13608
box -48 -56 538 834
use sg13g2_o21ai_1  _061_
timestamp 1685175443
transform -1 0 6432 0 -1 18144
box -48 -56 538 834
use sg13g2_mux4_1  _062_
timestamp 1677257233
transform 1 0 5376 0 -1 16632
box -48 -56 2064 834
use sg13g2_mux4_1  _063_
timestamp 1677257233
transform 1 0 6240 0 1 15120
box -48 -56 2064 834
use sg13g2_mux2_1  _064_
timestamp 1677247768
transform -1 0 9024 0 -1 15120
box -48 -56 1008 834
use sg13g2_nand2b_1  _065_
timestamp 1676567195
transform 1 0 6624 0 1 16632
box -48 -56 528 834
use sg13g2_o21ai_1  _066_
timestamp 1685175443
transform 1 0 6720 0 -1 13608
box -48 -56 538 834
use sg13g2_mux2_1  _067_
timestamp 1677247768
transform -1 0 5760 0 1 13608
box -48 -56 1008 834
use sg13g2_or2_1  _068_
timestamp 1684236171
transform 1 0 2976 0 -1 15120
box -48 -56 528 834
use sg13g2_a21oi_1  _069_
timestamp 1683973020
transform 1 0 4512 0 -1 13608
box -48 -56 528 834
use sg13g2_a221oi_1  _070_
timestamp 1685197497
transform -1 0 4704 0 -1 15120
box -48 -56 816 834
use sg13g2_nand2_1  _071_
timestamp 1676557249
transform 1 0 5856 0 1 12096
box -48 -56 432 834
use sg13g2_nand2b_1  _072_
timestamp 1676567195
transform 1 0 5376 0 1 12096
box -48 -56 528 834
use sg13g2_a21oi_1  _073_
timestamp 1683973020
transform 1 0 7584 0 1 16632
box -48 -56 528 834
use sg13g2_nor2b_1  _074_
timestamp 1685181386
transform 1 0 4992 0 -1 13608
box -54 -56 528 834
use sg13g2_o21ai_1  _075_
timestamp 1685175443
transform -1 0 5952 0 -1 13608
box -48 -56 538 834
use sg13g2_o21ai_1  _076_
timestamp 1685175443
transform 1 0 6048 0 1 13608
box -48 -56 538 834
use sg13g2_o21ai_1  _077_
timestamp 1685175443
transform -1 0 5376 0 1 12096
box -48 -56 538 834
use sg13g2_mux4_1  _078_
timestamp 1677257233
transform 1 0 4224 0 1 15120
box -48 -56 2064 834
use sg13g2_mux4_1  _079_
timestamp 1677257233
transform 1 0 6048 0 -1 15120
box -48 -56 2064 834
use sg13g2_mux2_1  _080_
timestamp 1677247768
transform 1 0 6720 0 1 13608
box -48 -56 1008 834
use sg13g2_nand2b_1  _081_
timestamp 1676567195
transform 1 0 7680 0 1 13608
box -48 -56 528 834
use sg13g2_o21ai_1  _082_
timestamp 1685175443
transform 1 0 8256 0 1 15120
box -48 -56 538 834
use sg13g2_mux4_1  _083_
timestamp 1677257233
transform 1 0 10272 0 1 19656
box -48 -56 2064 834
use sg13g2_mux4_1  _084_
timestamp 1677257233
transform 1 0 9600 0 1 12096
box -48 -56 2064 834
use sg13g2_mux4_1  _085_
timestamp 1677257233
transform 1 0 6912 0 1 34776
box -48 -56 2064 834
use sg13g2_mux4_1  _086_
timestamp 1677257233
transform 1 0 9696 0 1 28728
box -48 -56 2064 834
use sg13g2_mux4_1  _087_
timestamp 1677257233
transform 1 0 10368 0 -1 18144
box -48 -56 2064 834
use sg13g2_mux4_1  _088_
timestamp 1677257233
transform -1 0 11040 0 -1 12096
box -48 -56 2064 834
use sg13g2_mux4_1  _089_
timestamp 1677257233
transform 1 0 7488 0 1 4536
box -48 -56 2064 834
use sg13g2_mux4_1  _090_
timestamp 1677257233
transform 1 0 4032 0 1 22680
box -48 -56 2064 834
use sg13g2_mux4_1  _091_
timestamp 1677257233
transform 1 0 6912 0 -1 37800
box -48 -56 2064 834
use sg13g2_mux4_1  _092_
timestamp 1677257233
transform 1 0 7680 0 -1 24192
box -48 -56 2064 834
use sg13g2_mux4_1  _093_
timestamp 1677257233
transform 1 0 7872 0 -1 6048
box -48 -56 2064 834
use sg13g2_mux4_1  _094_
timestamp 1677257233
transform 1 0 4224 0 -1 27216
box -48 -56 2064 834
use sg13g2_mux4_1  _095_
timestamp 1677257233
transform 1 0 6528 0 1 18144
box -48 -56 2064 834
use sg13g2_mux4_1  _096_
timestamp 1677257233
transform 1 0 5664 0 -1 12096
box -48 -56 2064 834
use sg13g2_mux4_1  _097_
timestamp 1677257233
transform 1 0 4224 0 1 31752
box -48 -56 2064 834
use sg13g2_mux4_1  _098_
timestamp 1677257233
transform 1 0 3936 0 -1 30240
box -48 -56 2064 834
use sg13g2_mux4_1  _099_
timestamp 1677257233
transform -1 0 11904 0 -1 36288
box -48 -56 2064 834
use sg13g2_mux4_1  _100_
timestamp 1677257233
transform 1 0 9792 0 1 25704
box -48 -56 2064 834
use sg13g2_mux4_1  _101_
timestamp 1677257233
transform 1 0 4416 0 -1 31752
box -48 -56 2064 834
use sg13g2_mux4_1  _102_
timestamp 1677257233
transform 1 0 9504 0 -1 33264
box -48 -56 2064 834
use sg13g2_mux4_1  _103_
timestamp 1677257233
transform 1 0 7392 0 -1 16632
box -48 -56 2064 834
use sg13g2_mux4_1  _104_
timestamp 1677257233
transform 1 0 6816 0 1 12096
box -48 -56 2064 834
use sg13g2_mux4_1  _105_
timestamp 1677257233
transform 1 0 5472 0 1 9072
box -48 -56 2064 834
use sg13g2_mux4_1  _106_
timestamp 1677257233
transform 1 0 4704 0 1 21168
box -48 -56 2064 834
use sg13g2_mux4_1  _107_
timestamp 1677257233
transform 1 0 4416 0 -1 33264
box -48 -56 2064 834
use sg13g2_mux4_1  _108_
timestamp 1677257233
transform 1 0 5376 0 1 30240
box -48 -56 2064 834
use sg13g2_mux4_1  _109_
timestamp 1677257233
transform 1 0 9024 0 -1 37800
box -48 -56 2064 834
use sg13g2_mux4_1  _110_
timestamp 1677257233
transform 1 0 8640 0 1 27216
box -48 -56 2064 834
use sg13g2_mux4_1  _111_
timestamp 1677257233
transform 1 0 9120 0 1 18144
box -48 -56 2064 834
use sg13g2_mux4_1  _112_
timestamp 1677257233
transform 1 0 5856 0 -1 10584
box -48 -56 2064 834
use sg13g2_mux4_1  _113_
timestamp 1677257233
transform 1 0 5472 0 1 4536
box -48 -56 2064 834
use sg13g2_mux4_1  _114_
timestamp 1677257233
transform -1 0 5760 0 -1 21168
box -48 -56 2064 834
use sg13g2_mux4_1  _115_
timestamp 1677257233
transform 1 0 7680 0 -1 34776
box -48 -56 2064 834
use sg13g2_mux4_1  _116_
timestamp 1677257233
transform 1 0 9600 0 -1 27216
box -48 -56 2064 834
use sg13g2_mux4_1  _117_
timestamp 1677257233
transform 1 0 6528 0 -1 39312
box -48 -56 2064 834
use sg13g2_mux4_1  _118_
timestamp 1677257233
transform 1 0 7488 0 1 22680
box -48 -56 2064 834
use sg13g2_mux4_1  _119_
timestamp 1677257233
transform 1 0 9792 0 1 16632
box -48 -56 2064 834
use sg13g2_mux4_1  _120_
timestamp 1677257233
transform 1 0 8064 0 1 10584
box -48 -56 2064 834
use sg13g2_mux4_1  _121_
timestamp 1677257233
transform 1 0 7104 0 -1 4536
box -48 -56 2064 834
use sg13g2_mux4_1  _122_
timestamp 1677257233
transform 1 0 4416 0 -1 22680
box -48 -56 2064 834
use sg13g2_mux4_1  _123_
timestamp 1677257233
transform 1 0 6624 0 1 33264
box -48 -56 2064 834
use sg13g2_mux4_1  _124_
timestamp 1677257233
transform 1 0 8448 0 -1 28728
box -48 -56 2064 834
use sg13g2_mux4_1  _125_
timestamp 1677257233
transform 1 0 7008 0 1 37800
box -48 -56 2064 834
use sg13g2_mux4_1  _126_
timestamp 1677257233
transform 1 0 7200 0 -1 22680
box -48 -56 2064 834
use sg13g2_mux2_1  _127_
timestamp 1677247768
transform 1 0 9120 0 -1 21168
box -48 -56 1008 834
use sg13g2_mux2_1  _128_
timestamp 1677247768
transform 1 0 8832 0 1 7560
box -48 -56 1008 834
use sg13g2_mux2_1  _129_
timestamp 1677247768
transform 1 0 3936 0 1 12096
box -48 -56 1008 834
use sg13g2_mux2_1  _130_
timestamp 1677247768
transform 1 0 6528 0 1 6048
box -48 -56 1008 834
use sg13g2_nand2b_1  _131_
timestamp 1676567195
transform -1 0 6720 0 -1 9072
box -48 -56 528 834
use sg13g2_o21ai_1  _132_
timestamp 1685175443
transform -1 0 6432 0 1 10584
box -48 -56 538 834
use sg13g2_nand3_1  _133_
timestamp 1683988354
transform 1 0 5664 0 1 7560
box -48 -56 528 834
use sg13g2_o21ai_1  _134_
timestamp 1685175443
transform 1 0 5376 0 1 10584
box -48 -56 538 834
use sg13g2_nand3b_1  _135_
timestamp 1676573470
transform 1 0 4992 0 -1 9072
box -48 -56 720 834
use sg13g2_o21ai_1  _136_
timestamp 1685175443
transform 1 0 5088 0 -1 7560
box -48 -56 538 834
use sg13g2_nand2_1  _137_
timestamp 1676557249
transform 1 0 5088 0 1 9072
box -48 -56 432 834
use sg13g2_nand4_1  _138_
timestamp 1685201930
transform 1 0 5664 0 -1 9072
box -48 -56 624 834
use sg13g2_o21ai_1  _139_
timestamp 1685175443
transform 1 0 6720 0 -1 9072
box -48 -56 538 834
use sg13g2_nand2b_1  _140_
timestamp 1676567195
transform 1 0 8448 0 1 25704
box -48 -56 528 834
use sg13g2_mux4_1  _141_
timestamp 1677257233
transform 1 0 6720 0 1 24192
box -48 -56 2064 834
use sg13g2_o21ai_1  _142_
timestamp 1685175443
transform 1 0 7200 0 -1 27216
box -48 -56 538 834
use sg13g2_o21ai_1  _143_
timestamp 1685175443
transform 1 0 8448 0 -1 25704
box -48 -56 538 834
use sg13g2_nand2b_1  _144_
timestamp 1676567195
transform -1 0 8448 0 -1 25704
box -48 -56 528 834
use sg13g2_o21ai_1  _145_
timestamp 1685175443
transform 1 0 8928 0 -1 25704
box -48 -56 538 834
use sg13g2_dlhq_1  _146_
timestamp 1678805552
transform -1 0 12384 0 -1 24192
box -50 -56 1692 834
use sg13g2_dlhq_1  _147_
timestamp 1678805552
transform -1 0 12384 0 1 21168
box -50 -56 1692 834
use sg13g2_dlhq_1  _148_
timestamp 1678805552
transform -1 0 12384 0 -1 22680
box -50 -56 1692 834
use sg13g2_dlhq_1  _149_
timestamp 1678805552
transform -1 0 12384 0 1 22680
box -50 -56 1692 834
use sg13g2_dlhq_1  _150_
timestamp 1678805552
transform -1 0 3744 0 1 24192
box -50 -56 1692 834
use sg13g2_dlhq_1  _151_
timestamp 1678805552
transform -1 0 2784 0 1 25704
box -50 -56 1692 834
use sg13g2_dlhq_1  _152_
timestamp 1678805552
transform -1 0 4320 0 -1 25704
box -50 -56 1692 834
use sg13g2_dlhq_1  _153_
timestamp 1678805552
transform -1 0 4416 0 1 25704
box -50 -56 1692 834
use sg13g2_dlhq_1  _154_
timestamp 1678805552
transform 1 0 3840 0 1 4536
box -50 -56 1692 834
use sg13g2_dlhq_1  _155_
timestamp 1678805552
transform 1 0 2400 0 1 10584
box -50 -56 1692 834
use sg13g2_dlhq_1  _156_
timestamp 1678805552
transform 1 0 6720 0 -1 7560
box -50 -56 1692 834
use sg13g2_dlhq_1  _157_
timestamp 1678805552
transform 1 0 7872 0 1 19656
box -50 -56 1692 834
use sg13g2_dlhq_1  _158_
timestamp 1678805552
transform 1 0 5664 0 -1 24192
box -50 -56 1692 834
use sg13g2_dlhq_1  _159_
timestamp 1678805552
transform 1 0 6720 0 1 21168
box -50 -56 1692 834
use sg13g2_dlhq_1  _160_
timestamp 1678805552
transform 1 0 5856 0 1 39312
box -50 -56 1692 834
use sg13g2_dlhq_1  _161_
timestamp 1678805552
transform 1 0 5376 0 1 37800
box -50 -56 1692 834
use sg13g2_dlhq_1  _162_
timestamp 1678805552
transform 1 0 6336 0 1 28728
box -50 -56 1692 834
use sg13g2_dlhq_1  _163_
timestamp 1678805552
transform 1 0 7968 0 1 28728
box -50 -56 1692 834
use sg13g2_dlhq_1  _164_
timestamp 1678805552
transform 1 0 4416 0 -1 34776
box -50 -56 1692 834
use sg13g2_dlhq_1  _165_
timestamp 1678805552
transform 1 0 6048 0 -1 34776
box -50 -56 1692 834
use sg13g2_dlhq_1  _166_
timestamp 1678805552
transform 1 0 2400 0 1 22680
box -50 -56 1692 834
use sg13g2_dlhq_1  _167_
timestamp 1678805552
transform 1 0 2784 0 -1 22680
box -50 -56 1692 834
use sg13g2_dlhq_1  _168_
timestamp 1678805552
transform 1 0 5664 0 1 3024
box -50 -56 1692 834
use sg13g2_dlhq_1  _169_
timestamp 1678805552
transform -1 0 10752 0 -1 4536
box -50 -56 1692 834
use sg13g2_dlhq_1  _170_
timestamp 1678805552
transform 1 0 7392 0 -1 9072
box -50 -56 1692 834
use sg13g2_dlhq_1  _171_
timestamp 1678805552
transform 1 0 8256 0 1 9072
box -50 -56 1692 834
use sg13g2_dlhq_1  _172_
timestamp 1678805552
transform 1 0 8160 0 1 16632
box -50 -56 1692 834
use sg13g2_dlhq_1  _173_
timestamp 1678805552
transform 1 0 10560 0 1 13608
box -50 -56 1692 834
use sg13g2_dlhq_1  _174_
timestamp 1678805552
transform -1 0 8928 0 -1 31752
box -50 -56 1692 834
use sg13g2_dlhq_1  _175_
timestamp 1678805552
transform 1 0 7872 0 1 31752
box -50 -56 1692 834
use sg13g2_dlhq_1  _176_
timestamp 1678805552
transform 1 0 3744 0 1 37800
box -50 -56 1692 834
use sg13g2_dlhq_1  _177_
timestamp 1678805552
transform 1 0 4896 0 -1 39312
box -50 -56 1692 834
use sg13g2_dlhq_1  _178_
timestamp 1678805552
transform -1 0 11328 0 -1 25704
box -50 -56 1692 834
use sg13g2_dlhq_1  _179_
timestamp 1678805552
transform 1 0 10464 0 -1 28728
box -50 -56 1692 834
use sg13g2_dlhq_1  _180_
timestamp 1678805552
transform -1 0 11328 0 -1 34776
box -50 -56 1692 834
use sg13g2_dlhq_1  _181_
timestamp 1678805552
transform -1 0 10944 0 1 34776
box -50 -56 1692 834
use sg13g2_dlhq_1  _182_
timestamp 1678805552
transform 1 0 2112 0 -1 19656
box -50 -56 1692 834
use sg13g2_dlhq_1  _183_
timestamp 1678805552
transform 1 0 2592 0 1 19656
box -50 -56 1692 834
use sg13g2_dlhq_1  _184_
timestamp 1678805552
transform 1 0 2208 0 1 4536
box -50 -56 1692 834
use sg13g2_dlhq_1  _185_
timestamp 1678805552
transform 1 0 2976 0 -1 6048
box -50 -56 1692 834
use sg13g2_dlhq_1  _186_
timestamp 1678805552
transform 1 0 3840 0 -1 4536
box -50 -56 1692 834
use sg13g2_dlhq_1  _187_
timestamp 1678805552
transform 1 0 2976 0 -1 9072
box -50 -56 1692 834
use sg13g2_dlhq_1  _188_
timestamp 1678805552
transform 1 0 7584 0 -1 18144
box -50 -56 1692 834
use sg13g2_dlhq_1  _189_
timestamp 1678805552
transform 1 0 8160 0 -1 19656
box -50 -56 1692 834
use sg13g2_dlhq_1  _190_
timestamp 1678805552
transform 1 0 6816 0 -1 28728
box -50 -56 1692 834
use sg13g2_dlhq_1  _191_
timestamp 1678805552
transform 1 0 6720 0 1 27216
box -50 -56 1692 834
use sg13g2_dlhq_1  _192_
timestamp 1678805552
transform 1 0 9024 0 1 37800
box -50 -56 1692 834
use sg13g2_dlhq_1  _193_
timestamp 1678805552
transform 1 0 7488 0 1 39312
box -50 -56 1692 834
use sg13g2_dlhq_1  _194_
timestamp 1678805552
transform 1 0 5952 0 -1 30240
box -50 -56 1692 834
use sg13g2_dlhq_1  _195_
timestamp 1678805552
transform 1 0 3744 0 1 30240
box -50 -56 1692 834
use sg13g2_dlhq_1  _196_
timestamp 1678805552
transform 1 0 4224 0 1 34776
box -50 -56 1692 834
use sg13g2_dlhq_1  _197_
timestamp 1678805552
transform 1 0 3264 0 1 33264
box -50 -56 1692 834
use sg13g2_dlhq_1  _198_
timestamp 1678805552
transform 1 0 2112 0 -1 21168
box -50 -56 1692 834
use sg13g2_dlhq_1  _199_
timestamp 1678805552
transform 1 0 5760 0 -1 21168
box -50 -56 1692 834
use sg13g2_dlhq_1  _200_
timestamp 1678805552
transform 1 0 4032 0 1 3024
box -50 -56 1692 834
use sg13g2_dlhq_1  _201_
timestamp 1678805552
transform 1 0 6240 0 -1 6048
box -50 -56 1692 834
use sg13g2_dlhq_1  _202_
timestamp 1678805552
transform -1 0 9408 0 -1 13608
box -50 -56 1692 834
use sg13g2_dlhq_1  _203_
timestamp 1678805552
transform -1 0 9600 0 -1 10584
box -50 -56 1692 834
use sg13g2_dlhq_1  _204_
timestamp 1678805552
transform -1 0 10560 0 1 15120
box -50 -56 1692 834
use sg13g2_dlhq_1  _205_
timestamp 1678805552
transform -1 0 11040 0 -1 15120
box -50 -56 1692 834
use sg13g2_dlhq_1  _206_
timestamp 1678805552
transform 1 0 9504 0 1 33264
box -50 -56 1692 834
use sg13g2_dlhq_1  _207_
timestamp 1678805552
transform 1 0 7872 0 -1 33264
box -50 -56 1692 834
use sg13g2_dlhq_1  _208_
timestamp 1678805552
transform 1 0 3648 0 -1 37800
box -50 -56 1692 834
use sg13g2_dlhq_1  _209_
timestamp 1678805552
transform 1 0 3072 0 1 36288
box -50 -56 1692 834
use sg13g2_dlhq_1  _210_
timestamp 1678805552
transform 1 0 10560 0 1 24192
box -50 -56 1692 834
use sg13g2_dlhq_1  _211_
timestamp 1678805552
transform -1 0 12288 0 1 27216
box -50 -56 1692 834
use sg13g2_dlhq_1  _212_
timestamp 1678805552
transform -1 0 12192 0 1 36288
box -50 -56 1692 834
use sg13g2_dlhq_1  _213_
timestamp 1678805552
transform 1 0 10944 0 1 34776
box -50 -56 1692 834
use sg13g2_dlhq_1  _214_
timestamp 1678805552
transform 1 0 3072 0 1 28728
box -50 -56 1692 834
use sg13g2_dlhq_1  _215_
timestamp 1678805552
transform 1 0 2496 0 -1 28728
box -50 -56 1692 834
use sg13g2_dlhq_1  _216_
timestamp 1678805552
transform 1 0 2592 0 1 31752
box -50 -56 1692 834
use sg13g2_dlhq_1  _217_
timestamp 1678805552
transform 1 0 2784 0 -1 31752
box -50 -56 1692 834
use sg13g2_dlhq_1  _218_
timestamp 1678805552
transform 1 0 4608 0 -1 6048
box -50 -56 1692 834
use sg13g2_dlhq_1  _219_
timestamp 1678805552
transform 1 0 3456 0 1 9072
box -50 -56 1692 834
use sg13g2_dlhq_1  _220_
timestamp 1678805552
transform 1 0 6528 0 -1 19656
box -50 -56 1692 834
use sg13g2_dlhq_1  _221_
timestamp 1678805552
transform 1 0 3936 0 1 18144
box -50 -56 1692 834
use sg13g2_dlhq_1  _222_
timestamp 1678805552
transform 1 0 2592 0 -1 27216
box -50 -56 1692 834
use sg13g2_dlhq_1  _223_
timestamp 1678805552
transform 1 0 4224 0 1 27216
box -50 -56 1692 834
use sg13g2_dlhq_1  _224_
timestamp 1678805552
transform 1 0 6624 0 1 7560
box -50 -56 1692 834
use sg13g2_dlhq_1  _225_
timestamp 1678805552
transform 1 0 7488 0 1 6048
box -50 -56 1692 834
use sg13g2_dlhq_1  _226_
timestamp 1678805552
transform 1 0 4608 0 -1 25704
box -50 -56 1692 834
use sg13g2_dlhq_1  _227_
timestamp 1678805552
transform 1 0 8736 0 1 24192
box -50 -56 1692 834
use sg13g2_dlhq_1  _228_
timestamp 1678805552
transform 1 0 4800 0 -1 36288
box -50 -56 1692 834
use sg13g2_dlhq_1  _229_
timestamp 1678805552
transform 1 0 5280 0 -1 37800
box -50 -56 1692 834
use sg13g2_dlhq_1  _230_
timestamp 1678805552
transform 1 0 2592 0 1 21168
box -50 -56 1692 834
use sg13g2_dlhq_1  _231_
timestamp 1678805552
transform 1 0 4032 0 -1 24192
box -50 -56 1692 834
use sg13g2_dlhq_1  _232_
timestamp 1678805552
transform 1 0 5472 0 -1 4536
box -50 -56 1692 834
use sg13g2_dlhq_1  _233_
timestamp 1678805552
transform 1 0 7584 0 1 3024
box -50 -56 1692 834
use sg13g2_dlhq_1  _234_
timestamp 1678805552
transform 1 0 10080 0 1 10584
box -50 -56 1692 834
use sg13g2_dlhq_1  _235_
timestamp 1678805552
transform -1 0 11520 0 1 9072
box -50 -56 1692 834
use sg13g2_dlhq_1  _236_
timestamp 1678805552
transform 1 0 9888 0 -1 16632
box -50 -56 1692 834
use sg13g2_dlhq_1  _237_
timestamp 1678805552
transform 1 0 10752 0 1 15120
box -50 -56 1692 834
use sg13g2_dlhq_1  _238_
timestamp 1678805552
transform 1 0 8544 0 1 30240
box -50 -56 1692 834
use sg13g2_dlhq_1  _239_
timestamp 1678805552
transform 1 0 9504 0 -1 31752
box -50 -56 1692 834
use sg13g2_dlhq_1  _240_
timestamp 1678805552
transform 1 0 4704 0 1 36288
box -50 -56 1692 834
use sg13g2_dlhq_1  _241_
timestamp 1678805552
transform 1 0 6336 0 1 36288
box -50 -56 1692 834
use sg13g2_dlhq_1  _242_
timestamp 1678805552
transform -1 0 11424 0 -1 10584
box -50 -56 1692 834
use sg13g2_dlhq_1  _243_
timestamp 1678805552
transform 1 0 10464 0 -1 13608
box -50 -56 1692 834
use sg13g2_dlhq_1  _244_
timestamp 1678805552
transform -1 0 11712 0 -1 21168
box -50 -56 1692 834
use sg13g2_dlhq_1  _245_
timestamp 1678805552
transform 1 0 10656 0 -1 19656
box -50 -56 1692 834
use sg13g2_dlhq_1  _246_
timestamp 1678805552
transform 1 0 2400 0 1 15120
box -50 -56 1692 834
use sg13g2_dlhq_1  _247_
timestamp 1678805552
transform 1 0 2400 0 -1 18144
box -50 -56 1692 834
use sg13g2_dlhq_1  _248_
timestamp 1678805552
transform 1 0 2880 0 -1 13608
box -50 -56 1692 834
use sg13g2_dlhq_1  _249_
timestamp 1678805552
transform 1 0 3072 0 1 13608
box -50 -56 1692 834
use sg13g2_dlhq_1  _250_
timestamp 1678805552
transform 1 0 3648 0 1 6048
box -50 -56 1692 834
use sg13g2_dlhq_1  _251_
timestamp 1678805552
transform 1 0 2592 0 -1 10584
box -50 -56 1692 834
use sg13g2_dlhq_1  _252_
timestamp 1678805552
transform 1 0 4032 0 1 7560
box -50 -56 1692 834
use sg13g2_dlhq_1  _253_
timestamp 1678805552
transform 1 0 1824 0 -1 16632
box -50 -56 1692 834
use sg13g2_dlhq_1  _254_
timestamp 1678805552
transform 1 0 3072 0 1 16632
box -50 -56 1692 834
use sg13g2_dlhq_1  _255_
timestamp 1678805552
transform 1 0 3456 0 -1 16632
box -50 -56 1692 834
use sg13g2_dlhq_1  _256_
timestamp 1678805552
transform 1 0 4224 0 -1 10584
box -50 -56 1692 834
use sg13g2_dlhq_1  _257_
timestamp 1678805552
transform 1 0 6240 0 -1 25704
box -50 -56 1692 834
use sg13g2_dlhq_1  _258_
timestamp 1678805552
transform 1 0 5184 0 1 25704
box -50 -56 1692 834
use sg13g2_dlhq_1  _259_
timestamp 1678805552
transform 1 0 6816 0 1 25704
box -50 -56 1692 834
use sg13g2_tiehi  _260__196
timestamp 1680000651
transform 1 0 10560 0 1 30240
box -48 -56 432 834
use sg13g2_dfrbp_1  _260_
timestamp 1678705109
transform 1 0 10080 0 -1 30240
box -60 -56 2556 834
use sg13g2_tiehi  _261__197
timestamp 1680000651
transform -1 0 11520 0 1 33264
box -48 -56 432 834
use sg13g2_dfrbp_1  _261_
timestamp 1678705109
transform 1 0 10080 0 1 31752
box -60 -56 2556 834
use sg13g2_buf_1  _264_
timestamp 1676381911
transform -1 0 12480 0 -1 28728
box -48 -56 432 834
use sg13g2_buf_1  _265_
timestamp 1676381911
transform 1 0 8640 0 1 33264
box -48 -56 432 834
use sg13g2_buf_1  _266_
timestamp 1676381911
transform 1 0 6432 0 -1 22680
box -48 -56 432 834
use sg13g2_buf_1  _267_
timestamp 1676381911
transform -1 0 9984 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  _268_
timestamp 1676381911
transform -1 0 11808 0 -1 10584
box -48 -56 432 834
use sg13g2_buf_1  _269_
timestamp 1676381911
transform -1 0 11808 0 -1 15120
box -48 -56 432 834
use sg13g2_buf_1  _270_
timestamp 1676381911
transform 1 0 10272 0 1 22680
box -48 -56 432 834
use sg13g2_buf_1  _271_
timestamp 1676381911
transform 1 0 8544 0 -1 39312
box -48 -56 432 834
use sg13g2_buf_1  _272_
timestamp 1676381911
transform -1 0 12192 0 1 25704
box -48 -56 432 834
use sg13g2_buf_1  _273_
timestamp 1676381911
transform -1 0 11712 0 -1 34776
box -48 -56 432 834
use sg13g2_buf_1  _274_
timestamp 1676381911
transform 1 0 4320 0 1 21168
box -48 -56 432 834
use sg13g2_buf_1  _275_
timestamp 1676381911
transform 1 0 7872 0 -1 3024
box -48 -56 432 834
use sg13g2_buf_1  _276_
timestamp 1676381911
transform 1 0 7776 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  _277_
timestamp 1676381911
transform -1 0 12192 0 1 16632
box -48 -56 432 834
use sg13g2_buf_1  _278_
timestamp 1676381911
transform 1 0 6240 0 -1 27216
box -48 -56 432 834
use sg13g2_buf_1  _279_
timestamp 1676381911
transform 1 0 9888 0 -1 6048
box -48 -56 432 834
use sg13g2_buf_1  _280_
timestamp 1676381911
transform 1 0 9696 0 -1 24192
box -48 -56 432 834
use sg13g2_buf_1  _281_
timestamp 1676381911
transform 1 0 8928 0 -1 39312
box -48 -56 432 834
use sg13g2_buf_1  _282_
timestamp 1676381911
transform 1 0 6048 0 1 22680
box -48 -56 432 834
use sg13g2_buf_1  _283_
timestamp 1676381911
transform -1 0 10272 0 1 4536
box -48 -56 432 834
use sg13g2_buf_1  _284_
timestamp 1676381911
transform 1 0 9216 0 1 12096
box -48 -56 432 834
use sg13g2_buf_1  _285_
timestamp 1676381911
transform 1 0 11520 0 -1 16632
box -48 -56 432 834
use sg13g2_buf_1  _286_
timestamp 1676381911
transform 1 0 11328 0 1 30240
box -48 -56 432 834
use sg13g2_buf_1  _287_
timestamp 1676381911
transform 1 0 8928 0 1 34776
box -48 -56 432 834
use sg13g2_buf_1  _288_
timestamp 1676381911
transform 1 0 11520 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  _289_
timestamp 1676381911
transform 1 0 11328 0 1 18144
box -48 -56 432 834
use sg13g2_buf_1  _290_
timestamp 1676381911
transform 1 0 11616 0 -1 27216
box -48 -56 432 834
use sg13g2_buf_1  _291_
timestamp 1676381911
transform 1 0 10944 0 1 37800
box -48 -56 432 834
use sg13g2_buf_1  _292_
timestamp 1676381911
transform 1 0 7392 0 1 30240
box -48 -56 432 834
use sg13g2_buf_1  _293_
timestamp 1676381911
transform 1 0 6816 0 -1 33264
box -48 -56 432 834
use sg13g2_buf_1  _294_
timestamp 1676381911
transform 1 0 6816 0 -1 22680
box -48 -56 432 834
use sg13g2_buf_1  _295_
timestamp 1676381911
transform 1 0 8256 0 1 7560
box -48 -56 432 834
use sg13g2_buf_1  _296_
timestamp 1676381911
transform 1 0 9408 0 -1 13608
box -48 -56 432 834
use sg13g2_buf_1  _297_
timestamp 1676381911
transform 1 0 9408 0 -1 16632
box -48 -56 432 834
use sg13g2_buf_1  _298_
timestamp 1676381911
transform 1 0 9120 0 1 33264
box -48 -56 432 834
use sg13g2_buf_1  _299_
timestamp 1676381911
transform 1 0 6240 0 1 31752
box -48 -56 432 834
use sg13g2_buf_1  _300_
timestamp 1676381911
transform -1 0 12384 0 -1 27216
box -48 -56 432 834
use sg13g2_buf_1  _301_
timestamp 1676381911
transform -1 0 11424 0 -1 37800
box -48 -56 432 834
use sg13g2_buf_1  _302_
timestamp 1676381911
transform 1 0 5280 0 1 28728
box -48 -56 432 834
use sg13g2_buf_1  _303_
timestamp 1676381911
transform 1 0 6432 0 -1 33264
box -48 -56 432 834
use sg13g2_buf_1  _304_
timestamp 1676381911
transform 1 0 7680 0 -1 12096
box -48 -56 432 834
use sg13g2_buf_1  _305_
timestamp 1676381911
transform 1 0 8544 0 1 18144
box -48 -56 432 834
use sg13g2_buf_1  _306_
timestamp 1676381911
transform 1 0 4416 0 -1 36288
box -48 -56 432 834
use sg13g2_buf_1  _307_
timestamp 1676381911
transform 1 0 3840 0 1 34776
box -48 -56 432 834
use sg13g2_buf_1  _308_
timestamp 1676381911
transform 1 0 2208 0 1 21168
box -48 -56 432 834
use sg13g2_buf_1  _309_
timestamp 1676381911
transform 1 0 4416 0 1 24192
box -48 -56 432 834
use sg13g2_buf_1  _310_
timestamp 1676381911
transform 1 0 5088 0 -1 3024
box -48 -56 432 834
use sg13g2_buf_1  _311_
timestamp 1676381911
transform 1 0 6912 0 -1 3024
box -48 -56 432 834
use sg13g2_buf_1  _312_
timestamp 1676381911
transform 1 0 7680 0 1 10584
box -48 -56 432 834
use sg13g2_buf_1  _313_
timestamp 1676381911
transform 1 0 7296 0 1 10584
box -48 -56 432 834
use sg13g2_buf_1  _314_
timestamp 1676381911
transform 1 0 9600 0 -1 18144
box -48 -56 432 834
use sg13g2_buf_1  _315_
timestamp 1676381911
transform 1 0 11040 0 -1 15120
box -48 -56 432 834
use sg13g2_buf_1  _316_
timestamp 1676381911
transform 1 0 8928 0 -1 31752
box -48 -56 432 834
use sg13g2_buf_1  _317_
timestamp 1676381911
transform 1 0 9504 0 1 31752
box -48 -56 432 834
use sg13g2_buf_1  _318_
timestamp 1676381911
transform 1 0 4128 0 -1 39312
box -48 -56 432 834
use sg13g2_buf_1  _319_
timestamp 1676381911
transform 1 0 4512 0 -1 39312
box -48 -56 432 834
use sg13g2_buf_1  _320_
timestamp 1676381911
transform 1 0 11040 0 -1 12096
box -48 -56 432 834
use sg13g2_buf_1  _321_
timestamp 1676381911
transform 1 0 10176 0 1 13608
box -48 -56 432 834
use sg13g2_buf_1  _322_
timestamp 1676381911
transform 1 0 10176 0 1 36288
box -48 -56 432 834
use sg13g2_buf_1  _323_
timestamp 1676381911
transform 1 0 9504 0 -1 36288
box -48 -56 432 834
use sg13g2_buf_1  _324_
timestamp 1676381911
transform 1 0 2304 0 1 28728
box -48 -56 432 834
use sg13g2_buf_1  _325_
timestamp 1676381911
transform 1 0 2016 0 -1 18144
box -48 -56 432 834
use sg13g2_buf_1  _326_
timestamp 1676381911
transform 1 0 2880 0 -1 12096
box -48 -56 432 834
use sg13g2_buf_1  _327_
timestamp 1676381911
transform 1 0 3072 0 -1 4536
box -48 -56 432 834
use sg13g2_buf_1  _328_
timestamp 1676381911
transform 1 0 3456 0 -1 4536
box -48 -56 432 834
use sg13g2_buf_1  _329_
timestamp 1676381911
transform 1 0 2688 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  _330_
timestamp 1676381911
transform 1 0 4608 0 -1 7560
box -48 -56 432 834
use sg13g2_buf_1  _331_
timestamp 1676381911
transform 1 0 3072 0 1 18144
box -48 -56 432 834
use sg13g2_buf_1  _332_
timestamp 1676381911
transform 1 0 4032 0 -1 18144
box -48 -56 432 834
use sg13g2_buf_1  _333_
timestamp 1676381911
transform 1 0 4416 0 1 25704
box -48 -56 432 834
use sg13g2_buf_1  _334_
timestamp 1676381911
transform 1 0 6432 0 -1 36288
box -48 -56 432 834
use sg13g2_buf_1  _335_
timestamp 1676381911
transform 1 0 7584 0 -1 30240
box -48 -56 432 834
use sg13g2_buf_1  _336_
timestamp 1676381911
transform 1 0 5664 0 1 28728
box -48 -56 432 834
use sg13g2_buf_1  _337_
timestamp 1676381911
transform 1 0 7968 0 -1 30240
box -48 -56 432 834
use sg13g2_buf_1  _338_
timestamp 1676381911
transform -1 0 9792 0 1 13608
box -48 -56 432 834
use sg13g2_buf_1  _339_
timestamp 1676381911
transform -1 0 4416 0 -1 36288
box -48 -56 432 834
use sg13g2_buf_1  _340_
timestamp 1676381911
transform -1 0 7200 0 -1 31752
box -48 -56 432 834
use sg13g2_buf_1  _341_
timestamp 1676381911
transform -1 0 4224 0 -1 12096
box -48 -56 432 834
use sg13g2_buf_1  _342_
timestamp 1676381911
transform -1 0 12000 0 1 43848
box -48 -56 432 834
use sg13g2_buf_1  _343_
timestamp 1676381911
transform -1 0 11616 0 1 43848
box -48 -56 432 834
use sg13g2_buf_1  _344_
timestamp 1676381911
transform -1 0 11040 0 -1 45360
box -48 -56 432 834
use sg13g2_buf_1  _345_
timestamp 1676381911
transform 1 0 5376 0 -1 45360
box -48 -56 432 834
use sg13g2_buf_1  _346_
timestamp 1676381911
transform 1 0 4320 0 -1 45360
box -48 -56 432 834
use sg13g2_buf_1  _347_
timestamp 1676381911
transform -1 0 9024 0 -1 45360
box -48 -56 432 834
use sg13g2_buf_1  _348_
timestamp 1676381911
transform -1 0 8736 0 -1 43848
box -48 -56 432 834
use sg13g2_buf_1  _349_
timestamp 1676381911
transform -1 0 11232 0 1 43848
box -48 -56 432 834
use sg13g2_buf_1  _350_
timestamp 1676381911
transform -1 0 11616 0 -1 45360
box -48 -56 432 834
use sg13g2_buf_1  _351_
timestamp 1676381911
transform -1 0 10848 0 1 43848
box -48 -56 432 834
use sg13g2_buf_1  _352_
timestamp 1676381911
transform -1 0 12000 0 -1 45360
box -48 -56 432 834
use sg13g2_buf_1  _353_
timestamp 1676381911
transform -1 0 12384 0 -1 45360
box -48 -56 432 834
use sg13g2_buf_1  _354_
timestamp 1676381911
transform -1 0 11616 0 1 45360
box -48 -56 432 834
use sg13g2_buf_1  _355_
timestamp 1676381911
transform 1 0 10944 0 1 42336
box -48 -56 432 834
use sg13g2_buf_1  _356_
timestamp 1676381911
transform -1 0 11712 0 1 42336
box -48 -56 432 834
use sg13g2_buf_1  _357_
timestamp 1676381911
transform -1 0 12096 0 1 42336
box -48 -56 432 834
use sg13g2_buf_1  _358_
timestamp 1676381911
transform -1 0 10560 0 1 30240
box -48 -56 432 834
use sg13g2_buf_1  _359_
timestamp 1676381911
transform 1 0 9504 0 1 4536
box -48 -56 432 834
use sg13g2_buf_1  _360_
timestamp 1676381911
transform 1 0 4608 0 -1 12096
box -48 -56 432 834
use sg13g2_buf_1  _361_
timestamp 1676381911
transform 1 0 9792 0 1 7560
box -48 -56 432 834
use sg13g2_buf_1  _362_
timestamp 1676381911
transform -1 0 10272 0 1 19656
box -48 -56 432 834
use sg13g2_buf_1  _363_
timestamp 1676381911
transform 1 0 9888 0 1 22680
box -48 -56 432 834
use sg13g2_buf_1  _364_
timestamp 1676381911
transform 1 0 9312 0 -1 39312
box -48 -56 432 834
use sg13g2_buf_1  fanout66
timestamp 1676381911
transform 1 0 4704 0 -1 18144
box -48 -56 432 834
use sg13g2_buf_1  fanout67
timestamp 1676381911
transform 1 0 2016 0 1 15120
box -48 -56 432 834
use sg13g2_buf_1  fanout68
timestamp 1676381911
transform 1 0 9504 0 1 22680
box -48 -56 432 834
use sg13g2_buf_1  fanout69
timestamp 1676381911
transform -1 0 8064 0 -1 21168
box -48 -56 432 834
use sg13g2_buf_1  fanout70
timestamp 1676381911
transform -1 0 8736 0 -1 21168
box -48 -56 432 834
use sg13g2_buf_1  fanout71
timestamp 1676381911
transform 1 0 4224 0 -1 12096
box -48 -56 432 834
use sg13g2_buf_1  fanout72
timestamp 1676381911
transform -1 0 5664 0 1 19656
box -48 -56 432 834
use sg13g2_buf_1  fanout73
timestamp 1676381911
transform 1 0 6912 0 1 19656
box -48 -56 432 834
use sg13g2_buf_1  fanout74
timestamp 1676381911
transform 1 0 6240 0 1 33264
box -48 -56 432 834
use sg13g2_buf_1  fanout75
timestamp 1676381911
transform -1 0 6816 0 -1 31752
box -48 -56 432 834
use sg13g2_buf_1  fanout76
timestamp 1676381911
transform 1 0 7776 0 1 30240
box -48 -56 432 834
use sg13g2_buf_1  fanout77
timestamp 1676381911
transform -1 0 8544 0 1 30240
box -48 -56 432 834
use sg13g2_buf_1  fanout78
timestamp 1676381911
transform 1 0 9024 0 -1 9072
box -48 -56 432 834
use sg13g2_buf_1  fanout79
timestamp 1676381911
transform 1 0 4512 0 1 19656
box -48 -56 432 834
use sg13g2_buf_1  fanout80
timestamp 1676381911
transform 1 0 3360 0 1 30240
box -48 -56 432 834
use sg13g2_buf_1  fanout81
timestamp 1676381911
transform 1 0 4032 0 -1 33264
box -48 -56 432 834
use sg13g2_buf_1  fanout82
timestamp 1676381911
transform 1 0 3648 0 -1 33264
box -48 -56 432 834
use sg13g2_buf_1  fanout83
timestamp 1676381911
transform -1 0 3936 0 1 12096
box -48 -56 432 834
use sg13g2_buf_1  fanout84
timestamp 1676381911
transform -1 0 8448 0 -1 12096
box -48 -56 432 834
use sg13g2_buf_1  fanout85
timestamp 1676381911
transform -1 0 10368 0 1 21168
box -48 -56 432 834
use sg13g2_buf_1  fanout86
timestamp 1676381911
transform 1 0 9984 0 -1 18144
box -48 -56 432 834
use sg13g2_buf_1  fanout87
timestamp 1676381911
transform 1 0 8640 0 -1 12096
box -48 -56 432 834
use sg13g2_buf_1  fanout88
timestamp 1676381911
transform -1 0 9600 0 1 3024
box -48 -56 432 834
use sg13g2_decap_8  FILLER_0_4
timestamp 1679581782
transform 1 0 1536 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_11
timestamp 1679581782
transform 1 0 2208 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_18
timestamp 1679581782
transform 1 0 2880 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_25
timestamp 1679581782
transform 1 0 3552 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_32
timestamp 1679581782
transform 1 0 4224 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_39
timestamp 1679581782
transform 1 0 4896 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_46
timestamp 1679581782
transform 1 0 5568 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_53
timestamp 1679581782
transform 1 0 6240 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_60
timestamp 1679581782
transform 1 0 6912 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_67
timestamp 1679581782
transform 1 0 7584 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_74
timestamp 1679581782
transform 1 0 8256 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_81
timestamp 1679581782
transform 1 0 8928 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_88
timestamp 1679581782
transform 1 0 9600 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_95
timestamp 1679581782
transform 1 0 10272 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_102
timestamp 1679581782
transform 1 0 10944 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_109
timestamp 1679581782
transform 1 0 11616 0 1 1512
box -48 -56 720 834
use sg13g2_fill_2  FILLER_0_116
timestamp 1677580104
transform 1 0 12288 0 1 1512
box -48 -56 240 834
use sg13g2_fill_1  FILLER_0_118
timestamp 1677579658
transform 1 0 12480 0 1 1512
box -48 -56 144 834
use sg13g2_decap_8  FILLER_1_4
timestamp 1679581782
transform 1 0 1536 0 -1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_11
timestamp 1679581782
transform 1 0 2208 0 -1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_18
timestamp 1679581782
transform 1 0 2880 0 -1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_25
timestamp 1679581782
transform 1 0 3552 0 -1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_32
timestamp 1679581782
transform 1 0 4224 0 -1 3024
box -48 -56 720 834
use sg13g2_fill_2  FILLER_1_39
timestamp 1677580104
transform 1 0 4896 0 -1 3024
box -48 -56 240 834
use sg13g2_decap_8  FILLER_1_45
timestamp 1679581782
transform 1 0 5472 0 -1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_52
timestamp 1679581782
transform 1 0 6144 0 -1 3024
box -48 -56 720 834
use sg13g2_fill_1  FILLER_1_59
timestamp 1677579658
transform 1 0 6816 0 -1 3024
box -48 -56 144 834
use sg13g2_decap_4  FILLER_1_64
timestamp 1679577901
transform 1 0 7296 0 -1 3024
box -48 -56 432 834
use sg13g2_fill_2  FILLER_1_68
timestamp 1677580104
transform 1 0 7680 0 -1 3024
box -48 -56 240 834
use sg13g2_decap_8  FILLER_1_74
timestamp 1679581782
transform 1 0 8256 0 -1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_81
timestamp 1679581782
transform 1 0 8928 0 -1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_88
timestamp 1679581782
transform 1 0 9600 0 -1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_95
timestamp 1679581782
transform 1 0 10272 0 -1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_102
timestamp 1679581782
transform 1 0 10944 0 -1 3024
box -48 -56 720 834
use sg13g2_decap_4  FILLER_1_109
timestamp 1679577901
transform 1 0 11616 0 -1 3024
box -48 -56 432 834
use sg13g2_fill_2  FILLER_1_113
timestamp 1677580104
transform 1 0 12000 0 -1 3024
box -48 -56 240 834
use sg13g2_decap_8  FILLER_2_0
timestamp 1679581782
transform 1 0 1152 0 1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_7
timestamp 1679581782
transform 1 0 1824 0 1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_14
timestamp 1679581782
transform 1 0 2496 0 1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_21
timestamp 1679581782
transform 1 0 3168 0 1 3024
box -48 -56 720 834
use sg13g2_fill_2  FILLER_2_28
timestamp 1677580104
transform 1 0 3840 0 1 3024
box -48 -56 240 834
use sg13g2_fill_2  FILLER_2_64
timestamp 1677580104
transform 1 0 7296 0 1 3024
box -48 -56 240 834
use sg13g2_fill_1  FILLER_2_66
timestamp 1677579658
transform 1 0 7488 0 1 3024
box -48 -56 144 834
use sg13g2_decap_8  FILLER_2_92
timestamp 1679581782
transform 1 0 9984 0 1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_99
timestamp 1679581782
transform 1 0 10656 0 1 3024
box -48 -56 720 834
use sg13g2_decap_4  FILLER_2_106
timestamp 1679577901
transform 1 0 11328 0 1 3024
box -48 -56 432 834
use sg13g2_fill_1  FILLER_2_110
timestamp 1677579658
transform 1 0 11712 0 1 3024
box -48 -56 144 834
use sg13g2_decap_8  FILLER_3_4
timestamp 1679581782
transform 1 0 1536 0 -1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_11
timestamp 1679581782
transform 1 0 2208 0 -1 4536
box -48 -56 720 834
use sg13g2_fill_2  FILLER_3_18
timestamp 1677580104
transform 1 0 2880 0 -1 4536
box -48 -56 240 834
use sg13g2_decap_8  FILLER_3_100
timestamp 1679581782
transform 1 0 10752 0 -1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_4
timestamp 1679581782
transform 1 0 1536 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_95
timestamp 1679581782
transform 1 0 10272 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_102
timestamp 1679581782
transform 1 0 10944 0 1 4536
box -48 -56 720 834
use sg13g2_fill_2  FILLER_4_109
timestamp 1677580104
transform 1 0 11616 0 1 4536
box -48 -56 240 834
use sg13g2_decap_8  FILLER_5_4
timestamp 1679581782
transform 1 0 1536 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_11
timestamp 1679581782
transform 1 0 2208 0 -1 6048
box -48 -56 720 834
use sg13g2_fill_1  FILLER_5_18
timestamp 1677579658
transform 1 0 2880 0 -1 6048
box -48 -56 144 834
use sg13g2_decap_8  FILLER_5_95
timestamp 1679581782
transform 1 0 10272 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_102
timestamp 1679581782
transform 1 0 10944 0 -1 6048
box -48 -56 720 834
use sg13g2_fill_2  FILLER_5_109
timestamp 1677580104
transform 1 0 11616 0 -1 6048
box -48 -56 240 834
use sg13g2_decap_8  FILLER_6_0
timestamp 1679581782
transform 1 0 1152 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_7
timestamp 1679581782
transform 1 0 1824 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_14
timestamp 1679581782
transform 1 0 2496 0 1 6048
box -48 -56 720 834
use sg13g2_decap_4  FILLER_6_21
timestamp 1679577901
transform 1 0 3168 0 1 6048
box -48 -56 432 834
use sg13g2_fill_1  FILLER_6_25
timestamp 1677579658
transform 1 0 3552 0 1 6048
box -48 -56 144 834
use sg13g2_decap_8  FILLER_6_43
timestamp 1679581782
transform 1 0 5280 0 1 6048
box -48 -56 720 834
use sg13g2_decap_4  FILLER_6_50
timestamp 1679577901
transform 1 0 5952 0 1 6048
box -48 -56 432 834
use sg13g2_fill_2  FILLER_6_54
timestamp 1677580104
transform 1 0 6336 0 1 6048
box -48 -56 240 834
use sg13g2_decap_8  FILLER_6_83
timestamp 1679581782
transform 1 0 9120 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_90
timestamp 1679581782
transform 1 0 9792 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_97
timestamp 1679581782
transform 1 0 10464 0 1 6048
box -48 -56 720 834
use sg13g2_fill_2  FILLER_6_104
timestamp 1677580104
transform 1 0 11136 0 1 6048
box -48 -56 240 834
use sg13g2_fill_1  FILLER_6_106
timestamp 1677579658
transform 1 0 11328 0 1 6048
box -48 -56 144 834
use sg13g2_decap_8  FILLER_7_4
timestamp 1679581782
transform 1 0 1536 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_11
timestamp 1679581782
transform 1 0 2208 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_18
timestamp 1679581782
transform 1 0 2880 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_25
timestamp 1679581782
transform 1 0 3552 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_4  FILLER_7_32
timestamp 1679577901
transform 1 0 4224 0 -1 7560
box -48 -56 432 834
use sg13g2_fill_1  FILLER_7_40
timestamp 1677579658
transform 1 0 4992 0 -1 7560
box -48 -56 144 834
use sg13g2_decap_8  FILLER_7_46
timestamp 1679581782
transform 1 0 5568 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_4  FILLER_7_53
timestamp 1679577901
transform 1 0 6240 0 -1 7560
box -48 -56 432 834
use sg13g2_fill_1  FILLER_7_57
timestamp 1677579658
transform 1 0 6624 0 -1 7560
box -48 -56 144 834
use sg13g2_decap_8  FILLER_7_75
timestamp 1679581782
transform 1 0 8352 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_82
timestamp 1679581782
transform 1 0 9024 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_89
timestamp 1679581782
transform 1 0 9696 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_96
timestamp 1679581782
transform 1 0 10368 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_4
timestamp 1679581782
transform 1 0 1536 0 1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_11
timestamp 1679581782
transform 1 0 2208 0 1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_18
timestamp 1679581782
transform 1 0 2880 0 1 7560
box -48 -56 720 834
use sg13g2_decap_4  FILLER_8_25
timestamp 1679577901
transform 1 0 3552 0 1 7560
box -48 -56 432 834
use sg13g2_fill_1  FILLER_8_29
timestamp 1677579658
transform 1 0 3936 0 1 7560
box -48 -56 144 834
use sg13g2_decap_4  FILLER_8_52
timestamp 1679577901
transform 1 0 6144 0 1 7560
box -48 -56 432 834
use sg13g2_fill_1  FILLER_8_56
timestamp 1677579658
transform 1 0 6528 0 1 7560
box -48 -56 144 834
use sg13g2_fill_2  FILLER_8_78
timestamp 1677580104
transform 1 0 8640 0 1 7560
box -48 -56 240 834
use sg13g2_decap_8  FILLER_8_94
timestamp 1679581782
transform 1 0 10176 0 1 7560
box -48 -56 720 834
use sg13g2_fill_2  FILLER_8_101
timestamp 1677580104
transform 1 0 10848 0 1 7560
box -48 -56 240 834
use sg13g2_decap_8  FILLER_9_4
timestamp 1679581782
transform 1 0 1536 0 -1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_11
timestamp 1679581782
transform 1 0 2208 0 -1 9072
box -48 -56 720 834
use sg13g2_fill_1  FILLER_9_18
timestamp 1677579658
transform 1 0 2880 0 -1 9072
box -48 -56 144 834
use sg13g2_fill_1  FILLER_9_36
timestamp 1677579658
transform 1 0 4608 0 -1 9072
box -48 -56 144 834
use sg13g2_fill_2  FILLER_9_63
timestamp 1677580104
transform 1 0 7200 0 -1 9072
box -48 -56 240 834
use sg13g2_decap_8  FILLER_9_86
timestamp 1679581782
transform 1 0 9408 0 -1 9072
box -48 -56 720 834
use sg13g2_fill_2  FILLER_9_93
timestamp 1677580104
transform 1 0 10080 0 -1 9072
box -48 -56 240 834
use sg13g2_decap_8  FILLER_10_0
timestamp 1679581782
transform 1 0 1152 0 1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_7
timestamp 1679581782
transform 1 0 1824 0 1 9072
box -48 -56 720 834
use sg13g2_fill_2  FILLER_10_14
timestamp 1677580104
transform 1 0 2496 0 1 9072
box -48 -56 240 834
use sg13g2_decap_4  FILLER_10_20
timestamp 1679577901
transform 1 0 3072 0 1 9072
box -48 -56 432 834
use sg13g2_fill_2  FILLER_10_66
timestamp 1677580104
transform 1 0 7488 0 1 9072
box -48 -56 240 834
use sg13g2_fill_1  FILLER_10_68
timestamp 1677579658
transform 1 0 7680 0 1 9072
box -48 -56 144 834
use sg13g2_fill_1  FILLER_10_73
timestamp 1677579658
transform 1 0 8160 0 1 9072
box -48 -56 144 834
use sg13g2_fill_2  FILLER_10_112
timestamp 1677580104
transform 1 0 11904 0 1 9072
box -48 -56 240 834
use sg13g2_fill_1  FILLER_10_114
timestamp 1677579658
transform 1 0 12096 0 1 9072
box -48 -56 144 834
use sg13g2_decap_8  FILLER_11_4
timestamp 1679581782
transform 1 0 1536 0 -1 10584
box -48 -56 720 834
use sg13g2_decap_4  FILLER_11_11
timestamp 1679577901
transform 1 0 2208 0 -1 10584
box -48 -56 432 834
use sg13g2_fill_1  FILLER_11_70
timestamp 1677579658
transform 1 0 7872 0 -1 10584
box -48 -56 144 834
use sg13g2_fill_2  FILLER_11_88
timestamp 1677580104
transform 1 0 9600 0 -1 10584
box -48 -56 240 834
use sg13g2_decap_8  FILLER_12_4
timestamp 1679581782
transform 1 0 1536 0 1 10584
box -48 -56 720 834
use sg13g2_fill_2  FILLER_12_11
timestamp 1677580104
transform 1 0 2208 0 1 10584
box -48 -56 240 834
use sg13g2_decap_8  FILLER_12_30
timestamp 1679581782
transform 1 0 4032 0 1 10584
box -48 -56 720 834
use sg13g2_decap_4  FILLER_12_37
timestamp 1679577901
transform 1 0 4704 0 1 10584
box -48 -56 432 834
use sg13g2_fill_1  FILLER_12_49
timestamp 1677579658
transform 1 0 5856 0 1 10584
box -48 -56 144 834
use sg13g2_decap_8  FILLER_12_55
timestamp 1679581782
transform 1 0 6432 0 1 10584
box -48 -56 720 834
use sg13g2_fill_2  FILLER_12_62
timestamp 1677580104
transform 1 0 7104 0 1 10584
box -48 -56 240 834
use sg13g2_fill_1  FILLER_12_110
timestamp 1677579658
transform 1 0 11712 0 1 10584
box -48 -56 144 834
use sg13g2_decap_8  FILLER_13_4
timestamp 1679581782
transform 1 0 1536 0 -1 12096
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_11
timestamp 1679581782
transform 1 0 2208 0 -1 12096
box -48 -56 720 834
use sg13g2_decap_4  FILLER_13_22
timestamp 1679577901
transform 1 0 3264 0 -1 12096
box -48 -56 432 834
use sg13g2_fill_2  FILLER_13_26
timestamp 1677580104
transform 1 0 3648 0 -1 12096
box -48 -56 240 834
use sg13g2_decap_8  FILLER_13_40
timestamp 1679581782
transform 1 0 4992 0 -1 12096
box -48 -56 720 834
use sg13g2_fill_2  FILLER_13_76
timestamp 1677580104
transform 1 0 8448 0 -1 12096
box -48 -56 240 834
use sg13g2_decap_8  FILLER_14_0
timestamp 1679581782
transform 1 0 1152 0 1 12096
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_7
timestamp 1679581782
transform 1 0 1824 0 1 12096
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_14
timestamp 1679581782
transform 1 0 2496 0 1 12096
box -48 -56 720 834
use sg13g2_decap_4  FILLER_14_21
timestamp 1679577901
transform 1 0 3168 0 1 12096
box -48 -56 432 834
use sg13g2_decap_4  FILLER_14_53
timestamp 1679577901
transform 1 0 6240 0 1 12096
box -48 -56 432 834
use sg13g2_fill_2  FILLER_14_57
timestamp 1677580104
transform 1 0 6624 0 1 12096
box -48 -56 240 834
use sg13g2_fill_2  FILLER_14_109
timestamp 1677580104
transform 1 0 11616 0 1 12096
box -48 -56 240 834
use sg13g2_decap_8  FILLER_15_4
timestamp 1679581782
transform 1 0 1536 0 -1 13608
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_11
timestamp 1679581782
transform 1 0 2208 0 -1 13608
box -48 -56 720 834
use sg13g2_fill_1  FILLER_15_50
timestamp 1677579658
transform 1 0 5952 0 -1 13608
box -48 -56 144 834
use sg13g2_fill_2  FILLER_15_56
timestamp 1677580104
transform 1 0 6528 0 -1 13608
box -48 -56 240 834
use sg13g2_decap_4  FILLER_15_63
timestamp 1679577901
transform 1 0 7200 0 -1 13608
box -48 -56 432 834
use sg13g2_fill_2  FILLER_15_67
timestamp 1677580104
transform 1 0 7584 0 -1 13608
box -48 -56 240 834
use sg13g2_fill_2  FILLER_15_90
timestamp 1677580104
transform 1 0 9792 0 -1 13608
box -48 -56 240 834
use sg13g2_fill_1  FILLER_15_92
timestamp 1677579658
transform 1 0 9984 0 -1 13608
box -48 -56 144 834
use sg13g2_fill_1  FILLER_15_114
timestamp 1677579658
transform 1 0 12096 0 -1 13608
box -48 -56 144 834
use sg13g2_decap_8  FILLER_16_4
timestamp 1679581782
transform 1 0 1536 0 1 13608
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_11
timestamp 1679581782
transform 1 0 2208 0 1 13608
box -48 -56 720 834
use sg13g2_fill_2  FILLER_16_18
timestamp 1677580104
transform 1 0 2880 0 1 13608
box -48 -56 240 834
use sg13g2_fill_1  FILLER_16_37
timestamp 1677579658
transform 1 0 4704 0 1 13608
box -48 -56 144 834
use sg13g2_fill_2  FILLER_16_48
timestamp 1677580104
transform 1 0 5760 0 1 13608
box -48 -56 240 834
use sg13g2_fill_1  FILLER_16_50
timestamp 1677579658
transform 1 0 5952 0 1 13608
box -48 -56 144 834
use sg13g2_fill_2  FILLER_16_56
timestamp 1677580104
transform 1 0 6528 0 1 13608
box -48 -56 240 834
use sg13g2_decap_4  FILLER_16_73
timestamp 1679577901
transform 1 0 8160 0 1 13608
box -48 -56 432 834
use sg13g2_fill_1  FILLER_16_77
timestamp 1677579658
transform 1 0 8544 0 1 13608
box -48 -56 144 834
use sg13g2_decap_8  FILLER_17_4
timestamp 1679581782
transform 1 0 1536 0 -1 15120
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_11
timestamp 1679581782
transform 1 0 2208 0 -1 15120
box -48 -56 720 834
use sg13g2_fill_1  FILLER_17_18
timestamp 1677579658
transform 1 0 2880 0 -1 15120
box -48 -56 144 834
use sg13g2_decap_8  FILLER_18_0
timestamp 1679581782
transform 1 0 1152 0 1 15120
box -48 -56 720 834
use sg13g2_fill_2  FILLER_18_7
timestamp 1677580104
transform 1 0 1824 0 1 15120
box -48 -56 240 834
use sg13g2_fill_2  FILLER_18_30
timestamp 1677580104
transform 1 0 4032 0 1 15120
box -48 -56 240 834
use sg13g2_fill_2  FILLER_18_79
timestamp 1677580104
transform 1 0 8736 0 1 15120
box -48 -56 240 834
use sg13g2_fill_2  FILLER_18_98
timestamp 1677580104
transform 1 0 10560 0 1 15120
box -48 -56 240 834
use sg13g2_fill_2  FILLER_18_117
timestamp 1677580104
transform 1 0 12384 0 1 15120
box -48 -56 240 834
use sg13g2_fill_2  FILLER_19_4
timestamp 1677580104
transform 1 0 1536 0 -1 16632
box -48 -56 240 834
use sg13g2_fill_1  FILLER_19_6
timestamp 1677579658
transform 1 0 1728 0 -1 16632
box -48 -56 144 834
use sg13g2_fill_2  FILLER_19_41
timestamp 1677580104
transform 1 0 5088 0 -1 16632
box -48 -56 240 834
use sg13g2_fill_1  FILLER_19_43
timestamp 1677579658
transform 1 0 5280 0 -1 16632
box -48 -56 144 834
use sg13g2_fill_1  FILLER_19_90
timestamp 1677579658
transform 1 0 9792 0 -1 16632
box -48 -56 144 834
use sg13g2_fill_2  FILLER_19_112
timestamp 1677580104
transform 1 0 11904 0 -1 16632
box -48 -56 240 834
use sg13g2_fill_1  FILLER_19_114
timestamp 1677579658
transform 1 0 12096 0 -1 16632
box -48 -56 144 834
use sg13g2_decap_8  FILLER_20_4
timestamp 1679581782
transform 1 0 1536 0 1 16632
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_11
timestamp 1679581782
transform 1 0 2208 0 1 16632
box -48 -56 720 834
use sg13g2_fill_2  FILLER_20_18
timestamp 1677580104
transform 1 0 2880 0 1 16632
box -48 -56 240 834
use sg13g2_fill_1  FILLER_20_37
timestamp 1677579658
transform 1 0 4704 0 1 16632
box -48 -56 144 834
use sg13g2_fill_1  FILLER_20_56
timestamp 1677579658
transform 1 0 6528 0 1 16632
box -48 -56 144 834
use sg13g2_fill_1  FILLER_20_72
timestamp 1677579658
transform 1 0 8064 0 1 16632
box -48 -56 144 834
use sg13g2_decap_4  FILLER_21_4
timestamp 1679577901
transform 1 0 1536 0 -1 18144
box -48 -56 432 834
use sg13g2_fill_1  FILLER_21_8
timestamp 1677579658
transform 1 0 1920 0 -1 18144
box -48 -56 144 834
use sg13g2_fill_2  FILLER_21_34
timestamp 1677580104
transform 1 0 4416 0 -1 18144
box -48 -56 240 834
use sg13g2_fill_1  FILLER_21_36
timestamp 1677579658
transform 1 0 4608 0 -1 18144
box -48 -56 144 834
use sg13g2_fill_2  FILLER_21_41
timestamp 1677580104
transform 1 0 5088 0 -1 18144
box -48 -56 240 834
use sg13g2_fill_1  FILLER_21_43
timestamp 1677579658
transform 1 0 5280 0 -1 18144
box -48 -56 144 834
use sg13g2_fill_1  FILLER_21_49
timestamp 1677579658
transform 1 0 5856 0 -1 18144
box -48 -56 144 834
use sg13g2_decap_8  FILLER_21_60
timestamp 1679581782
transform 1 0 6912 0 -1 18144
box -48 -56 720 834
use sg13g2_fill_2  FILLER_21_117
timestamp 1677580104
transform 1 0 12384 0 -1 18144
box -48 -56 240 834
use sg13g2_decap_8  FILLER_22_0
timestamp 1679581782
transform 1 0 1152 0 1 18144
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_7
timestamp 1679581782
transform 1 0 1824 0 1 18144
box -48 -56 720 834
use sg13g2_decap_4  FILLER_22_14
timestamp 1679577901
transform 1 0 2496 0 1 18144
box -48 -56 432 834
use sg13g2_fill_2  FILLER_22_18
timestamp 1677580104
transform 1 0 2880 0 1 18144
box -48 -56 240 834
use sg13g2_decap_4  FILLER_22_24
timestamp 1679577901
transform 1 0 3456 0 1 18144
box -48 -56 432 834
use sg13g2_fill_1  FILLER_22_28
timestamp 1677579658
transform 1 0 3840 0 1 18144
box -48 -56 144 834
use sg13g2_decap_8  FILLER_22_46
timestamp 1679581782
transform 1 0 5568 0 1 18144
box -48 -56 720 834
use sg13g2_fill_2  FILLER_22_53
timestamp 1677580104
transform 1 0 6240 0 1 18144
box -48 -56 240 834
use sg13g2_fill_1  FILLER_22_55
timestamp 1677579658
transform 1 0 6432 0 1 18144
box -48 -56 144 834
use sg13g2_fill_2  FILLER_22_81
timestamp 1677580104
transform 1 0 8928 0 1 18144
box -48 -56 240 834
use sg13g2_fill_2  FILLER_22_104
timestamp 1677580104
transform 1 0 11136 0 1 18144
box -48 -56 240 834
use sg13g2_fill_1  FILLER_22_110
timestamp 1677579658
transform 1 0 11712 0 1 18144
box -48 -56 144 834
use sg13g2_decap_4  FILLER_23_4
timestamp 1679577901
transform 1 0 1536 0 -1 19656
box -48 -56 432 834
use sg13g2_fill_2  FILLER_23_8
timestamp 1677580104
transform 1 0 1920 0 -1 19656
box -48 -56 240 834
use sg13g2_decap_8  FILLER_23_27
timestamp 1679581782
transform 1 0 3744 0 -1 19656
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_34
timestamp 1679581782
transform 1 0 4416 0 -1 19656
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_41
timestamp 1679581782
transform 1 0 5088 0 -1 19656
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_48
timestamp 1679581782
transform 1 0 5760 0 -1 19656
box -48 -56 720 834
use sg13g2_fill_1  FILLER_23_55
timestamp 1677579658
transform 1 0 6432 0 -1 19656
box -48 -56 144 834
use sg13g2_fill_1  FILLER_23_90
timestamp 1677579658
transform 1 0 9792 0 -1 19656
box -48 -56 144 834
use sg13g2_fill_2  FILLER_23_116
timestamp 1677580104
transform 1 0 12288 0 -1 19656
box -48 -56 240 834
use sg13g2_fill_1  FILLER_23_118
timestamp 1677579658
transform 1 0 12480 0 -1 19656
box -48 -56 144 834
use sg13g2_decap_8  FILLER_24_4
timestamp 1679581782
transform 1 0 1536 0 1 19656
box -48 -56 720 834
use sg13g2_decap_4  FILLER_24_11
timestamp 1679577901
transform 1 0 2208 0 1 19656
box -48 -56 432 834
use sg13g2_fill_2  FILLER_24_32
timestamp 1677580104
transform 1 0 4224 0 1 19656
box -48 -56 240 834
use sg13g2_fill_1  FILLER_24_34
timestamp 1677579658
transform 1 0 4416 0 1 19656
box -48 -56 144 834
use sg13g2_decap_4  FILLER_24_39
timestamp 1679577901
transform 1 0 4896 0 1 19656
box -48 -56 432 834
use sg13g2_decap_8  FILLER_24_47
timestamp 1679581782
transform 1 0 5664 0 1 19656
box -48 -56 720 834
use sg13g2_decap_4  FILLER_24_54
timestamp 1679577901
transform 1 0 6336 0 1 19656
box -48 -56 432 834
use sg13g2_fill_2  FILLER_24_58
timestamp 1677580104
transform 1 0 6720 0 1 19656
box -48 -56 240 834
use sg13g2_decap_4  FILLER_24_64
timestamp 1679577901
transform 1 0 7296 0 1 19656
box -48 -56 432 834
use sg13g2_fill_2  FILLER_24_68
timestamp 1677580104
transform 1 0 7680 0 1 19656
box -48 -56 240 834
use sg13g2_fill_2  FILLER_24_116
timestamp 1677580104
transform 1 0 12288 0 1 19656
box -48 -56 240 834
use sg13g2_fill_1  FILLER_24_118
timestamp 1677579658
transform 1 0 12480 0 1 19656
box -48 -56 144 834
use sg13g2_decap_4  FILLER_25_4
timestamp 1679577901
transform 1 0 1536 0 -1 21168
box -48 -56 432 834
use sg13g2_fill_2  FILLER_25_8
timestamp 1677580104
transform 1 0 1920 0 -1 21168
box -48 -56 240 834
use sg13g2_fill_2  FILLER_25_65
timestamp 1677580104
transform 1 0 7392 0 -1 21168
box -48 -56 240 834
use sg13g2_fill_1  FILLER_25_67
timestamp 1677579658
transform 1 0 7584 0 -1 21168
box -48 -56 144 834
use sg13g2_fill_2  FILLER_25_72
timestamp 1677580104
transform 1 0 8064 0 -1 21168
box -48 -56 240 834
use sg13g2_fill_1  FILLER_25_74
timestamp 1677579658
transform 1 0 8256 0 -1 21168
box -48 -56 144 834
use sg13g2_decap_4  FILLER_25_79
timestamp 1679577901
transform 1 0 8736 0 -1 21168
box -48 -56 432 834
use sg13g2_fill_1  FILLER_25_110
timestamp 1677579658
transform 1 0 11712 0 -1 21168
box -48 -56 144 834
use sg13g2_decap_8  FILLER_26_0
timestamp 1679581782
transform 1 0 1152 0 1 21168
box -48 -56 720 834
use sg13g2_decap_4  FILLER_26_7
timestamp 1679577901
transform 1 0 1824 0 1 21168
box -48 -56 432 834
use sg13g2_fill_1  FILLER_26_32
timestamp 1677579658
transform 1 0 4224 0 1 21168
box -48 -56 144 834
use sg13g2_decap_4  FILLER_26_75
timestamp 1679577901
transform 1 0 8352 0 1 21168
box -48 -56 432 834
use sg13g2_fill_1  FILLER_26_79
timestamp 1677579658
transform 1 0 8736 0 1 21168
box -48 -56 144 834
use sg13g2_fill_2  FILLER_26_117
timestamp 1677580104
transform 1 0 12384 0 1 21168
box -48 -56 240 834
use sg13g2_decap_8  FILLER_27_4
timestamp 1679581782
transform 1 0 1536 0 -1 22680
box -48 -56 720 834
use sg13g2_decap_4  FILLER_27_11
timestamp 1679577901
transform 1 0 2208 0 -1 22680
box -48 -56 432 834
use sg13g2_fill_2  FILLER_27_15
timestamp 1677580104
transform 1 0 2592 0 -1 22680
box -48 -56 240 834
use sg13g2_fill_2  FILLER_27_117
timestamp 1677580104
transform 1 0 12384 0 -1 22680
box -48 -56 240 834
use sg13g2_decap_8  FILLER_28_4
timestamp 1679581782
transform 1 0 1536 0 1 22680
box -48 -56 720 834
use sg13g2_fill_2  FILLER_28_11
timestamp 1677580104
transform 1 0 2208 0 1 22680
box -48 -56 240 834
use sg13g2_decap_8  FILLER_28_55
timestamp 1679581782
transform 1 0 6432 0 1 22680
box -48 -56 720 834
use sg13g2_decap_4  FILLER_28_62
timestamp 1679577901
transform 1 0 7104 0 1 22680
box -48 -56 432 834
use sg13g2_fill_1  FILLER_28_99
timestamp 1677579658
transform 1 0 10656 0 1 22680
box -48 -56 144 834
use sg13g2_fill_2  FILLER_28_117
timestamp 1677580104
transform 1 0 12384 0 1 22680
box -48 -56 240 834
use sg13g2_decap_8  FILLER_29_4
timestamp 1679581782
transform 1 0 1536 0 -1 24192
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_11
timestamp 1679581782
transform 1 0 2208 0 -1 24192
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_18
timestamp 1679581782
transform 1 0 2880 0 -1 24192
box -48 -56 720 834
use sg13g2_decap_4  FILLER_29_25
timestamp 1679577901
transform 1 0 3552 0 -1 24192
box -48 -56 432 834
use sg13g2_fill_1  FILLER_29_29
timestamp 1677579658
transform 1 0 3936 0 -1 24192
box -48 -56 144 834
use sg13g2_decap_4  FILLER_29_64
timestamp 1679577901
transform 1 0 7296 0 -1 24192
box -48 -56 432 834
use sg13g2_fill_2  FILLER_29_93
timestamp 1677580104
transform 1 0 10080 0 -1 24192
box -48 -56 240 834
use sg13g2_fill_1  FILLER_29_95
timestamp 1677579658
transform 1 0 10272 0 -1 24192
box -48 -56 144 834
use sg13g2_fill_2  FILLER_29_117
timestamp 1677580104
transform 1 0 12384 0 -1 24192
box -48 -56 240 834
use sg13g2_decap_8  FILLER_30_0
timestamp 1679581782
transform 1 0 1152 0 1 24192
box -48 -56 720 834
use sg13g2_fill_2  FILLER_30_7
timestamp 1677580104
transform 1 0 1824 0 1 24192
box -48 -56 240 834
use sg13g2_fill_1  FILLER_30_9
timestamp 1677579658
transform 1 0 2016 0 1 24192
box -48 -56 144 834
use sg13g2_decap_8  FILLER_30_27
timestamp 1679581782
transform 1 0 3744 0 1 24192
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_38
timestamp 1679581782
transform 1 0 4800 0 1 24192
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_45
timestamp 1679581782
transform 1 0 5472 0 1 24192
box -48 -56 720 834
use sg13g2_decap_4  FILLER_30_52
timestamp 1679577901
transform 1 0 6144 0 1 24192
box -48 -56 432 834
use sg13g2_fill_2  FILLER_30_56
timestamp 1677580104
transform 1 0 6528 0 1 24192
box -48 -56 240 834
use sg13g2_fill_2  FILLER_30_96
timestamp 1677580104
transform 1 0 10368 0 1 24192
box -48 -56 240 834
use sg13g2_decap_8  FILLER_31_8
timestamp 1679581782
transform 1 0 1920 0 -1 25704
box -48 -56 720 834
use sg13g2_fill_1  FILLER_31_15
timestamp 1677579658
transform 1 0 2592 0 -1 25704
box -48 -56 144 834
use sg13g2_fill_2  FILLER_31_33
timestamp 1677580104
transform 1 0 4320 0 -1 25704
box -48 -56 240 834
use sg13g2_fill_1  FILLER_31_35
timestamp 1677579658
transform 1 0 4512 0 -1 25704
box -48 -56 144 834
use sg13g2_fill_1  FILLER_31_70
timestamp 1677579658
transform 1 0 7872 0 -1 25704
box -48 -56 144 834
use sg13g2_fill_2  FILLER_31_86
timestamp 1677580104
transform 1 0 9408 0 -1 25704
box -48 -56 240 834
use sg13g2_fill_1  FILLER_31_88
timestamp 1677579658
transform 1 0 9600 0 -1 25704
box -48 -56 144 834
use sg13g2_fill_1  FILLER_31_106
timestamp 1677579658
transform 1 0 11328 0 -1 25704
box -48 -56 144 834
use sg13g2_decap_4  FILLER_32_38
timestamp 1679577901
transform 1 0 4800 0 1 25704
box -48 -56 432 834
use sg13g2_decap_8  FILLER_32_81
timestamp 1679581782
transform 1 0 8928 0 1 25704
box -48 -56 720 834
use sg13g2_fill_2  FILLER_32_88
timestamp 1677580104
transform 1 0 9600 0 1 25704
box -48 -56 240 834
use sg13g2_decap_8  FILLER_33_4
timestamp 1679581782
transform 1 0 1536 0 -1 27216
box -48 -56 720 834
use sg13g2_decap_4  FILLER_33_11
timestamp 1679577901
transform 1 0 2208 0 -1 27216
box -48 -56 432 834
use sg13g2_decap_4  FILLER_33_57
timestamp 1679577901
transform 1 0 6624 0 -1 27216
box -48 -56 432 834
use sg13g2_fill_2  FILLER_33_61
timestamp 1677580104
transform 1 0 7008 0 -1 27216
box -48 -56 240 834
use sg13g2_decap_8  FILLER_33_68
timestamp 1679581782
transform 1 0 7680 0 -1 27216
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_75
timestamp 1679581782
transform 1 0 8352 0 -1 27216
box -48 -56 720 834
use sg13g2_decap_4  FILLER_33_82
timestamp 1679577901
transform 1 0 9024 0 -1 27216
box -48 -56 432 834
use sg13g2_fill_2  FILLER_33_86
timestamp 1677580104
transform 1 0 9408 0 -1 27216
box -48 -56 240 834
use sg13g2_fill_2  FILLER_33_117
timestamp 1677580104
transform 1 0 12384 0 -1 27216
box -48 -56 240 834
use sg13g2_decap_8  FILLER_34_0
timestamp 1679581782
transform 1 0 1152 0 1 27216
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_7
timestamp 1679581782
transform 1 0 1824 0 1 27216
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_14
timestamp 1679581782
transform 1 0 2496 0 1 27216
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_21
timestamp 1679581782
transform 1 0 3168 0 1 27216
box -48 -56 720 834
use sg13g2_decap_4  FILLER_34_28
timestamp 1679577901
transform 1 0 3840 0 1 27216
box -48 -56 432 834
use sg13g2_decap_8  FILLER_34_49
timestamp 1679581782
transform 1 0 5856 0 1 27216
box -48 -56 720 834
use sg13g2_fill_2  FILLER_34_56
timestamp 1677580104
transform 1 0 6528 0 1 27216
box -48 -56 240 834
use sg13g2_fill_2  FILLER_34_75
timestamp 1677580104
transform 1 0 8352 0 1 27216
box -48 -56 240 834
use sg13g2_fill_1  FILLER_34_77
timestamp 1677579658
transform 1 0 8544 0 1 27216
box -48 -56 144 834
use sg13g2_fill_2  FILLER_34_116
timestamp 1677580104
transform 1 0 12288 0 1 27216
box -48 -56 240 834
use sg13g2_fill_1  FILLER_34_118
timestamp 1677579658
transform 1 0 12480 0 1 27216
box -48 -56 144 834
use sg13g2_decap_8  FILLER_35_4
timestamp 1679581782
transform 1 0 1536 0 -1 28728
box -48 -56 720 834
use sg13g2_fill_2  FILLER_35_11
timestamp 1677580104
transform 1 0 2208 0 -1 28728
box -48 -56 240 834
use sg13g2_fill_1  FILLER_35_13
timestamp 1677579658
transform 1 0 2400 0 -1 28728
box -48 -56 144 834
use sg13g2_decap_8  FILLER_35_31
timestamp 1679581782
transform 1 0 4128 0 -1 28728
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_38
timestamp 1679581782
transform 1 0 4800 0 -1 28728
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_45
timestamp 1679581782
transform 1 0 5472 0 -1 28728
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_52
timestamp 1679581782
transform 1 0 6144 0 -1 28728
box -48 -56 720 834
use sg13g2_fill_1  FILLER_35_118
timestamp 1677579658
transform 1 0 12480 0 -1 28728
box -48 -56 144 834
use sg13g2_decap_8  FILLER_36_4
timestamp 1679581782
transform 1 0 1536 0 1 28728
box -48 -56 720 834
use sg13g2_fill_1  FILLER_36_11
timestamp 1677579658
transform 1 0 2208 0 1 28728
box -48 -56 144 834
use sg13g2_decap_4  FILLER_36_16
timestamp 1679577901
transform 1 0 2688 0 1 28728
box -48 -56 432 834
use sg13g2_decap_4  FILLER_36_37
timestamp 1679577901
transform 1 0 4704 0 1 28728
box -48 -56 432 834
use sg13g2_fill_2  FILLER_36_41
timestamp 1677580104
transform 1 0 5088 0 1 28728
box -48 -56 240 834
use sg13g2_fill_2  FILLER_36_51
timestamp 1677580104
transform 1 0 6048 0 1 28728
box -48 -56 240 834
use sg13g2_fill_1  FILLER_36_53
timestamp 1677579658
transform 1 0 6240 0 1 28728
box -48 -56 144 834
use sg13g2_fill_1  FILLER_36_88
timestamp 1677579658
transform 1 0 9600 0 1 28728
box -48 -56 144 834
use sg13g2_fill_1  FILLER_36_110
timestamp 1677579658
transform 1 0 11712 0 1 28728
box -48 -56 144 834
use sg13g2_decap_8  FILLER_37_4
timestamp 1679581782
transform 1 0 1536 0 -1 30240
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_11
timestamp 1679581782
transform 1 0 2208 0 -1 30240
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_18
timestamp 1679581782
transform 1 0 2880 0 -1 30240
box -48 -56 720 834
use sg13g2_decap_4  FILLER_37_25
timestamp 1679577901
transform 1 0 3552 0 -1 30240
box -48 -56 432 834
use sg13g2_decap_8  FILLER_37_75
timestamp 1679581782
transform 1 0 8352 0 -1 30240
box -48 -56 720 834
use sg13g2_fill_2  FILLER_37_82
timestamp 1677580104
transform 1 0 9024 0 -1 30240
box -48 -56 240 834
use sg13g2_fill_1  FILLER_37_84
timestamp 1677579658
transform 1 0 9216 0 -1 30240
box -48 -56 144 834
use sg13g2_decap_8  FILLER_38_0
timestamp 1679581782
transform 1 0 1152 0 1 30240
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_7
timestamp 1679581782
transform 1 0 1824 0 1 30240
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_14
timestamp 1679581782
transform 1 0 2496 0 1 30240
box -48 -56 720 834
use sg13g2_fill_2  FILLER_38_21
timestamp 1677580104
transform 1 0 3168 0 1 30240
box -48 -56 240 834
use sg13g2_fill_1  FILLER_38_110
timestamp 1677579658
transform 1 0 11712 0 1 30240
box -48 -56 144 834
use sg13g2_decap_8  FILLER_39_4
timestamp 1679581782
transform 1 0 1536 0 -1 31752
box -48 -56 720 834
use sg13g2_decap_4  FILLER_39_11
timestamp 1679577901
transform 1 0 2208 0 -1 31752
box -48 -56 432 834
use sg13g2_fill_2  FILLER_39_15
timestamp 1677580104
transform 1 0 2592 0 -1 31752
box -48 -56 240 834
use sg13g2_fill_1  FILLER_39_63
timestamp 1677579658
transform 1 0 7200 0 -1 31752
box -48 -56 144 834
use sg13g2_fill_2  FILLER_39_85
timestamp 1677580104
transform 1 0 9312 0 -1 31752
box -48 -56 240 834
use sg13g2_fill_2  FILLER_39_104
timestamp 1677580104
transform 1 0 11136 0 -1 31752
box -48 -56 240 834
use sg13g2_fill_1  FILLER_39_106
timestamp 1677579658
transform 1 0 11328 0 -1 31752
box -48 -56 144 834
use sg13g2_decap_8  FILLER_40_4
timestamp 1679581782
transform 1 0 1536 0 1 31752
box -48 -56 720 834
use sg13g2_decap_4  FILLER_40_11
timestamp 1679577901
transform 1 0 2208 0 1 31752
box -48 -56 432 834
use sg13g2_decap_8  FILLER_40_57
timestamp 1679581782
transform 1 0 6624 0 1 31752
box -48 -56 720 834
use sg13g2_decap_4  FILLER_40_64
timestamp 1679577901
transform 1 0 7296 0 1 31752
box -48 -56 432 834
use sg13g2_fill_2  FILLER_40_68
timestamp 1677580104
transform 1 0 7680 0 1 31752
box -48 -56 240 834
use sg13g2_fill_2  FILLER_40_91
timestamp 1677580104
transform 1 0 9888 0 1 31752
box -48 -56 240 834
use sg13g2_decap_8  FILLER_41_4
timestamp 1679581782
transform 1 0 1536 0 -1 33264
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_11
timestamp 1679581782
transform 1 0 2208 0 -1 33264
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_18
timestamp 1679581782
transform 1 0 2880 0 -1 33264
box -48 -56 720 834
use sg13g2_fill_1  FILLER_41_25
timestamp 1677579658
transform 1 0 3552 0 -1 33264
box -48 -56 144 834
use sg13g2_fill_2  FILLER_41_63
timestamp 1677580104
transform 1 0 7200 0 -1 33264
box -48 -56 240 834
use sg13g2_fill_1  FILLER_41_65
timestamp 1677579658
transform 1 0 7392 0 -1 33264
box -48 -56 144 834
use sg13g2_fill_2  FILLER_41_108
timestamp 1677580104
transform 1 0 11520 0 -1 33264
box -48 -56 240 834
use sg13g2_fill_1  FILLER_41_110
timestamp 1677579658
transform 1 0 11712 0 -1 33264
box -48 -56 144 834
use sg13g2_decap_8  FILLER_42_0
timestamp 1679581782
transform 1 0 1152 0 1 33264
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_7
timestamp 1679581782
transform 1 0 1824 0 1 33264
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_14
timestamp 1679581782
transform 1 0 2496 0 1 33264
box -48 -56 720 834
use sg13g2_fill_1  FILLER_42_21
timestamp 1677579658
transform 1 0 3168 0 1 33264
box -48 -56 144 834
use sg13g2_decap_8  FILLER_42_39
timestamp 1679581782
transform 1 0 4896 0 1 33264
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_46
timestamp 1679581782
transform 1 0 5568 0 1 33264
box -48 -56 720 834
use sg13g2_fill_1  FILLER_42_82
timestamp 1677579658
transform 1 0 9024 0 1 33264
box -48 -56 144 834
use sg13g2_fill_2  FILLER_42_108
timestamp 1677580104
transform 1 0 11520 0 1 33264
box -48 -56 240 834
use sg13g2_fill_1  FILLER_42_110
timestamp 1677579658
transform 1 0 11712 0 1 33264
box -48 -56 144 834
use sg13g2_decap_8  FILLER_43_4
timestamp 1679581782
transform 1 0 1536 0 -1 34776
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_11
timestamp 1679581782
transform 1 0 2208 0 -1 34776
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_18
timestamp 1679581782
transform 1 0 2880 0 -1 34776
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_25
timestamp 1679581782
transform 1 0 3552 0 -1 34776
box -48 -56 720 834
use sg13g2_fill_2  FILLER_43_32
timestamp 1677580104
transform 1 0 4224 0 -1 34776
box -48 -56 240 834
use sg13g2_fill_1  FILLER_43_110
timestamp 1677579658
transform 1 0 11712 0 -1 34776
box -48 -56 144 834
use sg13g2_decap_8  FILLER_44_4
timestamp 1679581782
transform 1 0 1536 0 1 34776
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_11
timestamp 1679581782
transform 1 0 2208 0 1 34776
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_18
timestamp 1679581782
transform 1 0 2880 0 1 34776
box -48 -56 720 834
use sg13g2_fill_2  FILLER_44_25
timestamp 1677580104
transform 1 0 3552 0 1 34776
box -48 -56 240 834
use sg13g2_fill_1  FILLER_44_27
timestamp 1677579658
transform 1 0 3744 0 1 34776
box -48 -56 144 834
use sg13g2_decap_8  FILLER_44_49
timestamp 1679581782
transform 1 0 5856 0 1 34776
box -48 -56 720 834
use sg13g2_decap_4  FILLER_44_56
timestamp 1679577901
transform 1 0 6528 0 1 34776
box -48 -56 432 834
use sg13g2_decap_8  FILLER_45_4
timestamp 1679581782
transform 1 0 1536 0 -1 36288
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_11
timestamp 1679581782
transform 1 0 2208 0 -1 36288
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_18
timestamp 1679581782
transform 1 0 2880 0 -1 36288
box -48 -56 720 834
use sg13g2_decap_4  FILLER_45_25
timestamp 1679577901
transform 1 0 3552 0 -1 36288
box -48 -56 432 834
use sg13g2_fill_1  FILLER_45_29
timestamp 1677579658
transform 1 0 3936 0 -1 36288
box -48 -56 144 834
use sg13g2_decap_8  FILLER_45_59
timestamp 1679581782
transform 1 0 6816 0 -1 36288
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_66
timestamp 1679581782
transform 1 0 7488 0 -1 36288
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_73
timestamp 1679581782
transform 1 0 8160 0 -1 36288
box -48 -56 720 834
use sg13g2_fill_2  FILLER_45_80
timestamp 1677580104
transform 1 0 8832 0 -1 36288
box -48 -56 240 834
use sg13g2_fill_1  FILLER_45_82
timestamp 1677579658
transform 1 0 9024 0 -1 36288
box -48 -56 144 834
use sg13g2_fill_2  FILLER_45_112
timestamp 1677580104
transform 1 0 11904 0 -1 36288
box -48 -56 240 834
use sg13g2_fill_1  FILLER_45_114
timestamp 1677579658
transform 1 0 12096 0 -1 36288
box -48 -56 144 834
use sg13g2_decap_8  FILLER_46_0
timestamp 1679581782
transform 1 0 1152 0 1 36288
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_7
timestamp 1679581782
transform 1 0 1824 0 1 36288
box -48 -56 720 834
use sg13g2_decap_4  FILLER_46_14
timestamp 1679577901
transform 1 0 2496 0 1 36288
box -48 -56 432 834
use sg13g2_fill_2  FILLER_46_18
timestamp 1677580104
transform 1 0 2880 0 1 36288
box -48 -56 240 834
use sg13g2_decap_8  FILLER_46_71
timestamp 1679581782
transform 1 0 7968 0 1 36288
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_78
timestamp 1679581782
transform 1 0 8640 0 1 36288
box -48 -56 720 834
use sg13g2_fill_1  FILLER_46_85
timestamp 1677579658
transform 1 0 9312 0 1 36288
box -48 -56 144 834
use sg13g2_decap_8  FILLER_47_4
timestamp 1679581782
transform 1 0 1536 0 -1 37800
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_11
timestamp 1679581782
transform 1 0 2208 0 -1 37800
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_18
timestamp 1679581782
transform 1 0 2880 0 -1 37800
box -48 -56 720 834
use sg13g2_fill_1  FILLER_47_25
timestamp 1677579658
transform 1 0 3552 0 -1 37800
box -48 -56 144 834
use sg13g2_fill_1  FILLER_47_81
timestamp 1677579658
transform 1 0 8928 0 -1 37800
box -48 -56 144 834
use sg13g2_decap_8  FILLER_48_4
timestamp 1679581782
transform 1 0 1536 0 1 37800
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_11
timestamp 1679581782
transform 1 0 2208 0 1 37800
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_18
timestamp 1679581782
transform 1 0 2880 0 1 37800
box -48 -56 720 834
use sg13g2_fill_2  FILLER_48_25
timestamp 1677580104
transform 1 0 3552 0 1 37800
box -48 -56 240 834
use sg13g2_fill_2  FILLER_48_99
timestamp 1677580104
transform 1 0 10656 0 1 37800
box -48 -56 240 834
use sg13g2_fill_1  FILLER_48_101
timestamp 1677579658
transform 1 0 10848 0 1 37800
box -48 -56 144 834
use sg13g2_fill_1  FILLER_48_106
timestamp 1677579658
transform 1 0 11328 0 1 37800
box -48 -56 144 834
use sg13g2_decap_8  FILLER_49_4
timestamp 1679581782
transform 1 0 1536 0 -1 39312
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_11
timestamp 1679581782
transform 1 0 2208 0 -1 39312
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_18
timestamp 1679581782
transform 1 0 2880 0 -1 39312
box -48 -56 720 834
use sg13g2_decap_4  FILLER_49_25
timestamp 1679577901
transform 1 0 3552 0 -1 39312
box -48 -56 432 834
use sg13g2_fill_2  FILLER_49_29
timestamp 1677580104
transform 1 0 3936 0 -1 39312
box -48 -56 240 834
use sg13g2_decap_8  FILLER_49_89
timestamp 1679581782
transform 1 0 9696 0 -1 39312
box -48 -56 720 834
use sg13g2_fill_2  FILLER_49_96
timestamp 1677580104
transform 1 0 10368 0 -1 39312
box -48 -56 240 834
use sg13g2_fill_1  FILLER_49_98
timestamp 1677579658
transform 1 0 10560 0 -1 39312
box -48 -56 144 834
use sg13g2_decap_8  FILLER_50_0
timestamp 1679581782
transform 1 0 1152 0 1 39312
box -48 -56 720 834
use sg13g2_decap_8  FILLER_50_7
timestamp 1679581782
transform 1 0 1824 0 1 39312
box -48 -56 720 834
use sg13g2_decap_8  FILLER_50_14
timestamp 1679581782
transform 1 0 2496 0 1 39312
box -48 -56 720 834
use sg13g2_decap_8  FILLER_50_21
timestamp 1679581782
transform 1 0 3168 0 1 39312
box -48 -56 720 834
use sg13g2_decap_8  FILLER_50_28
timestamp 1679581782
transform 1 0 3840 0 1 39312
box -48 -56 720 834
use sg13g2_decap_8  FILLER_50_35
timestamp 1679581782
transform 1 0 4512 0 1 39312
box -48 -56 720 834
use sg13g2_decap_8  FILLER_50_42
timestamp 1679581782
transform 1 0 5184 0 1 39312
box -48 -56 720 834
use sg13g2_decap_8  FILLER_50_83
timestamp 1679581782
transform 1 0 9120 0 1 39312
box -48 -56 720 834
use sg13g2_decap_8  FILLER_50_90
timestamp 1679581782
transform 1 0 9792 0 1 39312
box -48 -56 720 834
use sg13g2_decap_4  FILLER_50_97
timestamp 1679577901
transform 1 0 10464 0 1 39312
box -48 -56 432 834
use sg13g2_fill_2  FILLER_50_101
timestamp 1677580104
transform 1 0 10848 0 1 39312
box -48 -56 240 834
use sg13g2_decap_8  FILLER_51_4
timestamp 1679581782
transform 1 0 1536 0 -1 40824
box -48 -56 720 834
use sg13g2_decap_8  FILLER_51_11
timestamp 1679581782
transform 1 0 2208 0 -1 40824
box -48 -56 720 834
use sg13g2_decap_8  FILLER_51_18
timestamp 1679581782
transform 1 0 2880 0 -1 40824
box -48 -56 720 834
use sg13g2_decap_8  FILLER_51_25
timestamp 1679581782
transform 1 0 3552 0 -1 40824
box -48 -56 720 834
use sg13g2_decap_8  FILLER_51_32
timestamp 1679581782
transform 1 0 4224 0 -1 40824
box -48 -56 720 834
use sg13g2_decap_8  FILLER_51_39
timestamp 1679581782
transform 1 0 4896 0 -1 40824
box -48 -56 720 834
use sg13g2_decap_8  FILLER_51_46
timestamp 1679581782
transform 1 0 5568 0 -1 40824
box -48 -56 720 834
use sg13g2_decap_8  FILLER_51_53
timestamp 1679581782
transform 1 0 6240 0 -1 40824
box -48 -56 720 834
use sg13g2_decap_8  FILLER_51_60
timestamp 1679581782
transform 1 0 6912 0 -1 40824
box -48 -56 720 834
use sg13g2_decap_8  FILLER_51_67
timestamp 1679581782
transform 1 0 7584 0 -1 40824
box -48 -56 720 834
use sg13g2_decap_8  FILLER_51_74
timestamp 1679581782
transform 1 0 8256 0 -1 40824
box -48 -56 720 834
use sg13g2_decap_8  FILLER_51_81
timestamp 1679581782
transform 1 0 8928 0 -1 40824
box -48 -56 720 834
use sg13g2_decap_8  FILLER_51_88
timestamp 1679581782
transform 1 0 9600 0 -1 40824
box -48 -56 720 834
use sg13g2_decap_8  FILLER_51_95
timestamp 1679581782
transform 1 0 10272 0 -1 40824
box -48 -56 720 834
use sg13g2_decap_4  FILLER_51_102
timestamp 1679577901
transform 1 0 10944 0 -1 40824
box -48 -56 432 834
use sg13g2_fill_1  FILLER_51_106
timestamp 1677579658
transform 1 0 11328 0 -1 40824
box -48 -56 144 834
use sg13g2_decap_8  FILLER_52_4
timestamp 1679581782
transform 1 0 1536 0 1 40824
box -48 -56 720 834
use sg13g2_decap_8  FILLER_52_11
timestamp 1679581782
transform 1 0 2208 0 1 40824
box -48 -56 720 834
use sg13g2_decap_8  FILLER_52_18
timestamp 1679581782
transform 1 0 2880 0 1 40824
box -48 -56 720 834
use sg13g2_decap_8  FILLER_52_25
timestamp 1679581782
transform 1 0 3552 0 1 40824
box -48 -56 720 834
use sg13g2_decap_8  FILLER_52_32
timestamp 1679581782
transform 1 0 4224 0 1 40824
box -48 -56 720 834
use sg13g2_decap_8  FILLER_52_39
timestamp 1679581782
transform 1 0 4896 0 1 40824
box -48 -56 720 834
use sg13g2_decap_8  FILLER_52_46
timestamp 1679581782
transform 1 0 5568 0 1 40824
box -48 -56 720 834
use sg13g2_decap_8  FILLER_52_53
timestamp 1679581782
transform 1 0 6240 0 1 40824
box -48 -56 720 834
use sg13g2_decap_8  FILLER_52_60
timestamp 1679581782
transform 1 0 6912 0 1 40824
box -48 -56 720 834
use sg13g2_decap_8  FILLER_52_67
timestamp 1679581782
transform 1 0 7584 0 1 40824
box -48 -56 720 834
use sg13g2_decap_8  FILLER_52_74
timestamp 1679581782
transform 1 0 8256 0 1 40824
box -48 -56 720 834
use sg13g2_decap_8  FILLER_52_81
timestamp 1679581782
transform 1 0 8928 0 1 40824
box -48 -56 720 834
use sg13g2_decap_8  FILLER_52_88
timestamp 1679581782
transform 1 0 9600 0 1 40824
box -48 -56 720 834
use sg13g2_decap_8  FILLER_52_95
timestamp 1679581782
transform 1 0 10272 0 1 40824
box -48 -56 720 834
use sg13g2_decap_4  FILLER_52_102
timestamp 1679577901
transform 1 0 10944 0 1 40824
box -48 -56 432 834
use sg13g2_fill_1  FILLER_52_106
timestamp 1677579658
transform 1 0 11328 0 1 40824
box -48 -56 144 834
use sg13g2_decap_8  FILLER_53_4
timestamp 1679581782
transform 1 0 1536 0 -1 42336
box -48 -56 720 834
use sg13g2_decap_8  FILLER_53_11
timestamp 1679581782
transform 1 0 2208 0 -1 42336
box -48 -56 720 834
use sg13g2_decap_8  FILLER_53_18
timestamp 1679581782
transform 1 0 2880 0 -1 42336
box -48 -56 720 834
use sg13g2_decap_8  FILLER_53_25
timestamp 1679581782
transform 1 0 3552 0 -1 42336
box -48 -56 720 834
use sg13g2_decap_8  FILLER_53_32
timestamp 1679581782
transform 1 0 4224 0 -1 42336
box -48 -56 720 834
use sg13g2_decap_8  FILLER_53_39
timestamp 1679581782
transform 1 0 4896 0 -1 42336
box -48 -56 720 834
use sg13g2_decap_8  FILLER_53_46
timestamp 1679581782
transform 1 0 5568 0 -1 42336
box -48 -56 720 834
use sg13g2_decap_8  FILLER_53_53
timestamp 1679581782
transform 1 0 6240 0 -1 42336
box -48 -56 720 834
use sg13g2_decap_8  FILLER_53_60
timestamp 1679581782
transform 1 0 6912 0 -1 42336
box -48 -56 720 834
use sg13g2_decap_8  FILLER_53_67
timestamp 1679581782
transform 1 0 7584 0 -1 42336
box -48 -56 720 834
use sg13g2_decap_8  FILLER_53_74
timestamp 1679581782
transform 1 0 8256 0 -1 42336
box -48 -56 720 834
use sg13g2_decap_8  FILLER_53_81
timestamp 1679581782
transform 1 0 8928 0 -1 42336
box -48 -56 720 834
use sg13g2_decap_8  FILLER_53_88
timestamp 1679581782
transform 1 0 9600 0 -1 42336
box -48 -56 720 834
use sg13g2_decap_8  FILLER_53_95
timestamp 1679581782
transform 1 0 10272 0 -1 42336
box -48 -56 720 834
use sg13g2_decap_8  FILLER_53_102
timestamp 1679581782
transform 1 0 10944 0 -1 42336
box -48 -56 720 834
use sg13g2_fill_2  FILLER_53_109
timestamp 1677580104
transform 1 0 11616 0 -1 42336
box -48 -56 240 834
use sg13g2_decap_8  FILLER_54_0
timestamp 1679581782
transform 1 0 1152 0 1 42336
box -48 -56 720 834
use sg13g2_decap_8  FILLER_54_7
timestamp 1679581782
transform 1 0 1824 0 1 42336
box -48 -56 720 834
use sg13g2_decap_8  FILLER_54_14
timestamp 1679581782
transform 1 0 2496 0 1 42336
box -48 -56 720 834
use sg13g2_decap_8  FILLER_54_21
timestamp 1679581782
transform 1 0 3168 0 1 42336
box -48 -56 720 834
use sg13g2_decap_8  FILLER_54_28
timestamp 1679581782
transform 1 0 3840 0 1 42336
box -48 -56 720 834
use sg13g2_decap_8  FILLER_54_35
timestamp 1679581782
transform 1 0 4512 0 1 42336
box -48 -56 720 834
use sg13g2_decap_8  FILLER_54_42
timestamp 1679581782
transform 1 0 5184 0 1 42336
box -48 -56 720 834
use sg13g2_decap_8  FILLER_54_49
timestamp 1679581782
transform 1 0 5856 0 1 42336
box -48 -56 720 834
use sg13g2_decap_8  FILLER_54_56
timestamp 1679581782
transform 1 0 6528 0 1 42336
box -48 -56 720 834
use sg13g2_decap_8  FILLER_54_63
timestamp 1679581782
transform 1 0 7200 0 1 42336
box -48 -56 720 834
use sg13g2_decap_8  FILLER_54_70
timestamp 1679581782
transform 1 0 7872 0 1 42336
box -48 -56 720 834
use sg13g2_decap_8  FILLER_54_77
timestamp 1679581782
transform 1 0 8544 0 1 42336
box -48 -56 720 834
use sg13g2_decap_8  FILLER_54_84
timestamp 1679581782
transform 1 0 9216 0 1 42336
box -48 -56 720 834
use sg13g2_decap_8  FILLER_54_91
timestamp 1679581782
transform 1 0 9888 0 1 42336
box -48 -56 720 834
use sg13g2_decap_4  FILLER_54_98
timestamp 1679577901
transform 1 0 10560 0 1 42336
box -48 -56 432 834
use sg13g2_fill_1  FILLER_54_114
timestamp 1677579658
transform 1 0 12096 0 1 42336
box -48 -56 144 834
use sg13g2_decap_8  FILLER_55_4
timestamp 1679581782
transform 1 0 1536 0 -1 43848
box -48 -56 720 834
use sg13g2_decap_8  FILLER_55_11
timestamp 1679581782
transform 1 0 2208 0 -1 43848
box -48 -56 720 834
use sg13g2_decap_8  FILLER_55_18
timestamp 1679581782
transform 1 0 2880 0 -1 43848
box -48 -56 720 834
use sg13g2_decap_8  FILLER_55_25
timestamp 1679581782
transform 1 0 3552 0 -1 43848
box -48 -56 720 834
use sg13g2_decap_8  FILLER_55_32
timestamp 1679581782
transform 1 0 4224 0 -1 43848
box -48 -56 720 834
use sg13g2_decap_8  FILLER_55_39
timestamp 1679581782
transform 1 0 4896 0 -1 43848
box -48 -56 720 834
use sg13g2_decap_8  FILLER_55_46
timestamp 1679581782
transform 1 0 5568 0 -1 43848
box -48 -56 720 834
use sg13g2_decap_8  FILLER_55_53
timestamp 1679581782
transform 1 0 6240 0 -1 43848
box -48 -56 720 834
use sg13g2_decap_8  FILLER_55_60
timestamp 1679581782
transform 1 0 6912 0 -1 43848
box -48 -56 720 834
use sg13g2_decap_8  FILLER_55_67
timestamp 1679581782
transform 1 0 7584 0 -1 43848
box -48 -56 720 834
use sg13g2_fill_1  FILLER_55_74
timestamp 1677579658
transform 1 0 8256 0 -1 43848
box -48 -56 144 834
use sg13g2_decap_8  FILLER_55_79
timestamp 1679581782
transform 1 0 8736 0 -1 43848
box -48 -56 720 834
use sg13g2_decap_8  FILLER_55_86
timestamp 1679581782
transform 1 0 9408 0 -1 43848
box -48 -56 720 834
use sg13g2_decap_8  FILLER_55_93
timestamp 1679581782
transform 1 0 10080 0 -1 43848
box -48 -56 720 834
use sg13g2_fill_2  FILLER_55_100
timestamp 1677580104
transform 1 0 10752 0 -1 43848
box -48 -56 240 834
use sg13g2_fill_1  FILLER_55_102
timestamp 1677579658
transform 1 0 10944 0 -1 43848
box -48 -56 144 834
use sg13g2_decap_8  FILLER_56_4
timestamp 1679581782
transform 1 0 1536 0 1 43848
box -48 -56 720 834
use sg13g2_decap_8  FILLER_56_11
timestamp 1679581782
transform 1 0 2208 0 1 43848
box -48 -56 720 834
use sg13g2_decap_8  FILLER_56_18
timestamp 1679581782
transform 1 0 2880 0 1 43848
box -48 -56 720 834
use sg13g2_decap_8  FILLER_56_25
timestamp 1679581782
transform 1 0 3552 0 1 43848
box -48 -56 720 834
use sg13g2_decap_8  FILLER_56_32
timestamp 1679581782
transform 1 0 4224 0 1 43848
box -48 -56 720 834
use sg13g2_decap_8  FILLER_56_39
timestamp 1679581782
transform 1 0 4896 0 1 43848
box -48 -56 720 834
use sg13g2_decap_8  FILLER_56_46
timestamp 1679581782
transform 1 0 5568 0 1 43848
box -48 -56 720 834
use sg13g2_decap_8  FILLER_56_53
timestamp 1679581782
transform 1 0 6240 0 1 43848
box -48 -56 720 834
use sg13g2_decap_8  FILLER_56_60
timestamp 1679581782
transform 1 0 6912 0 1 43848
box -48 -56 720 834
use sg13g2_decap_8  FILLER_56_67
timestamp 1679581782
transform 1 0 7584 0 1 43848
box -48 -56 720 834
use sg13g2_decap_8  FILLER_56_74
timestamp 1679581782
transform 1 0 8256 0 1 43848
box -48 -56 720 834
use sg13g2_decap_8  FILLER_56_81
timestamp 1679581782
transform 1 0 8928 0 1 43848
box -48 -56 720 834
use sg13g2_decap_8  FILLER_56_88
timestamp 1679581782
transform 1 0 9600 0 1 43848
box -48 -56 720 834
use sg13g2_fill_2  FILLER_56_95
timestamp 1677580104
transform 1 0 10272 0 1 43848
box -48 -56 240 834
use sg13g2_fill_2  FILLER_56_113
timestamp 1677580104
transform 1 0 12000 0 1 43848
box -48 -56 240 834
use sg13g2_decap_8  FILLER_57_4
timestamp 1679581782
transform 1 0 1536 0 -1 45360
box -48 -56 720 834
use sg13g2_decap_8  FILLER_57_11
timestamp 1679581782
transform 1 0 2208 0 -1 45360
box -48 -56 720 834
use sg13g2_decap_8  FILLER_57_18
timestamp 1679581782
transform 1 0 2880 0 -1 45360
box -48 -56 720 834
use sg13g2_decap_8  FILLER_57_25
timestamp 1679581782
transform 1 0 3552 0 -1 45360
box -48 -56 720 834
use sg13g2_fill_1  FILLER_57_32
timestamp 1677579658
transform 1 0 4224 0 -1 45360
box -48 -56 144 834
use sg13g2_decap_8  FILLER_57_37
timestamp 1679581782
transform 1 0 4704 0 -1 45360
box -48 -56 720 834
use sg13g2_decap_8  FILLER_57_48
timestamp 1679581782
transform 1 0 5760 0 -1 45360
box -48 -56 720 834
use sg13g2_decap_8  FILLER_57_55
timestamp 1679581782
transform 1 0 6432 0 -1 45360
box -48 -56 720 834
use sg13g2_decap_8  FILLER_57_62
timestamp 1679581782
transform 1 0 7104 0 -1 45360
box -48 -56 720 834
use sg13g2_decap_8  FILLER_57_69
timestamp 1679581782
transform 1 0 7776 0 -1 45360
box -48 -56 720 834
use sg13g2_fill_2  FILLER_57_76
timestamp 1677580104
transform 1 0 8448 0 -1 45360
box -48 -56 240 834
use sg13g2_decap_8  FILLER_57_82
timestamp 1679581782
transform 1 0 9024 0 -1 45360
box -48 -56 720 834
use sg13g2_decap_4  FILLER_57_89
timestamp 1679577901
transform 1 0 9696 0 -1 45360
box -48 -56 432 834
use sg13g2_fill_2  FILLER_57_93
timestamp 1677580104
transform 1 0 10080 0 -1 45360
box -48 -56 240 834
use sg13g2_fill_2  FILLER_57_103
timestamp 1677580104
transform 1 0 11040 0 -1 45360
box -48 -56 240 834
use sg13g2_fill_2  FILLER_57_117
timestamp 1677580104
transform 1 0 12384 0 -1 45360
box -48 -56 240 834
use sg13g2_decap_8  FILLER_58_8
timestamp 1679581782
transform 1 0 1920 0 1 45360
box -48 -56 720 834
use sg13g2_decap_8  FILLER_58_15
timestamp 1679581782
transform 1 0 2592 0 1 45360
box -48 -56 720 834
use sg13g2_decap_8  FILLER_58_22
timestamp 1679581782
transform 1 0 3264 0 1 45360
box -48 -56 720 834
use sg13g2_decap_8  FILLER_58_29
timestamp 1679581782
transform 1 0 3936 0 1 45360
box -48 -56 720 834
use sg13g2_decap_8  FILLER_58_36
timestamp 1679581782
transform 1 0 4608 0 1 45360
box -48 -56 720 834
use sg13g2_decap_8  FILLER_58_43
timestamp 1679581782
transform 1 0 5280 0 1 45360
box -48 -56 720 834
use sg13g2_decap_8  FILLER_58_50
timestamp 1679581782
transform 1 0 5952 0 1 45360
box -48 -56 720 834
use sg13g2_decap_8  FILLER_58_57
timestamp 1679581782
transform 1 0 6624 0 1 45360
box -48 -56 720 834
use sg13g2_decap_8  FILLER_58_64
timestamp 1679581782
transform 1 0 7296 0 1 45360
box -48 -56 720 834
use sg13g2_decap_8  FILLER_58_71
timestamp 1679581782
transform 1 0 7968 0 1 45360
box -48 -56 720 834
use sg13g2_decap_8  FILLER_58_78
timestamp 1679581782
transform 1 0 8640 0 1 45360
box -48 -56 720 834
use sg13g2_decap_8  FILLER_58_85
timestamp 1679581782
transform 1 0 9312 0 1 45360
box -48 -56 720 834
use sg13g2_fill_1  FILLER_58_92
timestamp 1677579658
transform 1 0 9984 0 1 45360
box -48 -56 144 834
use sg13g2_fill_2  FILLER_58_109
timestamp 1677580104
transform 1 0 11616 0 1 45360
box -48 -56 240 834
use sg13g2_fill_1  FILLER_59_4
timestamp 1677579658
transform 1 0 1536 0 -1 46872
box -48 -56 144 834
use sg13g2_fill_2  FILLER_59_9
timestamp 1677580104
transform 1 0 2016 0 -1 46872
box -48 -56 240 834
use sg13g2_fill_2  FILLER_59_15
timestamp 1677580104
transform 1 0 2592 0 -1 46872
box -48 -56 240 834
use sg13g2_fill_2  FILLER_59_21
timestamp 1677580104
transform 1 0 3168 0 -1 46872
box -48 -56 240 834
use sg13g2_fill_2  FILLER_59_27
timestamp 1677580104
transform 1 0 3744 0 -1 46872
box -48 -56 240 834
use sg13g2_fill_2  FILLER_59_33
timestamp 1677580104
transform 1 0 4320 0 -1 46872
box -48 -56 240 834
use sg13g2_fill_2  FILLER_59_39
timestamp 1677580104
transform 1 0 4896 0 -1 46872
box -48 -56 240 834
use sg13g2_fill_2  FILLER_59_45
timestamp 1677580104
transform 1 0 5472 0 -1 46872
box -48 -56 240 834
use sg13g2_fill_2  FILLER_59_51
timestamp 1677580104
transform 1 0 6048 0 -1 46872
box -48 -56 240 834
use sg13g2_fill_2  FILLER_59_57
timestamp 1677580104
transform 1 0 6624 0 -1 46872
box -48 -56 240 834
use sg13g2_fill_2  FILLER_59_63
timestamp 1677580104
transform 1 0 7200 0 -1 46872
box -48 -56 240 834
use sg13g2_fill_2  FILLER_59_69
timestamp 1677580104
transform 1 0 7776 0 -1 46872
box -48 -56 240 834
use sg13g2_fill_2  FILLER_59_75
timestamp 1677580104
transform 1 0 8352 0 -1 46872
box -48 -56 240 834
use sg13g2_fill_2  FILLER_59_81
timestamp 1677580104
transform 1 0 8928 0 -1 46872
box -48 -56 240 834
use sg13g2_fill_2  FILLER_59_87
timestamp 1677580104
transform 1 0 9504 0 -1 46872
box -48 -56 240 834
use sg13g2_fill_2  FILLER_59_93
timestamp 1677580104
transform 1 0 10080 0 -1 46872
box -48 -56 240 834
use sg13g2_fill_2  FILLER_59_99
timestamp 1677580104
transform 1 0 10656 0 -1 46872
box -48 -56 240 834
use sg13g2_fill_2  FILLER_59_105
timestamp 1677580104
transform 1 0 11232 0 -1 46872
box -48 -56 240 834
use sg13g2_buf_1  input1
timestamp 1676381911
transform 1 0 1152 0 1 1512
box -48 -56 432 834
use sg13g2_buf_1  input2
timestamp 1676381911
transform 1 0 1152 0 1 4536
box -48 -56 432 834
use sg13g2_buf_1  input3
timestamp 1676381911
transform 1 0 1152 0 -1 16632
box -48 -56 432 834
use sg13g2_buf_1  input4
timestamp 1676381911
transform 1 0 1152 0 -1 25704
box -48 -56 432 834
use sg13g2_buf_1  input5
timestamp 1676381911
transform 1 0 1152 0 -1 27216
box -48 -56 432 834
use sg13g2_buf_1  input6
timestamp 1676381911
transform 1 0 1152 0 -1 28728
box -48 -56 432 834
use sg13g2_buf_1  input7
timestamp 1676381911
transform 1 0 1152 0 1 28728
box -48 -56 432 834
use sg13g2_buf_1  input8
timestamp 1676381911
transform 1 0 1152 0 -1 30240
box -48 -56 432 834
use sg13g2_buf_1  input9
timestamp 1676381911
transform 1 0 1152 0 -1 31752
box -48 -56 432 834
use sg13g2_buf_1  input10
timestamp 1676381911
transform 1 0 1152 0 1 31752
box -48 -56 432 834
use sg13g2_buf_1  input11
timestamp 1676381911
transform 1 0 1152 0 -1 33264
box -48 -56 432 834
use sg13g2_buf_1  input12
timestamp 1676381911
transform 1 0 1152 0 -1 34776
box -48 -56 432 834
use sg13g2_buf_1  input13
timestamp 1676381911
transform 1 0 1152 0 1 34776
box -48 -56 432 834
use sg13g2_buf_1  input14
timestamp 1676381911
transform 1 0 1152 0 1 16632
box -48 -56 432 834
use sg13g2_buf_1  input15
timestamp 1676381911
transform 1 0 1152 0 -1 36288
box -48 -56 432 834
use sg13g2_buf_1  input16
timestamp 1676381911
transform 1 0 1152 0 -1 37800
box -48 -56 432 834
use sg13g2_buf_1  input17
timestamp 1676381911
transform 1 0 1152 0 1 37800
box -48 -56 432 834
use sg13g2_buf_1  input18
timestamp 1676381911
transform 1 0 1152 0 -1 39312
box -48 -56 432 834
use sg13g2_buf_1  input19
timestamp 1676381911
transform 1 0 1152 0 -1 40824
box -48 -56 432 834
use sg13g2_buf_1  input20
timestamp 1676381911
transform 1 0 1152 0 1 40824
box -48 -56 432 834
use sg13g2_buf_1  input21
timestamp 1676381911
transform 1 0 1152 0 -1 42336
box -48 -56 432 834
use sg13g2_buf_1  input22
timestamp 1676381911
transform 1 0 1152 0 -1 43848
box -48 -56 432 834
use sg13g2_buf_1  input23
timestamp 1676381911
transform 1 0 1152 0 1 43848
box -48 -56 432 834
use sg13g2_buf_1  input24
timestamp 1676381911
transform 1 0 1152 0 -1 45360
box -48 -56 432 834
use sg13g2_buf_1  input25
timestamp 1676381911
transform 1 0 1152 0 -1 18144
box -48 -56 432 834
use sg13g2_buf_1  input26
timestamp 1676381911
transform 1 0 1152 0 -1 46872
box -48 -56 432 834
use sg13g2_buf_1  input27
timestamp 1676381911
transform 1 0 1152 0 1 45360
box -48 -56 432 834
use sg13g2_buf_1  input28
timestamp 1676381911
transform 1 0 1152 0 -1 19656
box -48 -56 432 834
use sg13g2_buf_1  input29
timestamp 1676381911
transform 1 0 1152 0 1 19656
box -48 -56 432 834
use sg13g2_buf_1  input30
timestamp 1676381911
transform 1 0 1152 0 -1 21168
box -48 -56 432 834
use sg13g2_buf_1  input31
timestamp 1676381911
transform 1 0 1152 0 -1 22680
box -48 -56 432 834
use sg13g2_buf_1  input32
timestamp 1676381911
transform 1 0 1152 0 1 22680
box -48 -56 432 834
use sg13g2_buf_1  input33
timestamp 1676381911
transform 1 0 1152 0 -1 24192
box -48 -56 432 834
use sg13g2_buf_1  input34
timestamp 1676381911
transform 1 0 1536 0 -1 25704
box -48 -56 432 834
use sg13g2_buf_1  input35
timestamp 1676381911
transform -1 0 12576 0 -1 3024
box -48 -56 432 834
use sg13g2_buf_1  input36
timestamp 1676381911
transform -1 0 12192 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  input37
timestamp 1676381911
transform -1 0 11808 0 -1 4536
box -48 -56 432 834
use sg13g2_buf_1  input38
timestamp 1676381911
transform -1 0 12576 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  input39
timestamp 1676381911
transform -1 0 12192 0 1 6048
box -48 -56 432 834
use sg13g2_buf_1  input40
timestamp 1676381911
transform -1 0 11808 0 -1 7560
box -48 -56 432 834
use sg13g2_buf_1  input41
timestamp 1676381911
transform -1 0 12576 0 1 6048
box -48 -56 432 834
use sg13g2_buf_1  input42
timestamp 1676381911
transform -1 0 11424 0 1 7560
box -48 -56 432 834
use sg13g2_buf_1  input43
timestamp 1676381911
transform -1 0 12192 0 -1 7560
box -48 -56 432 834
use sg13g2_buf_1  input44
timestamp 1676381911
transform -1 0 10656 0 -1 9072
box -48 -56 432 834
use sg13g2_buf_1  input45
timestamp 1676381911
transform -1 0 11040 0 -1 9072
box -48 -56 432 834
use sg13g2_buf_1  input46
timestamp 1676381911
transform -1 0 11808 0 1 7560
box -48 -56 432 834
use sg13g2_buf_1  input47
timestamp 1676381911
transform -1 0 12192 0 -1 4536
box -48 -56 432 834
use sg13g2_buf_1  input48
timestamp 1676381911
transform -1 0 12576 0 -1 4536
box -48 -56 432 834
use sg13g2_buf_1  input49
timestamp 1676381911
transform -1 0 12192 0 1 4536
box -48 -56 432 834
use sg13g2_buf_1  input50
timestamp 1676381911
transform -1 0 12576 0 1 4536
box -48 -56 432 834
use sg13g2_buf_1  input51
timestamp 1676381911
transform -1 0 12192 0 -1 6048
box -48 -56 432 834
use sg13g2_buf_1  input52
timestamp 1676381911
transform -1 0 11808 0 1 6048
box -48 -56 432 834
use sg13g2_buf_1  input53
timestamp 1676381911
transform -1 0 12576 0 -1 6048
box -48 -56 432 834
use sg13g2_buf_1  input54
timestamp 1676381911
transform -1 0 11424 0 -1 7560
box -48 -56 432 834
use sg13g2_buf_1  input55
timestamp 1676381911
transform -1 0 10464 0 -1 13608
box -48 -56 432 834
use sg13g2_buf_1  input56
timestamp 1676381911
transform -1 0 12576 0 -1 15120
box -48 -56 432 834
use sg13g2_buf_1  input57
timestamp 1676381911
transform -1 0 9600 0 -1 18144
box -48 -56 432 834
use sg13g2_buf_1  input58
timestamp 1676381911
transform -1 0 12192 0 -1 12096
box -48 -56 432 834
use sg13g2_buf_1  input59
timestamp 1676381911
transform -1 0 9408 0 -1 15120
box -48 -56 432 834
use sg13g2_buf_1  input60
timestamp 1676381911
transform -1 0 10176 0 1 13608
box -48 -56 432 834
use sg13g2_buf_1  input61
timestamp 1676381911
transform -1 0 12576 0 -1 12096
box -48 -56 432 834
use sg13g2_buf_1  input62
timestamp 1676381911
transform -1 0 12192 0 1 12096
box -48 -56 432 834
use sg13g2_buf_1  input63
timestamp 1676381911
transform -1 0 12576 0 1 12096
box -48 -56 432 834
use sg13g2_buf_1  input64
timestamp 1676381911
transform -1 0 12576 0 -1 13608
box -48 -56 432 834
use sg13g2_buf_1  input65
timestamp 1676381911
transform -1 0 12576 0 1 13608
box -48 -56 432 834
use sg13g2_buf_1  input66
timestamp 1676381911
transform -1 0 12192 0 -1 15120
box -48 -56 432 834
use sg13g2_buf_1  input67
timestamp 1676381911
transform -1 0 12576 0 -1 7560
box -48 -56 432 834
use sg13g2_buf_1  input68
timestamp 1676381911
transform -1 0 12576 0 -1 10584
box -48 -56 432 834
use sg13g2_buf_1  input69
timestamp 1676381911
transform -1 0 12192 0 1 10584
box -48 -56 432 834
use sg13g2_buf_1  input70
timestamp 1676381911
transform -1 0 9024 0 1 13608
box -48 -56 432 834
use sg13g2_buf_1  input71
timestamp 1676381911
transform -1 0 9408 0 1 13608
box -48 -56 432 834
use sg13g2_buf_1  input72
timestamp 1676381911
transform -1 0 11808 0 -1 12096
box -48 -56 432 834
use sg13g2_buf_1  input73
timestamp 1676381911
transform -1 0 12576 0 1 10584
box -48 -56 432 834
use sg13g2_buf_1  input74
timestamp 1676381911
transform -1 0 11424 0 -1 9072
box -48 -56 432 834
use sg13g2_buf_1  input75
timestamp 1676381911
transform -1 0 12192 0 1 7560
box -48 -56 432 834
use sg13g2_buf_1  input76
timestamp 1676381911
transform -1 0 11808 0 -1 9072
box -48 -56 432 834
use sg13g2_buf_1  input77
timestamp 1676381911
transform -1 0 12576 0 1 7560
box -48 -56 432 834
use sg13g2_buf_1  input78
timestamp 1676381911
transform -1 0 12192 0 -1 9072
box -48 -56 432 834
use sg13g2_buf_1  input79
timestamp 1676381911
transform -1 0 12576 0 -1 9072
box -48 -56 432 834
use sg13g2_buf_1  input80
timestamp 1676381911
transform -1 0 9216 0 1 12096
box -48 -56 432 834
use sg13g2_buf_1  input81
timestamp 1676381911
transform -1 0 12576 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  input82
timestamp 1676381911
transform -1 0 12192 0 -1 10584
box -48 -56 432 834
use sg13g2_buf_1  output83
timestamp 1676381911
transform -1 0 1536 0 -1 3024
box -48 -56 432 834
use sg13g2_buf_1  output84
timestamp 1676381911
transform -1 0 1536 0 -1 4536
box -48 -56 432 834
use sg13g2_buf_1  output85
timestamp 1676381911
transform -1 0 1536 0 1 7560
box -48 -56 432 834
use sg13g2_buf_1  output86
timestamp 1676381911
transform -1 0 1536 0 -1 9072
box -48 -56 432 834
use sg13g2_buf_1  output87
timestamp 1676381911
transform -1 0 1536 0 -1 10584
box -48 -56 432 834
use sg13g2_buf_1  output88
timestamp 1676381911
transform -1 0 1536 0 1 10584
box -48 -56 432 834
use sg13g2_buf_1  output89
timestamp 1676381911
transform -1 0 1536 0 -1 6048
box -48 -56 432 834
use sg13g2_buf_1  output90
timestamp 1676381911
transform -1 0 1536 0 -1 7560
box -48 -56 432 834
use sg13g2_buf_1  output91
timestamp 1676381911
transform -1 0 1536 0 -1 12096
box -48 -56 432 834
use sg13g2_buf_1  output92
timestamp 1676381911
transform -1 0 1536 0 -1 13608
box -48 -56 432 834
use sg13g2_buf_1  output93
timestamp 1676381911
transform -1 0 1536 0 1 13608
box -48 -56 432 834
use sg13g2_buf_1  output94
timestamp 1676381911
transform -1 0 1536 0 -1 15120
box -48 -56 432 834
use sg13g2_buf_1  output95
timestamp 1676381911
transform 1 0 12192 0 -1 16632
box -48 -56 432 834
use sg13g2_buf_1  output96
timestamp 1676381911
transform 1 0 9888 0 -1 19656
box -48 -56 432 834
use sg13g2_buf_1  output97
timestamp 1676381911
transform 1 0 12192 0 1 16632
box -48 -56 432 834
use sg13g2_buf_1  output98
timestamp 1676381911
transform 1 0 9504 0 1 19656
box -48 -56 432 834
use sg13g2_buf_1  output99
timestamp 1676381911
transform 1 0 10272 0 -1 19656
box -48 -56 432 834
use sg13g2_buf_1  output100
timestamp 1676381911
transform 1 0 11808 0 1 18144
box -48 -56 432 834
use sg13g2_buf_1  output101
timestamp 1676381911
transform 1 0 8832 0 1 21168
box -48 -56 432 834
use sg13g2_buf_1  output102
timestamp 1676381911
transform 1 0 12192 0 1 18144
box -48 -56 432 834
use sg13g2_buf_1  output103
timestamp 1676381911
transform 1 0 9216 0 1 21168
box -48 -56 432 834
use sg13g2_buf_1  output104
timestamp 1676381911
transform 1 0 9600 0 1 21168
box -48 -56 432 834
use sg13g2_buf_1  output105
timestamp 1676381911
transform 1 0 9216 0 -1 22680
box -48 -56 432 834
use sg13g2_buf_1  output106
timestamp 1676381911
transform 1 0 9600 0 -1 22680
box -48 -56 432 834
use sg13g2_buf_1  output107
timestamp 1676381911
transform 1 0 10368 0 1 21168
box -48 -56 432 834
use sg13g2_buf_1  output108
timestamp 1676381911
transform 1 0 9984 0 -1 22680
box -48 -56 432 834
use sg13g2_buf_1  output109
timestamp 1676381911
transform 1 0 11808 0 -1 21168
box -48 -56 432 834
use sg13g2_buf_1  output110
timestamp 1676381911
transform 1 0 10368 0 -1 22680
box -48 -56 432 834
use sg13g2_buf_1  output111
timestamp 1676381911
transform 1 0 12192 0 -1 21168
box -48 -56 432 834
use sg13g2_buf_1  output112
timestamp 1676381911
transform 1 0 10368 0 -1 24192
box -48 -56 432 834
use sg13g2_buf_1  output113
timestamp 1676381911
transform 1 0 11424 0 -1 25704
box -48 -56 432 834
use sg13g2_buf_1  output114
timestamp 1676381911
transform 1 0 11808 0 -1 25704
box -48 -56 432 834
use sg13g2_buf_1  output115
timestamp 1676381911
transform 1 0 11808 0 1 33264
box -48 -56 432 834
use sg13g2_buf_1  output116
timestamp 1676381911
transform 1 0 11808 0 1 37800
box -48 -56 432 834
use sg13g2_buf_1  output117
timestamp 1676381911
transform 1 0 12192 0 -1 39312
box -48 -56 432 834
use sg13g2_buf_1  output118
timestamp 1676381911
transform 1 0 12192 0 -1 34776
box -48 -56 432 834
use sg13g2_buf_1  output119
timestamp 1676381911
transform 1 0 11808 0 -1 34776
box -48 -56 432 834
use sg13g2_buf_1  output120
timestamp 1676381911
transform 1 0 12192 0 -1 36288
box -48 -56 432 834
use sg13g2_buf_1  output121
timestamp 1676381911
transform 1 0 12192 0 1 36288
box -48 -56 432 834
use sg13g2_buf_1  output122
timestamp 1676381911
transform 1 0 7488 0 -1 33264
box -48 -56 432 834
use sg13g2_buf_1  output123
timestamp 1676381911
transform 1 0 12192 0 -1 37800
box -48 -56 432 834
use sg13g2_buf_1  output124
timestamp 1676381911
transform 1 0 11808 0 -1 37800
box -48 -56 432 834
use sg13g2_buf_1  output125
timestamp 1676381911
transform 1 0 12192 0 1 37800
box -48 -56 432 834
use sg13g2_buf_1  output126
timestamp 1676381911
transform 1 0 11424 0 -1 37800
box -48 -56 432 834
use sg13g2_buf_1  output127
timestamp 1676381911
transform 1 0 12192 0 1 25704
box -48 -56 432 834
use sg13g2_buf_1  output128
timestamp 1676381911
transform 1 0 11424 0 -1 31752
box -48 -56 432 834
use sg13g2_buf_1  output129
timestamp 1676381911
transform 1 0 9696 0 -1 30240
box -48 -56 432 834
use sg13g2_buf_1  output130
timestamp 1676381911
transform 1 0 9312 0 -1 30240
box -48 -56 432 834
use sg13g2_buf_1  output131
timestamp 1676381911
transform 1 0 12192 0 -1 33264
box -48 -56 432 834
use sg13g2_buf_1  output132
timestamp 1676381911
transform 1 0 11808 0 -1 33264
box -48 -56 432 834
use sg13g2_buf_1  output133
timestamp 1676381911
transform 1 0 12192 0 1 33264
box -48 -56 432 834
use sg13g2_buf_1  output134
timestamp 1676381911
transform 1 0 12192 0 -1 25704
box -48 -56 432 834
use sg13g2_buf_1  output135
timestamp 1676381911
transform 1 0 12192 0 1 24192
box -48 -56 432 834
use sg13g2_buf_1  output136
timestamp 1676381911
transform 1 0 12192 0 1 28728
box -48 -56 432 834
use sg13g2_buf_1  output137
timestamp 1676381911
transform 1 0 11808 0 1 28728
box -48 -56 432 834
use sg13g2_buf_1  output138
timestamp 1676381911
transform 1 0 12192 0 1 30240
box -48 -56 432 834
use sg13g2_buf_1  output139
timestamp 1676381911
transform 1 0 11808 0 1 30240
box -48 -56 432 834
use sg13g2_buf_1  output140
timestamp 1676381911
transform 1 0 12192 0 -1 31752
box -48 -56 432 834
use sg13g2_buf_1  output141
timestamp 1676381911
transform 1 0 11808 0 -1 31752
box -48 -56 432 834
use sg13g2_buf_1  output142
timestamp 1676381911
transform 1 0 10944 0 1 30240
box -48 -56 432 834
use sg13g2_buf_1  output143
timestamp 1676381911
transform 1 0 11424 0 1 37800
box -48 -56 432 834
use sg13g2_buf_1  output144
timestamp 1676381911
transform 1 0 11424 0 1 39312
box -48 -56 432 834
use sg13g2_buf_1  output145
timestamp 1676381911
transform 1 0 10656 0 -1 39312
box -48 -56 432 834
use sg13g2_buf_1  output146
timestamp 1676381911
transform 1 0 11808 0 -1 40824
box -48 -56 432 834
use sg13g2_buf_1  output147
timestamp 1676381911
transform 1 0 11040 0 1 39312
box -48 -56 432 834
use sg13g2_buf_1  output148
timestamp 1676381911
transform 1 0 12192 0 1 40824
box -48 -56 432 834
use sg13g2_buf_1  output149
timestamp 1676381911
transform 1 0 11424 0 -1 40824
box -48 -56 432 834
use sg13g2_buf_1  output150
timestamp 1676381911
transform 1 0 11808 0 1 40824
box -48 -56 432 834
use sg13g2_buf_1  output151
timestamp 1676381911
transform 1 0 12192 0 -1 42336
box -48 -56 432 834
use sg13g2_buf_1  output152
timestamp 1676381911
transform 1 0 11424 0 1 40824
box -48 -56 432 834
use sg13g2_buf_1  output153
timestamp 1676381911
transform 1 0 11808 0 -1 42336
box -48 -56 432 834
use sg13g2_buf_1  output154
timestamp 1676381911
transform 1 0 9120 0 -1 36288
box -48 -56 432 834
use sg13g2_buf_1  output155
timestamp 1676381911
transform 1 0 12192 0 1 42336
box -48 -56 432 834
use sg13g2_buf_1  output156
timestamp 1676381911
transform 1 0 12192 0 -1 43848
box -48 -56 432 834
use sg13g2_buf_1  output157
timestamp 1676381911
transform 1 0 11808 0 -1 43848
box -48 -56 432 834
use sg13g2_buf_1  output158
timestamp 1676381911
transform 1 0 12192 0 1 43848
box -48 -56 432 834
use sg13g2_buf_1  output159
timestamp 1676381911
transform 1 0 11424 0 -1 43848
box -48 -56 432 834
use sg13g2_buf_1  output160
timestamp 1676381911
transform 1 0 11040 0 -1 43848
box -48 -56 432 834
use sg13g2_buf_1  output161
timestamp 1676381911
transform 1 0 12192 0 1 45360
box -48 -56 432 834
use sg13g2_buf_1  output162
timestamp 1676381911
transform 1 0 11808 0 1 45360
box -48 -56 432 834
use sg13g2_buf_1  output163
timestamp 1676381911
transform 1 0 12192 0 -1 46872
box -48 -56 432 834
use sg13g2_buf_1  output164
timestamp 1676381911
transform 1 0 10272 0 -1 45360
box -48 -56 432 834
use sg13g2_buf_1  output165
timestamp 1676381911
transform 1 0 9792 0 1 36288
box -48 -56 432 834
use sg13g2_buf_1  output166
timestamp 1676381911
transform 1 0 11808 0 -1 46872
box -48 -56 432 834
use sg13g2_buf_1  output167
timestamp 1676381911
transform 1 0 10848 0 1 45360
box -48 -56 432 834
use sg13g2_buf_1  output168
timestamp 1676381911
transform 1 0 9408 0 1 36288
box -48 -56 432 834
use sg13g2_buf_1  output169
timestamp 1676381911
transform 1 0 11808 0 -1 39312
box -48 -56 432 834
use sg13g2_buf_1  output170
timestamp 1676381911
transform 1 0 12192 0 1 39312
box -48 -56 432 834
use sg13g2_buf_1  output171
timestamp 1676381911
transform 1 0 11424 0 -1 39312
box -48 -56 432 834
use sg13g2_buf_1  output172
timestamp 1676381911
transform 1 0 11808 0 1 39312
box -48 -56 432 834
use sg13g2_buf_1  output173
timestamp 1676381911
transform 1 0 11040 0 -1 39312
box -48 -56 432 834
use sg13g2_buf_1  output174
timestamp 1676381911
transform 1 0 12192 0 -1 40824
box -48 -56 432 834
use sg13g2_buf_1  output175
timestamp 1676381911
transform -1 0 2016 0 -1 46872
box -48 -56 432 834
use sg13g2_buf_1  output176
timestamp 1676381911
transform -1 0 7776 0 -1 46872
box -48 -56 432 834
use sg13g2_buf_1  output177
timestamp 1676381911
transform -1 0 8352 0 -1 46872
box -48 -56 432 834
use sg13g2_buf_1  output178
timestamp 1676381911
transform -1 0 8928 0 -1 46872
box -48 -56 432 834
use sg13g2_buf_1  output179
timestamp 1676381911
transform -1 0 9504 0 -1 46872
box -48 -56 432 834
use sg13g2_buf_1  output180
timestamp 1676381911
transform -1 0 10080 0 -1 46872
box -48 -56 432 834
use sg13g2_buf_1  output181
timestamp 1676381911
transform -1 0 10656 0 -1 46872
box -48 -56 432 834
use sg13g2_buf_1  output182
timestamp 1676381911
transform -1 0 11232 0 -1 46872
box -48 -56 432 834
use sg13g2_buf_1  output183
timestamp 1676381911
transform -1 0 11808 0 -1 46872
box -48 -56 432 834
use sg13g2_buf_1  output184
timestamp 1676381911
transform 1 0 10464 0 1 45360
box -48 -56 432 834
use sg13g2_buf_1  output185
timestamp 1676381911
transform 1 0 10080 0 1 45360
box -48 -56 432 834
use sg13g2_buf_1  output186
timestamp 1676381911
transform -1 0 2592 0 -1 46872
box -48 -56 432 834
use sg13g2_buf_1  output187
timestamp 1676381911
transform -1 0 3168 0 -1 46872
box -48 -56 432 834
use sg13g2_buf_1  output188
timestamp 1676381911
transform -1 0 3744 0 -1 46872
box -48 -56 432 834
use sg13g2_buf_1  output189
timestamp 1676381911
transform -1 0 4320 0 -1 46872
box -48 -56 432 834
use sg13g2_buf_1  output190
timestamp 1676381911
transform -1 0 4896 0 -1 46872
box -48 -56 432 834
use sg13g2_buf_1  output191
timestamp 1676381911
transform -1 0 5472 0 -1 46872
box -48 -56 432 834
use sg13g2_buf_1  output192
timestamp 1676381911
transform -1 0 6048 0 -1 46872
box -48 -56 432 834
use sg13g2_buf_1  output193
timestamp 1676381911
transform -1 0 6624 0 -1 46872
box -48 -56 432 834
use sg13g2_buf_1  output194
timestamp 1676381911
transform -1 0 7200 0 -1 46872
box -48 -56 432 834
use sg13g2_buf_1  output195
timestamp 1676381911
transform -1 0 1920 0 1 45360
box -48 -56 432 834
<< labels >>
flabel metal2 s 0 2396 90 2476 0 FreeSans 320 0 0 0 A_I_top
port 0 nsew signal output
flabel metal2 s 0 1388 90 1468 0 FreeSans 320 0 0 0 A_O_top
port 1 nsew signal input
flabel metal2 s 0 3404 90 3484 0 FreeSans 320 0 0 0 A_T_top
port 2 nsew signal output
flabel metal2 s 0 7436 90 7516 0 FreeSans 320 0 0 0 A_config_C_bit0
port 3 nsew signal output
flabel metal2 s 0 8444 90 8524 0 FreeSans 320 0 0 0 A_config_C_bit1
port 4 nsew signal output
flabel metal2 s 0 9452 90 9532 0 FreeSans 320 0 0 0 A_config_C_bit2
port 5 nsew signal output
flabel metal2 s 0 10460 90 10540 0 FreeSans 320 0 0 0 A_config_C_bit3
port 6 nsew signal output
flabel metal2 s 0 5420 90 5500 0 FreeSans 320 0 0 0 B_I_top
port 7 nsew signal output
flabel metal2 s 0 4412 90 4492 0 FreeSans 320 0 0 0 B_O_top
port 8 nsew signal input
flabel metal2 s 0 6428 90 6508 0 FreeSans 320 0 0 0 B_T_top
port 9 nsew signal output
flabel metal2 s 0 11468 90 11548 0 FreeSans 320 0 0 0 B_config_C_bit0
port 10 nsew signal output
flabel metal2 s 0 12476 90 12556 0 FreeSans 320 0 0 0 B_config_C_bit1
port 11 nsew signal output
flabel metal2 s 0 13484 90 13564 0 FreeSans 320 0 0 0 B_config_C_bit2
port 12 nsew signal output
flabel metal2 s 0 14492 90 14572 0 FreeSans 320 0 0 0 B_config_C_bit3
port 13 nsew signal output
flabel metal2 s 13638 18860 13728 18940 0 FreeSans 320 0 0 0 E1BEG[0]
port 14 nsew signal output
flabel metal2 s 13638 19196 13728 19276 0 FreeSans 320 0 0 0 E1BEG[1]
port 15 nsew signal output
flabel metal2 s 13638 19532 13728 19612 0 FreeSans 320 0 0 0 E1BEG[2]
port 16 nsew signal output
flabel metal2 s 13638 19868 13728 19948 0 FreeSans 320 0 0 0 E1BEG[3]
port 17 nsew signal output
flabel metal2 s 13638 20204 13728 20284 0 FreeSans 320 0 0 0 E2BEG[0]
port 18 nsew signal output
flabel metal2 s 13638 20540 13728 20620 0 FreeSans 320 0 0 0 E2BEG[1]
port 19 nsew signal output
flabel metal2 s 13638 20876 13728 20956 0 FreeSans 320 0 0 0 E2BEG[2]
port 20 nsew signal output
flabel metal2 s 13638 21212 13728 21292 0 FreeSans 320 0 0 0 E2BEG[3]
port 21 nsew signal output
flabel metal2 s 13638 21548 13728 21628 0 FreeSans 320 0 0 0 E2BEG[4]
port 22 nsew signal output
flabel metal2 s 13638 21884 13728 21964 0 FreeSans 320 0 0 0 E2BEG[5]
port 23 nsew signal output
flabel metal2 s 13638 22220 13728 22300 0 FreeSans 320 0 0 0 E2BEG[6]
port 24 nsew signal output
flabel metal2 s 13638 22556 13728 22636 0 FreeSans 320 0 0 0 E2BEG[7]
port 25 nsew signal output
flabel metal2 s 13638 22892 13728 22972 0 FreeSans 320 0 0 0 E2BEGb[0]
port 26 nsew signal output
flabel metal2 s 13638 23228 13728 23308 0 FreeSans 320 0 0 0 E2BEGb[1]
port 27 nsew signal output
flabel metal2 s 13638 23564 13728 23644 0 FreeSans 320 0 0 0 E2BEGb[2]
port 28 nsew signal output
flabel metal2 s 13638 23900 13728 23980 0 FreeSans 320 0 0 0 E2BEGb[3]
port 29 nsew signal output
flabel metal2 s 13638 24236 13728 24316 0 FreeSans 320 0 0 0 E2BEGb[4]
port 30 nsew signal output
flabel metal2 s 13638 24572 13728 24652 0 FreeSans 320 0 0 0 E2BEGb[5]
port 31 nsew signal output
flabel metal2 s 13638 24908 13728 24988 0 FreeSans 320 0 0 0 E2BEGb[6]
port 32 nsew signal output
flabel metal2 s 13638 25244 13728 25324 0 FreeSans 320 0 0 0 E2BEGb[7]
port 33 nsew signal output
flabel metal2 s 13638 30956 13728 31036 0 FreeSans 320 0 0 0 E6BEG[0]
port 34 nsew signal output
flabel metal2 s 13638 34316 13728 34396 0 FreeSans 320 0 0 0 E6BEG[10]
port 35 nsew signal output
flabel metal2 s 13638 34652 13728 34732 0 FreeSans 320 0 0 0 E6BEG[11]
port 36 nsew signal output
flabel metal2 s 13638 31292 13728 31372 0 FreeSans 320 0 0 0 E6BEG[1]
port 37 nsew signal output
flabel metal2 s 13638 31628 13728 31708 0 FreeSans 320 0 0 0 E6BEG[2]
port 38 nsew signal output
flabel metal2 s 13638 31964 13728 32044 0 FreeSans 320 0 0 0 E6BEG[3]
port 39 nsew signal output
flabel metal2 s 13638 32300 13728 32380 0 FreeSans 320 0 0 0 E6BEG[4]
port 40 nsew signal output
flabel metal2 s 13638 32636 13728 32716 0 FreeSans 320 0 0 0 E6BEG[5]
port 41 nsew signal output
flabel metal2 s 13638 32972 13728 33052 0 FreeSans 320 0 0 0 E6BEG[6]
port 42 nsew signal output
flabel metal2 s 13638 33308 13728 33388 0 FreeSans 320 0 0 0 E6BEG[7]
port 43 nsew signal output
flabel metal2 s 13638 33644 13728 33724 0 FreeSans 320 0 0 0 E6BEG[8]
port 44 nsew signal output
flabel metal2 s 13638 33980 13728 34060 0 FreeSans 320 0 0 0 E6BEG[9]
port 45 nsew signal output
flabel metal2 s 13638 25580 13728 25660 0 FreeSans 320 0 0 0 EE4BEG[0]
port 46 nsew signal output
flabel metal2 s 13638 28940 13728 29020 0 FreeSans 320 0 0 0 EE4BEG[10]
port 47 nsew signal output
flabel metal2 s 13638 29276 13728 29356 0 FreeSans 320 0 0 0 EE4BEG[11]
port 48 nsew signal output
flabel metal2 s 13638 29612 13728 29692 0 FreeSans 320 0 0 0 EE4BEG[12]
port 49 nsew signal output
flabel metal2 s 13638 29948 13728 30028 0 FreeSans 320 0 0 0 EE4BEG[13]
port 50 nsew signal output
flabel metal2 s 13638 30284 13728 30364 0 FreeSans 320 0 0 0 EE4BEG[14]
port 51 nsew signal output
flabel metal2 s 13638 30620 13728 30700 0 FreeSans 320 0 0 0 EE4BEG[15]
port 52 nsew signal output
flabel metal2 s 13638 25916 13728 25996 0 FreeSans 320 0 0 0 EE4BEG[1]
port 53 nsew signal output
flabel metal2 s 13638 26252 13728 26332 0 FreeSans 320 0 0 0 EE4BEG[2]
port 54 nsew signal output
flabel metal2 s 13638 26588 13728 26668 0 FreeSans 320 0 0 0 EE4BEG[3]
port 55 nsew signal output
flabel metal2 s 13638 26924 13728 27004 0 FreeSans 320 0 0 0 EE4BEG[4]
port 56 nsew signal output
flabel metal2 s 13638 27260 13728 27340 0 FreeSans 320 0 0 0 EE4BEG[5]
port 57 nsew signal output
flabel metal2 s 13638 27596 13728 27676 0 FreeSans 320 0 0 0 EE4BEG[6]
port 58 nsew signal output
flabel metal2 s 13638 27932 13728 28012 0 FreeSans 320 0 0 0 EE4BEG[7]
port 59 nsew signal output
flabel metal2 s 13638 28268 13728 28348 0 FreeSans 320 0 0 0 EE4BEG[8]
port 60 nsew signal output
flabel metal2 s 13638 28604 13728 28684 0 FreeSans 320 0 0 0 EE4BEG[9]
port 61 nsew signal output
flabel metal2 s 0 15500 90 15580 0 FreeSans 320 0 0 0 FrameData[0]
port 62 nsew signal input
flabel metal2 s 0 25580 90 25660 0 FreeSans 320 0 0 0 FrameData[10]
port 63 nsew signal input
flabel metal2 s 0 26588 90 26668 0 FreeSans 320 0 0 0 FrameData[11]
port 64 nsew signal input
flabel metal2 s 0 27596 90 27676 0 FreeSans 320 0 0 0 FrameData[12]
port 65 nsew signal input
flabel metal2 s 0 28604 90 28684 0 FreeSans 320 0 0 0 FrameData[13]
port 66 nsew signal input
flabel metal2 s 0 29612 90 29692 0 FreeSans 320 0 0 0 FrameData[14]
port 67 nsew signal input
flabel metal2 s 0 30620 90 30700 0 FreeSans 320 0 0 0 FrameData[15]
port 68 nsew signal input
flabel metal2 s 0 31628 90 31708 0 FreeSans 320 0 0 0 FrameData[16]
port 69 nsew signal input
flabel metal2 s 0 32636 90 32716 0 FreeSans 320 0 0 0 FrameData[17]
port 70 nsew signal input
flabel metal2 s 0 33644 90 33724 0 FreeSans 320 0 0 0 FrameData[18]
port 71 nsew signal input
flabel metal2 s 0 34652 90 34732 0 FreeSans 320 0 0 0 FrameData[19]
port 72 nsew signal input
flabel metal2 s 0 16508 90 16588 0 FreeSans 320 0 0 0 FrameData[1]
port 73 nsew signal input
flabel metal2 s 0 35660 90 35740 0 FreeSans 320 0 0 0 FrameData[20]
port 74 nsew signal input
flabel metal2 s 0 36668 90 36748 0 FreeSans 320 0 0 0 FrameData[21]
port 75 nsew signal input
flabel metal2 s 0 37676 90 37756 0 FreeSans 320 0 0 0 FrameData[22]
port 76 nsew signal input
flabel metal2 s 0 38684 90 38764 0 FreeSans 320 0 0 0 FrameData[23]
port 77 nsew signal input
flabel metal2 s 0 39692 90 39772 0 FreeSans 320 0 0 0 FrameData[24]
port 78 nsew signal input
flabel metal2 s 0 40700 90 40780 0 FreeSans 320 0 0 0 FrameData[25]
port 79 nsew signal input
flabel metal2 s 0 41708 90 41788 0 FreeSans 320 0 0 0 FrameData[26]
port 80 nsew signal input
flabel metal2 s 0 42716 90 42796 0 FreeSans 320 0 0 0 FrameData[27]
port 81 nsew signal input
flabel metal2 s 0 43724 90 43804 0 FreeSans 320 0 0 0 FrameData[28]
port 82 nsew signal input
flabel metal2 s 0 44732 90 44812 0 FreeSans 320 0 0 0 FrameData[29]
port 83 nsew signal input
flabel metal2 s 0 17516 90 17596 0 FreeSans 320 0 0 0 FrameData[2]
port 84 nsew signal input
flabel metal2 s 0 45740 90 45820 0 FreeSans 320 0 0 0 FrameData[30]
port 85 nsew signal input
flabel metal2 s 0 46748 90 46828 0 FreeSans 320 0 0 0 FrameData[31]
port 86 nsew signal input
flabel metal2 s 0 18524 90 18604 0 FreeSans 320 0 0 0 FrameData[3]
port 87 nsew signal input
flabel metal2 s 0 19532 90 19612 0 FreeSans 320 0 0 0 FrameData[4]
port 88 nsew signal input
flabel metal2 s 0 20540 90 20620 0 FreeSans 320 0 0 0 FrameData[5]
port 89 nsew signal input
flabel metal2 s 0 21548 90 21628 0 FreeSans 320 0 0 0 FrameData[6]
port 90 nsew signal input
flabel metal2 s 0 22556 90 22636 0 FreeSans 320 0 0 0 FrameData[7]
port 91 nsew signal input
flabel metal2 s 0 23564 90 23644 0 FreeSans 320 0 0 0 FrameData[8]
port 92 nsew signal input
flabel metal2 s 0 24572 90 24652 0 FreeSans 320 0 0 0 FrameData[9]
port 93 nsew signal input
flabel metal2 s 13638 34988 13728 35068 0 FreeSans 320 0 0 0 FrameData_O[0]
port 94 nsew signal output
flabel metal2 s 13638 38348 13728 38428 0 FreeSans 320 0 0 0 FrameData_O[10]
port 95 nsew signal output
flabel metal2 s 13638 38684 13728 38764 0 FreeSans 320 0 0 0 FrameData_O[11]
port 96 nsew signal output
flabel metal2 s 13638 39020 13728 39100 0 FreeSans 320 0 0 0 FrameData_O[12]
port 97 nsew signal output
flabel metal2 s 13638 39356 13728 39436 0 FreeSans 320 0 0 0 FrameData_O[13]
port 98 nsew signal output
flabel metal2 s 13638 39692 13728 39772 0 FreeSans 320 0 0 0 FrameData_O[14]
port 99 nsew signal output
flabel metal2 s 13638 40028 13728 40108 0 FreeSans 320 0 0 0 FrameData_O[15]
port 100 nsew signal output
flabel metal2 s 13638 40364 13728 40444 0 FreeSans 320 0 0 0 FrameData_O[16]
port 101 nsew signal output
flabel metal2 s 13638 40700 13728 40780 0 FreeSans 320 0 0 0 FrameData_O[17]
port 102 nsew signal output
flabel metal2 s 13638 41036 13728 41116 0 FreeSans 320 0 0 0 FrameData_O[18]
port 103 nsew signal output
flabel metal2 s 13638 41372 13728 41452 0 FreeSans 320 0 0 0 FrameData_O[19]
port 104 nsew signal output
flabel metal2 s 13638 35324 13728 35404 0 FreeSans 320 0 0 0 FrameData_O[1]
port 105 nsew signal output
flabel metal2 s 13638 41708 13728 41788 0 FreeSans 320 0 0 0 FrameData_O[20]
port 106 nsew signal output
flabel metal2 s 13638 42044 13728 42124 0 FreeSans 320 0 0 0 FrameData_O[21]
port 107 nsew signal output
flabel metal2 s 13638 42380 13728 42460 0 FreeSans 320 0 0 0 FrameData_O[22]
port 108 nsew signal output
flabel metal2 s 13638 42716 13728 42796 0 FreeSans 320 0 0 0 FrameData_O[23]
port 109 nsew signal output
flabel metal2 s 13638 43052 13728 43132 0 FreeSans 320 0 0 0 FrameData_O[24]
port 110 nsew signal output
flabel metal2 s 13638 43388 13728 43468 0 FreeSans 320 0 0 0 FrameData_O[25]
port 111 nsew signal output
flabel metal2 s 13638 43724 13728 43804 0 FreeSans 320 0 0 0 FrameData_O[26]
port 112 nsew signal output
flabel metal2 s 13638 44060 13728 44140 0 FreeSans 320 0 0 0 FrameData_O[27]
port 113 nsew signal output
flabel metal2 s 13638 44396 13728 44476 0 FreeSans 320 0 0 0 FrameData_O[28]
port 114 nsew signal output
flabel metal2 s 13638 44732 13728 44812 0 FreeSans 320 0 0 0 FrameData_O[29]
port 115 nsew signal output
flabel metal2 s 13638 35660 13728 35740 0 FreeSans 320 0 0 0 FrameData_O[2]
port 116 nsew signal output
flabel metal2 s 13638 45068 13728 45148 0 FreeSans 320 0 0 0 FrameData_O[30]
port 117 nsew signal output
flabel metal2 s 13638 45404 13728 45484 0 FreeSans 320 0 0 0 FrameData_O[31]
port 118 nsew signal output
flabel metal2 s 13638 35996 13728 36076 0 FreeSans 320 0 0 0 FrameData_O[3]
port 119 nsew signal output
flabel metal2 s 13638 36332 13728 36412 0 FreeSans 320 0 0 0 FrameData_O[4]
port 120 nsew signal output
flabel metal2 s 13638 36668 13728 36748 0 FreeSans 320 0 0 0 FrameData_O[5]
port 121 nsew signal output
flabel metal2 s 13638 37004 13728 37084 0 FreeSans 320 0 0 0 FrameData_O[6]
port 122 nsew signal output
flabel metal2 s 13638 37340 13728 37420 0 FreeSans 320 0 0 0 FrameData_O[7]
port 123 nsew signal output
flabel metal2 s 13638 37676 13728 37756 0 FreeSans 320 0 0 0 FrameData_O[8]
port 124 nsew signal output
flabel metal2 s 13638 38012 13728 38092 0 FreeSans 320 0 0 0 FrameData_O[9]
port 125 nsew signal output
flabel metal3 s 1592 0 1672 80 0 FreeSans 320 0 0 0 FrameStrobe[0]
port 126 nsew signal input
flabel metal3 s 7352 0 7432 80 0 FreeSans 320 0 0 0 FrameStrobe[10]
port 127 nsew signal input
flabel metal3 s 7928 0 8008 80 0 FreeSans 320 0 0 0 FrameStrobe[11]
port 128 nsew signal input
flabel metal3 s 8504 0 8584 80 0 FreeSans 320 0 0 0 FrameStrobe[12]
port 129 nsew signal input
flabel metal3 s 9080 0 9160 80 0 FreeSans 320 0 0 0 FrameStrobe[13]
port 130 nsew signal input
flabel metal3 s 9656 0 9736 80 0 FreeSans 320 0 0 0 FrameStrobe[14]
port 131 nsew signal input
flabel metal3 s 10232 0 10312 80 0 FreeSans 320 0 0 0 FrameStrobe[15]
port 132 nsew signal input
flabel metal3 s 10808 0 10888 80 0 FreeSans 320 0 0 0 FrameStrobe[16]
port 133 nsew signal input
flabel metal3 s 11384 0 11464 80 0 FreeSans 320 0 0 0 FrameStrobe[17]
port 134 nsew signal input
flabel metal3 s 11960 0 12040 80 0 FreeSans 320 0 0 0 FrameStrobe[18]
port 135 nsew signal input
flabel metal3 s 12536 0 12616 80 0 FreeSans 320 0 0 0 FrameStrobe[19]
port 136 nsew signal input
flabel metal3 s 2168 0 2248 80 0 FreeSans 320 0 0 0 FrameStrobe[1]
port 137 nsew signal input
flabel metal3 s 2744 0 2824 80 0 FreeSans 320 0 0 0 FrameStrobe[2]
port 138 nsew signal input
flabel metal3 s 3320 0 3400 80 0 FreeSans 320 0 0 0 FrameStrobe[3]
port 139 nsew signal input
flabel metal3 s 3896 0 3976 80 0 FreeSans 320 0 0 0 FrameStrobe[4]
port 140 nsew signal input
flabel metal3 s 4472 0 4552 80 0 FreeSans 320 0 0 0 FrameStrobe[5]
port 141 nsew signal input
flabel metal3 s 5048 0 5128 80 0 FreeSans 320 0 0 0 FrameStrobe[6]
port 142 nsew signal input
flabel metal3 s 5624 0 5704 80 0 FreeSans 320 0 0 0 FrameStrobe[7]
port 143 nsew signal input
flabel metal3 s 6200 0 6280 80 0 FreeSans 320 0 0 0 FrameStrobe[8]
port 144 nsew signal input
flabel metal3 s 6776 0 6856 80 0 FreeSans 320 0 0 0 FrameStrobe[9]
port 145 nsew signal input
flabel metal3 s 1592 48304 1672 48384 0 FreeSans 320 0 0 0 FrameStrobe_O[0]
port 146 nsew signal output
flabel metal3 s 7352 48304 7432 48384 0 FreeSans 320 0 0 0 FrameStrobe_O[10]
port 147 nsew signal output
flabel metal3 s 7928 48304 8008 48384 0 FreeSans 320 0 0 0 FrameStrobe_O[11]
port 148 nsew signal output
flabel metal3 s 8504 48304 8584 48384 0 FreeSans 320 0 0 0 FrameStrobe_O[12]
port 149 nsew signal output
flabel metal3 s 9080 48304 9160 48384 0 FreeSans 320 0 0 0 FrameStrobe_O[13]
port 150 nsew signal output
flabel metal3 s 9656 48304 9736 48384 0 FreeSans 320 0 0 0 FrameStrobe_O[14]
port 151 nsew signal output
flabel metal3 s 10232 48304 10312 48384 0 FreeSans 320 0 0 0 FrameStrobe_O[15]
port 152 nsew signal output
flabel metal3 s 10808 48304 10888 48384 0 FreeSans 320 0 0 0 FrameStrobe_O[16]
port 153 nsew signal output
flabel metal3 s 11384 48304 11464 48384 0 FreeSans 320 0 0 0 FrameStrobe_O[17]
port 154 nsew signal output
flabel metal3 s 11960 48304 12040 48384 0 FreeSans 320 0 0 0 FrameStrobe_O[18]
port 155 nsew signal output
flabel metal3 s 12536 48304 12616 48384 0 FreeSans 320 0 0 0 FrameStrobe_O[19]
port 156 nsew signal output
flabel metal3 s 2168 48304 2248 48384 0 FreeSans 320 0 0 0 FrameStrobe_O[1]
port 157 nsew signal output
flabel metal3 s 2744 48304 2824 48384 0 FreeSans 320 0 0 0 FrameStrobe_O[2]
port 158 nsew signal output
flabel metal3 s 3320 48304 3400 48384 0 FreeSans 320 0 0 0 FrameStrobe_O[3]
port 159 nsew signal output
flabel metal3 s 3896 48304 3976 48384 0 FreeSans 320 0 0 0 FrameStrobe_O[4]
port 160 nsew signal output
flabel metal3 s 4472 48304 4552 48384 0 FreeSans 320 0 0 0 FrameStrobe_O[5]
port 161 nsew signal output
flabel metal3 s 5048 48304 5128 48384 0 FreeSans 320 0 0 0 FrameStrobe_O[6]
port 162 nsew signal output
flabel metal3 s 5624 48304 5704 48384 0 FreeSans 320 0 0 0 FrameStrobe_O[7]
port 163 nsew signal output
flabel metal3 s 6200 48304 6280 48384 0 FreeSans 320 0 0 0 FrameStrobe_O[8]
port 164 nsew signal output
flabel metal3 s 6776 48304 6856 48384 0 FreeSans 320 0 0 0 FrameStrobe_O[9]
port 165 nsew signal output
flabel metal3 s 1016 0 1096 80 0 FreeSans 320 0 0 0 UserCLK
port 166 nsew signal input
flabel metal3 s 1016 48304 1096 48384 0 FreeSans 320 0 0 0 UserCLKo
port 167 nsew signal output
flabel metal5 s 4892 0 5332 48384 0 FreeSans 2560 90 0 0 VGND
port 168 nsew ground bidirectional
flabel metal5 s 4892 0 5332 40 0 FreeSans 320 0 0 0 VGND
port 168 nsew ground bidirectional
flabel metal5 s 4892 48344 5332 48384 0 FreeSans 320 0 0 0 VGND
port 168 nsew ground bidirectional
flabel metal5 s 3652 0 4092 48384 0 FreeSans 2560 90 0 0 VPWR
port 169 nsew power bidirectional
flabel metal5 s 3652 0 4092 40 0 FreeSans 320 0 0 0 VPWR
port 169 nsew power bidirectional
flabel metal5 s 3652 48344 4092 48384 0 FreeSans 320 0 0 0 VPWR
port 169 nsew power bidirectional
flabel metal2 s 13638 2732 13728 2812 0 FreeSans 320 0 0 0 W1END[0]
port 170 nsew signal input
flabel metal2 s 13638 3068 13728 3148 0 FreeSans 320 0 0 0 W1END[1]
port 171 nsew signal input
flabel metal2 s 13638 3404 13728 3484 0 FreeSans 320 0 0 0 W1END[2]
port 172 nsew signal input
flabel metal2 s 13638 3740 13728 3820 0 FreeSans 320 0 0 0 W1END[3]
port 173 nsew signal input
flabel metal2 s 13638 6764 13728 6844 0 FreeSans 320 0 0 0 W2END[0]
port 174 nsew signal input
flabel metal2 s 13638 7100 13728 7180 0 FreeSans 320 0 0 0 W2END[1]
port 175 nsew signal input
flabel metal2 s 13638 7436 13728 7516 0 FreeSans 320 0 0 0 W2END[2]
port 176 nsew signal input
flabel metal2 s 13638 7772 13728 7852 0 FreeSans 320 0 0 0 W2END[3]
port 177 nsew signal input
flabel metal2 s 13638 8108 13728 8188 0 FreeSans 320 0 0 0 W2END[4]
port 178 nsew signal input
flabel metal2 s 13638 8444 13728 8524 0 FreeSans 320 0 0 0 W2END[5]
port 179 nsew signal input
flabel metal2 s 13638 8780 13728 8860 0 FreeSans 320 0 0 0 W2END[6]
port 180 nsew signal input
flabel metal2 s 13638 9116 13728 9196 0 FreeSans 320 0 0 0 W2END[7]
port 181 nsew signal input
flabel metal2 s 13638 4076 13728 4156 0 FreeSans 320 0 0 0 W2MID[0]
port 182 nsew signal input
flabel metal2 s 13638 4412 13728 4492 0 FreeSans 320 0 0 0 W2MID[1]
port 183 nsew signal input
flabel metal2 s 13638 4748 13728 4828 0 FreeSans 320 0 0 0 W2MID[2]
port 184 nsew signal input
flabel metal2 s 13638 5084 13728 5164 0 FreeSans 320 0 0 0 W2MID[3]
port 185 nsew signal input
flabel metal2 s 13638 5420 13728 5500 0 FreeSans 320 0 0 0 W2MID[4]
port 186 nsew signal input
flabel metal2 s 13638 5756 13728 5836 0 FreeSans 320 0 0 0 W2MID[5]
port 187 nsew signal input
flabel metal2 s 13638 6092 13728 6172 0 FreeSans 320 0 0 0 W2MID[6]
port 188 nsew signal input
flabel metal2 s 13638 6428 13728 6508 0 FreeSans 320 0 0 0 W2MID[7]
port 189 nsew signal input
flabel metal2 s 13638 14828 13728 14908 0 FreeSans 320 0 0 0 W6END[0]
port 190 nsew signal input
flabel metal2 s 13638 18188 13728 18268 0 FreeSans 320 0 0 0 W6END[10]
port 191 nsew signal input
flabel metal2 s 13638 18524 13728 18604 0 FreeSans 320 0 0 0 W6END[11]
port 192 nsew signal input
flabel metal2 s 13638 15164 13728 15244 0 FreeSans 320 0 0 0 W6END[1]
port 193 nsew signal input
flabel metal2 s 13638 15500 13728 15580 0 FreeSans 320 0 0 0 W6END[2]
port 194 nsew signal input
flabel metal2 s 13638 15836 13728 15916 0 FreeSans 320 0 0 0 W6END[3]
port 195 nsew signal input
flabel metal2 s 13638 16172 13728 16252 0 FreeSans 320 0 0 0 W6END[4]
port 196 nsew signal input
flabel metal2 s 13638 16508 13728 16588 0 FreeSans 320 0 0 0 W6END[5]
port 197 nsew signal input
flabel metal2 s 13638 16844 13728 16924 0 FreeSans 320 0 0 0 W6END[6]
port 198 nsew signal input
flabel metal2 s 13638 17180 13728 17260 0 FreeSans 320 0 0 0 W6END[7]
port 199 nsew signal input
flabel metal2 s 13638 17516 13728 17596 0 FreeSans 320 0 0 0 W6END[8]
port 200 nsew signal input
flabel metal2 s 13638 17852 13728 17932 0 FreeSans 320 0 0 0 W6END[9]
port 201 nsew signal input
flabel metal2 s 13638 9452 13728 9532 0 FreeSans 320 0 0 0 WW4END[0]
port 202 nsew signal input
flabel metal2 s 13638 12812 13728 12892 0 FreeSans 320 0 0 0 WW4END[10]
port 203 nsew signal input
flabel metal2 s 13638 13148 13728 13228 0 FreeSans 320 0 0 0 WW4END[11]
port 204 nsew signal input
flabel metal2 s 13638 13484 13728 13564 0 FreeSans 320 0 0 0 WW4END[12]
port 205 nsew signal input
flabel metal2 s 13638 13820 13728 13900 0 FreeSans 320 0 0 0 WW4END[13]
port 206 nsew signal input
flabel metal2 s 13638 14156 13728 14236 0 FreeSans 320 0 0 0 WW4END[14]
port 207 nsew signal input
flabel metal2 s 13638 14492 13728 14572 0 FreeSans 320 0 0 0 WW4END[15]
port 208 nsew signal input
flabel metal2 s 13638 9788 13728 9868 0 FreeSans 320 0 0 0 WW4END[1]
port 209 nsew signal input
flabel metal2 s 13638 10124 13728 10204 0 FreeSans 320 0 0 0 WW4END[2]
port 210 nsew signal input
flabel metal2 s 13638 10460 13728 10540 0 FreeSans 320 0 0 0 WW4END[3]
port 211 nsew signal input
flabel metal2 s 13638 10796 13728 10876 0 FreeSans 320 0 0 0 WW4END[4]
port 212 nsew signal input
flabel metal2 s 13638 11132 13728 11212 0 FreeSans 320 0 0 0 WW4END[5]
port 213 nsew signal input
flabel metal2 s 13638 11468 13728 11548 0 FreeSans 320 0 0 0 WW4END[6]
port 214 nsew signal input
flabel metal2 s 13638 11804 13728 11884 0 FreeSans 320 0 0 0 WW4END[7]
port 215 nsew signal input
flabel metal2 s 13638 12140 13728 12220 0 FreeSans 320 0 0 0 WW4END[8]
port 216 nsew signal input
flabel metal2 s 13638 12476 13728 12556 0 FreeSans 320 0 0 0 WW4END[9]
port 217 nsew signal input
rlabel metal1 6864 46872 6864 46872 0 VGND
rlabel metal1 6864 46116 6864 46116 0 VPWR
rlabel metal2 632 2436 632 2436 0 A_I_top
rlabel via2 80 1428 80 1428 0 A_O_top
rlabel via2 80 3444 80 3444 0 A_T_top
rlabel metal2 632 7476 632 7476 0 A_config_C_bit0
rlabel metal2 632 8484 632 8484 0 A_config_C_bit1
rlabel via2 80 9492 80 9492 0 A_config_C_bit2
rlabel metal2 632 10500 632 10500 0 A_config_C_bit3
rlabel metal2 632 5460 632 5460 0 B_I_top
rlabel metal2 656 4452 656 4452 0 B_O_top
rlabel metal2 320 6468 320 6468 0 B_T_top
rlabel metal2 632 11508 632 11508 0 B_config_C_bit0
rlabel metal2 622 13020 622 13020 0 B_config_C_bit1
rlabel via2 80 13524 80 13524 0 B_config_C_bit2
rlabel metal2 632 14532 632 14532 0 B_config_C_bit3
rlabel metal2 12648 16464 12648 16464 0 E1BEG[0]
rlabel metal2 13263 19236 13263 19236 0 E1BEG[1]
rlabel metal2 12696 17220 12696 17220 0 E1BEG[2]
rlabel metal2 10320 20118 10320 20118 0 E1BEG[3]
rlabel metal2 11112 19488 11112 19488 0 E2BEG[0]
rlabel metal2 12168 18564 12168 18564 0 E2BEG[1]
rlabel metal2 9456 21210 9456 21210 0 E2BEG[2]
rlabel metal2 12552 18648 12552 18648 0 E2BEG[3]
rlabel metal2 9552 21294 9552 21294 0 E2BEG[4]
rlabel metal2 10440 21420 10440 21420 0 E2BEG[5]
rlabel metal2 12639 22260 12639 22260 0 E2BEG[6]
rlabel metal2 10080 22512 10080 22512 0 E2BEG[7]
rlabel metal2 10824 21588 10824 21588 0 E2BEGb[0]
rlabel metal2 10392 22512 10392 22512 0 E2BEGb[1]
rlabel metal2 12168 21000 12168 21000 0 E2BEGb[2]
rlabel metal2 11112 22512 11112 22512 0 E2BEGb[3]
rlabel metal2 12696 21000 12696 21000 0 E2BEGb[4]
rlabel metal2 11592 24024 11592 24024 0 E2BEGb[5]
rlabel metal2 13023 24948 13023 24948 0 E2BEGb[6]
rlabel metal2 13311 25284 13311 25284 0 E2BEGb[7]
rlabel metal2 12216 33432 12216 33432 0 E6BEG[0]
rlabel metal2 13167 34356 13167 34356 0 E6BEG[10]
rlabel metal2 13359 34692 13359 34692 0 E6BEG[11]
rlabel metal2 12888 34188 12888 34188 0 E6BEG[1]
rlabel metal2 12456 34272 12456 34272 0 E6BEG[2]
rlabel metal4 12576 34104 12576 34104 0 E6BEG[3]
rlabel metal2 12936 36456 12936 36456 0 E6BEG[4]
rlabel metal2 13167 32676 13167 32676 0 E6BEG[5]
rlabel metal2 13080 37212 13080 37212 0 E6BEG[6]
rlabel metal2 13551 33348 13551 33348 0 E6BEG[7]
rlabel metal2 13263 33684 13263 33684 0 E6BEG[8]
rlabel metal2 12831 34020 12831 34020 0 E6BEG[9]
rlabel metal2 13095 25620 13095 25620 0 EE4BEG[0]
rlabel metal2 12831 28980 12831 28980 0 EE4BEG[10]
rlabel metal2 11919 29316 11919 29316 0 EE4BEG[11]
rlabel metal2 10272 29694 10272 29694 0 EE4BEG[12]
rlabel metal2 13119 29988 13119 29988 0 EE4BEG[13]
rlabel metal2 12975 30324 12975 30324 0 EE4BEG[14]
rlabel metal2 12792 33432 12792 33432 0 EE4BEG[15]
rlabel metal2 12840 25536 12840 25536 0 EE4BEG[1]
rlabel metal2 12792 24780 12792 24780 0 EE4BEG[2]
rlabel metal2 13407 26628 13407 26628 0 EE4BEG[3]
rlabel metal2 13023 26964 13023 26964 0 EE4BEG[4]
rlabel metal2 13359 27300 13359 27300 0 EE4BEG[5]
rlabel metal2 13215 27636 13215 27636 0 EE4BEG[6]
rlabel metal2 13455 27972 13455 27972 0 EE4BEG[7]
rlabel metal2 13503 28308 13503 28308 0 EE4BEG[8]
rlabel metal2 12783 28644 12783 28644 0 EE4BEG[9]
rlabel metal2 656 15540 656 15540 0 FrameData[0]
rlabel metal2 80 25620 80 25620 0 FrameData[10]
rlabel metal2 656 26628 656 26628 0 FrameData[11]
rlabel metal2 656 27636 656 27636 0 FrameData[12]
rlabel via2 80 28644 80 28644 0 FrameData[13]
rlabel via2 80 29652 80 29652 0 FrameData[14]
rlabel metal2 656 30660 656 30660 0 FrameData[15]
rlabel via2 80 31668 80 31668 0 FrameData[16]
rlabel via2 80 32676 80 32676 0 FrameData[17]
rlabel metal2 656 33684 656 33684 0 FrameData[18]
rlabel via2 80 34692 80 34692 0 FrameData[19]
rlabel via2 80 16548 80 16548 0 FrameData[1]
rlabel via2 80 35700 80 35700 0 FrameData[20]
rlabel metal2 656 36708 656 36708 0 FrameData[21]
rlabel via2 80 37716 80 37716 0 FrameData[22]
rlabel via2 80 38724 80 38724 0 FrameData[23]
rlabel metal2 656 39732 656 39732 0 FrameData[24]
rlabel via2 80 40740 80 40740 0 FrameData[25]
rlabel via2 80 41748 80 41748 0 FrameData[26]
rlabel metal2 656 42756 656 42756 0 FrameData[27]
rlabel via2 80 43764 80 43764 0 FrameData[28]
rlabel via2 80 44772 80 44772 0 FrameData[29]
rlabel via2 80 17556 80 17556 0 FrameData[2]
rlabel metal2 368 45780 368 45780 0 FrameData[30]
rlabel metal2 656 46788 656 46788 0 FrameData[31]
rlabel via2 80 18564 80 18564 0 FrameData[3]
rlabel via2 80 19572 80 19572 0 FrameData[4]
rlabel via2 80 20580 80 20580 0 FrameData[5]
rlabel metal2 656 21588 656 21588 0 FrameData[6]
rlabel metal2 646 23100 646 23100 0 FrameData[7]
rlabel metal2 656 23604 656 23604 0 FrameData[8]
rlabel metal2 80 24612 80 24612 0 FrameData[9]
rlabel metal2 13023 35028 13023 35028 0 FrameData_O[0]
rlabel metal2 12831 38388 12831 38388 0 FrameData_O[10]
rlabel via2 13647 38724 13647 38724 0 FrameData_O[11]
rlabel metal2 13647 39060 13647 39060 0 FrameData_O[12]
rlabel metal2 12519 39396 12519 39396 0 FrameData_O[13]
rlabel metal2 13407 39732 13407 39732 0 FrameData_O[14]
rlabel metal2 12711 40068 12711 40068 0 FrameData_O[15]
rlabel metal2 13263 40404 13263 40404 0 FrameData_O[16]
rlabel metal2 13311 40740 13311 40740 0 FrameData_O[17]
rlabel metal2 12711 41076 12711 41076 0 FrameData_O[18]
rlabel via2 13647 41412 13647 41412 0 FrameData_O[19]
rlabel metal2 13119 35364 13119 35364 0 FrameData_O[1]
rlabel metal2 13407 41748 13407 41748 0 FrameData_O[20]
rlabel metal2 13359 42084 13359 42084 0 FrameData_O[21]
rlabel metal2 13023 42420 13023 42420 0 FrameData_O[22]
rlabel metal2 13407 42756 13407 42756 0 FrameData_O[23]
rlabel metal2 12711 43092 12711 43092 0 FrameData_O[24]
rlabel metal2 13599 43428 13599 43428 0 FrameData_O[25]
rlabel metal2 13359 43764 13359 43764 0 FrameData_O[26]
rlabel metal2 12975 44100 12975 44100 0 FrameData_O[27]
rlabel metal2 13407 44436 13407 44436 0 FrameData_O[28]
rlabel metal2 12927 44772 12927 44772 0 FrameData_O[29]
rlabel metal2 13215 35700 13215 35700 0 FrameData_O[2]
rlabel metal2 13023 45108 13023 45108 0 FrameData_O[30]
rlabel metal2 12831 45444 12831 45444 0 FrameData_O[31]
rlabel metal2 13599 36036 13599 36036 0 FrameData_O[3]
rlabel metal2 13311 36372 13311 36372 0 FrameData_O[4]
rlabel metal2 13407 36708 13407 36708 0 FrameData_O[5]
rlabel metal2 12735 37044 12735 37044 0 FrameData_O[6]
rlabel metal2 13503 37380 13503 37380 0 FrameData_O[7]
rlabel metal2 12879 37716 12879 37716 0 FrameData_O[8]
rlabel metal2 13551 38052 13551 38052 0 FrameData_O[9]
rlabel metal3 1632 1626 1632 1626 0 FrameStrobe[0]
rlabel metal3 7392 156 7392 156 0 FrameStrobe[10]
rlabel metal3 7968 1470 7968 1470 0 FrameStrobe[11]
rlabel metal4 8928 7560 8928 7560 0 FrameStrobe[12]
rlabel metal3 9120 534 9120 534 0 FrameStrobe[13]
rlabel metal3 9696 534 9696 534 0 FrameStrobe[14]
rlabel metal3 10272 534 10272 534 0 FrameStrobe[15]
rlabel metal3 10848 534 10848 534 0 FrameStrobe[16]
rlabel metal3 11424 534 11424 534 0 FrameStrobe[17]
rlabel metal3 12000 366 12000 366 0 FrameStrobe[18]
rlabel metal4 11232 41916 11232 41916 0 FrameStrobe[19]
rlabel metal3 2208 744 2208 744 0 FrameStrobe[1]
rlabel metal3 2784 744 2784 744 0 FrameStrobe[2]
rlabel metal2 3840 11592 3840 11592 0 FrameStrobe[3]
rlabel via3 3936 72 3936 72 0 FrameStrobe[4]
rlabel metal3 4512 492 4512 492 0 FrameStrobe[5]
rlabel metal3 5088 114 5088 114 0 FrameStrobe[6]
rlabel metal3 5664 744 5664 744 0 FrameStrobe[7]
rlabel metal3 6240 744 6240 744 0 FrameStrobe[8]
rlabel metal3 6816 660 6816 660 0 FrameStrobe[9]
rlabel metal2 1656 46704 1656 46704 0 FrameStrobe_O[0]
rlabel metal2 7416 46704 7416 46704 0 FrameStrobe_O[10]
rlabel metal2 7992 46704 7992 46704 0 FrameStrobe_O[11]
rlabel metal2 8568 46704 8568 46704 0 FrameStrobe_O[12]
rlabel metal2 9144 46704 9144 46704 0 FrameStrobe_O[13]
rlabel metal2 9720 46704 9720 46704 0 FrameStrobe_O[14]
rlabel metal2 10296 46704 10296 46704 0 FrameStrobe_O[15]
rlabel metal2 10872 46704 10872 46704 0 FrameStrobe_O[16]
rlabel metal2 11448 46704 11448 46704 0 FrameStrobe_O[17]
rlabel metal2 11400 45864 11400 45864 0 FrameStrobe_O[18]
rlabel metal2 10728 45948 10728 45948 0 FrameStrobe_O[19]
rlabel metal2 2232 46704 2232 46704 0 FrameStrobe_O[1]
rlabel metal2 2808 46704 2808 46704 0 FrameStrobe_O[2]
rlabel metal2 3384 46704 3384 46704 0 FrameStrobe_O[3]
rlabel metal2 3960 46704 3960 46704 0 FrameStrobe_O[4]
rlabel metal2 4536 46704 4536 46704 0 FrameStrobe_O[5]
rlabel metal2 5256 46704 5256 46704 0 FrameStrobe_O[6]
rlabel metal2 5688 46704 5688 46704 0 FrameStrobe_O[7]
rlabel metal2 6264 46704 6264 46704 0 FrameStrobe_O[8]
rlabel metal2 6840 46704 6840 46704 0 FrameStrobe_O[9]
rlabel metal4 11136 16884 11136 16884 0 Inst_A_IO_1_bidirectional_frame_config_pass.Q
rlabel metal2 11520 20034 11520 20034 0 Inst_B_IO_1_bidirectional_frame_config_pass.Q
rlabel metal2 6672 36120 6672 36120 0 Inst_W_IO_ConfigMem.Inst_frame0_bit0.Q
rlabel metal2 8640 37380 8640 37380 0 Inst_W_IO_ConfigMem.Inst_frame0_bit1.Q
rlabel metal2 9888 29106 9888 29106 0 Inst_W_IO_ConfigMem.Inst_frame0_bit10.Q
rlabel metal2 11240 29064 11240 29064 0 Inst_W_IO_ConfigMem.Inst_frame0_bit11.Q
rlabel metal2 6672 35112 6672 35112 0 Inst_W_IO_ConfigMem.Inst_frame0_bit12.Q
rlabel via2 8648 35112 8648 35112 0 Inst_W_IO_ConfigMem.Inst_frame0_bit13.Q
rlabel metal3 9888 11382 9888 11382 0 Inst_W_IO_ConfigMem.Inst_frame0_bit14.Q
rlabel metal2 11712 13020 11712 13020 0 Inst_W_IO_ConfigMem.Inst_frame0_bit15.Q
rlabel metal2 10320 19992 10320 19992 0 Inst_W_IO_ConfigMem.Inst_frame0_bit16.Q
rlabel metal2 12144 19488 12144 19488 0 Inst_W_IO_ConfigMem.Inst_frame0_bit17.Q
rlabel metal2 2496 15540 2496 15540 0 Inst_W_IO_ConfigMem.Inst_frame0_bit18.Q
rlabel metal2 4224 14826 4224 14826 0 Inst_W_IO_ConfigMem.Inst_frame0_bit19.Q
rlabel metal3 4128 22386 4128 22386 0 Inst_W_IO_ConfigMem.Inst_frame0_bit2.Q
rlabel via2 4611 14784 4611 14784 0 Inst_W_IO_ConfigMem.Inst_frame0_bit20.Q
rlabel metal2 4848 13776 4848 13776 0 Inst_W_IO_ConfigMem.Inst_frame0_bit21.Q
rlabel metal2 5712 6720 5712 6720 0 Inst_W_IO_ConfigMem.Inst_frame0_bit22.Q
rlabel metal2 5400 10962 5400 10962 0 Inst_W_IO_ConfigMem.Inst_frame0_bit23.Q
rlabel metal2 5184 9492 5184 9492 0 Inst_W_IO_ConfigMem.Inst_frame0_bit24.Q
rlabel metal2 4080 16464 4080 16464 0 Inst_W_IO_ConfigMem.Inst_frame0_bit25.Q
rlabel metal3 4608 16254 4608 16254 0 Inst_W_IO_ConfigMem.Inst_frame0_bit26.Q
rlabel metal2 6336 13314 6336 13314 0 Inst_W_IO_ConfigMem.Inst_frame0_bit27.Q
rlabel via1 6151 17808 6151 17808 0 Inst_W_IO_ConfigMem.Inst_frame0_bit28.Q
rlabel metal3 7776 24906 7776 24906 0 Inst_W_IO_ConfigMem.Inst_frame0_bit29.Q
rlabel via2 5768 23016 5768 23016 0 Inst_W_IO_ConfigMem.Inst_frame0_bit3.Q
rlabel metal2 8448 26040 8448 26040 0 Inst_W_IO_ConfigMem.Inst_frame0_bit30.Q
rlabel metal3 8736 25662 8736 25662 0 Inst_W_IO_ConfigMem.Inst_frame0_bit31.Q
rlabel metal2 7248 4284 7248 4284 0 Inst_W_IO_ConfigMem.Inst_frame0_bit4.Q
rlabel metal2 9176 4872 9176 4872 0 Inst_W_IO_ConfigMem.Inst_frame0_bit5.Q
rlabel metal2 11568 11172 11568 11172 0 Inst_W_IO_ConfigMem.Inst_frame0_bit6.Q
rlabel metal2 9648 9576 9648 9576 0 Inst_W_IO_ConfigMem.Inst_frame0_bit7.Q
rlabel metal2 10992 16464 10992 16464 0 Inst_W_IO_ConfigMem.Inst_frame0_bit8.Q
rlabel metal3 12096 16758 12096 16758 0 Inst_W_IO_ConfigMem.Inst_frame0_bit9.Q
rlabel metal2 5952 34944 5952 34944 0 Inst_W_IO_ConfigMem.Inst_frame1_bit0.Q
rlabel metal2 4704 33012 4704 33012 0 Inst_W_IO_ConfigMem.Inst_frame1_bit1.Q
rlabel metal2 11136 33432 11136 33432 0 Inst_W_IO_ConfigMem.Inst_frame1_bit10.Q
rlabel metal2 9600 32928 9600 32928 0 Inst_W_IO_ConfigMem.Inst_frame1_bit11.Q
rlabel metal2 5472 37212 5472 37212 0 Inst_W_IO_ConfigMem.Inst_frame1_bit12.Q
rlabel metal2 4608 31458 4608 31458 0 Inst_W_IO_ConfigMem.Inst_frame1_bit13.Q
rlabel metal3 12096 25410 12096 25410 0 Inst_W_IO_ConfigMem.Inst_frame1_bit14.Q
rlabel metal2 9984 25998 9984 25998 0 Inst_W_IO_ConfigMem.Inst_frame1_bit15.Q
rlabel metal3 10176 36120 10176 36120 0 Inst_W_IO_ConfigMem.Inst_frame1_bit16.Q
rlabel metal2 12432 35364 12432 35364 0 Inst_W_IO_ConfigMem.Inst_frame1_bit17.Q
rlabel metal2 5136 29316 5136 29316 0 Inst_W_IO_ConfigMem.Inst_frame1_bit18.Q
rlabel metal2 4080 28560 4080 28560 0 Inst_W_IO_ConfigMem.Inst_frame1_bit19.Q
rlabel metal2 3936 20916 3936 20916 0 Inst_W_IO_ConfigMem.Inst_frame1_bit2.Q
rlabel metal2 5969 32004 5969 32004 0 Inst_W_IO_ConfigMem.Inst_frame1_bit20.Q
rlabel metal3 4320 31836 4320 31836 0 Inst_W_IO_ConfigMem.Inst_frame1_bit21.Q
rlabel metal2 6624 5544 6624 5544 0 Inst_W_IO_ConfigMem.Inst_frame1_bit22.Q
rlabel metal2 5184 9660 5184 9660 0 Inst_W_IO_ConfigMem.Inst_frame1_bit23.Q
rlabel metal2 8168 18480 8168 18480 0 Inst_W_IO_ConfigMem.Inst_frame1_bit24.Q
rlabel metal2 6096 18480 6096 18480 0 Inst_W_IO_ConfigMem.Inst_frame1_bit25.Q
rlabel metal2 4416 26922 4416 26922 0 Inst_W_IO_ConfigMem.Inst_frame1_bit26.Q
rlabel metal3 5952 27132 5952 27132 0 Inst_W_IO_ConfigMem.Inst_frame1_bit27.Q
rlabel metal2 8016 5712 8016 5712 0 Inst_W_IO_ConfigMem.Inst_frame1_bit28.Q
rlabel metal3 9600 5964 9600 5964 0 Inst_W_IO_ConfigMem.Inst_frame1_bit29.Q
rlabel metal2 6912 21000 6912 21000 0 Inst_W_IO_ConfigMem.Inst_frame1_bit3.Q
rlabel metal2 7680 23856 7680 23856 0 Inst_W_IO_ConfigMem.Inst_frame1_bit30.Q
rlabel metal2 9840 23856 9840 23856 0 Inst_W_IO_ConfigMem.Inst_frame1_bit31.Q
rlabel metal3 5568 6426 5568 6426 0 Inst_W_IO_ConfigMem.Inst_frame1_bit4.Q
rlabel metal2 7728 5544 7728 5544 0 Inst_W_IO_ConfigMem.Inst_frame1_bit5.Q
rlabel metal2 8456 12432 8456 12432 0 Inst_W_IO_ConfigMem.Inst_frame1_bit6.Q
rlabel metal2 7536 10332 7536 10332 0 Inst_W_IO_ConfigMem.Inst_frame1_bit7.Q
rlabel metal2 9072 15708 9072 15708 0 Inst_W_IO_ConfigMem.Inst_frame1_bit8.Q
rlabel metal3 9504 15414 9504 15414 0 Inst_W_IO_ConfigMem.Inst_frame1_bit9.Q
rlabel metal2 6384 33600 6384 33600 0 Inst_W_IO_ConfigMem.Inst_frame2_bit0.Q
rlabel metal2 8168 33600 8168 33600 0 Inst_W_IO_ConfigMem.Inst_frame2_bit1.Q
rlabel metal2 7536 23016 7536 23016 0 Inst_W_IO_ConfigMem.Inst_frame2_bit10.Q
rlabel via2 9224 23016 9224 23016 0 Inst_W_IO_ConfigMem.Inst_frame2_bit11.Q
rlabel metal2 5808 38388 5808 38388 0 Inst_W_IO_ConfigMem.Inst_frame2_bit12.Q
rlabel metal2 8256 39018 8256 39018 0 Inst_W_IO_ConfigMem.Inst_frame2_bit13.Q
rlabel metal3 9792 26166 9792 26166 0 Inst_W_IO_ConfigMem.Inst_frame2_bit14.Q
rlabel metal2 11664 26880 11664 26880 0 Inst_W_IO_ConfigMem.Inst_frame2_bit15.Q
rlabel metal2 7872 34482 7872 34482 0 Inst_W_IO_ConfigMem.Inst_frame2_bit16.Q
rlabel metal3 9408 34692 9408 34692 0 Inst_W_IO_ConfigMem.Inst_frame2_bit17.Q
rlabel metal2 4656 19488 4656 19488 0 Inst_W_IO_ConfigMem.Inst_frame2_bit18.Q
rlabel metal3 4128 20538 4128 20538 0 Inst_W_IO_ConfigMem.Inst_frame2_bit19.Q
rlabel metal2 4464 22344 4464 22344 0 Inst_W_IO_ConfigMem.Inst_frame2_bit2.Q
rlabel metal2 5472 4872 5472 4872 0 Inst_W_IO_ConfigMem.Inst_frame2_bit20.Q
rlabel metal2 7016 4872 7016 4872 0 Inst_W_IO_ConfigMem.Inst_frame2_bit21.Q
rlabel metal2 5664 4284 5664 4284 0 Inst_W_IO_ConfigMem.Inst_frame2_bit22.Q
rlabel metal2 4512 9030 4512 9030 0 Inst_W_IO_ConfigMem.Inst_frame2_bit23.Q
rlabel metal2 9216 17976 9216 17976 0 Inst_W_IO_ConfigMem.Inst_frame2_bit24.Q
rlabel metal2 10920 18480 10920 18480 0 Inst_W_IO_ConfigMem.Inst_frame2_bit25.Q
rlabel metal2 10184 27552 10184 27552 0 Inst_W_IO_ConfigMem.Inst_frame2_bit26.Q
rlabel metal2 8544 27552 8544 27552 0 Inst_W_IO_ConfigMem.Inst_frame2_bit27.Q
rlabel metal2 10656 37464 10656 37464 0 Inst_W_IO_ConfigMem.Inst_frame2_bit28.Q
rlabel metal2 9120 37464 9120 37464 0 Inst_W_IO_ConfigMem.Inst_frame2_bit29.Q
rlabel metal2 5952 22344 5952 22344 0 Inst_W_IO_ConfigMem.Inst_frame2_bit3.Q
rlabel metal3 7488 30324 7488 30324 0 Inst_W_IO_ConfigMem.Inst_frame2_bit30.Q
rlabel metal2 5424 30576 5424 30576 0 Inst_W_IO_ConfigMem.Inst_frame2_bit31.Q
rlabel metal2 7344 3612 7344 3612 0 Inst_W_IO_ConfigMem.Inst_frame2_bit4.Q
rlabel metal2 8832 4242 8832 4242 0 Inst_W_IO_ConfigMem.Inst_frame2_bit5.Q
rlabel metal3 8928 9870 8928 9870 0 Inst_W_IO_ConfigMem.Inst_frame2_bit6.Q
rlabel metal3 9792 10290 9792 10290 0 Inst_W_IO_ConfigMem.Inst_frame2_bit7.Q
rlabel metal2 9840 16968 9840 16968 0 Inst_W_IO_ConfigMem.Inst_frame2_bit8.Q
rlabel metal2 12000 14196 12000 14196 0 Inst_W_IO_ConfigMem.Inst_frame2_bit9.Q
rlabel metal3 6720 5754 6720 5754 0 Inst_W_IO_ConfigMem.Inst_frame3_bit22.Q
rlabel metal3 4128 11802 4128 11802 0 Inst_W_IO_ConfigMem.Inst_frame3_bit23.Q
rlabel metal3 9024 7476 9024 7476 0 Inst_W_IO_ConfigMem.Inst_frame3_bit24.Q
rlabel metal2 9360 20244 9360 20244 0 Inst_W_IO_ConfigMem.Inst_frame3_bit25.Q
rlabel metal2 7296 22344 7296 22344 0 Inst_W_IO_ConfigMem.Inst_frame3_bit26.Q
rlabel metal2 8592 21420 8592 21420 0 Inst_W_IO_ConfigMem.Inst_frame3_bit27.Q
rlabel metal2 7200 38178 7200 38178 0 Inst_W_IO_ConfigMem.Inst_frame3_bit28.Q
rlabel metal2 8736 38241 8736 38241 0 Inst_W_IO_ConfigMem.Inst_frame3_bit29.Q
rlabel metal2 8640 28434 8640 28434 0 Inst_W_IO_ConfigMem.Inst_frame3_bit30.Q
rlabel metal3 10176 28644 10176 28644 0 Inst_W_IO_ConfigMem.Inst_frame3_bit31.Q
rlabel metal2 9552 4956 9552 4956 0 Inst_W_IO_switch_matrix.E1BEG0
rlabel metal2 4704 11718 4704 11718 0 Inst_W_IO_switch_matrix.E1BEG1
rlabel metal2 9888 8022 9888 8022 0 Inst_W_IO_switch_matrix.E1BEG2
rlabel metal2 10128 20076 10128 20076 0 Inst_W_IO_switch_matrix.E1BEG3
rlabel metal2 9552 22596 9552 22596 0 Inst_W_IO_switch_matrix.E2BEG0
rlabel metal2 9168 37968 9168 37968 0 Inst_W_IO_switch_matrix.E2BEG1
rlabel metal2 12144 28308 12144 28308 0 Inst_W_IO_switch_matrix.E2BEG2
rlabel metal2 8664 33684 8664 33684 0 Inst_W_IO_switch_matrix.E2BEG3
rlabel metal2 6456 22260 6456 22260 0 Inst_W_IO_switch_matrix.E2BEG4
rlabel metal2 9384 3948 9384 3948 0 Inst_W_IO_switch_matrix.E2BEG5
rlabel metal2 11712 10290 11712 10290 0 Inst_W_IO_switch_matrix.E2BEG6
rlabel metal3 11712 15750 11712 15750 0 Inst_W_IO_switch_matrix.E2BEG7
rlabel metal2 10368 23142 10368 23142 0 Inst_W_IO_switch_matrix.E2BEGb0
rlabel metal2 8568 38892 8568 38892 0 Inst_W_IO_switch_matrix.E2BEGb1
rlabel metal2 11688 26628 11688 26628 0 Inst_W_IO_switch_matrix.E2BEGb2
rlabel metal2 11616 34314 11616 34314 0 Inst_W_IO_switch_matrix.E2BEGb3
rlabel metal2 4272 21588 4272 21588 0 Inst_W_IO_switch_matrix.E2BEGb4
rlabel metal2 7680 2604 7680 2604 0 Inst_W_IO_switch_matrix.E2BEGb5
rlabel metal3 7776 9954 7776 9954 0 Inst_W_IO_switch_matrix.E2BEGb6
rlabel metal2 11808 17052 11808 17052 0 Inst_W_IO_switch_matrix.E2BEGb7
rlabel metal2 6264 26796 6264 26796 0 Inst_W_IO_switch_matrix.E6BEG0
rlabel metal2 9912 5628 9912 5628 0 Inst_W_IO_switch_matrix.E6BEG1
rlabel metal3 11616 10878 11616 10878 0 Inst_W_IO_switch_matrix.E6BEG10
rlabel metal2 11424 18606 11424 18606 0 Inst_W_IO_switch_matrix.E6BEG11
rlabel metal2 9720 23772 9720 23772 0 Inst_W_IO_switch_matrix.E6BEG2
rlabel metal2 8928 38892 8928 38892 0 Inst_W_IO_switch_matrix.E6BEG3
rlabel metal2 6072 23100 6072 23100 0 Inst_W_IO_switch_matrix.E6BEG4
rlabel metal2 10176 4914 10176 4914 0 Inst_W_IO_switch_matrix.E6BEG5
rlabel metal2 9360 12516 9360 12516 0 Inst_W_IO_switch_matrix.E6BEG6
rlabel metal2 11952 17976 11952 17976 0 Inst_W_IO_switch_matrix.E6BEG7
rlabel metal3 11616 29778 11616 29778 0 Inst_W_IO_switch_matrix.E6BEG8
rlabel metal2 8952 35196 8952 35196 0 Inst_W_IO_switch_matrix.E6BEG9
rlabel metal3 11712 27006 11712 27006 0 Inst_W_IO_switch_matrix.EE4BEG0
rlabel metal3 11040 37926 11040 37926 0 Inst_W_IO_switch_matrix.EE4BEG1
rlabel metal2 11832 26292 11832 26292 0 Inst_W_IO_switch_matrix.EE4BEG10
rlabel metal3 11328 36750 11328 36750 0 Inst_W_IO_switch_matrix.EE4BEG11
rlabel metal2 5640 29652 5640 29652 0 Inst_W_IO_switch_matrix.EE4BEG12
rlabel metal2 6144 31962 6144 31962 0 Inst_W_IO_switch_matrix.EE4BEG13
rlabel metal2 7704 11676 7704 11676 0 Inst_W_IO_switch_matrix.EE4BEG14
rlabel metal2 8568 18564 8568 18564 0 Inst_W_IO_switch_matrix.EE4BEG15
rlabel metal2 7416 30660 7416 30660 0 Inst_W_IO_switch_matrix.EE4BEG2
rlabel metal2 6912 32886 6912 32886 0 Inst_W_IO_switch_matrix.EE4BEG3
rlabel metal2 6768 21336 6768 21336 0 Inst_W_IO_switch_matrix.EE4BEG4
rlabel metal3 8352 8568 8352 8568 0 Inst_W_IO_switch_matrix.EE4BEG5
rlabel metal2 9120 13188 9120 13188 0 Inst_W_IO_switch_matrix.EE4BEG6
rlabel metal2 9432 16212 9432 16212 0 Inst_W_IO_switch_matrix.EE4BEG7
rlabel metal3 10176 33432 10176 33432 0 Inst_W_IO_switch_matrix.EE4BEG8
rlabel metal3 6336 31878 6336 31878 0 Inst_W_IO_switch_matrix.EE4BEG9
rlabel metal2 1344 29736 1344 29736 0 UserCLK
rlabel metal2 1320 45948 1320 45948 0 UserCLKo
rlabel metal2 13599 2772 13599 2772 0 W1END[0]
rlabel metal2 13263 3108 13263 3108 0 W1END[1]
rlabel metal2 13167 3444 13167 3444 0 W1END[2]
rlabel metal2 13071 3780 13071 3780 0 W1END[3]
rlabel metal2 12879 6804 12879 6804 0 W2END[0]
rlabel metal2 13215 7140 13215 7140 0 W2END[1]
rlabel metal2 13071 7476 13071 7476 0 W2END[2]
rlabel metal2 12495 7812 12495 7812 0 W2END[3]
rlabel metal2 12879 8148 12879 8148 0 W2END[4]
rlabel metal2 13071 8484 13071 8484 0 W2END[5]
rlabel metal2 12303 8820 12303 8820 0 W2END[6]
rlabel metal2 12687 9156 12687 9156 0 W2END[7]
rlabel metal2 13263 4116 13263 4116 0 W2MID[0]
rlabel metal2 13071 4452 13071 4452 0 W2MID[1]
rlabel metal2 12879 4788 12879 4788 0 W2MID[2]
rlabel metal2 13071 5124 13071 5124 0 W2MID[3]
rlabel metal2 13263 5460 13263 5460 0 W2MID[4]
rlabel metal2 12687 5796 12687 5796 0 W2MID[5]
rlabel metal2 13071 6132 13071 6132 0 W2MID[6]
rlabel metal2 13119 6468 13119 6468 0 W2MID[7]
rlabel metal2 12015 14868 12015 14868 0 W6END[0]
rlabel metal2 13407 18228 13407 18228 0 W6END[10]
rlabel metal2 9504 17934 9504 17934 0 W6END[11]
rlabel metal3 12240 14112 12240 14112 0 W6END[1]
rlabel metal2 9312 14994 9312 14994 0 W6END[2]
rlabel metal2 11871 15876 11871 15876 0 W6END[3]
rlabel metal2 13263 16212 13263 16212 0 W6END[4]
rlabel metal2 13119 16548 13119 16548 0 W6END[5]
rlabel metal2 13311 16884 13311 16884 0 W6END[6]
rlabel metal2 13503 17220 13503 17220 0 W6END[7]
rlabel metal2 13071 17556 13071 17556 0 W6END[8]
rlabel metal2 12975 17892 12975 17892 0 W6END[9]
rlabel metal2 13119 9492 13119 9492 0 WW4END[0]
rlabel metal2 13071 12852 13071 12852 0 WW4END[10]
rlabel metal2 12336 13104 12336 13104 0 WW4END[11]
rlabel metal2 8928 13986 8928 13986 0 WW4END[12]
rlabel metal2 9312 14070 9312 14070 0 WW4END[13]
rlabel metal2 13215 14196 13215 14196 0 WW4END[14]
rlabel metal2 13407 14532 13407 14532 0 WW4END[15]
rlabel metal2 12495 9828 12495 9828 0 WW4END[1]
rlabel metal2 13263 10164 13263 10164 0 WW4END[2]
rlabel metal2 12783 10500 12783 10500 0 WW4END[3]
rlabel metal2 13407 10836 13407 10836 0 WW4END[4]
rlabel metal2 12975 11172 12975 11172 0 WW4END[5]
rlabel metal2 13551 11508 13551 11508 0 WW4END[6]
rlabel metal2 13599 11844 13599 11844 0 WW4END[7]
rlabel metal2 13359 12180 13359 12180 0 WW4END[8]
rlabel metal2 13503 12516 13503 12516 0 WW4END[9]
rlabel metal2 4752 13272 4752 13272 0 _000_
rlabel metal2 5448 8736 5448 8736 0 _001_
rlabel metal2 5712 14616 5712 14616 0 _002_
rlabel metal2 5424 17556 5424 17556 0 _003_
rlabel metal2 4608 14952 4608 14952 0 _004_
rlabel metal2 6597 13272 6597 13272 0 _005_
rlabel metal2 5808 14700 5808 14700 0 _006_
rlabel metal2 7008 17976 7008 17976 0 _007_
rlabel metal3 7488 17388 7488 17388 0 _008_
rlabel metal2 6091 13314 6091 13314 0 _009_
rlabel metal2 6264 13188 6264 13188 0 _010_
rlabel metal2 6432 13482 6432 13482 0 _011_
rlabel metal3 6912 14742 6912 14742 0 _012_
rlabel metal2 7584 16464 7584 16464 0 _013_
rlabel metal2 8304 14868 8304 14868 0 _014_
rlabel metal2 7920 14616 7920 14616 0 _015_
rlabel metal3 7008 15036 7008 15036 0 _016_
rlabel metal2 4065 14742 4065 14742 0 _017_
rlabel metal2 4368 14700 4368 14700 0 _018_
rlabel metal3 4704 14070 4704 14070 0 _019_
rlabel metal2 8277 15456 8277 15456 0 _020_
rlabel metal2 6384 12684 6384 12684 0 _021_
rlabel metal2 6528 12264 6528 12264 0 _022_
rlabel metal2 7776 16758 7776 16758 0 _023_
rlabel metal2 5280 13482 5280 13482 0 _024_
rlabel metal2 5760 13440 5760 13440 0 _025_
rlabel metal2 6384 13776 6384 13776 0 _026_
rlabel metal3 4992 12558 4992 12558 0 _027_
rlabel metal2 7176 13986 7176 13986 0 _028_
rlabel metal3 7296 14448 7296 14448 0 _029_
rlabel metal2 7893 13986 7893 13986 0 _030_
rlabel metal2 8304 13776 8304 13776 0 _031_
rlabel metal3 6144 9912 6144 9912 0 _032_
rlabel metal2 5808 11004 5808 11004 0 _033_
rlabel metal3 5856 9534 5856 9534 0 _034_
rlabel metal3 6912 9702 6912 9702 0 _035_
rlabel metal2 6000 8820 6000 8820 0 _036_
rlabel metal2 5760 7308 5760 7308 0 _037_
rlabel metal2 5712 8736 5712 8736 0 _038_
rlabel metal2 6528 8484 6528 8484 0 _039_
rlabel metal2 8640 25242 8640 25242 0 _040_
rlabel metal2 8904 24780 8904 24780 0 _041_
rlabel metal2 8184 25368 8184 25368 0 _042_
rlabel metal2 8352 25410 8352 25410 0 _043_
rlabel metal2 9216 25452 9216 25452 0 _044_
rlabel metal2 3144 2100 3144 2100 0 net1
rlabel metal2 1488 31878 1488 31878 0 net10
rlabel metal5 7344 18076 7344 18076 0 net100
rlabel metal2 12696 8904 12696 8904 0 net101
rlabel metal2 12216 8484 12216 8484 0 net102
rlabel metal3 8112 18312 8112 18312 0 net103
rlabel metal2 10512 16968 10512 16968 0 net104
rlabel metal2 8928 10920 8928 10920 0 net105
rlabel metal2 2016 2604 2016 2604 0 net106
rlabel metal2 1536 4116 1536 4116 0 net107
rlabel metal4 1488 7980 1488 7980 0 net108
rlabel metal3 1968 16128 1968 16128 0 net109
rlabel metal2 10992 19320 10992 19320 0 net11
rlabel metal4 1824 15960 1824 15960 0 net110
rlabel metal4 1584 11004 1584 11004 0 net111
rlabel metal2 4224 5544 4224 5544 0 net112
rlabel metal5 1440 15876 1440 15876 0 net113
rlabel metal2 2160 24612 2160 24612 0 net114
rlabel metal3 1296 25956 1296 25956 0 net115
rlabel metal2 2688 25116 2688 25116 0 net116
rlabel metal2 2592 14868 2592 14868 0 net117
rlabel metal2 11088 16128 11088 16128 0 net118
rlabel metal3 9168 16464 9168 16464 0 net119
rlabel metal2 2400 19320 2400 19320 0 net12
rlabel metal3 11856 14028 11856 14028 0 net120
rlabel metal2 9768 20076 9768 20076 0 net121
rlabel metal2 10296 23268 10296 23268 0 net122
rlabel metal4 10848 18648 10848 18648 0 net123
rlabel metal2 9216 21504 9216 21504 0 net124
rlabel metal4 9408 22512 9408 22512 0 net125
rlabel metal3 9312 21882 9312 21882 0 net126
rlabel metal3 9072 19320 9072 19320 0 net127
rlabel metal3 9264 17640 9264 17640 0 net128
rlabel metal2 10632 14616 10632 14616 0 net129
rlabel metal2 2592 26040 2592 26040 0 net13
rlabel metal2 10512 21588 10512 21588 0 net130
rlabel metal2 9744 38976 9744 38976 0 net131
rlabel metal2 11880 25956 11880 25956 0 net132
rlabel metal2 11064 34188 11064 34188 0 net133
rlabel metal2 12288 20790 12288 20790 0 net134
rlabel metal2 8232 2856 8232 2856 0 net135
rlabel metal4 9600 17892 9600 17892 0 net136
rlabel metal2 12024 17220 12024 17220 0 net137
rlabel metal2 6792 27048 6792 27048 0 net138
rlabel metal4 11472 38220 11472 38220 0 net139
rlabel metal2 2424 17136 2424 17136 0 net14
rlabel metal2 11688 18312 11688 18312 0 net140
rlabel metal4 11328 34356 11328 34356 0 net141
rlabel metal2 10944 34104 10944 34104 0 net142
rlabel metal2 12288 35826 12288 35826 0 net143
rlabel metal4 6336 34944 6336 34944 0 net144
rlabel metal3 7488 18564 7488 18564 0 net145
rlabel metal4 10512 37212 10512 37212 0 net146
rlabel metal2 11928 16464 11928 16464 0 net147
rlabel metal3 11664 33348 11664 33348 0 net148
rlabel metal2 9288 34944 9288 34944 0 net149
rlabel metal4 2832 17388 2832 17388 0 net15
rlabel metal2 12288 26376 12288 26376 0 net150
rlabel metal2 11784 27048 11784 27048 0 net151
rlabel metal2 10440 37212 10440 37212 0 net152
rlabel metal2 7512 29232 7512 29232 0 net153
rlabel metal2 7608 33012 7608 33012 0 net154
rlabel metal2 8040 11928 8040 11928 0 net155
rlabel metal4 12192 33684 12192 33684 0 net156
rlabel metal2 11208 37968 11208 37968 0 net157
rlabel metal2 12288 24654 12288 24654 0 net158
rlabel metal2 12288 29190 12288 29190 0 net159
rlabel metal2 3120 13944 3120 13944 0 net16
rlabel metal2 9624 22428 9624 22428 0 net160
rlabel metal2 8568 8148 8568 8148 0 net161
rlabel metal2 9768 13440 9768 13440 0 net162
rlabel metal2 9288 16464 9288 16464 0 net163
rlabel metal2 10944 33474 10944 33474 0 net164
rlabel metal2 10992 30660 10992 30660 0 net165
rlabel metal2 5496 35784 5496 35784 0 net166
rlabel metal4 9600 35616 9600 35616 0 net167
rlabel metal3 9936 38892 9936 38892 0 net168
rlabel metal2 5112 39060 5112 39060 0 net169
rlabel metal2 1512 37968 1512 37968 0 net17
rlabel metal2 7992 39144 7992 39144 0 net170
rlabel metal4 11904 18312 11904 18312 0 net171
rlabel metal2 10536 14196 10536 14196 0 net172
rlabel metal2 10680 36876 10680 36876 0 net173
rlabel metal2 9912 35700 9912 35700 0 net174
rlabel metal2 2616 29316 2616 29316 0 net175
rlabel metal3 5856 17976 5856 17976 0 net176
rlabel metal2 6696 35364 6696 35364 0 net177
rlabel metal4 3168 13776 3168 13776 0 net178
rlabel metal2 3432 4284 3432 4284 0 net179
rlabel metal2 2136 38892 2136 38892 0 net18
rlabel metal3 3312 13608 3312 13608 0 net180
rlabel metal4 4944 37968 4944 37968 0 net181
rlabel metal4 9024 40320 9024 40320 0 net182
rlabel metal2 3432 18648 3432 18648 0 net183
rlabel metal4 12912 29232 12912 29232 0 net184
rlabel metal4 12048 39396 12048 39396 0 net185
rlabel metal3 11904 35994 11904 35994 0 net186
rlabel metal2 10656 45024 10656 45024 0 net187
rlabel metal3 2304 27360 2304 27360 0 net188
rlabel metal2 6360 29316 6360 29316 0 net189
rlabel metal2 7344 17808 7344 17808 0 net19
rlabel metal2 10608 45696 10608 45696 0 net190
rlabel metal2 9552 36708 9552 36708 0 net191
rlabel metal2 5592 2436 5592 2436 0 net192
rlabel metal2 10248 2772 10248 2772 0 net193
rlabel metal4 13200 18648 13200 18648 0 net194
rlabel metal4 12240 13860 12240 13860 0 net195
rlabel metal2 9960 17976 9960 17976 0 net196
rlabel metal2 11784 14952 11784 14952 0 net197
rlabel metal5 1920 30156 1920 30156 0 net198
rlabel metal2 8040 43680 8040 43680 0 net199
rlabel metal2 10128 15792 10128 15792 0 net2
rlabel metal3 1920 16758 1920 16758 0 net20
rlabel metal2 10824 44436 10824 44436 0 net200
rlabel metal2 11256 44940 11256 44940 0 net201
rlabel metal2 9960 44436 9960 44436 0 net202
rlabel metal2 11016 45108 11016 45108 0 net203
rlabel metal2 11448 45192 11448 45192 0 net204
rlabel metal2 11208 45948 11208 45948 0 net205
rlabel metal2 11304 42924 11304 42924 0 net206
rlabel metal2 10968 42840 10968 42840 0 net207
rlabel metal2 11736 42924 11736 42924 0 net208
rlabel metal3 2496 41160 2496 41160 0 net209
rlabel metal2 1896 41832 1896 41832 0 net21
rlabel metal2 6888 31584 6888 31584 0 net210
rlabel metal3 4176 17976 4176 17976 0 net211
rlabel metal2 11352 44436 11352 44436 0 net212
rlabel metal2 10632 44352 10632 44352 0 net213
rlabel metal2 10392 45192 10392 45192 0 net214
rlabel metal2 5832 45192 5832 45192 0 net215
rlabel metal2 5592 45108 5592 45108 0 net216
rlabel metal2 8664 45192 8664 45192 0 net217
rlabel metal2 10176 30366 10176 30366 0 net218
rlabel metal3 10848 30492 10848 30492 0 net219
rlabel metal2 6384 16380 6384 16380 0 net22
rlabel metal2 11280 33768 11280 33768 0 net220
rlabel metal4 6336 18228 6336 18228 0 net23
rlabel metal3 2688 41370 2688 41370 0 net24
rlabel metal3 2208 19404 2208 19404 0 net25
rlabel metal4 5088 38304 5088 38304 0 net26
rlabel metal2 8064 29778 8064 29778 0 net27
rlabel metal2 3024 22344 3024 22344 0 net28
rlabel metal2 5280 2604 5280 2604 0 net29
rlabel metal3 4704 17136 4704 17136 0 net3
rlabel metal2 1608 20580 1608 20580 0 net30
rlabel metal2 2184 22092 2184 22092 0 net31
rlabel metal2 1656 23100 1656 23100 0 net32
rlabel metal2 1488 23562 1488 23562 0 net33
rlabel metal2 10848 15498 10848 15498 0 net34
rlabel metal2 12888 2856 12888 2856 0 net35
rlabel metal2 9696 7896 9696 7896 0 net36
rlabel metal4 4368 14364 4368 14364 0 net37
rlabel metal3 7776 4284 7776 4284 0 net38
rlabel via1 5289 8716 5289 8716 0 net39
rlabel metal2 9360 33600 9360 33600 0 net4
rlabel metal2 6081 7896 6081 7896 0 net40
rlabel metal2 5472 21588 5472 21588 0 net41
rlabel metal3 9408 8820 9408 8820 0 net42
rlabel metal2 5664 21504 5664 21504 0 net43
rlabel metal2 6432 9408 6432 9408 0 net44
rlabel metal2 5952 21546 5952 21546 0 net45
rlabel metal4 5376 21000 5376 21000 0 net46
rlabel metal2 5760 16296 5760 16296 0 net47
rlabel metal2 8592 4368 8592 4368 0 net48
rlabel metal2 6144 16170 6144 16170 0 net49
rlabel metal2 1488 27090 1488 27090 0 net5
rlabel metal2 6048 21672 6048 21672 0 net50
rlabel metal2 6672 33516 6672 33516 0 net51
rlabel metal2 10200 6300 10200 6300 0 net52
rlabel metal2 6960 14700 6960 14700 0 net53
rlabel metal2 7488 22302 7488 22302 0 net54
rlabel metal2 8928 27468 8928 27468 0 net55
rlabel metal2 11928 14616 11928 14616 0 net56
rlabel metal2 9144 17892 9144 17892 0 net57
rlabel metal4 6816 17976 6816 17976 0 net58
rlabel metal2 9384 14532 9384 14532 0 net59
rlabel metal2 3552 37464 3552 37464 0 net6
rlabel metal5 8448 14994 8448 14994 0 net60
rlabel metal4 12528 17976 12528 17976 0 net61
rlabel metal4 12000 16338 12000 16338 0 net62
rlabel metal4 12000 17052 12000 17052 0 net63
rlabel metal2 8544 22344 8544 22344 0 net64
rlabel metal2 12240 14238 12240 14238 0 net65
rlabel via1 5758 14784 5758 14784 0 net66
rlabel metal2 2813 14616 2813 14616 0 net67
rlabel metal2 2544 24528 2544 24528 0 net68
rlabel metal2 8232 20580 8232 20580 0 net69
rlabel metal2 3168 36582 3168 36582 0 net7
rlabel metal2 8712 21000 8712 21000 0 net70
rlabel metal2 9264 19992 9264 19992 0 net71
rlabel metal2 4032 19320 4032 19320 0 net72
rlabel metal2 8088 20076 8088 20076 0 net73
rlabel metal2 9552 16968 9552 16968 0 net74
rlabel metal2 6048 22848 6048 22848 0 net75
rlabel metal2 8880 39648 8880 39648 0 net76
rlabel metal2 6720 31290 6720 31290 0 net77
rlabel metal2 7680 20832 7680 20832 0 net78
rlabel metal2 4848 18480 4848 18480 0 net79
rlabel metal2 1488 29526 1488 29526 0 net8
rlabel metal2 4320 35826 4320 35826 0 net80
rlabel metal3 5568 27300 5568 27300 0 net81
rlabel metal2 3360 20832 3360 20832 0 net82
rlabel metal2 4320 13944 4320 13944 0 net83
rlabel metal2 7632 25368 7632 25368 0 net84
rlabel metal2 4176 21504 4176 21504 0 net85
rlabel metal2 10440 17976 10440 17976 0 net86
rlabel metal2 10224 17724 10224 17724 0 net87
rlabel metal2 8544 11676 8544 11676 0 net88
rlabel metal4 9312 13356 9312 13356 0 net89
rlabel metal2 1488 31122 1488 31122 0 net9
rlabel metal2 10656 17052 10656 17052 0 net90
rlabel metal2 8496 5712 8496 5712 0 net91
rlabel metal3 11328 18606 11328 18606 0 net92
rlabel metal2 8712 14196 8712 14196 0 net93
rlabel metal2 9528 14196 9528 14196 0 net94
rlabel metal4 8640 21672 8640 21672 0 net95
rlabel metal2 8016 22260 8016 22260 0 net96
rlabel metal2 10416 12516 10416 12516 0 net97
rlabel metal3 8160 6300 8160 6300 0 net98
rlabel metal4 4992 14784 4992 14784 0 net99
<< properties >>
string FIXED_BBOX 0 0 13728 48384
<< end >>
