VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO RegFile
  CLASS BLOCK ;
  FOREIGN RegFile ;
  ORIGIN 0.000 0.000 ;
  SIZE 266.400 BY 241.920 ;
  PIN E1BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 265.950 94.300 266.400 94.700 ;
    END
  END E1BEG[0]
  PIN E1BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 265.950 95.980 266.400 96.380 ;
    END
  END E1BEG[1]
  PIN E1BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 265.950 97.660 266.400 98.060 ;
    END
  END E1BEG[2]
  PIN E1BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 265.950 99.340 266.400 99.740 ;
    END
  END E1BEG[3]
  PIN E1END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 94.300 0.450 94.700 ;
    END
  END E1END[0]
  PIN E1END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.450800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 95.980 0.450 96.380 ;
    END
  END E1END[1]
  PIN E1END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 97.660 0.450 98.060 ;
    END
  END E1END[2]
  PIN E1END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 99.340 0.450 99.740 ;
    END
  END E1END[3]
  PIN E2BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 265.950 101.020 266.400 101.420 ;
    END
  END E2BEG[0]
  PIN E2BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 265.950 102.700 266.400 103.100 ;
    END
  END E2BEG[1]
  PIN E2BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 265.950 104.380 266.400 104.780 ;
    END
  END E2BEG[2]
  PIN E2BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 265.950 106.060 266.400 106.460 ;
    END
  END E2BEG[3]
  PIN E2BEG[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 265.950 107.740 266.400 108.140 ;
    END
  END E2BEG[4]
  PIN E2BEG[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.827200 ;
    PORT
      LAYER Metal2 ;
        RECT 265.950 109.420 266.400 109.820 ;
    END
  END E2BEG[5]
  PIN E2BEG[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 265.950 111.100 266.400 111.500 ;
    END
  END E2BEG[6]
  PIN E2BEG[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 265.950 112.780 266.400 113.180 ;
    END
  END E2BEG[7]
  PIN E2BEGb[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 265.950 114.460 266.400 114.860 ;
    END
  END E2BEGb[0]
  PIN E2BEGb[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 265.950 116.140 266.400 116.540 ;
    END
  END E2BEGb[1]
  PIN E2BEGb[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 265.950 117.820 266.400 118.220 ;
    END
  END E2BEGb[2]
  PIN E2BEGb[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 265.950 119.500 266.400 119.900 ;
    END
  END E2BEGb[3]
  PIN E2BEGb[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 265.950 121.180 266.400 121.580 ;
    END
  END E2BEGb[4]
  PIN E2BEGb[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 265.950 122.860 266.400 123.260 ;
    END
  END E2BEGb[5]
  PIN E2BEGb[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 265.950 124.540 266.400 124.940 ;
    END
  END E2BEGb[6]
  PIN E2BEGb[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 265.950 126.220 266.400 126.620 ;
    END
  END E2BEGb[7]
  PIN E2END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 114.460 0.450 114.860 ;
    END
  END E2END[0]
  PIN E2END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 116.140 0.450 116.540 ;
    END
  END E2END[1]
  PIN E2END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 117.820 0.450 118.220 ;
    END
  END E2END[2]
  PIN E2END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 119.500 0.450 119.900 ;
    END
  END E2END[3]
  PIN E2END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 121.180 0.450 121.580 ;
    END
  END E2END[4]
  PIN E2END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 122.860 0.450 123.260 ;
    END
  END E2END[5]
  PIN E2END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 124.540 0.450 124.940 ;
    END
  END E2END[6]
  PIN E2END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 126.220 0.450 126.620 ;
    END
  END E2END[7]
  PIN E2MID[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 101.020 0.450 101.420 ;
    END
  END E2MID[0]
  PIN E2MID[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 102.700 0.450 103.100 ;
    END
  END E2MID[1]
  PIN E2MID[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 104.380 0.450 104.780 ;
    END
  END E2MID[2]
  PIN E2MID[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 106.060 0.450 106.460 ;
    END
  END E2MID[3]
  PIN E2MID[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 107.740 0.450 108.140 ;
    END
  END E2MID[4]
  PIN E2MID[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 109.420 0.450 109.820 ;
    END
  END E2MID[5]
  PIN E2MID[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 111.100 0.450 111.500 ;
    END
  END E2MID[6]
  PIN E2MID[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 112.780 0.450 113.180 ;
    END
  END E2MID[7]
  PIN E6BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 265.950 154.780 266.400 155.180 ;
    END
  END E6BEG[0]
  PIN E6BEG[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 265.950 171.580 266.400 171.980 ;
    END
  END E6BEG[10]
  PIN E6BEG[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 265.950 173.260 266.400 173.660 ;
    END
  END E6BEG[11]
  PIN E6BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 265.950 156.460 266.400 156.860 ;
    END
  END E6BEG[1]
  PIN E6BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 265.950 158.140 266.400 158.540 ;
    END
  END E6BEG[2]
  PIN E6BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 265.950 159.820 266.400 160.220 ;
    END
  END E6BEG[3]
  PIN E6BEG[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 265.950 161.500 266.400 161.900 ;
    END
  END E6BEG[4]
  PIN E6BEG[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 265.950 163.180 266.400 163.580 ;
    END
  END E6BEG[5]
  PIN E6BEG[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 265.950 164.860 266.400 165.260 ;
    END
  END E6BEG[6]
  PIN E6BEG[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 265.950 166.540 266.400 166.940 ;
    END
  END E6BEG[7]
  PIN E6BEG[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 265.950 168.220 266.400 168.620 ;
    END
  END E6BEG[8]
  PIN E6BEG[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 265.950 169.900 266.400 170.300 ;
    END
  END E6BEG[9]
  PIN E6END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.361400 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 154.780 0.450 155.180 ;
    END
  END E6END[0]
  PIN E6END[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 171.580 0.450 171.980 ;
    END
  END E6END[10]
  PIN E6END[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 173.260 0.450 173.660 ;
    END
  END E6END[11]
  PIN E6END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.361400 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 156.460 0.450 156.860 ;
    END
  END E6END[1]
  PIN E6END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 158.140 0.450 158.540 ;
    END
  END E6END[2]
  PIN E6END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 159.820 0.450 160.220 ;
    END
  END E6END[3]
  PIN E6END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 161.500 0.450 161.900 ;
    END
  END E6END[4]
  PIN E6END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 163.180 0.450 163.580 ;
    END
  END E6END[5]
  PIN E6END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 164.860 0.450 165.260 ;
    END
  END E6END[6]
  PIN E6END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 166.540 0.450 166.940 ;
    END
  END E6END[7]
  PIN E6END[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 168.220 0.450 168.620 ;
    END
  END E6END[8]
  PIN E6END[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 169.900 0.450 170.300 ;
    END
  END E6END[9]
  PIN EE4BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 265.950 127.900 266.400 128.300 ;
    END
  END EE4BEG[0]
  PIN EE4BEG[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 265.950 144.700 266.400 145.100 ;
    END
  END EE4BEG[10]
  PIN EE4BEG[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 265.950 146.380 266.400 146.780 ;
    END
  END EE4BEG[11]
  PIN EE4BEG[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 265.950 148.060 266.400 148.460 ;
    END
  END EE4BEG[12]
  PIN EE4BEG[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 265.950 149.740 266.400 150.140 ;
    END
  END EE4BEG[13]
  PIN EE4BEG[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 265.950 151.420 266.400 151.820 ;
    END
  END EE4BEG[14]
  PIN EE4BEG[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 265.950 153.100 266.400 153.500 ;
    END
  END EE4BEG[15]
  PIN EE4BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 265.950 129.580 266.400 129.980 ;
    END
  END EE4BEG[1]
  PIN EE4BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 265.950 131.260 266.400 131.660 ;
    END
  END EE4BEG[2]
  PIN EE4BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 265.950 132.940 266.400 133.340 ;
    END
  END EE4BEG[3]
  PIN EE4BEG[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 265.950 134.620 266.400 135.020 ;
    END
  END EE4BEG[4]
  PIN EE4BEG[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 265.950 136.300 266.400 136.700 ;
    END
  END EE4BEG[5]
  PIN EE4BEG[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 265.950 137.980 266.400 138.380 ;
    END
  END EE4BEG[6]
  PIN EE4BEG[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 265.950 139.660 266.400 140.060 ;
    END
  END EE4BEG[7]
  PIN EE4BEG[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 265.950 141.340 266.400 141.740 ;
    END
  END EE4BEG[8]
  PIN EE4BEG[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 265.950 143.020 266.400 143.420 ;
    END
  END EE4BEG[9]
  PIN EE4END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 127.900 0.450 128.300 ;
    END
  END EE4END[0]
  PIN EE4END[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 144.700 0.450 145.100 ;
    END
  END EE4END[10]
  PIN EE4END[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 146.380 0.450 146.780 ;
    END
  END EE4END[11]
  PIN EE4END[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 148.060 0.450 148.460 ;
    END
  END EE4END[12]
  PIN EE4END[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 149.740 0.450 150.140 ;
    END
  END EE4END[13]
  PIN EE4END[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 151.420 0.450 151.820 ;
    END
  END EE4END[14]
  PIN EE4END[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 153.100 0.450 153.500 ;
    END
  END EE4END[15]
  PIN EE4END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 129.580 0.450 129.980 ;
    END
  END EE4END[1]
  PIN EE4END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 131.260 0.450 131.660 ;
    END
  END EE4END[2]
  PIN EE4END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 132.940 0.450 133.340 ;
    END
  END EE4END[3]
  PIN EE4END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 134.620 0.450 135.020 ;
    END
  END EE4END[4]
  PIN EE4END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 136.300 0.450 136.700 ;
    END
  END EE4END[5]
  PIN EE4END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 137.980 0.450 138.380 ;
    END
  END EE4END[6]
  PIN EE4END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 139.660 0.450 140.060 ;
    END
  END EE4END[7]
  PIN EE4END[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 141.340 0.450 141.740 ;
    END
  END EE4END[8]
  PIN EE4END[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 143.020 0.450 143.420 ;
    END
  END EE4END[9]
  PIN FrameData[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.361400 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 174.940 0.450 175.340 ;
    END
  END FrameData[0]
  PIN FrameData[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 191.740 0.450 192.140 ;
    END
  END FrameData[10]
  PIN FrameData[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 193.420 0.450 193.820 ;
    END
  END FrameData[11]
  PIN FrameData[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.361400 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 195.100 0.450 195.500 ;
    END
  END FrameData[12]
  PIN FrameData[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 196.780 0.450 197.180 ;
    END
  END FrameData[13]
  PIN FrameData[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 198.460 0.450 198.860 ;
    END
  END FrameData[14]
  PIN FrameData[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 200.140 0.450 200.540 ;
    END
  END FrameData[15]
  PIN FrameData[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 201.820 0.450 202.220 ;
    END
  END FrameData[16]
  PIN FrameData[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 203.500 0.450 203.900 ;
    END
  END FrameData[17]
  PIN FrameData[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 205.180 0.450 205.580 ;
    END
  END FrameData[18]
  PIN FrameData[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 206.860 0.450 207.260 ;
    END
  END FrameData[19]
  PIN FrameData[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.361400 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 176.620 0.450 177.020 ;
    END
  END FrameData[1]
  PIN FrameData[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.361400 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 208.540 0.450 208.940 ;
    END
  END FrameData[20]
  PIN FrameData[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.361400 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 210.220 0.450 210.620 ;
    END
  END FrameData[21]
  PIN FrameData[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.361400 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 211.900 0.450 212.300 ;
    END
  END FrameData[22]
  PIN FrameData[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 213.580 0.450 213.980 ;
    END
  END FrameData[23]
  PIN FrameData[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.361400 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 215.260 0.450 215.660 ;
    END
  END FrameData[24]
  PIN FrameData[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.361400 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 216.940 0.450 217.340 ;
    END
  END FrameData[25]
  PIN FrameData[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 218.620 0.450 219.020 ;
    END
  END FrameData[26]
  PIN FrameData[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.361400 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 220.300 0.450 220.700 ;
    END
  END FrameData[27]
  PIN FrameData[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 221.980 0.450 222.380 ;
    END
  END FrameData[28]
  PIN FrameData[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.361400 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 223.660 0.450 224.060 ;
    END
  END FrameData[29]
  PIN FrameData[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 178.300 0.450 178.700 ;
    END
  END FrameData[2]
  PIN FrameData[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 225.340 0.450 225.740 ;
    END
  END FrameData[30]
  PIN FrameData[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.361400 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 227.020 0.450 227.420 ;
    END
  END FrameData[31]
  PIN FrameData[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.361400 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 179.980 0.450 180.380 ;
    END
  END FrameData[3]
  PIN FrameData[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 181.660 0.450 182.060 ;
    END
  END FrameData[4]
  PIN FrameData[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 183.340 0.450 183.740 ;
    END
  END FrameData[5]
  PIN FrameData[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 185.020 0.450 185.420 ;
    END
  END FrameData[6]
  PIN FrameData[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 186.700 0.450 187.100 ;
    END
  END FrameData[7]
  PIN FrameData[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 188.380 0.450 188.780 ;
    END
  END FrameData[8]
  PIN FrameData[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 190.060 0.450 190.460 ;
    END
  END FrameData[9]
  PIN FrameData_O[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 265.950 174.940 266.400 175.340 ;
    END
  END FrameData_O[0]
  PIN FrameData_O[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 265.950 191.740 266.400 192.140 ;
    END
  END FrameData_O[10]
  PIN FrameData_O[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 265.950 193.420 266.400 193.820 ;
    END
  END FrameData_O[11]
  PIN FrameData_O[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 265.950 195.100 266.400 195.500 ;
    END
  END FrameData_O[12]
  PIN FrameData_O[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 265.950 196.780 266.400 197.180 ;
    END
  END FrameData_O[13]
  PIN FrameData_O[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 265.950 198.460 266.400 198.860 ;
    END
  END FrameData_O[14]
  PIN FrameData_O[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 265.950 200.140 266.400 200.540 ;
    END
  END FrameData_O[15]
  PIN FrameData_O[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 265.950 201.820 266.400 202.220 ;
    END
  END FrameData_O[16]
  PIN FrameData_O[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 265.950 203.500 266.400 203.900 ;
    END
  END FrameData_O[17]
  PIN FrameData_O[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 265.950 205.180 266.400 205.580 ;
    END
  END FrameData_O[18]
  PIN FrameData_O[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 265.950 206.860 266.400 207.260 ;
    END
  END FrameData_O[19]
  PIN FrameData_O[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 265.950 176.620 266.400 177.020 ;
    END
  END FrameData_O[1]
  PIN FrameData_O[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 265.950 208.540 266.400 208.940 ;
    END
  END FrameData_O[20]
  PIN FrameData_O[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 265.950 210.220 266.400 210.620 ;
    END
  END FrameData_O[21]
  PIN FrameData_O[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 265.950 211.900 266.400 212.300 ;
    END
  END FrameData_O[22]
  PIN FrameData_O[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 265.950 213.580 266.400 213.980 ;
    END
  END FrameData_O[23]
  PIN FrameData_O[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 265.950 215.260 266.400 215.660 ;
    END
  END FrameData_O[24]
  PIN FrameData_O[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 265.950 216.940 266.400 217.340 ;
    END
  END FrameData_O[25]
  PIN FrameData_O[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 265.950 218.620 266.400 219.020 ;
    END
  END FrameData_O[26]
  PIN FrameData_O[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 265.950 220.300 266.400 220.700 ;
    END
  END FrameData_O[27]
  PIN FrameData_O[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 265.950 221.980 266.400 222.380 ;
    END
  END FrameData_O[28]
  PIN FrameData_O[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 265.950 223.660 266.400 224.060 ;
    END
  END FrameData_O[29]
  PIN FrameData_O[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 265.950 178.300 266.400 178.700 ;
    END
  END FrameData_O[2]
  PIN FrameData_O[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 265.950 225.340 266.400 225.740 ;
    END
  END FrameData_O[30]
  PIN FrameData_O[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 265.950 227.020 266.400 227.420 ;
    END
  END FrameData_O[31]
  PIN FrameData_O[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 265.950 179.980 266.400 180.380 ;
    END
  END FrameData_O[3]
  PIN FrameData_O[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 265.950 181.660 266.400 182.060 ;
    END
  END FrameData_O[4]
  PIN FrameData_O[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 265.950 183.340 266.400 183.740 ;
    END
  END FrameData_O[5]
  PIN FrameData_O[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 265.950 185.020 266.400 185.420 ;
    END
  END FrameData_O[6]
  PIN FrameData_O[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 265.950 186.700 266.400 187.100 ;
    END
  END FrameData_O[7]
  PIN FrameData_O[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 265.950 188.380 266.400 188.780 ;
    END
  END FrameData_O[8]
  PIN FrameData_O[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 265.950 190.060 266.400 190.460 ;
    END
  END FrameData_O[9]
  PIN FrameStrobe[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 215.320 0.000 215.720 0.400 ;
    END
  END FrameStrobe[0]
  PIN FrameStrobe[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 234.520 0.000 234.920 0.400 ;
    END
  END FrameStrobe[10]
  PIN FrameStrobe[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 236.440 0.000 236.840 0.400 ;
    END
  END FrameStrobe[11]
  PIN FrameStrobe[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 238.360 0.000 238.760 0.400 ;
    END
  END FrameStrobe[12]
  PIN FrameStrobe[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 240.280 0.000 240.680 0.400 ;
    END
  END FrameStrobe[13]
  PIN FrameStrobe[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 242.200 0.000 242.600 0.400 ;
    END
  END FrameStrobe[14]
  PIN FrameStrobe[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 244.120 0.000 244.520 0.400 ;
    END
  END FrameStrobe[15]
  PIN FrameStrobe[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 246.040 0.000 246.440 0.400 ;
    END
  END FrameStrobe[16]
  PIN FrameStrobe[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 247.960 0.000 248.360 0.400 ;
    END
  END FrameStrobe[17]
  PIN FrameStrobe[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 249.880 0.000 250.280 0.400 ;
    END
  END FrameStrobe[18]
  PIN FrameStrobe[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 251.800 0.000 252.200 0.400 ;
    END
  END FrameStrobe[19]
  PIN FrameStrobe[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 217.240 0.000 217.640 0.400 ;
    END
  END FrameStrobe[1]
  PIN FrameStrobe[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 219.160 0.000 219.560 0.400 ;
    END
  END FrameStrobe[2]
  PIN FrameStrobe[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 221.080 0.000 221.480 0.400 ;
    END
  END FrameStrobe[3]
  PIN FrameStrobe[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 223.000 0.000 223.400 0.400 ;
    END
  END FrameStrobe[4]
  PIN FrameStrobe[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 224.920 0.000 225.320 0.400 ;
    END
  END FrameStrobe[5]
  PIN FrameStrobe[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 226.840 0.000 227.240 0.400 ;
    END
  END FrameStrobe[6]
  PIN FrameStrobe[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 228.760 0.000 229.160 0.400 ;
    END
  END FrameStrobe[7]
  PIN FrameStrobe[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.542100 ;
    PORT
      LAYER Metal3 ;
        RECT 230.680 0.000 231.080 0.400 ;
    END
  END FrameStrobe[8]
  PIN FrameStrobe[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 232.600 0.000 233.000 0.400 ;
    END
  END FrameStrobe[9]
  PIN FrameStrobe_O[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 215.320 241.520 215.720 241.920 ;
    END
  END FrameStrobe_O[0]
  PIN FrameStrobe_O[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 234.520 241.520 234.920 241.920 ;
    END
  END FrameStrobe_O[10]
  PIN FrameStrobe_O[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 236.440 241.520 236.840 241.920 ;
    END
  END FrameStrobe_O[11]
  PIN FrameStrobe_O[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 238.360 241.520 238.760 241.920 ;
    END
  END FrameStrobe_O[12]
  PIN FrameStrobe_O[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 240.280 241.520 240.680 241.920 ;
    END
  END FrameStrobe_O[13]
  PIN FrameStrobe_O[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 242.200 241.520 242.600 241.920 ;
    END
  END FrameStrobe_O[14]
  PIN FrameStrobe_O[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 244.120 241.520 244.520 241.920 ;
    END
  END FrameStrobe_O[15]
  PIN FrameStrobe_O[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 246.040 241.520 246.440 241.920 ;
    END
  END FrameStrobe_O[16]
  PIN FrameStrobe_O[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 247.960 241.520 248.360 241.920 ;
    END
  END FrameStrobe_O[17]
  PIN FrameStrobe_O[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 249.880 241.520 250.280 241.920 ;
    END
  END FrameStrobe_O[18]
  PIN FrameStrobe_O[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 251.800 241.520 252.200 241.920 ;
    END
  END FrameStrobe_O[19]
  PIN FrameStrobe_O[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 217.240 241.520 217.640 241.920 ;
    END
  END FrameStrobe_O[1]
  PIN FrameStrobe_O[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 219.160 241.520 219.560 241.920 ;
    END
  END FrameStrobe_O[2]
  PIN FrameStrobe_O[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 221.080 241.520 221.480 241.920 ;
    END
  END FrameStrobe_O[3]
  PIN FrameStrobe_O[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 223.000 241.520 223.400 241.920 ;
    END
  END FrameStrobe_O[4]
  PIN FrameStrobe_O[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 224.920 241.520 225.320 241.920 ;
    END
  END FrameStrobe_O[5]
  PIN FrameStrobe_O[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 226.840 241.520 227.240 241.920 ;
    END
  END FrameStrobe_O[6]
  PIN FrameStrobe_O[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 228.760 241.520 229.160 241.920 ;
    END
  END FrameStrobe_O[7]
  PIN FrameStrobe_O[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 230.680 241.520 231.080 241.920 ;
    END
  END FrameStrobe_O[8]
  PIN FrameStrobe_O[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 232.600 241.520 233.000 241.920 ;
    END
  END FrameStrobe_O[9]
  PIN N1BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 13.720 241.520 14.120 241.920 ;
    END
  END N1BEG[0]
  PIN N1BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 15.640 241.520 16.040 241.920 ;
    END
  END N1BEG[1]
  PIN N1BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 17.560 241.520 17.960 241.920 ;
    END
  END N1BEG[2]
  PIN N1BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 19.480 241.520 19.880 241.920 ;
    END
  END N1BEG[3]
  PIN N1END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 13.720 0.000 14.120 0.400 ;
    END
  END N1END[0]
  PIN N1END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.450800 ;
    PORT
      LAYER Metal3 ;
        RECT 15.640 0.000 16.040 0.400 ;
    END
  END N1END[1]
  PIN N1END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 17.560 0.000 17.960 0.400 ;
    END
  END N1END[2]
  PIN N1END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 19.480 0.000 19.880 0.400 ;
    END
  END N1END[3]
  PIN N2BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 21.400 241.520 21.800 241.920 ;
    END
  END N2BEG[0]
  PIN N2BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 23.320 241.520 23.720 241.920 ;
    END
  END N2BEG[1]
  PIN N2BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 25.240 241.520 25.640 241.920 ;
    END
  END N2BEG[2]
  PIN N2BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 27.160 241.520 27.560 241.920 ;
    END
  END N2BEG[3]
  PIN N2BEG[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 29.080 241.520 29.480 241.920 ;
    END
  END N2BEG[4]
  PIN N2BEG[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 31.000 241.520 31.400 241.920 ;
    END
  END N2BEG[5]
  PIN N2BEG[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 32.920 241.520 33.320 241.920 ;
    END
  END N2BEG[6]
  PIN N2BEG[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 34.840 241.520 35.240 241.920 ;
    END
  END N2BEG[7]
  PIN N2BEGb[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 36.760 241.520 37.160 241.920 ;
    END
  END N2BEGb[0]
  PIN N2BEGb[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 38.680 241.520 39.080 241.920 ;
    END
  END N2BEGb[1]
  PIN N2BEGb[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 40.600 241.520 41.000 241.920 ;
    END
  END N2BEGb[2]
  PIN N2BEGb[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 42.520 241.520 42.920 241.920 ;
    END
  END N2BEGb[3]
  PIN N2BEGb[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 44.440 241.520 44.840 241.920 ;
    END
  END N2BEGb[4]
  PIN N2BEGb[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 46.360 241.520 46.760 241.920 ;
    END
  END N2BEGb[5]
  PIN N2BEGb[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 48.280 241.520 48.680 241.920 ;
    END
  END N2BEGb[6]
  PIN N2BEGb[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 50.200 241.520 50.600 241.920 ;
    END
  END N2BEGb[7]
  PIN N2END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 36.760 0.000 37.160 0.400 ;
    END
  END N2END[0]
  PIN N2END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 38.680 0.000 39.080 0.400 ;
    END
  END N2END[1]
  PIN N2END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 40.600 0.000 41.000 0.400 ;
    END
  END N2END[2]
  PIN N2END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 42.520 0.000 42.920 0.400 ;
    END
  END N2END[3]
  PIN N2END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 44.440 0.000 44.840 0.400 ;
    END
  END N2END[4]
  PIN N2END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213200 ;
    PORT
      LAYER Metal3 ;
        RECT 46.360 0.000 46.760 0.400 ;
    END
  END N2END[5]
  PIN N2END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 48.280 0.000 48.680 0.400 ;
    END
  END N2END[6]
  PIN N2END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 50.200 0.000 50.600 0.400 ;
    END
  END N2END[7]
  PIN N2MID[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 21.400 0.000 21.800 0.400 ;
    END
  END N2MID[0]
  PIN N2MID[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 23.320 0.000 23.720 0.400 ;
    END
  END N2MID[1]
  PIN N2MID[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 25.240 0.000 25.640 0.400 ;
    END
  END N2MID[2]
  PIN N2MID[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 27.160 0.000 27.560 0.400 ;
    END
  END N2MID[3]
  PIN N2MID[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 29.080 0.000 29.480 0.400 ;
    END
  END N2MID[4]
  PIN N2MID[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 31.000 0.000 31.400 0.400 ;
    END
  END N2MID[5]
  PIN N2MID[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 32.920 0.000 33.320 0.400 ;
    END
  END N2MID[6]
  PIN N2MID[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 34.840 0.000 35.240 0.400 ;
    END
  END N2MID[7]
  PIN N4BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 52.120 241.520 52.520 241.920 ;
    END
  END N4BEG[0]
  PIN N4BEG[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 71.320 241.520 71.720 241.920 ;
    END
  END N4BEG[10]
  PIN N4BEG[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 73.240 241.520 73.640 241.920 ;
    END
  END N4BEG[11]
  PIN N4BEG[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 75.160 241.520 75.560 241.920 ;
    END
  END N4BEG[12]
  PIN N4BEG[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 77.080 241.520 77.480 241.920 ;
    END
  END N4BEG[13]
  PIN N4BEG[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 79.000 241.520 79.400 241.920 ;
    END
  END N4BEG[14]
  PIN N4BEG[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 80.920 241.520 81.320 241.920 ;
    END
  END N4BEG[15]
  PIN N4BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 54.040 241.520 54.440 241.920 ;
    END
  END N4BEG[1]
  PIN N4BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 55.960 241.520 56.360 241.920 ;
    END
  END N4BEG[2]
  PIN N4BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 57.880 241.520 58.280 241.920 ;
    END
  END N4BEG[3]
  PIN N4BEG[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 59.800 241.520 60.200 241.920 ;
    END
  END N4BEG[4]
  PIN N4BEG[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 61.720 241.520 62.120 241.920 ;
    END
  END N4BEG[5]
  PIN N4BEG[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 63.640 241.520 64.040 241.920 ;
    END
  END N4BEG[6]
  PIN N4BEG[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 65.560 241.520 65.960 241.920 ;
    END
  END N4BEG[7]
  PIN N4BEG[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 67.480 241.520 67.880 241.920 ;
    END
  END N4BEG[8]
  PIN N4BEG[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 69.400 241.520 69.800 241.920 ;
    END
  END N4BEG[9]
  PIN N4END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 52.120 0.000 52.520 0.400 ;
    END
  END N4END[0]
  PIN N4END[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 71.320 0.000 71.720 0.400 ;
    END
  END N4END[10]
  PIN N4END[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 73.240 0.000 73.640 0.400 ;
    END
  END N4END[11]
  PIN N4END[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 75.160 0.000 75.560 0.400 ;
    END
  END N4END[12]
  PIN N4END[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 77.080 0.000 77.480 0.400 ;
    END
  END N4END[13]
  PIN N4END[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 79.000 0.000 79.400 0.400 ;
    END
  END N4END[14]
  PIN N4END[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 80.920 0.000 81.320 0.400 ;
    END
  END N4END[15]
  PIN N4END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 54.040 0.000 54.440 0.400 ;
    END
  END N4END[1]
  PIN N4END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 55.960 0.000 56.360 0.400 ;
    END
  END N4END[2]
  PIN N4END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 57.880 0.000 58.280 0.400 ;
    END
  END N4END[3]
  PIN N4END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 59.800 0.000 60.200 0.400 ;
    END
  END N4END[4]
  PIN N4END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 61.720 0.000 62.120 0.400 ;
    END
  END N4END[5]
  PIN N4END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 63.640 0.000 64.040 0.400 ;
    END
  END N4END[6]
  PIN N4END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 65.560 0.000 65.960 0.400 ;
    END
  END N4END[7]
  PIN N4END[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 67.480 0.000 67.880 0.400 ;
    END
  END N4END[8]
  PIN N4END[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 69.400 0.000 69.800 0.400 ;
    END
  END N4END[9]
  PIN NN4BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 82.840 241.520 83.240 241.920 ;
    END
  END NN4BEG[0]
  PIN NN4BEG[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 102.040 241.520 102.440 241.920 ;
    END
  END NN4BEG[10]
  PIN NN4BEG[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 103.960 241.520 104.360 241.920 ;
    END
  END NN4BEG[11]
  PIN NN4BEG[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 105.880 241.520 106.280 241.920 ;
    END
  END NN4BEG[12]
  PIN NN4BEG[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 107.800 241.520 108.200 241.920 ;
    END
  END NN4BEG[13]
  PIN NN4BEG[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 109.720 241.520 110.120 241.920 ;
    END
  END NN4BEG[14]
  PIN NN4BEG[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 111.640 241.520 112.040 241.920 ;
    END
  END NN4BEG[15]
  PIN NN4BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 84.760 241.520 85.160 241.920 ;
    END
  END NN4BEG[1]
  PIN NN4BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 86.680 241.520 87.080 241.920 ;
    END
  END NN4BEG[2]
  PIN NN4BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 88.600 241.520 89.000 241.920 ;
    END
  END NN4BEG[3]
  PIN NN4BEG[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 90.520 241.520 90.920 241.920 ;
    END
  END NN4BEG[4]
  PIN NN4BEG[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 92.440 241.520 92.840 241.920 ;
    END
  END NN4BEG[5]
  PIN NN4BEG[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 94.360 241.520 94.760 241.920 ;
    END
  END NN4BEG[6]
  PIN NN4BEG[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 96.280 241.520 96.680 241.920 ;
    END
  END NN4BEG[7]
  PIN NN4BEG[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 98.200 241.520 98.600 241.920 ;
    END
  END NN4BEG[8]
  PIN NN4BEG[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 100.120 241.520 100.520 241.920 ;
    END
  END NN4BEG[9]
  PIN NN4END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 82.840 0.000 83.240 0.400 ;
    END
  END NN4END[0]
  PIN NN4END[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 102.040 0.000 102.440 0.400 ;
    END
  END NN4END[10]
  PIN NN4END[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 103.960 0.000 104.360 0.400 ;
    END
  END NN4END[11]
  PIN NN4END[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 105.880 0.000 106.280 0.400 ;
    END
  END NN4END[12]
  PIN NN4END[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 107.800 0.000 108.200 0.400 ;
    END
  END NN4END[13]
  PIN NN4END[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 109.720 0.000 110.120 0.400 ;
    END
  END NN4END[14]
  PIN NN4END[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 111.640 0.000 112.040 0.400 ;
    END
  END NN4END[15]
  PIN NN4END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 84.760 0.000 85.160 0.400 ;
    END
  END NN4END[1]
  PIN NN4END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 86.680 0.000 87.080 0.400 ;
    END
  END NN4END[2]
  PIN NN4END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.725400 ;
    PORT
      LAYER Metal3 ;
        RECT 88.600 0.000 89.000 0.400 ;
    END
  END NN4END[3]
  PIN NN4END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 90.520 0.000 90.920 0.400 ;
    END
  END NN4END[4]
  PIN NN4END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 92.440 0.000 92.840 0.400 ;
    END
  END NN4END[5]
  PIN NN4END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 94.360 0.000 94.760 0.400 ;
    END
  END NN4END[6]
  PIN NN4END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 96.280 0.000 96.680 0.400 ;
    END
  END NN4END[7]
  PIN NN4END[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 98.200 0.000 98.600 0.400 ;
    END
  END NN4END[8]
  PIN NN4END[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 100.120 0.000 100.520 0.400 ;
    END
  END NN4END[9]
  PIN S1BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 113.560 0.000 113.960 0.400 ;
    END
  END S1BEG[0]
  PIN S1BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 115.480 0.000 115.880 0.400 ;
    END
  END S1BEG[1]
  PIN S1BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 117.400 0.000 117.800 0.400 ;
    END
  END S1BEG[2]
  PIN S1BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 119.320 0.000 119.720 0.400 ;
    END
  END S1BEG[3]
  PIN S1END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 113.560 241.520 113.960 241.920 ;
    END
  END S1END[0]
  PIN S1END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213200 ;
    PORT
      LAYER Metal3 ;
        RECT 115.480 241.520 115.880 241.920 ;
    END
  END S1END[1]
  PIN S1END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 117.400 241.520 117.800 241.920 ;
    END
  END S1END[2]
  PIN S1END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 119.320 241.520 119.720 241.920 ;
    END
  END S1END[3]
  PIN S2BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 121.240 0.000 121.640 0.400 ;
    END
  END S2BEG[0]
  PIN S2BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 123.160 0.000 123.560 0.400 ;
    END
  END S2BEG[1]
  PIN S2BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 125.080 0.000 125.480 0.400 ;
    END
  END S2BEG[2]
  PIN S2BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 127.000 0.000 127.400 0.400 ;
    END
  END S2BEG[3]
  PIN S2BEG[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 128.920 0.000 129.320 0.400 ;
    END
  END S2BEG[4]
  PIN S2BEG[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 130.840 0.000 131.240 0.400 ;
    END
  END S2BEG[5]
  PIN S2BEG[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 132.760 0.000 133.160 0.400 ;
    END
  END S2BEG[6]
  PIN S2BEG[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 134.680 0.000 135.080 0.400 ;
    END
  END S2BEG[7]
  PIN S2BEGb[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 136.600 0.000 137.000 0.400 ;
    END
  END S2BEGb[0]
  PIN S2BEGb[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 138.520 0.000 138.920 0.400 ;
    END
  END S2BEGb[1]
  PIN S2BEGb[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 140.440 0.000 140.840 0.400 ;
    END
  END S2BEGb[2]
  PIN S2BEGb[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 142.360 0.000 142.760 0.400 ;
    END
  END S2BEGb[3]
  PIN S2BEGb[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 144.280 0.000 144.680 0.400 ;
    END
  END S2BEGb[4]
  PIN S2BEGb[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 146.200 0.000 146.600 0.400 ;
    END
  END S2BEGb[5]
  PIN S2BEGb[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 148.120 0.000 148.520 0.400 ;
    END
  END S2BEGb[6]
  PIN S2BEGb[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 150.040 0.000 150.440 0.400 ;
    END
  END S2BEGb[7]
  PIN S2END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 136.600 241.520 137.000 241.920 ;
    END
  END S2END[0]
  PIN S2END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 138.520 241.520 138.920 241.920 ;
    END
  END S2END[1]
  PIN S2END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 140.440 241.520 140.840 241.920 ;
    END
  END S2END[2]
  PIN S2END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 142.360 241.520 142.760 241.920 ;
    END
  END S2END[3]
  PIN S2END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 144.280 241.520 144.680 241.920 ;
    END
  END S2END[4]
  PIN S2END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 146.200 241.520 146.600 241.920 ;
    END
  END S2END[5]
  PIN S2END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 148.120 241.520 148.520 241.920 ;
    END
  END S2END[6]
  PIN S2END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 150.040 241.520 150.440 241.920 ;
    END
  END S2END[7]
  PIN S2MID[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 121.240 241.520 121.640 241.920 ;
    END
  END S2MID[0]
  PIN S2MID[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 123.160 241.520 123.560 241.920 ;
    END
  END S2MID[1]
  PIN S2MID[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 125.080 241.520 125.480 241.920 ;
    END
  END S2MID[2]
  PIN S2MID[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 127.000 241.520 127.400 241.920 ;
    END
  END S2MID[3]
  PIN S2MID[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 128.920 241.520 129.320 241.920 ;
    END
  END S2MID[4]
  PIN S2MID[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 130.840 241.520 131.240 241.920 ;
    END
  END S2MID[5]
  PIN S2MID[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 132.760 241.520 133.160 241.920 ;
    END
  END S2MID[6]
  PIN S2MID[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 134.680 241.520 135.080 241.920 ;
    END
  END S2MID[7]
  PIN S4BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 151.960 0.000 152.360 0.400 ;
    END
  END S4BEG[0]
  PIN S4BEG[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 171.160 0.000 171.560 0.400 ;
    END
  END S4BEG[10]
  PIN S4BEG[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 173.080 0.000 173.480 0.400 ;
    END
  END S4BEG[11]
  PIN S4BEG[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 175.000 0.000 175.400 0.400 ;
    END
  END S4BEG[12]
  PIN S4BEG[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 176.920 0.000 177.320 0.400 ;
    END
  END S4BEG[13]
  PIN S4BEG[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 178.840 0.000 179.240 0.400 ;
    END
  END S4BEG[14]
  PIN S4BEG[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 180.760 0.000 181.160 0.400 ;
    END
  END S4BEG[15]
  PIN S4BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 153.880 0.000 154.280 0.400 ;
    END
  END S4BEG[1]
  PIN S4BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 155.800 0.000 156.200 0.400 ;
    END
  END S4BEG[2]
  PIN S4BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 157.720 0.000 158.120 0.400 ;
    END
  END S4BEG[3]
  PIN S4BEG[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 159.640 0.000 160.040 0.400 ;
    END
  END S4BEG[4]
  PIN S4BEG[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 161.560 0.000 161.960 0.400 ;
    END
  END S4BEG[5]
  PIN S4BEG[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 163.480 0.000 163.880 0.400 ;
    END
  END S4BEG[6]
  PIN S4BEG[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 165.400 0.000 165.800 0.400 ;
    END
  END S4BEG[7]
  PIN S4BEG[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 167.320 0.000 167.720 0.400 ;
    END
  END S4BEG[8]
  PIN S4BEG[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 169.240 0.000 169.640 0.400 ;
    END
  END S4BEG[9]
  PIN S4END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 151.960 241.520 152.360 241.920 ;
    END
  END S4END[0]
  PIN S4END[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 171.160 241.520 171.560 241.920 ;
    END
  END S4END[10]
  PIN S4END[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 173.080 241.520 173.480 241.920 ;
    END
  END S4END[11]
  PIN S4END[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 175.000 241.520 175.400 241.920 ;
    END
  END S4END[12]
  PIN S4END[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 176.920 241.520 177.320 241.920 ;
    END
  END S4END[13]
  PIN S4END[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 178.840 241.520 179.240 241.920 ;
    END
  END S4END[14]
  PIN S4END[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 180.760 241.520 181.160 241.920 ;
    END
  END S4END[15]
  PIN S4END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 153.880 241.520 154.280 241.920 ;
    END
  END S4END[1]
  PIN S4END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 155.800 241.520 156.200 241.920 ;
    END
  END S4END[2]
  PIN S4END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 157.720 241.520 158.120 241.920 ;
    END
  END S4END[3]
  PIN S4END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 159.640 241.520 160.040 241.920 ;
    END
  END S4END[4]
  PIN S4END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 161.560 241.520 161.960 241.920 ;
    END
  END S4END[5]
  PIN S4END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 163.480 241.520 163.880 241.920 ;
    END
  END S4END[6]
  PIN S4END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 165.400 241.520 165.800 241.920 ;
    END
  END S4END[7]
  PIN S4END[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 167.320 241.520 167.720 241.920 ;
    END
  END S4END[8]
  PIN S4END[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 169.240 241.520 169.640 241.920 ;
    END
  END S4END[9]
  PIN SS4BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 182.680 0.000 183.080 0.400 ;
    END
  END SS4BEG[0]
  PIN SS4BEG[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 201.880 0.000 202.280 0.400 ;
    END
  END SS4BEG[10]
  PIN SS4BEG[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 203.800 0.000 204.200 0.400 ;
    END
  END SS4BEG[11]
  PIN SS4BEG[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 205.720 0.000 206.120 0.400 ;
    END
  END SS4BEG[12]
  PIN SS4BEG[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 207.640 0.000 208.040 0.400 ;
    END
  END SS4BEG[13]
  PIN SS4BEG[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 209.560 0.000 209.960 0.400 ;
    END
  END SS4BEG[14]
  PIN SS4BEG[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 211.480 0.000 211.880 0.400 ;
    END
  END SS4BEG[15]
  PIN SS4BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 184.600 0.000 185.000 0.400 ;
    END
  END SS4BEG[1]
  PIN SS4BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 186.520 0.000 186.920 0.400 ;
    END
  END SS4BEG[2]
  PIN SS4BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 188.440 0.000 188.840 0.400 ;
    END
  END SS4BEG[3]
  PIN SS4BEG[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 190.360 0.000 190.760 0.400 ;
    END
  END SS4BEG[4]
  PIN SS4BEG[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 192.280 0.000 192.680 0.400 ;
    END
  END SS4BEG[5]
  PIN SS4BEG[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 194.200 0.000 194.600 0.400 ;
    END
  END SS4BEG[6]
  PIN SS4BEG[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 196.120 0.000 196.520 0.400 ;
    END
  END SS4BEG[7]
  PIN SS4BEG[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 198.040 0.000 198.440 0.400 ;
    END
  END SS4BEG[8]
  PIN SS4BEG[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 199.960 0.000 200.360 0.400 ;
    END
  END SS4BEG[9]
  PIN SS4END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 182.680 241.520 183.080 241.920 ;
    END
  END SS4END[0]
  PIN SS4END[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 201.880 241.520 202.280 241.920 ;
    END
  END SS4END[10]
  PIN SS4END[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 203.800 241.520 204.200 241.920 ;
    END
  END SS4END[11]
  PIN SS4END[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 205.720 241.520 206.120 241.920 ;
    END
  END SS4END[12]
  PIN SS4END[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 207.640 241.520 208.040 241.920 ;
    END
  END SS4END[13]
  PIN SS4END[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 209.560 241.520 209.960 241.920 ;
    END
  END SS4END[14]
  PIN SS4END[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 211.480 241.520 211.880 241.920 ;
    END
  END SS4END[15]
  PIN SS4END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 184.600 241.520 185.000 241.920 ;
    END
  END SS4END[1]
  PIN SS4END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 186.520 241.520 186.920 241.920 ;
    END
  END SS4END[2]
  PIN SS4END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 188.440 241.520 188.840 241.920 ;
    END
  END SS4END[3]
  PIN SS4END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 190.360 241.520 190.760 241.920 ;
    END
  END SS4END[4]
  PIN SS4END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 192.280 241.520 192.680 241.920 ;
    END
  END SS4END[5]
  PIN SS4END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 194.200 241.520 194.600 241.920 ;
    END
  END SS4END[6]
  PIN SS4END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 196.120 241.520 196.520 241.920 ;
    END
  END SS4END[7]
  PIN SS4END[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 198.040 241.520 198.440 241.920 ;
    END
  END SS4END[8]
  PIN SS4END[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 199.960 241.520 200.360 241.920 ;
    END
  END SS4END[9]
  PIN UserCLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 30.943899 ;
    PORT
      LAYER Metal3 ;
        RECT 213.400 0.000 213.800 0.400 ;
    END
  END UserCLK
  PIN UserCLKo
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 213.400 241.520 213.800 241.920 ;
    END
  END UserCLKo
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal5 ;
        RECT 24.460 0.000 26.660 241.920 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 100.060 0.000 102.260 241.920 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 175.660 0.000 177.860 241.920 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 251.260 0.000 253.460 241.920 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal5 ;
        RECT 18.260 0.000 20.460 241.920 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 93.860 0.000 96.060 241.920 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 169.460 0.000 171.660 241.920 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 245.060 0.000 247.260 241.920 ;
    END
  END VPWR
  PIN W1BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 13.660 0.450 14.060 ;
    END
  END W1BEG[0]
  PIN W1BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 15.340 0.450 15.740 ;
    END
  END W1BEG[1]
  PIN W1BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 17.020 0.450 17.420 ;
    END
  END W1BEG[2]
  PIN W1BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 18.700 0.450 19.100 ;
    END
  END W1BEG[3]
  PIN W1END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 265.950 13.660 266.400 14.060 ;
    END
  END W1END[0]
  PIN W1END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.725400 ;
    PORT
      LAYER Metal2 ;
        RECT 265.950 15.340 266.400 15.740 ;
    END
  END W1END[1]
  PIN W1END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 265.950 17.020 266.400 17.420 ;
    END
  END W1END[2]
  PIN W1END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 265.950 18.700 266.400 19.100 ;
    END
  END W1END[3]
  PIN W2BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 20.380 0.450 20.780 ;
    END
  END W2BEG[0]
  PIN W2BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 22.060 0.450 22.460 ;
    END
  END W2BEG[1]
  PIN W2BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 23.740 0.450 24.140 ;
    END
  END W2BEG[2]
  PIN W2BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 25.420 0.450 25.820 ;
    END
  END W2BEG[3]
  PIN W2BEG[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 27.100 0.450 27.500 ;
    END
  END W2BEG[4]
  PIN W2BEG[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 28.780 0.450 29.180 ;
    END
  END W2BEG[5]
  PIN W2BEG[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 30.460 0.450 30.860 ;
    END
  END W2BEG[6]
  PIN W2BEG[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 32.140 0.450 32.540 ;
    END
  END W2BEG[7]
  PIN W2BEGb[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 33.820 0.450 34.220 ;
    END
  END W2BEGb[0]
  PIN W2BEGb[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 35.500 0.450 35.900 ;
    END
  END W2BEGb[1]
  PIN W2BEGb[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 37.180 0.450 37.580 ;
    END
  END W2BEGb[2]
  PIN W2BEGb[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 38.860 0.450 39.260 ;
    END
  END W2BEGb[3]
  PIN W2BEGb[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 40.540 0.450 40.940 ;
    END
  END W2BEGb[4]
  PIN W2BEGb[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 42.220 0.450 42.620 ;
    END
  END W2BEGb[5]
  PIN W2BEGb[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 43.900 0.450 44.300 ;
    END
  END W2BEGb[6]
  PIN W2BEGb[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 45.580 0.450 45.980 ;
    END
  END W2BEGb[7]
  PIN W2END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 265.950 33.820 266.400 34.220 ;
    END
  END W2END[0]
  PIN W2END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 265.950 35.500 266.400 35.900 ;
    END
  END W2END[1]
  PIN W2END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 265.950 37.180 266.400 37.580 ;
    END
  END W2END[2]
  PIN W2END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 265.950 38.860 266.400 39.260 ;
    END
  END W2END[3]
  PIN W2END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 265.950 40.540 266.400 40.940 ;
    END
  END W2END[4]
  PIN W2END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 265.950 42.220 266.400 42.620 ;
    END
  END W2END[5]
  PIN W2END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 265.950 43.900 266.400 44.300 ;
    END
  END W2END[6]
  PIN W2END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 265.950 45.580 266.400 45.980 ;
    END
  END W2END[7]
  PIN W2MID[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 265.950 20.380 266.400 20.780 ;
    END
  END W2MID[0]
  PIN W2MID[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 265.950 22.060 266.400 22.460 ;
    END
  END W2MID[1]
  PIN W2MID[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 265.950 23.740 266.400 24.140 ;
    END
  END W2MID[2]
  PIN W2MID[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 265.950 25.420 266.400 25.820 ;
    END
  END W2MID[3]
  PIN W2MID[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 265.950 27.100 266.400 27.500 ;
    END
  END W2MID[4]
  PIN W2MID[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 265.950 28.780 266.400 29.180 ;
    END
  END W2MID[5]
  PIN W2MID[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 265.950 30.460 266.400 30.860 ;
    END
  END W2MID[6]
  PIN W2MID[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 265.950 32.140 266.400 32.540 ;
    END
  END W2MID[7]
  PIN W6BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 74.140 0.450 74.540 ;
    END
  END W6BEG[0]
  PIN W6BEG[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 90.940 0.450 91.340 ;
    END
  END W6BEG[10]
  PIN W6BEG[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 92.620 0.450 93.020 ;
    END
  END W6BEG[11]
  PIN W6BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 75.820 0.450 76.220 ;
    END
  END W6BEG[1]
  PIN W6BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 77.500 0.450 77.900 ;
    END
  END W6BEG[2]
  PIN W6BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 79.180 0.450 79.580 ;
    END
  END W6BEG[3]
  PIN W6BEG[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 80.860 0.450 81.260 ;
    END
  END W6BEG[4]
  PIN W6BEG[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 82.540 0.450 82.940 ;
    END
  END W6BEG[5]
  PIN W6BEG[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 84.220 0.450 84.620 ;
    END
  END W6BEG[6]
  PIN W6BEG[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 85.900 0.450 86.300 ;
    END
  END W6BEG[7]
  PIN W6BEG[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 87.580 0.450 87.980 ;
    END
  END W6BEG[8]
  PIN W6BEG[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 89.260 0.450 89.660 ;
    END
  END W6BEG[9]
  PIN W6END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 265.950 74.140 266.400 74.540 ;
    END
  END W6END[0]
  PIN W6END[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 265.950 90.940 266.400 91.340 ;
    END
  END W6END[10]
  PIN W6END[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 265.950 92.620 266.400 93.020 ;
    END
  END W6END[11]
  PIN W6END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 265.950 75.820 266.400 76.220 ;
    END
  END W6END[1]
  PIN W6END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 265.950 77.500 266.400 77.900 ;
    END
  END W6END[2]
  PIN W6END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 265.950 79.180 266.400 79.580 ;
    END
  END W6END[3]
  PIN W6END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 265.950 80.860 266.400 81.260 ;
    END
  END W6END[4]
  PIN W6END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 265.950 82.540 266.400 82.940 ;
    END
  END W6END[5]
  PIN W6END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 265.950 84.220 266.400 84.620 ;
    END
  END W6END[6]
  PIN W6END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 265.950 85.900 266.400 86.300 ;
    END
  END W6END[7]
  PIN W6END[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 265.950 87.580 266.400 87.980 ;
    END
  END W6END[8]
  PIN W6END[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 265.950 89.260 266.400 89.660 ;
    END
  END W6END[9]
  PIN WW4BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 47.260 0.450 47.660 ;
    END
  END WW4BEG[0]
  PIN WW4BEG[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 64.060 0.450 64.460 ;
    END
  END WW4BEG[10]
  PIN WW4BEG[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 65.740 0.450 66.140 ;
    END
  END WW4BEG[11]
  PIN WW4BEG[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 67.420 0.450 67.820 ;
    END
  END WW4BEG[12]
  PIN WW4BEG[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 69.100 0.450 69.500 ;
    END
  END WW4BEG[13]
  PIN WW4BEG[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 70.780 0.450 71.180 ;
    END
  END WW4BEG[14]
  PIN WW4BEG[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 72.460 0.450 72.860 ;
    END
  END WW4BEG[15]
  PIN WW4BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 48.940 0.450 49.340 ;
    END
  END WW4BEG[1]
  PIN WW4BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 50.620 0.450 51.020 ;
    END
  END WW4BEG[2]
  PIN WW4BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 52.300 0.450 52.700 ;
    END
  END WW4BEG[3]
  PIN WW4BEG[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 53.980 0.450 54.380 ;
    END
  END WW4BEG[4]
  PIN WW4BEG[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 55.660 0.450 56.060 ;
    END
  END WW4BEG[5]
  PIN WW4BEG[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 57.340 0.450 57.740 ;
    END
  END WW4BEG[6]
  PIN WW4BEG[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 59.020 0.450 59.420 ;
    END
  END WW4BEG[7]
  PIN WW4BEG[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 60.700 0.450 61.100 ;
    END
  END WW4BEG[8]
  PIN WW4BEG[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 62.380 0.450 62.780 ;
    END
  END WW4BEG[9]
  PIN WW4END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 265.950 47.260 266.400 47.660 ;
    END
  END WW4END[0]
  PIN WW4END[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 265.950 64.060 266.400 64.460 ;
    END
  END WW4END[10]
  PIN WW4END[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 265.950 65.740 266.400 66.140 ;
    END
  END WW4END[11]
  PIN WW4END[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 265.950 67.420 266.400 67.820 ;
    END
  END WW4END[12]
  PIN WW4END[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 265.950 69.100 266.400 69.500 ;
    END
  END WW4END[13]
  PIN WW4END[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 265.950 70.780 266.400 71.180 ;
    END
  END WW4END[14]
  PIN WW4END[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 265.950 72.460 266.400 72.860 ;
    END
  END WW4END[15]
  PIN WW4END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 265.950 48.940 266.400 49.340 ;
    END
  END WW4END[1]
  PIN WW4END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 265.950 50.620 266.400 51.020 ;
    END
  END WW4END[2]
  PIN WW4END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 265.950 52.300 266.400 52.700 ;
    END
  END WW4END[3]
  PIN WW4END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 265.950 53.980 266.400 54.380 ;
    END
  END WW4END[4]
  PIN WW4END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 265.950 55.660 266.400 56.060 ;
    END
  END WW4END[5]
  PIN WW4END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 265.950 57.340 266.400 57.740 ;
    END
  END WW4END[6]
  PIN WW4END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 265.950 59.020 266.400 59.420 ;
    END
  END WW4END[7]
  PIN WW4END[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 265.950 60.700 266.400 61.100 ;
    END
  END WW4END[8]
  PIN WW4END[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 265.950 62.380 266.400 62.780 ;
    END
  END WW4END[9]
  OBS
      LAYER GatPoly ;
        RECT 5.760 7.410 260.640 234.510 ;
      LAYER Metal1 ;
        RECT 5.760 7.340 260.640 234.580 ;
      LAYER Metal2 ;
        RECT 0.335 227.630 266.065 241.600 ;
        RECT 0.660 226.810 265.740 227.630 ;
        RECT 0.335 225.950 266.065 226.810 ;
        RECT 0.660 225.130 265.740 225.950 ;
        RECT 0.335 224.270 266.065 225.130 ;
        RECT 0.660 223.450 265.740 224.270 ;
        RECT 0.335 222.590 266.065 223.450 ;
        RECT 0.660 221.770 265.740 222.590 ;
        RECT 0.335 220.910 266.065 221.770 ;
        RECT 0.660 220.090 265.740 220.910 ;
        RECT 0.335 219.230 266.065 220.090 ;
        RECT 0.660 218.410 265.740 219.230 ;
        RECT 0.335 217.550 266.065 218.410 ;
        RECT 0.660 216.730 265.740 217.550 ;
        RECT 0.335 215.870 266.065 216.730 ;
        RECT 0.660 215.050 265.740 215.870 ;
        RECT 0.335 214.190 266.065 215.050 ;
        RECT 0.660 213.370 265.740 214.190 ;
        RECT 0.335 212.510 266.065 213.370 ;
        RECT 0.660 211.690 265.740 212.510 ;
        RECT 0.335 210.830 266.065 211.690 ;
        RECT 0.660 210.010 265.740 210.830 ;
        RECT 0.335 209.150 266.065 210.010 ;
        RECT 0.660 208.330 265.740 209.150 ;
        RECT 0.335 207.470 266.065 208.330 ;
        RECT 0.660 206.650 265.740 207.470 ;
        RECT 0.335 205.790 266.065 206.650 ;
        RECT 0.660 204.970 265.740 205.790 ;
        RECT 0.335 204.110 266.065 204.970 ;
        RECT 0.660 203.290 265.740 204.110 ;
        RECT 0.335 202.430 266.065 203.290 ;
        RECT 0.660 201.610 265.740 202.430 ;
        RECT 0.335 200.750 266.065 201.610 ;
        RECT 0.660 199.930 265.740 200.750 ;
        RECT 0.335 199.070 266.065 199.930 ;
        RECT 0.660 198.250 265.740 199.070 ;
        RECT 0.335 197.390 266.065 198.250 ;
        RECT 0.660 196.570 265.740 197.390 ;
        RECT 0.335 195.710 266.065 196.570 ;
        RECT 0.660 194.890 265.740 195.710 ;
        RECT 0.335 194.030 266.065 194.890 ;
        RECT 0.660 193.210 265.740 194.030 ;
        RECT 0.335 192.350 266.065 193.210 ;
        RECT 0.660 191.530 265.740 192.350 ;
        RECT 0.335 190.670 266.065 191.530 ;
        RECT 0.660 189.850 265.740 190.670 ;
        RECT 0.335 188.990 266.065 189.850 ;
        RECT 0.660 188.170 265.740 188.990 ;
        RECT 0.335 187.310 266.065 188.170 ;
        RECT 0.660 186.490 265.740 187.310 ;
        RECT 0.335 185.630 266.065 186.490 ;
        RECT 0.660 184.810 265.740 185.630 ;
        RECT 0.335 183.950 266.065 184.810 ;
        RECT 0.660 183.130 265.740 183.950 ;
        RECT 0.335 182.270 266.065 183.130 ;
        RECT 0.660 181.450 265.740 182.270 ;
        RECT 0.335 180.590 266.065 181.450 ;
        RECT 0.660 179.770 265.740 180.590 ;
        RECT 0.335 178.910 266.065 179.770 ;
        RECT 0.660 178.090 265.740 178.910 ;
        RECT 0.335 177.230 266.065 178.090 ;
        RECT 0.660 176.410 265.740 177.230 ;
        RECT 0.335 175.550 266.065 176.410 ;
        RECT 0.660 174.730 265.740 175.550 ;
        RECT 0.335 173.870 266.065 174.730 ;
        RECT 0.660 173.050 265.740 173.870 ;
        RECT 0.335 172.190 266.065 173.050 ;
        RECT 0.660 171.370 265.740 172.190 ;
        RECT 0.335 170.510 266.065 171.370 ;
        RECT 0.660 169.690 265.740 170.510 ;
        RECT 0.335 168.830 266.065 169.690 ;
        RECT 0.660 168.010 265.740 168.830 ;
        RECT 0.335 167.150 266.065 168.010 ;
        RECT 0.660 166.330 265.740 167.150 ;
        RECT 0.335 165.470 266.065 166.330 ;
        RECT 0.660 164.650 265.740 165.470 ;
        RECT 0.335 163.790 266.065 164.650 ;
        RECT 0.660 162.970 265.740 163.790 ;
        RECT 0.335 162.110 266.065 162.970 ;
        RECT 0.660 161.290 265.740 162.110 ;
        RECT 0.335 160.430 266.065 161.290 ;
        RECT 0.660 159.610 265.740 160.430 ;
        RECT 0.335 158.750 266.065 159.610 ;
        RECT 0.660 157.930 265.740 158.750 ;
        RECT 0.335 157.070 266.065 157.930 ;
        RECT 0.660 156.250 265.740 157.070 ;
        RECT 0.335 155.390 266.065 156.250 ;
        RECT 0.660 154.570 265.740 155.390 ;
        RECT 0.335 153.710 266.065 154.570 ;
        RECT 0.660 152.890 265.740 153.710 ;
        RECT 0.335 152.030 266.065 152.890 ;
        RECT 0.660 151.210 265.740 152.030 ;
        RECT 0.335 150.350 266.065 151.210 ;
        RECT 0.660 149.530 265.740 150.350 ;
        RECT 0.335 148.670 266.065 149.530 ;
        RECT 0.660 147.850 265.740 148.670 ;
        RECT 0.335 146.990 266.065 147.850 ;
        RECT 0.660 146.170 265.740 146.990 ;
        RECT 0.335 145.310 266.065 146.170 ;
        RECT 0.660 144.490 265.740 145.310 ;
        RECT 0.335 143.630 266.065 144.490 ;
        RECT 0.660 142.810 265.740 143.630 ;
        RECT 0.335 141.950 266.065 142.810 ;
        RECT 0.660 141.130 265.740 141.950 ;
        RECT 0.335 140.270 266.065 141.130 ;
        RECT 0.660 139.450 265.740 140.270 ;
        RECT 0.335 138.590 266.065 139.450 ;
        RECT 0.660 137.770 265.740 138.590 ;
        RECT 0.335 136.910 266.065 137.770 ;
        RECT 0.660 136.090 265.740 136.910 ;
        RECT 0.335 135.230 266.065 136.090 ;
        RECT 0.660 134.410 265.740 135.230 ;
        RECT 0.335 133.550 266.065 134.410 ;
        RECT 0.660 132.730 265.740 133.550 ;
        RECT 0.335 131.870 266.065 132.730 ;
        RECT 0.660 131.050 265.740 131.870 ;
        RECT 0.335 130.190 266.065 131.050 ;
        RECT 0.660 129.370 265.740 130.190 ;
        RECT 0.335 128.510 266.065 129.370 ;
        RECT 0.660 127.690 265.740 128.510 ;
        RECT 0.335 126.830 266.065 127.690 ;
        RECT 0.660 126.010 265.740 126.830 ;
        RECT 0.335 125.150 266.065 126.010 ;
        RECT 0.660 124.330 265.740 125.150 ;
        RECT 0.335 123.470 266.065 124.330 ;
        RECT 0.660 122.650 265.740 123.470 ;
        RECT 0.335 121.790 266.065 122.650 ;
        RECT 0.660 120.970 265.740 121.790 ;
        RECT 0.335 120.110 266.065 120.970 ;
        RECT 0.660 119.290 265.740 120.110 ;
        RECT 0.335 118.430 266.065 119.290 ;
        RECT 0.660 117.610 265.740 118.430 ;
        RECT 0.335 116.750 266.065 117.610 ;
        RECT 0.660 115.930 265.740 116.750 ;
        RECT 0.335 115.070 266.065 115.930 ;
        RECT 0.660 114.250 265.740 115.070 ;
        RECT 0.335 113.390 266.065 114.250 ;
        RECT 0.660 112.570 265.740 113.390 ;
        RECT 0.335 111.710 266.065 112.570 ;
        RECT 0.660 110.890 265.740 111.710 ;
        RECT 0.335 110.030 266.065 110.890 ;
        RECT 0.660 109.210 265.740 110.030 ;
        RECT 0.335 108.350 266.065 109.210 ;
        RECT 0.660 107.530 265.740 108.350 ;
        RECT 0.335 106.670 266.065 107.530 ;
        RECT 0.660 105.850 265.740 106.670 ;
        RECT 0.335 104.990 266.065 105.850 ;
        RECT 0.660 104.170 265.740 104.990 ;
        RECT 0.335 103.310 266.065 104.170 ;
        RECT 0.660 102.490 265.740 103.310 ;
        RECT 0.335 101.630 266.065 102.490 ;
        RECT 0.660 100.810 265.740 101.630 ;
        RECT 0.335 99.950 266.065 100.810 ;
        RECT 0.660 99.130 265.740 99.950 ;
        RECT 0.335 98.270 266.065 99.130 ;
        RECT 0.660 97.450 265.740 98.270 ;
        RECT 0.335 96.590 266.065 97.450 ;
        RECT 0.660 95.770 265.740 96.590 ;
        RECT 0.335 94.910 266.065 95.770 ;
        RECT 0.660 94.090 265.740 94.910 ;
        RECT 0.335 93.230 266.065 94.090 ;
        RECT 0.660 92.410 265.740 93.230 ;
        RECT 0.335 91.550 266.065 92.410 ;
        RECT 0.660 90.730 265.740 91.550 ;
        RECT 0.335 89.870 266.065 90.730 ;
        RECT 0.660 89.050 265.740 89.870 ;
        RECT 0.335 88.190 266.065 89.050 ;
        RECT 0.660 87.370 265.740 88.190 ;
        RECT 0.335 86.510 266.065 87.370 ;
        RECT 0.660 85.690 265.740 86.510 ;
        RECT 0.335 84.830 266.065 85.690 ;
        RECT 0.660 84.010 265.740 84.830 ;
        RECT 0.335 83.150 266.065 84.010 ;
        RECT 0.660 82.330 265.740 83.150 ;
        RECT 0.335 81.470 266.065 82.330 ;
        RECT 0.660 80.650 265.740 81.470 ;
        RECT 0.335 79.790 266.065 80.650 ;
        RECT 0.660 78.970 265.740 79.790 ;
        RECT 0.335 78.110 266.065 78.970 ;
        RECT 0.660 77.290 265.740 78.110 ;
        RECT 0.335 76.430 266.065 77.290 ;
        RECT 0.660 75.610 265.740 76.430 ;
        RECT 0.335 74.750 266.065 75.610 ;
        RECT 0.660 73.930 265.740 74.750 ;
        RECT 0.335 73.070 266.065 73.930 ;
        RECT 0.660 72.250 265.740 73.070 ;
        RECT 0.335 71.390 266.065 72.250 ;
        RECT 0.660 70.570 265.740 71.390 ;
        RECT 0.335 69.710 266.065 70.570 ;
        RECT 0.660 68.890 265.740 69.710 ;
        RECT 0.335 68.030 266.065 68.890 ;
        RECT 0.660 67.210 265.740 68.030 ;
        RECT 0.335 66.350 266.065 67.210 ;
        RECT 0.660 65.530 265.740 66.350 ;
        RECT 0.335 64.670 266.065 65.530 ;
        RECT 0.660 63.850 265.740 64.670 ;
        RECT 0.335 62.990 266.065 63.850 ;
        RECT 0.660 62.170 265.740 62.990 ;
        RECT 0.335 61.310 266.065 62.170 ;
        RECT 0.660 60.490 265.740 61.310 ;
        RECT 0.335 59.630 266.065 60.490 ;
        RECT 0.660 58.810 265.740 59.630 ;
        RECT 0.335 57.950 266.065 58.810 ;
        RECT 0.660 57.130 265.740 57.950 ;
        RECT 0.335 56.270 266.065 57.130 ;
        RECT 0.660 55.450 265.740 56.270 ;
        RECT 0.335 54.590 266.065 55.450 ;
        RECT 0.660 53.770 265.740 54.590 ;
        RECT 0.335 52.910 266.065 53.770 ;
        RECT 0.660 52.090 265.740 52.910 ;
        RECT 0.335 51.230 266.065 52.090 ;
        RECT 0.660 50.410 265.740 51.230 ;
        RECT 0.335 49.550 266.065 50.410 ;
        RECT 0.660 48.730 265.740 49.550 ;
        RECT 0.335 47.870 266.065 48.730 ;
        RECT 0.660 47.050 265.740 47.870 ;
        RECT 0.335 46.190 266.065 47.050 ;
        RECT 0.660 45.370 265.740 46.190 ;
        RECT 0.335 44.510 266.065 45.370 ;
        RECT 0.660 43.690 265.740 44.510 ;
        RECT 0.335 42.830 266.065 43.690 ;
        RECT 0.660 42.010 265.740 42.830 ;
        RECT 0.335 41.150 266.065 42.010 ;
        RECT 0.660 40.330 265.740 41.150 ;
        RECT 0.335 39.470 266.065 40.330 ;
        RECT 0.660 38.650 265.740 39.470 ;
        RECT 0.335 37.790 266.065 38.650 ;
        RECT 0.660 36.970 265.740 37.790 ;
        RECT 0.335 36.110 266.065 36.970 ;
        RECT 0.660 35.290 265.740 36.110 ;
        RECT 0.335 34.430 266.065 35.290 ;
        RECT 0.660 33.610 265.740 34.430 ;
        RECT 0.335 32.750 266.065 33.610 ;
        RECT 0.660 31.930 265.740 32.750 ;
        RECT 0.335 31.070 266.065 31.930 ;
        RECT 0.660 30.250 265.740 31.070 ;
        RECT 0.335 29.390 266.065 30.250 ;
        RECT 0.660 28.570 265.740 29.390 ;
        RECT 0.335 27.710 266.065 28.570 ;
        RECT 0.660 26.890 265.740 27.710 ;
        RECT 0.335 26.030 266.065 26.890 ;
        RECT 0.660 25.210 265.740 26.030 ;
        RECT 0.335 24.350 266.065 25.210 ;
        RECT 0.660 23.530 265.740 24.350 ;
        RECT 0.335 22.670 266.065 23.530 ;
        RECT 0.660 21.850 265.740 22.670 ;
        RECT 0.335 20.990 266.065 21.850 ;
        RECT 0.660 20.170 265.740 20.990 ;
        RECT 0.335 19.310 266.065 20.170 ;
        RECT 0.660 18.490 265.740 19.310 ;
        RECT 0.335 17.630 266.065 18.490 ;
        RECT 0.660 16.810 265.740 17.630 ;
        RECT 0.335 15.950 266.065 16.810 ;
        RECT 0.660 15.130 265.740 15.950 ;
        RECT 0.335 14.270 266.065 15.130 ;
        RECT 0.660 13.450 265.740 14.270 ;
        RECT 0.335 0.320 266.065 13.450 ;
      LAYER Metal3 ;
        RECT 0.380 241.310 13.510 241.820 ;
        RECT 14.330 241.310 15.430 241.820 ;
        RECT 16.250 241.310 17.350 241.820 ;
        RECT 18.170 241.310 19.270 241.820 ;
        RECT 20.090 241.310 21.190 241.820 ;
        RECT 22.010 241.310 23.110 241.820 ;
        RECT 23.930 241.310 25.030 241.820 ;
        RECT 25.850 241.310 26.950 241.820 ;
        RECT 27.770 241.310 28.870 241.820 ;
        RECT 29.690 241.310 30.790 241.820 ;
        RECT 31.610 241.310 32.710 241.820 ;
        RECT 33.530 241.310 34.630 241.820 ;
        RECT 35.450 241.310 36.550 241.820 ;
        RECT 37.370 241.310 38.470 241.820 ;
        RECT 39.290 241.310 40.390 241.820 ;
        RECT 41.210 241.310 42.310 241.820 ;
        RECT 43.130 241.310 44.230 241.820 ;
        RECT 45.050 241.310 46.150 241.820 ;
        RECT 46.970 241.310 48.070 241.820 ;
        RECT 48.890 241.310 49.990 241.820 ;
        RECT 50.810 241.310 51.910 241.820 ;
        RECT 52.730 241.310 53.830 241.820 ;
        RECT 54.650 241.310 55.750 241.820 ;
        RECT 56.570 241.310 57.670 241.820 ;
        RECT 58.490 241.310 59.590 241.820 ;
        RECT 60.410 241.310 61.510 241.820 ;
        RECT 62.330 241.310 63.430 241.820 ;
        RECT 64.250 241.310 65.350 241.820 ;
        RECT 66.170 241.310 67.270 241.820 ;
        RECT 68.090 241.310 69.190 241.820 ;
        RECT 70.010 241.310 71.110 241.820 ;
        RECT 71.930 241.310 73.030 241.820 ;
        RECT 73.850 241.310 74.950 241.820 ;
        RECT 75.770 241.310 76.870 241.820 ;
        RECT 77.690 241.310 78.790 241.820 ;
        RECT 79.610 241.310 80.710 241.820 ;
        RECT 81.530 241.310 82.630 241.820 ;
        RECT 83.450 241.310 84.550 241.820 ;
        RECT 85.370 241.310 86.470 241.820 ;
        RECT 87.290 241.310 88.390 241.820 ;
        RECT 89.210 241.310 90.310 241.820 ;
        RECT 91.130 241.310 92.230 241.820 ;
        RECT 93.050 241.310 94.150 241.820 ;
        RECT 94.970 241.310 96.070 241.820 ;
        RECT 96.890 241.310 97.990 241.820 ;
        RECT 98.810 241.310 99.910 241.820 ;
        RECT 100.730 241.310 101.830 241.820 ;
        RECT 102.650 241.310 103.750 241.820 ;
        RECT 104.570 241.310 105.670 241.820 ;
        RECT 106.490 241.310 107.590 241.820 ;
        RECT 108.410 241.310 109.510 241.820 ;
        RECT 110.330 241.310 111.430 241.820 ;
        RECT 112.250 241.310 113.350 241.820 ;
        RECT 114.170 241.310 115.270 241.820 ;
        RECT 116.090 241.310 117.190 241.820 ;
        RECT 118.010 241.310 119.110 241.820 ;
        RECT 119.930 241.310 121.030 241.820 ;
        RECT 121.850 241.310 122.950 241.820 ;
        RECT 123.770 241.310 124.870 241.820 ;
        RECT 125.690 241.310 126.790 241.820 ;
        RECT 127.610 241.310 128.710 241.820 ;
        RECT 129.530 241.310 130.630 241.820 ;
        RECT 131.450 241.310 132.550 241.820 ;
        RECT 133.370 241.310 134.470 241.820 ;
        RECT 135.290 241.310 136.390 241.820 ;
        RECT 137.210 241.310 138.310 241.820 ;
        RECT 139.130 241.310 140.230 241.820 ;
        RECT 141.050 241.310 142.150 241.820 ;
        RECT 142.970 241.310 144.070 241.820 ;
        RECT 144.890 241.310 145.990 241.820 ;
        RECT 146.810 241.310 147.910 241.820 ;
        RECT 148.730 241.310 149.830 241.820 ;
        RECT 150.650 241.310 151.750 241.820 ;
        RECT 152.570 241.310 153.670 241.820 ;
        RECT 154.490 241.310 155.590 241.820 ;
        RECT 156.410 241.310 157.510 241.820 ;
        RECT 158.330 241.310 159.430 241.820 ;
        RECT 160.250 241.310 161.350 241.820 ;
        RECT 162.170 241.310 163.270 241.820 ;
        RECT 164.090 241.310 165.190 241.820 ;
        RECT 166.010 241.310 167.110 241.820 ;
        RECT 167.930 241.310 169.030 241.820 ;
        RECT 169.850 241.310 170.950 241.820 ;
        RECT 171.770 241.310 172.870 241.820 ;
        RECT 173.690 241.310 174.790 241.820 ;
        RECT 175.610 241.310 176.710 241.820 ;
        RECT 177.530 241.310 178.630 241.820 ;
        RECT 179.450 241.310 180.550 241.820 ;
        RECT 181.370 241.310 182.470 241.820 ;
        RECT 183.290 241.310 184.390 241.820 ;
        RECT 185.210 241.310 186.310 241.820 ;
        RECT 187.130 241.310 188.230 241.820 ;
        RECT 189.050 241.310 190.150 241.820 ;
        RECT 190.970 241.310 192.070 241.820 ;
        RECT 192.890 241.310 193.990 241.820 ;
        RECT 194.810 241.310 195.910 241.820 ;
        RECT 196.730 241.310 197.830 241.820 ;
        RECT 198.650 241.310 199.750 241.820 ;
        RECT 200.570 241.310 201.670 241.820 ;
        RECT 202.490 241.310 203.590 241.820 ;
        RECT 204.410 241.310 205.510 241.820 ;
        RECT 206.330 241.310 207.430 241.820 ;
        RECT 208.250 241.310 209.350 241.820 ;
        RECT 210.170 241.310 211.270 241.820 ;
        RECT 212.090 241.310 213.190 241.820 ;
        RECT 214.010 241.310 215.110 241.820 ;
        RECT 215.930 241.310 217.030 241.820 ;
        RECT 217.850 241.310 218.950 241.820 ;
        RECT 219.770 241.310 220.870 241.820 ;
        RECT 221.690 241.310 222.790 241.820 ;
        RECT 223.610 241.310 224.710 241.820 ;
        RECT 225.530 241.310 226.630 241.820 ;
        RECT 227.450 241.310 228.550 241.820 ;
        RECT 229.370 241.310 230.470 241.820 ;
        RECT 231.290 241.310 232.390 241.820 ;
        RECT 233.210 241.310 234.310 241.820 ;
        RECT 235.130 241.310 236.230 241.820 ;
        RECT 237.050 241.310 238.150 241.820 ;
        RECT 238.970 241.310 240.070 241.820 ;
        RECT 240.890 241.310 241.990 241.820 ;
        RECT 242.810 241.310 243.910 241.820 ;
        RECT 244.730 241.310 245.830 241.820 ;
        RECT 246.650 241.310 247.750 241.820 ;
        RECT 248.570 241.310 249.670 241.820 ;
        RECT 250.490 241.310 251.590 241.820 ;
        RECT 252.410 241.310 266.020 241.820 ;
        RECT 0.380 0.610 266.020 241.310 ;
        RECT 0.380 0.100 13.510 0.610 ;
        RECT 14.330 0.100 15.430 0.610 ;
        RECT 16.250 0.100 17.350 0.610 ;
        RECT 18.170 0.100 19.270 0.610 ;
        RECT 20.090 0.100 21.190 0.610 ;
        RECT 22.010 0.100 23.110 0.610 ;
        RECT 23.930 0.100 25.030 0.610 ;
        RECT 25.850 0.100 26.950 0.610 ;
        RECT 27.770 0.100 28.870 0.610 ;
        RECT 29.690 0.100 30.790 0.610 ;
        RECT 31.610 0.100 32.710 0.610 ;
        RECT 33.530 0.100 34.630 0.610 ;
        RECT 35.450 0.100 36.550 0.610 ;
        RECT 37.370 0.100 38.470 0.610 ;
        RECT 39.290 0.100 40.390 0.610 ;
        RECT 41.210 0.100 42.310 0.610 ;
        RECT 43.130 0.100 44.230 0.610 ;
        RECT 45.050 0.100 46.150 0.610 ;
        RECT 46.970 0.100 48.070 0.610 ;
        RECT 48.890 0.100 49.990 0.610 ;
        RECT 50.810 0.100 51.910 0.610 ;
        RECT 52.730 0.100 53.830 0.610 ;
        RECT 54.650 0.100 55.750 0.610 ;
        RECT 56.570 0.100 57.670 0.610 ;
        RECT 58.490 0.100 59.590 0.610 ;
        RECT 60.410 0.100 61.510 0.610 ;
        RECT 62.330 0.100 63.430 0.610 ;
        RECT 64.250 0.100 65.350 0.610 ;
        RECT 66.170 0.100 67.270 0.610 ;
        RECT 68.090 0.100 69.190 0.610 ;
        RECT 70.010 0.100 71.110 0.610 ;
        RECT 71.930 0.100 73.030 0.610 ;
        RECT 73.850 0.100 74.950 0.610 ;
        RECT 75.770 0.100 76.870 0.610 ;
        RECT 77.690 0.100 78.790 0.610 ;
        RECT 79.610 0.100 80.710 0.610 ;
        RECT 81.530 0.100 82.630 0.610 ;
        RECT 83.450 0.100 84.550 0.610 ;
        RECT 85.370 0.100 86.470 0.610 ;
        RECT 87.290 0.100 88.390 0.610 ;
        RECT 89.210 0.100 90.310 0.610 ;
        RECT 91.130 0.100 92.230 0.610 ;
        RECT 93.050 0.100 94.150 0.610 ;
        RECT 94.970 0.100 96.070 0.610 ;
        RECT 96.890 0.100 97.990 0.610 ;
        RECT 98.810 0.100 99.910 0.610 ;
        RECT 100.730 0.100 101.830 0.610 ;
        RECT 102.650 0.100 103.750 0.610 ;
        RECT 104.570 0.100 105.670 0.610 ;
        RECT 106.490 0.100 107.590 0.610 ;
        RECT 108.410 0.100 109.510 0.610 ;
        RECT 110.330 0.100 111.430 0.610 ;
        RECT 112.250 0.100 113.350 0.610 ;
        RECT 114.170 0.100 115.270 0.610 ;
        RECT 116.090 0.100 117.190 0.610 ;
        RECT 118.010 0.100 119.110 0.610 ;
        RECT 119.930 0.100 121.030 0.610 ;
        RECT 121.850 0.100 122.950 0.610 ;
        RECT 123.770 0.100 124.870 0.610 ;
        RECT 125.690 0.100 126.790 0.610 ;
        RECT 127.610 0.100 128.710 0.610 ;
        RECT 129.530 0.100 130.630 0.610 ;
        RECT 131.450 0.100 132.550 0.610 ;
        RECT 133.370 0.100 134.470 0.610 ;
        RECT 135.290 0.100 136.390 0.610 ;
        RECT 137.210 0.100 138.310 0.610 ;
        RECT 139.130 0.100 140.230 0.610 ;
        RECT 141.050 0.100 142.150 0.610 ;
        RECT 142.970 0.100 144.070 0.610 ;
        RECT 144.890 0.100 145.990 0.610 ;
        RECT 146.810 0.100 147.910 0.610 ;
        RECT 148.730 0.100 149.830 0.610 ;
        RECT 150.650 0.100 151.750 0.610 ;
        RECT 152.570 0.100 153.670 0.610 ;
        RECT 154.490 0.100 155.590 0.610 ;
        RECT 156.410 0.100 157.510 0.610 ;
        RECT 158.330 0.100 159.430 0.610 ;
        RECT 160.250 0.100 161.350 0.610 ;
        RECT 162.170 0.100 163.270 0.610 ;
        RECT 164.090 0.100 165.190 0.610 ;
        RECT 166.010 0.100 167.110 0.610 ;
        RECT 167.930 0.100 169.030 0.610 ;
        RECT 169.850 0.100 170.950 0.610 ;
        RECT 171.770 0.100 172.870 0.610 ;
        RECT 173.690 0.100 174.790 0.610 ;
        RECT 175.610 0.100 176.710 0.610 ;
        RECT 177.530 0.100 178.630 0.610 ;
        RECT 179.450 0.100 180.550 0.610 ;
        RECT 181.370 0.100 182.470 0.610 ;
        RECT 183.290 0.100 184.390 0.610 ;
        RECT 185.210 0.100 186.310 0.610 ;
        RECT 187.130 0.100 188.230 0.610 ;
        RECT 189.050 0.100 190.150 0.610 ;
        RECT 190.970 0.100 192.070 0.610 ;
        RECT 192.890 0.100 193.990 0.610 ;
        RECT 194.810 0.100 195.910 0.610 ;
        RECT 196.730 0.100 197.830 0.610 ;
        RECT 198.650 0.100 199.750 0.610 ;
        RECT 200.570 0.100 201.670 0.610 ;
        RECT 202.490 0.100 203.590 0.610 ;
        RECT 204.410 0.100 205.510 0.610 ;
        RECT 206.330 0.100 207.430 0.610 ;
        RECT 208.250 0.100 209.350 0.610 ;
        RECT 210.170 0.100 211.270 0.610 ;
        RECT 212.090 0.100 213.190 0.610 ;
        RECT 214.010 0.100 215.110 0.610 ;
        RECT 215.930 0.100 217.030 0.610 ;
        RECT 217.850 0.100 218.950 0.610 ;
        RECT 219.770 0.100 220.870 0.610 ;
        RECT 221.690 0.100 222.790 0.610 ;
        RECT 223.610 0.100 224.710 0.610 ;
        RECT 225.530 0.100 226.630 0.610 ;
        RECT 227.450 0.100 228.550 0.610 ;
        RECT 229.370 0.100 230.470 0.610 ;
        RECT 231.290 0.100 232.390 0.610 ;
        RECT 233.210 0.100 234.310 0.610 ;
        RECT 235.130 0.100 236.230 0.610 ;
        RECT 237.050 0.100 238.150 0.610 ;
        RECT 238.970 0.100 240.070 0.610 ;
        RECT 240.890 0.100 241.990 0.610 ;
        RECT 242.810 0.100 243.910 0.610 ;
        RECT 244.730 0.100 245.830 0.610 ;
        RECT 246.650 0.100 247.750 0.610 ;
        RECT 248.570 0.100 249.670 0.610 ;
        RECT 250.490 0.100 251.590 0.610 ;
        RECT 252.410 0.100 266.020 0.610 ;
      LAYER Metal4 ;
        RECT 0.335 0.320 266.065 241.600 ;
      LAYER Metal5 ;
        RECT 0.380 1.115 18.050 232.405 ;
        RECT 20.670 1.115 24.250 232.405 ;
        RECT 26.870 1.115 93.650 232.405 ;
        RECT 96.270 1.115 99.850 232.405 ;
        RECT 102.470 1.115 169.250 232.405 ;
        RECT 171.870 1.115 175.450 232.405 ;
        RECT 178.070 1.115 244.850 232.405 ;
        RECT 247.470 1.115 251.050 232.405 ;
        RECT 253.670 1.115 266.020 232.405 ;
  END
END RegFile
END LIBRARY

