magic
tech ihp-sg13g2
magscale 1 2
timestamp 1743692007
<< metal1 >>
rect 1152 10604 45216 10628
rect 1152 10564 4928 10604
rect 4968 10564 5010 10604
rect 5050 10564 5092 10604
rect 5132 10564 5174 10604
rect 5214 10564 5256 10604
rect 5296 10564 20048 10604
rect 20088 10564 20130 10604
rect 20170 10564 20212 10604
rect 20252 10564 20294 10604
rect 20334 10564 20376 10604
rect 20416 10564 35168 10604
rect 35208 10564 35250 10604
rect 35290 10564 35332 10604
rect 35372 10564 35414 10604
rect 35454 10564 35496 10604
rect 35536 10564 45216 10604
rect 1152 10540 45216 10564
rect 2043 10436 2085 10445
rect 2043 10396 2044 10436
rect 2084 10396 2085 10436
rect 2043 10387 2085 10396
rect 4155 10436 4197 10445
rect 4155 10396 4156 10436
rect 4196 10396 4197 10436
rect 4155 10387 4197 10396
rect 6267 10436 6309 10445
rect 6267 10396 6268 10436
rect 6308 10396 6309 10436
rect 6267 10387 6309 10396
rect 8379 10436 8421 10445
rect 8379 10396 8380 10436
rect 8420 10396 8421 10436
rect 8379 10387 8421 10396
rect 10491 10436 10533 10445
rect 10491 10396 10492 10436
rect 10532 10396 10533 10436
rect 10491 10387 10533 10396
rect 12603 10436 12645 10445
rect 12603 10396 12604 10436
rect 12644 10396 12645 10436
rect 12603 10387 12645 10396
rect 14715 10436 14757 10445
rect 14715 10396 14716 10436
rect 14756 10396 14757 10436
rect 14715 10387 14757 10396
rect 16827 10436 16869 10445
rect 16827 10396 16828 10436
rect 16868 10396 16869 10436
rect 16827 10387 16869 10396
rect 18939 10436 18981 10445
rect 18939 10396 18940 10436
rect 18980 10396 18981 10436
rect 18939 10387 18981 10396
rect 21051 10436 21093 10445
rect 21051 10396 21052 10436
rect 21092 10396 21093 10436
rect 21051 10387 21093 10396
rect 23163 10436 23205 10445
rect 23163 10396 23164 10436
rect 23204 10396 23205 10436
rect 23163 10387 23205 10396
rect 25275 10436 25317 10445
rect 25275 10396 25276 10436
rect 25316 10396 25317 10436
rect 25275 10387 25317 10396
rect 27387 10436 27429 10445
rect 27387 10396 27388 10436
rect 27428 10396 27429 10436
rect 27387 10387 27429 10396
rect 29499 10436 29541 10445
rect 29499 10396 29500 10436
rect 29540 10396 29541 10436
rect 29499 10387 29541 10396
rect 31611 10436 31653 10445
rect 31611 10396 31612 10436
rect 31652 10396 31653 10436
rect 31611 10387 31653 10396
rect 33723 10436 33765 10445
rect 33723 10396 33724 10436
rect 33764 10396 33765 10436
rect 33723 10387 33765 10396
rect 35835 10436 35877 10445
rect 35835 10396 35836 10436
rect 35876 10396 35877 10436
rect 35835 10387 35877 10396
rect 37947 10436 37989 10445
rect 37947 10396 37948 10436
rect 37988 10396 37989 10436
rect 37947 10387 37989 10396
rect 40059 10436 40101 10445
rect 40059 10396 40060 10436
rect 40100 10396 40101 10436
rect 40059 10387 40101 10396
rect 42171 10436 42213 10445
rect 42171 10396 42172 10436
rect 42212 10396 42213 10436
rect 42171 10387 42213 10396
rect 43419 10436 43461 10445
rect 43419 10396 43420 10436
rect 43460 10396 43461 10436
rect 43419 10387 43461 10396
rect 44283 10436 44325 10445
rect 44283 10396 44284 10436
rect 44324 10396 44325 10436
rect 44283 10387 44325 10396
rect 2283 10184 2325 10193
rect 2283 10144 2284 10184
rect 2324 10144 2325 10184
rect 2283 10135 2325 10144
rect 4395 10184 4437 10193
rect 4395 10144 4396 10184
rect 4436 10144 4437 10184
rect 4395 10135 4437 10144
rect 6507 10184 6549 10193
rect 6507 10144 6508 10184
rect 6548 10144 6549 10184
rect 6507 10135 6549 10144
rect 8619 10184 8661 10193
rect 8619 10144 8620 10184
rect 8660 10144 8661 10184
rect 8619 10135 8661 10144
rect 10731 10184 10773 10193
rect 10731 10144 10732 10184
rect 10772 10144 10773 10184
rect 10731 10135 10773 10144
rect 12843 10184 12885 10193
rect 12843 10144 12844 10184
rect 12884 10144 12885 10184
rect 12843 10135 12885 10144
rect 14955 10184 14997 10193
rect 14955 10144 14956 10184
rect 14996 10144 14997 10184
rect 14955 10135 14997 10144
rect 17067 10184 17109 10193
rect 17067 10144 17068 10184
rect 17108 10144 17109 10184
rect 17067 10135 17109 10144
rect 19179 10184 19221 10193
rect 19179 10144 19180 10184
rect 19220 10144 19221 10184
rect 19179 10135 19221 10144
rect 21291 10184 21333 10193
rect 21291 10144 21292 10184
rect 21332 10144 21333 10184
rect 21291 10135 21333 10144
rect 23451 10184 23493 10193
rect 23451 10144 23452 10184
rect 23492 10144 23493 10184
rect 23451 10135 23493 10144
rect 25515 10184 25557 10193
rect 25515 10144 25516 10184
rect 25556 10144 25557 10184
rect 25515 10135 25557 10144
rect 27627 10184 27669 10193
rect 27627 10144 27628 10184
rect 27668 10144 27669 10184
rect 27627 10135 27669 10144
rect 29739 10184 29781 10193
rect 29739 10144 29740 10184
rect 29780 10144 29781 10184
rect 29739 10135 29781 10144
rect 31851 10184 31893 10193
rect 31851 10144 31852 10184
rect 31892 10144 31893 10184
rect 31851 10135 31893 10144
rect 33963 10184 34005 10193
rect 33963 10144 33964 10184
rect 34004 10144 34005 10184
rect 33963 10135 34005 10144
rect 36075 10184 36117 10193
rect 36075 10144 36076 10184
rect 36116 10144 36117 10184
rect 36075 10135 36117 10144
rect 38187 10184 38229 10193
rect 38187 10144 38188 10184
rect 38228 10144 38229 10184
rect 38187 10135 38229 10144
rect 40299 10184 40341 10193
rect 40299 10144 40300 10184
rect 40340 10144 40341 10184
rect 40299 10135 40341 10144
rect 42411 10184 42453 10193
rect 42411 10144 42412 10184
rect 42452 10144 42453 10184
rect 42411 10135 42453 10144
rect 43179 10184 43221 10193
rect 43179 10144 43180 10184
rect 43220 10144 43221 10184
rect 43179 10135 43221 10144
rect 43563 10184 43605 10193
rect 43563 10144 43564 10184
rect 43604 10144 43605 10184
rect 43563 10135 43605 10144
rect 43947 10184 43989 10193
rect 43947 10144 43948 10184
rect 43988 10144 43989 10184
rect 43947 10135 43989 10144
rect 44523 10184 44565 10193
rect 44523 10144 44524 10184
rect 44564 10144 44565 10184
rect 44523 10135 44565 10144
rect 44907 10184 44949 10193
rect 44907 10144 44908 10184
rect 44948 10144 44949 10184
rect 44907 10135 44949 10144
rect 43803 10100 43845 10109
rect 43803 10060 43804 10100
rect 43844 10060 43845 10100
rect 43803 10051 43845 10060
rect 44187 10016 44229 10025
rect 44187 9976 44188 10016
rect 44228 9976 44229 10016
rect 44187 9967 44229 9976
rect 45147 10016 45189 10025
rect 45147 9976 45148 10016
rect 45188 9976 45189 10016
rect 45147 9967 45189 9976
rect 1152 9848 45216 9872
rect 1152 9808 3688 9848
rect 3728 9808 3770 9848
rect 3810 9808 3852 9848
rect 3892 9808 3934 9848
rect 3974 9808 4016 9848
rect 4056 9808 18808 9848
rect 18848 9808 18890 9848
rect 18930 9808 18972 9848
rect 19012 9808 19054 9848
rect 19094 9808 19136 9848
rect 19176 9808 33928 9848
rect 33968 9808 34010 9848
rect 34050 9808 34092 9848
rect 34132 9808 34174 9848
rect 34214 9808 34256 9848
rect 34296 9808 45216 9848
rect 1152 9784 45216 9808
rect 44379 9680 44421 9689
rect 44379 9640 44380 9680
rect 44420 9640 44421 9680
rect 44379 9631 44421 9640
rect 43995 9596 44037 9605
rect 43995 9556 43996 9596
rect 44036 9556 44037 9596
rect 43995 9547 44037 9556
rect 43755 9512 43797 9521
rect 43755 9472 43756 9512
rect 43796 9472 43797 9512
rect 43755 9463 43797 9472
rect 44139 9512 44181 9521
rect 44139 9472 44140 9512
rect 44180 9472 44181 9512
rect 44139 9463 44181 9472
rect 44523 9512 44565 9521
rect 44523 9472 44524 9512
rect 44564 9472 44565 9512
rect 44523 9463 44565 9472
rect 44907 9512 44949 9521
rect 44907 9472 44908 9512
rect 44948 9472 44949 9512
rect 44907 9463 44949 9472
rect 44763 9260 44805 9269
rect 44763 9220 44764 9260
rect 44804 9220 44805 9260
rect 44763 9211 44805 9220
rect 45147 9260 45189 9269
rect 45147 9220 45148 9260
rect 45188 9220 45189 9260
rect 45147 9211 45189 9220
rect 1152 9092 45216 9116
rect 1152 9052 4928 9092
rect 4968 9052 5010 9092
rect 5050 9052 5092 9092
rect 5132 9052 5174 9092
rect 5214 9052 5256 9092
rect 5296 9052 20048 9092
rect 20088 9052 20130 9092
rect 20170 9052 20212 9092
rect 20252 9052 20294 9092
rect 20334 9052 20376 9092
rect 20416 9052 35168 9092
rect 35208 9052 35250 9092
rect 35290 9052 35332 9092
rect 35372 9052 35414 9092
rect 35454 9052 35496 9092
rect 35536 9052 45216 9092
rect 1152 9028 45216 9052
rect 6171 8924 6213 8933
rect 6171 8884 6172 8924
rect 6212 8884 6213 8924
rect 6171 8875 6213 8884
rect 8571 8924 8613 8933
rect 8571 8884 8572 8924
rect 8612 8884 8613 8924
rect 8571 8875 8613 8884
rect 13083 8924 13125 8933
rect 13083 8884 13084 8924
rect 13124 8884 13125 8924
rect 13083 8875 13125 8884
rect 18747 8924 18789 8933
rect 18747 8884 18748 8924
rect 18788 8884 18789 8924
rect 18747 8875 18789 8884
rect 21531 8924 21573 8933
rect 21531 8884 21532 8924
rect 21572 8884 21573 8924
rect 21531 8875 21573 8884
rect 22299 8924 22341 8933
rect 22299 8884 22300 8924
rect 22340 8884 22341 8924
rect 22299 8875 22341 8884
rect 23067 8924 23109 8933
rect 23067 8884 23068 8924
rect 23108 8884 23109 8924
rect 23067 8875 23109 8884
rect 23451 8924 23493 8933
rect 23451 8884 23452 8924
rect 23492 8884 23493 8924
rect 23451 8875 23493 8884
rect 23835 8924 23877 8933
rect 23835 8884 23836 8924
rect 23876 8884 23877 8924
rect 23835 8875 23877 8884
rect 25851 8924 25893 8933
rect 25851 8884 25852 8924
rect 25892 8884 25893 8924
rect 25851 8875 25893 8884
rect 26907 8924 26949 8933
rect 26907 8884 26908 8924
rect 26948 8884 26949 8924
rect 26907 8875 26949 8884
rect 27291 8924 27333 8933
rect 27291 8884 27292 8924
rect 27332 8884 27333 8924
rect 27291 8875 27333 8884
rect 28059 8924 28101 8933
rect 28059 8884 28060 8924
rect 28100 8884 28101 8924
rect 28059 8875 28101 8884
rect 28731 8924 28773 8933
rect 28731 8884 28732 8924
rect 28772 8884 28773 8924
rect 28731 8875 28773 8884
rect 29115 8924 29157 8933
rect 29115 8884 29116 8924
rect 29156 8884 29157 8924
rect 29115 8875 29157 8884
rect 24411 8840 24453 8849
rect 24411 8800 24412 8840
rect 24452 8800 24453 8840
rect 24411 8791 24453 8800
rect 27963 8840 28005 8849
rect 27963 8800 27964 8840
rect 28004 8800 28005 8840
rect 27963 8791 28005 8800
rect 31227 8840 31269 8849
rect 31227 8800 31228 8840
rect 31268 8800 31269 8840
rect 31227 8791 31269 8800
rect 6411 8672 6453 8681
rect 6411 8632 6412 8672
rect 6452 8632 6453 8672
rect 6411 8623 6453 8632
rect 6651 8672 6693 8681
rect 6651 8632 6652 8672
rect 6692 8632 6693 8672
rect 6651 8623 6693 8632
rect 6891 8672 6933 8681
rect 6891 8632 6892 8672
rect 6932 8632 6933 8672
rect 6891 8623 6933 8632
rect 7467 8672 7509 8681
rect 7467 8632 7468 8672
rect 7508 8632 7509 8672
rect 7467 8623 7509 8632
rect 7707 8672 7749 8681
rect 7707 8632 7708 8672
rect 7748 8632 7749 8672
rect 7707 8623 7749 8632
rect 8811 8672 8853 8681
rect 8811 8632 8812 8672
rect 8852 8632 8853 8672
rect 8811 8623 8853 8632
rect 13323 8672 13365 8681
rect 13323 8632 13324 8672
rect 13364 8632 13365 8672
rect 13323 8623 13365 8632
rect 18987 8672 19029 8681
rect 18987 8632 18988 8672
rect 19028 8632 19029 8672
rect 18987 8623 19029 8632
rect 21291 8672 21333 8681
rect 21291 8632 21292 8672
rect 21332 8632 21333 8672
rect 21291 8623 21333 8632
rect 21675 8672 21717 8681
rect 21675 8632 21676 8672
rect 21716 8632 21717 8672
rect 21675 8623 21717 8632
rect 22059 8672 22101 8681
rect 22059 8632 22060 8672
rect 22100 8632 22101 8672
rect 22059 8623 22101 8632
rect 22443 8672 22485 8681
rect 22443 8632 22444 8672
rect 22484 8632 22485 8672
rect 22443 8623 22485 8632
rect 22858 8672 22916 8673
rect 22858 8632 22867 8672
rect 22907 8632 22916 8672
rect 22858 8631 22916 8632
rect 23211 8672 23253 8681
rect 23211 8632 23212 8672
rect 23252 8632 23253 8672
rect 23211 8623 23253 8632
rect 23595 8672 23637 8681
rect 23595 8632 23596 8672
rect 23636 8632 23637 8672
rect 23595 8623 23637 8632
rect 24171 8672 24213 8681
rect 24171 8632 24172 8672
rect 24212 8632 24213 8672
rect 24171 8623 24213 8632
rect 26091 8672 26133 8681
rect 26091 8632 26092 8672
rect 26132 8632 26133 8672
rect 26091 8623 26133 8632
rect 27147 8672 27189 8681
rect 27147 8632 27148 8672
rect 27188 8632 27189 8672
rect 27147 8623 27189 8632
rect 27531 8672 27573 8681
rect 27531 8632 27532 8672
rect 27572 8632 27573 8672
rect 27531 8623 27573 8632
rect 27723 8672 27765 8681
rect 27723 8632 27724 8672
rect 27764 8632 27765 8672
rect 27723 8623 27765 8632
rect 28299 8672 28341 8681
rect 28299 8632 28300 8672
rect 28340 8632 28341 8672
rect 28299 8623 28341 8632
rect 28491 8672 28533 8681
rect 28491 8632 28492 8672
rect 28532 8632 28533 8672
rect 28491 8623 28533 8632
rect 29355 8672 29397 8681
rect 29355 8632 29356 8672
rect 29396 8632 29397 8672
rect 29355 8623 29397 8632
rect 31467 8672 31509 8681
rect 31467 8632 31468 8672
rect 31508 8632 31509 8672
rect 31467 8623 31509 8632
rect 31851 8672 31893 8681
rect 31851 8632 31852 8672
rect 31892 8632 31893 8672
rect 31851 8623 31893 8632
rect 44523 8672 44565 8681
rect 44523 8632 44524 8672
rect 44564 8632 44565 8672
rect 44523 8623 44565 8632
rect 44907 8672 44949 8681
rect 44907 8632 44908 8672
rect 44948 8632 44949 8672
rect 44907 8623 44949 8632
rect 45147 8672 45189 8681
rect 45147 8632 45148 8672
rect 45188 8632 45189 8672
rect 45147 8623 45189 8632
rect 22683 8588 22725 8597
rect 22683 8548 22684 8588
rect 22724 8548 22725 8588
rect 22683 8539 22725 8548
rect 31611 8588 31653 8597
rect 31611 8548 31612 8588
rect 31652 8548 31653 8588
rect 31611 8539 31653 8548
rect 44763 8588 44805 8597
rect 44763 8548 44764 8588
rect 44804 8548 44805 8588
rect 44763 8539 44805 8548
rect 21915 8504 21957 8513
rect 21915 8464 21916 8504
rect 21956 8464 21957 8504
rect 21915 8455 21957 8464
rect 1152 8336 45216 8360
rect 1152 8296 3688 8336
rect 3728 8296 3770 8336
rect 3810 8296 3852 8336
rect 3892 8296 3934 8336
rect 3974 8296 4016 8336
rect 4056 8296 18808 8336
rect 18848 8296 18890 8336
rect 18930 8296 18972 8336
rect 19012 8296 19054 8336
rect 19094 8296 19136 8336
rect 19176 8296 33928 8336
rect 33968 8296 34010 8336
rect 34050 8296 34092 8336
rect 34132 8296 34174 8336
rect 34214 8296 34256 8336
rect 34296 8296 45216 8336
rect 1152 8272 45216 8296
rect 16827 8168 16869 8177
rect 16827 8128 16828 8168
rect 16868 8128 16869 8168
rect 16827 8119 16869 8128
rect 17979 8168 18021 8177
rect 17979 8128 17980 8168
rect 18020 8128 18021 8168
rect 17979 8119 18021 8128
rect 28059 8168 28101 8177
rect 28059 8128 28060 8168
rect 28100 8128 28101 8168
rect 28059 8119 28101 8128
rect 28827 8168 28869 8177
rect 28827 8128 28828 8168
rect 28868 8128 28869 8168
rect 28827 8119 28869 8128
rect 24987 8084 25029 8093
rect 24987 8044 24988 8084
rect 25028 8044 25029 8084
rect 24987 8035 25029 8044
rect 16203 8000 16245 8009
rect 16203 7960 16204 8000
rect 16244 7960 16245 8000
rect 16203 7951 16245 7960
rect 16587 8000 16629 8009
rect 16587 7960 16588 8000
rect 16628 7960 16629 8000
rect 16587 7951 16629 7960
rect 16971 8000 17013 8009
rect 16971 7960 16972 8000
rect 17012 7960 17013 8000
rect 16971 7951 17013 7960
rect 17355 8000 17397 8009
rect 17355 7960 17356 8000
rect 17396 7960 17397 8000
rect 17355 7951 17397 7960
rect 17739 8000 17781 8009
rect 17739 7960 17740 8000
rect 17780 7960 17781 8000
rect 17739 7951 17781 7960
rect 18411 8000 18453 8009
rect 18411 7960 18412 8000
rect 18452 7960 18453 8000
rect 18411 7951 18453 7960
rect 18795 8000 18837 8009
rect 18795 7960 18796 8000
rect 18836 7960 18837 8000
rect 18795 7951 18837 7960
rect 24747 8000 24789 8009
rect 24747 7960 24748 8000
rect 24788 7960 24789 8000
rect 24747 7951 24789 7960
rect 25419 8000 25461 8009
rect 25419 7960 25420 8000
rect 25460 7960 25461 8000
rect 25419 7951 25461 7960
rect 26283 8000 26325 8009
rect 26283 7960 26284 8000
rect 26324 7960 26325 8000
rect 26283 7951 26325 7960
rect 27819 8000 27861 8009
rect 27819 7960 27820 8000
rect 27860 7960 27861 8000
rect 27819 7951 27861 7960
rect 28587 8000 28629 8009
rect 28587 7960 28588 8000
rect 28628 7960 28629 8000
rect 28587 7951 28629 7960
rect 44523 8000 44565 8009
rect 44523 7960 44524 8000
rect 44564 7960 44565 8000
rect 44523 7951 44565 7960
rect 44907 8000 44949 8009
rect 44907 7960 44908 8000
rect 44948 7960 44949 8000
rect 44907 7951 44949 7960
rect 26523 7832 26565 7841
rect 26523 7792 26524 7832
rect 26564 7792 26565 7832
rect 26523 7783 26565 7792
rect 44763 7832 44805 7841
rect 44763 7792 44764 7832
rect 44804 7792 44805 7832
rect 44763 7783 44805 7792
rect 16443 7748 16485 7757
rect 16443 7708 16444 7748
rect 16484 7708 16485 7748
rect 16443 7699 16485 7708
rect 17211 7748 17253 7757
rect 17211 7708 17212 7748
rect 17252 7708 17253 7748
rect 17211 7699 17253 7708
rect 17595 7748 17637 7757
rect 17595 7708 17596 7748
rect 17636 7708 17637 7748
rect 17595 7699 17637 7708
rect 18651 7748 18693 7757
rect 18651 7708 18652 7748
rect 18692 7708 18693 7748
rect 18651 7699 18693 7708
rect 19035 7748 19077 7757
rect 19035 7708 19036 7748
rect 19076 7708 19077 7748
rect 19035 7699 19077 7708
rect 25659 7748 25701 7757
rect 25659 7708 25660 7748
rect 25700 7708 25701 7748
rect 25659 7699 25701 7708
rect 45147 7748 45189 7757
rect 45147 7708 45148 7748
rect 45188 7708 45189 7748
rect 45147 7699 45189 7708
rect 1152 7580 45216 7604
rect 1152 7540 4928 7580
rect 4968 7540 5010 7580
rect 5050 7540 5092 7580
rect 5132 7540 5174 7580
rect 5214 7540 5256 7580
rect 5296 7540 20048 7580
rect 20088 7540 20130 7580
rect 20170 7540 20212 7580
rect 20252 7540 20294 7580
rect 20334 7540 20376 7580
rect 20416 7540 35168 7580
rect 35208 7540 35250 7580
rect 35290 7540 35332 7580
rect 35372 7540 35414 7580
rect 35454 7540 35496 7580
rect 35536 7540 45216 7580
rect 1152 7516 45216 7540
rect 12459 7160 12501 7169
rect 12459 7120 12460 7160
rect 12500 7120 12501 7160
rect 12459 7111 12501 7120
rect 13899 7160 13941 7169
rect 13899 7120 13900 7160
rect 13940 7120 13941 7160
rect 13899 7111 13941 7120
rect 14955 7160 14997 7169
rect 14955 7120 14956 7160
rect 14996 7120 14997 7160
rect 14955 7111 14997 7120
rect 16107 7160 16149 7169
rect 16107 7120 16108 7160
rect 16148 7120 16149 7160
rect 16107 7111 16149 7120
rect 16875 7160 16917 7169
rect 16875 7120 16876 7160
rect 16916 7120 16917 7160
rect 16875 7111 16917 7120
rect 17355 7160 17397 7169
rect 17355 7120 17356 7160
rect 17396 7120 17397 7160
rect 17355 7111 17397 7120
rect 17739 7160 17781 7169
rect 17739 7120 17740 7160
rect 17780 7120 17781 7160
rect 17739 7111 17781 7120
rect 18123 7160 18165 7169
rect 18123 7120 18124 7160
rect 18164 7120 18165 7160
rect 18123 7111 18165 7120
rect 18507 7160 18549 7169
rect 18507 7120 18508 7160
rect 18548 7120 18549 7160
rect 18507 7111 18549 7120
rect 18891 7160 18933 7169
rect 18891 7120 18892 7160
rect 18932 7120 18933 7160
rect 18891 7111 18933 7120
rect 19275 7160 19317 7169
rect 19275 7120 19276 7160
rect 19316 7120 19317 7160
rect 19275 7111 19317 7120
rect 19659 7160 19701 7169
rect 19659 7120 19660 7160
rect 19700 7120 19701 7160
rect 19659 7111 19701 7120
rect 20043 7160 20085 7169
rect 20043 7120 20044 7160
rect 20084 7120 20085 7160
rect 20043 7111 20085 7120
rect 20427 7160 20469 7169
rect 20427 7120 20428 7160
rect 20468 7120 20469 7160
rect 20427 7111 20469 7120
rect 20811 7160 20853 7169
rect 20811 7120 20812 7160
rect 20852 7120 20853 7160
rect 20811 7111 20853 7120
rect 21051 7160 21093 7169
rect 21051 7120 21052 7160
rect 21092 7120 21093 7160
rect 21051 7111 21093 7120
rect 21195 7160 21237 7169
rect 21195 7120 21196 7160
rect 21236 7120 21237 7160
rect 21195 7111 21237 7120
rect 44523 7160 44565 7169
rect 44523 7120 44524 7160
rect 44564 7120 44565 7160
rect 44523 7111 44565 7120
rect 44907 7160 44949 7169
rect 44907 7120 44908 7160
rect 44948 7120 44949 7160
rect 44907 7111 44949 7120
rect 45147 7160 45189 7169
rect 45147 7120 45148 7160
rect 45188 7120 45189 7160
rect 45147 7111 45189 7120
rect 18747 7076 18789 7085
rect 18747 7036 18748 7076
rect 18788 7036 18789 7076
rect 18747 7027 18789 7036
rect 20667 7076 20709 7085
rect 20667 7036 20668 7076
rect 20708 7036 20709 7076
rect 20667 7027 20709 7036
rect 12699 6992 12741 7001
rect 12699 6952 12700 6992
rect 12740 6952 12741 6992
rect 12699 6943 12741 6952
rect 14139 6992 14181 7001
rect 14139 6952 14140 6992
rect 14180 6952 14181 6992
rect 14139 6943 14181 6952
rect 15195 6992 15237 7001
rect 15195 6952 15196 6992
rect 15236 6952 15237 6992
rect 15195 6943 15237 6952
rect 16347 6992 16389 7001
rect 16347 6952 16348 6992
rect 16388 6952 16389 6992
rect 16347 6943 16389 6952
rect 17115 6992 17157 7001
rect 17115 6952 17116 6992
rect 17156 6952 17157 6992
rect 17115 6943 17157 6952
rect 17595 6992 17637 7001
rect 17595 6952 17596 6992
rect 17636 6952 17637 6992
rect 17595 6943 17637 6952
rect 17979 6992 18021 7001
rect 17979 6952 17980 6992
rect 18020 6952 18021 6992
rect 17979 6943 18021 6952
rect 18363 6992 18405 7001
rect 18363 6952 18364 6992
rect 18404 6952 18405 6992
rect 18363 6943 18405 6952
rect 19131 6992 19173 7001
rect 19131 6952 19132 6992
rect 19172 6952 19173 6992
rect 19131 6943 19173 6952
rect 19515 6992 19557 7001
rect 19515 6952 19516 6992
rect 19556 6952 19557 6992
rect 19515 6943 19557 6952
rect 19899 6992 19941 7001
rect 19899 6952 19900 6992
rect 19940 6952 19941 6992
rect 19899 6943 19941 6952
rect 20283 6992 20325 7001
rect 20283 6952 20284 6992
rect 20324 6952 20325 6992
rect 20283 6943 20325 6952
rect 21435 6992 21477 7001
rect 21435 6952 21436 6992
rect 21476 6952 21477 6992
rect 21435 6943 21477 6952
rect 44763 6992 44805 7001
rect 44763 6952 44764 6992
rect 44804 6952 44805 6992
rect 44763 6943 44805 6952
rect 1152 6824 45216 6848
rect 1152 6784 3688 6824
rect 3728 6784 3770 6824
rect 3810 6784 3852 6824
rect 3892 6784 3934 6824
rect 3974 6784 4016 6824
rect 4056 6784 18808 6824
rect 18848 6784 18890 6824
rect 18930 6784 18972 6824
rect 19012 6784 19054 6824
rect 19094 6784 19136 6824
rect 19176 6784 33928 6824
rect 33968 6784 34010 6824
rect 34050 6784 34092 6824
rect 34132 6784 34174 6824
rect 34214 6784 34256 6824
rect 34296 6784 45216 6824
rect 1152 6760 45216 6784
rect 28347 6656 28389 6665
rect 28347 6616 28348 6656
rect 28388 6616 28389 6656
rect 28347 6607 28389 6616
rect 20187 6572 20229 6581
rect 20187 6532 20188 6572
rect 20228 6532 20229 6572
rect 20187 6523 20229 6532
rect 10827 6488 10869 6497
rect 10827 6448 10828 6488
rect 10868 6448 10869 6488
rect 10827 6439 10869 6448
rect 19947 6488 19989 6497
rect 19947 6448 19948 6488
rect 19988 6448 19989 6488
rect 19947 6439 19989 6448
rect 20379 6488 20421 6497
rect 20379 6448 20380 6488
rect 20420 6448 20421 6488
rect 20379 6439 20421 6448
rect 28107 6488 28149 6497
rect 28107 6448 28108 6488
rect 28148 6448 28149 6488
rect 28107 6439 28149 6448
rect 33195 6488 33237 6497
rect 33195 6448 33196 6488
rect 33236 6448 33237 6488
rect 33195 6439 33237 6448
rect 44523 6488 44565 6497
rect 44523 6448 44524 6488
rect 44564 6448 44565 6488
rect 44523 6439 44565 6448
rect 44907 6488 44949 6497
rect 44907 6448 44908 6488
rect 44948 6448 44949 6488
rect 44907 6439 44949 6448
rect 45147 6488 45189 6497
rect 45147 6448 45148 6488
rect 45188 6448 45189 6488
rect 45147 6439 45189 6448
rect 11067 6236 11109 6245
rect 11067 6196 11068 6236
rect 11108 6196 11109 6236
rect 11067 6187 11109 6196
rect 20667 6236 20709 6245
rect 20667 6196 20668 6236
rect 20708 6196 20709 6236
rect 20667 6187 20709 6196
rect 33435 6236 33477 6245
rect 33435 6196 33436 6236
rect 33476 6196 33477 6236
rect 33435 6187 33477 6196
rect 44763 6236 44805 6245
rect 44763 6196 44764 6236
rect 44804 6196 44805 6236
rect 44763 6187 44805 6196
rect 1152 6068 45216 6092
rect 1152 6028 4928 6068
rect 4968 6028 5010 6068
rect 5050 6028 5092 6068
rect 5132 6028 5174 6068
rect 5214 6028 5256 6068
rect 5296 6028 20048 6068
rect 20088 6028 20130 6068
rect 20170 6028 20212 6068
rect 20252 6028 20294 6068
rect 20334 6028 20376 6068
rect 20416 6028 35168 6068
rect 35208 6028 35250 6068
rect 35290 6028 35332 6068
rect 35372 6028 35414 6068
rect 35454 6028 35496 6068
rect 35536 6028 45216 6068
rect 1152 6004 45216 6028
rect 11739 5900 11781 5909
rect 11739 5860 11740 5900
rect 11780 5860 11781 5900
rect 11739 5851 11781 5860
rect 12507 5816 12549 5825
rect 12507 5776 12508 5816
rect 12548 5776 12549 5816
rect 12507 5767 12549 5776
rect 45147 5816 45189 5825
rect 45147 5776 45148 5816
rect 45188 5776 45189 5816
rect 45147 5767 45189 5776
rect 6699 5648 6741 5657
rect 6699 5608 6700 5648
rect 6740 5608 6741 5648
rect 6699 5599 6741 5608
rect 7563 5648 7605 5657
rect 7563 5608 7564 5648
rect 7604 5608 7605 5648
rect 7563 5599 7605 5608
rect 8715 5648 8757 5657
rect 8715 5608 8716 5648
rect 8756 5608 8757 5648
rect 8715 5599 8757 5608
rect 8955 5648 8997 5657
rect 8955 5608 8956 5648
rect 8996 5608 8997 5648
rect 8955 5599 8997 5608
rect 9867 5648 9909 5657
rect 9867 5608 9868 5648
rect 9908 5608 9909 5648
rect 9867 5599 9909 5608
rect 10827 5648 10869 5657
rect 10827 5608 10828 5648
rect 10868 5608 10869 5648
rect 10827 5599 10869 5608
rect 11499 5648 11541 5657
rect 11499 5608 11500 5648
rect 11540 5608 11541 5648
rect 11499 5599 11541 5608
rect 12267 5648 12309 5657
rect 12267 5608 12268 5648
rect 12308 5608 12309 5648
rect 12267 5599 12309 5608
rect 13515 5648 13557 5657
rect 13515 5608 13516 5648
rect 13556 5608 13557 5648
rect 13515 5599 13557 5608
rect 21003 5648 21045 5657
rect 21003 5608 21004 5648
rect 21044 5608 21045 5648
rect 21003 5599 21045 5608
rect 21387 5648 21429 5657
rect 21387 5608 21388 5648
rect 21428 5608 21429 5648
rect 21387 5599 21429 5608
rect 21771 5648 21813 5657
rect 21771 5608 21772 5648
rect 21812 5608 21813 5648
rect 21771 5599 21813 5608
rect 22011 5648 22053 5657
rect 22011 5608 22012 5648
rect 22052 5608 22053 5648
rect 22011 5599 22053 5608
rect 34155 5648 34197 5657
rect 34155 5608 34156 5648
rect 34196 5608 34197 5648
rect 34155 5599 34197 5608
rect 36939 5648 36981 5657
rect 36939 5608 36940 5648
rect 36980 5608 36981 5648
rect 36939 5599 36981 5608
rect 37515 5648 37557 5657
rect 37515 5608 37516 5648
rect 37556 5608 37557 5648
rect 37515 5599 37557 5608
rect 37899 5648 37941 5657
rect 37899 5608 37900 5648
rect 37940 5608 37941 5648
rect 37899 5599 37941 5608
rect 38091 5648 38133 5657
rect 38091 5608 38092 5648
rect 38132 5608 38133 5648
rect 38091 5599 38133 5608
rect 38475 5648 38517 5657
rect 38475 5608 38476 5648
rect 38516 5608 38517 5648
rect 38475 5599 38517 5608
rect 38715 5648 38757 5657
rect 38715 5608 38716 5648
rect 38756 5608 38757 5648
rect 38715 5599 38757 5608
rect 44523 5648 44565 5657
rect 44523 5608 44524 5648
rect 44564 5608 44565 5648
rect 44523 5599 44565 5608
rect 44907 5648 44949 5657
rect 44907 5608 44908 5648
rect 44948 5608 44949 5648
rect 44907 5599 44949 5608
rect 6939 5564 6981 5573
rect 6939 5524 6940 5564
rect 6980 5524 6981 5564
rect 6939 5515 6981 5524
rect 10107 5564 10149 5573
rect 10107 5524 10108 5564
rect 10148 5524 10149 5564
rect 10107 5515 10149 5524
rect 21627 5564 21669 5573
rect 21627 5524 21628 5564
rect 21668 5524 21669 5564
rect 21627 5515 21669 5524
rect 38331 5564 38373 5573
rect 38331 5524 38332 5564
rect 38372 5524 38373 5564
rect 38331 5515 38373 5524
rect 44763 5564 44805 5573
rect 44763 5524 44764 5564
rect 44804 5524 44805 5564
rect 44763 5515 44805 5524
rect 7803 5480 7845 5489
rect 7803 5440 7804 5480
rect 7844 5440 7845 5480
rect 7803 5431 7845 5440
rect 11067 5480 11109 5489
rect 11067 5440 11068 5480
rect 11108 5440 11109 5480
rect 11067 5431 11109 5440
rect 13755 5480 13797 5489
rect 13755 5440 13756 5480
rect 13796 5440 13797 5480
rect 13755 5431 13797 5440
rect 21243 5480 21285 5489
rect 21243 5440 21244 5480
rect 21284 5440 21285 5480
rect 21243 5431 21285 5440
rect 34395 5480 34437 5489
rect 34395 5440 34396 5480
rect 34436 5440 34437 5480
rect 34395 5431 34437 5440
rect 37179 5480 37221 5489
rect 37179 5440 37180 5480
rect 37220 5440 37221 5480
rect 37179 5431 37221 5440
rect 1152 5312 45216 5336
rect 1152 5272 3688 5312
rect 3728 5272 3770 5312
rect 3810 5272 3852 5312
rect 3892 5272 3934 5312
rect 3974 5272 4016 5312
rect 4056 5272 18808 5312
rect 18848 5272 18890 5312
rect 18930 5272 18972 5312
rect 19012 5272 19054 5312
rect 19094 5272 19136 5312
rect 19176 5272 33928 5312
rect 33968 5272 34010 5312
rect 34050 5272 34092 5312
rect 34132 5272 34174 5312
rect 34214 5272 34256 5312
rect 34296 5272 45216 5312
rect 1152 5248 45216 5272
rect 38907 5144 38949 5153
rect 38907 5104 38908 5144
rect 38948 5104 38949 5144
rect 38907 5095 38949 5104
rect 45147 5144 45189 5153
rect 45147 5104 45148 5144
rect 45188 5104 45189 5144
rect 45147 5095 45189 5104
rect 28347 5060 28389 5069
rect 28347 5020 28348 5060
rect 28388 5020 28389 5060
rect 28347 5011 28389 5020
rect 41019 5060 41061 5069
rect 41019 5020 41020 5060
rect 41060 5020 41061 5060
rect 41019 5011 41061 5020
rect 7179 4976 7221 4985
rect 7179 4936 7180 4976
rect 7220 4936 7221 4976
rect 7179 4927 7221 4936
rect 7419 4976 7461 4985
rect 7419 4936 7420 4976
rect 7460 4936 7461 4976
rect 7419 4927 7461 4936
rect 7563 4976 7605 4985
rect 7563 4936 7564 4976
rect 7604 4936 7605 4976
rect 7563 4927 7605 4936
rect 8331 4976 8373 4985
rect 8331 4936 8332 4976
rect 8372 4936 8373 4976
rect 8331 4927 8373 4936
rect 22059 4976 22101 4985
rect 22059 4936 22060 4976
rect 22100 4936 22101 4976
rect 22059 4927 22101 4936
rect 22299 4976 22341 4985
rect 22299 4936 22300 4976
rect 22340 4936 22341 4976
rect 22299 4927 22341 4936
rect 22474 4976 22532 4977
rect 22474 4936 22483 4976
rect 22523 4936 22532 4976
rect 22474 4935 22532 4936
rect 22923 4976 22965 4985
rect 22923 4936 22924 4976
rect 22964 4936 22965 4976
rect 22923 4927 22965 4936
rect 23403 4976 23445 4985
rect 23403 4936 23404 4976
rect 23444 4936 23445 4976
rect 23403 4927 23445 4936
rect 26859 4976 26901 4985
rect 26859 4936 26860 4976
rect 26900 4936 26901 4976
rect 26859 4927 26901 4936
rect 27723 4976 27765 4985
rect 27723 4936 27724 4976
rect 27764 4936 27765 4976
rect 27723 4927 27765 4936
rect 28107 4976 28149 4985
rect 28107 4936 28108 4976
rect 28148 4936 28149 4976
rect 28107 4927 28149 4936
rect 28491 4976 28533 4985
rect 28491 4936 28492 4976
rect 28532 4936 28533 4976
rect 28491 4927 28533 4936
rect 34155 4976 34197 4985
rect 34155 4936 34156 4976
rect 34196 4936 34197 4976
rect 34155 4927 34197 4936
rect 34443 4976 34485 4985
rect 34443 4936 34444 4976
rect 34484 4936 34485 4976
rect 34443 4927 34485 4936
rect 38667 4976 38709 4985
rect 38667 4936 38668 4976
rect 38708 4936 38709 4976
rect 38667 4927 38709 4936
rect 39627 4976 39669 4985
rect 39627 4936 39628 4976
rect 39668 4936 39669 4976
rect 39627 4927 39669 4936
rect 40491 4976 40533 4985
rect 40491 4936 40492 4976
rect 40532 4936 40533 4976
rect 40491 4927 40533 4936
rect 40779 4976 40821 4985
rect 40779 4936 40780 4976
rect 40820 4936 40821 4976
rect 40779 4927 40821 4936
rect 41163 4976 41205 4985
rect 41163 4936 41164 4976
rect 41204 4936 41205 4976
rect 41163 4927 41205 4936
rect 44523 4976 44565 4985
rect 44523 4936 44524 4976
rect 44564 4936 44565 4976
rect 44523 4927 44565 4936
rect 44907 4976 44949 4985
rect 44907 4936 44908 4976
rect 44948 4936 44949 4976
rect 44907 4927 44949 4936
rect 40107 4892 40149 4901
rect 40107 4852 40108 4892
rect 40148 4852 40149 4892
rect 40107 4843 40149 4852
rect 41547 4892 41589 4901
rect 41547 4852 41548 4892
rect 41588 4852 41589 4892
rect 41547 4843 41589 4852
rect 41835 4892 41877 4901
rect 41835 4852 41836 4892
rect 41876 4852 41877 4892
rect 41835 4843 41877 4852
rect 27963 4808 28005 4817
rect 27963 4768 27964 4808
rect 28004 4768 28005 4808
rect 27963 4759 28005 4768
rect 39867 4808 39909 4817
rect 39867 4768 39868 4808
rect 39908 4768 39909 4808
rect 39867 4759 39909 4768
rect 41403 4808 41445 4817
rect 41403 4768 41404 4808
rect 41444 4768 41445 4808
rect 41403 4759 41445 4768
rect 44763 4808 44805 4817
rect 44763 4768 44764 4808
rect 44804 4768 44805 4808
rect 44763 4759 44805 4768
rect 7803 4724 7845 4733
rect 7803 4684 7804 4724
rect 7844 4684 7845 4724
rect 7803 4675 7845 4684
rect 8571 4724 8613 4733
rect 8571 4684 8572 4724
rect 8612 4684 8613 4724
rect 8571 4675 8613 4684
rect 22683 4724 22725 4733
rect 22683 4684 22684 4724
rect 22724 4684 22725 4724
rect 22683 4675 22725 4684
rect 23163 4724 23205 4733
rect 23163 4684 23164 4724
rect 23204 4684 23205 4724
rect 23163 4675 23205 4684
rect 23643 4724 23685 4733
rect 23643 4684 23644 4724
rect 23684 4684 23685 4724
rect 23643 4675 23685 4684
rect 27099 4724 27141 4733
rect 27099 4684 27100 4724
rect 27140 4684 27141 4724
rect 27099 4675 27141 4684
rect 28731 4724 28773 4733
rect 28731 4684 28732 4724
rect 28772 4684 28773 4724
rect 28731 4675 28773 4684
rect 37690 4724 37748 4725
rect 37690 4684 37699 4724
rect 37739 4684 37748 4724
rect 37690 4683 37748 4684
rect 38362 4724 38420 4725
rect 38362 4684 38371 4724
rect 38411 4684 38420 4724
rect 38362 4683 38420 4684
rect 39034 4724 39092 4725
rect 39034 4684 39043 4724
rect 39083 4684 39092 4724
rect 39034 4683 39092 4684
rect 39322 4724 39380 4725
rect 39322 4684 39331 4724
rect 39371 4684 39380 4724
rect 39322 4683 39380 4684
rect 40090 4724 40148 4725
rect 40090 4684 40099 4724
rect 40139 4684 40148 4724
rect 40090 4683 40148 4684
rect 40474 4724 40532 4725
rect 40474 4684 40483 4724
rect 40523 4684 40532 4724
rect 40474 4683 40532 4684
rect 41818 4724 41876 4725
rect 41818 4684 41827 4724
rect 41867 4684 41876 4724
rect 41818 4683 41876 4684
rect 1152 4556 45216 4580
rect 1152 4516 4928 4556
rect 4968 4516 5010 4556
rect 5050 4516 5092 4556
rect 5132 4516 5174 4556
rect 5214 4516 5256 4556
rect 5296 4516 20048 4556
rect 20088 4516 20130 4556
rect 20170 4516 20212 4556
rect 20252 4516 20294 4556
rect 20334 4516 20376 4556
rect 20416 4516 35168 4556
rect 35208 4516 35250 4556
rect 35290 4516 35332 4556
rect 35372 4516 35414 4556
rect 35454 4516 35496 4556
rect 35536 4516 45216 4556
rect 1152 4492 45216 4516
rect 39322 4388 39380 4389
rect 39322 4348 39331 4388
rect 39371 4348 39380 4388
rect 39322 4347 39380 4348
rect 39994 4388 40052 4389
rect 39994 4348 40003 4388
rect 40043 4348 40052 4388
rect 39994 4347 40052 4348
rect 40474 4388 40532 4389
rect 40474 4348 40483 4388
rect 40523 4348 40532 4388
rect 40474 4347 40532 4348
rect 40762 4388 40820 4389
rect 40762 4348 40771 4388
rect 40811 4348 40820 4388
rect 40762 4347 40820 4348
rect 41050 4388 41108 4389
rect 41050 4348 41059 4388
rect 41099 4348 41108 4388
rect 41050 4347 41108 4348
rect 41338 4388 41396 4389
rect 41338 4348 41347 4388
rect 41387 4348 41396 4388
rect 41338 4347 41396 4348
rect 41626 4388 41684 4389
rect 41626 4348 41635 4388
rect 41675 4348 41684 4388
rect 41626 4347 41684 4348
rect 42202 4388 42260 4389
rect 42202 4348 42211 4388
rect 42251 4348 42260 4388
rect 42202 4347 42260 4348
rect 42778 4388 42836 4389
rect 42778 4348 42787 4388
rect 42827 4348 42836 4388
rect 42778 4347 42836 4348
rect 41931 4304 41973 4313
rect 41931 4264 41932 4304
rect 41972 4264 41973 4304
rect 41931 4255 41973 4264
rect 42507 4304 42549 4313
rect 42507 4264 42508 4304
rect 42548 4264 42549 4304
rect 42507 4255 42549 4264
rect 45147 4304 45189 4313
rect 45147 4264 45148 4304
rect 45188 4264 45189 4304
rect 45147 4255 45189 4264
rect 7083 4136 7125 4145
rect 7083 4096 7084 4136
rect 7124 4096 7125 4136
rect 7083 4087 7125 4096
rect 23979 4136 24021 4145
rect 23979 4096 23980 4136
rect 24020 4096 24021 4136
rect 23979 4087 24021 4096
rect 24459 4136 24501 4145
rect 24459 4096 24460 4136
rect 24500 4096 24501 4136
rect 24459 4087 24501 4096
rect 25323 4136 25365 4145
rect 25323 4096 25324 4136
rect 25364 4096 25365 4136
rect 25323 4087 25365 4096
rect 25563 4136 25605 4145
rect 25563 4096 25564 4136
rect 25604 4096 25605 4136
rect 25563 4087 25605 4096
rect 26187 4136 26229 4145
rect 26187 4096 26188 4136
rect 26228 4096 26229 4136
rect 26187 4087 26229 4096
rect 26427 4136 26469 4145
rect 26427 4096 26428 4136
rect 26468 4096 26469 4136
rect 26427 4087 26469 4096
rect 27627 4136 27669 4145
rect 27627 4096 27628 4136
rect 27668 4096 27669 4136
rect 27627 4087 27669 4096
rect 27867 4136 27909 4145
rect 27867 4096 27868 4136
rect 27908 4096 27909 4136
rect 27867 4087 27909 4096
rect 32619 4136 32661 4145
rect 32619 4096 32620 4136
rect 32660 4096 32661 4136
rect 32619 4087 32661 4096
rect 32859 4136 32901 4145
rect 32859 4096 32860 4136
rect 32900 4096 32901 4136
rect 32859 4087 32901 4096
rect 44139 4136 44181 4145
rect 44139 4096 44140 4136
rect 44180 4096 44181 4136
rect 44139 4087 44181 4096
rect 44523 4136 44565 4145
rect 44523 4096 44524 4136
rect 44564 4096 44565 4136
rect 44523 4087 44565 4096
rect 44907 4136 44949 4145
rect 44907 4096 44908 4136
rect 44948 4096 44949 4136
rect 44907 4087 44949 4096
rect 24699 4052 24741 4061
rect 24699 4012 24700 4052
rect 24740 4012 24741 4052
rect 24699 4003 24741 4012
rect 44763 4052 44805 4061
rect 44763 4012 44764 4052
rect 44804 4012 44805 4052
rect 44763 4003 44805 4012
rect 7323 3968 7365 3977
rect 7323 3928 7324 3968
rect 7364 3928 7365 3968
rect 7323 3919 7365 3928
rect 24219 3968 24261 3977
rect 24219 3928 24220 3968
rect 24260 3928 24261 3968
rect 24219 3919 24261 3928
rect 44379 3968 44421 3977
rect 44379 3928 44380 3968
rect 44420 3928 44421 3968
rect 44379 3919 44421 3928
rect 1152 3800 45216 3824
rect 1152 3760 3688 3800
rect 3728 3760 3770 3800
rect 3810 3760 3852 3800
rect 3892 3760 3934 3800
rect 3974 3760 4016 3800
rect 4056 3760 18808 3800
rect 18848 3760 18890 3800
rect 18930 3760 18972 3800
rect 19012 3760 19054 3800
rect 19094 3760 19136 3800
rect 19176 3760 33928 3800
rect 33968 3760 34010 3800
rect 34050 3760 34092 3800
rect 34132 3760 34174 3800
rect 34214 3760 34256 3800
rect 34296 3760 45216 3800
rect 1152 3736 45216 3760
rect 26907 3632 26949 3641
rect 26907 3592 26908 3632
rect 26948 3592 26949 3632
rect 26907 3583 26949 3592
rect 27291 3632 27333 3641
rect 27291 3592 27292 3632
rect 27332 3592 27333 3632
rect 27291 3583 27333 3592
rect 27675 3632 27717 3641
rect 27675 3592 27676 3632
rect 27716 3592 27717 3632
rect 27675 3583 27717 3592
rect 30939 3632 30981 3641
rect 30939 3592 30940 3632
rect 30980 3592 30981 3632
rect 30939 3583 30981 3592
rect 38139 3632 38181 3641
rect 38139 3592 38140 3632
rect 38180 3592 38181 3632
rect 38139 3583 38181 3592
rect 45147 3632 45189 3641
rect 45147 3592 45148 3632
rect 45188 3592 45189 3632
rect 45147 3583 45189 3592
rect 25899 3464 25941 3473
rect 25899 3424 25900 3464
rect 25940 3424 25941 3464
rect 25899 3415 25941 3424
rect 26283 3464 26325 3473
rect 26283 3424 26284 3464
rect 26324 3424 26325 3464
rect 26283 3415 26325 3424
rect 26667 3464 26709 3473
rect 26667 3424 26668 3464
rect 26708 3424 26709 3464
rect 26667 3415 26709 3424
rect 27051 3464 27093 3473
rect 27051 3424 27052 3464
rect 27092 3424 27093 3464
rect 27051 3415 27093 3424
rect 27435 3464 27477 3473
rect 27435 3424 27436 3464
rect 27476 3424 27477 3464
rect 27435 3415 27477 3424
rect 27819 3464 27861 3473
rect 27819 3424 27820 3464
rect 27860 3424 27861 3464
rect 27819 3415 27861 3424
rect 28203 3464 28245 3473
rect 28203 3424 28204 3464
rect 28244 3424 28245 3464
rect 28203 3415 28245 3424
rect 28443 3464 28485 3473
rect 28443 3424 28444 3464
rect 28484 3424 28485 3464
rect 28443 3415 28485 3424
rect 30027 3464 30069 3473
rect 30027 3424 30028 3464
rect 30068 3424 30069 3464
rect 30027 3415 30069 3424
rect 30699 3464 30741 3473
rect 30699 3424 30700 3464
rect 30740 3424 30741 3464
rect 30699 3415 30741 3424
rect 34827 3464 34869 3473
rect 34827 3424 34828 3464
rect 34868 3424 34869 3464
rect 34827 3415 34869 3424
rect 35067 3464 35109 3473
rect 35067 3424 35068 3464
rect 35108 3424 35109 3464
rect 35067 3415 35109 3424
rect 36555 3464 36597 3473
rect 36555 3424 36556 3464
rect 36596 3424 36597 3464
rect 36555 3415 36597 3424
rect 37899 3464 37941 3473
rect 37899 3424 37900 3464
rect 37940 3424 37941 3464
rect 37899 3415 37941 3424
rect 44523 3464 44565 3473
rect 44523 3424 44524 3464
rect 44564 3424 44565 3464
rect 44523 3415 44565 3424
rect 44907 3464 44949 3473
rect 44907 3424 44908 3464
rect 44948 3424 44949 3464
rect 44907 3415 44949 3424
rect 30267 3296 30309 3305
rect 30267 3256 30268 3296
rect 30308 3256 30309 3296
rect 30267 3247 30309 3256
rect 36795 3296 36837 3305
rect 36795 3256 36796 3296
rect 36836 3256 36837 3296
rect 36795 3247 36837 3256
rect 26139 3212 26181 3221
rect 26139 3172 26140 3212
rect 26180 3172 26181 3212
rect 26139 3163 26181 3172
rect 26523 3212 26565 3221
rect 26523 3172 26524 3212
rect 26564 3172 26565 3212
rect 26523 3163 26565 3172
rect 28059 3212 28101 3221
rect 28059 3172 28060 3212
rect 28100 3172 28101 3212
rect 28059 3163 28101 3172
rect 44763 3212 44805 3221
rect 44763 3172 44764 3212
rect 44804 3172 44805 3212
rect 44763 3163 44805 3172
rect 1152 3044 45216 3068
rect 1152 3004 4928 3044
rect 4968 3004 5010 3044
rect 5050 3004 5092 3044
rect 5132 3004 5174 3044
rect 5214 3004 5256 3044
rect 5296 3004 20048 3044
rect 20088 3004 20130 3044
rect 20170 3004 20212 3044
rect 20252 3004 20294 3044
rect 20334 3004 20376 3044
rect 20416 3004 35168 3044
rect 35208 3004 35250 3044
rect 35290 3004 35332 3044
rect 35372 3004 35414 3044
rect 35454 3004 35496 3044
rect 35536 3004 45216 3044
rect 1152 2980 45216 3004
rect 34827 2876 34869 2885
rect 34827 2836 34828 2876
rect 34868 2836 34869 2876
rect 34827 2827 34869 2836
rect 35098 2876 35156 2877
rect 35098 2836 35107 2876
rect 35147 2836 35156 2876
rect 35098 2835 35156 2836
rect 45147 2792 45189 2801
rect 45147 2752 45148 2792
rect 45188 2752 45189 2792
rect 45147 2743 45189 2752
rect 21483 2624 21525 2633
rect 21483 2584 21484 2624
rect 21524 2584 21525 2624
rect 21483 2575 21525 2584
rect 21867 2624 21909 2633
rect 21867 2584 21868 2624
rect 21908 2584 21909 2624
rect 21867 2575 21909 2584
rect 22251 2624 22293 2633
rect 22251 2584 22252 2624
rect 22292 2584 22293 2624
rect 22251 2575 22293 2584
rect 22635 2624 22677 2633
rect 22635 2584 22636 2624
rect 22676 2584 22677 2624
rect 22635 2575 22677 2584
rect 23019 2624 23061 2633
rect 23019 2584 23020 2624
rect 23060 2584 23061 2624
rect 23019 2575 23061 2584
rect 23403 2624 23445 2633
rect 23403 2584 23404 2624
rect 23444 2584 23445 2624
rect 23403 2575 23445 2584
rect 23787 2624 23829 2633
rect 23787 2584 23788 2624
rect 23828 2584 23829 2624
rect 23787 2575 23829 2584
rect 25515 2624 25557 2633
rect 25515 2584 25516 2624
rect 25556 2584 25557 2624
rect 25515 2575 25557 2584
rect 25899 2624 25941 2633
rect 25899 2584 25900 2624
rect 25940 2584 25941 2624
rect 25899 2575 25941 2584
rect 26283 2624 26325 2633
rect 26283 2584 26284 2624
rect 26324 2584 26325 2624
rect 26283 2575 26325 2584
rect 26667 2624 26709 2633
rect 26667 2584 26668 2624
rect 26708 2584 26709 2624
rect 26667 2575 26709 2584
rect 27051 2624 27093 2633
rect 27051 2584 27052 2624
rect 27092 2584 27093 2624
rect 27051 2575 27093 2584
rect 27435 2624 27477 2633
rect 27435 2584 27436 2624
rect 27476 2584 27477 2624
rect 27435 2575 27477 2584
rect 27819 2624 27861 2633
rect 27819 2584 27820 2624
rect 27860 2584 27861 2624
rect 27819 2575 27861 2584
rect 28203 2624 28245 2633
rect 28203 2584 28204 2624
rect 28244 2584 28245 2624
rect 28203 2575 28245 2584
rect 28587 2624 28629 2633
rect 28587 2584 28588 2624
rect 28628 2584 28629 2624
rect 28587 2575 28629 2584
rect 28971 2624 29013 2633
rect 28971 2584 28972 2624
rect 29012 2584 29013 2624
rect 28971 2575 29013 2584
rect 29355 2624 29397 2633
rect 29355 2584 29356 2624
rect 29396 2584 29397 2624
rect 29355 2575 29397 2584
rect 29739 2624 29781 2633
rect 29739 2584 29740 2624
rect 29780 2584 29781 2624
rect 29739 2575 29781 2584
rect 30123 2624 30165 2633
rect 30123 2584 30124 2624
rect 30164 2584 30165 2624
rect 30123 2575 30165 2584
rect 30507 2624 30549 2633
rect 30507 2584 30508 2624
rect 30548 2584 30549 2624
rect 30507 2575 30549 2584
rect 30891 2624 30933 2633
rect 30891 2584 30892 2624
rect 30932 2584 30933 2624
rect 30891 2575 30933 2584
rect 31275 2624 31317 2633
rect 31275 2584 31276 2624
rect 31316 2584 31317 2624
rect 31275 2575 31317 2584
rect 44139 2624 44181 2633
rect 44139 2584 44140 2624
rect 44180 2584 44181 2624
rect 44139 2575 44181 2584
rect 44523 2624 44565 2633
rect 44523 2584 44524 2624
rect 44564 2584 44565 2624
rect 44523 2575 44565 2584
rect 44907 2624 44949 2633
rect 44907 2584 44908 2624
rect 44948 2584 44949 2624
rect 44907 2575 44949 2584
rect 44763 2540 44805 2549
rect 44763 2500 44764 2540
rect 44804 2500 44805 2540
rect 44763 2491 44805 2500
rect 21243 2456 21285 2465
rect 21243 2416 21244 2456
rect 21284 2416 21285 2456
rect 21243 2407 21285 2416
rect 21627 2456 21669 2465
rect 21627 2416 21628 2456
rect 21668 2416 21669 2456
rect 21627 2407 21669 2416
rect 22011 2456 22053 2465
rect 22011 2416 22012 2456
rect 22052 2416 22053 2456
rect 22011 2407 22053 2416
rect 22395 2456 22437 2465
rect 22395 2416 22396 2456
rect 22436 2416 22437 2456
rect 22395 2407 22437 2416
rect 22779 2456 22821 2465
rect 22779 2416 22780 2456
rect 22820 2416 22821 2456
rect 22779 2407 22821 2416
rect 23163 2456 23205 2465
rect 23163 2416 23164 2456
rect 23204 2416 23205 2456
rect 23163 2407 23205 2416
rect 23547 2456 23589 2465
rect 23547 2416 23548 2456
rect 23588 2416 23589 2456
rect 23547 2407 23589 2416
rect 25275 2456 25317 2465
rect 25275 2416 25276 2456
rect 25316 2416 25317 2456
rect 25275 2407 25317 2416
rect 25659 2456 25701 2465
rect 25659 2416 25660 2456
rect 25700 2416 25701 2456
rect 25659 2407 25701 2416
rect 26043 2456 26085 2465
rect 26043 2416 26044 2456
rect 26084 2416 26085 2456
rect 26043 2407 26085 2416
rect 26427 2456 26469 2465
rect 26427 2416 26428 2456
rect 26468 2416 26469 2456
rect 26427 2407 26469 2416
rect 26811 2456 26853 2465
rect 26811 2416 26812 2456
rect 26852 2416 26853 2456
rect 26811 2407 26853 2416
rect 27195 2456 27237 2465
rect 27195 2416 27196 2456
rect 27236 2416 27237 2456
rect 27195 2407 27237 2416
rect 27579 2456 27621 2465
rect 27579 2416 27580 2456
rect 27620 2416 27621 2456
rect 27579 2407 27621 2416
rect 27963 2456 28005 2465
rect 27963 2416 27964 2456
rect 28004 2416 28005 2456
rect 27963 2407 28005 2416
rect 28347 2456 28389 2465
rect 28347 2416 28348 2456
rect 28388 2416 28389 2456
rect 28347 2407 28389 2416
rect 28731 2456 28773 2465
rect 28731 2416 28732 2456
rect 28772 2416 28773 2456
rect 28731 2407 28773 2416
rect 29115 2456 29157 2465
rect 29115 2416 29116 2456
rect 29156 2416 29157 2456
rect 29115 2407 29157 2416
rect 29499 2456 29541 2465
rect 29499 2416 29500 2456
rect 29540 2416 29541 2456
rect 29499 2407 29541 2416
rect 29883 2456 29925 2465
rect 29883 2416 29884 2456
rect 29924 2416 29925 2456
rect 29883 2407 29925 2416
rect 30267 2456 30309 2465
rect 30267 2416 30268 2456
rect 30308 2416 30309 2456
rect 30267 2407 30309 2416
rect 30651 2456 30693 2465
rect 30651 2416 30652 2456
rect 30692 2416 30693 2456
rect 30651 2407 30693 2416
rect 31035 2456 31077 2465
rect 31035 2416 31036 2456
rect 31076 2416 31077 2456
rect 31035 2407 31077 2416
rect 44379 2456 44421 2465
rect 44379 2416 44380 2456
rect 44420 2416 44421 2456
rect 44379 2407 44421 2416
rect 1152 2288 45216 2312
rect 1152 2248 3688 2288
rect 3728 2248 3770 2288
rect 3810 2248 3852 2288
rect 3892 2248 3934 2288
rect 3974 2248 4016 2288
rect 4056 2248 18808 2288
rect 18848 2248 18890 2288
rect 18930 2248 18972 2288
rect 19012 2248 19054 2288
rect 19094 2248 19136 2288
rect 19176 2248 33928 2288
rect 33968 2248 34010 2288
rect 34050 2248 34092 2288
rect 34132 2248 34174 2288
rect 34214 2248 34256 2288
rect 34296 2248 45216 2288
rect 1152 2224 45216 2248
rect 45147 2120 45189 2129
rect 45147 2080 45148 2120
rect 45188 2080 45189 2120
rect 45147 2071 45189 2080
rect 27003 2036 27045 2045
rect 27003 1996 27004 2036
rect 27044 1996 27045 2036
rect 27003 1987 27045 1996
rect 30075 2036 30117 2045
rect 30075 1996 30076 2036
rect 30116 1996 30117 2036
rect 30075 1987 30117 1996
rect 20907 1952 20949 1961
rect 20907 1912 20908 1952
rect 20948 1912 20949 1952
rect 20907 1903 20949 1912
rect 21291 1952 21333 1961
rect 21291 1912 21292 1952
rect 21332 1912 21333 1952
rect 21291 1903 21333 1912
rect 21675 1952 21717 1961
rect 21675 1912 21676 1952
rect 21716 1912 21717 1952
rect 21675 1903 21717 1912
rect 22059 1952 22101 1961
rect 22059 1912 22060 1952
rect 22100 1912 22101 1952
rect 22059 1903 22101 1912
rect 22443 1952 22485 1961
rect 22443 1912 22444 1952
rect 22484 1912 22485 1952
rect 22443 1903 22485 1912
rect 22827 1952 22869 1961
rect 22827 1912 22828 1952
rect 22868 1912 22869 1952
rect 22827 1903 22869 1912
rect 23211 1952 23253 1961
rect 23211 1912 23212 1952
rect 23252 1912 23253 1952
rect 23211 1903 23253 1912
rect 23595 1952 23637 1961
rect 23595 1912 23596 1952
rect 23636 1912 23637 1952
rect 23595 1903 23637 1912
rect 23979 1952 24021 1961
rect 23979 1912 23980 1952
rect 24020 1912 24021 1952
rect 23979 1903 24021 1912
rect 24555 1952 24597 1961
rect 24555 1912 24556 1952
rect 24596 1912 24597 1952
rect 24555 1903 24597 1912
rect 24939 1952 24981 1961
rect 24939 1912 24940 1952
rect 24980 1912 24981 1952
rect 24939 1903 24981 1912
rect 25323 1952 25365 1961
rect 25323 1912 25324 1952
rect 25364 1912 25365 1952
rect 25323 1903 25365 1912
rect 25707 1952 25749 1961
rect 25707 1912 25708 1952
rect 25748 1912 25749 1952
rect 25707 1903 25749 1912
rect 26091 1952 26133 1961
rect 26091 1912 26092 1952
rect 26132 1912 26133 1952
rect 26091 1903 26133 1912
rect 26475 1952 26517 1961
rect 26475 1912 26476 1952
rect 26516 1912 26517 1952
rect 26475 1903 26517 1912
rect 26859 1952 26901 1961
rect 26859 1912 26860 1952
rect 26900 1912 26901 1952
rect 26859 1903 26901 1912
rect 27243 1952 27285 1961
rect 27243 1912 27244 1952
rect 27284 1912 27285 1952
rect 27243 1903 27285 1912
rect 27627 1952 27669 1961
rect 27627 1912 27628 1952
rect 27668 1912 27669 1952
rect 27627 1903 27669 1912
rect 28011 1952 28053 1961
rect 28011 1912 28012 1952
rect 28052 1912 28053 1952
rect 28011 1903 28053 1912
rect 28395 1952 28437 1961
rect 28395 1912 28396 1952
rect 28436 1912 28437 1952
rect 28395 1903 28437 1912
rect 28779 1952 28821 1961
rect 28779 1912 28780 1952
rect 28820 1912 28821 1952
rect 28779 1903 28821 1912
rect 29163 1952 29205 1961
rect 29163 1912 29164 1952
rect 29204 1912 29205 1952
rect 29163 1903 29205 1912
rect 29547 1952 29589 1961
rect 29547 1912 29548 1952
rect 29588 1912 29589 1952
rect 29547 1903 29589 1912
rect 29931 1952 29973 1961
rect 29931 1912 29932 1952
rect 29972 1912 29973 1952
rect 29931 1903 29973 1912
rect 30315 1952 30357 1961
rect 30315 1912 30316 1952
rect 30356 1912 30357 1952
rect 30315 1903 30357 1912
rect 30699 1952 30741 1961
rect 30699 1912 30700 1952
rect 30740 1912 30741 1952
rect 30699 1903 30741 1912
rect 31083 1952 31125 1961
rect 31083 1912 31084 1952
rect 31124 1912 31125 1952
rect 31083 1903 31125 1912
rect 31467 1952 31509 1961
rect 31467 1912 31468 1952
rect 31508 1912 31509 1952
rect 31467 1903 31509 1912
rect 31851 1952 31893 1961
rect 31851 1912 31852 1952
rect 31892 1912 31893 1952
rect 31851 1903 31893 1912
rect 43755 1952 43797 1961
rect 43755 1912 43756 1952
rect 43796 1912 43797 1952
rect 43755 1903 43797 1912
rect 44139 1952 44181 1961
rect 44139 1912 44140 1952
rect 44180 1912 44181 1952
rect 44139 1903 44181 1912
rect 44523 1952 44565 1961
rect 44523 1912 44524 1952
rect 44564 1912 44565 1952
rect 44523 1903 44565 1912
rect 44907 1952 44949 1961
rect 44907 1912 44908 1952
rect 44948 1912 44949 1952
rect 44907 1903 44949 1912
rect 24219 1784 24261 1793
rect 24219 1744 24220 1784
rect 24260 1744 24261 1784
rect 24219 1735 24261 1744
rect 25083 1784 25125 1793
rect 25083 1744 25084 1784
rect 25124 1744 25125 1784
rect 25083 1735 25125 1744
rect 26235 1784 26277 1793
rect 26235 1744 26236 1784
rect 26276 1744 26277 1784
rect 26235 1735 26277 1744
rect 27771 1784 27813 1793
rect 27771 1744 27772 1784
rect 27812 1744 27813 1784
rect 27771 1735 27813 1744
rect 28923 1784 28965 1793
rect 28923 1744 28924 1784
rect 28964 1744 28965 1784
rect 28923 1735 28965 1744
rect 30843 1784 30885 1793
rect 30843 1744 30844 1784
rect 30884 1744 30885 1784
rect 30843 1735 30885 1744
rect 43995 1784 44037 1793
rect 43995 1744 43996 1784
rect 44036 1744 44037 1784
rect 43995 1735 44037 1744
rect 44763 1784 44805 1793
rect 44763 1744 44764 1784
rect 44804 1744 44805 1784
rect 44763 1735 44805 1744
rect 21147 1700 21189 1709
rect 21147 1660 21148 1700
rect 21188 1660 21189 1700
rect 21147 1651 21189 1660
rect 21531 1700 21573 1709
rect 21531 1660 21532 1700
rect 21572 1660 21573 1700
rect 21531 1651 21573 1660
rect 21915 1700 21957 1709
rect 21915 1660 21916 1700
rect 21956 1660 21957 1700
rect 21915 1651 21957 1660
rect 22299 1700 22341 1709
rect 22299 1660 22300 1700
rect 22340 1660 22341 1700
rect 22299 1651 22341 1660
rect 22683 1700 22725 1709
rect 22683 1660 22684 1700
rect 22724 1660 22725 1700
rect 22683 1651 22725 1660
rect 23067 1700 23109 1709
rect 23067 1660 23068 1700
rect 23108 1660 23109 1700
rect 23067 1651 23109 1660
rect 23451 1700 23493 1709
rect 23451 1660 23452 1700
rect 23492 1660 23493 1700
rect 23451 1651 23493 1660
rect 23835 1700 23877 1709
rect 23835 1660 23836 1700
rect 23876 1660 23877 1700
rect 23835 1651 23877 1660
rect 24315 1700 24357 1709
rect 24315 1660 24316 1700
rect 24356 1660 24357 1700
rect 24315 1651 24357 1660
rect 24699 1700 24741 1709
rect 24699 1660 24700 1700
rect 24740 1660 24741 1700
rect 24699 1651 24741 1660
rect 25467 1700 25509 1709
rect 25467 1660 25468 1700
rect 25508 1660 25509 1700
rect 25467 1651 25509 1660
rect 25851 1700 25893 1709
rect 25851 1660 25852 1700
rect 25892 1660 25893 1700
rect 25851 1651 25893 1660
rect 26619 1700 26661 1709
rect 26619 1660 26620 1700
rect 26660 1660 26661 1700
rect 26619 1651 26661 1660
rect 27387 1700 27429 1709
rect 27387 1660 27388 1700
rect 27428 1660 27429 1700
rect 27387 1651 27429 1660
rect 28155 1700 28197 1709
rect 28155 1660 28156 1700
rect 28196 1660 28197 1700
rect 28155 1651 28197 1660
rect 28539 1700 28581 1709
rect 28539 1660 28540 1700
rect 28580 1660 28581 1700
rect 28539 1651 28581 1660
rect 29307 1700 29349 1709
rect 29307 1660 29308 1700
rect 29348 1660 29349 1700
rect 29307 1651 29349 1660
rect 29691 1700 29733 1709
rect 29691 1660 29692 1700
rect 29732 1660 29733 1700
rect 29691 1651 29733 1660
rect 30459 1700 30501 1709
rect 30459 1660 30460 1700
rect 30500 1660 30501 1700
rect 30459 1651 30501 1660
rect 31227 1700 31269 1709
rect 31227 1660 31228 1700
rect 31268 1660 31269 1700
rect 31227 1651 31269 1660
rect 31611 1700 31653 1709
rect 31611 1660 31612 1700
rect 31652 1660 31653 1700
rect 31611 1651 31653 1660
rect 44379 1700 44421 1709
rect 44379 1660 44380 1700
rect 44420 1660 44421 1700
rect 44379 1651 44421 1660
rect 1152 1532 45216 1556
rect 1152 1492 4928 1532
rect 4968 1492 5010 1532
rect 5050 1492 5092 1532
rect 5132 1492 5174 1532
rect 5214 1492 5256 1532
rect 5296 1492 20048 1532
rect 20088 1492 20130 1532
rect 20170 1492 20212 1532
rect 20252 1492 20294 1532
rect 20334 1492 20376 1532
rect 20416 1492 35168 1532
rect 35208 1492 35250 1532
rect 35290 1492 35332 1532
rect 35372 1492 35414 1532
rect 35454 1492 35496 1532
rect 35536 1492 45216 1532
rect 1152 1468 45216 1492
<< via1 >>
rect 4928 10564 4968 10604
rect 5010 10564 5050 10604
rect 5092 10564 5132 10604
rect 5174 10564 5214 10604
rect 5256 10564 5296 10604
rect 20048 10564 20088 10604
rect 20130 10564 20170 10604
rect 20212 10564 20252 10604
rect 20294 10564 20334 10604
rect 20376 10564 20416 10604
rect 35168 10564 35208 10604
rect 35250 10564 35290 10604
rect 35332 10564 35372 10604
rect 35414 10564 35454 10604
rect 35496 10564 35536 10604
rect 2044 10396 2084 10436
rect 4156 10396 4196 10436
rect 6268 10396 6308 10436
rect 8380 10396 8420 10436
rect 10492 10396 10532 10436
rect 12604 10396 12644 10436
rect 14716 10396 14756 10436
rect 16828 10396 16868 10436
rect 18940 10396 18980 10436
rect 21052 10396 21092 10436
rect 23164 10396 23204 10436
rect 25276 10396 25316 10436
rect 27388 10396 27428 10436
rect 29500 10396 29540 10436
rect 31612 10396 31652 10436
rect 33724 10396 33764 10436
rect 35836 10396 35876 10436
rect 37948 10396 37988 10436
rect 40060 10396 40100 10436
rect 42172 10396 42212 10436
rect 43420 10396 43460 10436
rect 44284 10396 44324 10436
rect 2284 10144 2324 10184
rect 4396 10144 4436 10184
rect 6508 10144 6548 10184
rect 8620 10144 8660 10184
rect 10732 10144 10772 10184
rect 12844 10144 12884 10184
rect 14956 10144 14996 10184
rect 17068 10144 17108 10184
rect 19180 10144 19220 10184
rect 21292 10144 21332 10184
rect 23452 10144 23492 10184
rect 25516 10144 25556 10184
rect 27628 10144 27668 10184
rect 29740 10144 29780 10184
rect 31852 10144 31892 10184
rect 33964 10144 34004 10184
rect 36076 10144 36116 10184
rect 38188 10144 38228 10184
rect 40300 10144 40340 10184
rect 42412 10144 42452 10184
rect 43180 10144 43220 10184
rect 43564 10144 43604 10184
rect 43948 10144 43988 10184
rect 44524 10144 44564 10184
rect 44908 10144 44948 10184
rect 43804 10060 43844 10100
rect 44188 9976 44228 10016
rect 45148 9976 45188 10016
rect 3688 9808 3728 9848
rect 3770 9808 3810 9848
rect 3852 9808 3892 9848
rect 3934 9808 3974 9848
rect 4016 9808 4056 9848
rect 18808 9808 18848 9848
rect 18890 9808 18930 9848
rect 18972 9808 19012 9848
rect 19054 9808 19094 9848
rect 19136 9808 19176 9848
rect 33928 9808 33968 9848
rect 34010 9808 34050 9848
rect 34092 9808 34132 9848
rect 34174 9808 34214 9848
rect 34256 9808 34296 9848
rect 44380 9640 44420 9680
rect 43996 9556 44036 9596
rect 43756 9472 43796 9512
rect 44140 9472 44180 9512
rect 44524 9472 44564 9512
rect 44908 9472 44948 9512
rect 44764 9220 44804 9260
rect 45148 9220 45188 9260
rect 4928 9052 4968 9092
rect 5010 9052 5050 9092
rect 5092 9052 5132 9092
rect 5174 9052 5214 9092
rect 5256 9052 5296 9092
rect 20048 9052 20088 9092
rect 20130 9052 20170 9092
rect 20212 9052 20252 9092
rect 20294 9052 20334 9092
rect 20376 9052 20416 9092
rect 35168 9052 35208 9092
rect 35250 9052 35290 9092
rect 35332 9052 35372 9092
rect 35414 9052 35454 9092
rect 35496 9052 35536 9092
rect 6172 8884 6212 8924
rect 8572 8884 8612 8924
rect 13084 8884 13124 8924
rect 18748 8884 18788 8924
rect 21532 8884 21572 8924
rect 22300 8884 22340 8924
rect 23068 8884 23108 8924
rect 23452 8884 23492 8924
rect 23836 8884 23876 8924
rect 25852 8884 25892 8924
rect 26908 8884 26948 8924
rect 27292 8884 27332 8924
rect 28060 8884 28100 8924
rect 28732 8884 28772 8924
rect 29116 8884 29156 8924
rect 24412 8800 24452 8840
rect 27964 8800 28004 8840
rect 31228 8800 31268 8840
rect 6412 8632 6452 8672
rect 6652 8632 6692 8672
rect 6892 8632 6932 8672
rect 7468 8632 7508 8672
rect 7708 8632 7748 8672
rect 8812 8632 8852 8672
rect 13324 8632 13364 8672
rect 18988 8632 19028 8672
rect 21292 8632 21332 8672
rect 21676 8632 21716 8672
rect 22060 8632 22100 8672
rect 22444 8632 22484 8672
rect 22867 8632 22907 8672
rect 23212 8632 23252 8672
rect 23596 8632 23636 8672
rect 24172 8632 24212 8672
rect 26092 8632 26132 8672
rect 27148 8632 27188 8672
rect 27532 8632 27572 8672
rect 27724 8632 27764 8672
rect 28300 8632 28340 8672
rect 28492 8632 28532 8672
rect 29356 8632 29396 8672
rect 31468 8632 31508 8672
rect 31852 8632 31892 8672
rect 44524 8632 44564 8672
rect 44908 8632 44948 8672
rect 45148 8632 45188 8672
rect 22684 8548 22724 8588
rect 31612 8548 31652 8588
rect 44764 8548 44804 8588
rect 21916 8464 21956 8504
rect 3688 8296 3728 8336
rect 3770 8296 3810 8336
rect 3852 8296 3892 8336
rect 3934 8296 3974 8336
rect 4016 8296 4056 8336
rect 18808 8296 18848 8336
rect 18890 8296 18930 8336
rect 18972 8296 19012 8336
rect 19054 8296 19094 8336
rect 19136 8296 19176 8336
rect 33928 8296 33968 8336
rect 34010 8296 34050 8336
rect 34092 8296 34132 8336
rect 34174 8296 34214 8336
rect 34256 8296 34296 8336
rect 16828 8128 16868 8168
rect 17980 8128 18020 8168
rect 28060 8128 28100 8168
rect 28828 8128 28868 8168
rect 24988 8044 25028 8084
rect 16204 7960 16244 8000
rect 16588 7960 16628 8000
rect 16972 7960 17012 8000
rect 17356 7960 17396 8000
rect 17740 7960 17780 8000
rect 18412 7960 18452 8000
rect 18796 7960 18836 8000
rect 24748 7960 24788 8000
rect 25420 7960 25460 8000
rect 26284 7960 26324 8000
rect 27820 7960 27860 8000
rect 28588 7960 28628 8000
rect 44524 7960 44564 8000
rect 44908 7960 44948 8000
rect 26524 7792 26564 7832
rect 44764 7792 44804 7832
rect 16444 7708 16484 7748
rect 17212 7708 17252 7748
rect 17596 7708 17636 7748
rect 18652 7708 18692 7748
rect 19036 7708 19076 7748
rect 25660 7708 25700 7748
rect 45148 7708 45188 7748
rect 4928 7540 4968 7580
rect 5010 7540 5050 7580
rect 5092 7540 5132 7580
rect 5174 7540 5214 7580
rect 5256 7540 5296 7580
rect 20048 7540 20088 7580
rect 20130 7540 20170 7580
rect 20212 7540 20252 7580
rect 20294 7540 20334 7580
rect 20376 7540 20416 7580
rect 35168 7540 35208 7580
rect 35250 7540 35290 7580
rect 35332 7540 35372 7580
rect 35414 7540 35454 7580
rect 35496 7540 35536 7580
rect 12460 7120 12500 7160
rect 13900 7120 13940 7160
rect 14956 7120 14996 7160
rect 16108 7120 16148 7160
rect 16876 7120 16916 7160
rect 17356 7120 17396 7160
rect 17740 7120 17780 7160
rect 18124 7120 18164 7160
rect 18508 7120 18548 7160
rect 18892 7120 18932 7160
rect 19276 7120 19316 7160
rect 19660 7120 19700 7160
rect 20044 7120 20084 7160
rect 20428 7120 20468 7160
rect 20812 7120 20852 7160
rect 21052 7120 21092 7160
rect 21196 7120 21236 7160
rect 44524 7120 44564 7160
rect 44908 7120 44948 7160
rect 45148 7120 45188 7160
rect 18748 7036 18788 7076
rect 20668 7036 20708 7076
rect 12700 6952 12740 6992
rect 14140 6952 14180 6992
rect 15196 6952 15236 6992
rect 16348 6952 16388 6992
rect 17116 6952 17156 6992
rect 17596 6952 17636 6992
rect 17980 6952 18020 6992
rect 18364 6952 18404 6992
rect 19132 6952 19172 6992
rect 19516 6952 19556 6992
rect 19900 6952 19940 6992
rect 20284 6952 20324 6992
rect 21436 6952 21476 6992
rect 44764 6952 44804 6992
rect 3688 6784 3728 6824
rect 3770 6784 3810 6824
rect 3852 6784 3892 6824
rect 3934 6784 3974 6824
rect 4016 6784 4056 6824
rect 18808 6784 18848 6824
rect 18890 6784 18930 6824
rect 18972 6784 19012 6824
rect 19054 6784 19094 6824
rect 19136 6784 19176 6824
rect 33928 6784 33968 6824
rect 34010 6784 34050 6824
rect 34092 6784 34132 6824
rect 34174 6784 34214 6824
rect 34256 6784 34296 6824
rect 28348 6616 28388 6656
rect 20188 6532 20228 6572
rect 10828 6448 10868 6488
rect 19948 6448 19988 6488
rect 20380 6448 20420 6488
rect 28108 6448 28148 6488
rect 33196 6448 33236 6488
rect 44524 6448 44564 6488
rect 44908 6448 44948 6488
rect 45148 6448 45188 6488
rect 11068 6196 11108 6236
rect 20668 6196 20708 6236
rect 33436 6196 33476 6236
rect 44764 6196 44804 6236
rect 4928 6028 4968 6068
rect 5010 6028 5050 6068
rect 5092 6028 5132 6068
rect 5174 6028 5214 6068
rect 5256 6028 5296 6068
rect 20048 6028 20088 6068
rect 20130 6028 20170 6068
rect 20212 6028 20252 6068
rect 20294 6028 20334 6068
rect 20376 6028 20416 6068
rect 35168 6028 35208 6068
rect 35250 6028 35290 6068
rect 35332 6028 35372 6068
rect 35414 6028 35454 6068
rect 35496 6028 35536 6068
rect 11740 5860 11780 5900
rect 12508 5776 12548 5816
rect 45148 5776 45188 5816
rect 6700 5608 6740 5648
rect 7564 5608 7604 5648
rect 8716 5608 8756 5648
rect 8956 5608 8996 5648
rect 9868 5608 9908 5648
rect 10828 5608 10868 5648
rect 11500 5608 11540 5648
rect 12268 5608 12308 5648
rect 13516 5608 13556 5648
rect 21004 5608 21044 5648
rect 21388 5608 21428 5648
rect 21772 5608 21812 5648
rect 22012 5608 22052 5648
rect 34156 5608 34196 5648
rect 36940 5608 36980 5648
rect 37516 5608 37556 5648
rect 37900 5608 37940 5648
rect 38092 5608 38132 5648
rect 38476 5608 38516 5648
rect 38716 5608 38756 5648
rect 44524 5608 44564 5648
rect 44908 5608 44948 5648
rect 6940 5524 6980 5564
rect 10108 5524 10148 5564
rect 21628 5524 21668 5564
rect 38332 5524 38372 5564
rect 44764 5524 44804 5564
rect 7804 5440 7844 5480
rect 11068 5440 11108 5480
rect 13756 5440 13796 5480
rect 21244 5440 21284 5480
rect 34396 5440 34436 5480
rect 37180 5440 37220 5480
rect 3688 5272 3728 5312
rect 3770 5272 3810 5312
rect 3852 5272 3892 5312
rect 3934 5272 3974 5312
rect 4016 5272 4056 5312
rect 18808 5272 18848 5312
rect 18890 5272 18930 5312
rect 18972 5272 19012 5312
rect 19054 5272 19094 5312
rect 19136 5272 19176 5312
rect 33928 5272 33968 5312
rect 34010 5272 34050 5312
rect 34092 5272 34132 5312
rect 34174 5272 34214 5312
rect 34256 5272 34296 5312
rect 38908 5104 38948 5144
rect 45148 5104 45188 5144
rect 28348 5020 28388 5060
rect 41020 5020 41060 5060
rect 7180 4936 7220 4976
rect 7420 4936 7460 4976
rect 7564 4936 7604 4976
rect 8332 4936 8372 4976
rect 22060 4936 22100 4976
rect 22300 4936 22340 4976
rect 22483 4936 22523 4976
rect 22924 4936 22964 4976
rect 23404 4936 23444 4976
rect 26860 4936 26900 4976
rect 27724 4936 27764 4976
rect 28108 4936 28148 4976
rect 28492 4936 28532 4976
rect 34156 4936 34196 4976
rect 34444 4936 34484 4976
rect 38668 4936 38708 4976
rect 39628 4936 39668 4976
rect 40492 4936 40532 4976
rect 40780 4936 40820 4976
rect 41164 4936 41204 4976
rect 44524 4936 44564 4976
rect 44908 4936 44948 4976
rect 40108 4852 40148 4892
rect 41548 4852 41588 4892
rect 41836 4852 41876 4892
rect 27964 4768 28004 4808
rect 39868 4768 39908 4808
rect 41404 4768 41444 4808
rect 44764 4768 44804 4808
rect 7804 4684 7844 4724
rect 8572 4684 8612 4724
rect 22684 4684 22724 4724
rect 23164 4684 23204 4724
rect 23644 4684 23684 4724
rect 27100 4684 27140 4724
rect 28732 4684 28772 4724
rect 37699 4684 37739 4724
rect 38371 4684 38411 4724
rect 39043 4684 39083 4724
rect 39331 4684 39371 4724
rect 40099 4684 40139 4724
rect 40483 4684 40523 4724
rect 41827 4684 41867 4724
rect 4928 4516 4968 4556
rect 5010 4516 5050 4556
rect 5092 4516 5132 4556
rect 5174 4516 5214 4556
rect 5256 4516 5296 4556
rect 20048 4516 20088 4556
rect 20130 4516 20170 4556
rect 20212 4516 20252 4556
rect 20294 4516 20334 4556
rect 20376 4516 20416 4556
rect 35168 4516 35208 4556
rect 35250 4516 35290 4556
rect 35332 4516 35372 4556
rect 35414 4516 35454 4556
rect 35496 4516 35536 4556
rect 39331 4348 39371 4388
rect 40003 4348 40043 4388
rect 40483 4348 40523 4388
rect 40771 4348 40811 4388
rect 41059 4348 41099 4388
rect 41347 4348 41387 4388
rect 41635 4348 41675 4388
rect 42211 4348 42251 4388
rect 42787 4348 42827 4388
rect 41932 4264 41972 4304
rect 42508 4264 42548 4304
rect 45148 4264 45188 4304
rect 7084 4096 7124 4136
rect 23980 4096 24020 4136
rect 24460 4096 24500 4136
rect 25324 4096 25364 4136
rect 25564 4096 25604 4136
rect 26188 4096 26228 4136
rect 26428 4096 26468 4136
rect 27628 4096 27668 4136
rect 27868 4096 27908 4136
rect 32620 4096 32660 4136
rect 32860 4096 32900 4136
rect 44140 4096 44180 4136
rect 44524 4096 44564 4136
rect 44908 4096 44948 4136
rect 24700 4012 24740 4052
rect 44764 4012 44804 4052
rect 7324 3928 7364 3968
rect 24220 3928 24260 3968
rect 44380 3928 44420 3968
rect 3688 3760 3728 3800
rect 3770 3760 3810 3800
rect 3852 3760 3892 3800
rect 3934 3760 3974 3800
rect 4016 3760 4056 3800
rect 18808 3760 18848 3800
rect 18890 3760 18930 3800
rect 18972 3760 19012 3800
rect 19054 3760 19094 3800
rect 19136 3760 19176 3800
rect 33928 3760 33968 3800
rect 34010 3760 34050 3800
rect 34092 3760 34132 3800
rect 34174 3760 34214 3800
rect 34256 3760 34296 3800
rect 26908 3592 26948 3632
rect 27292 3592 27332 3632
rect 27676 3592 27716 3632
rect 30940 3592 30980 3632
rect 38140 3592 38180 3632
rect 45148 3592 45188 3632
rect 25900 3424 25940 3464
rect 26284 3424 26324 3464
rect 26668 3424 26708 3464
rect 27052 3424 27092 3464
rect 27436 3424 27476 3464
rect 27820 3424 27860 3464
rect 28204 3424 28244 3464
rect 28444 3424 28484 3464
rect 30028 3424 30068 3464
rect 30700 3424 30740 3464
rect 34828 3424 34868 3464
rect 35068 3424 35108 3464
rect 36556 3424 36596 3464
rect 37900 3424 37940 3464
rect 44524 3424 44564 3464
rect 44908 3424 44948 3464
rect 30268 3256 30308 3296
rect 36796 3256 36836 3296
rect 26140 3172 26180 3212
rect 26524 3172 26564 3212
rect 28060 3172 28100 3212
rect 44764 3172 44804 3212
rect 4928 3004 4968 3044
rect 5010 3004 5050 3044
rect 5092 3004 5132 3044
rect 5174 3004 5214 3044
rect 5256 3004 5296 3044
rect 20048 3004 20088 3044
rect 20130 3004 20170 3044
rect 20212 3004 20252 3044
rect 20294 3004 20334 3044
rect 20376 3004 20416 3044
rect 35168 3004 35208 3044
rect 35250 3004 35290 3044
rect 35332 3004 35372 3044
rect 35414 3004 35454 3044
rect 35496 3004 35536 3044
rect 34828 2836 34868 2876
rect 35107 2836 35147 2876
rect 45148 2752 45188 2792
rect 21484 2584 21524 2624
rect 21868 2584 21908 2624
rect 22252 2584 22292 2624
rect 22636 2584 22676 2624
rect 23020 2584 23060 2624
rect 23404 2584 23444 2624
rect 23788 2584 23828 2624
rect 25516 2584 25556 2624
rect 25900 2584 25940 2624
rect 26284 2584 26324 2624
rect 26668 2584 26708 2624
rect 27052 2584 27092 2624
rect 27436 2584 27476 2624
rect 27820 2584 27860 2624
rect 28204 2584 28244 2624
rect 28588 2584 28628 2624
rect 28972 2584 29012 2624
rect 29356 2584 29396 2624
rect 29740 2584 29780 2624
rect 30124 2584 30164 2624
rect 30508 2584 30548 2624
rect 30892 2584 30932 2624
rect 31276 2584 31316 2624
rect 44140 2584 44180 2624
rect 44524 2584 44564 2624
rect 44908 2584 44948 2624
rect 44764 2500 44804 2540
rect 21244 2416 21284 2456
rect 21628 2416 21668 2456
rect 22012 2416 22052 2456
rect 22396 2416 22436 2456
rect 22780 2416 22820 2456
rect 23164 2416 23204 2456
rect 23548 2416 23588 2456
rect 25276 2416 25316 2456
rect 25660 2416 25700 2456
rect 26044 2416 26084 2456
rect 26428 2416 26468 2456
rect 26812 2416 26852 2456
rect 27196 2416 27236 2456
rect 27580 2416 27620 2456
rect 27964 2416 28004 2456
rect 28348 2416 28388 2456
rect 28732 2416 28772 2456
rect 29116 2416 29156 2456
rect 29500 2416 29540 2456
rect 29884 2416 29924 2456
rect 30268 2416 30308 2456
rect 30652 2416 30692 2456
rect 31036 2416 31076 2456
rect 44380 2416 44420 2456
rect 3688 2248 3728 2288
rect 3770 2248 3810 2288
rect 3852 2248 3892 2288
rect 3934 2248 3974 2288
rect 4016 2248 4056 2288
rect 18808 2248 18848 2288
rect 18890 2248 18930 2288
rect 18972 2248 19012 2288
rect 19054 2248 19094 2288
rect 19136 2248 19176 2288
rect 33928 2248 33968 2288
rect 34010 2248 34050 2288
rect 34092 2248 34132 2288
rect 34174 2248 34214 2288
rect 34256 2248 34296 2288
rect 45148 2080 45188 2120
rect 27004 1996 27044 2036
rect 30076 1996 30116 2036
rect 20908 1912 20948 1952
rect 21292 1912 21332 1952
rect 21676 1912 21716 1952
rect 22060 1912 22100 1952
rect 22444 1912 22484 1952
rect 22828 1912 22868 1952
rect 23212 1912 23252 1952
rect 23596 1912 23636 1952
rect 23980 1912 24020 1952
rect 24556 1912 24596 1952
rect 24940 1912 24980 1952
rect 25324 1912 25364 1952
rect 25708 1912 25748 1952
rect 26092 1912 26132 1952
rect 26476 1912 26516 1952
rect 26860 1912 26900 1952
rect 27244 1912 27284 1952
rect 27628 1912 27668 1952
rect 28012 1912 28052 1952
rect 28396 1912 28436 1952
rect 28780 1912 28820 1952
rect 29164 1912 29204 1952
rect 29548 1912 29588 1952
rect 29932 1912 29972 1952
rect 30316 1912 30356 1952
rect 30700 1912 30740 1952
rect 31084 1912 31124 1952
rect 31468 1912 31508 1952
rect 31852 1912 31892 1952
rect 43756 1912 43796 1952
rect 44140 1912 44180 1952
rect 44524 1912 44564 1952
rect 44908 1912 44948 1952
rect 24220 1744 24260 1784
rect 25084 1744 25124 1784
rect 26236 1744 26276 1784
rect 27772 1744 27812 1784
rect 28924 1744 28964 1784
rect 30844 1744 30884 1784
rect 43996 1744 44036 1784
rect 44764 1744 44804 1784
rect 21148 1660 21188 1700
rect 21532 1660 21572 1700
rect 21916 1660 21956 1700
rect 22300 1660 22340 1700
rect 22684 1660 22724 1700
rect 23068 1660 23108 1700
rect 23452 1660 23492 1700
rect 23836 1660 23876 1700
rect 24316 1660 24356 1700
rect 24700 1660 24740 1700
rect 25468 1660 25508 1700
rect 25852 1660 25892 1700
rect 26620 1660 26660 1700
rect 27388 1660 27428 1700
rect 28156 1660 28196 1700
rect 28540 1660 28580 1700
rect 29308 1660 29348 1700
rect 29692 1660 29732 1700
rect 30460 1660 30500 1700
rect 31228 1660 31268 1700
rect 31612 1660 31652 1700
rect 44380 1660 44420 1700
rect 4928 1492 4968 1532
rect 5010 1492 5050 1532
rect 5092 1492 5132 1532
rect 5174 1492 5214 1532
rect 5256 1492 5296 1532
rect 20048 1492 20088 1532
rect 20130 1492 20170 1532
rect 20212 1492 20252 1532
rect 20294 1492 20334 1532
rect 20376 1492 20416 1532
rect 35168 1492 35208 1532
rect 35250 1492 35290 1532
rect 35332 1492 35372 1532
rect 35414 1492 35454 1532
rect 35496 1492 35536 1532
<< metal2 >>
rect 0 11192 90 11212
rect 46278 11192 46368 11212
rect 0 11152 364 11192
rect 404 11152 413 11192
rect 44035 11152 44044 11192
rect 44084 11152 46368 11192
rect 0 11132 90 11152
rect 46278 11132 46368 11152
rect 2860 10900 21484 10940
rect 21524 10900 21533 10940
rect 0 10856 90 10876
rect 2860 10856 2900 10900
rect 46278 10856 46368 10876
rect 0 10816 2900 10856
rect 16972 10816 21292 10856
rect 21332 10816 21341 10856
rect 26371 10816 26380 10856
rect 26420 10816 42412 10856
rect 42452 10816 42461 10856
rect 44140 10816 46368 10856
rect 0 10796 90 10816
rect 4919 10564 4928 10604
rect 4968 10564 5010 10604
rect 5050 10564 5092 10604
rect 5132 10564 5174 10604
rect 5214 10564 5256 10604
rect 5296 10564 5305 10604
rect 0 10520 90 10540
rect 16972 10520 17012 10816
rect 17059 10732 17068 10772
rect 17108 10732 31180 10772
rect 31220 10732 31229 10772
rect 19171 10648 19180 10688
rect 19220 10648 31468 10688
rect 31508 10648 31517 10688
rect 32044 10648 40204 10688
rect 40244 10648 40253 10688
rect 32044 10604 32084 10648
rect 20039 10564 20048 10604
rect 20088 10564 20130 10604
rect 20170 10564 20212 10604
rect 20252 10564 20294 10604
rect 20334 10564 20376 10604
rect 20416 10564 20425 10604
rect 26755 10564 26764 10604
rect 26804 10564 32084 10604
rect 35159 10564 35168 10604
rect 35208 10564 35250 10604
rect 35290 10564 35332 10604
rect 35372 10564 35414 10604
rect 35454 10564 35496 10604
rect 35536 10564 35545 10604
rect 0 10480 17012 10520
rect 23491 10480 23500 10520
rect 23540 10480 30220 10520
rect 30260 10480 30269 10520
rect 40291 10480 40300 10520
rect 40340 10480 43180 10520
rect 43220 10480 43229 10520
rect 0 10460 90 10480
rect 44140 10436 44180 10816
rect 46278 10796 46368 10816
rect 46278 10520 46368 10540
rect 44419 10480 44428 10520
rect 44468 10480 46368 10520
rect 46278 10460 46368 10480
rect 1987 10396 1996 10436
rect 2036 10396 2044 10436
rect 2084 10396 2167 10436
rect 4099 10396 4108 10436
rect 4148 10396 4156 10436
rect 4196 10396 4279 10436
rect 6211 10396 6220 10436
rect 6260 10396 6268 10436
rect 6308 10396 6391 10436
rect 8323 10396 8332 10436
rect 8372 10396 8380 10436
rect 8420 10396 8503 10436
rect 10435 10396 10444 10436
rect 10484 10396 10492 10436
rect 10532 10396 10615 10436
rect 12547 10396 12556 10436
rect 12596 10396 12604 10436
rect 12644 10396 12727 10436
rect 14659 10396 14668 10436
rect 14708 10396 14716 10436
rect 14756 10396 14839 10436
rect 16771 10396 16780 10436
rect 16820 10396 16828 10436
rect 16868 10396 16951 10436
rect 18883 10396 18892 10436
rect 18932 10396 18940 10436
rect 18980 10396 19063 10436
rect 20995 10396 21004 10436
rect 21044 10396 21052 10436
rect 21092 10396 21175 10436
rect 23107 10396 23116 10436
rect 23156 10396 23164 10436
rect 23204 10396 23287 10436
rect 25219 10396 25228 10436
rect 25268 10396 25276 10436
rect 25316 10396 25399 10436
rect 27331 10396 27340 10436
rect 27380 10396 27388 10436
rect 27428 10396 27511 10436
rect 29443 10396 29452 10436
rect 29492 10396 29500 10436
rect 29540 10396 29623 10436
rect 31555 10396 31564 10436
rect 31604 10396 31612 10436
rect 31652 10396 31735 10436
rect 33667 10396 33676 10436
rect 33716 10396 33724 10436
rect 33764 10396 33847 10436
rect 35779 10396 35788 10436
rect 35828 10396 35836 10436
rect 35876 10396 35959 10436
rect 37891 10396 37900 10436
rect 37940 10396 37948 10436
rect 37988 10396 38071 10436
rect 40003 10396 40012 10436
rect 40052 10396 40060 10436
rect 40100 10396 40183 10436
rect 42115 10396 42124 10436
rect 42164 10396 42172 10436
rect 42212 10396 42295 10436
rect 43411 10396 43420 10436
rect 43460 10396 44180 10436
rect 44227 10396 44236 10436
rect 44276 10396 44284 10436
rect 44324 10396 44407 10436
rect 172 10312 20524 10352
rect 20564 10312 20573 10352
rect 23299 10312 23308 10352
rect 23348 10312 25900 10352
rect 25940 10312 25949 10352
rect 28387 10312 28396 10352
rect 28436 10312 32084 10352
rect 0 10184 90 10204
rect 172 10184 212 10312
rect 32044 10268 32084 10312
rect 12940 10228 16972 10268
rect 17012 10228 17021 10268
rect 19276 10228 25036 10268
rect 25076 10228 25085 10268
rect 28867 10228 28876 10268
rect 28916 10228 31988 10268
rect 32044 10228 38324 10268
rect 12940 10184 12980 10228
rect 0 10144 212 10184
rect 2275 10144 2284 10184
rect 2324 10144 2333 10184
rect 4387 10144 4396 10184
rect 4436 10144 6220 10184
rect 6260 10144 6269 10184
rect 6377 10144 6508 10184
rect 6548 10144 6557 10184
rect 8489 10144 8620 10184
rect 8660 10144 8669 10184
rect 10723 10144 10732 10184
rect 10772 10144 10781 10184
rect 12835 10144 12844 10184
rect 12884 10144 12980 10184
rect 14947 10144 14956 10184
rect 14996 10144 15005 10184
rect 16937 10144 17068 10184
rect 17108 10144 17117 10184
rect 19049 10144 19180 10184
rect 19220 10144 19229 10184
rect 0 10124 90 10144
rect 2284 10100 2324 10144
rect 10732 10100 10772 10144
rect 14956 10100 14996 10144
rect 19276 10100 19316 10228
rect 31948 10184 31988 10228
rect 21283 10144 21292 10184
rect 21332 10144 23308 10184
rect 23348 10144 23357 10184
rect 23443 10144 23452 10184
rect 23492 10144 23540 10184
rect 25507 10144 25516 10184
rect 25556 10144 27244 10184
rect 27284 10144 27293 10184
rect 27497 10144 27628 10184
rect 27668 10144 27677 10184
rect 28771 10144 28780 10184
rect 28820 10144 29740 10184
rect 29780 10144 29789 10184
rect 31843 10144 31852 10184
rect 31892 10144 31901 10184
rect 31948 10144 33964 10184
rect 34004 10144 34013 10184
rect 34531 10144 34540 10184
rect 34580 10144 36076 10184
rect 36116 10144 36125 10184
rect 38179 10144 38188 10184
rect 38228 10144 38237 10184
rect 2284 10060 7180 10100
rect 7220 10060 7229 10100
rect 10732 10060 13036 10100
rect 13076 10060 13085 10100
rect 14956 10060 19316 10100
rect 23500 10100 23540 10144
rect 31852 10100 31892 10144
rect 38188 10100 38228 10144
rect 23500 10060 26860 10100
rect 26900 10060 26909 10100
rect 28099 10060 28108 10100
rect 28148 10060 31892 10100
rect 35587 10060 35596 10100
rect 35636 10060 38228 10100
rect 38284 10100 38324 10228
rect 46278 10184 46368 10204
rect 40169 10144 40204 10184
rect 40244 10144 40300 10184
rect 40340 10144 40349 10184
rect 42281 10144 42412 10184
rect 42452 10144 42461 10184
rect 43049 10144 43180 10184
rect 43220 10144 43229 10184
rect 43433 10144 43564 10184
rect 43604 10144 43613 10184
rect 43817 10144 43948 10184
rect 43988 10144 43997 10184
rect 44393 10144 44524 10184
rect 44564 10144 44573 10184
rect 44777 10144 44908 10184
rect 44948 10144 44957 10184
rect 45100 10144 46368 10184
rect 45100 10100 45140 10144
rect 46278 10124 46368 10144
rect 38284 10060 40396 10100
rect 40436 10060 40445 10100
rect 43795 10060 43804 10100
rect 43844 10060 45140 10100
rect 24547 9976 24556 10016
rect 24596 9976 33140 10016
rect 44179 9976 44188 10016
rect 44228 9976 45044 10016
rect 45139 9976 45148 10016
rect 45188 9976 45772 10016
rect 45812 9976 45821 10016
rect 33100 9932 33140 9976
rect 1315 9892 1324 9932
rect 1364 9892 27724 9932
rect 27764 9892 27773 9932
rect 27907 9892 27916 9932
rect 27956 9892 32140 9932
rect 32180 9892 32189 9932
rect 33100 9892 44948 9932
rect 0 9848 90 9868
rect 0 9808 2900 9848
rect 3679 9808 3688 9848
rect 3728 9808 3770 9848
rect 3810 9808 3852 9848
rect 3892 9808 3934 9848
rect 3974 9808 4016 9848
rect 4056 9808 4065 9848
rect 18799 9808 18808 9848
rect 18848 9808 18890 9848
rect 18930 9808 18972 9848
rect 19012 9808 19054 9848
rect 19094 9808 19136 9848
rect 19176 9808 19185 9848
rect 23107 9808 23116 9848
rect 23156 9808 30796 9848
rect 30836 9808 30845 9848
rect 33919 9808 33928 9848
rect 33968 9808 34010 9848
rect 34050 9808 34092 9848
rect 34132 9808 34174 9848
rect 34214 9808 34256 9848
rect 34296 9808 34305 9848
rect 0 9788 90 9808
rect 2860 9764 2900 9808
rect 2860 9724 22444 9764
rect 22484 9724 22493 9764
rect 27139 9724 27148 9764
rect 27188 9724 33100 9764
rect 33140 9724 33149 9764
rect 30211 9640 30220 9680
rect 30260 9640 44180 9680
rect 44297 9640 44380 9680
rect 44420 9640 44428 9680
rect 44468 9640 44477 9680
rect 23203 9556 23212 9596
rect 23252 9556 38092 9596
rect 38132 9556 38141 9596
rect 43913 9556 43996 9596
rect 44036 9556 44044 9596
rect 44084 9556 44093 9596
rect 0 9512 90 9532
rect 44140 9512 44180 9640
rect 44908 9512 44948 9892
rect 45004 9848 45044 9976
rect 46278 9848 46368 9868
rect 45004 9808 46368 9848
rect 46278 9788 46368 9808
rect 46278 9512 46368 9532
rect 0 9472 1228 9512
rect 1268 9472 1277 9512
rect 22627 9472 22636 9512
rect 22676 9472 30604 9512
rect 30644 9472 30653 9512
rect 30883 9472 30892 9512
rect 30932 9472 33484 9512
rect 33524 9472 33533 9512
rect 43625 9472 43756 9512
rect 43796 9472 43805 9512
rect 44131 9472 44140 9512
rect 44180 9472 44189 9512
rect 44515 9472 44524 9512
rect 44564 9472 44573 9512
rect 44899 9472 44908 9512
rect 44948 9472 44957 9512
rect 45763 9472 45772 9512
rect 45812 9472 46368 9512
rect 0 9452 90 9472
rect 18979 9388 18988 9428
rect 19028 9388 27916 9428
rect 27956 9388 27965 9428
rect 28291 9388 28300 9428
rect 28340 9388 33772 9428
rect 33812 9388 33821 9428
rect 38092 9388 43564 9428
rect 43604 9388 43613 9428
rect 38092 9344 38132 9388
rect 44524 9344 44564 9472
rect 46278 9452 46368 9472
rect 25891 9304 25900 9344
rect 25940 9304 29068 9344
rect 29108 9304 29117 9344
rect 30787 9304 30796 9344
rect 30836 9304 38132 9344
rect 38179 9304 38188 9344
rect 38228 9304 44564 9344
rect 28003 9220 28012 9260
rect 28052 9220 37996 9260
rect 38036 9220 38045 9260
rect 44755 9220 44764 9260
rect 44804 9220 44813 9260
rect 45139 9220 45148 9260
rect 45188 9220 45772 9260
rect 45812 9220 45821 9260
rect 0 9176 90 9196
rect 44764 9176 44804 9220
rect 46278 9176 46368 9196
rect 0 9136 23596 9176
rect 23636 9136 23645 9176
rect 26083 9136 26092 9176
rect 26132 9136 32332 9176
rect 32372 9136 32381 9176
rect 33100 9136 38036 9176
rect 44764 9136 46368 9176
rect 0 9116 90 9136
rect 33100 9092 33140 9136
rect 37996 9092 38036 9136
rect 46278 9116 46368 9136
rect 4919 9052 4928 9092
rect 4968 9052 5010 9092
rect 5050 9052 5092 9092
rect 5132 9052 5174 9092
rect 5214 9052 5256 9092
rect 5296 9052 5305 9092
rect 20039 9052 20048 9092
rect 20088 9052 20130 9092
rect 20170 9052 20212 9092
rect 20252 9052 20294 9092
rect 20334 9052 20376 9092
rect 20416 9052 20425 9092
rect 20515 9052 20524 9092
rect 20564 9052 22924 9092
rect 22964 9052 22973 9092
rect 23692 9052 33140 9092
rect 35159 9052 35168 9092
rect 35208 9052 35250 9092
rect 35290 9052 35332 9092
rect 35372 9052 35414 9092
rect 35454 9052 35496 9092
rect 35536 9052 35545 9092
rect 37996 9052 38324 9092
rect 22636 8968 23500 9008
rect 23540 8968 23549 9008
rect 22636 8924 22676 8968
rect 23692 8924 23732 9052
rect 38284 9008 38324 9052
rect 24940 8968 38188 9008
rect 38228 8968 38237 9008
rect 38284 8968 44524 9008
rect 44564 8968 44573 9008
rect 24940 8924 24980 8968
rect 6163 8884 6172 8924
rect 6212 8884 6508 8924
rect 6548 8884 6557 8924
rect 7171 8884 7180 8924
rect 7220 8884 8572 8924
rect 8612 8884 8621 8924
rect 13027 8884 13036 8924
rect 13076 8884 13084 8924
rect 13124 8884 13207 8924
rect 16963 8884 16972 8924
rect 17012 8884 18748 8924
rect 18788 8884 18797 8924
rect 21523 8884 21532 8924
rect 21572 8884 22156 8924
rect 22196 8884 22205 8924
rect 22291 8884 22300 8924
rect 22340 8884 22676 8924
rect 23059 8884 23068 8924
rect 23108 8884 23116 8924
rect 23156 8884 23239 8924
rect 23443 8884 23452 8924
rect 23492 8884 23732 8924
rect 23827 8884 23836 8924
rect 23876 8884 24980 8924
rect 25027 8884 25036 8924
rect 25076 8884 25852 8924
rect 25892 8884 25901 8924
rect 26851 8884 26860 8924
rect 26900 8884 26908 8924
rect 26948 8884 27031 8924
rect 27235 8884 27244 8924
rect 27284 8884 27292 8924
rect 27332 8884 27415 8924
rect 27619 8884 27628 8924
rect 27668 8884 28060 8924
rect 28100 8884 28109 8924
rect 28649 8884 28732 8924
rect 28772 8884 28780 8924
rect 28820 8884 28829 8924
rect 29059 8884 29068 8924
rect 29108 8884 29116 8924
rect 29156 8884 29239 8924
rect 30595 8884 30604 8924
rect 30644 8884 43948 8924
rect 43988 8884 43997 8924
rect 0 8840 90 8860
rect 46278 8840 46368 8860
rect 0 8800 76 8840
rect 116 8800 125 8840
rect 10051 8800 10060 8840
rect 10100 8800 24212 8840
rect 24403 8800 24412 8840
rect 24452 8800 24556 8840
rect 24596 8800 24605 8840
rect 27881 8800 27964 8840
rect 28004 8800 28012 8840
rect 28052 8800 28061 8840
rect 28396 8800 30892 8840
rect 30932 8800 30941 8840
rect 31171 8800 31180 8840
rect 31220 8800 31228 8840
rect 31268 8800 31351 8840
rect 45763 8800 45772 8840
rect 45812 8800 46368 8840
rect 0 8780 90 8800
rect 6211 8716 6220 8756
rect 6260 8716 6548 8756
rect 6508 8672 6548 8716
rect 8140 8716 8620 8756
rect 8660 8716 8669 8756
rect 8899 8716 8908 8756
rect 8948 8716 23060 8756
rect 8140 8672 8180 8716
rect 23020 8672 23060 8716
rect 24172 8672 24212 8800
rect 28396 8756 28436 8800
rect 46278 8780 46368 8800
rect 27532 8716 28436 8756
rect 28492 8716 33140 8756
rect 37987 8716 37996 8756
rect 38036 8716 44948 8756
rect 27532 8672 27572 8716
rect 28492 8672 28532 8716
rect 33100 8672 33140 8716
rect 44908 8672 44948 8716
rect 6281 8632 6412 8672
rect 6452 8632 6461 8672
rect 6508 8632 6652 8672
rect 6692 8632 6701 8672
rect 6761 8632 6892 8672
rect 6932 8632 6941 8672
rect 7337 8632 7468 8672
rect 7508 8632 7517 8672
rect 7699 8632 7708 8672
rect 7748 8632 8180 8672
rect 8681 8632 8812 8672
rect 8852 8632 8861 8672
rect 13315 8632 13324 8672
rect 13364 8632 14380 8672
rect 14420 8632 14429 8672
rect 18857 8632 18988 8672
rect 19028 8632 19037 8672
rect 21161 8632 21292 8672
rect 21332 8632 21341 8672
rect 21580 8632 21676 8672
rect 21716 8632 21725 8672
rect 21859 8632 21868 8672
rect 21908 8632 22060 8672
rect 22100 8632 22109 8672
rect 22313 8632 22444 8672
rect 22484 8632 22493 8672
rect 22627 8632 22636 8672
rect 22676 8632 22685 8672
rect 22793 8632 22867 8672
rect 22907 8632 22924 8672
rect 22964 8632 22973 8672
rect 23020 8632 23212 8672
rect 23252 8632 23261 8672
rect 23465 8632 23596 8672
rect 23636 8632 23645 8672
rect 24163 8632 24172 8672
rect 24212 8632 24221 8672
rect 25961 8632 26092 8672
rect 26132 8632 26141 8672
rect 27017 8632 27148 8672
rect 27188 8632 27197 8672
rect 27523 8632 27532 8672
rect 27572 8632 27581 8672
rect 27715 8632 27724 8672
rect 27764 8632 27895 8672
rect 28169 8632 28300 8672
rect 28340 8632 28349 8672
rect 28483 8632 28492 8672
rect 28532 8632 28541 8672
rect 29347 8632 29356 8672
rect 29396 8632 31316 8672
rect 31459 8632 31468 8672
rect 31508 8632 31796 8672
rect 31843 8632 31852 8672
rect 31892 8632 32716 8672
rect 32756 8632 32765 8672
rect 33100 8632 33388 8672
rect 33428 8632 33437 8672
rect 38083 8632 38092 8672
rect 38132 8632 44524 8672
rect 44564 8632 44573 8672
rect 44899 8632 44908 8672
rect 44948 8632 44957 8672
rect 45139 8632 45148 8672
rect 45188 8632 46252 8672
rect 46292 8632 46301 8672
rect 2860 8548 12980 8588
rect 0 8504 90 8524
rect 2860 8504 2900 8548
rect 0 8464 2900 8504
rect 12940 8504 12980 8548
rect 21580 8504 21620 8632
rect 22636 8588 22676 8632
rect 22636 8548 22684 8588
rect 22724 8548 22733 8588
rect 31276 8504 31316 8632
rect 31756 8588 31796 8632
rect 31459 8548 31468 8588
rect 31508 8548 31612 8588
rect 31652 8548 31661 8588
rect 31756 8548 32524 8588
rect 32564 8548 32573 8588
rect 44755 8548 44764 8588
rect 44804 8548 45620 8588
rect 45580 8504 45620 8548
rect 46278 8504 46368 8524
rect 12940 8464 21620 8504
rect 21907 8464 21916 8504
rect 21956 8464 23212 8504
rect 23252 8464 23261 8504
rect 31276 8464 32908 8504
rect 32948 8464 32957 8504
rect 45580 8464 46368 8504
rect 0 8444 90 8464
rect 46278 8444 46368 8464
rect 355 8380 364 8420
rect 404 8380 26284 8420
rect 26324 8380 26333 8420
rect 3679 8296 3688 8336
rect 3728 8296 3770 8336
rect 3810 8296 3852 8336
rect 3892 8296 3934 8336
rect 3974 8296 4016 8336
rect 4056 8296 4065 8336
rect 15811 8296 15820 8336
rect 15860 8296 18604 8336
rect 18644 8296 18653 8336
rect 18799 8296 18808 8336
rect 18848 8296 18890 8336
rect 18930 8296 18972 8336
rect 19012 8296 19054 8336
rect 19094 8296 19136 8336
rect 19176 8296 19185 8336
rect 19276 8296 26036 8336
rect 33919 8296 33928 8336
rect 33968 8296 34010 8336
rect 34050 8296 34092 8336
rect 34132 8296 34174 8336
rect 34214 8296 34256 8336
rect 34296 8296 34305 8336
rect 19276 8252 19316 8296
rect 25996 8252 26036 8296
rect 15619 8212 15628 8252
rect 15668 8212 17740 8252
rect 17780 8212 17789 8252
rect 17836 8212 19316 8252
rect 20524 8212 25900 8252
rect 25940 8212 25949 8252
rect 25996 8212 28780 8252
rect 28820 8212 28829 8252
rect 0 8168 90 8188
rect 17836 8168 17876 8212
rect 20524 8168 20564 8212
rect 46278 8168 46368 8188
rect 0 8128 1324 8168
rect 1364 8128 1373 8168
rect 15235 8128 15244 8168
rect 15284 8128 16724 8168
rect 16819 8128 16828 8168
rect 16868 8128 17876 8168
rect 17971 8128 17980 8168
rect 18020 8128 20564 8168
rect 27977 8128 28060 8168
rect 28100 8128 28108 8168
rect 28148 8128 28157 8168
rect 28745 8128 28828 8168
rect 28868 8128 28876 8168
rect 28916 8128 28925 8168
rect 46243 8128 46252 8168
rect 46292 8128 46368 8168
rect 0 8108 90 8128
rect 1219 8044 1228 8084
rect 1268 8044 16588 8084
rect 16628 8044 16637 8084
rect 16684 8000 16724 8128
rect 46278 8108 46368 8128
rect 16771 8044 16780 8084
rect 16820 8044 23060 8084
rect 24979 8044 24988 8084
rect 25028 8044 26228 8084
rect 23020 8000 23060 8044
rect 14851 7960 14860 8000
rect 14900 7960 16204 8000
rect 16244 7960 16253 8000
rect 16579 7960 16588 8000
rect 16628 7960 16637 8000
rect 16684 7960 16972 8000
rect 17012 7960 17021 8000
rect 17225 7960 17356 8000
rect 17396 7960 17405 8000
rect 17609 7960 17740 8000
rect 17780 7960 17789 8000
rect 18403 7960 18412 8000
rect 18452 7960 18461 8000
rect 18595 7960 18604 8000
rect 18644 7960 18796 8000
rect 18836 7960 18845 8000
rect 23020 7960 24748 8000
rect 24788 7960 24797 8000
rect 25411 7960 25420 8000
rect 25460 7960 25469 8000
rect 16588 7916 16628 7960
rect 18412 7916 18452 7960
rect 15043 7876 15052 7916
rect 15092 7876 16628 7916
rect 16684 7876 18452 7916
rect 0 7832 90 7852
rect 16684 7832 16724 7876
rect 25420 7832 25460 7960
rect 26188 7916 26228 8044
rect 27724 8044 30988 8084
rect 31028 8044 31037 8084
rect 43948 8044 44908 8084
rect 44948 8044 44957 8084
rect 26275 7960 26284 8000
rect 26324 7960 26455 8000
rect 27724 7916 27764 8044
rect 27811 7960 27820 8000
rect 27860 7960 27869 8000
rect 28579 7960 28588 8000
rect 28628 7960 33580 8000
rect 33620 7960 33629 8000
rect 26188 7876 27764 7916
rect 0 7792 8908 7832
rect 8948 7792 8957 7832
rect 16003 7792 16012 7832
rect 16052 7792 16724 7832
rect 17932 7792 25460 7832
rect 26515 7792 26524 7832
rect 26564 7792 27724 7832
rect 27764 7792 27773 7832
rect 0 7772 90 7792
rect 16435 7708 16444 7748
rect 16484 7708 17068 7748
rect 17108 7708 17117 7748
rect 17203 7708 17212 7748
rect 17252 7708 17452 7748
rect 17492 7708 17501 7748
rect 17587 7708 17596 7748
rect 17636 7708 17836 7748
rect 17876 7708 17885 7748
rect 17932 7664 17972 7792
rect 27820 7748 27860 7960
rect 27907 7876 27916 7916
rect 27956 7876 43756 7916
rect 43796 7876 43805 7916
rect 43948 7832 43988 8044
rect 44393 7960 44524 8000
rect 44564 7960 44573 8000
rect 44899 7960 44908 8000
rect 44948 7960 44957 8000
rect 44908 7916 44948 7960
rect 30979 7792 30988 7832
rect 31028 7792 43988 7832
rect 44044 7876 44948 7916
rect 18643 7708 18652 7748
rect 18692 7708 18932 7748
rect 19027 7708 19036 7748
rect 19076 7708 25556 7748
rect 25651 7708 25660 7748
rect 25700 7708 26420 7748
rect 27820 7708 33676 7748
rect 33716 7708 33725 7748
rect 2860 7624 17972 7664
rect 18892 7664 18932 7708
rect 18892 7624 25420 7664
rect 25460 7624 25469 7664
rect 0 7496 90 7516
rect 2860 7496 2900 7624
rect 25516 7580 25556 7708
rect 26380 7664 26420 7708
rect 44044 7664 44084 7876
rect 46278 7832 46368 7852
rect 44755 7792 44764 7832
rect 44804 7792 46368 7832
rect 46278 7772 46368 7792
rect 45139 7708 45148 7748
rect 45188 7708 45197 7748
rect 26380 7624 44084 7664
rect 45148 7664 45188 7708
rect 45148 7624 46252 7664
rect 46292 7624 46301 7664
rect 4919 7540 4928 7580
rect 4968 7540 5010 7580
rect 5050 7540 5092 7580
rect 5132 7540 5174 7580
rect 5214 7540 5256 7580
rect 5296 7540 5305 7580
rect 20039 7540 20048 7580
rect 20088 7540 20130 7580
rect 20170 7540 20212 7580
rect 20252 7540 20294 7580
rect 20334 7540 20376 7580
rect 20416 7540 20425 7580
rect 25516 7540 26668 7580
rect 26708 7540 26717 7580
rect 35159 7540 35168 7580
rect 35208 7540 35250 7580
rect 35290 7540 35332 7580
rect 35372 7540 35414 7580
rect 35454 7540 35496 7580
rect 35536 7540 35545 7580
rect 46278 7496 46368 7516
rect 0 7456 2900 7496
rect 17827 7456 17836 7496
rect 17876 7456 26860 7496
rect 26900 7456 26909 7496
rect 46243 7456 46252 7496
rect 46292 7456 46368 7496
rect 0 7436 90 7456
rect 46278 7436 46368 7456
rect 17443 7372 17452 7412
rect 17492 7372 25516 7412
rect 25556 7372 25565 7412
rect 25891 7372 25900 7412
rect 25940 7372 27244 7412
rect 27284 7372 27293 7412
rect 17059 7288 17068 7328
rect 17108 7288 25228 7328
rect 25268 7288 25277 7328
rect 15427 7204 15436 7244
rect 15476 7204 17356 7244
rect 17396 7204 17405 7244
rect 21100 7204 21524 7244
rect 0 7160 90 7180
rect 21100 7160 21140 7204
rect 21484 7160 21524 7204
rect 46278 7160 46368 7180
rect 0 7120 1420 7160
rect 1460 7120 1469 7160
rect 12451 7120 12460 7160
rect 12500 7120 13516 7160
rect 13556 7120 13565 7160
rect 13699 7120 13708 7160
rect 13748 7120 13900 7160
rect 13940 7120 13949 7160
rect 14947 7120 14956 7160
rect 14996 7120 15005 7160
rect 15052 7120 16108 7160
rect 16148 7120 16157 7160
rect 16204 7120 16876 7160
rect 16916 7120 16925 7160
rect 17059 7120 17068 7160
rect 17108 7120 17356 7160
rect 17396 7120 17405 7160
rect 17609 7120 17740 7160
rect 17780 7120 17789 7160
rect 18115 7120 18124 7160
rect 18164 7120 18173 7160
rect 18499 7120 18508 7160
rect 18548 7120 18557 7160
rect 18691 7120 18700 7160
rect 18740 7120 18892 7160
rect 18932 7120 18941 7160
rect 19145 7120 19276 7160
rect 19316 7120 19325 7160
rect 19529 7120 19660 7160
rect 19700 7120 19709 7160
rect 19843 7120 19852 7160
rect 19892 7120 20044 7160
rect 20084 7120 20093 7160
rect 20227 7120 20236 7160
rect 20276 7120 20428 7160
rect 20468 7120 20477 7160
rect 20681 7120 20716 7160
rect 20756 7120 20812 7160
rect 20852 7120 20861 7160
rect 21043 7120 21052 7160
rect 21092 7120 21140 7160
rect 21187 7120 21196 7160
rect 21236 7120 21367 7160
rect 21484 7120 23980 7160
rect 24020 7120 24029 7160
rect 27331 7120 27340 7160
rect 27380 7120 44524 7160
rect 44564 7120 44573 7160
rect 44899 7120 44908 7160
rect 44948 7120 44957 7160
rect 45139 7120 45148 7160
rect 45188 7120 46368 7160
rect 0 7100 90 7120
rect 14956 7076 14996 7120
rect 13891 7036 13900 7076
rect 13940 7036 14996 7076
rect 12691 6952 12700 6992
rect 12740 6952 13940 6992
rect 0 6824 90 6844
rect 0 6784 1132 6824
rect 1172 6784 1181 6824
rect 3679 6784 3688 6824
rect 3728 6784 3770 6824
rect 3810 6784 3852 6824
rect 3892 6784 3934 6824
rect 3974 6784 4016 6824
rect 4056 6784 4065 6824
rect 0 6764 90 6784
rect 0 6488 90 6508
rect 0 6448 940 6488
rect 980 6448 989 6488
rect 10819 6448 10828 6488
rect 10868 6448 13324 6488
rect 13364 6448 13373 6488
rect 0 6428 90 6448
rect 13900 6236 13940 6952
rect 13996 6952 14140 6992
rect 14180 6952 14189 6992
rect 13996 6320 14036 6952
rect 15052 6908 15092 7120
rect 15187 6952 15196 6992
rect 15236 6952 16108 6992
rect 16148 6952 16157 6992
rect 14083 6868 14092 6908
rect 14132 6868 15092 6908
rect 16204 6824 16244 7120
rect 18124 7076 18164 7120
rect 18508 7076 18548 7120
rect 44908 7076 44948 7120
rect 46278 7100 46368 7120
rect 16291 7036 16300 7076
rect 16340 7036 18164 7076
rect 18211 7036 18220 7076
rect 18260 7036 18548 7076
rect 18739 7036 18748 7076
rect 18788 7036 20180 7076
rect 20659 7036 20668 7076
rect 20708 7036 23212 7076
rect 23252 7036 23261 7076
rect 43171 7036 43180 7076
rect 43220 7036 44948 7076
rect 16339 6952 16348 6992
rect 16388 6952 17012 6992
rect 17107 6952 17116 6992
rect 17156 6952 17452 6992
rect 17492 6952 17501 6992
rect 17587 6952 17596 6992
rect 17636 6952 17836 6992
rect 17876 6952 17885 6992
rect 17971 6952 17980 6992
rect 18020 6952 18124 6992
rect 18164 6952 18173 6992
rect 18355 6952 18364 6992
rect 18404 6952 18604 6992
rect 18644 6952 18653 6992
rect 19123 6952 19132 6992
rect 19172 6952 19372 6992
rect 19412 6952 19421 6992
rect 19507 6952 19516 6992
rect 19556 6952 19796 6992
rect 19891 6952 19900 6992
rect 19940 6952 19948 6992
rect 19988 6952 20071 6992
rect 16972 6908 17012 6952
rect 16972 6868 19700 6908
rect 14275 6784 14284 6824
rect 14324 6784 16244 6824
rect 16387 6784 16396 6824
rect 16436 6784 18220 6824
rect 18260 6784 18269 6824
rect 18799 6784 18808 6824
rect 18848 6784 18890 6824
rect 18930 6784 18972 6824
rect 19012 6784 19054 6824
rect 19094 6784 19136 6824
rect 19176 6784 19185 6824
rect 19660 6740 19700 6868
rect 19756 6824 19796 6952
rect 20140 6908 20180 7036
rect 20275 6952 20284 6992
rect 20324 6952 20948 6992
rect 21427 6952 21436 6992
rect 21476 6952 24268 6992
rect 24308 6952 24317 6992
rect 44755 6952 44764 6992
rect 44804 6952 46252 6992
rect 46292 6952 46301 6992
rect 20908 6908 20948 6952
rect 20140 6868 20812 6908
rect 20852 6868 20861 6908
rect 20908 6868 24172 6908
rect 24212 6868 24221 6908
rect 46278 6824 46368 6844
rect 19756 6784 25804 6824
rect 25844 6784 25853 6824
rect 33919 6784 33928 6824
rect 33968 6784 34010 6824
rect 34050 6784 34092 6824
rect 34132 6784 34174 6824
rect 34214 6784 34256 6824
rect 34296 6784 34305 6824
rect 46243 6784 46252 6824
rect 46292 6784 46368 6824
rect 46278 6764 46368 6784
rect 14467 6700 14476 6740
rect 14516 6700 17068 6740
rect 17108 6700 17117 6740
rect 17827 6700 17836 6740
rect 17876 6700 19316 6740
rect 19660 6700 23788 6740
rect 23828 6700 23837 6740
rect 16579 6616 16588 6656
rect 16628 6616 18700 6656
rect 18740 6616 18749 6656
rect 19276 6572 19316 6700
rect 19363 6616 19372 6656
rect 19412 6616 25612 6656
rect 25652 6616 25661 6656
rect 28339 6616 28348 6656
rect 28388 6616 34540 6656
rect 34580 6616 34589 6656
rect 14659 6532 14668 6572
rect 14708 6532 17740 6572
rect 17780 6532 17789 6572
rect 19276 6532 20044 6572
rect 20084 6532 20093 6572
rect 20179 6532 20188 6572
rect 20228 6532 23308 6572
rect 23348 6532 23357 6572
rect 46278 6488 46368 6508
rect 16771 6448 16780 6488
rect 16820 6448 19276 6488
rect 19316 6448 19325 6488
rect 19939 6448 19948 6488
rect 19988 6448 19997 6488
rect 20249 6448 20332 6488
rect 20372 6448 20380 6488
rect 20420 6448 20429 6488
rect 20899 6448 20908 6488
rect 20948 6448 22540 6488
rect 22580 6448 22589 6488
rect 28099 6448 28108 6488
rect 28148 6448 28157 6488
rect 33187 6448 33196 6488
rect 33236 6448 33367 6488
rect 43180 6448 44524 6488
rect 44564 6448 44573 6488
rect 44899 6448 44908 6488
rect 44948 6448 44957 6488
rect 45139 6448 45148 6488
rect 45188 6448 46368 6488
rect 19948 6404 19988 6448
rect 16963 6364 16972 6404
rect 17012 6364 19660 6404
rect 19700 6364 19709 6404
rect 19948 6364 20812 6404
rect 20852 6364 20861 6404
rect 20908 6364 24844 6404
rect 24884 6364 24893 6404
rect 20908 6320 20948 6364
rect 28108 6320 28148 6448
rect 43180 6404 43220 6448
rect 44908 6404 44948 6448
rect 46278 6428 46368 6448
rect 28579 6364 28588 6404
rect 28628 6364 43220 6404
rect 44611 6364 44620 6404
rect 44660 6364 44948 6404
rect 13996 6280 18412 6320
rect 18452 6280 18461 6320
rect 18595 6280 18604 6320
rect 18644 6280 20948 6320
rect 20995 6280 21004 6320
rect 21044 6280 25708 6320
rect 25748 6280 25757 6320
rect 28108 6280 34444 6320
rect 34484 6280 34493 6320
rect 11059 6196 11068 6236
rect 11108 6196 12980 6236
rect 13900 6196 17548 6236
rect 17588 6196 17597 6236
rect 17731 6196 17740 6236
rect 17780 6196 20236 6236
rect 20276 6196 20285 6236
rect 20659 6196 20668 6236
rect 20708 6196 24076 6236
rect 24116 6196 24125 6236
rect 33427 6196 33436 6236
rect 33476 6196 41740 6236
rect 41780 6196 41789 6236
rect 44755 6196 44764 6236
rect 44804 6196 44813 6236
rect 0 6152 90 6172
rect 0 6112 556 6152
rect 596 6112 605 6152
rect 0 6092 90 6112
rect 4919 6028 4928 6068
rect 4968 6028 5010 6068
rect 5050 6028 5092 6068
rect 5132 6028 5174 6068
rect 5214 6028 5256 6068
rect 5296 6028 5305 6068
rect 12940 5984 12980 6196
rect 44764 6152 44804 6196
rect 46278 6152 46368 6172
rect 17443 6112 17452 6152
rect 17492 6112 23596 6152
rect 23636 6112 23645 6152
rect 44764 6112 46368 6152
rect 46278 6092 46368 6112
rect 17155 6028 17164 6068
rect 17204 6028 19852 6068
rect 19892 6028 19901 6068
rect 20039 6028 20048 6068
rect 20088 6028 20130 6068
rect 20170 6028 20212 6068
rect 20252 6028 20294 6068
rect 20334 6028 20376 6068
rect 20416 6028 20425 6068
rect 20515 6028 20524 6068
rect 20564 6028 21964 6068
rect 22004 6028 22013 6068
rect 35159 6028 35168 6068
rect 35208 6028 35250 6068
rect 35290 6028 35332 6068
rect 35372 6028 35414 6068
rect 35454 6028 35496 6068
rect 35536 6028 35545 6068
rect 12940 5944 18700 5984
rect 18740 5944 18749 5984
rect 19939 5944 19948 5984
rect 19988 5944 25132 5984
rect 25172 5944 25181 5984
rect 11731 5860 11740 5900
rect 11780 5860 15916 5900
rect 15956 5860 15965 5900
rect 17539 5860 17548 5900
rect 17588 5860 20716 5900
rect 20756 5860 20765 5900
rect 0 5816 90 5836
rect 46278 5816 46368 5836
rect 0 5776 1036 5816
rect 1076 5776 1085 5816
rect 9676 5776 11924 5816
rect 12499 5776 12508 5816
rect 12548 5776 16204 5816
rect 16244 5776 16253 5816
rect 17347 5776 17356 5816
rect 17396 5776 21196 5816
rect 21236 5776 21245 5816
rect 21571 5776 21580 5816
rect 21620 5776 22732 5816
rect 22772 5776 22781 5816
rect 45139 5776 45148 5816
rect 45188 5776 46368 5816
rect 0 5756 90 5776
rect 9676 5732 9716 5776
rect 11884 5732 11924 5776
rect 46278 5756 46368 5776
rect 7564 5692 9716 5732
rect 9772 5692 11788 5732
rect 11828 5692 11837 5732
rect 11884 5692 12076 5732
rect 12116 5692 12125 5732
rect 12172 5692 12556 5732
rect 12596 5692 12605 5732
rect 12739 5692 12748 5732
rect 12788 5692 30068 5732
rect 7564 5648 7604 5692
rect 9772 5648 9812 5692
rect 12172 5648 12212 5692
rect 6569 5608 6700 5648
rect 6740 5608 6749 5648
rect 7555 5608 7564 5648
rect 7604 5608 7613 5648
rect 8707 5608 8716 5648
rect 8756 5608 8765 5648
rect 8947 5608 8956 5648
rect 8996 5608 9812 5648
rect 9859 5608 9868 5648
rect 9908 5608 10540 5648
rect 10580 5608 10589 5648
rect 10697 5608 10828 5648
rect 10868 5608 10877 5648
rect 11491 5608 11500 5648
rect 11540 5608 12212 5648
rect 12259 5608 12268 5648
rect 12308 5608 12652 5648
rect 12692 5608 12701 5648
rect 13123 5608 13132 5648
rect 13172 5608 13516 5648
rect 13556 5608 13565 5648
rect 15907 5608 15916 5648
rect 15956 5608 20332 5648
rect 20372 5608 20381 5648
rect 20515 5608 20524 5648
rect 20564 5608 21004 5648
rect 21044 5608 21053 5648
rect 21379 5608 21388 5648
rect 21428 5608 21437 5648
rect 21484 5608 21772 5648
rect 21812 5608 21821 5648
rect 22003 5608 22012 5648
rect 22052 5608 29932 5648
rect 29972 5608 29981 5648
rect 8716 5564 8756 5608
rect 21388 5564 21428 5608
rect 21484 5564 21524 5608
rect 6931 5524 6940 5564
rect 6980 5524 8620 5564
rect 8660 5524 8669 5564
rect 8716 5524 9964 5564
rect 10004 5524 10013 5564
rect 10099 5524 10108 5564
rect 10148 5524 11500 5564
rect 11540 5524 11549 5564
rect 20707 5524 20716 5564
rect 20756 5524 21428 5564
rect 21475 5524 21484 5564
rect 21524 5524 21533 5564
rect 21619 5524 21628 5564
rect 21668 5524 28972 5564
rect 29012 5524 29021 5564
rect 0 5480 90 5500
rect 0 5440 844 5480
rect 884 5440 893 5480
rect 7795 5440 7804 5480
rect 7844 5440 8716 5480
rect 8756 5440 8765 5480
rect 11059 5440 11068 5480
rect 11108 5440 12172 5480
rect 12212 5440 12221 5480
rect 13747 5440 13756 5480
rect 13796 5440 20908 5480
rect 20948 5440 20957 5480
rect 21235 5440 21244 5480
rect 21284 5440 22196 5480
rect 23107 5440 23116 5480
rect 23156 5440 28876 5480
rect 28916 5440 28925 5480
rect 0 5420 90 5440
rect 8131 5356 8140 5396
rect 8180 5356 10060 5396
rect 10100 5356 10109 5396
rect 19939 5356 19948 5396
rect 19988 5356 21292 5396
rect 21332 5356 21341 5396
rect 22156 5312 22196 5440
rect 30028 5396 30068 5692
rect 37612 5692 38516 5732
rect 38563 5692 38572 5732
rect 38612 5692 43084 5732
rect 43124 5692 43133 5732
rect 37612 5648 37652 5692
rect 38476 5648 38516 5692
rect 34147 5608 34156 5648
rect 34196 5608 34348 5648
rect 34388 5608 34397 5648
rect 36809 5608 36940 5648
rect 36980 5608 36989 5648
rect 37481 5608 37516 5648
rect 37556 5608 37612 5648
rect 37652 5608 37661 5648
rect 37769 5608 37900 5648
rect 37940 5608 38092 5648
rect 38132 5608 38141 5648
rect 38467 5608 38476 5648
rect 38516 5608 38525 5648
rect 38707 5608 38716 5648
rect 38756 5608 41012 5648
rect 43843 5608 43852 5648
rect 43892 5608 44524 5648
rect 44564 5608 44573 5648
rect 44620 5608 44908 5648
rect 44948 5608 44957 5648
rect 37036 5524 38228 5564
rect 38323 5524 38332 5564
rect 38372 5524 40820 5564
rect 37036 5480 37076 5524
rect 38188 5480 38228 5524
rect 34387 5440 34396 5480
rect 34436 5440 37076 5480
rect 37171 5440 37180 5480
rect 37220 5440 38092 5480
rect 38132 5440 38141 5480
rect 38188 5440 38804 5480
rect 22243 5356 22252 5396
rect 22292 5356 29356 5396
rect 29396 5356 29405 5396
rect 30028 5356 30260 5396
rect 3679 5272 3688 5312
rect 3728 5272 3770 5312
rect 3810 5272 3852 5312
rect 3892 5272 3934 5312
rect 3974 5272 4016 5312
rect 4056 5272 4065 5312
rect 8611 5272 8620 5312
rect 8660 5272 9676 5312
rect 9716 5272 9725 5312
rect 9955 5272 9964 5312
rect 10004 5272 11692 5312
rect 11732 5272 11741 5312
rect 12076 5272 12748 5312
rect 12788 5272 12797 5312
rect 18799 5272 18808 5312
rect 18848 5272 18890 5312
rect 18930 5272 18972 5312
rect 19012 5272 19054 5312
rect 19094 5272 19136 5312
rect 19176 5272 19185 5312
rect 22156 5272 29548 5312
rect 29588 5272 29597 5312
rect 12076 5228 12116 5272
rect 30220 5228 30260 5356
rect 33919 5272 33928 5312
rect 33968 5272 34010 5312
rect 34050 5272 34092 5312
rect 34132 5272 34174 5312
rect 34214 5272 34256 5312
rect 34296 5272 34305 5312
rect 38764 5228 38804 5440
rect 40780 5396 40820 5524
rect 40972 5480 41012 5608
rect 44620 5564 44660 5608
rect 41059 5524 41068 5564
rect 41108 5524 44660 5564
rect 44755 5524 44764 5564
rect 44804 5524 45620 5564
rect 45580 5480 45620 5524
rect 46278 5480 46368 5500
rect 40972 5440 44140 5480
rect 44180 5440 44189 5480
rect 45580 5440 46368 5480
rect 46278 5420 46368 5440
rect 40780 5356 44332 5396
rect 44372 5356 44381 5396
rect 4771 5188 4780 5228
rect 4820 5188 12116 5228
rect 12163 5188 12172 5228
rect 12212 5188 21388 5228
rect 21428 5188 21437 5228
rect 30220 5188 38708 5228
rect 38764 5188 44716 5228
rect 44756 5188 44765 5228
rect 0 5144 90 5164
rect 0 5104 1324 5144
rect 1364 5104 1373 5144
rect 1420 5104 33140 5144
rect 0 5084 90 5104
rect 1420 5060 1460 5104
rect 739 5020 748 5060
rect 788 5020 1460 5060
rect 1612 5020 23060 5060
rect 23107 5020 23116 5060
rect 23156 5020 26900 5060
rect 26947 5020 26956 5060
rect 26996 5020 28148 5060
rect 28339 5020 28348 5060
rect 28388 5020 31660 5060
rect 31700 5020 31709 5060
rect 1612 4976 1652 5020
rect 1411 4936 1420 4976
rect 1460 4936 1652 4976
rect 7049 4936 7180 4976
rect 7220 4936 7229 4976
rect 7411 4936 7420 4976
rect 7460 4936 7508 4976
rect 7555 4936 7564 4976
rect 7604 4936 7735 4976
rect 8323 4936 8332 4976
rect 8372 4936 11596 4976
rect 11636 4936 11645 4976
rect 11779 4936 11788 4976
rect 11828 4936 15916 4976
rect 15956 4936 15965 4976
rect 19843 4936 19852 4976
rect 19892 4936 22060 4976
rect 22100 4936 22109 4976
rect 22243 4936 22252 4976
rect 22292 4936 22300 4976
rect 22340 4936 22423 4976
rect 22474 4936 22483 4976
rect 22523 4936 22580 4976
rect 22793 4936 22924 4976
rect 22964 4936 22973 4976
rect 7468 4892 7508 4936
rect 22540 4892 22580 4936
rect 7468 4852 11308 4892
rect 11348 4852 11357 4892
rect 11491 4852 11500 4892
rect 11540 4852 18700 4892
rect 18740 4852 18749 4892
rect 19651 4852 19660 4892
rect 19700 4852 22580 4892
rect 23020 4892 23060 5020
rect 26860 4976 26900 5020
rect 28108 4976 28148 5020
rect 33100 4976 33140 5104
rect 34540 5020 38572 5060
rect 38612 5020 38621 5060
rect 23273 4936 23404 4976
rect 23444 4936 23453 4976
rect 26851 4936 26860 4976
rect 26900 4936 26909 4976
rect 27715 4936 27724 4976
rect 27764 4936 27773 4976
rect 28099 4936 28108 4976
rect 28148 4936 28157 4976
rect 28483 4936 28492 4976
rect 28532 4936 28541 4976
rect 33100 4936 34156 4976
rect 34196 4936 34348 4976
rect 34388 4936 34444 4976
rect 34484 4936 34493 4976
rect 27724 4892 27764 4936
rect 28492 4892 28532 4936
rect 34540 4892 34580 5020
rect 38668 4976 38708 5188
rect 46278 5144 46368 5164
rect 38899 5104 38908 5144
rect 38948 5104 41068 5144
rect 41108 5104 41117 5144
rect 41347 5104 41356 5144
rect 41396 5104 44564 5144
rect 45139 5104 45148 5144
rect 45188 5104 46368 5144
rect 39148 5020 40876 5060
rect 40916 5020 40925 5060
rect 41011 5020 41020 5060
rect 41060 5020 44236 5060
rect 44276 5020 44285 5060
rect 38659 4936 38668 4976
rect 38708 4936 38717 4976
rect 23020 4852 27764 4892
rect 27811 4852 27820 4892
rect 27860 4852 28532 4892
rect 32428 4852 34580 4892
rect 38083 4852 38092 4892
rect 38132 4852 39052 4892
rect 39092 4852 39101 4892
rect 0 4808 90 4828
rect 32428 4808 32468 4852
rect 39148 4808 39188 5020
rect 44524 4976 44564 5104
rect 46278 5084 46368 5104
rect 0 4768 27860 4808
rect 27955 4768 27964 4808
rect 28004 4768 32468 4808
rect 33100 4768 39188 4808
rect 39436 4936 39628 4976
rect 39668 4936 39677 4976
rect 40483 4936 40492 4976
rect 40532 4936 40780 4976
rect 40820 4936 40829 4976
rect 41155 4936 41164 4976
rect 41204 4936 41213 4976
rect 44515 4936 44524 4976
rect 44564 4936 44573 4976
rect 44899 4936 44908 4976
rect 44948 4936 44957 4976
rect 0 4748 90 4768
rect 7795 4684 7804 4724
rect 7844 4684 8332 4724
rect 8372 4684 8381 4724
rect 8563 4684 8572 4724
rect 8612 4684 15148 4724
rect 15188 4684 15197 4724
rect 16195 4684 16204 4724
rect 16244 4684 21676 4724
rect 21716 4684 21725 4724
rect 22675 4684 22684 4724
rect 22724 4684 23020 4724
rect 23060 4684 23069 4724
rect 23155 4684 23164 4724
rect 23204 4684 23444 4724
rect 23635 4684 23644 4724
rect 23684 4684 26956 4724
rect 26996 4684 27005 4724
rect 27091 4684 27100 4724
rect 27140 4684 27764 4724
rect 10051 4600 10060 4640
rect 10100 4600 10636 4640
rect 10676 4600 10685 4640
rect 10819 4600 10828 4640
rect 10868 4600 12556 4640
rect 12596 4600 12605 4640
rect 19459 4600 19468 4640
rect 19508 4600 22924 4640
rect 22964 4600 22973 4640
rect 23404 4556 23444 4684
rect 27724 4556 27764 4684
rect 27820 4640 27860 4768
rect 28723 4684 28732 4724
rect 28772 4684 31276 4724
rect 31316 4684 31325 4724
rect 27820 4600 30796 4640
rect 30836 4600 30845 4640
rect 33100 4556 33140 4768
rect 37603 4684 37612 4724
rect 37652 4684 37699 4724
rect 37739 4684 37783 4724
rect 38362 4684 38371 4724
rect 38411 4684 38420 4724
rect 39034 4684 39043 4724
rect 39083 4684 39092 4724
rect 39209 4684 39331 4724
rect 39380 4684 39389 4724
rect 38380 4640 38420 4684
rect 39052 4640 39092 4684
rect 39436 4640 39476 4936
rect 41164 4892 41204 4936
rect 44908 4892 44948 4936
rect 40099 4852 40108 4892
rect 40148 4852 41548 4892
rect 41588 4852 41836 4892
rect 41876 4852 41885 4892
rect 44035 4852 44044 4892
rect 44084 4852 44948 4892
rect 46278 4808 46368 4828
rect 39859 4768 39868 4808
rect 39908 4768 41260 4808
rect 41300 4768 41309 4808
rect 41395 4768 41404 4808
rect 41444 4768 44428 4808
rect 44468 4768 44477 4808
rect 44755 4768 44764 4808
rect 44804 4768 46368 4808
rect 46278 4748 46368 4768
rect 39977 4684 40099 4724
rect 40148 4684 40157 4724
rect 40291 4684 40300 4724
rect 40340 4684 40483 4724
rect 40523 4684 40532 4724
rect 41818 4684 41827 4724
rect 41867 4684 41876 4724
rect 37411 4600 37420 4640
rect 37460 4600 39476 4640
rect 4919 4516 4928 4556
rect 4968 4516 5010 4556
rect 5050 4516 5092 4556
rect 5132 4516 5174 4556
rect 5214 4516 5256 4556
rect 5296 4516 5305 4556
rect 8419 4516 8428 4556
rect 8468 4516 18220 4556
rect 18260 4516 18269 4556
rect 18691 4516 18700 4556
rect 18740 4516 19756 4556
rect 19796 4516 19805 4556
rect 20039 4516 20048 4556
rect 20088 4516 20130 4556
rect 20170 4516 20212 4556
rect 20252 4516 20294 4556
rect 20334 4516 20376 4556
rect 20416 4516 20425 4556
rect 21571 4516 21580 4556
rect 21620 4516 22636 4556
rect 22676 4516 22685 4556
rect 23404 4516 27476 4556
rect 27724 4516 30220 4556
rect 30260 4516 30269 4556
rect 30316 4516 33140 4556
rect 35159 4516 35168 4556
rect 35208 4516 35250 4556
rect 35290 4516 35332 4556
rect 35372 4516 35414 4556
rect 35454 4516 35496 4556
rect 35536 4516 35545 4556
rect 35971 4516 35980 4556
rect 36020 4516 41356 4556
rect 41396 4516 41405 4556
rect 0 4472 90 4492
rect 27436 4472 27476 4516
rect 30316 4472 30356 4516
rect 0 4432 1420 4472
rect 1460 4432 1469 4472
rect 7555 4432 7564 4472
rect 7604 4432 11404 4472
rect 11444 4432 11453 4472
rect 19555 4432 19564 4472
rect 19604 4432 23404 4472
rect 23444 4432 23453 4472
rect 27436 4432 28012 4472
rect 28052 4432 28061 4472
rect 28195 4432 28204 4472
rect 28244 4432 30356 4472
rect 41836 4472 41876 4684
rect 46278 4472 46368 4492
rect 41836 4432 42260 4472
rect 0 4412 90 4432
rect 42220 4388 42260 4432
rect 45148 4432 46368 4472
rect 7171 4348 7180 4388
rect 7220 4348 11212 4388
rect 11252 4348 11261 4388
rect 18307 4348 18316 4388
rect 18356 4348 22828 4388
rect 22868 4348 22877 4388
rect 26947 4348 26956 4388
rect 26996 4348 30700 4388
rect 30740 4348 30749 4388
rect 30883 4348 30892 4388
rect 30932 4348 34828 4388
rect 34868 4348 34877 4388
rect 39209 4348 39331 4388
rect 39380 4348 40003 4388
rect 40043 4348 40300 4388
rect 40340 4348 40483 4388
rect 40523 4348 40771 4388
rect 40811 4348 41059 4388
rect 41099 4348 41347 4388
rect 41387 4348 41635 4388
rect 41675 4348 41876 4388
rect 42202 4348 42211 4388
rect 42251 4348 42787 4388
rect 42827 4348 42836 4388
rect 41836 4304 41876 4348
rect 45148 4304 45188 4432
rect 46278 4412 46368 4432
rect 1036 4264 37996 4304
rect 38036 4264 38045 4304
rect 41836 4264 41932 4304
rect 41972 4264 42508 4304
rect 42548 4264 42557 4304
rect 45139 4264 45148 4304
rect 45188 4264 45197 4304
rect 0 4136 90 4156
rect 1036 4136 1076 4264
rect 1123 4180 1132 4220
rect 1172 4180 23116 4220
rect 23156 4180 23165 4220
rect 24556 4180 27052 4220
rect 27092 4180 27101 4220
rect 27532 4180 28492 4220
rect 28532 4180 28541 4220
rect 30508 4180 35596 4220
rect 35636 4180 35645 4220
rect 37180 4180 38092 4220
rect 38132 4180 38141 4220
rect 41251 4180 41260 4220
rect 41300 4180 43220 4220
rect 0 4096 1076 4136
rect 7075 4096 7084 4136
rect 7124 4096 11020 4136
rect 11060 4096 11069 4136
rect 19363 4096 19372 4136
rect 19412 4096 23980 4136
rect 24020 4096 24029 4136
rect 24329 4096 24460 4136
rect 24500 4096 24509 4136
rect 0 4076 90 4096
rect 24556 4052 24596 4180
rect 27532 4136 27572 4180
rect 30508 4136 30548 4180
rect 37180 4136 37220 4180
rect 25193 4096 25324 4136
rect 25364 4096 25373 4136
rect 25555 4096 25564 4136
rect 25604 4096 25996 4136
rect 26036 4096 26045 4136
rect 26179 4096 26188 4136
rect 26228 4096 26237 4136
rect 26419 4096 26428 4136
rect 26468 4096 27572 4136
rect 27619 4096 27628 4136
rect 27668 4096 27677 4136
rect 27859 4096 27868 4136
rect 27908 4096 30548 4136
rect 32611 4096 32620 4136
rect 32660 4096 32669 4136
rect 32851 4096 32860 4136
rect 32900 4096 37220 4136
rect 43180 4136 43220 4180
rect 46278 4136 46368 4156
rect 43180 4096 44140 4136
rect 44180 4096 44189 4136
rect 44393 4096 44524 4136
rect 44564 4096 44573 4136
rect 44777 4096 44908 4136
rect 44948 4096 44957 4136
rect 45580 4096 46368 4136
rect 835 4012 844 4052
rect 884 4012 24596 4052
rect 24691 4012 24700 4052
rect 24740 4012 24940 4052
rect 24980 4012 24989 4052
rect 25516 4012 25900 4052
rect 25940 4012 25949 4052
rect 25516 3968 25556 4012
rect 26188 3968 26228 4096
rect 27628 4052 27668 4096
rect 26380 4012 27436 4052
rect 27476 4012 27485 4052
rect 27628 4012 30892 4052
rect 30932 4012 30941 4052
rect 931 3928 940 3968
rect 980 3928 5932 3968
rect 5972 3928 5981 3968
rect 7315 3928 7324 3968
rect 7364 3928 10156 3968
rect 10196 3928 10205 3968
rect 10339 3928 10348 3968
rect 10388 3928 19276 3968
rect 19316 3928 19325 3968
rect 24211 3928 24220 3968
rect 24260 3928 25556 3968
rect 26179 3928 26188 3968
rect 26228 3928 26237 3968
rect 26380 3884 26420 4012
rect 32620 3968 32660 4096
rect 45580 4052 45620 4096
rect 46278 4076 46368 4096
rect 37315 4012 37324 4052
rect 37364 4012 43852 4052
rect 43892 4012 43901 4052
rect 44755 4012 44764 4052
rect 44804 4012 45620 4052
rect 1027 3844 1036 3884
rect 1076 3844 10060 3884
rect 10100 3844 10109 3884
rect 10435 3844 10444 3884
rect 10484 3844 26420 3884
rect 27436 3928 32660 3968
rect 44371 3928 44380 3968
rect 44420 3928 45044 3968
rect 0 3800 90 3820
rect 27436 3800 27476 3928
rect 27523 3844 27532 3884
rect 27572 3844 37132 3884
rect 37172 3844 37181 3884
rect 38083 3844 38092 3884
rect 38132 3844 44948 3884
rect 0 3760 2900 3800
rect 3679 3760 3688 3800
rect 3728 3760 3770 3800
rect 3810 3760 3852 3800
rect 3892 3760 3934 3800
rect 3974 3760 4016 3800
rect 4056 3760 4065 3800
rect 4108 3760 10252 3800
rect 10292 3760 10301 3800
rect 18799 3760 18808 3800
rect 18848 3760 18890 3800
rect 18930 3760 18972 3800
rect 19012 3760 19054 3800
rect 19094 3760 19136 3800
rect 19176 3760 19185 3800
rect 19267 3760 19276 3800
rect 19316 3760 27476 3800
rect 27619 3760 27628 3800
rect 27668 3760 33140 3800
rect 33919 3760 33928 3800
rect 33968 3760 34010 3800
rect 34050 3760 34092 3800
rect 34132 3760 34174 3800
rect 34214 3760 34256 3800
rect 34296 3760 34305 3800
rect 0 3740 90 3760
rect 2860 3716 2900 3760
rect 4108 3716 4148 3760
rect 33100 3716 33140 3760
rect 2860 3676 4148 3716
rect 5923 3676 5932 3716
rect 5972 3676 28724 3716
rect 33100 3676 37420 3716
rect 37460 3676 37469 3716
rect 1315 3592 1324 3632
rect 1364 3592 26420 3632
rect 26755 3592 26764 3632
rect 26804 3592 26908 3632
rect 26948 3592 26957 3632
rect 27283 3592 27292 3632
rect 27332 3592 27532 3632
rect 27572 3592 27581 3632
rect 27667 3592 27676 3632
rect 27716 3592 28204 3632
rect 28244 3592 28253 3632
rect 1411 3508 1420 3548
rect 1460 3508 20140 3548
rect 20180 3508 20189 3548
rect 23107 3508 23116 3548
rect 23156 3508 26324 3548
rect 0 3464 90 3484
rect 26284 3464 26324 3508
rect 0 3424 24748 3464
rect 24788 3424 24797 3464
rect 25891 3424 25900 3464
rect 25940 3424 25996 3464
rect 26036 3424 26071 3464
rect 26275 3424 26284 3464
rect 26324 3424 26333 3464
rect 0 3404 90 3424
rect 26380 3380 26420 3592
rect 28684 3464 28724 3676
rect 30931 3592 30940 3632
rect 30980 3592 37844 3632
rect 38131 3592 38140 3632
rect 38180 3592 44524 3632
rect 44564 3592 44573 3632
rect 30115 3508 30124 3548
rect 30164 3508 36596 3548
rect 36556 3464 36596 3508
rect 26659 3424 26668 3464
rect 26708 3424 26764 3464
rect 26804 3424 26839 3464
rect 27043 3424 27052 3464
rect 27092 3424 27223 3464
rect 27427 3424 27436 3464
rect 27476 3424 27607 3464
rect 27811 3424 27820 3464
rect 27860 3424 27991 3464
rect 28073 3424 28204 3464
rect 28244 3424 28253 3464
rect 28435 3424 28444 3464
rect 28484 3424 28588 3464
rect 28628 3424 28637 3464
rect 28684 3424 30028 3464
rect 30068 3424 30077 3464
rect 30691 3424 30700 3464
rect 30740 3424 30749 3464
rect 30883 3424 30892 3464
rect 30932 3424 34444 3464
rect 34484 3424 34493 3464
rect 34697 3424 34828 3464
rect 34868 3424 34877 3464
rect 35059 3424 35068 3464
rect 35108 3424 35980 3464
rect 36020 3424 36029 3464
rect 36547 3424 36556 3464
rect 36596 3424 36605 3464
rect 30700 3380 30740 3424
rect 10147 3340 10156 3380
rect 10196 3340 18700 3380
rect 18740 3340 18749 3380
rect 26380 3340 30740 3380
rect 37804 3380 37844 3592
rect 44908 3464 44948 3844
rect 45004 3464 45044 3928
rect 46278 3800 46368 3820
rect 45148 3760 46368 3800
rect 45148 3632 45188 3760
rect 46278 3740 46368 3760
rect 45139 3592 45148 3632
rect 45188 3592 45197 3632
rect 46278 3464 46368 3484
rect 37891 3424 37900 3464
rect 37940 3424 37996 3464
rect 38036 3424 38071 3464
rect 41059 3424 41068 3464
rect 41108 3424 44524 3464
rect 44564 3424 44573 3464
rect 44899 3424 44908 3464
rect 44948 3424 44957 3464
rect 45004 3424 46368 3464
rect 46278 3404 46368 3424
rect 37804 3340 44044 3380
rect 44084 3340 44093 3380
rect 19555 3256 19564 3296
rect 19604 3256 24460 3296
rect 24500 3256 24509 3296
rect 27907 3256 27916 3296
rect 27956 3256 29588 3296
rect 30259 3256 30268 3296
rect 30308 3256 35252 3296
rect 36787 3256 36796 3296
rect 36836 3256 44908 3296
rect 44948 3256 44957 3296
rect 29548 3212 29588 3256
rect 18979 3172 18988 3212
rect 19028 3172 25324 3212
rect 25364 3172 25373 3212
rect 26131 3172 26140 3212
rect 26180 3172 26380 3212
rect 26420 3172 26429 3212
rect 26515 3172 26524 3212
rect 26564 3172 26804 3212
rect 28051 3172 28060 3212
rect 28100 3172 28396 3212
rect 28436 3172 28445 3212
rect 29548 3172 34732 3212
rect 34772 3172 34781 3212
rect 0 3128 90 3148
rect 26764 3128 26804 3172
rect 35212 3128 35252 3256
rect 44755 3172 44764 3212
rect 44804 3172 44813 3212
rect 44764 3128 44804 3172
rect 46278 3128 46368 3148
rect 0 3088 4780 3128
rect 4820 3088 4829 3128
rect 18499 3088 18508 3128
rect 18548 3088 26188 3128
rect 26228 3088 26237 3128
rect 26764 3088 27340 3128
rect 27380 3088 27389 3128
rect 27811 3088 27820 3128
rect 27860 3088 35020 3128
rect 35060 3088 35069 3128
rect 35212 3088 44620 3128
rect 44660 3088 44669 3128
rect 44764 3088 46368 3128
rect 0 3068 90 3088
rect 46278 3068 46368 3088
rect 4919 3004 4928 3044
rect 4968 3004 5010 3044
rect 5050 3004 5092 3044
rect 5132 3004 5174 3044
rect 5214 3004 5256 3044
rect 5296 3004 5305 3044
rect 20039 3004 20048 3044
rect 20088 3004 20130 3044
rect 20170 3004 20212 3044
rect 20252 3004 20294 3044
rect 20334 3004 20376 3044
rect 20416 3004 20425 3044
rect 24931 3004 24940 3044
rect 24980 3004 26092 3044
rect 26132 3004 26141 3044
rect 26755 3004 26764 3044
rect 26804 3004 34636 3044
rect 34676 3004 34685 3044
rect 35159 3004 35168 3044
rect 35208 3004 35250 3044
rect 35290 3004 35332 3044
rect 35372 3004 35414 3044
rect 35454 3004 35496 3044
rect 35536 3004 35545 3044
rect 547 2920 556 2960
rect 596 2920 28204 2960
rect 28244 2920 28253 2960
rect 9667 2836 9676 2876
rect 9716 2836 22828 2876
rect 22868 2836 22877 2876
rect 23011 2836 23020 2876
rect 23060 2836 23828 2876
rect 25123 2836 25132 2876
rect 25172 2836 25181 2876
rect 25507 2836 25516 2876
rect 25556 2836 27572 2876
rect 34697 2836 34828 2876
rect 34868 2836 35107 2876
rect 35147 2836 35156 2876
rect 0 2792 90 2812
rect 0 2752 1420 2792
rect 1460 2752 1469 2792
rect 8707 2752 8716 2792
rect 8756 2752 23444 2792
rect 0 2732 90 2752
rect 11299 2668 11308 2708
rect 11348 2668 21908 2708
rect 21955 2668 21964 2708
rect 22004 2668 23348 2708
rect 21868 2624 21908 2668
rect 15139 2584 15148 2624
rect 15188 2584 21484 2624
rect 21524 2584 21533 2624
rect 21859 2584 21868 2624
rect 21908 2584 21917 2624
rect 22243 2584 22252 2624
rect 22292 2584 22301 2624
rect 22505 2584 22636 2624
rect 22676 2584 22685 2624
rect 22924 2584 23020 2624
rect 23060 2584 23124 2624
rect 22252 2540 22292 2584
rect 19171 2500 19180 2540
rect 19220 2500 20044 2540
rect 20084 2500 20093 2540
rect 20899 2500 20908 2540
rect 20948 2500 22292 2540
rect 0 2456 90 2476
rect 0 2416 1420 2456
rect 1460 2416 1469 2456
rect 19075 2416 19084 2456
rect 19124 2416 19316 2456
rect 21113 2416 21196 2456
rect 21236 2416 21244 2456
rect 21284 2416 21293 2456
rect 21497 2416 21580 2456
rect 21620 2416 21628 2456
rect 21668 2416 21677 2456
rect 21881 2416 21964 2456
rect 22004 2416 22012 2456
rect 22052 2416 22061 2456
rect 22265 2416 22348 2456
rect 22388 2416 22396 2456
rect 22436 2416 22445 2456
rect 22649 2416 22732 2456
rect 22772 2416 22780 2456
rect 22820 2416 22829 2456
rect 0 2396 90 2416
rect 19276 2288 19316 2416
rect 22924 2372 22964 2584
rect 23308 2540 23348 2668
rect 23404 2624 23444 2752
rect 23788 2624 23828 2836
rect 25132 2792 25172 2836
rect 25132 2752 25420 2792
rect 25460 2752 25469 2792
rect 25699 2752 25708 2792
rect 25748 2752 26708 2792
rect 24451 2668 24460 2708
rect 24500 2668 25652 2708
rect 25795 2668 25804 2708
rect 25844 2668 26324 2708
rect 25612 2624 25652 2668
rect 26284 2624 26324 2668
rect 26668 2624 26708 2752
rect 27139 2668 27148 2708
rect 27188 2668 27197 2708
rect 27148 2624 27188 2668
rect 27532 2624 27572 2836
rect 46278 2792 46368 2812
rect 27907 2752 27916 2792
rect 27956 2752 30164 2792
rect 45139 2752 45148 2792
rect 45188 2752 46368 2792
rect 28003 2668 28012 2708
rect 28052 2668 29780 2708
rect 29740 2624 29780 2668
rect 30124 2624 30164 2752
rect 46278 2732 46368 2752
rect 30211 2668 30220 2708
rect 30260 2668 30932 2708
rect 44227 2668 44236 2708
rect 44276 2668 44948 2708
rect 30892 2624 30932 2668
rect 44908 2624 44948 2668
rect 23395 2584 23404 2624
rect 23444 2584 23453 2624
rect 23779 2584 23788 2624
rect 23828 2584 23837 2624
rect 23971 2584 23980 2624
rect 24020 2584 25516 2624
rect 25556 2584 25565 2624
rect 25612 2584 25900 2624
rect 25940 2584 25949 2624
rect 26275 2584 26284 2624
rect 26324 2584 26333 2624
rect 26659 2584 26668 2624
rect 26708 2584 26717 2624
rect 27043 2584 27052 2624
rect 27092 2584 27101 2624
rect 27148 2584 27436 2624
rect 27476 2584 27485 2624
rect 27532 2584 27820 2624
rect 27860 2584 27869 2624
rect 28195 2584 28204 2624
rect 28244 2584 28253 2624
rect 28387 2584 28396 2624
rect 28436 2584 28588 2624
rect 28628 2584 28637 2624
rect 28841 2584 28972 2624
rect 29012 2584 29021 2624
rect 29225 2584 29356 2624
rect 29396 2584 29405 2624
rect 29731 2584 29740 2624
rect 29780 2584 29789 2624
rect 30115 2584 30124 2624
rect 30164 2584 30173 2624
rect 30499 2584 30508 2624
rect 30548 2584 30557 2624
rect 30883 2584 30892 2624
rect 30932 2584 30941 2624
rect 31145 2584 31276 2624
rect 31316 2584 31325 2624
rect 44009 2584 44140 2624
rect 44180 2584 44189 2624
rect 44393 2584 44524 2624
rect 44564 2584 44573 2624
rect 44899 2584 44908 2624
rect 44948 2584 44957 2624
rect 27052 2540 27092 2584
rect 28204 2540 28244 2584
rect 30508 2540 30548 2584
rect 23308 2500 24940 2540
rect 24980 2500 24989 2540
rect 25315 2500 25324 2540
rect 25364 2500 27092 2540
rect 27292 2500 28244 2540
rect 29155 2500 29164 2540
rect 29204 2500 30548 2540
rect 44755 2500 44764 2540
rect 44804 2500 45812 2540
rect 23107 2416 23116 2456
rect 23156 2416 23164 2456
rect 23204 2416 23287 2456
rect 23417 2416 23500 2456
rect 23540 2416 23548 2456
rect 23588 2416 23597 2456
rect 25145 2416 25228 2456
rect 25268 2416 25276 2456
rect 25316 2416 25325 2456
rect 25529 2416 25612 2456
rect 25652 2416 25660 2456
rect 25700 2416 25709 2456
rect 25913 2416 25996 2456
rect 26036 2416 26044 2456
rect 26084 2416 26093 2456
rect 26297 2416 26380 2456
rect 26420 2416 26428 2456
rect 26468 2416 26477 2456
rect 26681 2416 26764 2456
rect 26804 2416 26812 2456
rect 26852 2416 26861 2456
rect 27065 2416 27148 2456
rect 27188 2416 27196 2456
rect 27236 2416 27245 2456
rect 27292 2372 27332 2500
rect 45772 2456 45812 2500
rect 46278 2456 46368 2476
rect 27449 2416 27532 2456
rect 27572 2416 27580 2456
rect 27620 2416 27629 2456
rect 27833 2416 27916 2456
rect 27956 2416 27964 2456
rect 28004 2416 28013 2456
rect 28217 2416 28300 2456
rect 28340 2416 28348 2456
rect 28388 2416 28397 2456
rect 28601 2416 28684 2456
rect 28724 2416 28732 2456
rect 28772 2416 28781 2456
rect 28985 2416 29068 2456
rect 29108 2416 29116 2456
rect 29156 2416 29165 2456
rect 29369 2416 29452 2456
rect 29492 2416 29500 2456
rect 29540 2416 29549 2456
rect 29753 2416 29836 2456
rect 29876 2416 29884 2456
rect 29924 2416 29933 2456
rect 30137 2416 30220 2456
rect 30260 2416 30268 2456
rect 30308 2416 30317 2456
rect 30521 2416 30604 2456
rect 30644 2416 30652 2456
rect 30692 2416 30701 2456
rect 30905 2416 30988 2456
rect 31028 2416 31036 2456
rect 31076 2416 31085 2456
rect 44371 2416 44380 2456
rect 44420 2416 45676 2456
rect 45716 2416 45725 2456
rect 45772 2416 46368 2456
rect 46278 2396 46368 2416
rect 19747 2332 19756 2372
rect 19796 2332 22964 2372
rect 23299 2332 23308 2372
rect 23348 2332 24788 2372
rect 25123 2332 25132 2372
rect 25172 2332 27332 2372
rect 24748 2288 24788 2332
rect 3679 2248 3688 2288
rect 3728 2248 3770 2288
rect 3810 2248 3852 2288
rect 3892 2248 3934 2288
rect 3974 2248 4016 2288
rect 4056 2248 4065 2288
rect 18799 2248 18808 2288
rect 18848 2248 18890 2288
rect 18930 2248 18972 2288
rect 19012 2248 19054 2288
rect 19094 2248 19136 2288
rect 19176 2248 19185 2288
rect 19276 2248 24556 2288
rect 24596 2248 24605 2288
rect 24748 2248 25460 2288
rect 33919 2248 33928 2288
rect 33968 2248 34010 2288
rect 34050 2248 34092 2288
rect 34132 2248 34174 2288
rect 34214 2248 34256 2288
rect 34296 2248 34305 2288
rect 16195 2164 16204 2204
rect 16244 2164 24116 2204
rect 0 2120 90 2140
rect 0 2080 748 2120
rect 788 2080 797 2120
rect 15907 2080 15916 2120
rect 15956 2080 22484 2120
rect 0 2060 90 2080
rect 18595 1996 18604 2036
rect 18644 1996 21332 2036
rect 21379 1996 21388 2036
rect 21428 1996 22100 2036
rect 21292 1952 21332 1996
rect 22060 1952 22100 1996
rect 22444 1952 22484 2080
rect 22531 1996 22540 2036
rect 22580 1996 23060 2036
rect 23020 1952 23060 1996
rect 24076 1952 24116 2164
rect 25420 2120 25460 2248
rect 25699 2164 25708 2204
rect 25748 2164 27052 2204
rect 27092 2164 27101 2204
rect 27331 2164 27340 2204
rect 27380 2164 31124 2204
rect 25420 2080 26132 2120
rect 26659 2080 26668 2120
rect 26708 2080 28052 2120
rect 28867 2080 28876 2120
rect 28916 2080 30356 2120
rect 24643 1996 24652 2036
rect 24692 1996 25364 2036
rect 25411 1996 25420 2036
rect 25460 1996 25844 2036
rect 25324 1952 25364 1996
rect 18211 1912 18220 1952
rect 18260 1912 20908 1952
rect 20948 1912 20957 1952
rect 21283 1912 21292 1952
rect 21332 1912 21341 1952
rect 21545 1912 21676 1952
rect 21716 1912 21725 1952
rect 22051 1912 22060 1952
rect 22100 1912 22109 1952
rect 22435 1912 22444 1952
rect 22484 1912 22493 1952
rect 22697 1912 22828 1952
rect 22868 1912 22877 1952
rect 23020 1912 23212 1952
rect 23252 1912 23261 1952
rect 23465 1912 23596 1952
rect 23636 1912 23645 1952
rect 23779 1912 23788 1952
rect 23828 1912 23980 1952
rect 24020 1912 24029 1952
rect 24076 1912 24556 1952
rect 24596 1912 24605 1952
rect 24809 1912 24940 1952
rect 24980 1912 24989 1952
rect 25315 1912 25324 1952
rect 25364 1912 25373 1952
rect 25699 1912 25708 1952
rect 25748 1912 25757 1952
rect 25708 1868 25748 1912
rect 24076 1828 25748 1868
rect 25804 1868 25844 1996
rect 26092 1952 26132 2080
rect 26179 1996 26188 2036
rect 26228 1996 27004 2036
rect 27044 1996 27053 2036
rect 28012 1952 28052 2080
rect 28099 1996 28108 2036
rect 28148 1996 29204 2036
rect 29251 1996 29260 2036
rect 29300 1996 30076 2036
rect 30116 1996 30125 2036
rect 29164 1952 29204 1996
rect 30316 1952 30356 2080
rect 31084 1952 31124 2164
rect 46278 2120 46368 2140
rect 45139 2080 45148 2120
rect 45188 2080 46368 2120
rect 46278 2060 46368 2080
rect 41731 1996 41740 2036
rect 41780 1996 44180 2036
rect 44140 1952 44180 1996
rect 26083 1912 26092 1952
rect 26132 1912 26141 1952
rect 26345 1912 26476 1952
rect 26516 1912 26525 1952
rect 26572 1912 26860 1952
rect 26900 1912 26909 1952
rect 27043 1912 27052 1952
rect 27092 1912 27244 1952
rect 27284 1912 27293 1952
rect 27427 1912 27436 1952
rect 27476 1912 27628 1952
rect 27668 1912 27677 1952
rect 28003 1912 28012 1952
rect 28052 1912 28061 1952
rect 28387 1912 28396 1952
rect 28436 1912 28445 1952
rect 28649 1912 28780 1952
rect 28820 1912 28829 1952
rect 29155 1912 29164 1952
rect 29204 1912 29213 1952
rect 29417 1912 29548 1952
rect 29588 1912 29597 1952
rect 29801 1912 29932 1952
rect 29972 1912 29981 1952
rect 30307 1912 30316 1952
rect 30356 1912 30365 1952
rect 30569 1912 30700 1952
rect 30740 1912 30749 1952
rect 31075 1912 31084 1952
rect 31124 1912 31133 1952
rect 31459 1912 31468 1952
rect 31508 1912 31517 1952
rect 31651 1912 31660 1952
rect 31700 1912 31852 1952
rect 31892 1912 31901 1952
rect 39043 1912 39052 1952
rect 39092 1912 43756 1952
rect 43796 1912 43805 1952
rect 44131 1912 44140 1952
rect 44180 1912 44189 1952
rect 44419 1912 44428 1952
rect 44468 1912 44524 1952
rect 44564 1912 44599 1952
rect 44707 1912 44716 1952
rect 44756 1912 44908 1952
rect 44948 1912 44957 1952
rect 26572 1868 26612 1912
rect 28396 1868 28436 1912
rect 31468 1868 31508 1912
rect 25804 1828 26612 1868
rect 26851 1828 26860 1868
rect 26900 1828 28436 1868
rect 28483 1828 28492 1868
rect 28532 1828 31508 1868
rect 0 1784 90 1804
rect 0 1744 1420 1784
rect 1460 1744 1469 1784
rect 0 1724 90 1744
rect 20035 1660 20044 1700
rect 20084 1660 20093 1700
rect 21139 1660 21148 1700
rect 21188 1660 21388 1700
rect 21428 1660 21437 1700
rect 21523 1660 21532 1700
rect 21572 1660 21772 1700
rect 21812 1660 21821 1700
rect 21907 1660 21916 1700
rect 21956 1660 22156 1700
rect 22196 1660 22205 1700
rect 22291 1660 22300 1700
rect 22340 1660 22540 1700
rect 22580 1660 22589 1700
rect 22675 1660 22684 1700
rect 22724 1660 22924 1700
rect 22964 1660 22973 1700
rect 23059 1660 23068 1700
rect 23108 1660 23308 1700
rect 23348 1660 23357 1700
rect 23443 1660 23452 1700
rect 23492 1660 23692 1700
rect 23732 1660 23741 1700
rect 23827 1660 23836 1700
rect 23876 1660 23884 1700
rect 23924 1660 24007 1700
rect 20044 1616 20084 1660
rect 24076 1616 24116 1828
rect 46278 1784 46368 1804
rect 24163 1744 24172 1784
rect 24212 1744 24220 1784
rect 24260 1744 24343 1784
rect 24643 1744 24652 1784
rect 24692 1744 25084 1784
rect 25124 1744 25133 1784
rect 25411 1744 25420 1784
rect 25460 1744 26236 1784
rect 26276 1744 26285 1784
rect 26947 1744 26956 1784
rect 26996 1744 27772 1784
rect 27812 1744 27821 1784
rect 28099 1744 28108 1784
rect 28148 1744 28924 1784
rect 28964 1744 28973 1784
rect 30019 1744 30028 1784
rect 30068 1744 30844 1784
rect 30884 1744 30893 1784
rect 43987 1744 43996 1784
rect 44036 1744 44620 1784
rect 44660 1744 44669 1784
rect 44755 1744 44764 1784
rect 44804 1744 46368 1784
rect 46278 1724 46368 1744
rect 24185 1660 24268 1700
rect 24308 1660 24316 1700
rect 24356 1660 24365 1700
rect 24451 1660 24460 1700
rect 24500 1660 24700 1700
rect 24740 1660 24749 1700
rect 24835 1660 24844 1700
rect 24884 1660 25468 1700
rect 25508 1660 25517 1700
rect 25612 1660 25852 1700
rect 25892 1660 25901 1700
rect 26188 1660 26620 1700
rect 26660 1660 26669 1700
rect 26764 1660 27388 1700
rect 27428 1660 27437 1700
rect 27532 1660 28156 1700
rect 28196 1660 28205 1700
rect 28300 1660 28540 1700
rect 28580 1660 28589 1700
rect 28684 1660 29308 1700
rect 29348 1660 29357 1700
rect 29452 1660 29692 1700
rect 29732 1660 29741 1700
rect 29836 1660 30460 1700
rect 30500 1660 30509 1700
rect 30604 1660 31228 1700
rect 31268 1660 31277 1700
rect 31372 1660 31612 1700
rect 31652 1660 31661 1700
rect 44371 1660 44380 1700
rect 44420 1660 45388 1700
rect 45428 1660 45437 1700
rect 25612 1616 25652 1660
rect 26188 1616 26228 1660
rect 26764 1616 26804 1660
rect 27532 1616 27572 1660
rect 28300 1616 28340 1660
rect 28684 1616 28724 1660
rect 29452 1616 29492 1660
rect 29836 1616 29876 1660
rect 30604 1616 30644 1660
rect 31372 1616 31412 1660
rect 20044 1576 24116 1616
rect 25027 1576 25036 1616
rect 25076 1576 25652 1616
rect 25795 1576 25804 1616
rect 25844 1576 26228 1616
rect 26563 1576 26572 1616
rect 26612 1576 26804 1616
rect 27331 1576 27340 1616
rect 27380 1576 27572 1616
rect 27715 1576 27724 1616
rect 27764 1576 28340 1616
rect 28483 1576 28492 1616
rect 28532 1576 28724 1616
rect 28867 1576 28876 1616
rect 28916 1576 29492 1616
rect 29635 1576 29644 1616
rect 29684 1576 29876 1616
rect 30403 1576 30412 1616
rect 30452 1576 30644 1616
rect 30787 1576 30796 1616
rect 30836 1576 31412 1616
rect 4919 1492 4928 1532
rect 4968 1492 5010 1532
rect 5050 1492 5092 1532
rect 5132 1492 5174 1532
rect 5214 1492 5256 1532
rect 5296 1492 5305 1532
rect 20039 1492 20048 1532
rect 20088 1492 20130 1532
rect 20170 1492 20212 1532
rect 20252 1492 20294 1532
rect 20334 1492 20376 1532
rect 20416 1492 20425 1532
rect 24355 1492 24364 1532
rect 24404 1492 26476 1532
rect 26516 1492 26525 1532
rect 35159 1492 35168 1532
rect 35208 1492 35250 1532
rect 35290 1492 35332 1532
rect 35372 1492 35414 1532
rect 35454 1492 35496 1532
rect 35536 1492 35545 1532
rect 0 1448 90 1468
rect 46278 1448 46368 1468
rect 0 1408 1420 1448
rect 1460 1408 1469 1448
rect 45667 1408 45676 1448
rect 45716 1408 46368 1448
rect 0 1388 90 1408
rect 46278 1388 46368 1408
rect 0 1112 90 1132
rect 46278 1112 46368 1132
rect 0 1072 8140 1112
rect 8180 1072 8189 1112
rect 44611 1072 44620 1112
rect 44660 1072 46368 1112
rect 0 1052 90 1072
rect 46278 1052 46368 1072
rect 0 776 90 796
rect 46278 776 46368 796
rect 0 736 460 776
rect 500 736 509 776
rect 45379 736 45388 776
rect 45428 736 46368 776
rect 0 716 90 736
rect 46278 716 46368 736
<< via2 >>
rect 364 11152 404 11192
rect 44044 11152 44084 11192
rect 21484 10900 21524 10940
rect 21292 10816 21332 10856
rect 26380 10816 26420 10856
rect 42412 10816 42452 10856
rect 4928 10564 4968 10604
rect 5010 10564 5050 10604
rect 5092 10564 5132 10604
rect 5174 10564 5214 10604
rect 5256 10564 5296 10604
rect 17068 10732 17108 10772
rect 31180 10732 31220 10772
rect 19180 10648 19220 10688
rect 31468 10648 31508 10688
rect 40204 10648 40244 10688
rect 20048 10564 20088 10604
rect 20130 10564 20170 10604
rect 20212 10564 20252 10604
rect 20294 10564 20334 10604
rect 20376 10564 20416 10604
rect 26764 10564 26804 10604
rect 35168 10564 35208 10604
rect 35250 10564 35290 10604
rect 35332 10564 35372 10604
rect 35414 10564 35454 10604
rect 35496 10564 35536 10604
rect 23500 10480 23540 10520
rect 30220 10480 30260 10520
rect 40300 10480 40340 10520
rect 43180 10480 43220 10520
rect 44428 10480 44468 10520
rect 1996 10396 2036 10436
rect 4108 10396 4148 10436
rect 6220 10396 6260 10436
rect 8332 10396 8372 10436
rect 10444 10396 10484 10436
rect 12556 10396 12596 10436
rect 14668 10396 14708 10436
rect 16780 10396 16820 10436
rect 18892 10396 18932 10436
rect 21004 10396 21044 10436
rect 23116 10396 23156 10436
rect 25228 10396 25268 10436
rect 27340 10396 27380 10436
rect 29452 10396 29492 10436
rect 31564 10396 31604 10436
rect 33676 10396 33716 10436
rect 35788 10396 35828 10436
rect 37900 10396 37940 10436
rect 40012 10396 40052 10436
rect 42124 10396 42164 10436
rect 44236 10396 44276 10436
rect 20524 10312 20564 10352
rect 23308 10312 23348 10352
rect 25900 10312 25940 10352
rect 28396 10312 28436 10352
rect 16972 10228 17012 10268
rect 25036 10228 25076 10268
rect 28876 10228 28916 10268
rect 6220 10144 6260 10184
rect 6508 10144 6548 10184
rect 8620 10144 8660 10184
rect 17068 10144 17108 10184
rect 19180 10144 19220 10184
rect 23308 10144 23348 10184
rect 27244 10144 27284 10184
rect 27628 10144 27668 10184
rect 28780 10144 28820 10184
rect 34540 10144 34580 10184
rect 7180 10060 7220 10100
rect 13036 10060 13076 10100
rect 26860 10060 26900 10100
rect 28108 10060 28148 10100
rect 35596 10060 35636 10100
rect 40204 10144 40244 10184
rect 42412 10144 42452 10184
rect 43180 10144 43220 10184
rect 43564 10144 43604 10184
rect 43948 10144 43988 10184
rect 44524 10144 44564 10184
rect 44908 10144 44948 10184
rect 40396 10060 40436 10100
rect 24556 9976 24596 10016
rect 45772 9976 45812 10016
rect 1324 9892 1364 9932
rect 27724 9892 27764 9932
rect 27916 9892 27956 9932
rect 32140 9892 32180 9932
rect 3688 9808 3728 9848
rect 3770 9808 3810 9848
rect 3852 9808 3892 9848
rect 3934 9808 3974 9848
rect 4016 9808 4056 9848
rect 18808 9808 18848 9848
rect 18890 9808 18930 9848
rect 18972 9808 19012 9848
rect 19054 9808 19094 9848
rect 19136 9808 19176 9848
rect 23116 9808 23156 9848
rect 30796 9808 30836 9848
rect 33928 9808 33968 9848
rect 34010 9808 34050 9848
rect 34092 9808 34132 9848
rect 34174 9808 34214 9848
rect 34256 9808 34296 9848
rect 22444 9724 22484 9764
rect 27148 9724 27188 9764
rect 33100 9724 33140 9764
rect 30220 9640 30260 9680
rect 44428 9640 44468 9680
rect 23212 9556 23252 9596
rect 38092 9556 38132 9596
rect 44044 9556 44084 9596
rect 1228 9472 1268 9512
rect 22636 9472 22676 9512
rect 30604 9472 30644 9512
rect 30892 9472 30932 9512
rect 33484 9472 33524 9512
rect 43756 9472 43796 9512
rect 45772 9472 45812 9512
rect 18988 9388 19028 9428
rect 27916 9388 27956 9428
rect 28300 9388 28340 9428
rect 33772 9388 33812 9428
rect 43564 9388 43604 9428
rect 25900 9304 25940 9344
rect 29068 9304 29108 9344
rect 30796 9304 30836 9344
rect 38188 9304 38228 9344
rect 28012 9220 28052 9260
rect 37996 9220 38036 9260
rect 45772 9220 45812 9260
rect 23596 9136 23636 9176
rect 26092 9136 26132 9176
rect 32332 9136 32372 9176
rect 4928 9052 4968 9092
rect 5010 9052 5050 9092
rect 5092 9052 5132 9092
rect 5174 9052 5214 9092
rect 5256 9052 5296 9092
rect 20048 9052 20088 9092
rect 20130 9052 20170 9092
rect 20212 9052 20252 9092
rect 20294 9052 20334 9092
rect 20376 9052 20416 9092
rect 20524 9052 20564 9092
rect 22924 9052 22964 9092
rect 35168 9052 35208 9092
rect 35250 9052 35290 9092
rect 35332 9052 35372 9092
rect 35414 9052 35454 9092
rect 35496 9052 35536 9092
rect 23500 8968 23540 9008
rect 38188 8968 38228 9008
rect 44524 8968 44564 9008
rect 6508 8884 6548 8924
rect 7180 8884 7220 8924
rect 13036 8884 13076 8924
rect 16972 8884 17012 8924
rect 22156 8884 22196 8924
rect 23116 8884 23156 8924
rect 25036 8884 25076 8924
rect 26860 8884 26900 8924
rect 27244 8884 27284 8924
rect 27628 8884 27668 8924
rect 28780 8884 28820 8924
rect 29068 8884 29108 8924
rect 30604 8884 30644 8924
rect 43948 8884 43988 8924
rect 76 8800 116 8840
rect 10060 8800 10100 8840
rect 24556 8800 24596 8840
rect 28012 8800 28052 8840
rect 30892 8800 30932 8840
rect 31180 8800 31220 8840
rect 45772 8800 45812 8840
rect 6220 8716 6260 8756
rect 8620 8716 8660 8756
rect 8908 8716 8948 8756
rect 37996 8716 38036 8756
rect 6412 8632 6452 8672
rect 6892 8632 6932 8672
rect 7468 8632 7508 8672
rect 8812 8632 8852 8672
rect 14380 8632 14420 8672
rect 18988 8632 19028 8672
rect 21292 8632 21332 8672
rect 21868 8632 21908 8672
rect 22444 8632 22484 8672
rect 22636 8632 22676 8672
rect 22924 8632 22964 8672
rect 23596 8632 23636 8672
rect 26092 8632 26132 8672
rect 27148 8632 27188 8672
rect 27724 8632 27764 8672
rect 28300 8632 28340 8672
rect 32716 8632 32756 8672
rect 33388 8632 33428 8672
rect 38092 8632 38132 8672
rect 46252 8632 46292 8672
rect 31468 8548 31508 8588
rect 32524 8548 32564 8588
rect 23212 8464 23252 8504
rect 32908 8464 32948 8504
rect 364 8380 404 8420
rect 26284 8380 26324 8420
rect 3688 8296 3728 8336
rect 3770 8296 3810 8336
rect 3852 8296 3892 8336
rect 3934 8296 3974 8336
rect 4016 8296 4056 8336
rect 15820 8296 15860 8336
rect 18604 8296 18644 8336
rect 18808 8296 18848 8336
rect 18890 8296 18930 8336
rect 18972 8296 19012 8336
rect 19054 8296 19094 8336
rect 19136 8296 19176 8336
rect 33928 8296 33968 8336
rect 34010 8296 34050 8336
rect 34092 8296 34132 8336
rect 34174 8296 34214 8336
rect 34256 8296 34296 8336
rect 15628 8212 15668 8252
rect 17740 8212 17780 8252
rect 25900 8212 25940 8252
rect 28780 8212 28820 8252
rect 1324 8128 1364 8168
rect 15244 8128 15284 8168
rect 28108 8128 28148 8168
rect 28876 8128 28916 8168
rect 46252 8128 46292 8168
rect 1228 8044 1268 8084
rect 16588 8044 16628 8084
rect 16780 8044 16820 8084
rect 14860 7960 14900 8000
rect 17356 7960 17396 8000
rect 17740 7960 17780 8000
rect 18604 7960 18644 8000
rect 15052 7876 15092 7916
rect 30988 8044 31028 8084
rect 44908 8044 44948 8084
rect 26284 7960 26324 8000
rect 33580 7960 33620 8000
rect 8908 7792 8948 7832
rect 16012 7792 16052 7832
rect 27724 7792 27764 7832
rect 17068 7708 17108 7748
rect 17452 7708 17492 7748
rect 17836 7708 17876 7748
rect 27916 7876 27956 7916
rect 43756 7876 43796 7916
rect 44524 7960 44564 8000
rect 30988 7792 31028 7832
rect 33676 7708 33716 7748
rect 25420 7624 25460 7664
rect 46252 7624 46292 7664
rect 4928 7540 4968 7580
rect 5010 7540 5050 7580
rect 5092 7540 5132 7580
rect 5174 7540 5214 7580
rect 5256 7540 5296 7580
rect 20048 7540 20088 7580
rect 20130 7540 20170 7580
rect 20212 7540 20252 7580
rect 20294 7540 20334 7580
rect 20376 7540 20416 7580
rect 26668 7540 26708 7580
rect 35168 7540 35208 7580
rect 35250 7540 35290 7580
rect 35332 7540 35372 7580
rect 35414 7540 35454 7580
rect 35496 7540 35536 7580
rect 17836 7456 17876 7496
rect 26860 7456 26900 7496
rect 46252 7456 46292 7496
rect 17452 7372 17492 7412
rect 25516 7372 25556 7412
rect 25900 7372 25940 7412
rect 27244 7372 27284 7412
rect 17068 7288 17108 7328
rect 25228 7288 25268 7328
rect 15436 7204 15476 7244
rect 17356 7204 17396 7244
rect 1420 7120 1460 7160
rect 13516 7120 13556 7160
rect 13708 7120 13748 7160
rect 17068 7120 17108 7160
rect 17740 7120 17780 7160
rect 18700 7120 18740 7160
rect 19276 7120 19316 7160
rect 19660 7120 19700 7160
rect 19852 7120 19892 7160
rect 20236 7120 20276 7160
rect 20716 7120 20756 7160
rect 21196 7120 21236 7160
rect 23980 7120 24020 7160
rect 27340 7120 27380 7160
rect 13900 7036 13940 7076
rect 1132 6784 1172 6824
rect 3688 6784 3728 6824
rect 3770 6784 3810 6824
rect 3852 6784 3892 6824
rect 3934 6784 3974 6824
rect 4016 6784 4056 6824
rect 940 6448 980 6488
rect 13324 6448 13364 6488
rect 16108 6952 16148 6992
rect 14092 6868 14132 6908
rect 16300 7036 16340 7076
rect 18220 7036 18260 7076
rect 23212 7036 23252 7076
rect 43180 7036 43220 7076
rect 17452 6952 17492 6992
rect 17836 6952 17876 6992
rect 18124 6952 18164 6992
rect 18604 6952 18644 6992
rect 19372 6952 19412 6992
rect 19948 6952 19988 6992
rect 14284 6784 14324 6824
rect 16396 6784 16436 6824
rect 18220 6784 18260 6824
rect 18808 6784 18848 6824
rect 18890 6784 18930 6824
rect 18972 6784 19012 6824
rect 19054 6784 19094 6824
rect 19136 6784 19176 6824
rect 24268 6952 24308 6992
rect 46252 6952 46292 6992
rect 20812 6868 20852 6908
rect 24172 6868 24212 6908
rect 25804 6784 25844 6824
rect 33928 6784 33968 6824
rect 34010 6784 34050 6824
rect 34092 6784 34132 6824
rect 34174 6784 34214 6824
rect 34256 6784 34296 6824
rect 46252 6784 46292 6824
rect 14476 6700 14516 6740
rect 17068 6700 17108 6740
rect 17836 6700 17876 6740
rect 23788 6700 23828 6740
rect 16588 6616 16628 6656
rect 18700 6616 18740 6656
rect 19372 6616 19412 6656
rect 25612 6616 25652 6656
rect 34540 6616 34580 6656
rect 14668 6532 14708 6572
rect 17740 6532 17780 6572
rect 20044 6532 20084 6572
rect 23308 6532 23348 6572
rect 16780 6448 16820 6488
rect 19276 6448 19316 6488
rect 20332 6448 20372 6488
rect 20908 6448 20948 6488
rect 22540 6448 22580 6488
rect 33196 6448 33236 6488
rect 16972 6364 17012 6404
rect 19660 6364 19700 6404
rect 20812 6364 20852 6404
rect 24844 6364 24884 6404
rect 28588 6364 28628 6404
rect 44620 6364 44660 6404
rect 18412 6280 18452 6320
rect 18604 6280 18644 6320
rect 21004 6280 21044 6320
rect 25708 6280 25748 6320
rect 34444 6280 34484 6320
rect 17548 6196 17588 6236
rect 17740 6196 17780 6236
rect 20236 6196 20276 6236
rect 24076 6196 24116 6236
rect 41740 6196 41780 6236
rect 556 6112 596 6152
rect 4928 6028 4968 6068
rect 5010 6028 5050 6068
rect 5092 6028 5132 6068
rect 5174 6028 5214 6068
rect 5256 6028 5296 6068
rect 17452 6112 17492 6152
rect 23596 6112 23636 6152
rect 17164 6028 17204 6068
rect 19852 6028 19892 6068
rect 20048 6028 20088 6068
rect 20130 6028 20170 6068
rect 20212 6028 20252 6068
rect 20294 6028 20334 6068
rect 20376 6028 20416 6068
rect 20524 6028 20564 6068
rect 21964 6028 22004 6068
rect 35168 6028 35208 6068
rect 35250 6028 35290 6068
rect 35332 6028 35372 6068
rect 35414 6028 35454 6068
rect 35496 6028 35536 6068
rect 18700 5944 18740 5984
rect 19948 5944 19988 5984
rect 25132 5944 25172 5984
rect 15916 5860 15956 5900
rect 17548 5860 17588 5900
rect 20716 5860 20756 5900
rect 1036 5776 1076 5816
rect 16204 5776 16244 5816
rect 17356 5776 17396 5816
rect 21196 5776 21236 5816
rect 21580 5776 21620 5816
rect 22732 5776 22772 5816
rect 11788 5692 11828 5732
rect 12076 5692 12116 5732
rect 12556 5692 12596 5732
rect 12748 5692 12788 5732
rect 6700 5608 6740 5648
rect 10540 5608 10580 5648
rect 10828 5608 10868 5648
rect 12652 5608 12692 5648
rect 13132 5608 13172 5648
rect 15916 5608 15956 5648
rect 20332 5608 20372 5648
rect 20524 5608 20564 5648
rect 29932 5608 29972 5648
rect 8620 5524 8660 5564
rect 9964 5524 10004 5564
rect 11500 5524 11540 5564
rect 20716 5524 20756 5564
rect 21484 5524 21524 5564
rect 28972 5524 29012 5564
rect 844 5440 884 5480
rect 8716 5440 8756 5480
rect 12172 5440 12212 5480
rect 20908 5440 20948 5480
rect 23116 5440 23156 5480
rect 28876 5440 28916 5480
rect 8140 5356 8180 5396
rect 10060 5356 10100 5396
rect 19948 5356 19988 5396
rect 21292 5356 21332 5396
rect 38572 5692 38612 5732
rect 43084 5692 43124 5732
rect 34348 5608 34388 5648
rect 36940 5608 36980 5648
rect 37612 5608 37652 5648
rect 37900 5608 37940 5648
rect 43852 5608 43892 5648
rect 38092 5440 38132 5480
rect 22252 5356 22292 5396
rect 29356 5356 29396 5396
rect 3688 5272 3728 5312
rect 3770 5272 3810 5312
rect 3852 5272 3892 5312
rect 3934 5272 3974 5312
rect 4016 5272 4056 5312
rect 8620 5272 8660 5312
rect 9676 5272 9716 5312
rect 9964 5272 10004 5312
rect 11692 5272 11732 5312
rect 12748 5272 12788 5312
rect 18808 5272 18848 5312
rect 18890 5272 18930 5312
rect 18972 5272 19012 5312
rect 19054 5272 19094 5312
rect 19136 5272 19176 5312
rect 29548 5272 29588 5312
rect 33928 5272 33968 5312
rect 34010 5272 34050 5312
rect 34092 5272 34132 5312
rect 34174 5272 34214 5312
rect 34256 5272 34296 5312
rect 41068 5524 41108 5564
rect 44140 5440 44180 5480
rect 44332 5356 44372 5396
rect 4780 5188 4820 5228
rect 12172 5188 12212 5228
rect 21388 5188 21428 5228
rect 44716 5188 44756 5228
rect 1324 5104 1364 5144
rect 748 5020 788 5060
rect 23116 5020 23156 5060
rect 26956 5020 26996 5060
rect 31660 5020 31700 5060
rect 1420 4936 1460 4976
rect 7180 4936 7220 4976
rect 7564 4936 7604 4976
rect 11596 4936 11636 4976
rect 11788 4936 11828 4976
rect 15916 4936 15956 4976
rect 19852 4936 19892 4976
rect 22252 4936 22292 4976
rect 22924 4936 22964 4976
rect 11308 4852 11348 4892
rect 11500 4852 11540 4892
rect 18700 4852 18740 4892
rect 19660 4852 19700 4892
rect 38572 5020 38612 5060
rect 23404 4936 23444 4976
rect 34348 4936 34388 4976
rect 41068 5104 41108 5144
rect 41356 5104 41396 5144
rect 40876 5020 40916 5060
rect 44236 5020 44276 5060
rect 27820 4852 27860 4892
rect 38092 4852 38132 4892
rect 39052 4852 39092 4892
rect 8332 4684 8372 4724
rect 15148 4684 15188 4724
rect 16204 4684 16244 4724
rect 21676 4684 21716 4724
rect 23020 4684 23060 4724
rect 26956 4684 26996 4724
rect 10060 4600 10100 4640
rect 10636 4600 10676 4640
rect 10828 4600 10868 4640
rect 12556 4600 12596 4640
rect 19468 4600 19508 4640
rect 22924 4600 22964 4640
rect 31276 4684 31316 4724
rect 30796 4600 30836 4640
rect 37612 4684 37652 4724
rect 39340 4684 39371 4724
rect 39371 4684 39380 4724
rect 44044 4852 44084 4892
rect 41260 4768 41300 4808
rect 44428 4768 44468 4808
rect 40108 4684 40139 4724
rect 40139 4684 40148 4724
rect 40300 4684 40340 4724
rect 37420 4600 37460 4640
rect 4928 4516 4968 4556
rect 5010 4516 5050 4556
rect 5092 4516 5132 4556
rect 5174 4516 5214 4556
rect 5256 4516 5296 4556
rect 8428 4516 8468 4556
rect 18220 4516 18260 4556
rect 18700 4516 18740 4556
rect 19756 4516 19796 4556
rect 20048 4516 20088 4556
rect 20130 4516 20170 4556
rect 20212 4516 20252 4556
rect 20294 4516 20334 4556
rect 20376 4516 20416 4556
rect 21580 4516 21620 4556
rect 22636 4516 22676 4556
rect 30220 4516 30260 4556
rect 35168 4516 35208 4556
rect 35250 4516 35290 4556
rect 35332 4516 35372 4556
rect 35414 4516 35454 4556
rect 35496 4516 35536 4556
rect 35980 4516 36020 4556
rect 41356 4516 41396 4556
rect 1420 4432 1460 4472
rect 7564 4432 7604 4472
rect 11404 4432 11444 4472
rect 19564 4432 19604 4472
rect 23404 4432 23444 4472
rect 28012 4432 28052 4472
rect 28204 4432 28244 4472
rect 7180 4348 7220 4388
rect 11212 4348 11252 4388
rect 18316 4348 18356 4388
rect 22828 4348 22868 4388
rect 26956 4348 26996 4388
rect 30700 4348 30740 4388
rect 30892 4348 30932 4388
rect 34828 4348 34868 4388
rect 39340 4348 39371 4388
rect 39371 4348 39380 4388
rect 40300 4348 40340 4388
rect 37996 4264 38036 4304
rect 1132 4180 1172 4220
rect 23116 4180 23156 4220
rect 27052 4180 27092 4220
rect 28492 4180 28532 4220
rect 35596 4180 35636 4220
rect 38092 4180 38132 4220
rect 41260 4180 41300 4220
rect 11020 4096 11060 4136
rect 19372 4096 19412 4136
rect 24460 4096 24500 4136
rect 25324 4096 25364 4136
rect 25996 4096 26036 4136
rect 44524 4096 44564 4136
rect 44908 4096 44948 4136
rect 844 4012 884 4052
rect 24940 4012 24980 4052
rect 25900 4012 25940 4052
rect 27436 4012 27476 4052
rect 30892 4012 30932 4052
rect 940 3928 980 3968
rect 5932 3928 5972 3968
rect 10156 3928 10196 3968
rect 10348 3928 10388 3968
rect 19276 3928 19316 3968
rect 26188 3928 26228 3968
rect 37324 4012 37364 4052
rect 43852 4012 43892 4052
rect 1036 3844 1076 3884
rect 10060 3844 10100 3884
rect 10444 3844 10484 3884
rect 27532 3844 27572 3884
rect 37132 3844 37172 3884
rect 38092 3844 38132 3884
rect 3688 3760 3728 3800
rect 3770 3760 3810 3800
rect 3852 3760 3892 3800
rect 3934 3760 3974 3800
rect 4016 3760 4056 3800
rect 10252 3760 10292 3800
rect 18808 3760 18848 3800
rect 18890 3760 18930 3800
rect 18972 3760 19012 3800
rect 19054 3760 19094 3800
rect 19136 3760 19176 3800
rect 19276 3760 19316 3800
rect 27628 3760 27668 3800
rect 33928 3760 33968 3800
rect 34010 3760 34050 3800
rect 34092 3760 34132 3800
rect 34174 3760 34214 3800
rect 34256 3760 34296 3800
rect 5932 3676 5972 3716
rect 37420 3676 37460 3716
rect 1324 3592 1364 3632
rect 26764 3592 26804 3632
rect 27532 3592 27572 3632
rect 28204 3592 28244 3632
rect 1420 3508 1460 3548
rect 20140 3508 20180 3548
rect 23116 3508 23156 3548
rect 24748 3424 24788 3464
rect 25996 3424 26036 3464
rect 44524 3592 44564 3632
rect 30124 3508 30164 3548
rect 26764 3424 26804 3464
rect 27052 3424 27092 3464
rect 27436 3424 27476 3464
rect 27820 3424 27860 3464
rect 28204 3424 28244 3464
rect 28588 3424 28628 3464
rect 30892 3424 30932 3464
rect 34444 3424 34484 3464
rect 34828 3424 34868 3464
rect 35980 3424 36020 3464
rect 10156 3340 10196 3380
rect 18700 3340 18740 3380
rect 37996 3424 38036 3464
rect 41068 3424 41108 3464
rect 44044 3340 44084 3380
rect 19564 3256 19604 3296
rect 24460 3256 24500 3296
rect 27916 3256 27956 3296
rect 44908 3256 44948 3296
rect 18988 3172 19028 3212
rect 25324 3172 25364 3212
rect 26380 3172 26420 3212
rect 28396 3172 28436 3212
rect 34732 3172 34772 3212
rect 4780 3088 4820 3128
rect 18508 3088 18548 3128
rect 26188 3088 26228 3128
rect 27340 3088 27380 3128
rect 27820 3088 27860 3128
rect 35020 3088 35060 3128
rect 44620 3088 44660 3128
rect 4928 3004 4968 3044
rect 5010 3004 5050 3044
rect 5092 3004 5132 3044
rect 5174 3004 5214 3044
rect 5256 3004 5296 3044
rect 20048 3004 20088 3044
rect 20130 3004 20170 3044
rect 20212 3004 20252 3044
rect 20294 3004 20334 3044
rect 20376 3004 20416 3044
rect 24940 3004 24980 3044
rect 26092 3004 26132 3044
rect 26764 3004 26804 3044
rect 34636 3004 34676 3044
rect 35168 3004 35208 3044
rect 35250 3004 35290 3044
rect 35332 3004 35372 3044
rect 35414 3004 35454 3044
rect 35496 3004 35536 3044
rect 556 2920 596 2960
rect 28204 2920 28244 2960
rect 9676 2836 9716 2876
rect 22828 2836 22868 2876
rect 23020 2836 23060 2876
rect 25132 2836 25172 2876
rect 25516 2836 25556 2876
rect 34828 2836 34868 2876
rect 1420 2752 1460 2792
rect 8716 2752 8756 2792
rect 11308 2668 11348 2708
rect 21964 2668 22004 2708
rect 15148 2584 15188 2624
rect 22636 2584 22676 2624
rect 19180 2500 19220 2540
rect 20044 2500 20084 2540
rect 20908 2500 20948 2540
rect 1420 2416 1460 2456
rect 19084 2416 19124 2456
rect 21196 2416 21236 2456
rect 21580 2416 21620 2456
rect 21964 2416 22004 2456
rect 22348 2416 22388 2456
rect 22732 2416 22772 2456
rect 25420 2752 25460 2792
rect 25708 2752 25748 2792
rect 24460 2668 24500 2708
rect 25804 2668 25844 2708
rect 27148 2668 27188 2708
rect 27916 2752 27956 2792
rect 28012 2668 28052 2708
rect 30220 2668 30260 2708
rect 44236 2668 44276 2708
rect 23980 2584 24020 2624
rect 28396 2584 28436 2624
rect 28972 2584 29012 2624
rect 29356 2584 29396 2624
rect 31276 2584 31316 2624
rect 44140 2584 44180 2624
rect 44524 2584 44564 2624
rect 24940 2500 24980 2540
rect 25324 2500 25364 2540
rect 29164 2500 29204 2540
rect 23116 2416 23156 2456
rect 23500 2416 23540 2456
rect 25228 2416 25268 2456
rect 25612 2416 25652 2456
rect 25996 2416 26036 2456
rect 26380 2416 26420 2456
rect 26764 2416 26804 2456
rect 27148 2416 27188 2456
rect 27532 2416 27572 2456
rect 27916 2416 27956 2456
rect 28300 2416 28340 2456
rect 28684 2416 28724 2456
rect 29068 2416 29108 2456
rect 29452 2416 29492 2456
rect 29836 2416 29876 2456
rect 30220 2416 30260 2456
rect 30604 2416 30644 2456
rect 30988 2416 31028 2456
rect 45676 2416 45716 2456
rect 19756 2332 19796 2372
rect 23308 2332 23348 2372
rect 25132 2332 25172 2372
rect 3688 2248 3728 2288
rect 3770 2248 3810 2288
rect 3852 2248 3892 2288
rect 3934 2248 3974 2288
rect 4016 2248 4056 2288
rect 18808 2248 18848 2288
rect 18890 2248 18930 2288
rect 18972 2248 19012 2288
rect 19054 2248 19094 2288
rect 19136 2248 19176 2288
rect 24556 2248 24596 2288
rect 33928 2248 33968 2288
rect 34010 2248 34050 2288
rect 34092 2248 34132 2288
rect 34174 2248 34214 2288
rect 34256 2248 34296 2288
rect 16204 2164 16244 2204
rect 748 2080 788 2120
rect 15916 2080 15956 2120
rect 18604 1996 18644 2036
rect 21388 1996 21428 2036
rect 22540 1996 22580 2036
rect 25708 2164 25748 2204
rect 27052 2164 27092 2204
rect 27340 2164 27380 2204
rect 26668 2080 26708 2120
rect 28876 2080 28916 2120
rect 24652 1996 24692 2036
rect 25420 1996 25460 2036
rect 18220 1912 18260 1952
rect 21676 1912 21716 1952
rect 22828 1912 22868 1952
rect 23596 1912 23636 1952
rect 23788 1912 23828 1952
rect 24940 1912 24980 1952
rect 26188 1996 26228 2036
rect 28108 1996 28148 2036
rect 29260 1996 29300 2036
rect 41740 1996 41780 2036
rect 26476 1912 26516 1952
rect 27052 1912 27092 1952
rect 27436 1912 27476 1952
rect 28780 1912 28820 1952
rect 29548 1912 29588 1952
rect 29932 1912 29972 1952
rect 30700 1912 30740 1952
rect 31660 1912 31700 1952
rect 39052 1912 39092 1952
rect 44428 1912 44468 1952
rect 44716 1912 44756 1952
rect 26860 1828 26900 1868
rect 28492 1828 28532 1868
rect 1420 1744 1460 1784
rect 20044 1660 20084 1700
rect 21388 1660 21428 1700
rect 21772 1660 21812 1700
rect 22156 1660 22196 1700
rect 22540 1660 22580 1700
rect 22924 1660 22964 1700
rect 23308 1660 23348 1700
rect 23692 1660 23732 1700
rect 23884 1660 23924 1700
rect 24172 1744 24212 1784
rect 24652 1744 24692 1784
rect 25420 1744 25460 1784
rect 26956 1744 26996 1784
rect 28108 1744 28148 1784
rect 30028 1744 30068 1784
rect 44620 1744 44660 1784
rect 24268 1660 24308 1700
rect 24460 1660 24500 1700
rect 24844 1660 24884 1700
rect 45388 1660 45428 1700
rect 25036 1576 25076 1616
rect 25804 1576 25844 1616
rect 26572 1576 26612 1616
rect 27340 1576 27380 1616
rect 27724 1576 27764 1616
rect 28492 1576 28532 1616
rect 28876 1576 28916 1616
rect 29644 1576 29684 1616
rect 30412 1576 30452 1616
rect 30796 1576 30836 1616
rect 4928 1492 4968 1532
rect 5010 1492 5050 1532
rect 5092 1492 5132 1532
rect 5174 1492 5214 1532
rect 5256 1492 5296 1532
rect 20048 1492 20088 1532
rect 20130 1492 20170 1532
rect 20212 1492 20252 1532
rect 20294 1492 20334 1532
rect 20376 1492 20416 1532
rect 24364 1492 24404 1532
rect 26476 1492 26516 1532
rect 35168 1492 35208 1532
rect 35250 1492 35290 1532
rect 35332 1492 35372 1532
rect 35414 1492 35454 1532
rect 35496 1492 35536 1532
rect 1420 1408 1460 1448
rect 45676 1408 45716 1448
rect 8140 1072 8180 1112
rect 44620 1072 44660 1112
rect 460 736 500 776
rect 45388 736 45428 776
<< metal3 >>
rect 1976 12100 2056 12180
rect 4088 12100 4168 12180
rect 6200 12100 6280 12180
rect 8312 12100 8392 12180
rect 10424 12100 10504 12180
rect 12536 12100 12616 12180
rect 14648 12100 14728 12180
rect 16760 12100 16840 12180
rect 18872 12100 18952 12180
rect 20984 12100 21064 12180
rect 23096 12100 23176 12180
rect 25208 12100 25288 12180
rect 27320 12100 27400 12180
rect 29432 12100 29512 12180
rect 31544 12100 31624 12180
rect 33656 12100 33736 12180
rect 35768 12100 35848 12180
rect 37880 12100 37960 12180
rect 39992 12100 40072 12180
rect 42104 12100 42184 12180
rect 44216 12100 44296 12180
rect 364 11192 404 11201
rect 76 8840 116 8849
rect 76 8705 116 8800
rect 364 8420 404 11152
rect 1996 10436 2036 12100
rect 1996 10387 2036 10396
rect 4108 10436 4148 12100
rect 4928 10604 5296 10613
rect 4968 10564 5010 10604
rect 5050 10564 5092 10604
rect 5132 10564 5174 10604
rect 5214 10564 5256 10604
rect 4928 10555 5296 10564
rect 4108 10387 4148 10396
rect 6220 10436 6260 12100
rect 6220 10387 6260 10396
rect 8332 10436 8372 12100
rect 8332 10387 8372 10396
rect 10444 10436 10484 12100
rect 10444 10387 10484 10396
rect 12556 10436 12596 12100
rect 12556 10387 12596 10396
rect 14668 10436 14708 12100
rect 14668 10387 14708 10396
rect 16780 10436 16820 12100
rect 16780 10387 16820 10396
rect 17068 10772 17108 10781
rect 16972 10268 17012 10277
rect 6220 10184 6260 10193
rect 1324 9932 1364 9941
rect 364 8371 404 8380
rect 1228 9512 1268 9521
rect 1228 8084 1268 9472
rect 1324 8168 1364 9892
rect 3688 9848 4056 9857
rect 3728 9808 3770 9848
rect 3810 9808 3852 9848
rect 3892 9808 3934 9848
rect 3974 9808 4016 9848
rect 3688 9799 4056 9808
rect 4928 9092 5296 9101
rect 4968 9052 5010 9092
rect 5050 9052 5092 9092
rect 5132 9052 5174 9092
rect 5214 9052 5256 9092
rect 4928 9043 5296 9052
rect 6220 8756 6260 10144
rect 6508 10184 6548 10193
rect 6508 8924 6548 10144
rect 8620 10184 8660 10193
rect 6508 8875 6548 8884
rect 7180 10100 7220 10109
rect 7180 8924 7220 10060
rect 7180 8875 7220 8884
rect 6220 8707 6260 8716
rect 8620 8756 8660 10144
rect 13036 10100 13076 10109
rect 13036 8924 13076 10060
rect 13036 8875 13076 8884
rect 16972 8924 17012 10228
rect 17068 10184 17108 10732
rect 18892 10436 18932 12100
rect 18892 10387 18932 10396
rect 19180 10688 19220 10697
rect 17068 10135 17108 10144
rect 19180 10184 19220 10648
rect 20048 10604 20416 10613
rect 20088 10564 20130 10604
rect 20170 10564 20212 10604
rect 20252 10564 20294 10604
rect 20334 10564 20376 10604
rect 20048 10555 20416 10564
rect 21004 10436 21044 12100
rect 21484 10940 21524 10949
rect 21004 10387 21044 10396
rect 21292 10856 21332 10865
rect 19180 10135 19220 10144
rect 20524 10352 20564 10361
rect 18808 9848 19176 9857
rect 18848 9808 18890 9848
rect 18930 9808 18972 9848
rect 19012 9808 19054 9848
rect 19094 9808 19136 9848
rect 18808 9799 19176 9808
rect 16972 8875 17012 8884
rect 18988 9428 19028 9437
rect 10060 8840 10100 8849
rect 8620 8707 8660 8716
rect 8908 8756 8948 8765
rect 6412 8672 6452 8681
rect 3688 8336 4056 8345
rect 3728 8296 3770 8336
rect 3810 8296 3852 8336
rect 3892 8296 3934 8336
rect 3974 8296 4016 8336
rect 3688 8287 4056 8296
rect 1324 8119 1364 8128
rect 1228 8035 1268 8044
rect 4928 7580 5296 7589
rect 4968 7540 5010 7580
rect 5050 7540 5092 7580
rect 5132 7540 5174 7580
rect 5214 7540 5256 7580
rect 4928 7531 5296 7540
rect 1420 7160 1460 7169
rect 1132 6824 1172 6833
rect 460 6488 500 6497
rect 460 776 500 6448
rect 940 6488 980 6497
rect 556 6152 596 6161
rect 556 2960 596 6112
rect 844 5480 884 5489
rect 556 2911 596 2920
rect 748 5060 788 5069
rect 748 2120 788 5020
rect 844 4052 884 5440
rect 844 4003 884 4012
rect 940 3968 980 6448
rect 940 3919 980 3928
rect 1036 5816 1076 5825
rect 1036 3884 1076 5776
rect 1132 4220 1172 6784
rect 1132 4171 1172 4180
rect 1324 5144 1364 5153
rect 1036 3835 1076 3844
rect 1324 3632 1364 5104
rect 1420 4976 1460 7120
rect 3688 6824 4056 6833
rect 3728 6784 3770 6824
rect 3810 6784 3852 6824
rect 3892 6784 3934 6824
rect 3974 6784 4016 6824
rect 3688 6775 4056 6784
rect 4928 6068 5296 6077
rect 4968 6028 5010 6068
rect 5050 6028 5092 6068
rect 5132 6028 5174 6068
rect 5214 6028 5256 6068
rect 4928 6019 5296 6028
rect 3688 5312 4056 5321
rect 3728 5272 3770 5312
rect 3810 5272 3852 5312
rect 3892 5272 3934 5312
rect 3974 5272 4016 5312
rect 3688 5263 4056 5272
rect 1420 4927 1460 4936
rect 4780 5228 4820 5237
rect 1324 3583 1364 3592
rect 1420 4472 1460 4481
rect 1420 3548 1460 4432
rect 3688 3800 4056 3809
rect 3728 3760 3770 3800
rect 3810 3760 3852 3800
rect 3892 3760 3934 3800
rect 3974 3760 4016 3800
rect 3688 3751 4056 3760
rect 1420 3499 1460 3508
rect 4780 3128 4820 5188
rect 4928 4556 5296 4565
rect 4968 4516 5010 4556
rect 5050 4516 5092 4556
rect 5132 4516 5174 4556
rect 5214 4516 5256 4556
rect 4928 4507 5296 4516
rect 5932 3968 5972 3977
rect 5932 3716 5972 3928
rect 5932 3667 5972 3676
rect 4780 3079 4820 3088
rect 4928 3044 5296 3053
rect 4968 3004 5010 3044
rect 5050 3004 5092 3044
rect 5132 3004 5174 3044
rect 5214 3004 5256 3044
rect 4928 2995 5296 3004
rect 1420 2792 1460 2801
rect 1420 2657 1460 2752
rect 1420 2456 1460 2465
rect 1420 2321 1460 2416
rect 3688 2288 4056 2297
rect 3728 2248 3770 2288
rect 3810 2248 3852 2288
rect 3892 2248 3934 2288
rect 3974 2248 4016 2288
rect 3688 2239 4056 2248
rect 748 2071 788 2080
rect 1420 1784 1460 1793
rect 1420 1649 1460 1744
rect 4928 1532 5296 1541
rect 4968 1492 5010 1532
rect 5050 1492 5092 1532
rect 5132 1492 5174 1532
rect 5214 1492 5256 1532
rect 4928 1483 5296 1492
rect 1420 1448 1460 1457
rect 1420 1313 1460 1408
rect 460 727 500 736
rect 6412 188 6452 8632
rect 6892 8672 6932 8681
rect 6700 5648 6740 5657
rect 6700 4640 6740 5608
rect 6700 4591 6740 4600
rect 6892 272 6932 8632
rect 7468 8672 7508 8681
rect 7180 4976 7220 4985
rect 7180 4388 7220 4936
rect 7180 4339 7220 4348
rect 7468 356 7508 8632
rect 8812 8672 8852 8681
rect 8620 5564 8660 5573
rect 8140 5396 8180 5405
rect 7564 4976 7604 4985
rect 7564 4472 7604 4936
rect 7564 4423 7604 4432
rect 8140 1112 8180 5356
rect 8620 5312 8660 5524
rect 8620 5263 8660 5272
rect 8716 5480 8756 5489
rect 8332 4724 8372 4733
rect 8332 4556 8372 4684
rect 8428 4556 8468 4565
rect 8332 4516 8428 4556
rect 8428 4507 8468 4516
rect 8716 2792 8756 5440
rect 8716 2743 8756 2752
rect 8140 1063 8180 1072
rect 7468 307 7508 316
rect 6892 223 6932 232
rect 6412 139 6452 148
rect 8812 104 8852 8632
rect 8908 7832 8948 8716
rect 10060 8705 10100 8800
rect 8908 7783 8948 7792
rect 14380 8672 14420 8681
rect 13516 7160 13556 7169
rect 13324 6488 13364 6497
rect 11788 5732 11828 5741
rect 10540 5648 10580 5657
rect 9964 5564 10004 5573
rect 9676 5312 9716 5321
rect 9676 2876 9716 5272
rect 9964 5312 10004 5524
rect 10540 5513 10580 5608
rect 10828 5648 10868 5657
rect 9964 5263 10004 5272
rect 10060 5396 10100 5405
rect 10060 5261 10100 5356
rect 10060 4640 10100 4649
rect 10060 4505 10100 4600
rect 10636 4640 10676 4649
rect 10636 4052 10676 4600
rect 10828 4640 10868 5608
rect 11500 5564 11540 5573
rect 10828 4591 10868 4600
rect 11308 4892 11348 4901
rect 11212 4388 11252 4397
rect 10636 4003 10676 4012
rect 11020 4136 11060 4145
rect 10156 3968 10196 3977
rect 10060 3884 10100 3893
rect 10060 3749 10100 3844
rect 10156 3380 10196 3928
rect 10348 3968 10388 3977
rect 10252 3800 10292 3809
rect 10348 3800 10388 3928
rect 10292 3760 10388 3800
rect 10444 3884 10484 3893
rect 10252 3751 10292 3760
rect 10444 3749 10484 3844
rect 10156 3331 10196 3340
rect 9676 2827 9716 2836
rect 11020 80 11060 4096
rect 11212 80 11252 4348
rect 11308 2708 11348 4852
rect 11500 4892 11540 5524
rect 11692 5312 11732 5321
rect 11500 4843 11540 4852
rect 11596 4976 11636 4985
rect 11308 2659 11348 2668
rect 11404 4472 11444 4481
rect 11404 80 11444 4432
rect 11596 80 11636 4936
rect 11692 4220 11732 5272
rect 11788 4976 11828 5692
rect 12076 5732 12116 5741
rect 11788 4927 11828 4936
rect 11980 5648 12020 5657
rect 11692 4171 11732 4180
rect 11884 4136 11924 4145
rect 11692 4052 11732 4061
rect 11692 2624 11732 4012
rect 11788 3968 11828 3977
rect 11788 2708 11828 3928
rect 11884 2792 11924 4096
rect 11980 2876 12020 5608
rect 12076 3968 12116 5692
rect 12556 5732 12596 5741
rect 12172 5480 12212 5489
rect 12172 5228 12212 5440
rect 12172 5179 12212 5188
rect 12556 4808 12596 5692
rect 12748 5732 12788 5741
rect 12652 5648 12692 5657
rect 12652 5513 12692 5608
rect 12748 5312 12788 5692
rect 12940 5648 12980 5657
rect 13132 5648 13172 5657
rect 12980 5608 13076 5648
rect 12940 5580 12980 5608
rect 12748 5263 12788 5272
rect 12556 4768 12788 4808
rect 12076 3919 12116 3928
rect 12556 4640 12596 4649
rect 11980 2836 12404 2876
rect 11884 2752 12212 2792
rect 11788 2668 12020 2708
rect 11692 2584 11828 2624
rect 11788 80 11828 2584
rect 11980 80 12020 2668
rect 12172 80 12212 2752
rect 12364 80 12404 2836
rect 12556 80 12596 4600
rect 12748 80 12788 4768
rect 13036 440 13076 5608
rect 12940 400 13076 440
rect 12940 80 12980 400
rect 13132 80 13172 5608
rect 13324 80 13364 6448
rect 13516 80 13556 7120
rect 13708 7160 13748 7169
rect 13708 80 13748 7120
rect 13900 7076 13940 7085
rect 13900 80 13940 7036
rect 14092 6908 14132 6917
rect 14092 80 14132 6868
rect 14284 6824 14324 6833
rect 14284 80 14324 6784
rect 14380 440 14420 8632
rect 18988 8672 19028 9388
rect 20048 9092 20416 9101
rect 20088 9052 20130 9092
rect 20170 9052 20212 9092
rect 20252 9052 20294 9092
rect 20334 9052 20376 9092
rect 20048 9043 20416 9052
rect 20524 9092 20564 10312
rect 20524 9043 20564 9052
rect 18988 8623 19028 8632
rect 21292 8672 21332 10816
rect 21484 8672 21524 10900
rect 23116 10436 23156 12100
rect 23116 10387 23156 10396
rect 23500 10520 23540 10529
rect 23308 10352 23348 10361
rect 23308 10184 23348 10312
rect 23308 10135 23348 10144
rect 23116 9848 23156 9857
rect 22444 9764 22484 9773
rect 22156 9680 22196 9689
rect 22156 8924 22196 9640
rect 22156 8875 22196 8884
rect 21868 8672 21908 8681
rect 21484 8632 21868 8672
rect 21292 8623 21332 8632
rect 21868 8623 21908 8632
rect 22444 8672 22484 9724
rect 22444 8623 22484 8632
rect 22636 9512 22676 9521
rect 22636 8672 22676 9472
rect 22636 8623 22676 8632
rect 22924 9092 22964 9101
rect 22924 8672 22964 9052
rect 23116 8924 23156 9808
rect 23116 8875 23156 8884
rect 23212 9596 23252 9605
rect 22924 8623 22964 8632
rect 23212 8504 23252 9556
rect 23500 9008 23540 10480
rect 25228 10436 25268 12100
rect 25228 10387 25268 10396
rect 26380 10856 26420 10865
rect 25900 10352 25940 10361
rect 25036 10268 25076 10277
rect 24556 10016 24596 10025
rect 23500 8959 23540 8968
rect 23596 9176 23636 9185
rect 23596 8672 23636 9136
rect 24556 8840 24596 9976
rect 25036 8924 25076 10228
rect 25900 9344 25940 10312
rect 25900 9295 25940 9304
rect 25036 8875 25076 8884
rect 26092 9176 26132 9185
rect 24556 8791 24596 8800
rect 23596 8623 23636 8632
rect 26092 8672 26132 9136
rect 26092 8623 26132 8632
rect 23212 8455 23252 8464
rect 26284 8420 26324 8429
rect 15820 8336 15860 8345
rect 15628 8252 15668 8261
rect 15244 8168 15284 8177
rect 14860 8000 14900 8009
rect 14380 391 14420 400
rect 14476 6740 14516 6749
rect 14476 80 14516 6700
rect 14668 6572 14708 6581
rect 14668 80 14708 6532
rect 14860 80 14900 7960
rect 15052 7916 15092 7925
rect 15052 80 15092 7876
rect 15148 4724 15188 4733
rect 15148 2624 15188 4684
rect 15148 2575 15188 2584
rect 15244 80 15284 8128
rect 15436 7244 15476 7253
rect 15436 80 15476 7204
rect 15628 80 15668 8212
rect 15820 80 15860 8296
rect 18604 8336 18644 8345
rect 17740 8252 17780 8261
rect 16588 8084 16628 8093
rect 16780 8084 16820 8093
rect 16628 8044 16780 8084
rect 16588 8035 16628 8044
rect 16780 8035 16820 8044
rect 17356 8000 17396 8009
rect 16012 7832 16052 7841
rect 15916 5900 15956 5909
rect 15916 5648 15956 5860
rect 15916 5599 15956 5608
rect 15916 4976 15956 4985
rect 15916 2120 15956 4936
rect 15916 2071 15956 2080
rect 16012 80 16052 7792
rect 17068 7748 17108 7757
rect 17068 7328 17108 7708
rect 17068 7279 17108 7288
rect 17356 7244 17396 7960
rect 17740 8000 17780 8212
rect 17740 7951 17780 7960
rect 18604 8000 18644 8296
rect 18808 8336 19176 8345
rect 18848 8296 18890 8336
rect 18930 8296 18972 8336
rect 19012 8296 19054 8336
rect 19094 8296 19136 8336
rect 18808 8287 19176 8296
rect 18604 7951 18644 7960
rect 25900 8252 25940 8261
rect 17452 7748 17492 7757
rect 17452 7412 17492 7708
rect 17836 7748 17876 7757
rect 17836 7496 17876 7708
rect 25420 7664 25460 7673
rect 20048 7580 20416 7589
rect 20088 7540 20130 7580
rect 20170 7540 20212 7580
rect 20252 7540 20294 7580
rect 20334 7540 20376 7580
rect 20048 7531 20416 7540
rect 17836 7447 17876 7456
rect 17452 7363 17492 7372
rect 17356 7195 17396 7204
rect 25228 7328 25268 7337
rect 17068 7160 17108 7169
rect 16300 7076 16340 7085
rect 16108 6992 16148 7001
rect 16108 2900 16148 6952
rect 16204 5816 16244 5825
rect 16204 4724 16244 5776
rect 16204 4675 16244 4684
rect 16108 2860 16244 2900
rect 16204 2204 16244 2860
rect 16204 2155 16244 2164
rect 16300 440 16340 7036
rect 16204 400 16340 440
rect 16396 6824 16436 6833
rect 16204 80 16244 400
rect 16396 80 16436 6784
rect 17068 6740 17108 7120
rect 17740 7160 17780 7169
rect 17068 6691 17108 6700
rect 17452 6992 17492 7001
rect 16588 6656 16628 6665
rect 16588 80 16628 6616
rect 16780 6488 16820 6497
rect 16780 80 16820 6448
rect 16972 6404 17012 6413
rect 16972 80 17012 6364
rect 17452 6152 17492 6952
rect 17740 6572 17780 7120
rect 18700 7160 18740 7169
rect 18220 7076 18260 7085
rect 17836 6992 17876 7001
rect 17836 6740 17876 6952
rect 18124 6992 18164 7001
rect 18124 6857 18164 6952
rect 18220 6824 18260 7036
rect 18220 6775 18260 6784
rect 18604 6992 18644 7001
rect 17836 6691 17876 6700
rect 17740 6523 17780 6532
rect 18412 6320 18452 6329
rect 17548 6236 17588 6245
rect 17740 6236 17780 6245
rect 17588 6196 17684 6236
rect 17548 6187 17588 6196
rect 17452 6103 17492 6112
rect 17164 6068 17204 6077
rect 17164 80 17204 6028
rect 17548 5900 17588 5909
rect 17356 5816 17396 5825
rect 17356 80 17396 5776
rect 17548 80 17588 5860
rect 17644 3464 17684 6196
rect 17644 3415 17684 3424
rect 17740 80 17780 6196
rect 18412 6185 18452 6280
rect 18604 6320 18644 6952
rect 18700 6656 18740 7120
rect 19276 7160 19316 7169
rect 18808 6824 19176 6833
rect 18848 6784 18890 6824
rect 18930 6784 18972 6824
rect 19012 6784 19054 6824
rect 19094 6784 19136 6824
rect 18808 6775 19176 6784
rect 18700 6607 18740 6616
rect 19276 6488 19316 7120
rect 19660 7160 19700 7169
rect 19372 6992 19412 7001
rect 19372 6656 19412 6952
rect 19372 6607 19412 6616
rect 19276 6439 19316 6448
rect 19660 6404 19700 7120
rect 19660 6355 19700 6364
rect 19852 7160 19892 7169
rect 18604 6271 18644 6280
rect 19852 6068 19892 7120
rect 20236 7160 20276 7169
rect 19852 6019 19892 6028
rect 19948 6992 19988 7001
rect 18700 5984 18740 5993
rect 18700 5144 18740 5944
rect 19948 5984 19988 6952
rect 20044 6572 20084 6581
rect 20044 6437 20084 6532
rect 20236 6236 20276 7120
rect 20716 7160 20756 7169
rect 20332 6532 20660 6572
rect 20332 6488 20372 6532
rect 20332 6439 20372 6448
rect 20236 6187 20276 6196
rect 20524 6320 20564 6329
rect 20048 6068 20416 6077
rect 20088 6028 20130 6068
rect 20170 6028 20212 6068
rect 20252 6028 20294 6068
rect 20334 6028 20376 6068
rect 20048 6019 20416 6028
rect 20524 6068 20564 6280
rect 20524 6019 20564 6028
rect 19948 5935 19988 5944
rect 20332 5648 20372 5657
rect 20332 5513 20372 5608
rect 20524 5648 20564 5657
rect 19948 5396 19988 5405
rect 18808 5312 19176 5321
rect 18848 5272 18890 5312
rect 18930 5272 18972 5312
rect 19012 5272 19054 5312
rect 19094 5272 19136 5312
rect 18808 5263 19176 5272
rect 18700 5104 18836 5144
rect 18124 4892 18164 4901
rect 17932 4640 17972 4649
rect 17932 80 17972 4600
rect 18124 80 18164 4852
rect 18700 4892 18740 4901
rect 18220 4556 18260 4565
rect 18220 1952 18260 4516
rect 18700 4556 18740 4852
rect 18700 4507 18740 4516
rect 18220 1903 18260 1912
rect 18316 4388 18356 4397
rect 18796 4388 18836 5104
rect 19852 4976 19892 4985
rect 19660 4892 19700 4901
rect 18316 80 18356 4348
rect 18700 4348 18836 4388
rect 19468 4640 19508 4649
rect 18700 3632 18740 4348
rect 19372 4136 19412 4145
rect 19276 3968 19316 3977
rect 18808 3800 19176 3809
rect 18848 3760 18890 3800
rect 18930 3760 18972 3800
rect 19012 3760 19054 3800
rect 19094 3760 19136 3800
rect 18808 3751 19176 3760
rect 19276 3800 19316 3928
rect 19276 3751 19316 3760
rect 19276 3632 19316 3641
rect 18700 3592 19220 3632
rect 18796 3464 18836 3473
rect 18700 3380 18740 3389
rect 18508 3128 18548 3137
rect 18508 2876 18548 3088
rect 18508 2827 18548 2836
rect 18700 2540 18740 3340
rect 18796 2624 18836 3424
rect 18796 2575 18836 2584
rect 18988 3212 19028 3221
rect 18604 2500 18740 2540
rect 18604 2036 18644 2500
rect 18988 2456 19028 3172
rect 18604 1987 18644 1996
rect 18700 2416 19028 2456
rect 19084 2624 19124 2633
rect 19084 2456 19124 2584
rect 19180 2540 19220 3592
rect 19180 2491 19220 2500
rect 18508 1616 18548 1625
rect 18508 80 18548 1576
rect 18700 80 18740 2416
rect 19084 2407 19124 2416
rect 18808 2288 19176 2297
rect 18848 2248 18890 2288
rect 18930 2248 18972 2288
rect 19012 2248 19054 2288
rect 19094 2248 19136 2288
rect 18808 2239 19176 2248
rect 19084 1532 19124 1541
rect 18892 1364 18932 1373
rect 18892 80 18932 1324
rect 19084 80 19124 1492
rect 19276 80 19316 3592
rect 19372 1532 19412 4096
rect 19372 1483 19412 1492
rect 19468 80 19508 4600
rect 19564 4472 19604 4481
rect 19564 3632 19604 4432
rect 19564 3583 19604 3592
rect 19564 3296 19604 3305
rect 19564 1364 19604 3256
rect 19564 1315 19604 1324
rect 19660 80 19700 4852
rect 19756 4556 19796 4565
rect 19756 2372 19796 4516
rect 19756 2323 19796 2332
rect 19852 80 19892 4936
rect 19948 1364 19988 5356
rect 20048 4556 20416 4565
rect 20088 4516 20130 4556
rect 20170 4516 20212 4556
rect 20252 4516 20294 4556
rect 20334 4516 20376 4556
rect 20048 4507 20416 4516
rect 20140 3548 20180 3557
rect 20140 3413 20180 3508
rect 20048 3044 20416 3053
rect 20088 3004 20130 3044
rect 20170 3004 20212 3044
rect 20252 3004 20294 3044
rect 20334 3004 20376 3044
rect 20048 2995 20416 3004
rect 20044 2540 20084 2549
rect 20044 1700 20084 2500
rect 20044 1651 20084 1660
rect 20048 1532 20416 1541
rect 20088 1492 20130 1532
rect 20170 1492 20212 1532
rect 20252 1492 20294 1532
rect 20334 1492 20376 1532
rect 20048 1483 20416 1492
rect 20236 1364 20276 1373
rect 20524 1364 20564 5608
rect 19948 1324 20084 1364
rect 20044 80 20084 1324
rect 20236 80 20276 1324
rect 20428 1324 20564 1364
rect 20428 80 20468 1324
rect 20620 80 20660 6532
rect 20716 5900 20756 7120
rect 21196 7160 21236 7169
rect 20812 6908 20852 6917
rect 20852 6868 21044 6908
rect 20812 6859 20852 6868
rect 20908 6572 20948 6581
rect 20908 6488 20948 6532
rect 20908 6437 20948 6448
rect 20716 5851 20756 5860
rect 20812 6404 20852 6413
rect 20716 5564 20756 5573
rect 20716 1364 20756 5524
rect 20716 1315 20756 1324
rect 20812 80 20852 6364
rect 21004 6320 21044 6868
rect 21004 6271 21044 6280
rect 21196 5816 21236 7120
rect 23980 7160 24020 7169
rect 23212 7076 23252 7085
rect 21196 5767 21236 5776
rect 21580 6992 21620 7001
rect 21580 5816 21620 6952
rect 22540 6488 22580 6497
rect 21580 5767 21620 5776
rect 21964 6068 22004 6077
rect 21580 5648 21620 5657
rect 21484 5564 21524 5573
rect 21292 5524 21484 5564
rect 20908 5480 20948 5489
rect 20908 2540 20948 5440
rect 21292 5396 21332 5524
rect 21484 5515 21524 5524
rect 21292 5347 21332 5356
rect 20908 2491 20948 2500
rect 21388 5228 21428 5237
rect 21196 2456 21236 2465
rect 21196 80 21236 2416
rect 21388 2036 21428 5188
rect 21580 4556 21620 5608
rect 21580 4507 21620 4516
rect 21676 4724 21716 4733
rect 21388 1987 21428 1996
rect 21580 2456 21620 2465
rect 21388 1700 21428 1709
rect 21388 80 21428 1660
rect 21580 80 21620 2416
rect 21676 1952 21716 4684
rect 21964 2708 22004 6028
rect 22252 5396 22292 5405
rect 22252 4976 22292 5356
rect 22252 4927 22292 4936
rect 21964 2659 22004 2668
rect 21676 1903 21716 1912
rect 21964 2456 22004 2465
rect 21772 1700 21812 1709
rect 21772 80 21812 1660
rect 21964 80 22004 2416
rect 22348 2456 22388 2465
rect 22156 1700 22196 1709
rect 22156 80 22196 1660
rect 22348 80 22388 2416
rect 22540 2036 22580 6448
rect 22732 5816 22772 5825
rect 22636 4556 22676 4565
rect 22636 2624 22676 4516
rect 22732 3044 22772 5776
rect 23116 5480 23156 5489
rect 23116 5228 23156 5440
rect 23020 5188 23156 5228
rect 22828 4976 22868 4985
rect 22828 4388 22868 4936
rect 22924 4976 22964 4985
rect 22924 4640 22964 4936
rect 23020 4724 23060 5188
rect 23116 5060 23156 5069
rect 23116 4976 23156 5020
rect 23116 4925 23156 4936
rect 23020 4675 23060 4684
rect 22924 4591 22964 4600
rect 22828 4339 22868 4348
rect 23116 4220 23156 4229
rect 23116 3548 23156 4180
rect 23116 3499 23156 3508
rect 22732 3004 22964 3044
rect 22924 2900 22964 3004
rect 23212 2900 23252 7036
rect 23788 6740 23828 6749
rect 23308 6572 23348 6581
rect 23308 4304 23348 6532
rect 23596 6152 23636 6161
rect 23404 4976 23444 4985
rect 23404 4472 23444 4936
rect 23404 4423 23444 4432
rect 23308 4264 23444 4304
rect 22636 2575 22676 2584
rect 22828 2876 22868 2885
rect 22924 2876 23060 2900
rect 22924 2860 23020 2876
rect 22540 1987 22580 1996
rect 22732 2456 22772 2465
rect 22540 1700 22580 1709
rect 22540 80 22580 1660
rect 22732 80 22772 2416
rect 22828 1952 22868 2836
rect 23212 2860 23348 2900
rect 23020 2827 23060 2836
rect 22828 1903 22868 1912
rect 23116 2456 23156 2465
rect 22924 1700 22964 1709
rect 22924 80 22964 1660
rect 23116 80 23156 2416
rect 23308 2372 23348 2860
rect 23308 2323 23348 2332
rect 23404 2036 23444 4264
rect 23404 1987 23444 1996
rect 23500 2456 23540 2465
rect 23308 1700 23348 1709
rect 23308 80 23348 1660
rect 23500 80 23540 2416
rect 23596 1952 23636 6112
rect 23596 1903 23636 1912
rect 23788 1952 23828 6700
rect 23980 2624 24020 7120
rect 24268 6992 24308 7001
rect 24172 6908 24212 6917
rect 23980 2575 24020 2584
rect 24076 6236 24116 6245
rect 24076 2624 24116 6196
rect 24172 3128 24212 6868
rect 24172 3079 24212 3088
rect 24268 2900 24308 6952
rect 24844 6404 24884 6413
rect 24460 4136 24500 4145
rect 24460 3296 24500 4096
rect 24748 3800 24788 3809
rect 24748 3464 24788 3760
rect 24748 3415 24788 3424
rect 24460 3247 24500 3256
rect 24460 3128 24500 3137
rect 24268 2860 24404 2900
rect 24076 2575 24116 2584
rect 23788 1903 23828 1912
rect 24172 1784 24212 1793
rect 24076 1744 24172 1784
rect 23692 1700 23732 1709
rect 23692 80 23732 1660
rect 23884 1700 23924 1709
rect 23884 80 23924 1660
rect 24076 80 24116 1744
rect 24172 1735 24212 1744
rect 24268 1700 24308 1709
rect 24268 80 24308 1660
rect 24364 1532 24404 2860
rect 24460 2708 24500 3088
rect 24460 2659 24500 2668
rect 24556 2288 24596 2297
rect 24596 2248 24692 2288
rect 24556 2239 24596 2248
rect 24652 2036 24692 2248
rect 24652 1987 24692 1996
rect 24844 1952 24884 6364
rect 25132 5984 25172 5993
rect 24940 4052 24980 4061
rect 24940 3044 24980 4012
rect 24940 2995 24980 3004
rect 25132 2876 25172 5944
rect 25132 2827 25172 2836
rect 25228 2708 25268 7288
rect 25324 4136 25364 4145
rect 25324 3212 25364 4096
rect 25324 3163 25364 3172
rect 25420 2900 25460 7624
rect 25132 2668 25268 2708
rect 25324 2860 25460 2900
rect 25516 7412 25556 7421
rect 25516 2876 25556 7372
rect 25900 7412 25940 8212
rect 26284 8000 26324 8380
rect 26284 7951 26324 7960
rect 25900 7363 25940 7372
rect 25804 6824 25844 6833
rect 24844 1903 24884 1912
rect 24940 2540 24980 2549
rect 24940 1952 24980 2500
rect 25132 2372 25172 2668
rect 25324 2540 25364 2860
rect 25516 2827 25556 2836
rect 25612 6656 25652 6665
rect 25324 2491 25364 2500
rect 25420 2792 25460 2801
rect 25132 2323 25172 2332
rect 25228 2456 25268 2465
rect 24940 1903 24980 1912
rect 24652 1784 24692 1793
rect 24364 1483 24404 1492
rect 24460 1700 24500 1709
rect 24460 80 24500 1660
rect 24652 80 24692 1744
rect 24844 1700 24884 1709
rect 24844 80 24884 1660
rect 25036 1616 25076 1625
rect 25036 80 25076 1576
rect 25228 80 25268 2416
rect 25420 2036 25460 2752
rect 25612 2624 25652 6616
rect 25708 6320 25748 6329
rect 25708 2792 25748 6280
rect 25708 2743 25748 2752
rect 25804 2708 25844 6784
rect 25996 4136 26036 4145
rect 25900 4052 25940 4061
rect 25900 2876 25940 4012
rect 25996 4001 26036 4096
rect 26188 3968 26228 3977
rect 25996 3464 26036 3473
rect 25996 3329 26036 3424
rect 26188 3128 26228 3928
rect 26380 3212 26420 10816
rect 26764 10604 26804 10613
rect 26380 3163 26420 3172
rect 26668 7580 26708 7589
rect 26188 3079 26228 3088
rect 25900 2827 25940 2836
rect 26092 3044 26132 3053
rect 25804 2659 25844 2668
rect 25612 2584 25748 2624
rect 25420 1987 25460 1996
rect 25612 2456 25652 2465
rect 25420 1784 25460 1793
rect 25420 80 25460 1744
rect 25612 80 25652 2416
rect 25708 2204 25748 2584
rect 25708 2155 25748 2164
rect 25996 2456 26036 2465
rect 25804 1616 25844 1625
rect 25804 80 25844 1576
rect 25996 80 26036 2416
rect 26092 2204 26132 3004
rect 26092 2155 26132 2164
rect 26380 2456 26420 2465
rect 26188 2036 26228 2045
rect 26188 80 26228 1996
rect 26380 80 26420 2416
rect 26668 2120 26708 7540
rect 26764 3632 26804 10564
rect 27340 10436 27380 12100
rect 27340 10387 27380 10396
rect 29452 10436 29492 12100
rect 31180 10772 31220 10781
rect 29452 10387 29492 10396
rect 30220 10520 30260 10529
rect 30220 10385 30260 10480
rect 28396 10352 28436 10361
rect 27244 10184 27284 10193
rect 26860 10100 26900 10109
rect 26860 8924 26900 10060
rect 26860 8875 26900 8884
rect 27148 9764 27188 9773
rect 27148 8672 27188 9724
rect 27244 8924 27284 10144
rect 27244 8875 27284 8884
rect 27628 10184 27668 10193
rect 27628 8924 27668 10144
rect 28108 10100 28148 10109
rect 27628 8875 27668 8884
rect 27724 9932 27764 9941
rect 27148 8623 27188 8632
rect 27724 8672 27764 9892
rect 27916 9932 27956 9941
rect 27916 9428 27956 9892
rect 27916 9379 27956 9388
rect 28012 9260 28052 9269
rect 28012 8840 28052 9220
rect 28012 8791 28052 8800
rect 27724 8623 27764 8632
rect 28108 8168 28148 10060
rect 28300 9428 28340 9437
rect 28300 8672 28340 9388
rect 28300 8623 28340 8632
rect 28108 8119 28148 8128
rect 27916 7916 27956 7925
rect 27724 7876 27916 7916
rect 27724 7832 27764 7876
rect 27916 7867 27956 7876
rect 27724 7783 27764 7792
rect 26764 3583 26804 3592
rect 26860 7496 26900 7505
rect 26764 3464 26804 3473
rect 26764 3044 26804 3424
rect 26764 2995 26804 3004
rect 26668 2071 26708 2080
rect 26764 2456 26804 2465
rect 26476 1952 26516 1961
rect 26476 1532 26516 1912
rect 26476 1483 26516 1492
rect 26572 1616 26612 1625
rect 26572 80 26612 1576
rect 26764 80 26804 2416
rect 26860 1868 26900 7456
rect 27244 7412 27284 7421
rect 26956 5060 26996 5069
rect 26956 4892 26996 5020
rect 26956 4843 26996 4852
rect 26956 4724 26996 4733
rect 26956 4388 26996 4684
rect 26956 4339 26996 4348
rect 27052 4220 27092 4229
rect 27052 3464 27092 4180
rect 27052 3415 27092 3424
rect 27244 2900 27284 7372
rect 27340 7160 27380 7169
rect 27340 3128 27380 7120
rect 27820 4892 27860 4901
rect 27820 4640 27860 4852
rect 27820 4591 27860 4600
rect 28012 4472 28052 4481
rect 27436 4052 27476 4061
rect 27436 3464 27476 4012
rect 27532 3884 27572 3893
rect 27532 3632 27572 3844
rect 27628 3800 27668 3809
rect 27628 3665 27668 3760
rect 27532 3583 27572 3592
rect 27436 3415 27476 3424
rect 27820 3464 27860 3473
rect 27340 3079 27380 3088
rect 27820 3128 27860 3424
rect 27916 3464 27956 3473
rect 27916 3296 27956 3424
rect 27916 3247 27956 3256
rect 27820 3079 27860 3088
rect 27148 2860 27284 2900
rect 27916 2876 27956 2885
rect 27148 2708 27188 2860
rect 27916 2792 27956 2836
rect 27916 2741 27956 2752
rect 27148 2659 27188 2668
rect 28012 2708 28052 4432
rect 28204 4472 28244 4481
rect 28204 3632 28244 4432
rect 28204 3583 28244 3592
rect 28204 3464 28244 3473
rect 28204 2960 28244 3424
rect 28396 3212 28436 10312
rect 28876 10268 28916 10277
rect 28780 10184 28820 10193
rect 28780 8924 28820 10144
rect 28780 8875 28820 8884
rect 28780 8252 28820 8261
rect 28588 6404 28628 6413
rect 28396 3163 28436 3172
rect 28492 4220 28532 4229
rect 28204 2911 28244 2920
rect 28012 2659 28052 2668
rect 28396 2624 28436 2633
rect 28396 2489 28436 2584
rect 27148 2456 27188 2465
rect 27052 2204 27092 2213
rect 27052 1952 27092 2164
rect 27052 1903 27092 1912
rect 26860 1819 26900 1828
rect 26956 1784 26996 1793
rect 26956 80 26996 1744
rect 27148 80 27188 2416
rect 27532 2456 27572 2465
rect 27340 2204 27380 2213
rect 27340 2069 27380 2164
rect 27436 1952 27476 1961
rect 27436 1817 27476 1912
rect 27340 1616 27380 1625
rect 27340 80 27380 1576
rect 27532 80 27572 2416
rect 27916 2456 27956 2465
rect 27724 1616 27764 1625
rect 27724 80 27764 1576
rect 27916 80 27956 2416
rect 28300 2456 28340 2465
rect 28108 2036 28148 2131
rect 28108 1987 28148 1996
rect 28108 1784 28148 1793
rect 28108 80 28148 1744
rect 28300 80 28340 2416
rect 28492 1868 28532 4180
rect 28588 3464 28628 6364
rect 28588 3415 28628 3424
rect 28492 1819 28532 1828
rect 28684 2456 28724 2465
rect 28492 1616 28532 1625
rect 28492 80 28532 1576
rect 28684 80 28724 2416
rect 28780 1952 28820 8212
rect 28876 8168 28916 10228
rect 30796 9848 30836 9857
rect 30220 9680 30260 9689
rect 30220 9545 30260 9640
rect 30604 9512 30644 9521
rect 29068 9344 29108 9353
rect 29068 8924 29108 9304
rect 29068 8875 29108 8884
rect 30604 8924 30644 9472
rect 30796 9344 30836 9808
rect 30796 9295 30836 9304
rect 30892 9512 30932 9521
rect 30604 8875 30644 8884
rect 30892 8840 30932 9472
rect 30892 8791 30932 8800
rect 31180 8840 31220 10732
rect 31180 8791 31220 8800
rect 31468 10688 31508 10697
rect 31468 8588 31508 10648
rect 31564 10436 31604 12100
rect 31564 10387 31604 10396
rect 33676 10436 33716 12100
rect 35168 10604 35536 10613
rect 35208 10564 35250 10604
rect 35290 10564 35332 10604
rect 35372 10564 35414 10604
rect 35454 10564 35496 10604
rect 35168 10555 35536 10564
rect 33676 10387 33716 10396
rect 35788 10436 35828 12100
rect 35788 10387 35828 10396
rect 37900 10436 37940 12100
rect 37900 10387 37940 10396
rect 40012 10436 40052 12100
rect 40012 10387 40052 10396
rect 40204 10688 40244 10697
rect 34540 10184 34580 10193
rect 31468 8539 31508 8548
rect 32140 9932 32180 9941
rect 28876 8119 28916 8128
rect 30988 8084 31028 8093
rect 30988 7832 31028 8044
rect 30988 7783 31028 7792
rect 29932 5648 29972 5657
rect 28972 5564 29012 5573
rect 28876 5480 28916 5489
rect 28876 2120 28916 5440
rect 28972 2624 29012 5524
rect 29356 5396 29396 5405
rect 28972 2575 29012 2584
rect 29164 4136 29204 4145
rect 29164 2540 29204 4096
rect 29356 2624 29396 5356
rect 29356 2575 29396 2584
rect 29548 5312 29588 5321
rect 29164 2491 29204 2500
rect 28876 2071 28916 2080
rect 29068 2456 29108 2465
rect 28780 1903 28820 1912
rect 28876 1616 28916 1625
rect 28876 80 28916 1576
rect 29068 80 29108 2416
rect 29452 2456 29492 2465
rect 29260 2036 29300 2045
rect 29260 80 29300 1996
rect 29452 80 29492 2416
rect 29548 1952 29588 5272
rect 29548 1903 29588 1912
rect 29836 2456 29876 2465
rect 29644 1616 29684 1625
rect 29644 80 29684 1576
rect 29836 80 29876 2416
rect 29932 1952 29972 5608
rect 31660 5060 31700 5069
rect 31276 4724 31316 4733
rect 30796 4640 30836 4649
rect 30836 4600 30932 4640
rect 30796 4591 30836 4600
rect 30220 4556 30260 4565
rect 30124 3548 30164 3557
rect 30124 3413 30164 3508
rect 30220 2708 30260 4516
rect 30220 2659 30260 2668
rect 30700 4388 30740 4397
rect 29932 1903 29972 1912
rect 30220 2456 30260 2465
rect 30028 1784 30068 1793
rect 30028 80 30068 1744
rect 30220 80 30260 2416
rect 30604 2456 30644 2465
rect 30412 1616 30452 1625
rect 30412 80 30452 1576
rect 30604 80 30644 2416
rect 30700 1952 30740 4348
rect 30892 4388 30932 4600
rect 30892 4339 30932 4348
rect 30892 4052 30932 4061
rect 30892 3464 30932 4012
rect 30892 3415 30932 3424
rect 31276 2624 31316 4684
rect 31276 2575 31316 2584
rect 30700 1903 30740 1912
rect 30988 2456 31028 2465
rect 30796 1616 30836 1625
rect 30796 80 30836 1576
rect 30988 80 31028 2416
rect 31660 1952 31700 5020
rect 31660 1903 31700 1912
rect 31948 440 31988 449
rect 31756 356 31796 365
rect 31372 272 31412 281
rect 31180 104 31220 113
rect 8812 55 8852 64
rect 11000 0 11080 80
rect 11192 0 11272 80
rect 11384 0 11464 80
rect 11576 0 11656 80
rect 11768 0 11848 80
rect 11960 0 12040 80
rect 12152 0 12232 80
rect 12344 0 12424 80
rect 12536 0 12616 80
rect 12728 0 12808 80
rect 12920 0 13000 80
rect 13112 0 13192 80
rect 13304 0 13384 80
rect 13496 0 13576 80
rect 13688 0 13768 80
rect 13880 0 13960 80
rect 14072 0 14152 80
rect 14264 0 14344 80
rect 14456 0 14536 80
rect 14648 0 14728 80
rect 14840 0 14920 80
rect 15032 0 15112 80
rect 15224 0 15304 80
rect 15416 0 15496 80
rect 15608 0 15688 80
rect 15800 0 15880 80
rect 15992 0 16072 80
rect 16184 0 16264 80
rect 16376 0 16456 80
rect 16568 0 16648 80
rect 16760 0 16840 80
rect 16952 0 17032 80
rect 17144 0 17224 80
rect 17336 0 17416 80
rect 17528 0 17608 80
rect 17720 0 17800 80
rect 17912 0 17992 80
rect 18104 0 18184 80
rect 18296 0 18376 80
rect 18488 0 18568 80
rect 18680 0 18760 80
rect 18872 0 18952 80
rect 19064 0 19144 80
rect 19256 0 19336 80
rect 19448 0 19528 80
rect 19640 0 19720 80
rect 19832 0 19912 80
rect 20024 0 20104 80
rect 20216 0 20296 80
rect 20408 0 20488 80
rect 20600 0 20680 80
rect 20792 0 20872 80
rect 20984 0 21064 80
rect 21176 0 21256 80
rect 21368 0 21448 80
rect 21560 0 21640 80
rect 21752 0 21832 80
rect 21944 0 22024 80
rect 22136 0 22216 80
rect 22328 0 22408 80
rect 22520 0 22600 80
rect 22712 0 22792 80
rect 22904 0 22984 80
rect 23096 0 23176 80
rect 23288 0 23368 80
rect 23480 0 23560 80
rect 23672 0 23752 80
rect 23864 0 23944 80
rect 24056 0 24136 80
rect 24248 0 24328 80
rect 24440 0 24520 80
rect 24632 0 24712 80
rect 24824 0 24904 80
rect 25016 0 25096 80
rect 25208 0 25288 80
rect 25400 0 25480 80
rect 25592 0 25672 80
rect 25784 0 25864 80
rect 25976 0 26056 80
rect 26168 0 26248 80
rect 26360 0 26440 80
rect 26552 0 26632 80
rect 26744 0 26824 80
rect 26936 0 27016 80
rect 27128 0 27208 80
rect 27320 0 27400 80
rect 27512 0 27592 80
rect 27704 0 27784 80
rect 27896 0 27976 80
rect 28088 0 28168 80
rect 28280 0 28360 80
rect 28472 0 28552 80
rect 28664 0 28744 80
rect 28856 0 28936 80
rect 29048 0 29128 80
rect 29240 0 29320 80
rect 29432 0 29512 80
rect 29624 0 29704 80
rect 29816 0 29896 80
rect 30008 0 30088 80
rect 30200 0 30280 80
rect 30392 0 30472 80
rect 30584 0 30664 80
rect 30776 0 30856 80
rect 30968 0 31048 80
rect 31160 64 31180 80
rect 31372 80 31412 232
rect 31564 188 31604 197
rect 31564 80 31604 148
rect 31756 80 31796 316
rect 31948 80 31988 400
rect 32140 80 32180 9892
rect 33928 9848 34296 9857
rect 33968 9808 34010 9848
rect 34050 9808 34092 9848
rect 34132 9808 34174 9848
rect 34214 9808 34256 9848
rect 33928 9799 34296 9808
rect 33100 9764 33140 9773
rect 33100 9596 33140 9724
rect 33100 9547 33140 9556
rect 33292 9596 33332 9605
rect 32332 9176 32372 9185
rect 32332 80 32372 9136
rect 32716 8672 32756 8681
rect 32524 8588 32564 8597
rect 32524 80 32564 8548
rect 32716 80 32756 8632
rect 32908 8504 32948 8513
rect 32908 80 32948 8464
rect 33196 6488 33236 6497
rect 33196 6353 33236 6448
rect 33292 3044 33332 9556
rect 33484 9512 33524 9521
rect 33196 3004 33332 3044
rect 33388 8672 33428 8681
rect 33196 2900 33236 3004
rect 33004 2860 33236 2900
rect 33292 2900 33332 2909
rect 33004 440 33044 2860
rect 33004 400 33140 440
rect 33100 80 33140 400
rect 33292 80 33332 2860
rect 33388 1952 33428 8632
rect 33484 3044 33524 9472
rect 33772 9428 33812 9437
rect 33484 2995 33524 3004
rect 33580 8000 33620 8009
rect 33388 1903 33428 1912
rect 33484 2900 33524 2909
rect 33484 80 33524 2860
rect 33580 2120 33620 7960
rect 33676 7748 33716 7757
rect 33676 2120 33716 7708
rect 33772 3044 33812 9388
rect 33928 8336 34296 8345
rect 33968 8296 34010 8336
rect 34050 8296 34092 8336
rect 34132 8296 34174 8336
rect 34214 8296 34256 8336
rect 33928 8287 34296 8296
rect 33928 6824 34296 6833
rect 33968 6784 34010 6824
rect 34050 6784 34092 6824
rect 34132 6784 34174 6824
rect 34214 6784 34256 6824
rect 33928 6775 34296 6784
rect 34540 6656 34580 10144
rect 40204 10184 40244 10648
rect 40300 10520 40340 10615
rect 40300 10471 40340 10480
rect 42124 10436 42164 12100
rect 44044 11192 44084 11201
rect 42124 10387 42164 10396
rect 42412 10856 42452 10865
rect 40204 10135 40244 10144
rect 40396 10184 40436 10195
rect 35596 10100 35636 10109
rect 35168 9092 35536 9101
rect 35208 9052 35250 9092
rect 35290 9052 35332 9092
rect 35372 9052 35414 9092
rect 35454 9052 35496 9092
rect 35168 9043 35536 9052
rect 35168 7580 35536 7589
rect 35208 7540 35250 7580
rect 35290 7540 35332 7580
rect 35372 7540 35414 7580
rect 35454 7540 35496 7580
rect 35168 7531 35536 7540
rect 34540 6607 34580 6616
rect 34444 6320 34484 6329
rect 34348 5648 34388 5657
rect 33928 5312 34296 5321
rect 33968 5272 34010 5312
rect 34050 5272 34092 5312
rect 34132 5272 34174 5312
rect 34214 5272 34256 5312
rect 33928 5263 34296 5272
rect 34348 4976 34388 5608
rect 34348 4927 34388 4936
rect 34444 4724 34484 6280
rect 35168 6068 35536 6077
rect 35208 6028 35250 6068
rect 35290 6028 35332 6068
rect 35372 6028 35414 6068
rect 35454 6028 35496 6068
rect 35168 6019 35536 6028
rect 34348 4684 34484 4724
rect 33928 3800 34296 3809
rect 33968 3760 34010 3800
rect 34050 3760 34092 3800
rect 34132 3760 34174 3800
rect 34214 3760 34256 3800
rect 33928 3751 34296 3760
rect 33772 2995 33812 3004
rect 33928 2288 34296 2297
rect 33968 2248 34010 2288
rect 34050 2248 34092 2288
rect 34132 2248 34174 2288
rect 34214 2248 34256 2288
rect 33928 2239 34296 2248
rect 34060 2120 34100 2129
rect 34348 2120 34388 4684
rect 35168 4556 35536 4565
rect 35208 4516 35250 4556
rect 35290 4516 35332 4556
rect 35372 4516 35414 4556
rect 35454 4516 35496 4556
rect 35168 4507 35536 4516
rect 34828 4388 34868 4397
rect 33676 2080 33908 2120
rect 33580 2071 33620 2080
rect 33676 1952 33716 1961
rect 33676 80 33716 1912
rect 33868 80 33908 2080
rect 34060 80 34100 2080
rect 34252 2080 34388 2120
rect 34444 3464 34484 3473
rect 34252 80 34292 2080
rect 34444 80 34484 3424
rect 34828 3464 34868 4348
rect 35596 4220 35636 10060
rect 40396 10100 40436 10144
rect 42412 10184 42452 10816
rect 42412 10135 42452 10144
rect 43180 10520 43220 10529
rect 43180 10184 43220 10480
rect 43180 10135 43220 10144
rect 43564 10184 43604 10193
rect 40396 10051 40436 10060
rect 38092 9596 38132 9605
rect 37996 9260 38036 9269
rect 37996 8756 38036 9220
rect 37996 8707 38036 8716
rect 38092 8672 38132 9556
rect 43564 9428 43604 10144
rect 43948 10184 43988 10193
rect 43564 9379 43604 9388
rect 43756 9512 43796 9521
rect 38188 9344 38228 9353
rect 38188 9008 38228 9304
rect 38188 8959 38228 8968
rect 38092 8623 38132 8632
rect 43756 7916 43796 9472
rect 43948 8924 43988 10144
rect 44044 9596 44084 11152
rect 44236 10436 44276 12100
rect 44236 10387 44276 10396
rect 44428 10520 44468 10529
rect 44428 9680 44468 10480
rect 44524 10184 44564 10279
rect 44524 10135 44564 10144
rect 44908 10184 44948 10193
rect 44428 9631 44468 9640
rect 44044 9547 44084 9556
rect 43948 8875 43988 8884
rect 44524 9008 44564 9017
rect 44524 8000 44564 8968
rect 44908 8084 44948 10144
rect 45772 10016 45812 10025
rect 45772 9512 45812 9976
rect 45772 9463 45812 9472
rect 45772 9260 45812 9269
rect 45772 8840 45812 9220
rect 45772 8791 45812 8800
rect 46252 8672 46292 8681
rect 46252 8168 46292 8632
rect 46252 8119 46292 8128
rect 44908 8035 44948 8044
rect 44524 7951 44564 7960
rect 43756 7867 43796 7876
rect 46252 7664 46292 7673
rect 46252 7496 46292 7624
rect 46252 7447 46292 7456
rect 43180 7076 43220 7085
rect 43084 7036 43180 7076
rect 41740 6236 41780 6245
rect 38572 5732 38612 5741
rect 36940 5648 36980 5657
rect 36940 5396 36980 5608
rect 36940 5347 36980 5356
rect 37612 5648 37652 5657
rect 37612 4724 37652 5608
rect 37420 4640 37460 4649
rect 35596 4171 35636 4180
rect 35980 4556 36020 4565
rect 34732 3212 34772 3221
rect 34636 3044 34676 3053
rect 34636 80 34676 3004
rect 34732 2120 34772 3172
rect 34828 2876 34868 3424
rect 35980 3464 36020 4516
rect 37324 4052 37364 4061
rect 37132 3884 37172 3893
rect 37324 3884 37364 4012
rect 37172 3844 37364 3884
rect 37132 3835 37172 3844
rect 37420 3716 37460 4600
rect 37420 3667 37460 3676
rect 35980 3415 36020 3424
rect 34828 2827 34868 2836
rect 35020 3128 35060 3137
rect 34732 2080 34868 2120
rect 34828 80 34868 2080
rect 35020 80 35060 3088
rect 35168 3044 35536 3053
rect 35208 3004 35250 3044
rect 35290 3004 35332 3044
rect 35372 3004 35414 3044
rect 35454 3004 35496 3044
rect 35168 2995 35536 3004
rect 35168 1532 35536 1541
rect 35208 1492 35250 1532
rect 35290 1492 35332 1532
rect 35372 1492 35414 1532
rect 35454 1492 35496 1532
rect 35168 1483 35536 1492
rect 37612 1448 37652 4684
rect 37900 5648 37940 5657
rect 37900 1784 37940 5608
rect 38092 5480 38132 5489
rect 38092 4892 38132 5440
rect 38572 5060 38612 5692
rect 41068 5564 41108 5573
rect 38572 5011 38612 5020
rect 40876 5524 41068 5564
rect 40876 5060 40916 5524
rect 41068 5515 41108 5524
rect 40876 5011 40916 5020
rect 41068 5144 41108 5153
rect 38092 4843 38132 4852
rect 39052 4892 39092 4901
rect 37996 4304 38036 4313
rect 37996 3464 38036 4264
rect 38092 4220 38132 4229
rect 38092 3884 38132 4180
rect 38092 3835 38132 3844
rect 37996 3415 38036 3424
rect 39052 1952 39092 4852
rect 39340 4724 39380 4733
rect 39340 4388 39380 4684
rect 39340 2792 39380 4348
rect 39340 2743 39380 2752
rect 40108 4724 40148 4733
rect 40108 2456 40148 4684
rect 40300 4724 40340 4733
rect 40300 4388 40340 4684
rect 40300 4339 40340 4348
rect 41068 3464 41108 5104
rect 41356 5144 41396 5153
rect 41260 4808 41300 4817
rect 41260 4220 41300 4768
rect 41356 4556 41396 5104
rect 41356 4507 41396 4516
rect 41260 4171 41300 4180
rect 41068 3415 41108 3424
rect 40108 2407 40148 2416
rect 41740 2036 41780 6196
rect 43084 5732 43124 7036
rect 43180 7008 43220 7036
rect 46252 6992 46292 7001
rect 46252 6824 46292 6952
rect 46252 6775 46292 6784
rect 43084 5683 43124 5692
rect 44620 6404 44660 6413
rect 43852 5648 43892 5657
rect 43852 4052 43892 5608
rect 44140 5480 44180 5489
rect 43852 4003 43892 4012
rect 44044 4892 44084 4901
rect 44044 3380 44084 4852
rect 44044 3331 44084 3340
rect 44140 2624 44180 5440
rect 44332 5396 44372 5405
rect 44236 5060 44276 5069
rect 44236 2708 44276 5020
rect 44332 2900 44372 5356
rect 44428 4808 44468 4817
rect 44428 3464 44468 4768
rect 44524 4136 44564 4145
rect 44524 3632 44564 4096
rect 44524 3583 44564 3592
rect 44428 3424 44564 3464
rect 44332 2860 44468 2900
rect 44236 2659 44276 2668
rect 44140 2575 44180 2584
rect 41740 1987 41780 1996
rect 39052 1903 39092 1912
rect 44428 1952 44468 2860
rect 44524 2624 44564 3424
rect 44620 3128 44660 6364
rect 44620 3079 44660 3088
rect 44716 5228 44756 5237
rect 44524 2575 44564 2584
rect 44428 1903 44468 1912
rect 44716 1952 44756 5188
rect 44908 4136 44948 4145
rect 44908 3296 44948 4096
rect 44908 3247 44948 3256
rect 44716 1903 44756 1912
rect 45676 2456 45716 2465
rect 37900 1735 37940 1744
rect 44620 1784 44660 1793
rect 37612 1399 37652 1408
rect 44620 1112 44660 1744
rect 44620 1063 44660 1072
rect 45388 1700 45428 1709
rect 45388 776 45428 1660
rect 45676 1448 45716 2416
rect 45676 1399 45716 1408
rect 45388 727 45428 736
rect 31220 64 31240 80
rect 31160 0 31240 64
rect 31352 0 31432 80
rect 31544 0 31624 80
rect 31736 0 31816 80
rect 31928 0 32008 80
rect 32120 0 32200 80
rect 32312 0 32392 80
rect 32504 0 32584 80
rect 32696 0 32776 80
rect 32888 0 32968 80
rect 33080 0 33160 80
rect 33272 0 33352 80
rect 33464 0 33544 80
rect 33656 0 33736 80
rect 33848 0 33928 80
rect 34040 0 34120 80
rect 34232 0 34312 80
rect 34424 0 34504 80
rect 34616 0 34696 80
rect 34808 0 34888 80
rect 35000 0 35080 80
<< via3 >>
rect 76 8800 116 8840
rect 4928 10564 4968 10604
rect 5010 10564 5050 10604
rect 5092 10564 5132 10604
rect 5174 10564 5214 10604
rect 5256 10564 5296 10604
rect 3688 9808 3728 9848
rect 3770 9808 3810 9848
rect 3852 9808 3892 9848
rect 3934 9808 3974 9848
rect 4016 9808 4056 9848
rect 4928 9052 4968 9092
rect 5010 9052 5050 9092
rect 5092 9052 5132 9092
rect 5174 9052 5214 9092
rect 5256 9052 5296 9092
rect 20048 10564 20088 10604
rect 20130 10564 20170 10604
rect 20212 10564 20252 10604
rect 20294 10564 20334 10604
rect 20376 10564 20416 10604
rect 18808 9808 18848 9848
rect 18890 9808 18930 9848
rect 18972 9808 19012 9848
rect 19054 9808 19094 9848
rect 19136 9808 19176 9848
rect 10060 8800 10100 8840
rect 3688 8296 3728 8336
rect 3770 8296 3810 8336
rect 3852 8296 3892 8336
rect 3934 8296 3974 8336
rect 4016 8296 4056 8336
rect 4928 7540 4968 7580
rect 5010 7540 5050 7580
rect 5092 7540 5132 7580
rect 5174 7540 5214 7580
rect 5256 7540 5296 7580
rect 460 6448 500 6488
rect 3688 6784 3728 6824
rect 3770 6784 3810 6824
rect 3852 6784 3892 6824
rect 3934 6784 3974 6824
rect 4016 6784 4056 6824
rect 4928 6028 4968 6068
rect 5010 6028 5050 6068
rect 5092 6028 5132 6068
rect 5174 6028 5214 6068
rect 5256 6028 5296 6068
rect 3688 5272 3728 5312
rect 3770 5272 3810 5312
rect 3852 5272 3892 5312
rect 3934 5272 3974 5312
rect 4016 5272 4056 5312
rect 3688 3760 3728 3800
rect 3770 3760 3810 3800
rect 3852 3760 3892 3800
rect 3934 3760 3974 3800
rect 4016 3760 4056 3800
rect 4928 4516 4968 4556
rect 5010 4516 5050 4556
rect 5092 4516 5132 4556
rect 5174 4516 5214 4556
rect 5256 4516 5296 4556
rect 4928 3004 4968 3044
rect 5010 3004 5050 3044
rect 5092 3004 5132 3044
rect 5174 3004 5214 3044
rect 5256 3004 5296 3044
rect 1420 2752 1460 2792
rect 1420 2416 1460 2456
rect 3688 2248 3728 2288
rect 3770 2248 3810 2288
rect 3852 2248 3892 2288
rect 3934 2248 3974 2288
rect 4016 2248 4056 2288
rect 1420 1744 1460 1784
rect 4928 1492 4968 1532
rect 5010 1492 5050 1532
rect 5092 1492 5132 1532
rect 5174 1492 5214 1532
rect 5256 1492 5296 1532
rect 1420 1408 1460 1448
rect 6700 4600 6740 4640
rect 7468 316 7508 356
rect 6892 232 6932 272
rect 6412 148 6452 188
rect 10540 5608 10580 5648
rect 10060 5356 10100 5396
rect 10060 4600 10100 4640
rect 10636 4012 10676 4052
rect 10060 3844 10100 3884
rect 10444 3844 10484 3884
rect 8812 64 8852 104
rect 11980 5608 12020 5648
rect 11692 4180 11732 4220
rect 11884 4096 11924 4136
rect 11692 4012 11732 4052
rect 11788 3928 11828 3968
rect 12652 5608 12692 5648
rect 12940 5608 12980 5648
rect 12076 3928 12116 3968
rect 20048 9052 20088 9092
rect 20130 9052 20170 9092
rect 20212 9052 20252 9092
rect 20294 9052 20334 9092
rect 20376 9052 20416 9092
rect 22156 9640 22196 9680
rect 14380 400 14420 440
rect 18808 8296 18848 8336
rect 18890 8296 18930 8336
rect 18972 8296 19012 8336
rect 19054 8296 19094 8336
rect 19136 8296 19176 8336
rect 20048 7540 20088 7580
rect 20130 7540 20170 7580
rect 20212 7540 20252 7580
rect 20294 7540 20334 7580
rect 20376 7540 20416 7580
rect 18124 6952 18164 6992
rect 18412 6280 18452 6320
rect 17644 3424 17684 3464
rect 18808 6784 18848 6824
rect 18890 6784 18930 6824
rect 18972 6784 19012 6824
rect 19054 6784 19094 6824
rect 19136 6784 19176 6824
rect 20044 6532 20084 6572
rect 20524 6280 20564 6320
rect 20048 6028 20088 6068
rect 20130 6028 20170 6068
rect 20212 6028 20252 6068
rect 20294 6028 20334 6068
rect 20376 6028 20416 6068
rect 20332 5608 20372 5648
rect 18808 5272 18848 5312
rect 18890 5272 18930 5312
rect 18972 5272 19012 5312
rect 19054 5272 19094 5312
rect 19136 5272 19176 5312
rect 18124 4852 18164 4892
rect 17932 4600 17972 4640
rect 18808 3760 18848 3800
rect 18890 3760 18930 3800
rect 18972 3760 19012 3800
rect 19054 3760 19094 3800
rect 19136 3760 19176 3800
rect 18796 3424 18836 3464
rect 18508 2836 18548 2876
rect 18796 2584 18836 2624
rect 19084 2584 19124 2624
rect 19276 3592 19316 3632
rect 18508 1576 18548 1616
rect 18808 2248 18848 2288
rect 18890 2248 18930 2288
rect 18972 2248 19012 2288
rect 19054 2248 19094 2288
rect 19136 2248 19176 2288
rect 19084 1492 19124 1532
rect 18892 1324 18932 1364
rect 19372 1492 19412 1532
rect 19564 3592 19604 3632
rect 19564 1324 19604 1364
rect 20048 4516 20088 4556
rect 20130 4516 20170 4556
rect 20212 4516 20252 4556
rect 20294 4516 20334 4556
rect 20376 4516 20416 4556
rect 20140 3508 20180 3548
rect 20048 3004 20088 3044
rect 20130 3004 20170 3044
rect 20212 3004 20252 3044
rect 20294 3004 20334 3044
rect 20376 3004 20416 3044
rect 20048 1492 20088 1532
rect 20130 1492 20170 1532
rect 20212 1492 20252 1532
rect 20294 1492 20334 1532
rect 20376 1492 20416 1532
rect 20236 1324 20276 1364
rect 20908 6532 20948 6572
rect 20716 1324 20756 1364
rect 21580 6952 21620 6992
rect 21580 5608 21620 5648
rect 22828 4936 22868 4976
rect 23116 4936 23156 4976
rect 23404 1996 23444 2036
rect 24172 3088 24212 3128
rect 24748 3760 24788 3800
rect 24460 3088 24500 3128
rect 24076 2584 24116 2624
rect 24844 1912 24884 1952
rect 25996 4096 26036 4136
rect 25996 3424 26036 3464
rect 25900 2836 25940 2876
rect 26092 2164 26132 2204
rect 30220 10480 30260 10520
rect 26956 4852 26996 4892
rect 27820 4600 27860 4640
rect 27628 3760 27668 3800
rect 27916 3424 27956 3464
rect 27916 2836 27956 2876
rect 28396 2584 28436 2624
rect 27340 2164 27380 2204
rect 27436 1912 27476 1952
rect 28108 1996 28148 2036
rect 30220 9640 30260 9680
rect 35168 10564 35208 10604
rect 35250 10564 35290 10604
rect 35332 10564 35372 10604
rect 35414 10564 35454 10604
rect 35496 10564 35536 10604
rect 29164 4096 29204 4136
rect 30124 3508 30164 3548
rect 31948 400 31988 440
rect 31756 316 31796 356
rect 31372 232 31412 272
rect 31180 64 31220 104
rect 31564 148 31604 188
rect 33928 9808 33968 9848
rect 34010 9808 34050 9848
rect 34092 9808 34132 9848
rect 34174 9808 34214 9848
rect 34256 9808 34296 9848
rect 33100 9556 33140 9596
rect 33292 9556 33332 9596
rect 33196 6448 33236 6488
rect 33292 2860 33332 2900
rect 33484 3004 33524 3044
rect 33388 1912 33428 1952
rect 33484 2860 33524 2900
rect 33580 2080 33620 2120
rect 33928 8296 33968 8336
rect 34010 8296 34050 8336
rect 34092 8296 34132 8336
rect 34174 8296 34214 8336
rect 34256 8296 34296 8336
rect 33928 6784 33968 6824
rect 34010 6784 34050 6824
rect 34092 6784 34132 6824
rect 34174 6784 34214 6824
rect 34256 6784 34296 6824
rect 40300 10480 40340 10520
rect 40396 10144 40436 10184
rect 35168 9052 35208 9092
rect 35250 9052 35290 9092
rect 35332 9052 35372 9092
rect 35414 9052 35454 9092
rect 35496 9052 35536 9092
rect 35168 7540 35208 7580
rect 35250 7540 35290 7580
rect 35332 7540 35372 7580
rect 35414 7540 35454 7580
rect 35496 7540 35536 7580
rect 33928 5272 33968 5312
rect 34010 5272 34050 5312
rect 34092 5272 34132 5312
rect 34174 5272 34214 5312
rect 34256 5272 34296 5312
rect 35168 6028 35208 6068
rect 35250 6028 35290 6068
rect 35332 6028 35372 6068
rect 35414 6028 35454 6068
rect 35496 6028 35536 6068
rect 33928 3760 33968 3800
rect 34010 3760 34050 3800
rect 34092 3760 34132 3800
rect 34174 3760 34214 3800
rect 34256 3760 34296 3800
rect 33772 3004 33812 3044
rect 33928 2248 33968 2288
rect 34010 2248 34050 2288
rect 34092 2248 34132 2288
rect 34174 2248 34214 2288
rect 34256 2248 34296 2288
rect 35168 4516 35208 4556
rect 35250 4516 35290 4556
rect 35332 4516 35372 4556
rect 35414 4516 35454 4556
rect 35496 4516 35536 4556
rect 33676 1912 33716 1952
rect 34060 2080 34100 2120
rect 44524 10144 44564 10184
rect 36940 5356 36980 5396
rect 35168 3004 35208 3044
rect 35250 3004 35290 3044
rect 35332 3004 35372 3044
rect 35414 3004 35454 3044
rect 35496 3004 35536 3044
rect 35168 1492 35208 1532
rect 35250 1492 35290 1532
rect 35332 1492 35372 1532
rect 35414 1492 35454 1532
rect 35496 1492 35536 1532
rect 39340 2752 39380 2792
rect 40108 2416 40148 2456
rect 37900 1744 37940 1784
rect 37612 1408 37652 1448
<< metal4 >>
rect 4919 10564 4928 10604
rect 4968 10564 5010 10604
rect 5050 10564 5092 10604
rect 5132 10564 5174 10604
rect 5214 10564 5256 10604
rect 5296 10564 5305 10604
rect 20039 10564 20048 10604
rect 20088 10564 20130 10604
rect 20170 10564 20212 10604
rect 20252 10564 20294 10604
rect 20334 10564 20376 10604
rect 20416 10564 20425 10604
rect 35159 10564 35168 10604
rect 35208 10564 35250 10604
rect 35290 10564 35332 10604
rect 35372 10564 35414 10604
rect 35454 10564 35496 10604
rect 35536 10564 35545 10604
rect 30211 10480 30220 10520
rect 30260 10480 40300 10520
rect 40340 10480 40349 10520
rect 40387 10144 40396 10184
rect 40436 10144 44524 10184
rect 44564 10144 44573 10184
rect 3679 9808 3688 9848
rect 3728 9808 3770 9848
rect 3810 9808 3852 9848
rect 3892 9808 3934 9848
rect 3974 9808 4016 9848
rect 4056 9808 4065 9848
rect 18799 9808 18808 9848
rect 18848 9808 18890 9848
rect 18930 9808 18972 9848
rect 19012 9808 19054 9848
rect 19094 9808 19136 9848
rect 19176 9808 19185 9848
rect 33919 9808 33928 9848
rect 33968 9808 34010 9848
rect 34050 9808 34092 9848
rect 34132 9808 34174 9848
rect 34214 9808 34256 9848
rect 34296 9808 34305 9848
rect 22147 9640 22156 9680
rect 22196 9640 30220 9680
rect 30260 9640 30269 9680
rect 33091 9556 33100 9596
rect 33140 9556 33292 9596
rect 33332 9556 33341 9596
rect 4919 9052 4928 9092
rect 4968 9052 5010 9092
rect 5050 9052 5092 9092
rect 5132 9052 5174 9092
rect 5214 9052 5256 9092
rect 5296 9052 5305 9092
rect 20039 9052 20048 9092
rect 20088 9052 20130 9092
rect 20170 9052 20212 9092
rect 20252 9052 20294 9092
rect 20334 9052 20376 9092
rect 20416 9052 20425 9092
rect 35159 9052 35168 9092
rect 35208 9052 35250 9092
rect 35290 9052 35332 9092
rect 35372 9052 35414 9092
rect 35454 9052 35496 9092
rect 35536 9052 35545 9092
rect 67 8800 76 8840
rect 116 8800 10060 8840
rect 10100 8800 10109 8840
rect 3679 8296 3688 8336
rect 3728 8296 3770 8336
rect 3810 8296 3852 8336
rect 3892 8296 3934 8336
rect 3974 8296 4016 8336
rect 4056 8296 4065 8336
rect 18799 8296 18808 8336
rect 18848 8296 18890 8336
rect 18930 8296 18972 8336
rect 19012 8296 19054 8336
rect 19094 8296 19136 8336
rect 19176 8296 19185 8336
rect 33919 8296 33928 8336
rect 33968 8296 34010 8336
rect 34050 8296 34092 8336
rect 34132 8296 34174 8336
rect 34214 8296 34256 8336
rect 34296 8296 34305 8336
rect 4919 7540 4928 7580
rect 4968 7540 5010 7580
rect 5050 7540 5092 7580
rect 5132 7540 5174 7580
rect 5214 7540 5256 7580
rect 5296 7540 5305 7580
rect 20039 7540 20048 7580
rect 20088 7540 20130 7580
rect 20170 7540 20212 7580
rect 20252 7540 20294 7580
rect 20334 7540 20376 7580
rect 20416 7540 20425 7580
rect 35159 7540 35168 7580
rect 35208 7540 35250 7580
rect 35290 7540 35332 7580
rect 35372 7540 35414 7580
rect 35454 7540 35496 7580
rect 35536 7540 35545 7580
rect 18115 6952 18124 6992
rect 18164 6952 21580 6992
rect 21620 6952 21629 6992
rect 3679 6784 3688 6824
rect 3728 6784 3770 6824
rect 3810 6784 3852 6824
rect 3892 6784 3934 6824
rect 3974 6784 4016 6824
rect 4056 6784 4065 6824
rect 18799 6784 18808 6824
rect 18848 6784 18890 6824
rect 18930 6784 18972 6824
rect 19012 6784 19054 6824
rect 19094 6784 19136 6824
rect 19176 6784 19185 6824
rect 33919 6784 33928 6824
rect 33968 6784 34010 6824
rect 34050 6784 34092 6824
rect 34132 6784 34174 6824
rect 34214 6784 34256 6824
rect 34296 6784 34305 6824
rect 20035 6532 20044 6572
rect 20084 6532 20908 6572
rect 20948 6532 20957 6572
rect 451 6448 460 6488
rect 500 6448 33196 6488
rect 33236 6448 33245 6488
rect 18403 6280 18412 6320
rect 18452 6280 20524 6320
rect 20564 6280 20573 6320
rect 4919 6028 4928 6068
rect 4968 6028 5010 6068
rect 5050 6028 5092 6068
rect 5132 6028 5174 6068
rect 5214 6028 5256 6068
rect 5296 6028 5305 6068
rect 20039 6028 20048 6068
rect 20088 6028 20130 6068
rect 20170 6028 20212 6068
rect 20252 6028 20294 6068
rect 20334 6028 20376 6068
rect 20416 6028 20425 6068
rect 35159 6028 35168 6068
rect 35208 6028 35250 6068
rect 35290 6028 35332 6068
rect 35372 6028 35414 6068
rect 35454 6028 35496 6068
rect 35536 6028 35545 6068
rect 10531 5608 10540 5648
rect 10580 5608 11980 5648
rect 12020 5608 12029 5648
rect 12643 5608 12652 5648
rect 12692 5608 12940 5648
rect 12980 5608 12989 5648
rect 20323 5608 20332 5648
rect 20372 5608 21580 5648
rect 21620 5608 21629 5648
rect 10051 5356 10060 5396
rect 10100 5356 20180 5396
rect 20140 5312 20180 5356
rect 30220 5356 36940 5396
rect 36980 5356 36989 5396
rect 30220 5312 30260 5356
rect 3679 5272 3688 5312
rect 3728 5272 3770 5312
rect 3810 5272 3852 5312
rect 3892 5272 3934 5312
rect 3974 5272 4016 5312
rect 4056 5272 4065 5312
rect 18799 5272 18808 5312
rect 18848 5272 18890 5312
rect 18930 5272 18972 5312
rect 19012 5272 19054 5312
rect 19094 5272 19136 5312
rect 19176 5272 19185 5312
rect 20140 5272 30260 5312
rect 33919 5272 33928 5312
rect 33968 5272 34010 5312
rect 34050 5272 34092 5312
rect 34132 5272 34174 5312
rect 34214 5272 34256 5312
rect 34296 5272 34305 5312
rect 22819 4936 22828 4976
rect 22868 4936 23116 4976
rect 23156 4936 23165 4976
rect 18115 4852 18124 4892
rect 18164 4852 26956 4892
rect 26996 4852 27005 4892
rect 6691 4600 6700 4640
rect 6740 4600 10060 4640
rect 10100 4600 10109 4640
rect 17923 4600 17932 4640
rect 17972 4600 27820 4640
rect 27860 4600 27869 4640
rect 4919 4516 4928 4556
rect 4968 4516 5010 4556
rect 5050 4516 5092 4556
rect 5132 4516 5174 4556
rect 5214 4516 5256 4556
rect 5296 4516 5305 4556
rect 20039 4516 20048 4556
rect 20088 4516 20130 4556
rect 20170 4516 20212 4556
rect 20252 4516 20294 4556
rect 20334 4516 20376 4556
rect 20416 4516 20425 4556
rect 35159 4516 35168 4556
rect 35208 4516 35250 4556
rect 35290 4516 35332 4556
rect 35372 4516 35414 4556
rect 35454 4516 35496 4556
rect 35536 4516 35545 4556
rect 11683 4180 11692 4220
rect 11732 4180 11924 4220
rect 11884 4136 11924 4180
rect 11875 4096 11884 4136
rect 11924 4096 11933 4136
rect 25987 4096 25996 4136
rect 26036 4096 29164 4136
rect 29204 4096 29213 4136
rect 10627 4012 10636 4052
rect 10676 4012 11692 4052
rect 11732 4012 11741 4052
rect 11779 3928 11788 3968
rect 11828 3928 12076 3968
rect 12116 3928 12125 3968
rect 10051 3844 10060 3884
rect 10100 3844 10444 3884
rect 10484 3844 10493 3884
rect 3679 3760 3688 3800
rect 3728 3760 3770 3800
rect 3810 3760 3852 3800
rect 3892 3760 3934 3800
rect 3974 3760 4016 3800
rect 4056 3760 4065 3800
rect 18799 3760 18808 3800
rect 18848 3760 18890 3800
rect 18930 3760 18972 3800
rect 19012 3760 19054 3800
rect 19094 3760 19136 3800
rect 19176 3760 19185 3800
rect 24739 3760 24748 3800
rect 24788 3760 27628 3800
rect 27668 3760 27677 3800
rect 33919 3760 33928 3800
rect 33968 3760 34010 3800
rect 34050 3760 34092 3800
rect 34132 3760 34174 3800
rect 34214 3760 34256 3800
rect 34296 3760 34305 3800
rect 19267 3592 19276 3632
rect 19316 3592 19564 3632
rect 19604 3592 19613 3632
rect 20131 3508 20140 3548
rect 20180 3508 30124 3548
rect 30164 3508 30173 3548
rect 17635 3424 17644 3464
rect 17684 3424 18796 3464
rect 18836 3424 18845 3464
rect 25987 3424 25996 3464
rect 26036 3424 27916 3464
rect 27956 3424 27965 3464
rect 24163 3088 24172 3128
rect 24212 3088 24460 3128
rect 24500 3088 24509 3128
rect 4919 3004 4928 3044
rect 4968 3004 5010 3044
rect 5050 3004 5092 3044
rect 5132 3004 5174 3044
rect 5214 3004 5256 3044
rect 5296 3004 5305 3044
rect 20039 3004 20048 3044
rect 20088 3004 20130 3044
rect 20170 3004 20212 3044
rect 20252 3004 20294 3044
rect 20334 3004 20376 3044
rect 20416 3004 20425 3044
rect 33292 3004 33484 3044
rect 33524 3004 33533 3044
rect 33580 3004 33772 3044
rect 33812 3004 33821 3044
rect 35159 3004 35168 3044
rect 35208 3004 35250 3044
rect 35290 3004 35332 3044
rect 35372 3004 35414 3044
rect 35454 3004 35496 3044
rect 35536 3004 35545 3044
rect 33292 2900 33332 3004
rect 33580 2900 33620 3004
rect 18413 2836 18508 2876
rect 18548 2836 18557 2876
rect 25891 2836 25900 2876
rect 25940 2836 27916 2876
rect 27956 2836 27965 2876
rect 33283 2860 33292 2900
rect 33332 2860 33341 2900
rect 33475 2860 33484 2900
rect 33524 2860 33620 2900
rect 1411 2752 1420 2792
rect 1460 2752 39340 2792
rect 39380 2752 39389 2792
rect 18787 2584 18796 2624
rect 18836 2584 19084 2624
rect 19124 2584 19133 2624
rect 24067 2584 24076 2624
rect 24116 2584 28396 2624
rect 28436 2584 28445 2624
rect 1411 2416 1420 2456
rect 1460 2416 40108 2456
rect 40148 2416 40157 2456
rect 3679 2248 3688 2288
rect 3728 2248 3770 2288
rect 3810 2248 3852 2288
rect 3892 2248 3934 2288
rect 3974 2248 4016 2288
rect 4056 2248 4065 2288
rect 18799 2248 18808 2288
rect 18848 2248 18890 2288
rect 18930 2248 18972 2288
rect 19012 2248 19054 2288
rect 19094 2248 19136 2288
rect 19176 2248 19185 2288
rect 33919 2248 33928 2288
rect 33968 2248 34010 2288
rect 34050 2248 34092 2288
rect 34132 2248 34174 2288
rect 34214 2248 34256 2288
rect 34296 2248 34305 2288
rect 26083 2164 26092 2204
rect 26132 2164 27340 2204
rect 27380 2164 27389 2204
rect 33571 2080 33580 2120
rect 33620 2080 34060 2120
rect 34100 2080 34109 2120
rect 23395 1996 23404 2036
rect 23444 1996 28108 2036
rect 28148 1996 28157 2036
rect 24835 1912 24844 1952
rect 24884 1912 27436 1952
rect 27476 1912 27485 1952
rect 33379 1912 33388 1952
rect 33428 1912 33676 1952
rect 33716 1912 33725 1952
rect 1411 1744 1420 1784
rect 1460 1744 37900 1784
rect 37940 1744 37949 1784
rect 18413 1576 18508 1616
rect 18548 1576 18557 1616
rect 4919 1492 4928 1532
rect 4968 1492 5010 1532
rect 5050 1492 5092 1532
rect 5132 1492 5174 1532
rect 5214 1492 5256 1532
rect 5296 1492 5305 1532
rect 19075 1492 19084 1532
rect 19124 1492 19372 1532
rect 19412 1492 19421 1532
rect 20039 1492 20048 1532
rect 20088 1492 20130 1532
rect 20170 1492 20212 1532
rect 20252 1492 20294 1532
rect 20334 1492 20376 1532
rect 20416 1492 20425 1532
rect 35159 1492 35168 1532
rect 35208 1492 35250 1532
rect 35290 1492 35332 1532
rect 35372 1492 35414 1532
rect 35454 1492 35496 1532
rect 35536 1492 35545 1532
rect 1411 1408 1420 1448
rect 1460 1408 37612 1448
rect 37652 1408 37661 1448
rect 18883 1324 18892 1364
rect 18932 1324 19564 1364
rect 19604 1324 19613 1364
rect 20227 1324 20236 1364
rect 20276 1324 20716 1364
rect 20756 1324 20765 1364
rect 14371 400 14380 440
rect 14420 400 31948 440
rect 31988 400 31997 440
rect 7459 316 7468 356
rect 7508 316 31756 356
rect 31796 316 31805 356
rect 6883 232 6892 272
rect 6932 232 31372 272
rect 31412 232 31421 272
rect 6403 148 6412 188
rect 6452 148 31564 188
rect 31604 148 31613 188
rect 8803 64 8812 104
rect 8852 64 31180 104
rect 31220 64 31229 104
<< via4 >>
rect 4928 10564 4968 10604
rect 5010 10564 5050 10604
rect 5092 10564 5132 10604
rect 5174 10564 5214 10604
rect 5256 10564 5296 10604
rect 20048 10564 20088 10604
rect 20130 10564 20170 10604
rect 20212 10564 20252 10604
rect 20294 10564 20334 10604
rect 20376 10564 20416 10604
rect 35168 10564 35208 10604
rect 35250 10564 35290 10604
rect 35332 10564 35372 10604
rect 35414 10564 35454 10604
rect 35496 10564 35536 10604
rect 3688 9808 3728 9848
rect 3770 9808 3810 9848
rect 3852 9808 3892 9848
rect 3934 9808 3974 9848
rect 4016 9808 4056 9848
rect 18808 9808 18848 9848
rect 18890 9808 18930 9848
rect 18972 9808 19012 9848
rect 19054 9808 19094 9848
rect 19136 9808 19176 9848
rect 33928 9808 33968 9848
rect 34010 9808 34050 9848
rect 34092 9808 34132 9848
rect 34174 9808 34214 9848
rect 34256 9808 34296 9848
rect 4928 9052 4968 9092
rect 5010 9052 5050 9092
rect 5092 9052 5132 9092
rect 5174 9052 5214 9092
rect 5256 9052 5296 9092
rect 20048 9052 20088 9092
rect 20130 9052 20170 9092
rect 20212 9052 20252 9092
rect 20294 9052 20334 9092
rect 20376 9052 20416 9092
rect 35168 9052 35208 9092
rect 35250 9052 35290 9092
rect 35332 9052 35372 9092
rect 35414 9052 35454 9092
rect 35496 9052 35536 9092
rect 3688 8296 3728 8336
rect 3770 8296 3810 8336
rect 3852 8296 3892 8336
rect 3934 8296 3974 8336
rect 4016 8296 4056 8336
rect 18808 8296 18848 8336
rect 18890 8296 18930 8336
rect 18972 8296 19012 8336
rect 19054 8296 19094 8336
rect 19136 8296 19176 8336
rect 33928 8296 33968 8336
rect 34010 8296 34050 8336
rect 34092 8296 34132 8336
rect 34174 8296 34214 8336
rect 34256 8296 34296 8336
rect 4928 7540 4968 7580
rect 5010 7540 5050 7580
rect 5092 7540 5132 7580
rect 5174 7540 5214 7580
rect 5256 7540 5296 7580
rect 20048 7540 20088 7580
rect 20130 7540 20170 7580
rect 20212 7540 20252 7580
rect 20294 7540 20334 7580
rect 20376 7540 20416 7580
rect 35168 7540 35208 7580
rect 35250 7540 35290 7580
rect 35332 7540 35372 7580
rect 35414 7540 35454 7580
rect 35496 7540 35536 7580
rect 3688 6784 3728 6824
rect 3770 6784 3810 6824
rect 3852 6784 3892 6824
rect 3934 6784 3974 6824
rect 4016 6784 4056 6824
rect 18808 6784 18848 6824
rect 18890 6784 18930 6824
rect 18972 6784 19012 6824
rect 19054 6784 19094 6824
rect 19136 6784 19176 6824
rect 33928 6784 33968 6824
rect 34010 6784 34050 6824
rect 34092 6784 34132 6824
rect 34174 6784 34214 6824
rect 34256 6784 34296 6824
rect 4928 6028 4968 6068
rect 5010 6028 5050 6068
rect 5092 6028 5132 6068
rect 5174 6028 5214 6068
rect 5256 6028 5296 6068
rect 20048 6028 20088 6068
rect 20130 6028 20170 6068
rect 20212 6028 20252 6068
rect 20294 6028 20334 6068
rect 20376 6028 20416 6068
rect 35168 6028 35208 6068
rect 35250 6028 35290 6068
rect 35332 6028 35372 6068
rect 35414 6028 35454 6068
rect 35496 6028 35536 6068
rect 3688 5272 3728 5312
rect 3770 5272 3810 5312
rect 3852 5272 3892 5312
rect 3934 5272 3974 5312
rect 4016 5272 4056 5312
rect 18808 5272 18848 5312
rect 18890 5272 18930 5312
rect 18972 5272 19012 5312
rect 19054 5272 19094 5312
rect 19136 5272 19176 5312
rect 33928 5272 33968 5312
rect 34010 5272 34050 5312
rect 34092 5272 34132 5312
rect 34174 5272 34214 5312
rect 34256 5272 34296 5312
rect 4928 4516 4968 4556
rect 5010 4516 5050 4556
rect 5092 4516 5132 4556
rect 5174 4516 5214 4556
rect 5256 4516 5296 4556
rect 20048 4516 20088 4556
rect 20130 4516 20170 4556
rect 20212 4516 20252 4556
rect 20294 4516 20334 4556
rect 20376 4516 20416 4556
rect 35168 4516 35208 4556
rect 35250 4516 35290 4556
rect 35332 4516 35372 4556
rect 35414 4516 35454 4556
rect 35496 4516 35536 4556
rect 3688 3760 3728 3800
rect 3770 3760 3810 3800
rect 3852 3760 3892 3800
rect 3934 3760 3974 3800
rect 4016 3760 4056 3800
rect 18808 3760 18848 3800
rect 18890 3760 18930 3800
rect 18972 3760 19012 3800
rect 19054 3760 19094 3800
rect 19136 3760 19176 3800
rect 33928 3760 33968 3800
rect 34010 3760 34050 3800
rect 34092 3760 34132 3800
rect 34174 3760 34214 3800
rect 34256 3760 34296 3800
rect 4928 3004 4968 3044
rect 5010 3004 5050 3044
rect 5092 3004 5132 3044
rect 5174 3004 5214 3044
rect 5256 3004 5296 3044
rect 20048 3004 20088 3044
rect 20130 3004 20170 3044
rect 20212 3004 20252 3044
rect 20294 3004 20334 3044
rect 20376 3004 20416 3044
rect 35168 3004 35208 3044
rect 35250 3004 35290 3044
rect 35332 3004 35372 3044
rect 35414 3004 35454 3044
rect 35496 3004 35536 3044
rect 18508 2836 18548 2876
rect 3688 2248 3728 2288
rect 3770 2248 3810 2288
rect 3852 2248 3892 2288
rect 3934 2248 3974 2288
rect 4016 2248 4056 2288
rect 18808 2248 18848 2288
rect 18890 2248 18930 2288
rect 18972 2248 19012 2288
rect 19054 2248 19094 2288
rect 19136 2248 19176 2288
rect 33928 2248 33968 2288
rect 34010 2248 34050 2288
rect 34092 2248 34132 2288
rect 34174 2248 34214 2288
rect 34256 2248 34296 2288
rect 18508 1576 18548 1616
rect 4928 1492 4968 1532
rect 5010 1492 5050 1532
rect 5092 1492 5132 1532
rect 5174 1492 5214 1532
rect 5256 1492 5296 1532
rect 20048 1492 20088 1532
rect 20130 1492 20170 1532
rect 20212 1492 20252 1532
rect 20294 1492 20334 1532
rect 20376 1492 20416 1532
rect 35168 1492 35208 1532
rect 35250 1492 35290 1532
rect 35332 1492 35372 1532
rect 35414 1492 35454 1532
rect 35496 1492 35536 1532
<< metal5 >>
rect 3652 9848 4092 12180
rect 3652 9808 3688 9848
rect 3728 9808 3770 9848
rect 3810 9808 3852 9848
rect 3892 9808 3934 9848
rect 3974 9808 4016 9848
rect 4056 9808 4092 9848
rect 3652 8336 4092 9808
rect 3652 8296 3688 8336
rect 3728 8296 3770 8336
rect 3810 8296 3852 8336
rect 3892 8296 3934 8336
rect 3974 8296 4016 8336
rect 4056 8296 4092 8336
rect 3652 6824 4092 8296
rect 3652 6784 3688 6824
rect 3728 6784 3770 6824
rect 3810 6784 3852 6824
rect 3892 6784 3934 6824
rect 3974 6784 4016 6824
rect 4056 6784 4092 6824
rect 3652 5312 4092 6784
rect 3652 5272 3688 5312
rect 3728 5272 3770 5312
rect 3810 5272 3852 5312
rect 3892 5272 3934 5312
rect 3974 5272 4016 5312
rect 4056 5272 4092 5312
rect 3652 3800 4092 5272
rect 3652 3760 3688 3800
rect 3728 3760 3770 3800
rect 3810 3760 3852 3800
rect 3892 3760 3934 3800
rect 3974 3760 4016 3800
rect 4056 3760 4092 3800
rect 3652 2288 4092 3760
rect 3652 2248 3688 2288
rect 3728 2248 3770 2288
rect 3810 2248 3852 2288
rect 3892 2248 3934 2288
rect 3974 2248 4016 2288
rect 4056 2248 4092 2288
rect 3652 0 4092 2248
rect 4892 10604 5332 12180
rect 4892 10564 4928 10604
rect 4968 10564 5010 10604
rect 5050 10564 5092 10604
rect 5132 10564 5174 10604
rect 5214 10564 5256 10604
rect 5296 10564 5332 10604
rect 4892 9092 5332 10564
rect 4892 9052 4928 9092
rect 4968 9052 5010 9092
rect 5050 9052 5092 9092
rect 5132 9052 5174 9092
rect 5214 9052 5256 9092
rect 5296 9052 5332 9092
rect 4892 7580 5332 9052
rect 4892 7540 4928 7580
rect 4968 7540 5010 7580
rect 5050 7540 5092 7580
rect 5132 7540 5174 7580
rect 5214 7540 5256 7580
rect 5296 7540 5332 7580
rect 4892 6068 5332 7540
rect 4892 6028 4928 6068
rect 4968 6028 5010 6068
rect 5050 6028 5092 6068
rect 5132 6028 5174 6068
rect 5214 6028 5256 6068
rect 5296 6028 5332 6068
rect 4892 4556 5332 6028
rect 4892 4516 4928 4556
rect 4968 4516 5010 4556
rect 5050 4516 5092 4556
rect 5132 4516 5174 4556
rect 5214 4516 5256 4556
rect 5296 4516 5332 4556
rect 4892 3044 5332 4516
rect 4892 3004 4928 3044
rect 4968 3004 5010 3044
rect 5050 3004 5092 3044
rect 5132 3004 5174 3044
rect 5214 3004 5256 3044
rect 5296 3004 5332 3044
rect 4892 1532 5332 3004
rect 18772 9848 19212 12180
rect 18772 9808 18808 9848
rect 18848 9808 18890 9848
rect 18930 9808 18972 9848
rect 19012 9808 19054 9848
rect 19094 9808 19136 9848
rect 19176 9808 19212 9848
rect 18772 8336 19212 9808
rect 18772 8296 18808 8336
rect 18848 8296 18890 8336
rect 18930 8296 18972 8336
rect 19012 8296 19054 8336
rect 19094 8296 19136 8336
rect 19176 8296 19212 8336
rect 18772 6824 19212 8296
rect 18772 6784 18808 6824
rect 18848 6784 18890 6824
rect 18930 6784 18972 6824
rect 19012 6784 19054 6824
rect 19094 6784 19136 6824
rect 19176 6784 19212 6824
rect 18772 5312 19212 6784
rect 18772 5272 18808 5312
rect 18848 5272 18890 5312
rect 18930 5272 18972 5312
rect 19012 5272 19054 5312
rect 19094 5272 19136 5312
rect 19176 5272 19212 5312
rect 18772 3800 19212 5272
rect 18772 3760 18808 3800
rect 18848 3760 18890 3800
rect 18930 3760 18972 3800
rect 19012 3760 19054 3800
rect 19094 3760 19136 3800
rect 19176 3760 19212 3800
rect 18508 2876 18548 2885
rect 18508 1616 18548 2836
rect 18508 1567 18548 1576
rect 18772 2288 19212 3760
rect 18772 2248 18808 2288
rect 18848 2248 18890 2288
rect 18930 2248 18972 2288
rect 19012 2248 19054 2288
rect 19094 2248 19136 2288
rect 19176 2248 19212 2288
rect 4892 1492 4928 1532
rect 4968 1492 5010 1532
rect 5050 1492 5092 1532
rect 5132 1492 5174 1532
rect 5214 1492 5256 1532
rect 5296 1492 5332 1532
rect 4892 0 5332 1492
rect 18772 0 19212 2248
rect 20012 10604 20452 12180
rect 20012 10564 20048 10604
rect 20088 10564 20130 10604
rect 20170 10564 20212 10604
rect 20252 10564 20294 10604
rect 20334 10564 20376 10604
rect 20416 10564 20452 10604
rect 20012 9092 20452 10564
rect 20012 9052 20048 9092
rect 20088 9052 20130 9092
rect 20170 9052 20212 9092
rect 20252 9052 20294 9092
rect 20334 9052 20376 9092
rect 20416 9052 20452 9092
rect 20012 7580 20452 9052
rect 20012 7540 20048 7580
rect 20088 7540 20130 7580
rect 20170 7540 20212 7580
rect 20252 7540 20294 7580
rect 20334 7540 20376 7580
rect 20416 7540 20452 7580
rect 20012 6068 20452 7540
rect 20012 6028 20048 6068
rect 20088 6028 20130 6068
rect 20170 6028 20212 6068
rect 20252 6028 20294 6068
rect 20334 6028 20376 6068
rect 20416 6028 20452 6068
rect 20012 4556 20452 6028
rect 20012 4516 20048 4556
rect 20088 4516 20130 4556
rect 20170 4516 20212 4556
rect 20252 4516 20294 4556
rect 20334 4516 20376 4556
rect 20416 4516 20452 4556
rect 20012 3044 20452 4516
rect 20012 3004 20048 3044
rect 20088 3004 20130 3044
rect 20170 3004 20212 3044
rect 20252 3004 20294 3044
rect 20334 3004 20376 3044
rect 20416 3004 20452 3044
rect 20012 1532 20452 3004
rect 20012 1492 20048 1532
rect 20088 1492 20130 1532
rect 20170 1492 20212 1532
rect 20252 1492 20294 1532
rect 20334 1492 20376 1532
rect 20416 1492 20452 1532
rect 20012 0 20452 1492
rect 33892 9848 34332 12180
rect 33892 9808 33928 9848
rect 33968 9808 34010 9848
rect 34050 9808 34092 9848
rect 34132 9808 34174 9848
rect 34214 9808 34256 9848
rect 34296 9808 34332 9848
rect 33892 8336 34332 9808
rect 33892 8296 33928 8336
rect 33968 8296 34010 8336
rect 34050 8296 34092 8336
rect 34132 8296 34174 8336
rect 34214 8296 34256 8336
rect 34296 8296 34332 8336
rect 33892 6824 34332 8296
rect 33892 6784 33928 6824
rect 33968 6784 34010 6824
rect 34050 6784 34092 6824
rect 34132 6784 34174 6824
rect 34214 6784 34256 6824
rect 34296 6784 34332 6824
rect 33892 5312 34332 6784
rect 33892 5272 33928 5312
rect 33968 5272 34010 5312
rect 34050 5272 34092 5312
rect 34132 5272 34174 5312
rect 34214 5272 34256 5312
rect 34296 5272 34332 5312
rect 33892 3800 34332 5272
rect 33892 3760 33928 3800
rect 33968 3760 34010 3800
rect 34050 3760 34092 3800
rect 34132 3760 34174 3800
rect 34214 3760 34256 3800
rect 34296 3760 34332 3800
rect 33892 2288 34332 3760
rect 33892 2248 33928 2288
rect 33968 2248 34010 2288
rect 34050 2248 34092 2288
rect 34132 2248 34174 2288
rect 34214 2248 34256 2288
rect 34296 2248 34332 2288
rect 33892 0 34332 2248
rect 35132 10604 35572 12180
rect 35132 10564 35168 10604
rect 35208 10564 35250 10604
rect 35290 10564 35332 10604
rect 35372 10564 35414 10604
rect 35454 10564 35496 10604
rect 35536 10564 35572 10604
rect 35132 9092 35572 10564
rect 35132 9052 35168 9092
rect 35208 9052 35250 9092
rect 35290 9052 35332 9092
rect 35372 9052 35414 9092
rect 35454 9052 35496 9092
rect 35536 9052 35572 9092
rect 35132 7580 35572 9052
rect 35132 7540 35168 7580
rect 35208 7540 35250 7580
rect 35290 7540 35332 7580
rect 35372 7540 35414 7580
rect 35454 7540 35496 7580
rect 35536 7540 35572 7580
rect 35132 6068 35572 7540
rect 35132 6028 35168 6068
rect 35208 6028 35250 6068
rect 35290 6028 35332 6068
rect 35372 6028 35414 6068
rect 35454 6028 35496 6068
rect 35536 6028 35572 6068
rect 35132 4556 35572 6028
rect 35132 4516 35168 4556
rect 35208 4516 35250 4556
rect 35290 4516 35332 4556
rect 35372 4516 35414 4556
rect 35454 4516 35496 4556
rect 35536 4516 35572 4556
rect 35132 3044 35572 4516
rect 35132 3004 35168 3044
rect 35208 3004 35250 3044
rect 35290 3004 35332 3044
rect 35372 3004 35414 3044
rect 35454 3004 35496 3044
rect 35536 3004 35572 3044
rect 35132 1532 35572 3004
rect 35132 1492 35168 1532
rect 35208 1492 35250 1532
rect 35290 1492 35332 1532
rect 35372 1492 35414 1532
rect 35454 1492 35496 1532
rect 35536 1492 35572 1532
rect 35132 0 35572 1492
use sg13g2_buf_1  _000_
timestamp 1676381911
transform 1 0 33120 0 1 6048
box -48 -56 432 834
use sg13g2_buf_1  _001_
timestamp 1676381911
transform 1 0 36864 0 -1 6048
box -48 -56 432 834
use sg13g2_buf_1  _002_
timestamp 1676381911
transform 1 0 38400 0 -1 6048
box -48 -56 432 834
use sg13g2_buf_1  _003_
timestamp 1676381911
transform 1 0 38016 0 -1 6048
box -48 -56 432 834
use sg13g2_buf_1  _004_
timestamp 1676381911
transform 1 0 34080 0 -1 6048
box -48 -56 432 834
use sg13g2_buf_1  _005_
timestamp 1676381911
transform 1 0 41088 0 1 4536
box -48 -56 432 834
use sg13g2_buf_1  _006_
timestamp 1676381911
transform 1 0 40704 0 1 4536
box -48 -56 432 834
use sg13g2_buf_1  _007_
timestamp 1676381911
transform 1 0 38592 0 1 4536
box -48 -56 432 834
use sg13g2_buf_1  _008_
timestamp 1676381911
transform 1 0 39552 0 1 4536
box -48 -56 432 834
use sg13g2_buf_1  _009_
timestamp 1676381911
transform 1 0 32544 0 -1 4536
box -48 -56 432 834
use sg13g2_buf_1  _010_
timestamp 1676381911
transform 1 0 37824 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  _011_
timestamp 1676381911
transform 1 0 36480 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  _012_
timestamp 1676381911
transform 1 0 34752 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  _013_
timestamp 1676381911
transform 1 0 30624 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  _014_
timestamp 1676381911
transform 1 0 26976 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  _015_
timestamp 1676381911
transform 1 0 27360 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  _016_
timestamp 1676381911
transform 1 0 28128 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  _017_
timestamp 1676381911
transform 1 0 29952 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  _018_
timestamp 1676381911
transform 1 0 26208 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  _019_
timestamp 1676381911
transform 1 0 27648 0 1 4536
box -48 -56 432 834
use sg13g2_buf_1  _020_
timestamp 1676381911
transform 1 0 25344 0 1 7560
box -48 -56 432 834
use sg13g2_buf_1  _021_
timestamp 1676381911
transform 1 0 23136 0 -1 9072
box -48 -56 432 834
use sg13g2_buf_1  _022_
timestamp 1676381911
transform 1 0 27648 0 -1 9072
box -48 -56 432 834
use sg13g2_buf_1  _023_
timestamp 1676381911
transform 1 0 21600 0 -1 9072
box -48 -56 432 834
use sg13g2_buf_1  _024_
timestamp 1676381911
transform 1 0 24096 0 -1 9072
box -48 -56 432 834
use sg13g2_buf_1  _025_
timestamp 1676381911
transform 1 0 23520 0 -1 9072
box -48 -56 432 834
use sg13g2_buf_1  _026_
timestamp 1676381911
transform 1 0 24672 0 1 7560
box -48 -56 432 834
use sg13g2_buf_1  _027_
timestamp 1676381911
transform 1 0 22368 0 -1 9072
box -48 -56 432 834
use sg13g2_buf_1  _028_
timestamp 1676381911
transform 1 0 22752 0 -1 9072
box -48 -56 432 834
use sg13g2_buf_1  _029_
timestamp 1676381911
transform 1 0 21216 0 -1 9072
box -48 -56 432 834
use sg13g2_buf_1  _030_
timestamp 1676381911
transform 1 0 21984 0 -1 9072
box -48 -56 432 834
use sg13g2_buf_1  _031_
timestamp 1676381911
transform 1 0 26208 0 1 7560
box -48 -56 432 834
use sg13g2_buf_1  _032_
timestamp 1676381911
transform -1 0 7008 0 -1 9072
box -48 -56 432 834
use sg13g2_buf_1  _033_
timestamp 1676381911
transform -1 0 6528 0 -1 9072
box -48 -56 432 834
use sg13g2_buf_1  _034_
timestamp 1676381911
transform 1 0 7392 0 -1 9072
box -48 -56 432 834
use sg13g2_buf_1  _035_
timestamp 1676381911
transform -1 0 13440 0 -1 9072
box -48 -56 432 834
use sg13g2_buf_1  _036_
timestamp 1676381911
transform -1 0 19104 0 -1 9072
box -48 -56 432 834
use sg13g2_buf_1  _037_
timestamp 1676381911
transform -1 0 26208 0 -1 9072
box -48 -56 432 834
use sg13g2_buf_1  _038_
timestamp 1676381911
transform -1 0 31584 0 -1 9072
box -48 -56 432 834
use sg13g2_buf_1  _039_
timestamp 1676381911
transform -1 0 31968 0 -1 9072
box -48 -56 432 834
use sg13g2_buf_1  _040_
timestamp 1676381911
transform -1 0 29472 0 -1 9072
box -48 -56 432 834
use sg13g2_buf_1  _041_
timestamp 1676381911
transform -1 0 27264 0 -1 9072
box -48 -56 432 834
use sg13g2_buf_1  _042_
timestamp 1676381911
transform -1 0 27648 0 -1 9072
box -48 -56 432 834
use sg13g2_buf_1  _043_
timestamp 1676381911
transform -1 0 28416 0 -1 9072
box -48 -56 432 834
use sg13g2_buf_1  _044_
timestamp 1676381911
transform 1 0 28416 0 -1 9072
box -48 -56 432 834
use sg13g2_buf_1  _045_
timestamp 1676381911
transform 1 0 27744 0 1 7560
box -48 -56 432 834
use sg13g2_buf_1  _046_
timestamp 1676381911
transform 1 0 28512 0 1 7560
box -48 -56 432 834
use sg13g2_buf_1  _047_
timestamp 1676381911
transform 1 0 28032 0 1 6048
box -48 -56 432 834
use sg13g2_buf_1  _048_
timestamp 1676381911
transform 1 0 27552 0 -1 4536
box -48 -56 432 834
use sg13g2_buf_1  _049_
timestamp 1676381911
transform 1 0 26592 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  _050_
timestamp 1676381911
transform 1 0 25824 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  _051_
timestamp 1676381911
transform 1 0 27744 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  _052_
timestamp 1676381911
transform 1 0 8256 0 1 4536
box -48 -56 432 834
use sg13g2_buf_1  _053_
timestamp 1676381911
transform 1 0 7488 0 1 4536
box -48 -56 432 834
use sg13g2_buf_1  _054_
timestamp 1676381911
transform 1 0 7104 0 1 4536
box -48 -56 432 834
use sg13g2_buf_1  _055_
timestamp 1676381911
transform 1 0 7008 0 -1 4536
box -48 -56 432 834
use sg13g2_buf_1  _056_
timestamp 1676381911
transform 1 0 13440 0 -1 6048
box -48 -56 432 834
use sg13g2_buf_1  _057_
timestamp 1676381911
transform 1 0 12192 0 -1 6048
box -48 -56 432 834
use sg13g2_buf_1  _058_
timestamp 1676381911
transform 1 0 11424 0 -1 6048
box -48 -56 432 834
use sg13g2_buf_1  _059_
timestamp 1676381911
transform 1 0 10752 0 -1 6048
box -48 -56 432 834
use sg13g2_buf_1  _060_
timestamp 1676381911
transform 1 0 9792 0 -1 6048
box -48 -56 432 834
use sg13g2_buf_1  _061_
timestamp 1676381911
transform 1 0 8640 0 -1 6048
box -48 -56 432 834
use sg13g2_buf_1  _062_
timestamp 1676381911
transform 1 0 7488 0 -1 6048
box -48 -56 432 834
use sg13g2_buf_1  _063_
timestamp 1676381911
transform 1 0 6624 0 -1 6048
box -48 -56 432 834
use sg13g2_buf_1  _064_
timestamp 1676381911
transform 1 0 17664 0 -1 7560
box -48 -56 432 834
use sg13g2_buf_1  _065_
timestamp 1676381911
transform 1 0 17280 0 -1 7560
box -48 -56 432 834
use sg13g2_buf_1  _066_
timestamp 1676381911
transform 1 0 16800 0 -1 7560
box -48 -56 432 834
use sg13g2_buf_1  _067_
timestamp 1676381911
transform 1 0 16032 0 -1 7560
box -48 -56 432 834
use sg13g2_buf_1  _068_
timestamp 1676381911
transform 1 0 14880 0 -1 7560
box -48 -56 432 834
use sg13g2_buf_1  _069_
timestamp 1676381911
transform 1 0 13824 0 -1 7560
box -48 -56 432 834
use sg13g2_buf_1  _070_
timestamp 1676381911
transform 1 0 12384 0 -1 7560
box -48 -56 432 834
use sg13g2_buf_1  _071_
timestamp 1676381911
transform 1 0 10752 0 1 6048
box -48 -56 432 834
use sg13g2_buf_1  _072_
timestamp 1676381911
transform 1 0 20352 0 -1 7560
box -48 -56 432 834
use sg13g2_buf_1  _073_
timestamp 1676381911
transform 1 0 20736 0 -1 7560
box -48 -56 432 834
use sg13g2_buf_1  _074_
timestamp 1676381911
transform 1 0 21120 0 -1 7560
box -48 -56 432 834
use sg13g2_buf_1  _075_
timestamp 1676381911
transform 1 0 19968 0 -1 7560
box -48 -56 432 834
use sg13g2_buf_1  _076_
timestamp 1676381911
transform 1 0 19584 0 -1 7560
box -48 -56 432 834
use sg13g2_buf_1  _077_
timestamp 1676381911
transform 1 0 19200 0 -1 7560
box -48 -56 432 834
use sg13g2_buf_1  _078_
timestamp 1676381911
transform 1 0 18816 0 -1 7560
box -48 -56 432 834
use sg13g2_buf_1  _079_
timestamp 1676381911
transform 1 0 18432 0 -1 7560
box -48 -56 432 834
use sg13g2_buf_1  _080_
timestamp 1676381911
transform 1 0 18048 0 -1 7560
box -48 -56 432 834
use sg13g2_buf_1  _081_
timestamp 1676381911
transform 1 0 18336 0 1 7560
box -48 -56 432 834
use sg13g2_buf_1  _082_
timestamp 1676381911
transform 1 0 18720 0 1 7560
box -48 -56 432 834
use sg13g2_buf_1  _083_
timestamp 1676381911
transform 1 0 17664 0 1 7560
box -48 -56 432 834
use sg13g2_buf_1  _084_
timestamp 1676381911
transform 1 0 17280 0 1 7560
box -48 -56 432 834
use sg13g2_buf_1  _085_
timestamp 1676381911
transform 1 0 16896 0 1 7560
box -48 -56 432 834
use sg13g2_buf_1  _086_
timestamp 1676381911
transform 1 0 16512 0 1 7560
box -48 -56 432 834
use sg13g2_buf_1  _087_
timestamp 1676381911
transform 1 0 16128 0 1 7560
box -48 -56 432 834
use sg13g2_buf_1  _088_
timestamp 1676381911
transform 1 0 19872 0 1 6048
box -48 -56 432 834
use sg13g2_buf_1  _089_
timestamp 1676381911
transform 1 0 20352 0 1 6048
box -48 -56 432 834
use sg13g2_buf_1  _090_
timestamp 1676381911
transform 1 0 20928 0 -1 6048
box -48 -56 432 834
use sg13g2_buf_1  _091_
timestamp 1676381911
transform 1 0 21312 0 -1 6048
box -48 -56 432 834
use sg13g2_buf_1  _092_
timestamp 1676381911
transform 1 0 21696 0 -1 6048
box -48 -56 432 834
use sg13g2_buf_1  _093_
timestamp 1676381911
transform 1 0 21984 0 1 4536
box -48 -56 432 834
use sg13g2_buf_1  _094_
timestamp 1676381911
transform 1 0 22368 0 1 4536
box -48 -56 432 834
use sg13g2_buf_1  _095_
timestamp 1676381911
transform 1 0 22848 0 1 4536
box -48 -56 432 834
use sg13g2_buf_1  _096_
timestamp 1676381911
transform 1 0 23328 0 1 4536
box -48 -56 432 834
use sg13g2_buf_1  _097_
timestamp 1676381911
transform 1 0 23904 0 -1 4536
box -48 -56 432 834
use sg13g2_buf_1  _098_
timestamp 1676381911
transform 1 0 24384 0 -1 4536
box -48 -56 432 834
use sg13g2_buf_1  _099_
timestamp 1676381911
transform 1 0 25248 0 -1 4536
box -48 -56 432 834
use sg13g2_buf_1  _100_
timestamp 1676381911
transform 1 0 26112 0 -1 4536
box -48 -56 432 834
use sg13g2_buf_1  _101_
timestamp 1676381911
transform 1 0 26784 0 1 4536
box -48 -56 432 834
use sg13g2_buf_1  _102_
timestamp 1676381911
transform 1 0 28032 0 1 4536
box -48 -56 432 834
use sg13g2_buf_1  _103_
timestamp 1676381911
transform 1 0 28416 0 1 4536
box -48 -56 432 834
use sg13g2_buf_1  _104_
timestamp 1676381911
transform -1 0 8928 0 -1 9072
box -48 -56 432 834
use sg13g2_antennanp  ANTENNA_1
timestamp 1679999689
transform 1 0 35040 0 -1 3024
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_2
timestamp 1679999689
transform -1 0 37632 0 -1 6048
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_3
timestamp 1679999689
transform 1 0 37632 0 1 4536
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_4
timestamp 1679999689
transform 1 0 34368 0 1 4536
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_5
timestamp 1679999689
transform 1 0 41760 0 1 4536
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_6
timestamp 1679999689
transform 1 0 42720 0 -1 4536
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_7
timestamp 1679999689
transform 1 0 39264 0 -1 4536
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_8
timestamp 1679999689
transform 1 0 42432 0 -1 4536
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_9
timestamp 1679999689
transform 1 0 38304 0 1 4536
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_10
timestamp 1679999689
transform -1 0 35040 0 -1 3024
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_11
timestamp 1679999689
transform -1 0 38016 0 -1 6048
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_12
timestamp 1679999689
transform 1 0 34080 0 1 4536
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_13
timestamp 1679999689
transform 1 0 41472 0 1 4536
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_14
timestamp 1679999689
transform 1 0 42144 0 -1 4536
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_15
timestamp 1679999689
transform 1 0 39264 0 1 4536
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_16
timestamp 1679999689
transform 1 0 39936 0 -1 4536
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_17
timestamp 1679999689
transform 1 0 38976 0 1 4536
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_18
timestamp 1679999689
transform 1 0 40032 0 1 4536
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_19
timestamp 1679999689
transform 1 0 41856 0 -1 4536
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_20
timestamp 1679999689
transform 1 0 41568 0 -1 4536
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_21
timestamp 1679999689
transform 1 0 41280 0 -1 4536
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_22
timestamp 1679999689
transform 1 0 40992 0 -1 4536
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_23
timestamp 1679999689
transform 1 0 40704 0 -1 4536
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_24
timestamp 1679999689
transform 1 0 40416 0 -1 4536
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_25
timestamp 1679999689
transform 1 0 40416 0 1 4536
box -48 -56 336 834
use sg13g2_decap_8  FILLER_0_0
timestamp 1679581782
transform 1 0 1152 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_7
timestamp 1679581782
transform 1 0 1824 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_14
timestamp 1679581782
transform 1 0 2496 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_21
timestamp 1679581782
transform 1 0 3168 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_28
timestamp 1679581782
transform 1 0 3840 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_35
timestamp 1679581782
transform 1 0 4512 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_42
timestamp 1679581782
transform 1 0 5184 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_49
timestamp 1679581782
transform 1 0 5856 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_56
timestamp 1679581782
transform 1 0 6528 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_63
timestamp 1679581782
transform 1 0 7200 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_70
timestamp 1679581782
transform 1 0 7872 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_77
timestamp 1679581782
transform 1 0 8544 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_84
timestamp 1679581782
transform 1 0 9216 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_91
timestamp 1679581782
transform 1 0 9888 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_98
timestamp 1679581782
transform 1 0 10560 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_105
timestamp 1679581782
transform 1 0 11232 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_112
timestamp 1679581782
transform 1 0 11904 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_119
timestamp 1679581782
transform 1 0 12576 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_126
timestamp 1679581782
transform 1 0 13248 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_133
timestamp 1679581782
transform 1 0 13920 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_140
timestamp 1679581782
transform 1 0 14592 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_147
timestamp 1679581782
transform 1 0 15264 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_154
timestamp 1679581782
transform 1 0 15936 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_161
timestamp 1679581782
transform 1 0 16608 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_168
timestamp 1679581782
transform 1 0 17280 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_175
timestamp 1679581782
transform 1 0 17952 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_182
timestamp 1679581782
transform 1 0 18624 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_189
timestamp 1679581782
transform 1 0 19296 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_196
timestamp 1679581782
transform 1 0 19968 0 1 1512
box -48 -56 720 834
use sg13g2_fill_2  FILLER_0_203
timestamp 1677580104
transform 1 0 20640 0 1 1512
box -48 -56 240 834
use sg13g2_decap_8  FILLER_0_321
timestamp 1679581782
transform 1 0 31968 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_328
timestamp 1679581782
transform 1 0 32640 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_335
timestamp 1679581782
transform 1 0 33312 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_342
timestamp 1679581782
transform 1 0 33984 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_349
timestamp 1679581782
transform 1 0 34656 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_356
timestamp 1679581782
transform 1 0 35328 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_363
timestamp 1679581782
transform 1 0 36000 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_370
timestamp 1679581782
transform 1 0 36672 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_377
timestamp 1679581782
transform 1 0 37344 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_384
timestamp 1679581782
transform 1 0 38016 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_391
timestamp 1679581782
transform 1 0 38688 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_398
timestamp 1679581782
transform 1 0 39360 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_405
timestamp 1679581782
transform 1 0 40032 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_412
timestamp 1679581782
transform 1 0 40704 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_419
timestamp 1679581782
transform 1 0 41376 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_426
timestamp 1679581782
transform 1 0 42048 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_433
timestamp 1679581782
transform 1 0 42720 0 1 1512
box -48 -56 720 834
use sg13g2_fill_2  FILLER_0_440
timestamp 1677580104
transform 1 0 43392 0 1 1512
box -48 -56 240 834
use sg13g2_fill_1  FILLER_0_442
timestamp 1677579658
transform 1 0 43584 0 1 1512
box -48 -56 144 834
use sg13g2_decap_8  FILLER_1_0
timestamp 1679581782
transform 1 0 1152 0 -1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_7
timestamp 1679581782
transform 1 0 1824 0 -1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_14
timestamp 1679581782
transform 1 0 2496 0 -1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_21
timestamp 1679581782
transform 1 0 3168 0 -1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_28
timestamp 1679581782
transform 1 0 3840 0 -1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_35
timestamp 1679581782
transform 1 0 4512 0 -1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_42
timestamp 1679581782
transform 1 0 5184 0 -1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_49
timestamp 1679581782
transform 1 0 5856 0 -1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_56
timestamp 1679581782
transform 1 0 6528 0 -1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_63
timestamp 1679581782
transform 1 0 7200 0 -1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_70
timestamp 1679581782
transform 1 0 7872 0 -1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_77
timestamp 1679581782
transform 1 0 8544 0 -1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_84
timestamp 1679581782
transform 1 0 9216 0 -1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_91
timestamp 1679581782
transform 1 0 9888 0 -1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_98
timestamp 1679581782
transform 1 0 10560 0 -1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_105
timestamp 1679581782
transform 1 0 11232 0 -1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_112
timestamp 1679581782
transform 1 0 11904 0 -1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_119
timestamp 1679581782
transform 1 0 12576 0 -1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_126
timestamp 1679581782
transform 1 0 13248 0 -1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_133
timestamp 1679581782
transform 1 0 13920 0 -1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_140
timestamp 1679581782
transform 1 0 14592 0 -1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_147
timestamp 1679581782
transform 1 0 15264 0 -1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_154
timestamp 1679581782
transform 1 0 15936 0 -1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_161
timestamp 1679581782
transform 1 0 16608 0 -1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_168
timestamp 1679581782
transform 1 0 17280 0 -1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_175
timestamp 1679581782
transform 1 0 17952 0 -1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_182
timestamp 1679581782
transform 1 0 18624 0 -1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_189
timestamp 1679581782
transform 1 0 19296 0 -1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_196
timestamp 1679581782
transform 1 0 19968 0 -1 3024
box -48 -56 720 834
use sg13g2_decap_4  FILLER_1_203
timestamp 1679577901
transform 1 0 20640 0 -1 3024
box -48 -56 432 834
use sg13g2_fill_2  FILLER_1_207
timestamp 1677580104
transform 1 0 21024 0 -1 3024
box -48 -56 240 834
use sg13g2_decap_8  FILLER_1_237
timestamp 1679581782
transform 1 0 23904 0 -1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_244
timestamp 1679581782
transform 1 0 24576 0 -1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_315
timestamp 1679581782
transform 1 0 31392 0 -1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_322
timestamp 1679581782
transform 1 0 32064 0 -1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_329
timestamp 1679581782
transform 1 0 32736 0 -1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_336
timestamp 1679581782
transform 1 0 33408 0 -1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_343
timestamp 1679581782
transform 1 0 34080 0 -1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_356
timestamp 1679581782
transform 1 0 35328 0 -1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_363
timestamp 1679581782
transform 1 0 36000 0 -1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_370
timestamp 1679581782
transform 1 0 36672 0 -1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_377
timestamp 1679581782
transform 1 0 37344 0 -1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_384
timestamp 1679581782
transform 1 0 38016 0 -1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_391
timestamp 1679581782
transform 1 0 38688 0 -1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_398
timestamp 1679581782
transform 1 0 39360 0 -1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_405
timestamp 1679581782
transform 1 0 40032 0 -1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_412
timestamp 1679581782
transform 1 0 40704 0 -1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_419
timestamp 1679581782
transform 1 0 41376 0 -1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_426
timestamp 1679581782
transform 1 0 42048 0 -1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_433
timestamp 1679581782
transform 1 0 42720 0 -1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_440
timestamp 1679581782
transform 1 0 43392 0 -1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_0
timestamp 1679581782
transform 1 0 1152 0 1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_7
timestamp 1679581782
transform 1 0 1824 0 1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_14
timestamp 1679581782
transform 1 0 2496 0 1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_21
timestamp 1679581782
transform 1 0 3168 0 1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_28
timestamp 1679581782
transform 1 0 3840 0 1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_35
timestamp 1679581782
transform 1 0 4512 0 1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_42
timestamp 1679581782
transform 1 0 5184 0 1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_49
timestamp 1679581782
transform 1 0 5856 0 1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_56
timestamp 1679581782
transform 1 0 6528 0 1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_63
timestamp 1679581782
transform 1 0 7200 0 1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_70
timestamp 1679581782
transform 1 0 7872 0 1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_77
timestamp 1679581782
transform 1 0 8544 0 1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_84
timestamp 1679581782
transform 1 0 9216 0 1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_91
timestamp 1679581782
transform 1 0 9888 0 1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_98
timestamp 1679581782
transform 1 0 10560 0 1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_105
timestamp 1679581782
transform 1 0 11232 0 1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_112
timestamp 1679581782
transform 1 0 11904 0 1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_119
timestamp 1679581782
transform 1 0 12576 0 1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_126
timestamp 1679581782
transform 1 0 13248 0 1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_133
timestamp 1679581782
transform 1 0 13920 0 1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_140
timestamp 1679581782
transform 1 0 14592 0 1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_147
timestamp 1679581782
transform 1 0 15264 0 1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_154
timestamp 1679581782
transform 1 0 15936 0 1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_161
timestamp 1679581782
transform 1 0 16608 0 1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_168
timestamp 1679581782
transform 1 0 17280 0 1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_175
timestamp 1679581782
transform 1 0 17952 0 1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_182
timestamp 1679581782
transform 1 0 18624 0 1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_189
timestamp 1679581782
transform 1 0 19296 0 1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_196
timestamp 1679581782
transform 1 0 19968 0 1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_203
timestamp 1679581782
transform 1 0 20640 0 1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_210
timestamp 1679581782
transform 1 0 21312 0 1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_217
timestamp 1679581782
transform 1 0 21984 0 1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_224
timestamp 1679581782
transform 1 0 22656 0 1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_231
timestamp 1679581782
transform 1 0 23328 0 1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_238
timestamp 1679581782
transform 1 0 24000 0 1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_245
timestamp 1679581782
transform 1 0 24672 0 1 3024
box -48 -56 720 834
use sg13g2_decap_4  FILLER_2_252
timestamp 1679577901
transform 1 0 25344 0 1 3024
box -48 -56 432 834
use sg13g2_fill_1  FILLER_2_256
timestamp 1677579658
transform 1 0 25728 0 1 3024
box -48 -56 144 834
use sg13g2_decap_8  FILLER_2_285
timestamp 1679581782
transform 1 0 28512 0 1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_292
timestamp 1679581782
transform 1 0 29184 0 1 3024
box -48 -56 720 834
use sg13g2_fill_1  FILLER_2_299
timestamp 1677579658
transform 1 0 29856 0 1 3024
box -48 -56 144 834
use sg13g2_fill_2  FILLER_2_304
timestamp 1677580104
transform 1 0 30336 0 1 3024
box -48 -56 240 834
use sg13g2_fill_1  FILLER_2_306
timestamp 1677579658
transform 1 0 30528 0 1 3024
box -48 -56 144 834
use sg13g2_decap_8  FILLER_2_311
timestamp 1679581782
transform 1 0 31008 0 1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_318
timestamp 1679581782
transform 1 0 31680 0 1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_325
timestamp 1679581782
transform 1 0 32352 0 1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_332
timestamp 1679581782
transform 1 0 33024 0 1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_339
timestamp 1679581782
transform 1 0 33696 0 1 3024
box -48 -56 720 834
use sg13g2_decap_4  FILLER_2_346
timestamp 1679577901
transform 1 0 34368 0 1 3024
box -48 -56 432 834
use sg13g2_decap_8  FILLER_2_354
timestamp 1679581782
transform 1 0 35136 0 1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_361
timestamp 1679581782
transform 1 0 35808 0 1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_372
timestamp 1679581782
transform 1 0 36864 0 1 3024
box -48 -56 720 834
use sg13g2_fill_2  FILLER_2_379
timestamp 1677580104
transform 1 0 37536 0 1 3024
box -48 -56 240 834
use sg13g2_fill_1  FILLER_2_381
timestamp 1677579658
transform 1 0 37728 0 1 3024
box -48 -56 144 834
use sg13g2_decap_8  FILLER_2_386
timestamp 1679581782
transform 1 0 38208 0 1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_393
timestamp 1679581782
transform 1 0 38880 0 1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_400
timestamp 1679581782
transform 1 0 39552 0 1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_407
timestamp 1679581782
transform 1 0 40224 0 1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_414
timestamp 1679581782
transform 1 0 40896 0 1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_421
timestamp 1679581782
transform 1 0 41568 0 1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_428
timestamp 1679581782
transform 1 0 42240 0 1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_435
timestamp 1679581782
transform 1 0 42912 0 1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_442
timestamp 1679581782
transform 1 0 43584 0 1 3024
box -48 -56 720 834
use sg13g2_fill_2  FILLER_2_449
timestamp 1677580104
transform 1 0 44256 0 1 3024
box -48 -56 240 834
use sg13g2_decap_8  FILLER_3_0
timestamp 1679581782
transform 1 0 1152 0 -1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_7
timestamp 1679581782
transform 1 0 1824 0 -1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_14
timestamp 1679581782
transform 1 0 2496 0 -1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_21
timestamp 1679581782
transform 1 0 3168 0 -1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_28
timestamp 1679581782
transform 1 0 3840 0 -1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_35
timestamp 1679581782
transform 1 0 4512 0 -1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_42
timestamp 1679581782
transform 1 0 5184 0 -1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_49
timestamp 1679581782
transform 1 0 5856 0 -1 4536
box -48 -56 720 834
use sg13g2_decap_4  FILLER_3_56
timestamp 1679577901
transform 1 0 6528 0 -1 4536
box -48 -56 432 834
use sg13g2_fill_1  FILLER_3_60
timestamp 1677579658
transform 1 0 6912 0 -1 4536
box -48 -56 144 834
use sg13g2_decap_8  FILLER_3_65
timestamp 1679581782
transform 1 0 7392 0 -1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_72
timestamp 1679581782
transform 1 0 8064 0 -1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_79
timestamp 1679581782
transform 1 0 8736 0 -1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_86
timestamp 1679581782
transform 1 0 9408 0 -1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_93
timestamp 1679581782
transform 1 0 10080 0 -1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_100
timestamp 1679581782
transform 1 0 10752 0 -1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_107
timestamp 1679581782
transform 1 0 11424 0 -1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_114
timestamp 1679581782
transform 1 0 12096 0 -1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_121
timestamp 1679581782
transform 1 0 12768 0 -1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_128
timestamp 1679581782
transform 1 0 13440 0 -1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_135
timestamp 1679581782
transform 1 0 14112 0 -1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_142
timestamp 1679581782
transform 1 0 14784 0 -1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_149
timestamp 1679581782
transform 1 0 15456 0 -1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_156
timestamp 1679581782
transform 1 0 16128 0 -1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_163
timestamp 1679581782
transform 1 0 16800 0 -1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_170
timestamp 1679581782
transform 1 0 17472 0 -1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_177
timestamp 1679581782
transform 1 0 18144 0 -1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_184
timestamp 1679581782
transform 1 0 18816 0 -1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_191
timestamp 1679581782
transform 1 0 19488 0 -1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_198
timestamp 1679581782
transform 1 0 20160 0 -1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_205
timestamp 1679581782
transform 1 0 20832 0 -1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_212
timestamp 1679581782
transform 1 0 21504 0 -1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_219
timestamp 1679581782
transform 1 0 22176 0 -1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_226
timestamp 1679581782
transform 1 0 22848 0 -1 4536
box -48 -56 720 834
use sg13g2_decap_4  FILLER_3_233
timestamp 1679577901
transform 1 0 23520 0 -1 4536
box -48 -56 432 834
use sg13g2_fill_1  FILLER_3_241
timestamp 1677579658
transform 1 0 24288 0 -1 4536
box -48 -56 144 834
use sg13g2_decap_4  FILLER_3_246
timestamp 1679577901
transform 1 0 24768 0 -1 4536
box -48 -56 432 834
use sg13g2_fill_1  FILLER_3_250
timestamp 1677579658
transform 1 0 25152 0 -1 4536
box -48 -56 144 834
use sg13g2_decap_4  FILLER_3_255
timestamp 1679577901
transform 1 0 25632 0 -1 4536
box -48 -56 432 834
use sg13g2_fill_1  FILLER_3_259
timestamp 1677579658
transform 1 0 26016 0 -1 4536
box -48 -56 144 834
use sg13g2_decap_8  FILLER_3_264
timestamp 1679581782
transform 1 0 26496 0 -1 4536
box -48 -56 720 834
use sg13g2_decap_4  FILLER_3_271
timestamp 1679577901
transform 1 0 27168 0 -1 4536
box -48 -56 432 834
use sg13g2_decap_8  FILLER_3_279
timestamp 1679581782
transform 1 0 27936 0 -1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_286
timestamp 1679581782
transform 1 0 28608 0 -1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_293
timestamp 1679581782
transform 1 0 29280 0 -1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_300
timestamp 1679581782
transform 1 0 29952 0 -1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_307
timestamp 1679581782
transform 1 0 30624 0 -1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_314
timestamp 1679581782
transform 1 0 31296 0 -1 4536
box -48 -56 720 834
use sg13g2_decap_4  FILLER_3_321
timestamp 1679577901
transform 1 0 31968 0 -1 4536
box -48 -56 432 834
use sg13g2_fill_2  FILLER_3_325
timestamp 1677580104
transform 1 0 32352 0 -1 4536
box -48 -56 240 834
use sg13g2_decap_8  FILLER_3_331
timestamp 1679581782
transform 1 0 32928 0 -1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_338
timestamp 1679581782
transform 1 0 33600 0 -1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_345
timestamp 1679581782
transform 1 0 34272 0 -1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_352
timestamp 1679581782
transform 1 0 34944 0 -1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_359
timestamp 1679581782
transform 1 0 35616 0 -1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_366
timestamp 1679581782
transform 1 0 36288 0 -1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_373
timestamp 1679581782
transform 1 0 36960 0 -1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_380
timestamp 1679581782
transform 1 0 37632 0 -1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_387
timestamp 1679581782
transform 1 0 38304 0 -1 4536
box -48 -56 720 834
use sg13g2_fill_2  FILLER_3_394
timestamp 1677580104
transform 1 0 38976 0 -1 4536
box -48 -56 240 834
use sg13g2_fill_1  FILLER_3_396
timestamp 1677579658
transform 1 0 39168 0 -1 4536
box -48 -56 144 834
use sg13g2_decap_4  FILLER_3_400
timestamp 1679577901
transform 1 0 39552 0 -1 4536
box -48 -56 432 834
use sg13g2_fill_2  FILLER_3_407
timestamp 1677580104
transform 1 0 40224 0 -1 4536
box -48 -56 240 834
use sg13g2_decap_8  FILLER_3_436
timestamp 1679581782
transform 1 0 43008 0 -1 4536
box -48 -56 720 834
use sg13g2_decap_4  FILLER_3_443
timestamp 1679577901
transform 1 0 43680 0 -1 4536
box -48 -56 432 834
use sg13g2_decap_8  FILLER_4_0
timestamp 1679581782
transform 1 0 1152 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_7
timestamp 1679581782
transform 1 0 1824 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_14
timestamp 1679581782
transform 1 0 2496 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_21
timestamp 1679581782
transform 1 0 3168 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_28
timestamp 1679581782
transform 1 0 3840 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_35
timestamp 1679581782
transform 1 0 4512 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_42
timestamp 1679581782
transform 1 0 5184 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_49
timestamp 1679581782
transform 1 0 5856 0 1 4536
box -48 -56 720 834
use sg13g2_decap_4  FILLER_4_56
timestamp 1679577901
transform 1 0 6528 0 1 4536
box -48 -56 432 834
use sg13g2_fill_2  FILLER_4_60
timestamp 1677580104
transform 1 0 6912 0 1 4536
box -48 -56 240 834
use sg13g2_decap_4  FILLER_4_70
timestamp 1679577901
transform 1 0 7872 0 1 4536
box -48 -56 432 834
use sg13g2_decap_8  FILLER_4_78
timestamp 1679581782
transform 1 0 8640 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_85
timestamp 1679581782
transform 1 0 9312 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_92
timestamp 1679581782
transform 1 0 9984 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_99
timestamp 1679581782
transform 1 0 10656 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_106
timestamp 1679581782
transform 1 0 11328 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_113
timestamp 1679581782
transform 1 0 12000 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_120
timestamp 1679581782
transform 1 0 12672 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_127
timestamp 1679581782
transform 1 0 13344 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_134
timestamp 1679581782
transform 1 0 14016 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_141
timestamp 1679581782
transform 1 0 14688 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_148
timestamp 1679581782
transform 1 0 15360 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_155
timestamp 1679581782
transform 1 0 16032 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_162
timestamp 1679581782
transform 1 0 16704 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_169
timestamp 1679581782
transform 1 0 17376 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_176
timestamp 1679581782
transform 1 0 18048 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_183
timestamp 1679581782
transform 1 0 18720 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_190
timestamp 1679581782
transform 1 0 19392 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_197
timestamp 1679581782
transform 1 0 20064 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_204
timestamp 1679581782
transform 1 0 20736 0 1 4536
box -48 -56 720 834
use sg13g2_decap_4  FILLER_4_211
timestamp 1679577901
transform 1 0 21408 0 1 4536
box -48 -56 432 834
use sg13g2_fill_2  FILLER_4_215
timestamp 1677580104
transform 1 0 21792 0 1 4536
box -48 -56 240 834
use sg13g2_fill_1  FILLER_4_225
timestamp 1677579658
transform 1 0 22752 0 1 4536
box -48 -56 144 834
use sg13g2_fill_1  FILLER_4_230
timestamp 1677579658
transform 1 0 23232 0 1 4536
box -48 -56 144 834
use sg13g2_decap_8  FILLER_4_235
timestamp 1679581782
transform 1 0 23712 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_242
timestamp 1679581782
transform 1 0 24384 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_249
timestamp 1679581782
transform 1 0 25056 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_256
timestamp 1679581782
transform 1 0 25728 0 1 4536
box -48 -56 720 834
use sg13g2_decap_4  FILLER_4_263
timestamp 1679577901
transform 1 0 26400 0 1 4536
box -48 -56 432 834
use sg13g2_decap_4  FILLER_4_271
timestamp 1679577901
transform 1 0 27168 0 1 4536
box -48 -56 432 834
use sg13g2_fill_1  FILLER_4_275
timestamp 1677579658
transform 1 0 27552 0 1 4536
box -48 -56 144 834
use sg13g2_decap_8  FILLER_4_288
timestamp 1679581782
transform 1 0 28800 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_295
timestamp 1679581782
transform 1 0 29472 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_302
timestamp 1679581782
transform 1 0 30144 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_309
timestamp 1679581782
transform 1 0 30816 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_316
timestamp 1679581782
transform 1 0 31488 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_323
timestamp 1679581782
transform 1 0 32160 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_330
timestamp 1679581782
transform 1 0 32832 0 1 4536
box -48 -56 720 834
use sg13g2_decap_4  FILLER_4_337
timestamp 1679577901
transform 1 0 33504 0 1 4536
box -48 -56 432 834
use sg13g2_fill_2  FILLER_4_341
timestamp 1677580104
transform 1 0 33888 0 1 4536
box -48 -56 240 834
use sg13g2_decap_8  FILLER_4_349
timestamp 1679581782
transform 1 0 34656 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_356
timestamp 1679581782
transform 1 0 35328 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_363
timestamp 1679581782
transform 1 0 36000 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_370
timestamp 1679581782
transform 1 0 36672 0 1 4536
box -48 -56 720 834
use sg13g2_fill_2  FILLER_4_377
timestamp 1677580104
transform 1 0 37344 0 1 4536
box -48 -56 240 834
use sg13g2_fill_1  FILLER_4_379
timestamp 1677579658
transform 1 0 37536 0 1 4536
box -48 -56 144 834
use sg13g2_decap_4  FILLER_4_383
timestamp 1679577901
transform 1 0 37920 0 1 4536
box -48 -56 432 834
use sg13g2_fill_1  FILLER_4_404
timestamp 1677579658
transform 1 0 39936 0 1 4536
box -48 -56 144 834
use sg13g2_fill_1  FILLER_4_408
timestamp 1677579658
transform 1 0 40320 0 1 4536
box -48 -56 144 834
use sg13g2_decap_8  FILLER_4_426
timestamp 1679581782
transform 1 0 42048 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_433
timestamp 1679581782
transform 1 0 42720 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_440
timestamp 1679581782
transform 1 0 43392 0 1 4536
box -48 -56 720 834
use sg13g2_decap_4  FILLER_4_447
timestamp 1679577901
transform 1 0 44064 0 1 4536
box -48 -56 432 834
use sg13g2_decap_8  FILLER_5_0
timestamp 1679581782
transform 1 0 1152 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_7
timestamp 1679581782
transform 1 0 1824 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_14
timestamp 1679581782
transform 1 0 2496 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_21
timestamp 1679581782
transform 1 0 3168 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_28
timestamp 1679581782
transform 1 0 3840 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_35
timestamp 1679581782
transform 1 0 4512 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_42
timestamp 1679581782
transform 1 0 5184 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_49
timestamp 1679581782
transform 1 0 5856 0 -1 6048
box -48 -56 720 834
use sg13g2_fill_1  FILLER_5_56
timestamp 1677579658
transform 1 0 6528 0 -1 6048
box -48 -56 144 834
use sg13g2_decap_4  FILLER_5_61
timestamp 1679577901
transform 1 0 7008 0 -1 6048
box -48 -56 432 834
use sg13g2_fill_1  FILLER_5_65
timestamp 1677579658
transform 1 0 7392 0 -1 6048
box -48 -56 144 834
use sg13g2_decap_8  FILLER_5_70
timestamp 1679581782
transform 1 0 7872 0 -1 6048
box -48 -56 720 834
use sg13g2_fill_1  FILLER_5_77
timestamp 1677579658
transform 1 0 8544 0 -1 6048
box -48 -56 144 834
use sg13g2_decap_8  FILLER_5_82
timestamp 1679581782
transform 1 0 9024 0 -1 6048
box -48 -56 720 834
use sg13g2_fill_1  FILLER_5_89
timestamp 1677579658
transform 1 0 9696 0 -1 6048
box -48 -56 144 834
use sg13g2_decap_4  FILLER_5_94
timestamp 1679577901
transform 1 0 10176 0 -1 6048
box -48 -56 432 834
use sg13g2_fill_2  FILLER_5_98
timestamp 1677580104
transform 1 0 10560 0 -1 6048
box -48 -56 240 834
use sg13g2_fill_2  FILLER_5_104
timestamp 1677580104
transform 1 0 11136 0 -1 6048
box -48 -56 240 834
use sg13g2_fill_1  FILLER_5_106
timestamp 1677579658
transform 1 0 11328 0 -1 6048
box -48 -56 144 834
use sg13g2_decap_4  FILLER_5_111
timestamp 1679577901
transform 1 0 11808 0 -1 6048
box -48 -56 432 834
use sg13g2_decap_8  FILLER_5_119
timestamp 1679581782
transform 1 0 12576 0 -1 6048
box -48 -56 720 834
use sg13g2_fill_2  FILLER_5_126
timestamp 1677580104
transform 1 0 13248 0 -1 6048
box -48 -56 240 834
use sg13g2_decap_8  FILLER_5_132
timestamp 1679581782
transform 1 0 13824 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_139
timestamp 1679581782
transform 1 0 14496 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_146
timestamp 1679581782
transform 1 0 15168 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_153
timestamp 1679581782
transform 1 0 15840 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_160
timestamp 1679581782
transform 1 0 16512 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_167
timestamp 1679581782
transform 1 0 17184 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_174
timestamp 1679581782
transform 1 0 17856 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_181
timestamp 1679581782
transform 1 0 18528 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_188
timestamp 1679581782
transform 1 0 19200 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_195
timestamp 1679581782
transform 1 0 19872 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_4  FILLER_5_202
timestamp 1679577901
transform 1 0 20544 0 -1 6048
box -48 -56 432 834
use sg13g2_decap_8  FILLER_5_218
timestamp 1679581782
transform 1 0 22080 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_225
timestamp 1679581782
transform 1 0 22752 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_232
timestamp 1679581782
transform 1 0 23424 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_239
timestamp 1679581782
transform 1 0 24096 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_246
timestamp 1679581782
transform 1 0 24768 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_253
timestamp 1679581782
transform 1 0 25440 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_260
timestamp 1679581782
transform 1 0 26112 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_267
timestamp 1679581782
transform 1 0 26784 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_274
timestamp 1679581782
transform 1 0 27456 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_281
timestamp 1679581782
transform 1 0 28128 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_288
timestamp 1679581782
transform 1 0 28800 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_295
timestamp 1679581782
transform 1 0 29472 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_302
timestamp 1679581782
transform 1 0 30144 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_309
timestamp 1679581782
transform 1 0 30816 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_316
timestamp 1679581782
transform 1 0 31488 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_323
timestamp 1679581782
transform 1 0 32160 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_330
timestamp 1679581782
transform 1 0 32832 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_4  FILLER_5_337
timestamp 1679577901
transform 1 0 33504 0 -1 6048
box -48 -56 432 834
use sg13g2_fill_2  FILLER_5_341
timestamp 1677580104
transform 1 0 33888 0 -1 6048
box -48 -56 240 834
use sg13g2_decap_8  FILLER_5_347
timestamp 1679581782
transform 1 0 34464 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_354
timestamp 1679581782
transform 1 0 35136 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_361
timestamp 1679581782
transform 1 0 35808 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_4  FILLER_5_368
timestamp 1679577901
transform 1 0 36480 0 -1 6048
box -48 -56 432 834
use sg13g2_fill_1  FILLER_5_376
timestamp 1677579658
transform 1 0 37248 0 -1 6048
box -48 -56 144 834
use sg13g2_fill_1  FILLER_5_380
timestamp 1677579658
transform 1 0 37632 0 -1 6048
box -48 -56 144 834
use sg13g2_decap_8  FILLER_5_392
timestamp 1679581782
transform 1 0 38784 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_399
timestamp 1679581782
transform 1 0 39456 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_406
timestamp 1679581782
transform 1 0 40128 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_413
timestamp 1679581782
transform 1 0 40800 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_420
timestamp 1679581782
transform 1 0 41472 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_427
timestamp 1679581782
transform 1 0 42144 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_434
timestamp 1679581782
transform 1 0 42816 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_441
timestamp 1679581782
transform 1 0 43488 0 -1 6048
box -48 -56 720 834
use sg13g2_fill_2  FILLER_5_448
timestamp 1677580104
transform 1 0 44160 0 -1 6048
box -48 -56 240 834
use sg13g2_fill_1  FILLER_5_450
timestamp 1677579658
transform 1 0 44352 0 -1 6048
box -48 -56 144 834
use sg13g2_decap_8  FILLER_6_0
timestamp 1679581782
transform 1 0 1152 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_7
timestamp 1679581782
transform 1 0 1824 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_14
timestamp 1679581782
transform 1 0 2496 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_21
timestamp 1679581782
transform 1 0 3168 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_28
timestamp 1679581782
transform 1 0 3840 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_35
timestamp 1679581782
transform 1 0 4512 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_42
timestamp 1679581782
transform 1 0 5184 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_49
timestamp 1679581782
transform 1 0 5856 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_56
timestamp 1679581782
transform 1 0 6528 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_63
timestamp 1679581782
transform 1 0 7200 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_70
timestamp 1679581782
transform 1 0 7872 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_77
timestamp 1679581782
transform 1 0 8544 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_84
timestamp 1679581782
transform 1 0 9216 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_91
timestamp 1679581782
transform 1 0 9888 0 1 6048
box -48 -56 720 834
use sg13g2_fill_2  FILLER_6_98
timestamp 1677580104
transform 1 0 10560 0 1 6048
box -48 -56 240 834
use sg13g2_decap_8  FILLER_6_104
timestamp 1679581782
transform 1 0 11136 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_111
timestamp 1679581782
transform 1 0 11808 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_118
timestamp 1679581782
transform 1 0 12480 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_125
timestamp 1679581782
transform 1 0 13152 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_132
timestamp 1679581782
transform 1 0 13824 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_139
timestamp 1679581782
transform 1 0 14496 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_146
timestamp 1679581782
transform 1 0 15168 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_153
timestamp 1679581782
transform 1 0 15840 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_160
timestamp 1679581782
transform 1 0 16512 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_167
timestamp 1679581782
transform 1 0 17184 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_174
timestamp 1679581782
transform 1 0 17856 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_181
timestamp 1679581782
transform 1 0 18528 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_188
timestamp 1679581782
transform 1 0 19200 0 1 6048
box -48 -56 720 834
use sg13g2_fill_1  FILLER_6_199
timestamp 1677579658
transform 1 0 20256 0 1 6048
box -48 -56 144 834
use sg13g2_decap_8  FILLER_6_204
timestamp 1679581782
transform 1 0 20736 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_211
timestamp 1679581782
transform 1 0 21408 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_218
timestamp 1679581782
transform 1 0 22080 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_225
timestamp 1679581782
transform 1 0 22752 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_232
timestamp 1679581782
transform 1 0 23424 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_239
timestamp 1679581782
transform 1 0 24096 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_246
timestamp 1679581782
transform 1 0 24768 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_253
timestamp 1679581782
transform 1 0 25440 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_260
timestamp 1679581782
transform 1 0 26112 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_267
timestamp 1679581782
transform 1 0 26784 0 1 6048
box -48 -56 720 834
use sg13g2_decap_4  FILLER_6_274
timestamp 1679577901
transform 1 0 27456 0 1 6048
box -48 -56 432 834
use sg13g2_fill_2  FILLER_6_278
timestamp 1677580104
transform 1 0 27840 0 1 6048
box -48 -56 240 834
use sg13g2_decap_8  FILLER_6_284
timestamp 1679581782
transform 1 0 28416 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_291
timestamp 1679581782
transform 1 0 29088 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_298
timestamp 1679581782
transform 1 0 29760 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_305
timestamp 1679581782
transform 1 0 30432 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_312
timestamp 1679581782
transform 1 0 31104 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_319
timestamp 1679581782
transform 1 0 31776 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_326
timestamp 1679581782
transform 1 0 32448 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_337
timestamp 1679581782
transform 1 0 33504 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_344
timestamp 1679581782
transform 1 0 34176 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_351
timestamp 1679581782
transform 1 0 34848 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_358
timestamp 1679581782
transform 1 0 35520 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_365
timestamp 1679581782
transform 1 0 36192 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_372
timestamp 1679581782
transform 1 0 36864 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_379
timestamp 1679581782
transform 1 0 37536 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_386
timestamp 1679581782
transform 1 0 38208 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_393
timestamp 1679581782
transform 1 0 38880 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_400
timestamp 1679581782
transform 1 0 39552 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_407
timestamp 1679581782
transform 1 0 40224 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_414
timestamp 1679581782
transform 1 0 40896 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_421
timestamp 1679581782
transform 1 0 41568 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_428
timestamp 1679581782
transform 1 0 42240 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_435
timestamp 1679581782
transform 1 0 42912 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_442
timestamp 1679581782
transform 1 0 43584 0 1 6048
box -48 -56 720 834
use sg13g2_fill_2  FILLER_6_449
timestamp 1677580104
transform 1 0 44256 0 1 6048
box -48 -56 240 834
use sg13g2_decap_8  FILLER_7_0
timestamp 1679581782
transform 1 0 1152 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_7
timestamp 1679581782
transform 1 0 1824 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_14
timestamp 1679581782
transform 1 0 2496 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_21
timestamp 1679581782
transform 1 0 3168 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_28
timestamp 1679581782
transform 1 0 3840 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_35
timestamp 1679581782
transform 1 0 4512 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_42
timestamp 1679581782
transform 1 0 5184 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_49
timestamp 1679581782
transform 1 0 5856 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_56
timestamp 1679581782
transform 1 0 6528 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_63
timestamp 1679581782
transform 1 0 7200 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_70
timestamp 1679581782
transform 1 0 7872 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_77
timestamp 1679581782
transform 1 0 8544 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_84
timestamp 1679581782
transform 1 0 9216 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_91
timestamp 1679581782
transform 1 0 9888 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_98
timestamp 1679581782
transform 1 0 10560 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_105
timestamp 1679581782
transform 1 0 11232 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_4  FILLER_7_112
timestamp 1679577901
transform 1 0 11904 0 -1 7560
box -48 -56 432 834
use sg13g2_fill_1  FILLER_7_116
timestamp 1677579658
transform 1 0 12288 0 -1 7560
box -48 -56 144 834
use sg13g2_decap_8  FILLER_7_121
timestamp 1679581782
transform 1 0 12768 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_4  FILLER_7_128
timestamp 1679577901
transform 1 0 13440 0 -1 7560
box -48 -56 432 834
use sg13g2_decap_8  FILLER_7_136
timestamp 1679581782
transform 1 0 14208 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_147
timestamp 1679581782
transform 1 0 15264 0 -1 7560
box -48 -56 720 834
use sg13g2_fill_1  FILLER_7_154
timestamp 1677579658
transform 1 0 15936 0 -1 7560
box -48 -56 144 834
use sg13g2_decap_4  FILLER_7_159
timestamp 1679577901
transform 1 0 16416 0 -1 7560
box -48 -56 432 834
use sg13g2_fill_1  FILLER_7_167
timestamp 1677579658
transform 1 0 17184 0 -1 7560
box -48 -56 144 834
use sg13g2_decap_8  FILLER_7_212
timestamp 1679581782
transform 1 0 21504 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_219
timestamp 1679581782
transform 1 0 22176 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_226
timestamp 1679581782
transform 1 0 22848 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_233
timestamp 1679581782
transform 1 0 23520 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_240
timestamp 1679581782
transform 1 0 24192 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_247
timestamp 1679581782
transform 1 0 24864 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_254
timestamp 1679581782
transform 1 0 25536 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_261
timestamp 1679581782
transform 1 0 26208 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_268
timestamp 1679581782
transform 1 0 26880 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_275
timestamp 1679581782
transform 1 0 27552 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_282
timestamp 1679581782
transform 1 0 28224 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_289
timestamp 1679581782
transform 1 0 28896 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_296
timestamp 1679581782
transform 1 0 29568 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_303
timestamp 1679581782
transform 1 0 30240 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_310
timestamp 1679581782
transform 1 0 30912 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_317
timestamp 1679581782
transform 1 0 31584 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_324
timestamp 1679581782
transform 1 0 32256 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_331
timestamp 1679581782
transform 1 0 32928 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_338
timestamp 1679581782
transform 1 0 33600 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_345
timestamp 1679581782
transform 1 0 34272 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_352
timestamp 1679581782
transform 1 0 34944 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_359
timestamp 1679581782
transform 1 0 35616 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_366
timestamp 1679581782
transform 1 0 36288 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_373
timestamp 1679581782
transform 1 0 36960 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_380
timestamp 1679581782
transform 1 0 37632 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_387
timestamp 1679581782
transform 1 0 38304 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_394
timestamp 1679581782
transform 1 0 38976 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_401
timestamp 1679581782
transform 1 0 39648 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_408
timestamp 1679581782
transform 1 0 40320 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_415
timestamp 1679581782
transform 1 0 40992 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_422
timestamp 1679581782
transform 1 0 41664 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_429
timestamp 1679581782
transform 1 0 42336 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_436
timestamp 1679581782
transform 1 0 43008 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_443
timestamp 1679581782
transform 1 0 43680 0 -1 7560
box -48 -56 720 834
use sg13g2_fill_1  FILLER_7_450
timestamp 1677579658
transform 1 0 44352 0 -1 7560
box -48 -56 144 834
use sg13g2_decap_8  FILLER_8_0
timestamp 1679581782
transform 1 0 1152 0 1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_7
timestamp 1679581782
transform 1 0 1824 0 1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_14
timestamp 1679581782
transform 1 0 2496 0 1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_21
timestamp 1679581782
transform 1 0 3168 0 1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_28
timestamp 1679581782
transform 1 0 3840 0 1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_35
timestamp 1679581782
transform 1 0 4512 0 1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_42
timestamp 1679581782
transform 1 0 5184 0 1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_49
timestamp 1679581782
transform 1 0 5856 0 1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_56
timestamp 1679581782
transform 1 0 6528 0 1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_63
timestamp 1679581782
transform 1 0 7200 0 1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_70
timestamp 1679581782
transform 1 0 7872 0 1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_77
timestamp 1679581782
transform 1 0 8544 0 1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_84
timestamp 1679581782
transform 1 0 9216 0 1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_91
timestamp 1679581782
transform 1 0 9888 0 1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_98
timestamp 1679581782
transform 1 0 10560 0 1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_105
timestamp 1679581782
transform 1 0 11232 0 1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_112
timestamp 1679581782
transform 1 0 11904 0 1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_119
timestamp 1679581782
transform 1 0 12576 0 1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_126
timestamp 1679581782
transform 1 0 13248 0 1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_133
timestamp 1679581782
transform 1 0 13920 0 1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_140
timestamp 1679581782
transform 1 0 14592 0 1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_147
timestamp 1679581782
transform 1 0 15264 0 1 7560
box -48 -56 720 834
use sg13g2_fill_2  FILLER_8_154
timestamp 1677580104
transform 1 0 15936 0 1 7560
box -48 -56 240 834
use sg13g2_fill_2  FILLER_8_176
timestamp 1677580104
transform 1 0 18048 0 1 7560
box -48 -56 240 834
use sg13g2_fill_1  FILLER_8_178
timestamp 1677579658
transform 1 0 18240 0 1 7560
box -48 -56 144 834
use sg13g2_decap_8  FILLER_8_187
timestamp 1679581782
transform 1 0 19104 0 1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_194
timestamp 1679581782
transform 1 0 19776 0 1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_201
timestamp 1679581782
transform 1 0 20448 0 1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_208
timestamp 1679581782
transform 1 0 21120 0 1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_215
timestamp 1679581782
transform 1 0 21792 0 1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_222
timestamp 1679581782
transform 1 0 22464 0 1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_229
timestamp 1679581782
transform 1 0 23136 0 1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_236
timestamp 1679581782
transform 1 0 23808 0 1 7560
box -48 -56 720 834
use sg13g2_fill_2  FILLER_8_243
timestamp 1677580104
transform 1 0 24480 0 1 7560
box -48 -56 240 834
use sg13g2_fill_2  FILLER_8_249
timestamp 1677580104
transform 1 0 25056 0 1 7560
box -48 -56 240 834
use sg13g2_fill_1  FILLER_8_251
timestamp 1677579658
transform 1 0 25248 0 1 7560
box -48 -56 144 834
use sg13g2_decap_4  FILLER_8_256
timestamp 1679577901
transform 1 0 25728 0 1 7560
box -48 -56 432 834
use sg13g2_fill_1  FILLER_8_260
timestamp 1677579658
transform 1 0 26112 0 1 7560
box -48 -56 144 834
use sg13g2_decap_8  FILLER_8_265
timestamp 1679581782
transform 1 0 26592 0 1 7560
box -48 -56 720 834
use sg13g2_decap_4  FILLER_8_272
timestamp 1679577901
transform 1 0 27264 0 1 7560
box -48 -56 432 834
use sg13g2_fill_1  FILLER_8_276
timestamp 1677579658
transform 1 0 27648 0 1 7560
box -48 -56 144 834
use sg13g2_decap_4  FILLER_8_281
timestamp 1679577901
transform 1 0 28128 0 1 7560
box -48 -56 432 834
use sg13g2_decap_8  FILLER_8_289
timestamp 1679581782
transform 1 0 28896 0 1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_296
timestamp 1679581782
transform 1 0 29568 0 1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_303
timestamp 1679581782
transform 1 0 30240 0 1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_310
timestamp 1679581782
transform 1 0 30912 0 1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_317
timestamp 1679581782
transform 1 0 31584 0 1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_324
timestamp 1679581782
transform 1 0 32256 0 1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_331
timestamp 1679581782
transform 1 0 32928 0 1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_338
timestamp 1679581782
transform 1 0 33600 0 1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_345
timestamp 1679581782
transform 1 0 34272 0 1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_352
timestamp 1679581782
transform 1 0 34944 0 1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_359
timestamp 1679581782
transform 1 0 35616 0 1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_366
timestamp 1679581782
transform 1 0 36288 0 1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_373
timestamp 1679581782
transform 1 0 36960 0 1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_380
timestamp 1679581782
transform 1 0 37632 0 1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_387
timestamp 1679581782
transform 1 0 38304 0 1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_394
timestamp 1679581782
transform 1 0 38976 0 1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_401
timestamp 1679581782
transform 1 0 39648 0 1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_408
timestamp 1679581782
transform 1 0 40320 0 1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_415
timestamp 1679581782
transform 1 0 40992 0 1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_422
timestamp 1679581782
transform 1 0 41664 0 1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_429
timestamp 1679581782
transform 1 0 42336 0 1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_436
timestamp 1679581782
transform 1 0 43008 0 1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_443
timestamp 1679581782
transform 1 0 43680 0 1 7560
box -48 -56 720 834
use sg13g2_fill_1  FILLER_8_450
timestamp 1677579658
transform 1 0 44352 0 1 7560
box -48 -56 144 834
use sg13g2_decap_8  FILLER_9_0
timestamp 1679581782
transform 1 0 1152 0 -1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_7
timestamp 1679581782
transform 1 0 1824 0 -1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_14
timestamp 1679581782
transform 1 0 2496 0 -1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_21
timestamp 1679581782
transform 1 0 3168 0 -1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_28
timestamp 1679581782
transform 1 0 3840 0 -1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_35
timestamp 1679581782
transform 1 0 4512 0 -1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_42
timestamp 1679581782
transform 1 0 5184 0 -1 9072
box -48 -56 720 834
use sg13g2_fill_2  FILLER_9_49
timestamp 1677580104
transform 1 0 5856 0 -1 9072
box -48 -56 240 834
use sg13g2_fill_1  FILLER_9_51
timestamp 1677579658
transform 1 0 6048 0 -1 9072
box -48 -56 144 834
use sg13g2_fill_1  FILLER_9_56
timestamp 1677579658
transform 1 0 6528 0 -1 9072
box -48 -56 144 834
use sg13g2_decap_4  FILLER_9_61
timestamp 1679577901
transform 1 0 7008 0 -1 9072
box -48 -56 432 834
use sg13g2_decap_8  FILLER_9_69
timestamp 1679581782
transform 1 0 7776 0 -1 9072
box -48 -56 720 834
use sg13g2_fill_1  FILLER_9_76
timestamp 1677579658
transform 1 0 8448 0 -1 9072
box -48 -56 144 834
use sg13g2_decap_8  FILLER_9_81
timestamp 1679581782
transform 1 0 8928 0 -1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_88
timestamp 1679581782
transform 1 0 9600 0 -1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_95
timestamp 1679581782
transform 1 0 10272 0 -1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_102
timestamp 1679581782
transform 1 0 10944 0 -1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_109
timestamp 1679581782
transform 1 0 11616 0 -1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_116
timestamp 1679581782
transform 1 0 12288 0 -1 9072
box -48 -56 720 834
use sg13g2_fill_1  FILLER_9_123
timestamp 1677579658
transform 1 0 12960 0 -1 9072
box -48 -56 144 834
use sg13g2_decap_8  FILLER_9_128
timestamp 1679581782
transform 1 0 13440 0 -1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_135
timestamp 1679581782
transform 1 0 14112 0 -1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_142
timestamp 1679581782
transform 1 0 14784 0 -1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_149
timestamp 1679581782
transform 1 0 15456 0 -1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_156
timestamp 1679581782
transform 1 0 16128 0 -1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_163
timestamp 1679581782
transform 1 0 16800 0 -1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_170
timestamp 1679581782
transform 1 0 17472 0 -1 9072
box -48 -56 720 834
use sg13g2_decap_4  FILLER_9_177
timestamp 1679577901
transform 1 0 18144 0 -1 9072
box -48 -56 432 834
use sg13g2_fill_2  FILLER_9_181
timestamp 1677580104
transform 1 0 18528 0 -1 9072
box -48 -56 240 834
use sg13g2_decap_8  FILLER_9_187
timestamp 1679581782
transform 1 0 19104 0 -1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_194
timestamp 1679581782
transform 1 0 19776 0 -1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_201
timestamp 1679581782
transform 1 0 20448 0 -1 9072
box -48 -56 720 834
use sg13g2_fill_1  FILLER_9_208
timestamp 1677579658
transform 1 0 21120 0 -1 9072
box -48 -56 144 834
use sg13g2_fill_2  FILLER_9_237
timestamp 1677580104
transform 1 0 23904 0 -1 9072
box -48 -56 240 834
use sg13g2_decap_8  FILLER_9_243
timestamp 1679581782
transform 1 0 24480 0 -1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_250
timestamp 1679581782
transform 1 0 25152 0 -1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_261
timestamp 1679581782
transform 1 0 26208 0 -1 9072
box -48 -56 720 834
use sg13g2_fill_2  FILLER_9_288
timestamp 1677580104
transform 1 0 28800 0 -1 9072
box -48 -56 240 834
use sg13g2_fill_1  FILLER_9_290
timestamp 1677579658
transform 1 0 28992 0 -1 9072
box -48 -56 144 834
use sg13g2_decap_8  FILLER_9_295
timestamp 1679581782
transform 1 0 29472 0 -1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_302
timestamp 1679581782
transform 1 0 30144 0 -1 9072
box -48 -56 720 834
use sg13g2_decap_4  FILLER_9_309
timestamp 1679577901
transform 1 0 30816 0 -1 9072
box -48 -56 432 834
use sg13g2_decap_8  FILLER_9_321
timestamp 1679581782
transform 1 0 31968 0 -1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_328
timestamp 1679581782
transform 1 0 32640 0 -1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_335
timestamp 1679581782
transform 1 0 33312 0 -1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_342
timestamp 1679581782
transform 1 0 33984 0 -1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_349
timestamp 1679581782
transform 1 0 34656 0 -1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_356
timestamp 1679581782
transform 1 0 35328 0 -1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_363
timestamp 1679581782
transform 1 0 36000 0 -1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_370
timestamp 1679581782
transform 1 0 36672 0 -1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_377
timestamp 1679581782
transform 1 0 37344 0 -1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_384
timestamp 1679581782
transform 1 0 38016 0 -1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_391
timestamp 1679581782
transform 1 0 38688 0 -1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_398
timestamp 1679581782
transform 1 0 39360 0 -1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_405
timestamp 1679581782
transform 1 0 40032 0 -1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_412
timestamp 1679581782
transform 1 0 40704 0 -1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_419
timestamp 1679581782
transform 1 0 41376 0 -1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_426
timestamp 1679581782
transform 1 0 42048 0 -1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_433
timestamp 1679581782
transform 1 0 42720 0 -1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_440
timestamp 1679581782
transform 1 0 43392 0 -1 9072
box -48 -56 720 834
use sg13g2_decap_4  FILLER_9_447
timestamp 1679577901
transform 1 0 44064 0 -1 9072
box -48 -56 432 834
use sg13g2_decap_8  FILLER_10_0
timestamp 1679581782
transform 1 0 1152 0 1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_7
timestamp 1679581782
transform 1 0 1824 0 1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_14
timestamp 1679581782
transform 1 0 2496 0 1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_21
timestamp 1679581782
transform 1 0 3168 0 1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_28
timestamp 1679581782
transform 1 0 3840 0 1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_35
timestamp 1679581782
transform 1 0 4512 0 1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_42
timestamp 1679581782
transform 1 0 5184 0 1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_49
timestamp 1679581782
transform 1 0 5856 0 1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_56
timestamp 1679581782
transform 1 0 6528 0 1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_63
timestamp 1679581782
transform 1 0 7200 0 1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_70
timestamp 1679581782
transform 1 0 7872 0 1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_77
timestamp 1679581782
transform 1 0 8544 0 1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_84
timestamp 1679581782
transform 1 0 9216 0 1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_91
timestamp 1679581782
transform 1 0 9888 0 1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_98
timestamp 1679581782
transform 1 0 10560 0 1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_105
timestamp 1679581782
transform 1 0 11232 0 1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_112
timestamp 1679581782
transform 1 0 11904 0 1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_119
timestamp 1679581782
transform 1 0 12576 0 1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_126
timestamp 1679581782
transform 1 0 13248 0 1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_133
timestamp 1679581782
transform 1 0 13920 0 1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_140
timestamp 1679581782
transform 1 0 14592 0 1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_147
timestamp 1679581782
transform 1 0 15264 0 1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_154
timestamp 1679581782
transform 1 0 15936 0 1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_161
timestamp 1679581782
transform 1 0 16608 0 1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_168
timestamp 1679581782
transform 1 0 17280 0 1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_175
timestamp 1679581782
transform 1 0 17952 0 1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_182
timestamp 1679581782
transform 1 0 18624 0 1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_189
timestamp 1679581782
transform 1 0 19296 0 1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_196
timestamp 1679581782
transform 1 0 19968 0 1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_203
timestamp 1679581782
transform 1 0 20640 0 1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_210
timestamp 1679581782
transform 1 0 21312 0 1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_217
timestamp 1679581782
transform 1 0 21984 0 1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_224
timestamp 1679581782
transform 1 0 22656 0 1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_231
timestamp 1679581782
transform 1 0 23328 0 1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_238
timestamp 1679581782
transform 1 0 24000 0 1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_245
timestamp 1679581782
transform 1 0 24672 0 1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_252
timestamp 1679581782
transform 1 0 25344 0 1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_259
timestamp 1679581782
transform 1 0 26016 0 1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_266
timestamp 1679581782
transform 1 0 26688 0 1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_273
timestamp 1679581782
transform 1 0 27360 0 1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_280
timestamp 1679581782
transform 1 0 28032 0 1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_287
timestamp 1679581782
transform 1 0 28704 0 1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_294
timestamp 1679581782
transform 1 0 29376 0 1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_301
timestamp 1679581782
transform 1 0 30048 0 1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_308
timestamp 1679581782
transform 1 0 30720 0 1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_315
timestamp 1679581782
transform 1 0 31392 0 1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_322
timestamp 1679581782
transform 1 0 32064 0 1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_329
timestamp 1679581782
transform 1 0 32736 0 1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_336
timestamp 1679581782
transform 1 0 33408 0 1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_343
timestamp 1679581782
transform 1 0 34080 0 1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_350
timestamp 1679581782
transform 1 0 34752 0 1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_357
timestamp 1679581782
transform 1 0 35424 0 1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_364
timestamp 1679581782
transform 1 0 36096 0 1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_371
timestamp 1679581782
transform 1 0 36768 0 1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_378
timestamp 1679581782
transform 1 0 37440 0 1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_385
timestamp 1679581782
transform 1 0 38112 0 1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_392
timestamp 1679581782
transform 1 0 38784 0 1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_399
timestamp 1679581782
transform 1 0 39456 0 1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_406
timestamp 1679581782
transform 1 0 40128 0 1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_413
timestamp 1679581782
transform 1 0 40800 0 1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_420
timestamp 1679581782
transform 1 0 41472 0 1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_427
timestamp 1679581782
transform 1 0 42144 0 1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_434
timestamp 1679581782
transform 1 0 42816 0 1 9072
box -48 -56 720 834
use sg13g2_fill_2  FILLER_10_441
timestamp 1677580104
transform 1 0 43488 0 1 9072
box -48 -56 240 834
use sg13g2_decap_8  FILLER_11_0
timestamp 1679581782
transform 1 0 1152 0 -1 10584
box -48 -56 720 834
use sg13g2_fill_2  FILLER_11_7
timestamp 1677580104
transform 1 0 1824 0 -1 10584
box -48 -56 240 834
use sg13g2_decap_8  FILLER_11_13
timestamp 1679581782
transform 1 0 2400 0 -1 10584
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_20
timestamp 1679581782
transform 1 0 3072 0 -1 10584
box -48 -56 720 834
use sg13g2_decap_4  FILLER_11_27
timestamp 1679577901
transform 1 0 3744 0 -1 10584
box -48 -56 432 834
use sg13g2_decap_8  FILLER_11_35
timestamp 1679581782
transform 1 0 4512 0 -1 10584
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_42
timestamp 1679581782
transform 1 0 5184 0 -1 10584
box -48 -56 720 834
use sg13g2_decap_4  FILLER_11_49
timestamp 1679577901
transform 1 0 5856 0 -1 10584
box -48 -56 432 834
use sg13g2_decap_8  FILLER_11_57
timestamp 1679581782
transform 1 0 6624 0 -1 10584
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_64
timestamp 1679581782
transform 1 0 7296 0 -1 10584
box -48 -56 720 834
use sg13g2_decap_4  FILLER_11_71
timestamp 1679577901
transform 1 0 7968 0 -1 10584
box -48 -56 432 834
use sg13g2_decap_8  FILLER_11_79
timestamp 1679581782
transform 1 0 8736 0 -1 10584
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_86
timestamp 1679581782
transform 1 0 9408 0 -1 10584
box -48 -56 720 834
use sg13g2_decap_4  FILLER_11_93
timestamp 1679577901
transform 1 0 10080 0 -1 10584
box -48 -56 432 834
use sg13g2_decap_8  FILLER_11_101
timestamp 1679581782
transform 1 0 10848 0 -1 10584
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_108
timestamp 1679581782
transform 1 0 11520 0 -1 10584
box -48 -56 720 834
use sg13g2_decap_4  FILLER_11_115
timestamp 1679577901
transform 1 0 12192 0 -1 10584
box -48 -56 432 834
use sg13g2_decap_8  FILLER_11_123
timestamp 1679581782
transform 1 0 12960 0 -1 10584
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_130
timestamp 1679581782
transform 1 0 13632 0 -1 10584
box -48 -56 720 834
use sg13g2_decap_4  FILLER_11_137
timestamp 1679577901
transform 1 0 14304 0 -1 10584
box -48 -56 432 834
use sg13g2_decap_8  FILLER_11_145
timestamp 1679581782
transform 1 0 15072 0 -1 10584
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_152
timestamp 1679581782
transform 1 0 15744 0 -1 10584
box -48 -56 720 834
use sg13g2_decap_4  FILLER_11_159
timestamp 1679577901
transform 1 0 16416 0 -1 10584
box -48 -56 432 834
use sg13g2_decap_8  FILLER_11_167
timestamp 1679581782
transform 1 0 17184 0 -1 10584
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_174
timestamp 1679581782
transform 1 0 17856 0 -1 10584
box -48 -56 720 834
use sg13g2_decap_4  FILLER_11_181
timestamp 1679577901
transform 1 0 18528 0 -1 10584
box -48 -56 432 834
use sg13g2_decap_8  FILLER_11_189
timestamp 1679581782
transform 1 0 19296 0 -1 10584
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_196
timestamp 1679581782
transform 1 0 19968 0 -1 10584
box -48 -56 720 834
use sg13g2_decap_4  FILLER_11_203
timestamp 1679577901
transform 1 0 20640 0 -1 10584
box -48 -56 432 834
use sg13g2_decap_8  FILLER_11_211
timestamp 1679581782
transform 1 0 21408 0 -1 10584
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_218
timestamp 1679581782
transform 1 0 22080 0 -1 10584
box -48 -56 720 834
use sg13g2_decap_4  FILLER_11_225
timestamp 1679577901
transform 1 0 22752 0 -1 10584
box -48 -56 432 834
use sg13g2_decap_8  FILLER_11_233
timestamp 1679581782
transform 1 0 23520 0 -1 10584
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_240
timestamp 1679581782
transform 1 0 24192 0 -1 10584
box -48 -56 720 834
use sg13g2_decap_4  FILLER_11_247
timestamp 1679577901
transform 1 0 24864 0 -1 10584
box -48 -56 432 834
use sg13g2_decap_8  FILLER_11_255
timestamp 1679581782
transform 1 0 25632 0 -1 10584
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_262
timestamp 1679581782
transform 1 0 26304 0 -1 10584
box -48 -56 720 834
use sg13g2_decap_4  FILLER_11_269
timestamp 1679577901
transform 1 0 26976 0 -1 10584
box -48 -56 432 834
use sg13g2_decap_8  FILLER_11_277
timestamp 1679581782
transform 1 0 27744 0 -1 10584
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_284
timestamp 1679581782
transform 1 0 28416 0 -1 10584
box -48 -56 720 834
use sg13g2_decap_4  FILLER_11_291
timestamp 1679577901
transform 1 0 29088 0 -1 10584
box -48 -56 432 834
use sg13g2_decap_8  FILLER_11_299
timestamp 1679581782
transform 1 0 29856 0 -1 10584
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_306
timestamp 1679581782
transform 1 0 30528 0 -1 10584
box -48 -56 720 834
use sg13g2_decap_4  FILLER_11_313
timestamp 1679577901
transform 1 0 31200 0 -1 10584
box -48 -56 432 834
use sg13g2_decap_8  FILLER_11_321
timestamp 1679581782
transform 1 0 31968 0 -1 10584
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_328
timestamp 1679581782
transform 1 0 32640 0 -1 10584
box -48 -56 720 834
use sg13g2_decap_4  FILLER_11_335
timestamp 1679577901
transform 1 0 33312 0 -1 10584
box -48 -56 432 834
use sg13g2_decap_8  FILLER_11_343
timestamp 1679581782
transform 1 0 34080 0 -1 10584
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_350
timestamp 1679581782
transform 1 0 34752 0 -1 10584
box -48 -56 720 834
use sg13g2_decap_4  FILLER_11_357
timestamp 1679577901
transform 1 0 35424 0 -1 10584
box -48 -56 432 834
use sg13g2_decap_8  FILLER_11_365
timestamp 1679581782
transform 1 0 36192 0 -1 10584
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_372
timestamp 1679581782
transform 1 0 36864 0 -1 10584
box -48 -56 720 834
use sg13g2_decap_4  FILLER_11_379
timestamp 1679577901
transform 1 0 37536 0 -1 10584
box -48 -56 432 834
use sg13g2_decap_8  FILLER_11_387
timestamp 1679581782
transform 1 0 38304 0 -1 10584
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_394
timestamp 1679581782
transform 1 0 38976 0 -1 10584
box -48 -56 720 834
use sg13g2_decap_4  FILLER_11_401
timestamp 1679577901
transform 1 0 39648 0 -1 10584
box -48 -56 432 834
use sg13g2_decap_8  FILLER_11_409
timestamp 1679581782
transform 1 0 40416 0 -1 10584
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_416
timestamp 1679581782
transform 1 0 41088 0 -1 10584
box -48 -56 720 834
use sg13g2_decap_4  FILLER_11_423
timestamp 1679577901
transform 1 0 41760 0 -1 10584
box -48 -56 432 834
use sg13g2_decap_4  FILLER_11_431
timestamp 1679577901
transform 1 0 42528 0 -1 10584
box -48 -56 432 834
use sg13g2_fill_2  FILLER_11_435
timestamp 1677580104
transform 1 0 42912 0 -1 10584
box -48 -56 240 834
use sg13g2_fill_2  FILLER_11_453
timestamp 1677580104
transform 1 0 44640 0 -1 10584
box -48 -56 240 834
use sg13g2_buf_1  output1
timestamp 1676381911
transform 1 0 44064 0 1 1512
box -48 -56 432 834
use sg13g2_buf_1  output2
timestamp 1676381911
transform 1 0 44448 0 -1 4536
box -48 -56 432 834
use sg13g2_buf_1  output3
timestamp 1676381911
transform 1 0 44832 0 -1 4536
box -48 -56 432 834
use sg13g2_buf_1  output4
timestamp 1676381911
transform 1 0 44448 0 1 4536
box -48 -56 432 834
use sg13g2_buf_1  output5
timestamp 1676381911
transform 1 0 44832 0 1 4536
box -48 -56 432 834
use sg13g2_buf_1  output6
timestamp 1676381911
transform 1 0 44448 0 -1 6048
box -48 -56 432 834
use sg13g2_buf_1  output7
timestamp 1676381911
transform 1 0 44832 0 -1 6048
box -48 -56 432 834
use sg13g2_buf_1  output8
timestamp 1676381911
transform 1 0 44448 0 1 6048
box -48 -56 432 834
use sg13g2_buf_1  output9
timestamp 1676381911
transform 1 0 44832 0 1 6048
box -48 -56 432 834
use sg13g2_buf_1  output10
timestamp 1676381911
transform 1 0 44448 0 -1 7560
box -48 -56 432 834
use sg13g2_buf_1  output11
timestamp 1676381911
transform 1 0 44832 0 -1 7560
box -48 -56 432 834
use sg13g2_buf_1  output12
timestamp 1676381911
transform 1 0 43680 0 1 1512
box -48 -56 432 834
use sg13g2_buf_1  output13
timestamp 1676381911
transform 1 0 44832 0 1 7560
box -48 -56 432 834
use sg13g2_buf_1  output14
timestamp 1676381911
transform 1 0 44448 0 1 7560
box -48 -56 432 834
use sg13g2_buf_1  output15
timestamp 1676381911
transform 1 0 44832 0 -1 9072
box -48 -56 432 834
use sg13g2_buf_1  output16
timestamp 1676381911
transform 1 0 44448 0 -1 9072
box -48 -56 432 834
use sg13g2_buf_1  output17
timestamp 1676381911
transform 1 0 44832 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  output18
timestamp 1676381911
transform 1 0 44448 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  output19
timestamp 1676381911
transform 1 0 44832 0 -1 10584
box -48 -56 432 834
use sg13g2_buf_1  output20
timestamp 1676381911
transform 1 0 43872 0 -1 10584
box -48 -56 432 834
use sg13g2_buf_1  output21
timestamp 1676381911
transform 1 0 43488 0 -1 10584
box -48 -56 432 834
use sg13g2_buf_1  output22
timestamp 1676381911
transform 1 0 44064 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  output23
timestamp 1676381911
transform 1 0 44064 0 -1 3024
box -48 -56 432 834
use sg13g2_buf_1  output24
timestamp 1676381911
transform 1 0 43104 0 -1 10584
box -48 -56 432 834
use sg13g2_buf_1  output25
timestamp 1676381911
transform 1 0 43680 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  output26
timestamp 1676381911
transform 1 0 44448 0 1 1512
box -48 -56 432 834
use sg13g2_buf_1  output27
timestamp 1676381911
transform 1 0 44832 0 1 1512
box -48 -56 432 834
use sg13g2_buf_1  output28
timestamp 1676381911
transform 1 0 44448 0 -1 3024
box -48 -56 432 834
use sg13g2_buf_1  output29
timestamp 1676381911
transform 1 0 44832 0 -1 3024
box -48 -56 432 834
use sg13g2_buf_1  output30
timestamp 1676381911
transform 1 0 44448 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  output31
timestamp 1676381911
transform 1 0 44064 0 -1 4536
box -48 -56 432 834
use sg13g2_buf_1  output32
timestamp 1676381911
transform 1 0 44832 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  output33
timestamp 1676381911
transform -1 0 4512 0 -1 10584
box -48 -56 432 834
use sg13g2_buf_1  output34
timestamp 1676381911
transform -1 0 25632 0 -1 10584
box -48 -56 432 834
use sg13g2_buf_1  output35
timestamp 1676381911
transform -1 0 27744 0 -1 10584
box -48 -56 432 834
use sg13g2_buf_1  output36
timestamp 1676381911
transform -1 0 29856 0 -1 10584
box -48 -56 432 834
use sg13g2_buf_1  output37
timestamp 1676381911
transform -1 0 31968 0 -1 10584
box -48 -56 432 834
use sg13g2_buf_1  output38
timestamp 1676381911
transform -1 0 34080 0 -1 10584
box -48 -56 432 834
use sg13g2_buf_1  output39
timestamp 1676381911
transform -1 0 36192 0 -1 10584
box -48 -56 432 834
use sg13g2_buf_1  output40
timestamp 1676381911
transform -1 0 38304 0 -1 10584
box -48 -56 432 834
use sg13g2_buf_1  output41
timestamp 1676381911
transform -1 0 40416 0 -1 10584
box -48 -56 432 834
use sg13g2_buf_1  output42
timestamp 1676381911
transform -1 0 42528 0 -1 10584
box -48 -56 432 834
use sg13g2_buf_1  output43
timestamp 1676381911
transform -1 0 44640 0 -1 10584
box -48 -56 432 834
use sg13g2_buf_1  output44
timestamp 1676381911
transform -1 0 6624 0 -1 10584
box -48 -56 432 834
use sg13g2_buf_1  output45
timestamp 1676381911
transform -1 0 8736 0 -1 10584
box -48 -56 432 834
use sg13g2_buf_1  output46
timestamp 1676381911
transform -1 0 10848 0 -1 10584
box -48 -56 432 834
use sg13g2_buf_1  output47
timestamp 1676381911
transform -1 0 12960 0 -1 10584
box -48 -56 432 834
use sg13g2_buf_1  output48
timestamp 1676381911
transform -1 0 15072 0 -1 10584
box -48 -56 432 834
use sg13g2_buf_1  output49
timestamp 1676381911
transform -1 0 17184 0 -1 10584
box -48 -56 432 834
use sg13g2_buf_1  output50
timestamp 1676381911
transform -1 0 19296 0 -1 10584
box -48 -56 432 834
use sg13g2_buf_1  output51
timestamp 1676381911
transform -1 0 21408 0 -1 10584
box -48 -56 432 834
use sg13g2_buf_1  output52
timestamp 1676381911
transform -1 0 23520 0 -1 10584
box -48 -56 432 834
use sg13g2_buf_1  output53
timestamp 1676381911
transform -1 0 21600 0 -1 3024
box -48 -56 432 834
use sg13g2_buf_1  output54
timestamp 1676381911
transform 1 0 20832 0 1 1512
box -48 -56 432 834
use sg13g2_buf_1  output55
timestamp 1676381911
transform -1 0 21984 0 -1 3024
box -48 -56 432 834
use sg13g2_buf_1  output56
timestamp 1676381911
transform 1 0 21216 0 1 1512
box -48 -56 432 834
use sg13g2_buf_1  output57
timestamp 1676381911
transform -1 0 22368 0 -1 3024
box -48 -56 432 834
use sg13g2_buf_1  output58
timestamp 1676381911
transform 1 0 21600 0 1 1512
box -48 -56 432 834
use sg13g2_buf_1  output59
timestamp 1676381911
transform -1 0 22752 0 -1 3024
box -48 -56 432 834
use sg13g2_buf_1  output60
timestamp 1676381911
transform 1 0 21984 0 1 1512
box -48 -56 432 834
use sg13g2_buf_1  output61
timestamp 1676381911
transform -1 0 23136 0 -1 3024
box -48 -56 432 834
use sg13g2_buf_1  output62
timestamp 1676381911
transform 1 0 22368 0 1 1512
box -48 -56 432 834
use sg13g2_buf_1  output63
timestamp 1676381911
transform -1 0 23520 0 -1 3024
box -48 -56 432 834
use sg13g2_buf_1  output64
timestamp 1676381911
transform 1 0 22752 0 1 1512
box -48 -56 432 834
use sg13g2_buf_1  output65
timestamp 1676381911
transform -1 0 23904 0 -1 3024
box -48 -56 432 834
use sg13g2_buf_1  output66
timestamp 1676381911
transform 1 0 23136 0 1 1512
box -48 -56 432 834
use sg13g2_buf_1  output67
timestamp 1676381911
transform 1 0 23520 0 1 1512
box -48 -56 432 834
use sg13g2_buf_1  output68
timestamp 1676381911
transform 1 0 23904 0 1 1512
box -48 -56 432 834
use sg13g2_buf_1  output69
timestamp 1676381911
transform -1 0 24672 0 1 1512
box -48 -56 432 834
use sg13g2_buf_1  output70
timestamp 1676381911
transform -1 0 25056 0 1 1512
box -48 -56 432 834
use sg13g2_buf_1  output71
timestamp 1676381911
transform -1 0 25440 0 1 1512
box -48 -56 432 834
use sg13g2_buf_1  output72
timestamp 1676381911
transform -1 0 25824 0 1 1512
box -48 -56 432 834
use sg13g2_buf_1  output73
timestamp 1676381911
transform -1 0 26208 0 1 1512
box -48 -56 432 834
use sg13g2_buf_1  output74
timestamp 1676381911
transform -1 0 28128 0 1 1512
box -48 -56 432 834
use sg13g2_buf_1  output75
timestamp 1676381911
transform -1 0 27552 0 -1 3024
box -48 -56 432 834
use sg13g2_buf_1  output76
timestamp 1676381911
transform -1 0 28512 0 1 1512
box -48 -56 432 834
use sg13g2_buf_1  output77
timestamp 1676381911
transform -1 0 27936 0 -1 3024
box -48 -56 432 834
use sg13g2_buf_1  output78
timestamp 1676381911
transform -1 0 28896 0 1 1512
box -48 -56 432 834
use sg13g2_buf_1  output79
timestamp 1676381911
transform -1 0 28320 0 -1 3024
box -48 -56 432 834
use sg13g2_buf_1  output80
timestamp 1676381911
transform -1 0 25632 0 -1 3024
box -48 -56 432 834
use sg13g2_buf_1  output81
timestamp 1676381911
transform -1 0 26592 0 1 1512
box -48 -56 432 834
use sg13g2_buf_1  output82
timestamp 1676381911
transform -1 0 26016 0 -1 3024
box -48 -56 432 834
use sg13g2_buf_1  output83
timestamp 1676381911
transform -1 0 26976 0 1 1512
box -48 -56 432 834
use sg13g2_buf_1  output84
timestamp 1676381911
transform -1 0 26400 0 -1 3024
box -48 -56 432 834
use sg13g2_buf_1  output85
timestamp 1676381911
transform -1 0 27360 0 1 1512
box -48 -56 432 834
use sg13g2_buf_1  output86
timestamp 1676381911
transform -1 0 26784 0 -1 3024
box -48 -56 432 834
use sg13g2_buf_1  output87
timestamp 1676381911
transform -1 0 27744 0 1 1512
box -48 -56 432 834
use sg13g2_buf_1  output88
timestamp 1676381911
transform -1 0 27168 0 -1 3024
box -48 -56 432 834
use sg13g2_buf_1  output89
timestamp 1676381911
transform -1 0 29280 0 1 1512
box -48 -56 432 834
use sg13g2_buf_1  output90
timestamp 1676381911
transform -1 0 31200 0 1 1512
box -48 -56 432 834
use sg13g2_buf_1  output91
timestamp 1676381911
transform -1 0 30624 0 -1 3024
box -48 -56 432 834
use sg13g2_buf_1  output92
timestamp 1676381911
transform -1 0 31584 0 1 1512
box -48 -56 432 834
use sg13g2_buf_1  output93
timestamp 1676381911
transform -1 0 31008 0 -1 3024
box -48 -56 432 834
use sg13g2_buf_1  output94
timestamp 1676381911
transform -1 0 31968 0 1 1512
box -48 -56 432 834
use sg13g2_buf_1  output95
timestamp 1676381911
transform -1 0 31392 0 -1 3024
box -48 -56 432 834
use sg13g2_buf_1  output96
timestamp 1676381911
transform -1 0 28704 0 -1 3024
box -48 -56 432 834
use sg13g2_buf_1  output97
timestamp 1676381911
transform -1 0 29664 0 1 1512
box -48 -56 432 834
use sg13g2_buf_1  output98
timestamp 1676381911
transform -1 0 29088 0 -1 3024
box -48 -56 432 834
use sg13g2_buf_1  output99
timestamp 1676381911
transform -1 0 30048 0 1 1512
box -48 -56 432 834
use sg13g2_buf_1  output100
timestamp 1676381911
transform -1 0 29472 0 -1 3024
box -48 -56 432 834
use sg13g2_buf_1  output101
timestamp 1676381911
transform -1 0 30432 0 1 1512
box -48 -56 432 834
use sg13g2_buf_1  output102
timestamp 1676381911
transform -1 0 29856 0 -1 3024
box -48 -56 432 834
use sg13g2_buf_1  output103
timestamp 1676381911
transform -1 0 30816 0 1 1512
box -48 -56 432 834
use sg13g2_buf_1  output104
timestamp 1676381911
transform -1 0 30240 0 -1 3024
box -48 -56 432 834
use sg13g2_buf_1  output105
timestamp 1676381911
transform -1 0 2400 0 -1 10584
box -48 -56 432 834
<< labels >>
flabel metal3 s 20984 0 21064 80 0 FreeSans 320 0 0 0 Ci
port 0 nsew signal input
flabel metal2 s 0 716 90 796 0 FreeSans 320 0 0 0 FrameData[0]
port 1 nsew signal input
flabel metal2 s 0 4076 90 4156 0 FreeSans 320 0 0 0 FrameData[10]
port 2 nsew signal input
flabel metal2 s 0 4412 90 4492 0 FreeSans 320 0 0 0 FrameData[11]
port 3 nsew signal input
flabel metal2 s 0 4748 90 4828 0 FreeSans 320 0 0 0 FrameData[12]
port 4 nsew signal input
flabel metal2 s 0 5084 90 5164 0 FreeSans 320 0 0 0 FrameData[13]
port 5 nsew signal input
flabel metal2 s 0 5420 90 5500 0 FreeSans 320 0 0 0 FrameData[14]
port 6 nsew signal input
flabel metal2 s 0 5756 90 5836 0 FreeSans 320 0 0 0 FrameData[15]
port 7 nsew signal input
flabel metal2 s 0 6092 90 6172 0 FreeSans 320 0 0 0 FrameData[16]
port 8 nsew signal input
flabel metal2 s 0 6428 90 6508 0 FreeSans 320 0 0 0 FrameData[17]
port 9 nsew signal input
flabel metal2 s 0 6764 90 6844 0 FreeSans 320 0 0 0 FrameData[18]
port 10 nsew signal input
flabel metal2 s 0 7100 90 7180 0 FreeSans 320 0 0 0 FrameData[19]
port 11 nsew signal input
flabel metal2 s 0 1052 90 1132 0 FreeSans 320 0 0 0 FrameData[1]
port 12 nsew signal input
flabel metal2 s 0 7436 90 7516 0 FreeSans 320 0 0 0 FrameData[20]
port 13 nsew signal input
flabel metal2 s 0 7772 90 7852 0 FreeSans 320 0 0 0 FrameData[21]
port 14 nsew signal input
flabel metal2 s 0 8108 90 8188 0 FreeSans 320 0 0 0 FrameData[22]
port 15 nsew signal input
flabel metal2 s 0 8444 90 8524 0 FreeSans 320 0 0 0 FrameData[23]
port 16 nsew signal input
flabel metal2 s 0 8780 90 8860 0 FreeSans 320 0 0 0 FrameData[24]
port 17 nsew signal input
flabel metal2 s 0 9116 90 9196 0 FreeSans 320 0 0 0 FrameData[25]
port 18 nsew signal input
flabel metal2 s 0 9452 90 9532 0 FreeSans 320 0 0 0 FrameData[26]
port 19 nsew signal input
flabel metal2 s 0 9788 90 9868 0 FreeSans 320 0 0 0 FrameData[27]
port 20 nsew signal input
flabel metal2 s 0 10124 90 10204 0 FreeSans 320 0 0 0 FrameData[28]
port 21 nsew signal input
flabel metal2 s 0 10460 90 10540 0 FreeSans 320 0 0 0 FrameData[29]
port 22 nsew signal input
flabel metal2 s 0 1388 90 1468 0 FreeSans 320 0 0 0 FrameData[2]
port 23 nsew signal input
flabel metal2 s 0 10796 90 10876 0 FreeSans 320 0 0 0 FrameData[30]
port 24 nsew signal input
flabel metal2 s 0 11132 90 11212 0 FreeSans 320 0 0 0 FrameData[31]
port 25 nsew signal input
flabel metal2 s 0 1724 90 1804 0 FreeSans 320 0 0 0 FrameData[3]
port 26 nsew signal input
flabel metal2 s 0 2060 90 2140 0 FreeSans 320 0 0 0 FrameData[4]
port 27 nsew signal input
flabel metal2 s 0 2396 90 2476 0 FreeSans 320 0 0 0 FrameData[5]
port 28 nsew signal input
flabel metal2 s 0 2732 90 2812 0 FreeSans 320 0 0 0 FrameData[6]
port 29 nsew signal input
flabel metal2 s 0 3068 90 3148 0 FreeSans 320 0 0 0 FrameData[7]
port 30 nsew signal input
flabel metal2 s 0 3404 90 3484 0 FreeSans 320 0 0 0 FrameData[8]
port 31 nsew signal input
flabel metal2 s 0 3740 90 3820 0 FreeSans 320 0 0 0 FrameData[9]
port 32 nsew signal input
flabel metal2 s 46278 716 46368 796 0 FreeSans 320 0 0 0 FrameData_O[0]
port 33 nsew signal output
flabel metal2 s 46278 4076 46368 4156 0 FreeSans 320 0 0 0 FrameData_O[10]
port 34 nsew signal output
flabel metal2 s 46278 4412 46368 4492 0 FreeSans 320 0 0 0 FrameData_O[11]
port 35 nsew signal output
flabel metal2 s 46278 4748 46368 4828 0 FreeSans 320 0 0 0 FrameData_O[12]
port 36 nsew signal output
flabel metal2 s 46278 5084 46368 5164 0 FreeSans 320 0 0 0 FrameData_O[13]
port 37 nsew signal output
flabel metal2 s 46278 5420 46368 5500 0 FreeSans 320 0 0 0 FrameData_O[14]
port 38 nsew signal output
flabel metal2 s 46278 5756 46368 5836 0 FreeSans 320 0 0 0 FrameData_O[15]
port 39 nsew signal output
flabel metal2 s 46278 6092 46368 6172 0 FreeSans 320 0 0 0 FrameData_O[16]
port 40 nsew signal output
flabel metal2 s 46278 6428 46368 6508 0 FreeSans 320 0 0 0 FrameData_O[17]
port 41 nsew signal output
flabel metal2 s 46278 6764 46368 6844 0 FreeSans 320 0 0 0 FrameData_O[18]
port 42 nsew signal output
flabel metal2 s 46278 7100 46368 7180 0 FreeSans 320 0 0 0 FrameData_O[19]
port 43 nsew signal output
flabel metal2 s 46278 1052 46368 1132 0 FreeSans 320 0 0 0 FrameData_O[1]
port 44 nsew signal output
flabel metal2 s 46278 7436 46368 7516 0 FreeSans 320 0 0 0 FrameData_O[20]
port 45 nsew signal output
flabel metal2 s 46278 7772 46368 7852 0 FreeSans 320 0 0 0 FrameData_O[21]
port 46 nsew signal output
flabel metal2 s 46278 8108 46368 8188 0 FreeSans 320 0 0 0 FrameData_O[22]
port 47 nsew signal output
flabel metal2 s 46278 8444 46368 8524 0 FreeSans 320 0 0 0 FrameData_O[23]
port 48 nsew signal output
flabel metal2 s 46278 8780 46368 8860 0 FreeSans 320 0 0 0 FrameData_O[24]
port 49 nsew signal output
flabel metal2 s 46278 9116 46368 9196 0 FreeSans 320 0 0 0 FrameData_O[25]
port 50 nsew signal output
flabel metal2 s 46278 9452 46368 9532 0 FreeSans 320 0 0 0 FrameData_O[26]
port 51 nsew signal output
flabel metal2 s 46278 9788 46368 9868 0 FreeSans 320 0 0 0 FrameData_O[27]
port 52 nsew signal output
flabel metal2 s 46278 10124 46368 10204 0 FreeSans 320 0 0 0 FrameData_O[28]
port 53 nsew signal output
flabel metal2 s 46278 10460 46368 10540 0 FreeSans 320 0 0 0 FrameData_O[29]
port 54 nsew signal output
flabel metal2 s 46278 1388 46368 1468 0 FreeSans 320 0 0 0 FrameData_O[2]
port 55 nsew signal output
flabel metal2 s 46278 10796 46368 10876 0 FreeSans 320 0 0 0 FrameData_O[30]
port 56 nsew signal output
flabel metal2 s 46278 11132 46368 11212 0 FreeSans 320 0 0 0 FrameData_O[31]
port 57 nsew signal output
flabel metal2 s 46278 1724 46368 1804 0 FreeSans 320 0 0 0 FrameData_O[3]
port 58 nsew signal output
flabel metal2 s 46278 2060 46368 2140 0 FreeSans 320 0 0 0 FrameData_O[4]
port 59 nsew signal output
flabel metal2 s 46278 2396 46368 2476 0 FreeSans 320 0 0 0 FrameData_O[5]
port 60 nsew signal output
flabel metal2 s 46278 2732 46368 2812 0 FreeSans 320 0 0 0 FrameData_O[6]
port 61 nsew signal output
flabel metal2 s 46278 3068 46368 3148 0 FreeSans 320 0 0 0 FrameData_O[7]
port 62 nsew signal output
flabel metal2 s 46278 3404 46368 3484 0 FreeSans 320 0 0 0 FrameData_O[8]
port 63 nsew signal output
flabel metal2 s 46278 3740 46368 3820 0 FreeSans 320 0 0 0 FrameData_O[9]
port 64 nsew signal output
flabel metal3 s 31352 0 31432 80 0 FreeSans 320 0 0 0 FrameStrobe[0]
port 65 nsew signal input
flabel metal3 s 33272 0 33352 80 0 FreeSans 320 0 0 0 FrameStrobe[10]
port 66 nsew signal input
flabel metal3 s 33464 0 33544 80 0 FreeSans 320 0 0 0 FrameStrobe[11]
port 67 nsew signal input
flabel metal3 s 33656 0 33736 80 0 FreeSans 320 0 0 0 FrameStrobe[12]
port 68 nsew signal input
flabel metal3 s 33848 0 33928 80 0 FreeSans 320 0 0 0 FrameStrobe[13]
port 69 nsew signal input
flabel metal3 s 34040 0 34120 80 0 FreeSans 320 0 0 0 FrameStrobe[14]
port 70 nsew signal input
flabel metal3 s 34232 0 34312 80 0 FreeSans 320 0 0 0 FrameStrobe[15]
port 71 nsew signal input
flabel metal3 s 34424 0 34504 80 0 FreeSans 320 0 0 0 FrameStrobe[16]
port 72 nsew signal input
flabel metal3 s 34616 0 34696 80 0 FreeSans 320 0 0 0 FrameStrobe[17]
port 73 nsew signal input
flabel metal3 s 34808 0 34888 80 0 FreeSans 320 0 0 0 FrameStrobe[18]
port 74 nsew signal input
flabel metal3 s 35000 0 35080 80 0 FreeSans 320 0 0 0 FrameStrobe[19]
port 75 nsew signal input
flabel metal3 s 31544 0 31624 80 0 FreeSans 320 0 0 0 FrameStrobe[1]
port 76 nsew signal input
flabel metal3 s 31736 0 31816 80 0 FreeSans 320 0 0 0 FrameStrobe[2]
port 77 nsew signal input
flabel metal3 s 31928 0 32008 80 0 FreeSans 320 0 0 0 FrameStrobe[3]
port 78 nsew signal input
flabel metal3 s 32120 0 32200 80 0 FreeSans 320 0 0 0 FrameStrobe[4]
port 79 nsew signal input
flabel metal3 s 32312 0 32392 80 0 FreeSans 320 0 0 0 FrameStrobe[5]
port 80 nsew signal input
flabel metal3 s 32504 0 32584 80 0 FreeSans 320 0 0 0 FrameStrobe[6]
port 81 nsew signal input
flabel metal3 s 32696 0 32776 80 0 FreeSans 320 0 0 0 FrameStrobe[7]
port 82 nsew signal input
flabel metal3 s 32888 0 32968 80 0 FreeSans 320 0 0 0 FrameStrobe[8]
port 83 nsew signal input
flabel metal3 s 33080 0 33160 80 0 FreeSans 320 0 0 0 FrameStrobe[9]
port 84 nsew signal input
flabel metal3 s 4088 12100 4168 12180 0 FreeSans 320 0 0 0 FrameStrobe_O[0]
port 85 nsew signal output
flabel metal3 s 25208 12100 25288 12180 0 FreeSans 320 0 0 0 FrameStrobe_O[10]
port 86 nsew signal output
flabel metal3 s 27320 12100 27400 12180 0 FreeSans 320 0 0 0 FrameStrobe_O[11]
port 87 nsew signal output
flabel metal3 s 29432 12100 29512 12180 0 FreeSans 320 0 0 0 FrameStrobe_O[12]
port 88 nsew signal output
flabel metal3 s 31544 12100 31624 12180 0 FreeSans 320 0 0 0 FrameStrobe_O[13]
port 89 nsew signal output
flabel metal3 s 33656 12100 33736 12180 0 FreeSans 320 0 0 0 FrameStrobe_O[14]
port 90 nsew signal output
flabel metal3 s 35768 12100 35848 12180 0 FreeSans 320 0 0 0 FrameStrobe_O[15]
port 91 nsew signal output
flabel metal3 s 37880 12100 37960 12180 0 FreeSans 320 0 0 0 FrameStrobe_O[16]
port 92 nsew signal output
flabel metal3 s 39992 12100 40072 12180 0 FreeSans 320 0 0 0 FrameStrobe_O[17]
port 93 nsew signal output
flabel metal3 s 42104 12100 42184 12180 0 FreeSans 320 0 0 0 FrameStrobe_O[18]
port 94 nsew signal output
flabel metal3 s 44216 12100 44296 12180 0 FreeSans 320 0 0 0 FrameStrobe_O[19]
port 95 nsew signal output
flabel metal3 s 6200 12100 6280 12180 0 FreeSans 320 0 0 0 FrameStrobe_O[1]
port 96 nsew signal output
flabel metal3 s 8312 12100 8392 12180 0 FreeSans 320 0 0 0 FrameStrobe_O[2]
port 97 nsew signal output
flabel metal3 s 10424 12100 10504 12180 0 FreeSans 320 0 0 0 FrameStrobe_O[3]
port 98 nsew signal output
flabel metal3 s 12536 12100 12616 12180 0 FreeSans 320 0 0 0 FrameStrobe_O[4]
port 99 nsew signal output
flabel metal3 s 14648 12100 14728 12180 0 FreeSans 320 0 0 0 FrameStrobe_O[5]
port 100 nsew signal output
flabel metal3 s 16760 12100 16840 12180 0 FreeSans 320 0 0 0 FrameStrobe_O[6]
port 101 nsew signal output
flabel metal3 s 18872 12100 18952 12180 0 FreeSans 320 0 0 0 FrameStrobe_O[7]
port 102 nsew signal output
flabel metal3 s 20984 12100 21064 12180 0 FreeSans 320 0 0 0 FrameStrobe_O[8]
port 103 nsew signal output
flabel metal3 s 23096 12100 23176 12180 0 FreeSans 320 0 0 0 FrameStrobe_O[9]
port 104 nsew signal output
flabel metal3 s 11000 0 11080 80 0 FreeSans 320 0 0 0 N1END[0]
port 105 nsew signal input
flabel metal3 s 11192 0 11272 80 0 FreeSans 320 0 0 0 N1END[1]
port 106 nsew signal input
flabel metal3 s 11384 0 11464 80 0 FreeSans 320 0 0 0 N1END[2]
port 107 nsew signal input
flabel metal3 s 11576 0 11656 80 0 FreeSans 320 0 0 0 N1END[3]
port 108 nsew signal input
flabel metal3 s 13304 0 13384 80 0 FreeSans 320 0 0 0 N2END[0]
port 109 nsew signal input
flabel metal3 s 13496 0 13576 80 0 FreeSans 320 0 0 0 N2END[1]
port 110 nsew signal input
flabel metal3 s 13688 0 13768 80 0 FreeSans 320 0 0 0 N2END[2]
port 111 nsew signal input
flabel metal3 s 13880 0 13960 80 0 FreeSans 320 0 0 0 N2END[3]
port 112 nsew signal input
flabel metal3 s 14072 0 14152 80 0 FreeSans 320 0 0 0 N2END[4]
port 113 nsew signal input
flabel metal3 s 14264 0 14344 80 0 FreeSans 320 0 0 0 N2END[5]
port 114 nsew signal input
flabel metal3 s 14456 0 14536 80 0 FreeSans 320 0 0 0 N2END[6]
port 115 nsew signal input
flabel metal3 s 14648 0 14728 80 0 FreeSans 320 0 0 0 N2END[7]
port 116 nsew signal input
flabel metal3 s 11768 0 11848 80 0 FreeSans 320 0 0 0 N2MID[0]
port 117 nsew signal input
flabel metal3 s 11960 0 12040 80 0 FreeSans 320 0 0 0 N2MID[1]
port 118 nsew signal input
flabel metal3 s 12152 0 12232 80 0 FreeSans 320 0 0 0 N2MID[2]
port 119 nsew signal input
flabel metal3 s 12344 0 12424 80 0 FreeSans 320 0 0 0 N2MID[3]
port 120 nsew signal input
flabel metal3 s 12536 0 12616 80 0 FreeSans 320 0 0 0 N2MID[4]
port 121 nsew signal input
flabel metal3 s 12728 0 12808 80 0 FreeSans 320 0 0 0 N2MID[5]
port 122 nsew signal input
flabel metal3 s 12920 0 13000 80 0 FreeSans 320 0 0 0 N2MID[6]
port 123 nsew signal input
flabel metal3 s 13112 0 13192 80 0 FreeSans 320 0 0 0 N2MID[7]
port 124 nsew signal input
flabel metal3 s 14840 0 14920 80 0 FreeSans 320 0 0 0 N4END[0]
port 125 nsew signal input
flabel metal3 s 16760 0 16840 80 0 FreeSans 320 0 0 0 N4END[10]
port 126 nsew signal input
flabel metal3 s 16952 0 17032 80 0 FreeSans 320 0 0 0 N4END[11]
port 127 nsew signal input
flabel metal3 s 17144 0 17224 80 0 FreeSans 320 0 0 0 N4END[12]
port 128 nsew signal input
flabel metal3 s 17336 0 17416 80 0 FreeSans 320 0 0 0 N4END[13]
port 129 nsew signal input
flabel metal3 s 17528 0 17608 80 0 FreeSans 320 0 0 0 N4END[14]
port 130 nsew signal input
flabel metal3 s 17720 0 17800 80 0 FreeSans 320 0 0 0 N4END[15]
port 131 nsew signal input
flabel metal3 s 15032 0 15112 80 0 FreeSans 320 0 0 0 N4END[1]
port 132 nsew signal input
flabel metal3 s 15224 0 15304 80 0 FreeSans 320 0 0 0 N4END[2]
port 133 nsew signal input
flabel metal3 s 15416 0 15496 80 0 FreeSans 320 0 0 0 N4END[3]
port 134 nsew signal input
flabel metal3 s 15608 0 15688 80 0 FreeSans 320 0 0 0 N4END[4]
port 135 nsew signal input
flabel metal3 s 15800 0 15880 80 0 FreeSans 320 0 0 0 N4END[5]
port 136 nsew signal input
flabel metal3 s 15992 0 16072 80 0 FreeSans 320 0 0 0 N4END[6]
port 137 nsew signal input
flabel metal3 s 16184 0 16264 80 0 FreeSans 320 0 0 0 N4END[7]
port 138 nsew signal input
flabel metal3 s 16376 0 16456 80 0 FreeSans 320 0 0 0 N4END[8]
port 139 nsew signal input
flabel metal3 s 16568 0 16648 80 0 FreeSans 320 0 0 0 N4END[9]
port 140 nsew signal input
flabel metal3 s 17912 0 17992 80 0 FreeSans 320 0 0 0 NN4END[0]
port 141 nsew signal input
flabel metal3 s 19832 0 19912 80 0 FreeSans 320 0 0 0 NN4END[10]
port 142 nsew signal input
flabel metal3 s 20024 0 20104 80 0 FreeSans 320 0 0 0 NN4END[11]
port 143 nsew signal input
flabel metal3 s 20216 0 20296 80 0 FreeSans 320 0 0 0 NN4END[12]
port 144 nsew signal input
flabel metal3 s 20408 0 20488 80 0 FreeSans 320 0 0 0 NN4END[13]
port 145 nsew signal input
flabel metal3 s 20600 0 20680 80 0 FreeSans 320 0 0 0 NN4END[14]
port 146 nsew signal input
flabel metal3 s 20792 0 20872 80 0 FreeSans 320 0 0 0 NN4END[15]
port 147 nsew signal input
flabel metal3 s 18104 0 18184 80 0 FreeSans 320 0 0 0 NN4END[1]
port 148 nsew signal input
flabel metal3 s 18296 0 18376 80 0 FreeSans 320 0 0 0 NN4END[2]
port 149 nsew signal input
flabel metal3 s 18488 0 18568 80 0 FreeSans 320 0 0 0 NN4END[3]
port 150 nsew signal input
flabel metal3 s 18680 0 18760 80 0 FreeSans 320 0 0 0 NN4END[4]
port 151 nsew signal input
flabel metal3 s 18872 0 18952 80 0 FreeSans 320 0 0 0 NN4END[5]
port 152 nsew signal input
flabel metal3 s 19064 0 19144 80 0 FreeSans 320 0 0 0 NN4END[6]
port 153 nsew signal input
flabel metal3 s 19256 0 19336 80 0 FreeSans 320 0 0 0 NN4END[7]
port 154 nsew signal input
flabel metal3 s 19448 0 19528 80 0 FreeSans 320 0 0 0 NN4END[8]
port 155 nsew signal input
flabel metal3 s 19640 0 19720 80 0 FreeSans 320 0 0 0 NN4END[9]
port 156 nsew signal input
flabel metal3 s 21176 0 21256 80 0 FreeSans 320 0 0 0 S1BEG[0]
port 157 nsew signal output
flabel metal3 s 21368 0 21448 80 0 FreeSans 320 0 0 0 S1BEG[1]
port 158 nsew signal output
flabel metal3 s 21560 0 21640 80 0 FreeSans 320 0 0 0 S1BEG[2]
port 159 nsew signal output
flabel metal3 s 21752 0 21832 80 0 FreeSans 320 0 0 0 S1BEG[3]
port 160 nsew signal output
flabel metal3 s 21944 0 22024 80 0 FreeSans 320 0 0 0 S2BEG[0]
port 161 nsew signal output
flabel metal3 s 22136 0 22216 80 0 FreeSans 320 0 0 0 S2BEG[1]
port 162 nsew signal output
flabel metal3 s 22328 0 22408 80 0 FreeSans 320 0 0 0 S2BEG[2]
port 163 nsew signal output
flabel metal3 s 22520 0 22600 80 0 FreeSans 320 0 0 0 S2BEG[3]
port 164 nsew signal output
flabel metal3 s 22712 0 22792 80 0 FreeSans 320 0 0 0 S2BEG[4]
port 165 nsew signal output
flabel metal3 s 22904 0 22984 80 0 FreeSans 320 0 0 0 S2BEG[5]
port 166 nsew signal output
flabel metal3 s 23096 0 23176 80 0 FreeSans 320 0 0 0 S2BEG[6]
port 167 nsew signal output
flabel metal3 s 23288 0 23368 80 0 FreeSans 320 0 0 0 S2BEG[7]
port 168 nsew signal output
flabel metal3 s 23480 0 23560 80 0 FreeSans 320 0 0 0 S2BEGb[0]
port 169 nsew signal output
flabel metal3 s 23672 0 23752 80 0 FreeSans 320 0 0 0 S2BEGb[1]
port 170 nsew signal output
flabel metal3 s 23864 0 23944 80 0 FreeSans 320 0 0 0 S2BEGb[2]
port 171 nsew signal output
flabel metal3 s 24056 0 24136 80 0 FreeSans 320 0 0 0 S2BEGb[3]
port 172 nsew signal output
flabel metal3 s 24248 0 24328 80 0 FreeSans 320 0 0 0 S2BEGb[4]
port 173 nsew signal output
flabel metal3 s 24440 0 24520 80 0 FreeSans 320 0 0 0 S2BEGb[5]
port 174 nsew signal output
flabel metal3 s 24632 0 24712 80 0 FreeSans 320 0 0 0 S2BEGb[6]
port 175 nsew signal output
flabel metal3 s 24824 0 24904 80 0 FreeSans 320 0 0 0 S2BEGb[7]
port 176 nsew signal output
flabel metal3 s 25016 0 25096 80 0 FreeSans 320 0 0 0 S4BEG[0]
port 177 nsew signal output
flabel metal3 s 26936 0 27016 80 0 FreeSans 320 0 0 0 S4BEG[10]
port 178 nsew signal output
flabel metal3 s 27128 0 27208 80 0 FreeSans 320 0 0 0 S4BEG[11]
port 179 nsew signal output
flabel metal3 s 27320 0 27400 80 0 FreeSans 320 0 0 0 S4BEG[12]
port 180 nsew signal output
flabel metal3 s 27512 0 27592 80 0 FreeSans 320 0 0 0 S4BEG[13]
port 181 nsew signal output
flabel metal3 s 27704 0 27784 80 0 FreeSans 320 0 0 0 S4BEG[14]
port 182 nsew signal output
flabel metal3 s 27896 0 27976 80 0 FreeSans 320 0 0 0 S4BEG[15]
port 183 nsew signal output
flabel metal3 s 25208 0 25288 80 0 FreeSans 320 0 0 0 S4BEG[1]
port 184 nsew signal output
flabel metal3 s 25400 0 25480 80 0 FreeSans 320 0 0 0 S4BEG[2]
port 185 nsew signal output
flabel metal3 s 25592 0 25672 80 0 FreeSans 320 0 0 0 S4BEG[3]
port 186 nsew signal output
flabel metal3 s 25784 0 25864 80 0 FreeSans 320 0 0 0 S4BEG[4]
port 187 nsew signal output
flabel metal3 s 25976 0 26056 80 0 FreeSans 320 0 0 0 S4BEG[5]
port 188 nsew signal output
flabel metal3 s 26168 0 26248 80 0 FreeSans 320 0 0 0 S4BEG[6]
port 189 nsew signal output
flabel metal3 s 26360 0 26440 80 0 FreeSans 320 0 0 0 S4BEG[7]
port 190 nsew signal output
flabel metal3 s 26552 0 26632 80 0 FreeSans 320 0 0 0 S4BEG[8]
port 191 nsew signal output
flabel metal3 s 26744 0 26824 80 0 FreeSans 320 0 0 0 S4BEG[9]
port 192 nsew signal output
flabel metal3 s 28088 0 28168 80 0 FreeSans 320 0 0 0 SS4BEG[0]
port 193 nsew signal output
flabel metal3 s 30008 0 30088 80 0 FreeSans 320 0 0 0 SS4BEG[10]
port 194 nsew signal output
flabel metal3 s 30200 0 30280 80 0 FreeSans 320 0 0 0 SS4BEG[11]
port 195 nsew signal output
flabel metal3 s 30392 0 30472 80 0 FreeSans 320 0 0 0 SS4BEG[12]
port 196 nsew signal output
flabel metal3 s 30584 0 30664 80 0 FreeSans 320 0 0 0 SS4BEG[13]
port 197 nsew signal output
flabel metal3 s 30776 0 30856 80 0 FreeSans 320 0 0 0 SS4BEG[14]
port 198 nsew signal output
flabel metal3 s 30968 0 31048 80 0 FreeSans 320 0 0 0 SS4BEG[15]
port 199 nsew signal output
flabel metal3 s 28280 0 28360 80 0 FreeSans 320 0 0 0 SS4BEG[1]
port 200 nsew signal output
flabel metal3 s 28472 0 28552 80 0 FreeSans 320 0 0 0 SS4BEG[2]
port 201 nsew signal output
flabel metal3 s 28664 0 28744 80 0 FreeSans 320 0 0 0 SS4BEG[3]
port 202 nsew signal output
flabel metal3 s 28856 0 28936 80 0 FreeSans 320 0 0 0 SS4BEG[4]
port 203 nsew signal output
flabel metal3 s 29048 0 29128 80 0 FreeSans 320 0 0 0 SS4BEG[5]
port 204 nsew signal output
flabel metal3 s 29240 0 29320 80 0 FreeSans 320 0 0 0 SS4BEG[6]
port 205 nsew signal output
flabel metal3 s 29432 0 29512 80 0 FreeSans 320 0 0 0 SS4BEG[7]
port 206 nsew signal output
flabel metal3 s 29624 0 29704 80 0 FreeSans 320 0 0 0 SS4BEG[8]
port 207 nsew signal output
flabel metal3 s 29816 0 29896 80 0 FreeSans 320 0 0 0 SS4BEG[9]
port 208 nsew signal output
flabel metal3 s 31160 0 31240 80 0 FreeSans 320 0 0 0 UserCLK
port 209 nsew signal input
flabel metal3 s 1976 12100 2056 12180 0 FreeSans 320 0 0 0 UserCLKo
port 210 nsew signal output
flabel metal5 s 4892 0 5332 12180 0 FreeSans 2560 90 0 0 VGND
port 211 nsew ground bidirectional
flabel metal5 s 4892 0 5332 40 0 FreeSans 320 0 0 0 VGND
port 211 nsew ground bidirectional
flabel metal5 s 4892 12140 5332 12180 0 FreeSans 320 0 0 0 VGND
port 211 nsew ground bidirectional
flabel metal5 s 20012 0 20452 12180 0 FreeSans 2560 90 0 0 VGND
port 211 nsew ground bidirectional
flabel metal5 s 20012 0 20452 40 0 FreeSans 320 0 0 0 VGND
port 211 nsew ground bidirectional
flabel metal5 s 20012 12140 20452 12180 0 FreeSans 320 0 0 0 VGND
port 211 nsew ground bidirectional
flabel metal5 s 35132 0 35572 12180 0 FreeSans 2560 90 0 0 VGND
port 211 nsew ground bidirectional
flabel metal5 s 35132 0 35572 40 0 FreeSans 320 0 0 0 VGND
port 211 nsew ground bidirectional
flabel metal5 s 35132 12140 35572 12180 0 FreeSans 320 0 0 0 VGND
port 211 nsew ground bidirectional
flabel metal5 s 3652 0 4092 12180 0 FreeSans 2560 90 0 0 VPWR
port 212 nsew power bidirectional
flabel metal5 s 3652 0 4092 40 0 FreeSans 320 0 0 0 VPWR
port 212 nsew power bidirectional
flabel metal5 s 3652 12140 4092 12180 0 FreeSans 320 0 0 0 VPWR
port 212 nsew power bidirectional
flabel metal5 s 18772 0 19212 12180 0 FreeSans 2560 90 0 0 VPWR
port 212 nsew power bidirectional
flabel metal5 s 18772 0 19212 40 0 FreeSans 320 0 0 0 VPWR
port 212 nsew power bidirectional
flabel metal5 s 18772 12140 19212 12180 0 FreeSans 320 0 0 0 VPWR
port 212 nsew power bidirectional
flabel metal5 s 33892 0 34332 12180 0 FreeSans 2560 90 0 0 VPWR
port 212 nsew power bidirectional
flabel metal5 s 33892 0 34332 40 0 FreeSans 320 0 0 0 VPWR
port 212 nsew power bidirectional
flabel metal5 s 33892 12140 34332 12180 0 FreeSans 320 0 0 0 VPWR
port 212 nsew power bidirectional
rlabel metal1 23184 10584 23184 10584 0 VGND
rlabel metal1 23184 9828 23184 9828 0 VPWR
rlabel metal2 272 756 272 756 0 FrameData[0]
rlabel metal2 560 4116 560 4116 0 FrameData[10]
rlabel metal2 752 4452 752 4452 0 FrameData[11]
rlabel metal2 34992 2856 34992 2856 0 FrameData[12]
rlabel metal2 704 5124 704 5124 0 FrameData[13]
rlabel metal2 464 5460 464 5460 0 FrameData[14]
rlabel metal2 560 5796 560 5796 0 FrameData[15]
rlabel metal2 320 6132 320 6132 0 FrameData[16]
rlabel metal2 512 6468 512 6468 0 FrameData[17]
rlabel metal2 608 6804 608 6804 0 FrameData[18]
rlabel metal2 752 7140 752 7140 0 FrameData[19]
rlabel metal2 4112 1092 4112 1092 0 FrameData[1]
rlabel metal2 17952 7728 17952 7728 0 FrameData[20]
rlabel metal2 23040 8694 23040 8694 0 FrameData[21]
rlabel metal2 704 8148 704 8148 0 FrameData[22]
rlabel metal2 21600 8568 21600 8568 0 FrameData[23]
rlabel metal2 24192 8736 24192 8736 0 FrameData[24]
rlabel metal3 23616 8904 23616 8904 0 FrameData[25]
rlabel metal2 656 9492 656 9492 0 FrameData[26]
rlabel metal3 22464 9198 22464 9198 0 FrameData[27]
rlabel metal2 128 10164 128 10164 0 FrameData[28]
rlabel metal2 16992 10668 16992 10668 0 FrameData[29]
rlabel metal2 752 1428 752 1428 0 FrameData[2]
rlabel metal3 21504 9786 21504 9786 0 FrameData[30]
rlabel metal2 224 11172 224 11172 0 FrameData[31]
rlabel metal2 752 1764 752 1764 0 FrameData[3]
rlabel metal2 416 2100 416 2100 0 FrameData[4]
rlabel metal2 752 2436 752 2436 0 FrameData[5]
rlabel metal2 752 2772 752 2772 0 FrameData[6]
rlabel metal2 30048 5544 30048 5544 0 FrameData[7]
rlabel metal2 38400 4662 38400 4662 0 FrameData[8]
rlabel metal3 19296 3864 19296 3864 0 FrameData[9]
rlabel metal2 45855 756 45855 756 0 FrameData_O[0]
rlabel metal2 45951 4116 45951 4116 0 FrameData_O[10]
rlabel metal2 45168 4368 45168 4368 0 FrameData_O[11]
rlabel metal2 45543 4788 45543 4788 0 FrameData_O[12]
rlabel metal2 45735 5124 45735 5124 0 FrameData_O[13]
rlabel metal2 45951 5460 45951 5460 0 FrameData_O[14]
rlabel metal2 45735 5796 45735 5796 0 FrameData_O[15]
rlabel metal2 45543 6132 45543 6132 0 FrameData_O[16]
rlabel metal2 45735 6468 45735 6468 0 FrameData_O[17]
rlabel via2 46287 6804 46287 6804 0 FrameData_O[18]
rlabel metal2 45735 7140 45735 7140 0 FrameData_O[19]
rlabel metal2 45471 1092 45471 1092 0 FrameData_O[1]
rlabel via2 46287 7476 46287 7476 0 FrameData_O[20]
rlabel metal2 45543 7812 45543 7812 0 FrameData_O[21]
rlabel via2 46287 8148 46287 8148 0 FrameData_O[22]
rlabel metal2 45951 8484 45951 8484 0 FrameData_O[23]
rlabel metal2 46047 8820 46047 8820 0 FrameData_O[24]
rlabel metal2 45543 9156 45543 9156 0 FrameData_O[25]
rlabel metal2 46047 9492 46047 9492 0 FrameData_O[26]
rlabel metal2 45663 9828 45663 9828 0 FrameData_O[27]
rlabel metal2 45711 10164 45711 10164 0 FrameData_O[28]
rlabel metal2 44424 9660 44424 9660 0 FrameData_O[29]
rlabel metal2 45999 1428 45999 1428 0 FrameData_O[2]
rlabel metal2 43800 10416 43800 10416 0 FrameData_O[30]
rlabel metal2 44040 9576 44040 9576 0 FrameData_O[31]
rlabel metal2 45543 1764 45543 1764 0 FrameData_O[3]
rlabel metal2 45735 2100 45735 2100 0 FrameData_O[4]
rlabel metal2 46047 2436 46047 2436 0 FrameData_O[5]
rlabel metal2 45735 2772 45735 2772 0 FrameData_O[6]
rlabel metal2 45543 3108 45543 3108 0 FrameData_O[7]
rlabel metal2 45663 3444 45663 3444 0 FrameData_O[8]
rlabel metal2 45168 3696 45168 3696 0 FrameData_O[9]
rlabel metal3 31392 156 31392 156 0 FrameStrobe[0]
rlabel metal3 33312 1470 33312 1470 0 FrameStrobe[10]
rlabel metal3 33504 1470 33504 1470 0 FrameStrobe[11]
rlabel metal3 33696 996 33696 996 0 FrameStrobe[12]
rlabel metal3 33888 1080 33888 1080 0 FrameStrobe[13]
rlabel metal3 34080 1080 34080 1080 0 FrameStrobe[14]
rlabel metal3 34272 1080 34272 1080 0 FrameStrobe[15]
rlabel metal3 34464 1752 34464 1752 0 FrameStrobe[16]
rlabel metal3 34656 1542 34656 1542 0 FrameStrobe[17]
rlabel metal3 34848 1080 34848 1080 0 FrameStrobe[18]
rlabel metal3 35040 1584 35040 1584 0 FrameStrobe[19]
rlabel metal3 31584 114 31584 114 0 FrameStrobe[1]
rlabel metal3 31776 198 31776 198 0 FrameStrobe[2]
rlabel metal2 13872 8652 13872 8652 0 FrameStrobe[3]
rlabel metal3 19008 9030 19008 9030 0 FrameStrobe[4]
rlabel metal2 29232 9156 29232 9156 0 FrameStrobe[5]
rlabel metal2 32160 8568 32160 8568 0 FrameStrobe[6]
rlabel metal2 32304 8652 32304 8652 0 FrameStrobe[7]
rlabel metal2 32112 8484 32112 8484 0 FrameStrobe[8]
rlabel metal3 33216 2952 33216 2952 0 FrameStrobe[9]
rlabel metal2 4152 10416 4152 10416 0 FrameStrobe_O[0]
rlabel metal2 25272 10416 25272 10416 0 FrameStrobe_O[10]
rlabel metal2 27384 10416 27384 10416 0 FrameStrobe_O[11]
rlabel metal2 29496 10416 29496 10416 0 FrameStrobe_O[12]
rlabel metal2 31608 10416 31608 10416 0 FrameStrobe_O[13]
rlabel metal2 33720 10416 33720 10416 0 FrameStrobe_O[14]
rlabel metal2 35832 10416 35832 10416 0 FrameStrobe_O[15]
rlabel metal2 37944 10416 37944 10416 0 FrameStrobe_O[16]
rlabel metal2 40056 10416 40056 10416 0 FrameStrobe_O[17]
rlabel metal2 42168 10416 42168 10416 0 FrameStrobe_O[18]
rlabel metal2 44280 10416 44280 10416 0 FrameStrobe_O[19]
rlabel metal2 6264 10416 6264 10416 0 FrameStrobe_O[1]
rlabel metal2 8376 10416 8376 10416 0 FrameStrobe_O[2]
rlabel metal2 10488 10416 10488 10416 0 FrameStrobe_O[3]
rlabel metal2 12600 10416 12600 10416 0 FrameStrobe_O[4]
rlabel metal2 14712 10416 14712 10416 0 FrameStrobe_O[5]
rlabel metal2 16824 10416 16824 10416 0 FrameStrobe_O[6]
rlabel metal2 18936 10416 18936 10416 0 FrameStrobe_O[7]
rlabel metal2 21048 10416 21048 10416 0 FrameStrobe_O[8]
rlabel metal2 23160 10416 23160 10416 0 FrameStrobe_O[9]
rlabel metal2 9072 4116 9072 4116 0 N1END[0]
rlabel metal2 9216 4368 9216 4368 0 N1END[1]
rlabel metal2 9504 4452 9504 4452 0 N1END[2]
rlabel metal2 9984 4956 9984 4956 0 N1END[3]
rlabel metal3 13344 3264 13344 3264 0 N2END[0]
rlabel metal3 13536 3600 13536 3600 0 N2END[1]
rlabel metal2 13824 7140 13824 7140 0 N2END[2]
rlabel metal2 14448 7056 14448 7056 0 N2END[3]
rlabel metal2 14592 6888 14592 6888 0 N2END[4]
rlabel metal2 15264 6804 15264 6804 0 N2END[5]
rlabel metal2 15792 6720 15792 6720 0 N2END[6]
rlabel metal2 16224 6552 16224 6552 0 N2END[7]
rlabel metal3 11808 1332 11808 1332 0 N2MID[0]
rlabel metal3 12000 1374 12000 1374 0 N2MID[1]
rlabel metal3 12192 1416 12192 1416 0 N2MID[2]
rlabel metal3 12384 1458 12384 1458 0 N2MID[3]
rlabel metal2 11712 4620 11712 4620 0 N2MID[4]
rlabel metal3 12672 4788 12672 4788 0 N2MID[5]
rlabel metal3 12960 240 12960 240 0 N2MID[6]
rlabel metal2 13344 5628 13344 5628 0 N2MID[7]
rlabel metal2 15552 7980 15552 7980 0 N4END[0]
rlabel metal2 18048 6468 18048 6468 0 N4END[10]
rlabel metal2 18336 6384 18336 6384 0 N4END[11]
rlabel metal2 18528 6048 18528 6048 0 N4END[12]
rlabel metal2 19296 5796 19296 5796 0 N4END[13]
rlabel metal2 19152 5880 19152 5880 0 N4END[14]
rlabel metal2 19008 6216 19008 6216 0 N4END[15]
rlabel metal2 15840 7896 15840 7896 0 N4END[1]
rlabel metal2 15984 8148 15984 8148 0 N4END[2]
rlabel metal2 16416 7224 16416 7224 0 N4END[3]
rlabel metal2 16704 8232 16704 8232 0 N4END[4]
rlabel metal2 17232 8316 17232 8316 0 N4END[5]
rlabel metal2 16368 7812 16368 7812 0 N4END[6]
rlabel metal3 16224 240 16224 240 0 N4END[7]
rlabel metal2 17328 6804 17328 6804 0 N4END[8]
rlabel metal2 17664 6636 17664 6636 0 N4END[9]
rlabel metal3 17952 2340 17952 2340 0 NN4END[0]
rlabel metal2 20976 4956 20976 4956 0 NN4END[10]
rlabel metal3 20064 702 20064 702 0 NN4END[11]
rlabel metal3 20256 702 20256 702 0 NN4END[12]
rlabel metal3 20448 702 20448 702 0 NN4END[13]
rlabel metal3 20496 6552 20496 6552 0 NN4END[14]
rlabel metal2 20400 6384 20400 6384 0 NN4END[15]
rlabel metal3 18144 2466 18144 2466 0 NN4END[1]
rlabel metal2 20592 4368 20592 4368 0 NN4END[2]
rlabel metal3 26208 3528 26208 3528 0 NN4END[3]
rlabel metal3 18720 1248 18720 1248 0 NN4END[4]
rlabel metal3 18912 702 18912 702 0 NN4END[5]
rlabel metal3 19104 786 19104 786 0 NN4END[6]
rlabel metal4 19440 3612 19440 3612 0 NN4END[7]
rlabel metal2 21216 4620 21216 4620 0 NN4END[8]
rlabel metal2 21120 4872 21120 4872 0 NN4END[9]
rlabel metal3 21216 1248 21216 1248 0 S1BEG[0]
rlabel metal3 21408 870 21408 870 0 S1BEG[1]
rlabel metal3 21600 1248 21600 1248 0 S1BEG[2]
rlabel metal3 21792 870 21792 870 0 S1BEG[3]
rlabel metal3 21984 1248 21984 1248 0 S2BEG[0]
rlabel metal3 22176 870 22176 870 0 S2BEG[1]
rlabel metal3 22368 1248 22368 1248 0 S2BEG[2]
rlabel metal3 22560 870 22560 870 0 S2BEG[3]
rlabel metal3 22752 1248 22752 1248 0 S2BEG[4]
rlabel metal3 22944 870 22944 870 0 S2BEG[5]
rlabel metal3 23136 1248 23136 1248 0 S2BEG[6]
rlabel metal3 23328 870 23328 870 0 S2BEG[7]
rlabel metal3 23520 1248 23520 1248 0 S2BEGb[0]
rlabel metal3 23712 870 23712 870 0 S2BEGb[1]
rlabel metal3 23904 870 23904 870 0 S2BEGb[2]
rlabel metal3 24096 912 24096 912 0 S2BEGb[3]
rlabel metal3 24288 870 24288 870 0 S2BEGb[4]
rlabel metal3 24480 870 24480 870 0 S2BEGb[5]
rlabel metal3 24672 912 24672 912 0 S2BEGb[6]
rlabel metal3 24864 870 24864 870 0 S2BEGb[7]
rlabel metal3 25056 828 25056 828 0 S4BEG[0]
rlabel metal3 26976 912 26976 912 0 S4BEG[10]
rlabel metal3 27168 1248 27168 1248 0 S4BEG[11]
rlabel metal3 27360 828 27360 828 0 S4BEG[12]
rlabel metal3 27552 1248 27552 1248 0 S4BEG[13]
rlabel metal3 27744 828 27744 828 0 S4BEG[14]
rlabel metal3 27936 1248 27936 1248 0 S4BEG[15]
rlabel metal3 25248 1248 25248 1248 0 S4BEG[1]
rlabel metal3 25440 912 25440 912 0 S4BEG[2]
rlabel metal3 25632 1248 25632 1248 0 S4BEG[3]
rlabel metal3 25824 828 25824 828 0 S4BEG[4]
rlabel metal3 26016 1248 26016 1248 0 S4BEG[5]
rlabel metal3 26208 1038 26208 1038 0 S4BEG[6]
rlabel metal3 26400 1248 26400 1248 0 S4BEG[7]
rlabel metal3 26592 828 26592 828 0 S4BEG[8]
rlabel metal3 26784 1248 26784 1248 0 S4BEG[9]
rlabel metal3 28128 912 28128 912 0 SS4BEG[0]
rlabel metal3 30048 912 30048 912 0 SS4BEG[10]
rlabel metal3 30240 1248 30240 1248 0 SS4BEG[11]
rlabel metal3 30432 828 30432 828 0 SS4BEG[12]
rlabel metal3 30624 1248 30624 1248 0 SS4BEG[13]
rlabel metal3 30816 828 30816 828 0 SS4BEG[14]
rlabel metal3 31008 1248 31008 1248 0 SS4BEG[15]
rlabel metal3 28320 1248 28320 1248 0 SS4BEG[1]
rlabel metal3 28512 828 28512 828 0 SS4BEG[2]
rlabel metal3 28704 1248 28704 1248 0 SS4BEG[3]
rlabel metal3 28896 828 28896 828 0 SS4BEG[4]
rlabel metal3 29088 1248 29088 1248 0 SS4BEG[5]
rlabel metal3 29280 1038 29280 1038 0 SS4BEG[6]
rlabel metal3 29472 1248 29472 1248 0 SS4BEG[7]
rlabel metal3 29664 828 29664 828 0 SS4BEG[8]
rlabel metal3 29856 1248 29856 1248 0 SS4BEG[9]
rlabel via3 31200 72 31200 72 0 UserCLK
rlabel metal2 2040 10416 2040 10416 0 UserCLKo
rlabel metal2 42960 2016 42960 2016 0 net1
rlabel metal2 26664 3192 26664 3192 0 net10
rlabel metal2 22296 4956 22296 4956 0 net100
rlabel metal2 29616 2100 29616 2100 0 net101
rlabel metal2 28896 2688 28896 2688 0 net102
rlabel metal2 28848 4368 28848 4368 0 net103
rlabel metal4 26928 2856 26928 2856 0 net104
rlabel metal2 2304 10122 2304 10122 0 net105
rlabel metal2 34560 4956 34560 4956 0 net11
rlabel metal2 41424 1932 41424 1932 0 net12
rlabel metal2 26400 7686 26400 7686 0 net13
rlabel metal2 38016 9114 38016 9114 0 net14
rlabel metal3 38016 8988 38016 8988 0 net15
rlabel metal3 38112 9114 38112 9114 0 net16
rlabel metal2 24504 8820 24504 8820 0 net17
rlabel metal3 38208 9156 38208 9156 0 net18
rlabel metal3 31008 7938 31008 7938 0 net19
rlabel metal3 44544 3864 44544 3864 0 net2
rlabel metal2 22680 8568 22680 8568 0 net20
rlabel metal2 38112 9366 38112 9366 0 net21
rlabel metal2 44160 9576 44160 9576 0 net22
rlabel metal2 40992 5544 40992 5544 0 net23
rlabel metal2 22488 8904 22488 8904 0 net24
rlabel metal3 27840 7896 27840 7896 0 net25
rlabel metal2 44496 1932 44496 1932 0 net26
rlabel metal2 44832 1932 44832 1932 0 net27
rlabel metal3 44448 4116 44448 4116 0 net28
rlabel metal2 44928 2646 44928 2646 0 net29
rlabel metal3 44928 3696 44928 3696 0 net3
rlabel metal3 41088 4284 41088 4284 0 net30
rlabel metal3 41280 4494 41280 4494 0 net31
rlabel metal2 44928 3654 44928 3654 0 net32
rlabel metal2 6600 8652 6600 8652 0 net33
rlabel metal2 27288 8904 27288 8904 0 net34
rlabel metal2 27864 8904 27864 8904 0 net35
rlabel metal2 28776 8904 28776 8904 0 net36
rlabel metal2 28104 8148 28104 8148 0 net37
rlabel metal2 28872 8148 28872 8148 0 net38
rlabel metal3 34560 8400 34560 8400 0 net39
rlabel metal2 35544 3444 35544 3444 0 net4
rlabel metal3 35616 7140 35616 7140 0 net40
rlabel metal2 26856 3612 26856 3612 0 net41
rlabel metal3 42432 10500 42432 10500 0 net42
rlabel metal2 38304 10164 38304 10164 0 net43
rlabel metal2 6360 8904 6360 8904 0 net44
rlabel metal2 7944 8652 7944 8652 0 net45
rlabel metal2 13080 8904 13080 8904 0 net46
rlabel metal2 17880 8904 17880 8904 0 net47
rlabel metal2 19296 10164 19296 10164 0 net48
rlabel metal3 17088 10458 17088 10458 0 net49
rlabel metal2 37824 3486 37824 3486 0 net5
rlabel metal3 19200 10416 19200 10416 0 net50
rlabel metal2 29112 8904 29112 8904 0 net51
rlabel metal2 26904 8904 26904 8904 0 net52
rlabel metal3 15168 3654 15168 3654 0 net53
rlabel metal2 19584 1932 19584 1932 0 net54
rlabel metal2 21888 2646 21888 2646 0 net55
rlabel metal3 18672 2520 18672 2520 0 net56
rlabel metal2 21600 2520 21600 2520 0 net57
rlabel metal3 21696 3318 21696 3318 0 net58
rlabel metal4 20976 5628 20976 5628 0 net59
rlabel metal2 27432 3612 27432 3612 0 net6
rlabel metal2 21744 2016 21744 2016 0 net60
rlabel metal2 22944 2478 22944 2478 0 net61
rlabel metal2 19200 2100 19200 2100 0 net62
rlabel metal2 23424 2688 23424 2688 0 net63
rlabel metal3 22848 2394 22848 2394 0 net64
rlabel metal3 22944 2952 22944 2952 0 net65
rlabel metal2 21744 6468 21744 6468 0 net66
rlabel metal3 17472 6552 17472 6552 0 net67
rlabel metal2 19680 6804 19680 6804 0 net68
rlabel metal3 16224 2532 16224 2532 0 net69
rlabel metal2 39168 4914 39168 4914 0 net7
rlabel metal2 21264 6048 21264 6048 0 net70
rlabel metal4 18960 2604 18960 2604 0 net71
rlabel metal2 19632 2520 19632 2520 0 net72
rlabel metal2 24048 2352 24048 2352 0 net73
rlabel metal2 27360 2100 27360 2100 0 net74
rlabel metal2 19272 8148 19272 8148 0 net75
rlabel metal3 17856 7602 17856 7602 0 net76
rlabel metal3 17472 7560 17472 7560 0 net77
rlabel metal2 17352 8148 17352 8148 0 net78
rlabel metal3 17088 7518 17088 7518 0 net79
rlabel metal2 28536 3444 28536 3444 0 net8
rlabel metal2 21504 7182 21504 7182 0 net80
rlabel metal2 25440 1512 25440 1512 0 net81
rlabel metal2 20928 6930 20928 6930 0 net82
rlabel metal3 19968 6468 19968 6468 0 net83
rlabel metal2 19776 6888 19776 6888 0 net84
rlabel metal3 19392 6804 19392 6804 0 net85
rlabel metal3 21024 6594 21024 6594 0 net86
rlabel metal2 20928 6342 20928 6342 0 net87
rlabel metal2 18912 7686 18912 7686 0 net88
rlabel metal4 25776 2016 25776 2016 0 net89
rlabel metal2 35232 3192 35232 3192 0 net9
rlabel metal4 26736 2184 26736 2184 0 net90
rlabel metal2 30528 2562 30528 2562 0 net91
rlabel metal2 30000 1848 30000 1848 0 net92
rlabel metal2 30576 2688 30576 2688 0 net93
rlabel metal2 31776 1932 31776 1932 0 net94
rlabel metal2 30024 4704 30024 4704 0 net95
rlabel metal4 26256 2604 26256 2604 0 net96
rlabel metal3 29568 3612 29568 3612 0 net97
rlabel metal2 25320 5544 25320 5544 0 net98
rlabel metal2 25992 5628 25992 5628 0 net99
<< properties >>
string FIXED_BBOX 0 0 46368 12180
<< end >>
