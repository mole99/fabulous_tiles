module N_term_single2 (UserCLK,
    UserCLKo,
    FrameData,
    FrameData_O,
    FrameStrobe,
    FrameStrobe_O,
    N1END,
    N2END,
    N2MID,
    N4END,
    NN4END,
    S1BEG,
    S2BEG,
    S2BEGb,
    S4BEG,
    SS4BEG);
 input UserCLK;
 output UserCLKo;
 input [31:0] FrameData;
 output [31:0] FrameData_O;
 input [19:0] FrameStrobe;
 output [19:0] FrameStrobe_O;
 input [3:0] N1END;
 input [7:0] N2END;
 input [7:0] N2MID;
 input [15:0] N4END;
 input [15:0] NN4END;
 output [3:0] S1BEG;
 output [7:0] S2BEG;
 output [7:0] S2BEGb;
 output [15:0] S4BEG;
 output [15:0] SS4BEG;

 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;

 sg13g2_buf_1 _000_ (.A(FrameData[0]),
    .X(net1));
 sg13g2_buf_1 _001_ (.A(FrameData[1]),
    .X(net12));
 sg13g2_buf_1 _002_ (.A(FrameData[2]),
    .X(net23));
 sg13g2_buf_1 _003_ (.A(FrameData[3]),
    .X(net26));
 sg13g2_buf_1 _004_ (.A(FrameData[4]),
    .X(net27));
 sg13g2_buf_1 _005_ (.A(FrameData[5]),
    .X(net28));
 sg13g2_buf_1 _006_ (.A(FrameData[6]),
    .X(net29));
 sg13g2_buf_1 _007_ (.A(FrameData[7]),
    .X(net30));
 sg13g2_buf_1 _008_ (.A(FrameData[8]),
    .X(net31));
 sg13g2_buf_1 _009_ (.A(FrameData[9]),
    .X(net32));
 sg13g2_buf_1 _010_ (.A(FrameData[10]),
    .X(net2));
 sg13g2_buf_1 _011_ (.A(FrameData[11]),
    .X(net3));
 sg13g2_buf_1 _012_ (.A(FrameData[12]),
    .X(net4));
 sg13g2_buf_1 _013_ (.A(FrameData[13]),
    .X(net5));
 sg13g2_buf_1 _014_ (.A(FrameData[14]),
    .X(net6));
 sg13g2_buf_1 _015_ (.A(FrameData[15]),
    .X(net7));
 sg13g2_buf_1 _016_ (.A(FrameData[16]),
    .X(net8));
 sg13g2_buf_1 _017_ (.A(FrameData[17]),
    .X(net9));
 sg13g2_buf_1 _018_ (.A(FrameData[18]),
    .X(net10));
 sg13g2_buf_1 _019_ (.A(FrameData[19]),
    .X(net11));
 sg13g2_buf_1 _020_ (.A(FrameData[20]),
    .X(net13));
 sg13g2_buf_1 _021_ (.A(FrameData[21]),
    .X(net14));
 sg13g2_buf_1 _022_ (.A(FrameData[22]),
    .X(net15));
 sg13g2_buf_1 _023_ (.A(FrameData[23]),
    .X(net16));
 sg13g2_buf_1 _024_ (.A(FrameData[24]),
    .X(net17));
 sg13g2_buf_1 _025_ (.A(FrameData[25]),
    .X(net18));
 sg13g2_buf_1 _026_ (.A(FrameData[26]),
    .X(net19));
 sg13g2_buf_1 _027_ (.A(FrameData[27]),
    .X(net20));
 sg13g2_buf_1 _028_ (.A(FrameData[28]),
    .X(net21));
 sg13g2_buf_1 _029_ (.A(FrameData[29]),
    .X(net22));
 sg13g2_buf_1 _030_ (.A(FrameData[30]),
    .X(net24));
 sg13g2_buf_1 _031_ (.A(FrameData[31]),
    .X(net25));
 sg13g2_buf_1 _032_ (.A(FrameStrobe[0]),
    .X(net33));
 sg13g2_buf_1 _033_ (.A(FrameStrobe[1]),
    .X(net44));
 sg13g2_buf_1 _034_ (.A(FrameStrobe[2]),
    .X(net45));
 sg13g2_buf_1 _035_ (.A(FrameStrobe[3]),
    .X(net46));
 sg13g2_buf_1 _036_ (.A(FrameStrobe[4]),
    .X(net47));
 sg13g2_buf_1 _037_ (.A(FrameStrobe[5]),
    .X(net48));
 sg13g2_buf_1 _038_ (.A(FrameStrobe[6]),
    .X(net49));
 sg13g2_buf_1 _039_ (.A(FrameStrobe[7]),
    .X(net50));
 sg13g2_buf_1 _040_ (.A(FrameStrobe[8]),
    .X(net51));
 sg13g2_buf_1 _041_ (.A(FrameStrobe[9]),
    .X(net52));
 sg13g2_buf_1 _042_ (.A(FrameStrobe[10]),
    .X(net34));
 sg13g2_buf_1 _043_ (.A(FrameStrobe[11]),
    .X(net35));
 sg13g2_buf_1 _044_ (.A(FrameStrobe[12]),
    .X(net36));
 sg13g2_buf_1 _045_ (.A(FrameStrobe[13]),
    .X(net37));
 sg13g2_buf_1 _046_ (.A(FrameStrobe[14]),
    .X(net38));
 sg13g2_buf_1 _047_ (.A(FrameStrobe[15]),
    .X(net39));
 sg13g2_buf_1 _048_ (.A(FrameStrobe[16]),
    .X(net40));
 sg13g2_buf_1 _049_ (.A(FrameStrobe[17]),
    .X(net41));
 sg13g2_buf_1 _050_ (.A(FrameStrobe[18]),
    .X(net42));
 sg13g2_buf_1 _051_ (.A(FrameStrobe[19]),
    .X(net43));
 sg13g2_buf_1 _052_ (.A(N1END[3]),
    .X(net53));
 sg13g2_buf_1 _053_ (.A(N1END[2]),
    .X(net54));
 sg13g2_buf_1 _054_ (.A(N1END[1]),
    .X(net55));
 sg13g2_buf_1 _055_ (.A(N1END[0]),
    .X(net56));
 sg13g2_buf_1 _056_ (.A(N2MID[7]),
    .X(net57));
 sg13g2_buf_1 _057_ (.A(N2MID[6]),
    .X(net58));
 sg13g2_buf_1 _058_ (.A(N2MID[5]),
    .X(net59));
 sg13g2_buf_1 _059_ (.A(N2MID[4]),
    .X(net60));
 sg13g2_buf_1 _060_ (.A(N2MID[3]),
    .X(net61));
 sg13g2_buf_1 _061_ (.A(N2MID[2]),
    .X(net62));
 sg13g2_buf_1 _062_ (.A(N2MID[1]),
    .X(net63));
 sg13g2_buf_1 _063_ (.A(N2MID[0]),
    .X(net64));
 sg13g2_buf_1 _064_ (.A(N2END[7]),
    .X(net65));
 sg13g2_buf_1 _065_ (.A(N2END[6]),
    .X(net66));
 sg13g2_buf_1 _066_ (.A(N2END[5]),
    .X(net67));
 sg13g2_buf_1 _067_ (.A(N2END[4]),
    .X(net68));
 sg13g2_buf_1 _068_ (.A(N2END[3]),
    .X(net69));
 sg13g2_buf_1 _069_ (.A(N2END[2]),
    .X(net70));
 sg13g2_buf_1 _070_ (.A(N2END[1]),
    .X(net71));
 sg13g2_buf_1 _071_ (.A(N2END[0]),
    .X(net72));
 sg13g2_buf_1 _072_ (.A(N4END[15]),
    .X(net73));
 sg13g2_buf_1 _073_ (.A(N4END[14]),
    .X(net80));
 sg13g2_buf_1 _074_ (.A(N4END[13]),
    .X(net81));
 sg13g2_buf_1 _075_ (.A(N4END[12]),
    .X(net82));
 sg13g2_buf_1 _076_ (.A(N4END[11]),
    .X(net83));
 sg13g2_buf_1 _077_ (.A(N4END[10]),
    .X(net84));
 sg13g2_buf_1 _078_ (.A(N4END[9]),
    .X(net85));
 sg13g2_buf_1 _079_ (.A(N4END[8]),
    .X(net86));
 sg13g2_buf_1 _080_ (.A(N4END[7]),
    .X(net87));
 sg13g2_buf_1 _081_ (.A(N4END[6]),
    .X(net88));
 sg13g2_buf_1 _082_ (.A(N4END[5]),
    .X(net74));
 sg13g2_buf_1 _083_ (.A(N4END[4]),
    .X(net75));
 sg13g2_buf_1 _084_ (.A(N4END[3]),
    .X(net76));
 sg13g2_buf_1 _085_ (.A(N4END[2]),
    .X(net77));
 sg13g2_buf_1 _086_ (.A(N4END[1]),
    .X(net78));
 sg13g2_buf_1 _087_ (.A(N4END[0]),
    .X(net79));
 sg13g2_buf_1 _088_ (.A(NN4END[15]),
    .X(net89));
 sg13g2_buf_1 _089_ (.A(NN4END[14]),
    .X(net96));
 sg13g2_buf_1 _090_ (.A(NN4END[13]),
    .X(net97));
 sg13g2_buf_1 _091_ (.A(NN4END[12]),
    .X(net98));
 sg13g2_buf_1 _092_ (.A(NN4END[11]),
    .X(net99));
 sg13g2_buf_1 _093_ (.A(NN4END[10]),
    .X(net100));
 sg13g2_buf_1 _094_ (.A(NN4END[9]),
    .X(net101));
 sg13g2_buf_1 _095_ (.A(NN4END[8]),
    .X(net102));
 sg13g2_buf_1 _096_ (.A(NN4END[7]),
    .X(net103));
 sg13g2_buf_1 _097_ (.A(NN4END[6]),
    .X(net104));
 sg13g2_buf_1 _098_ (.A(NN4END[5]),
    .X(net90));
 sg13g2_buf_1 _099_ (.A(NN4END[4]),
    .X(net91));
 sg13g2_buf_1 _100_ (.A(NN4END[3]),
    .X(net92));
 sg13g2_buf_1 _101_ (.A(NN4END[2]),
    .X(net93));
 sg13g2_buf_1 _102_ (.A(NN4END[1]),
    .X(net94));
 sg13g2_buf_1 _103_ (.A(NN4END[0]),
    .X(net95));
 sg13g2_buf_1 _104_ (.A(UserCLK),
    .X(net105));
 sg13g2_buf_1 output1 (.A(net1),
    .X(FrameData_O[0]));
 sg13g2_buf_1 output2 (.A(net2),
    .X(FrameData_O[10]));
 sg13g2_buf_1 output3 (.A(net3),
    .X(FrameData_O[11]));
 sg13g2_buf_1 output4 (.A(net4),
    .X(FrameData_O[12]));
 sg13g2_buf_1 output5 (.A(net5),
    .X(FrameData_O[13]));
 sg13g2_buf_1 output6 (.A(net6),
    .X(FrameData_O[14]));
 sg13g2_buf_1 output7 (.A(net7),
    .X(FrameData_O[15]));
 sg13g2_buf_1 output8 (.A(net8),
    .X(FrameData_O[16]));
 sg13g2_buf_1 output9 (.A(net9),
    .X(FrameData_O[17]));
 sg13g2_buf_1 output10 (.A(net10),
    .X(FrameData_O[18]));
 sg13g2_buf_1 output11 (.A(net11),
    .X(FrameData_O[19]));
 sg13g2_buf_1 output12 (.A(net12),
    .X(FrameData_O[1]));
 sg13g2_buf_1 output13 (.A(net13),
    .X(FrameData_O[20]));
 sg13g2_buf_1 output14 (.A(net14),
    .X(FrameData_O[21]));
 sg13g2_buf_1 output15 (.A(net15),
    .X(FrameData_O[22]));
 sg13g2_buf_1 output16 (.A(net16),
    .X(FrameData_O[23]));
 sg13g2_buf_1 output17 (.A(net17),
    .X(FrameData_O[24]));
 sg13g2_buf_1 output18 (.A(net18),
    .X(FrameData_O[25]));
 sg13g2_buf_1 output19 (.A(net19),
    .X(FrameData_O[26]));
 sg13g2_buf_1 output20 (.A(net20),
    .X(FrameData_O[27]));
 sg13g2_buf_1 output21 (.A(net21),
    .X(FrameData_O[28]));
 sg13g2_buf_1 output22 (.A(net22),
    .X(FrameData_O[29]));
 sg13g2_buf_1 output23 (.A(net23),
    .X(FrameData_O[2]));
 sg13g2_buf_1 output24 (.A(net24),
    .X(FrameData_O[30]));
 sg13g2_buf_1 output25 (.A(net25),
    .X(FrameData_O[31]));
 sg13g2_buf_1 output26 (.A(net26),
    .X(FrameData_O[3]));
 sg13g2_buf_1 output27 (.A(net27),
    .X(FrameData_O[4]));
 sg13g2_buf_1 output28 (.A(net28),
    .X(FrameData_O[5]));
 sg13g2_buf_1 output29 (.A(net29),
    .X(FrameData_O[6]));
 sg13g2_buf_1 output30 (.A(net30),
    .X(FrameData_O[7]));
 sg13g2_buf_1 output31 (.A(net31),
    .X(FrameData_O[8]));
 sg13g2_buf_1 output32 (.A(net32),
    .X(FrameData_O[9]));
 sg13g2_buf_1 output33 (.A(net33),
    .X(FrameStrobe_O[0]));
 sg13g2_buf_1 output34 (.A(net34),
    .X(FrameStrobe_O[10]));
 sg13g2_buf_1 output35 (.A(net35),
    .X(FrameStrobe_O[11]));
 sg13g2_buf_1 output36 (.A(net36),
    .X(FrameStrobe_O[12]));
 sg13g2_buf_1 output37 (.A(net37),
    .X(FrameStrobe_O[13]));
 sg13g2_buf_1 output38 (.A(net38),
    .X(FrameStrobe_O[14]));
 sg13g2_buf_1 output39 (.A(net39),
    .X(FrameStrobe_O[15]));
 sg13g2_buf_1 output40 (.A(net40),
    .X(FrameStrobe_O[16]));
 sg13g2_buf_1 output41 (.A(net41),
    .X(FrameStrobe_O[17]));
 sg13g2_buf_1 output42 (.A(net42),
    .X(FrameStrobe_O[18]));
 sg13g2_buf_1 output43 (.A(net43),
    .X(FrameStrobe_O[19]));
 sg13g2_buf_1 output44 (.A(net44),
    .X(FrameStrobe_O[1]));
 sg13g2_buf_1 output45 (.A(net45),
    .X(FrameStrobe_O[2]));
 sg13g2_buf_1 output46 (.A(net46),
    .X(FrameStrobe_O[3]));
 sg13g2_buf_1 output47 (.A(net47),
    .X(FrameStrobe_O[4]));
 sg13g2_buf_1 output48 (.A(net48),
    .X(FrameStrobe_O[5]));
 sg13g2_buf_1 output49 (.A(net49),
    .X(FrameStrobe_O[6]));
 sg13g2_buf_1 output50 (.A(net50),
    .X(FrameStrobe_O[7]));
 sg13g2_buf_1 output51 (.A(net51),
    .X(FrameStrobe_O[8]));
 sg13g2_buf_1 output52 (.A(net52),
    .X(FrameStrobe_O[9]));
 sg13g2_buf_1 output53 (.A(net53),
    .X(S1BEG[0]));
 sg13g2_buf_1 output54 (.A(net54),
    .X(S1BEG[1]));
 sg13g2_buf_1 output55 (.A(net55),
    .X(S1BEG[2]));
 sg13g2_buf_1 output56 (.A(net56),
    .X(S1BEG[3]));
 sg13g2_buf_1 output57 (.A(net57),
    .X(S2BEG[0]));
 sg13g2_buf_1 output58 (.A(net58),
    .X(S2BEG[1]));
 sg13g2_buf_1 output59 (.A(net59),
    .X(S2BEG[2]));
 sg13g2_buf_1 output60 (.A(net60),
    .X(S2BEG[3]));
 sg13g2_buf_1 output61 (.A(net61),
    .X(S2BEG[4]));
 sg13g2_buf_1 output62 (.A(net62),
    .X(S2BEG[5]));
 sg13g2_buf_1 output63 (.A(net63),
    .X(S2BEG[6]));
 sg13g2_buf_1 output64 (.A(net64),
    .X(S2BEG[7]));
 sg13g2_buf_1 output65 (.A(net65),
    .X(S2BEGb[0]));
 sg13g2_buf_1 output66 (.A(net66),
    .X(S2BEGb[1]));
 sg13g2_buf_1 output67 (.A(net67),
    .X(S2BEGb[2]));
 sg13g2_buf_1 output68 (.A(net68),
    .X(S2BEGb[3]));
 sg13g2_buf_1 output69 (.A(net69),
    .X(S2BEGb[4]));
 sg13g2_buf_1 output70 (.A(net70),
    .X(S2BEGb[5]));
 sg13g2_buf_1 output71 (.A(net71),
    .X(S2BEGb[6]));
 sg13g2_buf_1 output72 (.A(net72),
    .X(S2BEGb[7]));
 sg13g2_buf_1 output73 (.A(net73),
    .X(S4BEG[0]));
 sg13g2_buf_1 output74 (.A(net74),
    .X(S4BEG[10]));
 sg13g2_buf_1 output75 (.A(net75),
    .X(S4BEG[11]));
 sg13g2_buf_1 output76 (.A(net76),
    .X(S4BEG[12]));
 sg13g2_buf_1 output77 (.A(net77),
    .X(S4BEG[13]));
 sg13g2_buf_1 output78 (.A(net78),
    .X(S4BEG[14]));
 sg13g2_buf_1 output79 (.A(net79),
    .X(S4BEG[15]));
 sg13g2_buf_1 output80 (.A(net80),
    .X(S4BEG[1]));
 sg13g2_buf_1 output81 (.A(net81),
    .X(S4BEG[2]));
 sg13g2_buf_1 output82 (.A(net82),
    .X(S4BEG[3]));
 sg13g2_buf_1 output83 (.A(net83),
    .X(S4BEG[4]));
 sg13g2_buf_1 output84 (.A(net84),
    .X(S4BEG[5]));
 sg13g2_buf_1 output85 (.A(net85),
    .X(S4BEG[6]));
 sg13g2_buf_1 output86 (.A(net86),
    .X(S4BEG[7]));
 sg13g2_buf_1 output87 (.A(net87),
    .X(S4BEG[8]));
 sg13g2_buf_1 output88 (.A(net88),
    .X(S4BEG[9]));
 sg13g2_buf_1 output89 (.A(net89),
    .X(SS4BEG[0]));
 sg13g2_buf_1 output90 (.A(net90),
    .X(SS4BEG[10]));
 sg13g2_buf_1 output91 (.A(net91),
    .X(SS4BEG[11]));
 sg13g2_buf_1 output92 (.A(net92),
    .X(SS4BEG[12]));
 sg13g2_buf_1 output93 (.A(net93),
    .X(SS4BEG[13]));
 sg13g2_buf_1 output94 (.A(net94),
    .X(SS4BEG[14]));
 sg13g2_buf_1 output95 (.A(net95),
    .X(SS4BEG[15]));
 sg13g2_buf_1 output96 (.A(net96),
    .X(SS4BEG[1]));
 sg13g2_buf_1 output97 (.A(net97),
    .X(SS4BEG[2]));
 sg13g2_buf_1 output98 (.A(net98),
    .X(SS4BEG[3]));
 sg13g2_buf_1 output99 (.A(net99),
    .X(SS4BEG[4]));
 sg13g2_buf_1 output100 (.A(net100),
    .X(SS4BEG[5]));
 sg13g2_buf_1 output101 (.A(net101),
    .X(SS4BEG[6]));
 sg13g2_buf_1 output102 (.A(net102),
    .X(SS4BEG[7]));
 sg13g2_buf_1 output103 (.A(net103),
    .X(SS4BEG[8]));
 sg13g2_buf_1 output104 (.A(net104),
    .X(SS4BEG[9]));
 sg13g2_buf_1 output105 (.A(net105),
    .X(UserCLKo));
 sg13g2_antennanp ANTENNA_1 (.A(FrameData[10]));
 sg13g2_antennanp ANTENNA_2 (.A(FrameData[5]));
 sg13g2_antennanp ANTENNA_3 (.A(FrameData[6]));
 sg13g2_antennanp ANTENNA_4 (.A(FrameData[7]));
 sg13g2_antennanp ANTENNA_5 (.A(net1));
 sg13g2_antennanp ANTENNA_6 (.A(net27));
 sg13g2_antennanp ANTENNA_7 (.A(FrameStrobe[3]));
 sg13g2_antennanp ANTENNA_8 (.A(FrameStrobe[4]));
 sg13g2_antennanp ANTENNA_9 (.A(FrameData[10]));
 sg13g2_antennanp ANTENNA_10 (.A(FrameData[5]));
 sg13g2_antennanp ANTENNA_11 (.A(FrameData[6]));
 sg13g2_antennanp ANTENNA_12 (.A(FrameData[7]));
 sg13g2_antennanp ANTENNA_13 (.A(net1));
 sg13g2_antennanp ANTENNA_14 (.A(net22));
 sg13g2_antennanp ANTENNA_15 (.A(net27));
 sg13g2_antennanp ANTENNA_16 (.A(FrameData[5]));
 sg13g2_antennanp ANTENNA_17 (.A(FrameData[6]));
 sg13g2_antennanp ANTENNA_18 (.A(FrameData[7]));
 sg13g2_antennanp ANTENNA_19 (.A(net1));
 sg13g2_antennanp ANTENNA_20 (.A(net22));
 sg13g2_antennanp ANTENNA_21 (.A(net27));
 sg13g2_antennanp ANTENNA_22 (.A(FrameData[5]));
 sg13g2_antennanp ANTENNA_23 (.A(FrameData[6]));
 sg13g2_antennanp ANTENNA_24 (.A(FrameData[7]));
 sg13g2_antennanp ANTENNA_25 (.A(net1));
 sg13g2_antennanp ANTENNA_26 (.A(net27));
 sg13g2_antennanp ANTENNA_27 (.A(FrameData[5]));
 sg13g2_antennanp ANTENNA_28 (.A(FrameData[6]));
 sg13g2_antennanp ANTENNA_29 (.A(FrameData[7]));
 sg13g2_antennanp ANTENNA_30 (.A(net1));
 sg13g2_antennanp ANTENNA_31 (.A(net27));
 sg13g2_antennanp ANTENNA_32 (.A(FrameData[5]));
 sg13g2_antennanp ANTENNA_33 (.A(FrameData[6]));
 sg13g2_antennanp ANTENNA_34 (.A(FrameData[7]));
 sg13g2_antennanp ANTENNA_35 (.A(net1));
 sg13g2_antennanp ANTENNA_36 (.A(net27));
 sg13g2_antennanp ANTENNA_37 (.A(FrameData[5]));
 sg13g2_antennanp ANTENNA_38 (.A(FrameData[6]));
 sg13g2_antennanp ANTENNA_39 (.A(FrameData[7]));
 sg13g2_antennanp ANTENNA_40 (.A(net1));
 sg13g2_antennanp ANTENNA_41 (.A(net27));
 sg13g2_antennanp ANTENNA_42 (.A(FrameData[5]));
 sg13g2_antennanp ANTENNA_43 (.A(FrameData[6]));
 sg13g2_antennanp ANTENNA_44 (.A(FrameData[7]));
 sg13g2_antennanp ANTENNA_45 (.A(net1));
 sg13g2_antennanp ANTENNA_46 (.A(net27));
 sg13g2_antennanp ANTENNA_47 (.A(FrameData[5]));
 sg13g2_antennanp ANTENNA_48 (.A(FrameData[6]));
 sg13g2_antennanp ANTENNA_49 (.A(FrameData[7]));
 sg13g2_antennanp ANTENNA_50 (.A(net1));
 sg13g2_antennanp ANTENNA_51 (.A(net27));
 sg13g2_antennanp ANTENNA_52 (.A(FrameData[5]));
 sg13g2_antennanp ANTENNA_53 (.A(FrameData[6]));
 sg13g2_antennanp ANTENNA_54 (.A(FrameData[7]));
 sg13g2_antennanp ANTENNA_55 (.A(net1));
 sg13g2_antennanp ANTENNA_56 (.A(net27));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_decap_8 FILLER_0_21 ();
 sg13g2_decap_8 FILLER_0_28 ();
 sg13g2_decap_8 FILLER_0_35 ();
 sg13g2_decap_8 FILLER_0_42 ();
 sg13g2_decap_8 FILLER_0_49 ();
 sg13g2_decap_8 FILLER_0_56 ();
 sg13g2_decap_8 FILLER_0_63 ();
 sg13g2_decap_8 FILLER_0_70 ();
 sg13g2_decap_8 FILLER_0_77 ();
 sg13g2_decap_8 FILLER_0_84 ();
 sg13g2_decap_8 FILLER_0_91 ();
 sg13g2_decap_8 FILLER_0_98 ();
 sg13g2_decap_8 FILLER_0_105 ();
 sg13g2_decap_8 FILLER_0_112 ();
 sg13g2_decap_8 FILLER_0_119 ();
 sg13g2_decap_8 FILLER_0_126 ();
 sg13g2_decap_8 FILLER_0_133 ();
 sg13g2_decap_8 FILLER_0_140 ();
 sg13g2_decap_8 FILLER_0_147 ();
 sg13g2_decap_8 FILLER_0_154 ();
 sg13g2_decap_8 FILLER_0_161 ();
 sg13g2_decap_8 FILLER_0_168 ();
 sg13g2_decap_8 FILLER_0_175 ();
 sg13g2_decap_8 FILLER_0_182 ();
 sg13g2_decap_8 FILLER_0_189 ();
 sg13g2_decap_8 FILLER_0_196 ();
 sg13g2_decap_8 FILLER_0_203 ();
 sg13g2_decap_8 FILLER_0_210 ();
 sg13g2_decap_8 FILLER_0_217 ();
 sg13g2_fill_1 FILLER_0_224 ();
 sg13g2_decap_8 FILLER_0_433 ();
 sg13g2_decap_8 FILLER_0_440 ();
 sg13g2_decap_8 FILLER_0_447 ();
 sg13g2_decap_8 FILLER_0_454 ();
 sg13g2_decap_8 FILLER_0_461 ();
 sg13g2_decap_8 FILLER_0_468 ();
 sg13g2_decap_8 FILLER_0_475 ();
 sg13g2_decap_8 FILLER_0_482 ();
 sg13g2_decap_4 FILLER_0_489 ();
 sg13g2_fill_1 FILLER_0_523 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_fill_2 FILLER_1_7 ();
 sg13g2_fill_1 FILLER_1_9 ();
 sg13g2_decap_8 FILLER_1_14 ();
 sg13g2_decap_8 FILLER_1_21 ();
 sg13g2_decap_8 FILLER_1_28 ();
 sg13g2_decap_8 FILLER_1_35 ();
 sg13g2_decap_8 FILLER_1_42 ();
 sg13g2_decap_8 FILLER_1_49 ();
 sg13g2_decap_8 FILLER_1_56 ();
 sg13g2_decap_8 FILLER_1_67 ();
 sg13g2_decap_8 FILLER_1_74 ();
 sg13g2_decap_8 FILLER_1_81 ();
 sg13g2_decap_8 FILLER_1_88 ();
 sg13g2_decap_8 FILLER_1_95 ();
 sg13g2_decap_8 FILLER_1_102 ();
 sg13g2_fill_1 FILLER_1_109 ();
 sg13g2_decap_8 FILLER_1_114 ();
 sg13g2_fill_2 FILLER_1_121 ();
 sg13g2_fill_1 FILLER_1_123 ();
 sg13g2_decap_4 FILLER_1_128 ();
 sg13g2_fill_2 FILLER_1_132 ();
 sg13g2_fill_2 FILLER_1_138 ();
 sg13g2_decap_8 FILLER_1_144 ();
 sg13g2_decap_8 FILLER_1_151 ();
 sg13g2_decap_8 FILLER_1_158 ();
 sg13g2_decap_8 FILLER_1_165 ();
 sg13g2_decap_4 FILLER_1_172 ();
 sg13g2_fill_1 FILLER_1_176 ();
 sg13g2_decap_8 FILLER_1_185 ();
 sg13g2_decap_8 FILLER_1_192 ();
 sg13g2_fill_2 FILLER_1_199 ();
 sg13g2_decap_8 FILLER_1_209 ();
 sg13g2_decap_8 FILLER_1_216 ();
 sg13g2_decap_4 FILLER_1_223 ();
 sg13g2_fill_1 FILLER_1_231 ();
 sg13g2_fill_2 FILLER_1_236 ();
 sg13g2_fill_1 FILLER_1_242 ();
 sg13g2_fill_2 FILLER_1_251 ();
 sg13g2_fill_1 FILLER_1_253 ();
 sg13g2_decap_8 FILLER_1_258 ();
 sg13g2_decap_4 FILLER_1_265 ();
 sg13g2_decap_8 FILLER_1_273 ();
 sg13g2_fill_2 FILLER_1_280 ();
 sg13g2_fill_1 FILLER_1_282 ();
 sg13g2_decap_8 FILLER_1_291 ();
 sg13g2_decap_8 FILLER_1_298 ();
 sg13g2_decap_8 FILLER_1_305 ();
 sg13g2_decap_8 FILLER_1_312 ();
 sg13g2_decap_8 FILLER_1_319 ();
 sg13g2_decap_8 FILLER_1_326 ();
 sg13g2_fill_2 FILLER_1_333 ();
 sg13g2_decap_4 FILLER_1_339 ();
 sg13g2_fill_1 FILLER_1_343 ();
 sg13g2_decap_8 FILLER_1_352 ();
 sg13g2_decap_8 FILLER_1_359 ();
 sg13g2_decap_8 FILLER_1_366 ();
 sg13g2_decap_8 FILLER_1_373 ();
 sg13g2_decap_8 FILLER_1_380 ();
 sg13g2_decap_8 FILLER_1_387 ();
 sg13g2_fill_2 FILLER_1_394 ();
 sg13g2_fill_1 FILLER_1_396 ();
 sg13g2_fill_1 FILLER_1_401 ();
 sg13g2_decap_8 FILLER_1_406 ();
 sg13g2_decap_8 FILLER_1_413 ();
 sg13g2_decap_8 FILLER_1_420 ();
 sg13g2_decap_8 FILLER_1_427 ();
 sg13g2_decap_8 FILLER_1_434 ();
 sg13g2_decap_8 FILLER_1_441 ();
 sg13g2_decap_8 FILLER_1_448 ();
 sg13g2_decap_8 FILLER_1_455 ();
 sg13g2_decap_8 FILLER_1_462 ();
 sg13g2_decap_8 FILLER_1_469 ();
 sg13g2_decap_8 FILLER_1_476 ();
 sg13g2_decap_8 FILLER_1_483 ();
 sg13g2_decap_8 FILLER_1_490 ();
 sg13g2_fill_1 FILLER_1_497 ();
 sg13g2_decap_8 FILLER_2_0 ();
 sg13g2_decap_8 FILLER_2_7 ();
 sg13g2_decap_8 FILLER_2_14 ();
 sg13g2_decap_8 FILLER_2_21 ();
 sg13g2_decap_8 FILLER_2_28 ();
 sg13g2_decap_8 FILLER_2_35 ();
 sg13g2_decap_8 FILLER_2_42 ();
 sg13g2_decap_8 FILLER_2_49 ();
 sg13g2_decap_8 FILLER_2_56 ();
 sg13g2_decap_8 FILLER_2_63 ();
 sg13g2_decap_8 FILLER_2_70 ();
 sg13g2_decap_8 FILLER_2_77 ();
 sg13g2_decap_8 FILLER_2_84 ();
 sg13g2_decap_8 FILLER_2_91 ();
 sg13g2_decap_8 FILLER_2_98 ();
 sg13g2_decap_8 FILLER_2_105 ();
 sg13g2_decap_8 FILLER_2_112 ();
 sg13g2_decap_8 FILLER_2_119 ();
 sg13g2_decap_8 FILLER_2_126 ();
 sg13g2_fill_2 FILLER_2_133 ();
 sg13g2_fill_1 FILLER_2_139 ();
 sg13g2_decap_8 FILLER_2_144 ();
 sg13g2_decap_8 FILLER_2_151 ();
 sg13g2_decap_8 FILLER_2_158 ();
 sg13g2_fill_1 FILLER_2_165 ();
 sg13g2_decap_8 FILLER_2_170 ();
 sg13g2_decap_8 FILLER_2_177 ();
 sg13g2_decap_8 FILLER_2_184 ();
 sg13g2_decap_8 FILLER_2_195 ();
 sg13g2_decap_8 FILLER_2_202 ();
 sg13g2_decap_4 FILLER_2_217 ();
 sg13g2_fill_1 FILLER_2_221 ();
 sg13g2_decap_8 FILLER_2_226 ();
 sg13g2_decap_8 FILLER_2_233 ();
 sg13g2_decap_8 FILLER_2_240 ();
 sg13g2_decap_8 FILLER_2_247 ();
 sg13g2_decap_8 FILLER_2_254 ();
 sg13g2_decap_8 FILLER_2_261 ();
 sg13g2_decap_8 FILLER_2_268 ();
 sg13g2_decap_4 FILLER_2_275 ();
 sg13g2_fill_2 FILLER_2_279 ();
 sg13g2_decap_8 FILLER_2_285 ();
 sg13g2_decap_4 FILLER_2_292 ();
 sg13g2_decap_4 FILLER_2_300 ();
 sg13g2_fill_1 FILLER_2_316 ();
 sg13g2_decap_4 FILLER_2_321 ();
 sg13g2_fill_1 FILLER_2_329 ();
 sg13g2_decap_4 FILLER_2_334 ();
 sg13g2_fill_1 FILLER_2_338 ();
 sg13g2_decap_8 FILLER_2_343 ();
 sg13g2_fill_2 FILLER_2_350 ();
 sg13g2_fill_2 FILLER_2_356 ();
 sg13g2_fill_1 FILLER_2_362 ();
 sg13g2_fill_2 FILLER_2_367 ();
 sg13g2_fill_1 FILLER_2_369 ();
 sg13g2_decap_4 FILLER_2_374 ();
 sg13g2_decap_8 FILLER_2_382 ();
 sg13g2_decap_8 FILLER_2_389 ();
 sg13g2_decap_8 FILLER_2_396 ();
 sg13g2_decap_8 FILLER_2_403 ();
 sg13g2_decap_8 FILLER_2_410 ();
 sg13g2_decap_4 FILLER_2_417 ();
 sg13g2_fill_1 FILLER_2_421 ();
 sg13g2_decap_8 FILLER_2_456 ();
 sg13g2_decap_8 FILLER_2_463 ();
 sg13g2_decap_8 FILLER_2_470 ();
 sg13g2_decap_8 FILLER_2_477 ();
 sg13g2_decap_8 FILLER_2_484 ();
 sg13g2_decap_8 FILLER_2_491 ();
 sg13g2_decap_8 FILLER_2_498 ();
 sg13g2_fill_2 FILLER_2_505 ();
 sg13g2_fill_1 FILLER_2_519 ();
 sg13g2_decap_8 FILLER_3_0 ();
 sg13g2_decap_8 FILLER_3_7 ();
 sg13g2_decap_8 FILLER_3_14 ();
 sg13g2_decap_8 FILLER_3_21 ();
 sg13g2_decap_8 FILLER_3_28 ();
 sg13g2_decap_8 FILLER_3_35 ();
 sg13g2_decap_8 FILLER_3_42 ();
 sg13g2_decap_8 FILLER_3_49 ();
 sg13g2_decap_8 FILLER_3_56 ();
 sg13g2_decap_8 FILLER_3_63 ();
 sg13g2_decap_8 FILLER_3_70 ();
 sg13g2_decap_8 FILLER_3_77 ();
 sg13g2_decap_8 FILLER_3_84 ();
 sg13g2_decap_8 FILLER_3_91 ();
 sg13g2_decap_8 FILLER_3_98 ();
 sg13g2_decap_8 FILLER_3_105 ();
 sg13g2_decap_8 FILLER_3_112 ();
 sg13g2_decap_8 FILLER_3_119 ();
 sg13g2_fill_1 FILLER_3_126 ();
 sg13g2_decap_8 FILLER_3_131 ();
 sg13g2_decap_8 FILLER_3_138 ();
 sg13g2_decap_8 FILLER_3_145 ();
 sg13g2_decap_4 FILLER_3_152 ();
 sg13g2_fill_2 FILLER_3_156 ();
 sg13g2_fill_1 FILLER_3_162 ();
 sg13g2_decap_8 FILLER_3_167 ();
 sg13g2_decap_8 FILLER_3_174 ();
 sg13g2_decap_4 FILLER_3_181 ();
 sg13g2_fill_2 FILLER_3_185 ();
 sg13g2_decap_8 FILLER_3_191 ();
 sg13g2_decap_8 FILLER_3_198 ();
 sg13g2_decap_8 FILLER_3_205 ();
 sg13g2_decap_8 FILLER_3_212 ();
 sg13g2_decap_8 FILLER_3_219 ();
 sg13g2_fill_1 FILLER_3_226 ();
 sg13g2_decap_8 FILLER_3_231 ();
 sg13g2_decap_8 FILLER_3_238 ();
 sg13g2_decap_8 FILLER_3_245 ();
 sg13g2_decap_8 FILLER_3_252 ();
 sg13g2_decap_8 FILLER_3_259 ();
 sg13g2_decap_8 FILLER_3_266 ();
 sg13g2_decap_4 FILLER_3_273 ();
 sg13g2_fill_2 FILLER_3_277 ();
 sg13g2_decap_8 FILLER_3_283 ();
 sg13g2_decap_8 FILLER_3_290 ();
 sg13g2_decap_8 FILLER_3_297 ();
 sg13g2_decap_8 FILLER_3_304 ();
 sg13g2_decap_8 FILLER_3_311 ();
 sg13g2_decap_8 FILLER_3_318 ();
 sg13g2_decap_8 FILLER_3_325 ();
 sg13g2_decap_8 FILLER_3_332 ();
 sg13g2_decap_8 FILLER_3_339 ();
 sg13g2_decap_8 FILLER_3_346 ();
 sg13g2_decap_8 FILLER_3_353 ();
 sg13g2_decap_8 FILLER_3_360 ();
 sg13g2_decap_8 FILLER_3_367 ();
 sg13g2_decap_8 FILLER_3_374 ();
 sg13g2_decap_8 FILLER_3_381 ();
 sg13g2_fill_2 FILLER_3_388 ();
 sg13g2_decap_8 FILLER_3_394 ();
 sg13g2_decap_8 FILLER_3_401 ();
 sg13g2_decap_8 FILLER_3_408 ();
 sg13g2_decap_8 FILLER_3_415 ();
 sg13g2_decap_8 FILLER_3_422 ();
 sg13g2_decap_8 FILLER_3_429 ();
 sg13g2_decap_8 FILLER_3_436 ();
 sg13g2_decap_8 FILLER_3_443 ();
 sg13g2_decap_8 FILLER_3_450 ();
 sg13g2_decap_8 FILLER_3_457 ();
 sg13g2_decap_8 FILLER_3_464 ();
 sg13g2_decap_8 FILLER_3_471 ();
 sg13g2_decap_8 FILLER_3_478 ();
 sg13g2_decap_8 FILLER_3_485 ();
 sg13g2_decap_8 FILLER_3_492 ();
 sg13g2_decap_8 FILLER_3_499 ();
 sg13g2_decap_8 FILLER_3_506 ();
 sg13g2_fill_2 FILLER_3_513 ();
 sg13g2_fill_1 FILLER_3_515 ();
 sg13g2_decap_8 FILLER_4_0 ();
 sg13g2_decap_8 FILLER_4_7 ();
 sg13g2_decap_8 FILLER_4_14 ();
 sg13g2_decap_8 FILLER_4_21 ();
 sg13g2_decap_8 FILLER_4_28 ();
 sg13g2_decap_8 FILLER_4_35 ();
 sg13g2_decap_8 FILLER_4_42 ();
 sg13g2_decap_8 FILLER_4_49 ();
 sg13g2_decap_8 FILLER_4_56 ();
 sg13g2_decap_8 FILLER_4_63 ();
 sg13g2_decap_8 FILLER_4_70 ();
 sg13g2_decap_8 FILLER_4_77 ();
 sg13g2_decap_8 FILLER_4_84 ();
 sg13g2_decap_8 FILLER_4_91 ();
 sg13g2_decap_8 FILLER_4_98 ();
 sg13g2_decap_8 FILLER_4_105 ();
 sg13g2_decap_8 FILLER_4_112 ();
 sg13g2_decap_8 FILLER_4_119 ();
 sg13g2_decap_8 FILLER_4_126 ();
 sg13g2_decap_8 FILLER_4_133 ();
 sg13g2_fill_2 FILLER_4_144 ();
 sg13g2_decap_8 FILLER_4_150 ();
 sg13g2_decap_8 FILLER_4_157 ();
 sg13g2_decap_8 FILLER_4_164 ();
 sg13g2_decap_8 FILLER_4_171 ();
 sg13g2_decap_8 FILLER_4_178 ();
 sg13g2_decap_8 FILLER_4_185 ();
 sg13g2_decap_8 FILLER_4_192 ();
 sg13g2_decap_8 FILLER_4_199 ();
 sg13g2_decap_8 FILLER_4_206 ();
 sg13g2_decap_8 FILLER_4_213 ();
 sg13g2_decap_8 FILLER_4_220 ();
 sg13g2_decap_8 FILLER_4_227 ();
 sg13g2_decap_4 FILLER_4_234 ();
 sg13g2_fill_1 FILLER_4_238 ();
 sg13g2_fill_2 FILLER_4_243 ();
 sg13g2_fill_1 FILLER_4_245 ();
 sg13g2_decap_8 FILLER_4_254 ();
 sg13g2_decap_8 FILLER_4_261 ();
 sg13g2_decap_8 FILLER_4_268 ();
 sg13g2_decap_8 FILLER_4_275 ();
 sg13g2_decap_8 FILLER_4_282 ();
 sg13g2_decap_8 FILLER_4_289 ();
 sg13g2_decap_4 FILLER_4_296 ();
 sg13g2_decap_8 FILLER_4_304 ();
 sg13g2_decap_8 FILLER_4_311 ();
 sg13g2_decap_8 FILLER_4_318 ();
 sg13g2_decap_8 FILLER_4_325 ();
 sg13g2_decap_8 FILLER_4_332 ();
 sg13g2_decap_8 FILLER_4_339 ();
 sg13g2_decap_8 FILLER_4_346 ();
 sg13g2_decap_8 FILLER_4_353 ();
 sg13g2_decap_8 FILLER_4_360 ();
 sg13g2_decap_8 FILLER_4_367 ();
 sg13g2_decap_8 FILLER_4_374 ();
 sg13g2_decap_8 FILLER_4_381 ();
 sg13g2_decap_8 FILLER_4_388 ();
 sg13g2_decap_8 FILLER_4_395 ();
 sg13g2_decap_8 FILLER_4_402 ();
 sg13g2_decap_8 FILLER_4_409 ();
 sg13g2_decap_8 FILLER_4_416 ();
 sg13g2_decap_8 FILLER_4_423 ();
 sg13g2_decap_8 FILLER_4_430 ();
 sg13g2_decap_8 FILLER_4_437 ();
 sg13g2_decap_8 FILLER_4_444 ();
 sg13g2_decap_8 FILLER_4_451 ();
 sg13g2_decap_8 FILLER_4_458 ();
 sg13g2_decap_8 FILLER_4_465 ();
 sg13g2_decap_8 FILLER_4_472 ();
 sg13g2_decap_8 FILLER_4_479 ();
 sg13g2_decap_8 FILLER_4_486 ();
 sg13g2_decap_8 FILLER_4_493 ();
 sg13g2_decap_8 FILLER_4_500 ();
 sg13g2_decap_8 FILLER_4_507 ();
 sg13g2_decap_8 FILLER_4_514 ();
 sg13g2_fill_2 FILLER_4_521 ();
 sg13g2_decap_8 FILLER_5_0 ();
 sg13g2_decap_8 FILLER_5_7 ();
 sg13g2_decap_8 FILLER_5_14 ();
 sg13g2_decap_8 FILLER_5_21 ();
 sg13g2_decap_8 FILLER_5_28 ();
 sg13g2_decap_8 FILLER_5_35 ();
 sg13g2_decap_8 FILLER_5_42 ();
 sg13g2_decap_8 FILLER_5_49 ();
 sg13g2_decap_8 FILLER_5_56 ();
 sg13g2_decap_8 FILLER_5_63 ();
 sg13g2_decap_8 FILLER_5_70 ();
 sg13g2_decap_8 FILLER_5_77 ();
 sg13g2_decap_8 FILLER_5_84 ();
 sg13g2_decap_8 FILLER_5_91 ();
 sg13g2_decap_8 FILLER_5_98 ();
 sg13g2_decap_8 FILLER_5_105 ();
 sg13g2_decap_8 FILLER_5_112 ();
 sg13g2_decap_8 FILLER_5_119 ();
 sg13g2_decap_8 FILLER_5_126 ();
 sg13g2_decap_8 FILLER_5_133 ();
 sg13g2_decap_8 FILLER_5_140 ();
 sg13g2_decap_8 FILLER_5_147 ();
 sg13g2_decap_8 FILLER_5_154 ();
 sg13g2_decap_8 FILLER_5_161 ();
 sg13g2_decap_8 FILLER_5_168 ();
 sg13g2_decap_8 FILLER_5_175 ();
 sg13g2_decap_8 FILLER_5_182 ();
 sg13g2_decap_8 FILLER_5_189 ();
 sg13g2_decap_8 FILLER_5_196 ();
 sg13g2_decap_8 FILLER_5_203 ();
 sg13g2_decap_8 FILLER_5_210 ();
 sg13g2_decap_8 FILLER_5_217 ();
 sg13g2_decap_8 FILLER_5_224 ();
 sg13g2_decap_4 FILLER_5_231 ();
 sg13g2_fill_1 FILLER_5_235 ();
 sg13g2_decap_8 FILLER_5_240 ();
 sg13g2_decap_8 FILLER_5_247 ();
 sg13g2_decap_8 FILLER_5_254 ();
 sg13g2_decap_8 FILLER_5_261 ();
 sg13g2_decap_8 FILLER_5_268 ();
 sg13g2_fill_2 FILLER_5_275 ();
 sg13g2_decap_8 FILLER_5_281 ();
 sg13g2_decap_8 FILLER_5_288 ();
 sg13g2_decap_8 FILLER_5_295 ();
 sg13g2_decap_8 FILLER_5_302 ();
 sg13g2_decap_8 FILLER_5_309 ();
 sg13g2_decap_8 FILLER_5_316 ();
 sg13g2_decap_8 FILLER_5_323 ();
 sg13g2_decap_8 FILLER_5_330 ();
 sg13g2_decap_8 FILLER_5_337 ();
 sg13g2_decap_8 FILLER_5_344 ();
 sg13g2_decap_8 FILLER_5_351 ();
 sg13g2_fill_2 FILLER_5_358 ();
 sg13g2_decap_8 FILLER_5_366 ();
 sg13g2_decap_8 FILLER_5_373 ();
 sg13g2_decap_8 FILLER_5_380 ();
 sg13g2_decap_8 FILLER_5_387 ();
 sg13g2_decap_8 FILLER_5_394 ();
 sg13g2_decap_8 FILLER_5_401 ();
 sg13g2_decap_8 FILLER_5_408 ();
 sg13g2_decap_8 FILLER_5_415 ();
 sg13g2_decap_8 FILLER_5_422 ();
 sg13g2_decap_8 FILLER_5_429 ();
 sg13g2_decap_8 FILLER_5_436 ();
 sg13g2_decap_8 FILLER_5_443 ();
 sg13g2_decap_8 FILLER_5_450 ();
 sg13g2_decap_8 FILLER_5_457 ();
 sg13g2_decap_8 FILLER_5_464 ();
 sg13g2_decap_8 FILLER_5_471 ();
 sg13g2_decap_8 FILLER_5_478 ();
 sg13g2_decap_8 FILLER_5_485 ();
 sg13g2_decap_8 FILLER_5_492 ();
 sg13g2_decap_8 FILLER_5_499 ();
 sg13g2_decap_8 FILLER_5_506 ();
 sg13g2_decap_8 FILLER_5_513 ();
 sg13g2_fill_2 FILLER_5_520 ();
 sg13g2_fill_1 FILLER_5_522 ();
 sg13g2_decap_8 FILLER_6_0 ();
 sg13g2_decap_8 FILLER_6_7 ();
 sg13g2_decap_8 FILLER_6_14 ();
 sg13g2_decap_8 FILLER_6_21 ();
 sg13g2_decap_8 FILLER_6_28 ();
 sg13g2_decap_8 FILLER_6_35 ();
 sg13g2_decap_8 FILLER_6_42 ();
 sg13g2_decap_8 FILLER_6_49 ();
 sg13g2_decap_8 FILLER_6_56 ();
 sg13g2_decap_8 FILLER_6_63 ();
 sg13g2_decap_8 FILLER_6_70 ();
 sg13g2_decap_8 FILLER_6_77 ();
 sg13g2_decap_8 FILLER_6_84 ();
 sg13g2_decap_8 FILLER_6_91 ();
 sg13g2_decap_8 FILLER_6_98 ();
 sg13g2_decap_8 FILLER_6_105 ();
 sg13g2_decap_8 FILLER_6_112 ();
 sg13g2_decap_8 FILLER_6_119 ();
 sg13g2_decap_8 FILLER_6_126 ();
 sg13g2_decap_8 FILLER_6_133 ();
 sg13g2_decap_8 FILLER_6_140 ();
 sg13g2_decap_8 FILLER_6_147 ();
 sg13g2_decap_8 FILLER_6_154 ();
 sg13g2_decap_8 FILLER_6_161 ();
 sg13g2_decap_8 FILLER_6_168 ();
 sg13g2_decap_8 FILLER_6_175 ();
 sg13g2_decap_8 FILLER_6_182 ();
 sg13g2_decap_8 FILLER_6_189 ();
 sg13g2_decap_8 FILLER_6_196 ();
 sg13g2_decap_8 FILLER_6_203 ();
 sg13g2_decap_8 FILLER_6_210 ();
 sg13g2_decap_8 FILLER_6_217 ();
 sg13g2_decap_8 FILLER_6_228 ();
 sg13g2_decap_8 FILLER_6_235 ();
 sg13g2_decap_8 FILLER_6_242 ();
 sg13g2_fill_2 FILLER_6_249 ();
 sg13g2_fill_1 FILLER_6_251 ();
 sg13g2_decap_8 FILLER_6_260 ();
 sg13g2_decap_8 FILLER_6_267 ();
 sg13g2_decap_8 FILLER_6_274 ();
 sg13g2_decap_8 FILLER_6_281 ();
 sg13g2_decap_8 FILLER_6_288 ();
 sg13g2_decap_8 FILLER_6_295 ();
 sg13g2_decap_8 FILLER_6_302 ();
 sg13g2_decap_8 FILLER_6_309 ();
 sg13g2_decap_8 FILLER_6_316 ();
 sg13g2_decap_8 FILLER_6_323 ();
 sg13g2_decap_8 FILLER_6_330 ();
 sg13g2_decap_8 FILLER_6_337 ();
 sg13g2_decap_8 FILLER_6_344 ();
 sg13g2_decap_4 FILLER_6_351 ();
 sg13g2_fill_2 FILLER_6_355 ();
 sg13g2_fill_1 FILLER_6_385 ();
 sg13g2_decap_8 FILLER_6_390 ();
 sg13g2_decap_8 FILLER_6_397 ();
 sg13g2_decap_8 FILLER_6_404 ();
 sg13g2_decap_8 FILLER_6_411 ();
 sg13g2_decap_8 FILLER_6_418 ();
 sg13g2_decap_8 FILLER_6_425 ();
 sg13g2_decap_8 FILLER_6_432 ();
 sg13g2_decap_8 FILLER_6_439 ();
 sg13g2_decap_8 FILLER_6_446 ();
 sg13g2_decap_8 FILLER_6_453 ();
 sg13g2_decap_8 FILLER_6_460 ();
 sg13g2_decap_8 FILLER_6_467 ();
 sg13g2_decap_8 FILLER_6_474 ();
 sg13g2_decap_8 FILLER_6_481 ();
 sg13g2_decap_8 FILLER_6_488 ();
 sg13g2_decap_8 FILLER_6_495 ();
 sg13g2_decap_8 FILLER_6_502 ();
 sg13g2_decap_8 FILLER_6_509 ();
 sg13g2_decap_8 FILLER_6_516 ();
 sg13g2_decap_8 FILLER_7_0 ();
 sg13g2_decap_8 FILLER_7_7 ();
 sg13g2_decap_8 FILLER_7_14 ();
 sg13g2_decap_8 FILLER_7_21 ();
 sg13g2_decap_8 FILLER_7_28 ();
 sg13g2_decap_8 FILLER_7_35 ();
 sg13g2_decap_8 FILLER_7_42 ();
 sg13g2_decap_8 FILLER_7_49 ();
 sg13g2_decap_8 FILLER_7_56 ();
 sg13g2_decap_8 FILLER_7_63 ();
 sg13g2_decap_8 FILLER_7_70 ();
 sg13g2_decap_8 FILLER_7_77 ();
 sg13g2_decap_8 FILLER_7_84 ();
 sg13g2_decap_8 FILLER_7_91 ();
 sg13g2_decap_8 FILLER_7_98 ();
 sg13g2_decap_8 FILLER_7_105 ();
 sg13g2_decap_8 FILLER_7_112 ();
 sg13g2_decap_8 FILLER_7_119 ();
 sg13g2_decap_8 FILLER_7_126 ();
 sg13g2_decap_8 FILLER_7_133 ();
 sg13g2_decap_8 FILLER_7_140 ();
 sg13g2_decap_8 FILLER_7_147 ();
 sg13g2_decap_8 FILLER_7_154 ();
 sg13g2_decap_8 FILLER_7_161 ();
 sg13g2_decap_8 FILLER_7_168 ();
 sg13g2_decap_8 FILLER_7_175 ();
 sg13g2_fill_2 FILLER_7_182 ();
 sg13g2_decap_8 FILLER_7_188 ();
 sg13g2_decap_8 FILLER_7_195 ();
 sg13g2_decap_8 FILLER_7_202 ();
 sg13g2_decap_8 FILLER_7_209 ();
 sg13g2_decap_8 FILLER_7_216 ();
 sg13g2_decap_8 FILLER_7_223 ();
 sg13g2_fill_2 FILLER_7_230 ();
 sg13g2_fill_1 FILLER_7_232 ();
 sg13g2_decap_8 FILLER_7_237 ();
 sg13g2_decap_8 FILLER_7_244 ();
 sg13g2_decap_8 FILLER_7_251 ();
 sg13g2_decap_8 FILLER_7_258 ();
 sg13g2_decap_8 FILLER_7_265 ();
 sg13g2_decap_8 FILLER_7_272 ();
 sg13g2_decap_8 FILLER_7_279 ();
 sg13g2_decap_8 FILLER_7_286 ();
 sg13g2_decap_4 FILLER_7_293 ();
 sg13g2_fill_1 FILLER_7_301 ();
 sg13g2_decap_8 FILLER_7_306 ();
 sg13g2_decap_8 FILLER_7_313 ();
 sg13g2_decap_8 FILLER_7_320 ();
 sg13g2_decap_8 FILLER_7_327 ();
 sg13g2_decap_8 FILLER_7_334 ();
 sg13g2_decap_8 FILLER_7_341 ();
 sg13g2_decap_4 FILLER_7_348 ();
 sg13g2_fill_2 FILLER_7_352 ();
 sg13g2_decap_8 FILLER_7_360 ();
 sg13g2_decap_8 FILLER_7_367 ();
 sg13g2_decap_8 FILLER_7_374 ();
 sg13g2_decap_8 FILLER_7_381 ();
 sg13g2_decap_8 FILLER_7_388 ();
 sg13g2_decap_8 FILLER_7_395 ();
 sg13g2_decap_8 FILLER_7_402 ();
 sg13g2_decap_8 FILLER_7_409 ();
 sg13g2_decap_8 FILLER_7_416 ();
 sg13g2_decap_8 FILLER_7_423 ();
 sg13g2_decap_8 FILLER_7_430 ();
 sg13g2_decap_8 FILLER_7_437 ();
 sg13g2_decap_8 FILLER_7_444 ();
 sg13g2_decap_8 FILLER_7_451 ();
 sg13g2_decap_8 FILLER_7_458 ();
 sg13g2_decap_8 FILLER_7_465 ();
 sg13g2_decap_8 FILLER_7_472 ();
 sg13g2_decap_8 FILLER_7_479 ();
 sg13g2_decap_8 FILLER_7_486 ();
 sg13g2_decap_8 FILLER_7_493 ();
 sg13g2_decap_8 FILLER_7_500 ();
 sg13g2_decap_8 FILLER_7_507 ();
 sg13g2_decap_8 FILLER_7_514 ();
 sg13g2_fill_2 FILLER_7_521 ();
 sg13g2_decap_8 FILLER_8_0 ();
 sg13g2_decap_8 FILLER_8_7 ();
 sg13g2_decap_8 FILLER_8_14 ();
 sg13g2_decap_8 FILLER_8_21 ();
 sg13g2_decap_8 FILLER_8_28 ();
 sg13g2_decap_8 FILLER_8_35 ();
 sg13g2_decap_8 FILLER_8_42 ();
 sg13g2_decap_8 FILLER_8_49 ();
 sg13g2_decap_8 FILLER_8_56 ();
 sg13g2_decap_8 FILLER_8_63 ();
 sg13g2_decap_8 FILLER_8_70 ();
 sg13g2_decap_8 FILLER_8_77 ();
 sg13g2_decap_8 FILLER_8_84 ();
 sg13g2_decap_8 FILLER_8_91 ();
 sg13g2_decap_8 FILLER_8_98 ();
 sg13g2_decap_8 FILLER_8_105 ();
 sg13g2_decap_8 FILLER_8_112 ();
 sg13g2_decap_8 FILLER_8_119 ();
 sg13g2_decap_8 FILLER_8_126 ();
 sg13g2_decap_8 FILLER_8_133 ();
 sg13g2_decap_8 FILLER_8_140 ();
 sg13g2_decap_8 FILLER_8_147 ();
 sg13g2_decap_8 FILLER_8_154 ();
 sg13g2_decap_8 FILLER_8_161 ();
 sg13g2_decap_8 FILLER_8_168 ();
 sg13g2_decap_8 FILLER_8_175 ();
 sg13g2_decap_8 FILLER_8_182 ();
 sg13g2_decap_8 FILLER_8_189 ();
 sg13g2_decap_8 FILLER_8_196 ();
 sg13g2_decap_8 FILLER_8_203 ();
 sg13g2_decap_8 FILLER_8_210 ();
 sg13g2_decap_8 FILLER_8_217 ();
 sg13g2_decap_4 FILLER_8_224 ();
 sg13g2_fill_2 FILLER_8_228 ();
 sg13g2_decap_8 FILLER_8_234 ();
 sg13g2_decap_8 FILLER_8_241 ();
 sg13g2_decap_8 FILLER_8_248 ();
 sg13g2_decap_8 FILLER_8_255 ();
 sg13g2_decap_8 FILLER_8_262 ();
 sg13g2_decap_8 FILLER_8_269 ();
 sg13g2_fill_2 FILLER_8_276 ();
 sg13g2_fill_1 FILLER_8_278 ();
 sg13g2_decap_8 FILLER_8_283 ();
 sg13g2_decap_8 FILLER_8_290 ();
 sg13g2_decap_8 FILLER_8_297 ();
 sg13g2_decap_8 FILLER_8_304 ();
 sg13g2_decap_4 FILLER_8_311 ();
 sg13g2_decap_8 FILLER_8_319 ();
 sg13g2_decap_8 FILLER_8_326 ();
 sg13g2_fill_2 FILLER_8_333 ();
 sg13g2_fill_1 FILLER_8_335 ();
 sg13g2_decap_8 FILLER_8_339 ();
 sg13g2_decap_8 FILLER_8_346 ();
 sg13g2_fill_1 FILLER_8_353 ();
 sg13g2_decap_8 FILLER_8_358 ();
 sg13g2_decap_8 FILLER_8_365 ();
 sg13g2_decap_8 FILLER_8_372 ();
 sg13g2_decap_8 FILLER_8_379 ();
 sg13g2_decap_8 FILLER_8_386 ();
 sg13g2_decap_8 FILLER_8_393 ();
 sg13g2_decap_8 FILLER_8_400 ();
 sg13g2_decap_8 FILLER_8_407 ();
 sg13g2_decap_8 FILLER_8_414 ();
 sg13g2_decap_8 FILLER_8_421 ();
 sg13g2_decap_8 FILLER_8_428 ();
 sg13g2_decap_8 FILLER_8_435 ();
 sg13g2_decap_8 FILLER_8_442 ();
 sg13g2_decap_8 FILLER_8_449 ();
 sg13g2_decap_8 FILLER_8_456 ();
 sg13g2_decap_8 FILLER_8_463 ();
 sg13g2_decap_8 FILLER_8_470 ();
 sg13g2_decap_8 FILLER_8_477 ();
 sg13g2_decap_8 FILLER_8_484 ();
 sg13g2_decap_8 FILLER_8_491 ();
 sg13g2_decap_8 FILLER_8_498 ();
 sg13g2_decap_8 FILLER_8_505 ();
 sg13g2_decap_8 FILLER_8_512 ();
 sg13g2_decap_4 FILLER_8_519 ();
 sg13g2_decap_8 FILLER_9_0 ();
 sg13g2_decap_8 FILLER_9_7 ();
 sg13g2_decap_8 FILLER_9_14 ();
 sg13g2_decap_8 FILLER_9_21 ();
 sg13g2_decap_8 FILLER_9_28 ();
 sg13g2_decap_8 FILLER_9_35 ();
 sg13g2_decap_8 FILLER_9_42 ();
 sg13g2_decap_8 FILLER_9_49 ();
 sg13g2_decap_8 FILLER_9_56 ();
 sg13g2_decap_8 FILLER_9_63 ();
 sg13g2_decap_8 FILLER_9_70 ();
 sg13g2_decap_8 FILLER_9_77 ();
 sg13g2_decap_8 FILLER_9_84 ();
 sg13g2_decap_8 FILLER_9_91 ();
 sg13g2_decap_8 FILLER_9_98 ();
 sg13g2_decap_8 FILLER_9_105 ();
 sg13g2_decap_8 FILLER_9_112 ();
 sg13g2_decap_8 FILLER_9_119 ();
 sg13g2_decap_8 FILLER_9_126 ();
 sg13g2_decap_8 FILLER_9_133 ();
 sg13g2_decap_8 FILLER_9_140 ();
 sg13g2_decap_8 FILLER_9_147 ();
 sg13g2_decap_8 FILLER_9_154 ();
 sg13g2_decap_8 FILLER_9_161 ();
 sg13g2_decap_8 FILLER_9_168 ();
 sg13g2_decap_8 FILLER_9_175 ();
 sg13g2_decap_8 FILLER_9_182 ();
 sg13g2_decap_8 FILLER_9_189 ();
 sg13g2_decap_8 FILLER_9_196 ();
 sg13g2_decap_8 FILLER_9_203 ();
 sg13g2_decap_8 FILLER_9_210 ();
 sg13g2_decap_8 FILLER_9_217 ();
 sg13g2_decap_8 FILLER_9_224 ();
 sg13g2_decap_8 FILLER_9_231 ();
 sg13g2_decap_8 FILLER_9_238 ();
 sg13g2_decap_8 FILLER_9_245 ();
 sg13g2_fill_2 FILLER_9_252 ();
 sg13g2_decap_8 FILLER_9_258 ();
 sg13g2_decap_8 FILLER_9_265 ();
 sg13g2_decap_4 FILLER_9_272 ();
 sg13g2_decap_8 FILLER_9_284 ();
 sg13g2_decap_8 FILLER_9_291 ();
 sg13g2_decap_8 FILLER_9_298 ();
 sg13g2_decap_8 FILLER_9_305 ();
 sg13g2_decap_8 FILLER_9_312 ();
 sg13g2_decap_8 FILLER_9_319 ();
 sg13g2_decap_8 FILLER_9_326 ();
 sg13g2_decap_8 FILLER_9_364 ();
 sg13g2_decap_8 FILLER_9_371 ();
 sg13g2_decap_8 FILLER_9_378 ();
 sg13g2_decap_8 FILLER_9_385 ();
 sg13g2_decap_8 FILLER_9_392 ();
 sg13g2_decap_8 FILLER_9_399 ();
 sg13g2_decap_8 FILLER_9_406 ();
 sg13g2_decap_8 FILLER_9_413 ();
 sg13g2_decap_8 FILLER_9_420 ();
 sg13g2_decap_8 FILLER_9_427 ();
 sg13g2_decap_8 FILLER_9_434 ();
 sg13g2_decap_8 FILLER_9_441 ();
 sg13g2_decap_8 FILLER_9_448 ();
 sg13g2_decap_8 FILLER_9_455 ();
 sg13g2_decap_8 FILLER_9_462 ();
 sg13g2_decap_8 FILLER_9_469 ();
 sg13g2_decap_8 FILLER_9_476 ();
 sg13g2_decap_8 FILLER_9_483 ();
 sg13g2_decap_8 FILLER_9_490 ();
 sg13g2_decap_8 FILLER_9_497 ();
 sg13g2_decap_8 FILLER_9_504 ();
 sg13g2_decap_8 FILLER_9_511 ();
 sg13g2_decap_4 FILLER_9_518 ();
 sg13g2_fill_1 FILLER_9_522 ();
 sg13g2_decap_8 FILLER_10_0 ();
 sg13g2_decap_8 FILLER_10_7 ();
 sg13g2_decap_8 FILLER_10_14 ();
 sg13g2_decap_8 FILLER_10_21 ();
 sg13g2_decap_8 FILLER_10_28 ();
 sg13g2_decap_8 FILLER_10_35 ();
 sg13g2_decap_8 FILLER_10_42 ();
 sg13g2_decap_8 FILLER_10_49 ();
 sg13g2_decap_8 FILLER_10_56 ();
 sg13g2_decap_8 FILLER_10_63 ();
 sg13g2_decap_8 FILLER_10_70 ();
 sg13g2_decap_8 FILLER_10_77 ();
 sg13g2_decap_8 FILLER_10_84 ();
 sg13g2_decap_8 FILLER_10_91 ();
 sg13g2_decap_8 FILLER_10_98 ();
 sg13g2_decap_8 FILLER_10_105 ();
 sg13g2_decap_8 FILLER_10_112 ();
 sg13g2_decap_8 FILLER_10_119 ();
 sg13g2_fill_2 FILLER_10_126 ();
 sg13g2_fill_1 FILLER_10_128 ();
 sg13g2_decap_8 FILLER_10_140 ();
 sg13g2_fill_2 FILLER_10_147 ();
 sg13g2_decap_8 FILLER_10_156 ();
 sg13g2_decap_8 FILLER_10_163 ();
 sg13g2_decap_8 FILLER_10_170 ();
 sg13g2_fill_2 FILLER_10_177 ();
 sg13g2_fill_1 FILLER_10_179 ();
 sg13g2_decap_8 FILLER_10_184 ();
 sg13g2_decap_8 FILLER_10_191 ();
 sg13g2_decap_8 FILLER_10_198 ();
 sg13g2_decap_8 FILLER_10_209 ();
 sg13g2_decap_8 FILLER_10_216 ();
 sg13g2_decap_4 FILLER_10_223 ();
 sg13g2_fill_2 FILLER_10_227 ();
 sg13g2_fill_2 FILLER_10_233 ();
 sg13g2_decap_8 FILLER_10_239 ();
 sg13g2_decap_4 FILLER_10_246 ();
 sg13g2_fill_2 FILLER_10_250 ();
 sg13g2_decap_4 FILLER_10_256 ();
 sg13g2_fill_1 FILLER_10_264 ();
 sg13g2_decap_8 FILLER_10_269 ();
 sg13g2_fill_2 FILLER_10_276 ();
 sg13g2_decap_4 FILLER_10_282 ();
 sg13g2_fill_2 FILLER_10_286 ();
 sg13g2_decap_4 FILLER_10_292 ();
 sg13g2_fill_1 FILLER_10_296 ();
 sg13g2_fill_1 FILLER_10_301 ();
 sg13g2_decap_8 FILLER_10_306 ();
 sg13g2_decap_8 FILLER_10_313 ();
 sg13g2_decap_8 FILLER_10_320 ();
 sg13g2_decap_8 FILLER_10_327 ();
 sg13g2_decap_8 FILLER_10_334 ();
 sg13g2_decap_8 FILLER_10_341 ();
 sg13g2_decap_8 FILLER_10_348 ();
 sg13g2_decap_8 FILLER_10_355 ();
 sg13g2_decap_8 FILLER_10_362 ();
 sg13g2_decap_8 FILLER_10_369 ();
 sg13g2_decap_8 FILLER_10_376 ();
 sg13g2_decap_8 FILLER_10_383 ();
 sg13g2_decap_8 FILLER_10_390 ();
 sg13g2_decap_8 FILLER_10_397 ();
 sg13g2_fill_1 FILLER_10_404 ();
 sg13g2_fill_2 FILLER_10_409 ();
 sg13g2_decap_4 FILLER_10_415 ();
 sg13g2_fill_2 FILLER_10_419 ();
 sg13g2_decap_4 FILLER_10_425 ();
 sg13g2_fill_2 FILLER_10_429 ();
 sg13g2_decap_4 FILLER_10_435 ();
 sg13g2_fill_1 FILLER_10_439 ();
 sg13g2_fill_2 FILLER_10_444 ();
 sg13g2_decap_4 FILLER_10_450 ();
 sg13g2_fill_2 FILLER_10_454 ();
 sg13g2_decap_8 FILLER_10_460 ();
 sg13g2_fill_2 FILLER_10_467 ();
 sg13g2_fill_1 FILLER_10_473 ();
 sg13g2_decap_8 FILLER_10_482 ();
 sg13g2_fill_1 FILLER_10_489 ();
 sg13g2_decap_8 FILLER_10_498 ();
 sg13g2_decap_4 FILLER_10_505 ();
 sg13g2_fill_2 FILLER_10_509 ();
 sg13g2_fill_1 FILLER_10_522 ();
 sg13g2_decap_4 FILLER_11_0 ();
 sg13g2_fill_1 FILLER_11_4 ();
 sg13g2_decap_8 FILLER_11_9 ();
 sg13g2_decap_8 FILLER_11_16 ();
 sg13g2_decap_8 FILLER_11_23 ();
 sg13g2_fill_1 FILLER_11_30 ();
 sg13g2_decap_8 FILLER_11_35 ();
 sg13g2_decap_8 FILLER_11_42 ();
 sg13g2_decap_8 FILLER_11_49 ();
 sg13g2_fill_1 FILLER_11_56 ();
 sg13g2_decap_8 FILLER_11_61 ();
 sg13g2_decap_8 FILLER_11_68 ();
 sg13g2_decap_8 FILLER_11_75 ();
 sg13g2_fill_1 FILLER_11_82 ();
 sg13g2_decap_8 FILLER_11_87 ();
 sg13g2_decap_8 FILLER_11_94 ();
 sg13g2_decap_8 FILLER_11_101 ();
 sg13g2_fill_1 FILLER_11_108 ();
 sg13g2_decap_8 FILLER_11_113 ();
 sg13g2_decap_8 FILLER_11_120 ();
 sg13g2_decap_8 FILLER_11_127 ();
 sg13g2_fill_1 FILLER_11_134 ();
 sg13g2_decap_8 FILLER_11_139 ();
 sg13g2_decap_8 FILLER_11_146 ();
 sg13g2_decap_8 FILLER_11_153 ();
 sg13g2_fill_1 FILLER_11_160 ();
 sg13g2_decap_8 FILLER_11_165 ();
 sg13g2_decap_8 FILLER_11_172 ();
 sg13g2_decap_8 FILLER_11_179 ();
 sg13g2_fill_1 FILLER_11_186 ();
 sg13g2_decap_8 FILLER_11_191 ();
 sg13g2_decap_8 FILLER_11_198 ();
 sg13g2_decap_8 FILLER_11_205 ();
 sg13g2_fill_1 FILLER_11_212 ();
 sg13g2_decap_8 FILLER_11_217 ();
 sg13g2_decap_8 FILLER_11_224 ();
 sg13g2_decap_8 FILLER_11_231 ();
 sg13g2_fill_1 FILLER_11_238 ();
 sg13g2_decap_8 FILLER_11_243 ();
 sg13g2_decap_8 FILLER_11_250 ();
 sg13g2_decap_8 FILLER_11_257 ();
 sg13g2_fill_1 FILLER_11_264 ();
 sg13g2_decap_8 FILLER_11_269 ();
 sg13g2_decap_8 FILLER_11_276 ();
 sg13g2_decap_8 FILLER_11_283 ();
 sg13g2_fill_1 FILLER_11_290 ();
 sg13g2_decap_8 FILLER_11_295 ();
 sg13g2_decap_8 FILLER_11_302 ();
 sg13g2_decap_8 FILLER_11_309 ();
 sg13g2_fill_1 FILLER_11_316 ();
 sg13g2_decap_8 FILLER_11_321 ();
 sg13g2_decap_8 FILLER_11_328 ();
 sg13g2_decap_8 FILLER_11_335 ();
 sg13g2_fill_1 FILLER_11_342 ();
 sg13g2_decap_8 FILLER_11_347 ();
 sg13g2_decap_8 FILLER_11_354 ();
 sg13g2_decap_8 FILLER_11_361 ();
 sg13g2_fill_1 FILLER_11_368 ();
 sg13g2_decap_8 FILLER_11_373 ();
 sg13g2_decap_8 FILLER_11_380 ();
 sg13g2_decap_8 FILLER_11_387 ();
 sg13g2_fill_1 FILLER_11_394 ();
 sg13g2_decap_8 FILLER_11_399 ();
 sg13g2_decap_8 FILLER_11_406 ();
 sg13g2_decap_8 FILLER_11_413 ();
 sg13g2_fill_1 FILLER_11_420 ();
 sg13g2_decap_8 FILLER_11_425 ();
 sg13g2_decap_8 FILLER_11_432 ();
 sg13g2_decap_8 FILLER_11_439 ();
 sg13g2_fill_1 FILLER_11_446 ();
 sg13g2_decap_8 FILLER_11_451 ();
 sg13g2_decap_8 FILLER_11_458 ();
 sg13g2_decap_8 FILLER_11_465 ();
 sg13g2_fill_1 FILLER_11_472 ();
 sg13g2_decap_8 FILLER_11_477 ();
 sg13g2_decap_8 FILLER_11_484 ();
 sg13g2_decap_8 FILLER_11_491 ();
 sg13g2_fill_1 FILLER_11_498 ();
 sg13g2_fill_1 FILLER_11_503 ();
endmodule
