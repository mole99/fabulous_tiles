* NGSPICE file created from N_term_single2.ext - technology: sky130A

* Black-box entry subcircuit for sky130_ef_sc_hd__decap_12 abstract view
.subckt sky130_ef_sc_hd__decap_12 VPWR VGND VPB VNB
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_2 abstract view
.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_1 abstract view
.subckt sky130_fd_sc_hd__buf_1 A VGND VNB VPB VPWR X
.ends

.subckt N_term_single2 FrameData[0] FrameData[10] FrameData[11] FrameData[12] FrameData[13]
+ FrameData[14] FrameData[15] FrameData[16] FrameData[17] FrameData[18] FrameData[19]
+ FrameData[1] FrameData[20] FrameData[21] FrameData[22] FrameData[23] FrameData[24]
+ FrameData[25] FrameData[26] FrameData[27] FrameData[28] FrameData[29] FrameData[2]
+ FrameData[30] FrameData[31] FrameData[3] FrameData[4] FrameData[5] FrameData[6]
+ FrameData[7] FrameData[8] FrameData[9] FrameData_O[0] FrameData_O[10] FrameData_O[11]
+ FrameData_O[12] FrameData_O[13] FrameData_O[14] FrameData_O[15] FrameData_O[16]
+ FrameData_O[17] FrameData_O[18] FrameData_O[19] FrameData_O[1] FrameData_O[20] FrameData_O[21]
+ FrameData_O[22] FrameData_O[23] FrameData_O[24] FrameData_O[25] FrameData_O[26]
+ FrameData_O[27] FrameData_O[28] FrameData_O[29] FrameData_O[2] FrameData_O[30] FrameData_O[31]
+ FrameData_O[3] FrameData_O[4] FrameData_O[5] FrameData_O[6] FrameData_O[7] FrameData_O[8]
+ FrameData_O[9] FrameStrobe[0] FrameStrobe[10] FrameStrobe[11] FrameStrobe[12] FrameStrobe[13]
+ FrameStrobe[14] FrameStrobe[15] FrameStrobe[16] FrameStrobe[17] FrameStrobe[18]
+ FrameStrobe[19] FrameStrobe[1] FrameStrobe[2] FrameStrobe[3] FrameStrobe[4] FrameStrobe[5]
+ FrameStrobe[6] FrameStrobe[7] FrameStrobe[8] FrameStrobe[9] FrameStrobe_O[0] FrameStrobe_O[10]
+ FrameStrobe_O[11] FrameStrobe_O[12] FrameStrobe_O[13] FrameStrobe_O[14] FrameStrobe_O[15]
+ FrameStrobe_O[16] FrameStrobe_O[17] FrameStrobe_O[18] FrameStrobe_O[19] FrameStrobe_O[1]
+ FrameStrobe_O[2] FrameStrobe_O[3] FrameStrobe_O[4] FrameStrobe_O[5] FrameStrobe_O[6]
+ FrameStrobe_O[7] FrameStrobe_O[8] FrameStrobe_O[9] N1END[0] N1END[1] N1END[2] N1END[3]
+ N2END[0] N2END[1] N2END[2] N2END[3] N2END[4] N2END[5] N2END[6] N2END[7] N2MID[0]
+ N2MID[1] N2MID[2] N2MID[3] N2MID[4] N2MID[5] N2MID[6] N2MID[7] N4END[0] N4END[10]
+ N4END[11] N4END[12] N4END[13] N4END[14] N4END[15] N4END[1] N4END[2] N4END[3] N4END[4]
+ N4END[5] N4END[6] N4END[7] N4END[8] N4END[9] NN4END[0] NN4END[10] NN4END[11] NN4END[12]
+ NN4END[13] NN4END[14] NN4END[15] NN4END[1] NN4END[2] NN4END[3] NN4END[4] NN4END[5]
+ NN4END[6] NN4END[7] NN4END[8] NN4END[9] S1BEG[0] S1BEG[1] S1BEG[2] S1BEG[3] S2BEG[0]
+ S2BEG[1] S2BEG[2] S2BEG[3] S2BEG[4] S2BEG[5] S2BEG[6] S2BEG[7] S2BEGb[0] S2BEGb[1]
+ S2BEGb[2] S2BEGb[3] S2BEGb[4] S2BEGb[5] S2BEGb[6] S2BEGb[7] S4BEG[0] S4BEG[10] S4BEG[11]
+ S4BEG[12] S4BEG[13] S4BEG[14] S4BEG[15] S4BEG[1] S4BEG[2] S4BEG[3] S4BEG[4] S4BEG[5]
+ S4BEG[6] S4BEG[7] S4BEG[8] S4BEG[9] SS4BEG[0] SS4BEG[10] SS4BEG[11] SS4BEG[12] SS4BEG[13]
+ SS4BEG[14] SS4BEG[15] SS4BEG[1] SS4BEG[2] SS4BEG[3] SS4BEG[4] SS4BEG[5] SS4BEG[6]
+ SS4BEG[7] SS4BEG[8] SS4BEG[9] UserCLK UserCLKo VGND VPWR
XFILLER_10_339 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_9_115 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_0_Left_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_11_142 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_140 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_11_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_062_ N2MID[1] VGND VGND VPWR VPWR net63 sky130_fd_sc_hd__clkbuf_1
XFILLER_9_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_045_ FrameStrobe[13] VGND VGND VPWR VPWR net37 sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_5_78 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_028_ FrameData[28] VGND VGND VPWR VPWR net21 sky130_fd_sc_hd__clkbuf_2
XANTENNA_5 FrameData[14] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput42 net42 VGND VGND VPWR VPWR FrameStrobe_O[18] sky130_fd_sc_hd__buf_2
Xoutput20 net20 VGND VGND VPWR VPWR FrameData_O[27] sky130_fd_sc_hd__buf_2
XFILLER_8_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput7 net7 VGND VGND VPWR VPWR FrameData_O[15] sky130_fd_sc_hd__buf_2
Xoutput64 net64 VGND VGND VPWR VPWR S2BEG[7] sky130_fd_sc_hd__buf_2
Xoutput53 net53 VGND VGND VPWR VPWR S1BEG[0] sky130_fd_sc_hd__buf_2
Xoutput86 net86 VGND VGND VPWR VPWR S4BEG[7] sky130_fd_sc_hd__buf_2
Xoutput75 net75 VGND VGND VPWR VPWR S4BEG[11] sky130_fd_sc_hd__buf_2
Xoutput97 net97 VGND VGND VPWR VPWR SS4BEG[2] sky130_fd_sc_hd__buf_2
Xoutput31 net31 VGND VGND VPWR VPWR FrameData_O[8] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_2_57 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_9_116 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_11_143 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_11_132 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_061_ N2MID[2] VGND VGND VPWR VPWR net62 sky130_fd_sc_hd__clkbuf_1
XFILLER_7_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_044_ FrameStrobe[12] VGND VGND VPWR VPWR net36 sky130_fd_sc_hd__buf_1
XFILLER_7_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_5_79 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_027_ FrameData[27] VGND VGND VPWR VPWR net20 sky130_fd_sc_hd__buf_1
XANTENNA_6 FrameData[15] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_6_Right_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput43 net43 VGND VGND VPWR VPWR FrameStrobe_O[19] sky130_fd_sc_hd__buf_2
Xoutput21 net21 VGND VGND VPWR VPWR FrameData_O[28] sky130_fd_sc_hd__buf_2
Xoutput8 net8 VGND VGND VPWR VPWR FrameData_O[16] sky130_fd_sc_hd__buf_2
Xoutput10 net10 VGND VGND VPWR VPWR FrameData_O[18] sky130_fd_sc_hd__buf_2
Xoutput65 net65 VGND VGND VPWR VPWR S2BEGb[0] sky130_fd_sc_hd__buf_2
XFILLER_0_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput54 net54 VGND VGND VPWR VPWR S1BEG[1] sky130_fd_sc_hd__buf_2
Xoutput87 net87 VGND VGND VPWR VPWR S4BEG[8] sky130_fd_sc_hd__buf_2
Xoutput76 net76 VGND VGND VPWR VPWR S4BEG[12] sky130_fd_sc_hd__buf_2
Xoutput98 net98 VGND VGND VPWR VPWR SS4BEG[3] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_2_58 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput32 net32 VGND VGND VPWR VPWR FrameData_O[9] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_9_117 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_301 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_8_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_11_144 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_11_133 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_370 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_11_458 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_060_ N2MID[3] VGND VGND VPWR VPWR net61 sky130_fd_sc_hd__clkbuf_1
XFILLER_7_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_11_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_043_ FrameStrobe[11] VGND VGND VPWR VPWR net35 sky130_fd_sc_hd__clkbuf_1
XFILLER_3_454 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_026_ FrameData[26] VGND VGND VPWR VPWR net19 sky130_fd_sc_hd__buf_1
XANTENNA_7 FrameData[16] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_6_90 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput44 net44 VGND VGND VPWR VPWR FrameStrobe_O[1] sky130_fd_sc_hd__buf_2
Xoutput33 net33 VGND VGND VPWR VPWR FrameStrobe_O[0] sky130_fd_sc_hd__buf_2
Xoutput22 net22 VGND VGND VPWR VPWR FrameData_O[29] sky130_fd_sc_hd__buf_2
Xoutput11 net11 VGND VGND VPWR VPWR FrameData_O[19] sky130_fd_sc_hd__buf_2
Xoutput9 net9 VGND VGND VPWR VPWR FrameData_O[17] sky130_fd_sc_hd__buf_2
Xoutput66 net66 VGND VGND VPWR VPWR S2BEGb[1] sky130_fd_sc_hd__buf_2
Xoutput55 net55 VGND VGND VPWR VPWR S1BEG[2] sky130_fd_sc_hd__buf_2
Xoutput88 net88 VGND VGND VPWR VPWR S4BEG[9] sky130_fd_sc_hd__buf_2
Xoutput77 net77 VGND VGND VPWR VPWR S4BEG[13] sky130_fd_sc_hd__buf_2
Xoutput99 net99 VGND VGND VPWR VPWR SS4BEG[4] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_2_59 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_009_ FrameData[9] VGND VGND VPWR VPWR net32 sky130_fd_sc_hd__buf_1
XFILLER_8_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_8_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_9_118 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_313 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_3_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_10_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_11_145 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_11_134 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_4_Left_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_11_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_042_ FrameStrobe[10] VGND VGND VPWR VPWR net34 sky130_fd_sc_hd__buf_1
XFILLER_7_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_3_466 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_025_ FrameData[25] VGND VGND VPWR VPWR net18 sky130_fd_sc_hd__clkbuf_1
XFILLER_6_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_8 FrameData[18] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_6_91 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput34 net34 VGND VGND VPWR VPWR FrameStrobe_O[10] sky130_fd_sc_hd__buf_2
Xoutput45 net45 VGND VGND VPWR VPWR FrameStrobe_O[2] sky130_fd_sc_hd__buf_2
Xoutput56 net56 VGND VGND VPWR VPWR S1BEG[3] sky130_fd_sc_hd__buf_2
Xoutput67 net67 VGND VGND VPWR VPWR S2BEGb[2] sky130_fd_sc_hd__buf_2
Xoutput78 net78 VGND VGND VPWR VPWR S4BEG[14] sky130_fd_sc_hd__buf_2
Xoutput89 net89 VGND VGND VPWR VPWR SS4BEG[0] sky130_fd_sc_hd__buf_2
Xoutput23 net23 VGND VGND VPWR VPWR FrameData_O[2] sky130_fd_sc_hd__buf_2
Xoutput12 net12 VGND VGND VPWR VPWR FrameData_O[1] sky130_fd_sc_hd__buf_2
XFILLER_11_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_8_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_008_ FrameData[8] VGND VGND VPWR VPWR net31 sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_9_119 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_8_163 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_8_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_11_146 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_11_135 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_11_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_6_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_041_ FrameStrobe[9] VGND VGND VPWR VPWR net52 sky130_fd_sc_hd__clkbuf_1
XFILLER_7_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_478 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_024_ FrameData[24] VGND VGND VPWR VPWR net17 sky130_fd_sc_hd__buf_1
XTAP_TAPCELL_ROW_6_92 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_9 FrameData[19] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xoutput35 net35 VGND VGND VPWR VPWR FrameStrobe_O[11] sky130_fd_sc_hd__buf_2
Xoutput46 net46 VGND VGND VPWR VPWR FrameStrobe_O[3] sky130_fd_sc_hd__buf_2
Xoutput24 net24 VGND VGND VPWR VPWR FrameData_O[30] sky130_fd_sc_hd__buf_2
Xoutput13 net13 VGND VGND VPWR VPWR FrameData_O[20] sky130_fd_sc_hd__buf_2
Xoutput57 net57 VGND VGND VPWR VPWR S2BEG[0] sky130_fd_sc_hd__buf_2
XFILLER_8_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_8_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput68 net68 VGND VGND VPWR VPWR S2BEGb[3] sky130_fd_sc_hd__buf_2
Xoutput79 net79 VGND VGND VPWR VPWR S4BEG[15] sky130_fd_sc_hd__buf_2
X_007_ FrameData[7] VGND VGND VPWR VPWR net30 sky130_fd_sc_hd__clkbuf_1
XFILLER_7_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_5_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_3_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_8_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_8_175 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_8_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_3_60 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_11_147 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_11_136 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_71 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_9_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_6_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_9_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_11_258 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_11_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_040_ FrameStrobe[8] VGND VGND VPWR VPWR net51 sky130_fd_sc_hd__clkbuf_1
XFILLER_1_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_023_ FrameData[23] VGND VGND VPWR VPWR net16 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_6_93 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput36 net36 VGND VGND VPWR VPWR FrameStrobe_O[12] sky130_fd_sc_hd__buf_2
Xoutput47 net47 VGND VGND VPWR VPWR FrameStrobe_O[4] sky130_fd_sc_hd__buf_2
Xoutput25 net25 VGND VGND VPWR VPWR FrameData_O[31] sky130_fd_sc_hd__buf_2
Xoutput14 net14 VGND VGND VPWR VPWR FrameData_O[21] sky130_fd_sc_hd__buf_2
XFILLER_8_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xoutput58 net58 VGND VGND VPWR VPWR S2BEG[1] sky130_fd_sc_hd__buf_2
Xoutput69 net69 VGND VGND VPWR VPWR S2BEGb[4] sky130_fd_sc_hd__buf_2
X_006_ FrameData[6] VGND VGND VPWR VPWR net29 sky130_fd_sc_hd__clkbuf_1
XFILLER_7_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_8_110 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_8_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_3_61 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_11_148 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_11_137 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_6_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_9_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_6_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_0_40 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_099_ NN4END[4] VGND VGND VPWR VPWR net91 sky130_fd_sc_hd__buf_1
XFILLER_1_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_022_ FrameData[22] VGND VGND VPWR VPWR net15 sky130_fd_sc_hd__buf_1
XFILLER_6_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_6_94 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput37 net37 VGND VGND VPWR VPWR FrameStrobe_O[13] sky130_fd_sc_hd__buf_2
Xoutput48 net48 VGND VGND VPWR VPWR FrameStrobe_O[5] sky130_fd_sc_hd__buf_2
Xoutput15 net15 VGND VGND VPWR VPWR FrameData_O[22] sky130_fd_sc_hd__buf_2
Xoutput59 net59 VGND VGND VPWR VPWR S2BEG[2] sky130_fd_sc_hd__buf_2
XFILLER_0_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput26 net26 VGND VGND VPWR VPWR FrameData_O[3] sky130_fd_sc_hd__buf_2
XPHY_EDGE_ROW_1_Right_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_005_ FrameData[5] VGND VGND VPWR VPWR net28 sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_8_111 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_3_62 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_11_149 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_11_138 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_408 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_430 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_6_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_6_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_0_30 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_41 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_098_ NN4END[5] VGND VGND VPWR VPWR net90 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_10_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_021_ FrameData[21] VGND VGND VPWR VPWR net14 sky130_fd_sc_hd__clkbuf_2
XPHY_EDGE_ROW_11_Left_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_6_95 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput38 net38 VGND VGND VPWR VPWR FrameStrobe_O[14] sky130_fd_sc_hd__buf_2
Xoutput49 net49 VGND VGND VPWR VPWR FrameStrobe_O[6] sky130_fd_sc_hd__buf_2
Xoutput16 net16 VGND VGND VPWR VPWR FrameData_O[23] sky130_fd_sc_hd__buf_2
Xoutput27 net27 VGND VGND VPWR VPWR FrameData_O[4] sky130_fd_sc_hd__buf_2
XFILLER_11_7 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_004_ FrameData[4] VGND VGND VPWR VPWR net27 sky130_fd_sc_hd__buf_1
XFILLER_7_370 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_7_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_8_112 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_3_63 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_11_139 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_10_442 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_6_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_6_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_0_31 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_6_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_097_ NN4END[6] VGND VGND VPWR VPWR net104 sky130_fd_sc_hd__buf_1
XFILLER_10_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_020_ FrameData[20] VGND VGND VPWR VPWR net13 sky130_fd_sc_hd__buf_1
XFILLER_3_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput17 net17 VGND VGND VPWR VPWR FrameData_O[24] sky130_fd_sc_hd__buf_2
Xoutput39 net39 VGND VGND VPWR VPWR FrameStrobe_O[15] sky130_fd_sc_hd__buf_2
Xoutput28 net28 VGND VGND VPWR VPWR FrameData_O[5] sky130_fd_sc_hd__buf_2
X_003_ FrameData[3] VGND VGND VPWR VPWR net26 sky130_fd_sc_hd__buf_1
XFILLER_7_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_7_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_8_113 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_3_64 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_10_454 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_10_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_0_32 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_428 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_10_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_096_ NN4END[7] VGND VGND VPWR VPWR net103 sky130_fd_sc_hd__buf_1
XFILLER_10_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_10_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_3_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput18 net18 VGND VGND VPWR VPWR FrameData_O[25] sky130_fd_sc_hd__buf_2
X_079_ N4END[8] VGND VGND VPWR VPWR net86 sky130_fd_sc_hd__buf_1
Xoutput29 net29 VGND VGND VPWR VPWR FrameData_O[6] sky130_fd_sc_hd__buf_2
XFILLER_2_280 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_002_ FrameData[2] VGND VGND VPWR VPWR net23 sky130_fd_sc_hd__buf_1
XPHY_EDGE_ROW_5_Right_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_3_65 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_10_130 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_434 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_9_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_0_33 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_242 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_11_208 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_095_ NN4END[8] VGND VGND VPWR VPWR net102 sky130_fd_sc_hd__clkbuf_1
XFILLER_6_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_6_87 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_078_ N4END[9] VGND VGND VPWR VPWR net85 sky130_fd_sc_hd__buf_1
XFILLER_2_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput19 net19 VGND VGND VPWR VPWR FrameData_O[26] sky130_fd_sc_hd__buf_2
XFILLER_8_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_001_ FrameData[1] VGND VGND VPWR VPWR net12 sky130_fd_sc_hd__buf_1
XFILLER_11_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_11_Right_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_3_66 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_5_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_10_131 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_254 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_9_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_0_34 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_3_Left_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_094_ NN4END[9] VGND VGND VPWR VPWR net101 sky130_fd_sc_hd__buf_1
XFILLER_10_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_077_ N4END[10] VGND VGND VPWR VPWR net84 sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_6_88 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_000_ FrameData[0] VGND VGND VPWR VPWR net1 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_8_105 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_3_67 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_5_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_358 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_10_402 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_9_266 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_8_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_0_24 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_35 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_093_ NN4END[10] VGND VGND VPWR VPWR net100 sky130_fd_sc_hd__clkbuf_1
XFILLER_10_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_206 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_6_89 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_076_ N4END[11] VGND VGND VPWR VPWR net83 sky130_fd_sc_hd__buf_1
XFILLER_0_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_11_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_059_ N2MID[4] VGND VGND VPWR VPWR net60 sky130_fd_sc_hd__buf_1
XFILLER_8_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_8_106 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_3_68 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_9_Right_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_10_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_0_25 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_36 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_10_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_092_ NN4END[11] VGND VGND VPWR VPWR net99 sky130_fd_sc_hd__clkbuf_1
XFILLER_1_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_3_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_075_ N4END[12] VGND VGND VPWR VPWR net82 sky130_fd_sc_hd__clkbuf_1
XANTENNA_40 net81 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_058_ N2MID[5] VGND VGND VPWR VPWR net59 sky130_fd_sc_hd__buf_1
XTAP_TAPCELL_ROW_8_107 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_10_123 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_9_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_0_26 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_37 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_6_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_091_ NN4END[12] VGND VGND VPWR VPWR net98 sky130_fd_sc_hd__buf_1
XFILLER_1_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_7_Left_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_13 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_074_ N4END[13] VGND VGND VPWR VPWR net81 sky130_fd_sc_hd__buf_1
XFILLER_2_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_30 FrameStrobe[8] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_41 net83 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_057_ N2MID[6] VGND VGND VPWR VPWR net58 sky130_fd_sc_hd__buf_1
XTAP_TAPCELL_ROW_8_108 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_0_Right_0 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_10_124 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_59 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_147 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_0_27 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_38 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_5_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_090_ NN4END[13] VGND VGND VPWR VPWR net97 sky130_fd_sc_hd__clkbuf_1
XFILLER_6_217 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_6_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_10_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_073_ N4END[14] VGND VGND VPWR VPWR net80 sky130_fd_sc_hd__buf_1
XANTENNA_20 FrameData[31] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_31 N2END[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_42 net85 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_056_ N2MID[7] VGND VGND VPWR VPWR net57 sky130_fd_sc_hd__buf_1
XPHY_EDGE_ROW_10_Left_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_8_109 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_039_ FrameStrobe[7] VGND VGND VPWR VPWR net50 sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_10_125 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_440 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_4_70 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_0_28 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_0_39 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_10_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_229 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_5_262 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_5_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_072_ N4END[15] VGND VGND VPWR VPWR net73 sky130_fd_sc_hd__clkbuf_1
XFILLER_2_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_21 FrameData[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_10 FrameData[20] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_43 net86 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_32 N4END[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_055_ N1END[0] VGND VGND VPWR VPWR net56 sky130_fd_sc_hd__clkbuf_1
XFILLER_7_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_11_183 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_038_ FrameStrobe[6] VGND VGND VPWR VPWR net49 sky130_fd_sc_hd__clkbuf_1
XFILLER_3_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_10_126 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_452 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_4_71 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_29 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_1_50 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_071_ N2END[0] VGND VGND VPWR VPWR net72 sky130_fd_sc_hd__clkbuf_1
XFILLER_2_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_44 FrameStrobe[9] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_11 FrameData[21] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_22 FrameData[4] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_33 N4END[6] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_054_ N1END[1] VGND VGND VPWR VPWR net55 sky130_fd_sc_hd__buf_1
XFILLER_7_358 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_7_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_11_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_037_ FrameStrobe[5] VGND VGND VPWR VPWR net48 sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_7_100 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_4_Right_4 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_10_127 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_4_72 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_283 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_5_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_256 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_070_ N2END[1] VGND VGND VPWR VPWR net71 sky130_fd_sc_hd__clkbuf_1
XFILLER_4_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_12 FrameData[22] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_45 N2END[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_34 N4END[7] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_23 FrameData[5] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_053_ N1END[2] VGND VGND VPWR VPWR net54 sky130_fd_sc_hd__buf_1
XFILLER_11_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_7_101 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_036_ FrameStrobe[4] VGND VGND VPWR VPWR net47 sky130_fd_sc_hd__clkbuf_1
XFILLER_8_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_10_128 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_019_ FrameData[19] VGND VGND VPWR VPWR net11 sky130_fd_sc_hd__buf_1
XTAP_TAPCELL_ROW_4_73 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_295 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_8_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_2_Left_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_268 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_35 NN4END[11] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_13 FrameData[23] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_46 N4END[12] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_24 FrameData[6] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_61 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_7_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_052_ N1END[3] VGND VGND VPWR VPWR net53 sky130_fd_sc_hd__buf_1
XTAP_TAPCELL_ROW_7_102 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_104_ UserCLK VGND VGND VPWR VPWR net105 sky130_fd_sc_hd__buf_2
X_035_ FrameStrobe[3] VGND VGND VPWR VPWR net46 sky130_fd_sc_hd__clkbuf_1
XFILLER_7_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_3_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_10_129 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_4_74 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_018_ FrameData[18] VGND VGND VPWR VPWR net10 sky130_fd_sc_hd__clkbuf_2
XFILLER_5_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_10_229 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_10_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_1_42 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_10_Right_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_14 FrameData[24] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_36 NN4END[13] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_25 FrameData[7] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_051_ FrameStrobe[19] VGND VGND VPWR VPWR net43 sky130_fd_sc_hd__clkbuf_1
XFILLER_7_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_6_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_7_96 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_7_103 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_034_ FrameStrobe[2] VGND VGND VPWR VPWR net45 sky130_fd_sc_hd__clkbuf_1
XFILLER_7_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_7_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_103_ NN4END[0] VGND VGND VPWR VPWR net95 sky130_fd_sc_hd__clkbuf_2
XFILLER_8_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_8_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_8_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_8_Right_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_017_ FrameData[17] VGND VGND VPWR VPWR net9 sky130_fd_sc_hd__buf_1
XTAP_TAPCELL_ROW_4_75 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_194 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_9_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_8_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_5_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_5_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_5_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_1_43 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_15 FrameData[25] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_37 NN4END[14] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_26 FrameData[8] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_050_ FrameStrobe[18] VGND VGND VPWR VPWR net42 sky130_fd_sc_hd__clkbuf_1
XFILLER_7_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xoutput100 net100 VGND VGND VPWR VPWR SS4BEG[5] sky130_fd_sc_hd__buf_2
XFILLER_11_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_7_97 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_7_104 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_033_ FrameStrobe[1] VGND VGND VPWR VPWR net44 sky130_fd_sc_hd__clkbuf_2
XFILLER_7_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_102_ NN4END[1] VGND VGND VPWR VPWR net94 sky130_fd_sc_hd__buf_1
XFILLER_8_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_8_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_6_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_4_76 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_016_ FrameData[16] VGND VGND VPWR VPWR net8 sky130_fd_sc_hd__clkbuf_2
XFILLER_8_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_5_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_5_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_1_44 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_38 NN4END[8] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_16 FrameData[26] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_27 net10 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_6_Left_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput101 net101 VGND VGND VPWR VPWR SS4BEG[6] sky130_fd_sc_hd__buf_2
XFILLER_11_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_7_98 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_032_ FrameStrobe[0] VGND VGND VPWR VPWR net33 sky130_fd_sc_hd__clkbuf_2
XFILLER_7_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_7_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_101_ NN4END[2] VGND VGND VPWR VPWR net93 sky130_fd_sc_hd__buf_1
XFILLER_8_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_9_Left_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_4_77 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_015_ FrameData[15] VGND VGND VPWR VPWR net7 sky130_fd_sc_hd__clkbuf_2
XFILLER_5_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_10_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_5_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_1_45 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_39 NN4END[9] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_17 FrameData[27] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_28 FrameStrobe[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xoutput102 net102 VGND VGND VPWR VPWR SS4BEG[7] sky130_fd_sc_hd__buf_2
XFILLER_11_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_7_99 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_031_ FrameData[31] VGND VGND VPWR VPWR net25 sky130_fd_sc_hd__clkbuf_1
X_100_ NN4END[3] VGND VGND VPWR VPWR net92 sky130_fd_sc_hd__buf_1
XFILLER_8_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_161 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_8_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_014_ FrameData[14] VGND VGND VPWR VPWR net6 sky130_fd_sc_hd__clkbuf_2
XFILLER_5_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_8_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_1_46 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_29 FrameStrobe[4] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_18 FrameData[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xoutput103 net103 VGND VGND VPWR VPWR SS4BEG[8] sky130_fd_sc_hd__buf_2
XFILLER_11_33 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_6_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_6_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_11_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_030_ FrameData[30] VGND VGND VPWR VPWR net24 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_3_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_013_ FrameData[13] VGND VGND VPWR VPWR net5 sky130_fd_sc_hd__buf_1
XFILLER_0_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_5_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_5_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_1_47 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_352 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_19 FrameData[30] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_230 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput104 net104 VGND VGND VPWR VPWR SS4BEG[9] sky130_fd_sc_hd__buf_2
XFILLER_11_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_351 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_6_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_6_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_089_ NN4END[14] VGND VGND VPWR VPWR net96 sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_4_69 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_012_ FrameData[12] VGND VGND VPWR VPWR net4 sky130_fd_sc_hd__buf_1
XPHY_EDGE_ROW_3_Right_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_5_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_1_48 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_283 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_9_364 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_242 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_297 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput105 net105 VGND VGND VPWR VPWR UserCLKo sky130_fd_sc_hd__buf_1
XFILLER_10_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_6_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_6_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_088_ NN4END[15] VGND VGND VPWR VPWR net89 sky130_fd_sc_hd__clkbuf_1
X_011_ FrameData[11] VGND VGND VPWR VPWR net3 sky130_fd_sc_hd__buf_1
XFILLER_3_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_462 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_5_80 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_1_49 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_295 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_9_376 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_10_375 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_1_Left_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_3_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_8_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_6_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_087_ N4END[0] VGND VGND VPWR VPWR net79 sky130_fd_sc_hd__clkbuf_1
XFILLER_8_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_010_ FrameData[10] VGND VGND VPWR VPWR net2 sky130_fd_sc_hd__clkbuf_1
XFILLER_11_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_474 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_7_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_5_81 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_7_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_414 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_9_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_9_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_152 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_9_185 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_5_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_086_ N4END[1] VGND VGND VPWR VPWR net78 sky130_fd_sc_hd__clkbuf_1
XFILLER_3_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_3_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_3_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_7_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_069_ N2END[2] VGND VGND VPWR VPWR net70 sky130_fd_sc_hd__clkbuf_1
XFILLER_9_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_5_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_7_Right_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_5_82 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_426 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_9_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput90 net90 VGND VGND VPWR VPWR SS4BEG[10] sky130_fd_sc_hd__buf_2
XFILLER_2_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_11_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_9_120 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_9_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_3_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_085_ N4END[2] VGND VGND VPWR VPWR net77 sky130_fd_sc_hd__clkbuf_1
XFILLER_2_351 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_3_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_11_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_068_ N2END[3] VGND VGND VPWR VPWR net69 sky130_fd_sc_hd__clkbuf_1
XFILLER_9_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_5_83 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_6_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput1 net1 VGND VGND VPWR VPWR FrameData_O[0] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_2_51 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput80 net80 VGND VGND VPWR VPWR S4BEG[1] sky130_fd_sc_hd__buf_2
Xoutput91 net91 VGND VGND VPWR VPWR SS4BEG[11] sky130_fd_sc_hd__buf_2
XFILLER_10_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_9_121 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_5_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_3_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_5_Left_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_164 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_10_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_084_ N4END[3] VGND VGND VPWR VPWR net76 sky130_fd_sc_hd__clkbuf_1
XFILLER_2_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_067_ N2END[4] VGND VGND VPWR VPWR net68 sky130_fd_sc_hd__buf_1
XPHY_EDGE_ROW_8_Left_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_230 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_5_84 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_200 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput70 net70 VGND VGND VPWR VPWR S2BEGb[5] sky130_fd_sc_hd__buf_2
Xoutput81 net81 VGND VGND VPWR VPWR S4BEG[2] sky130_fd_sc_hd__buf_2
Xoutput92 net92 VGND VGND VPWR VPWR SS4BEG[12] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_2_52 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput2 net2 VGND VGND VPWR VPWR FrameData_O[10] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_9_122 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_9_122 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_9_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_10_176 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_10_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_083_ N4END[4] VGND VGND VPWR VPWR net75 sky130_fd_sc_hd__clkbuf_1
XFILLER_2_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_066_ N2END[5] VGND VGND VPWR VPWR net67 sky130_fd_sc_hd__buf_1
XFILLER_8_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_049_ FrameStrobe[17] VGND VGND VPWR VPWR net41 sky130_fd_sc_hd__clkbuf_1
XFILLER_7_242 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_5_85 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_6_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_1 FrameData[10] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_204 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_9_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xoutput3 net3 VGND VGND VPWR VPWR FrameData_O[11] sky130_fd_sc_hd__buf_2
Xoutput60 net60 VGND VGND VPWR VPWR S2BEG[3] sky130_fd_sc_hd__buf_2
Xoutput71 net71 VGND VGND VPWR VPWR S2BEGb[6] sky130_fd_sc_hd__buf_2
Xoutput82 net82 VGND VGND VPWR VPWR S4BEG[3] sky130_fd_sc_hd__buf_2
Xoutput93 net93 VGND VGND VPWR VPWR SS4BEG[13] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_2_53 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_134 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_5_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_86 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_10_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_100 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_082_ N4END[5] VGND VGND VPWR VPWR net74 sky130_fd_sc_hd__clkbuf_1
XFILLER_2_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_5_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_11_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_065_ N2END[6] VGND VGND VPWR VPWR net66 sky130_fd_sc_hd__buf_1
XFILLER_7_254 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_5_86 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_048_ FrameStrobe[16] VGND VGND VPWR VPWR net40 sky130_fd_sc_hd__clkbuf_1
XANTENNA_2 FrameData[11] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_6_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xoutput50 net50 VGND VGND VPWR VPWR FrameStrobe_O[7] sky130_fd_sc_hd__buf_2
XFILLER_9_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput4 net4 VGND VGND VPWR VPWR FrameData_O[12] sky130_fd_sc_hd__buf_2
Xoutput61 net61 VGND VGND VPWR VPWR S2BEG[4] sky130_fd_sc_hd__buf_2
Xoutput72 net72 VGND VGND VPWR VPWR S2BEGb[7] sky130_fd_sc_hd__buf_2
Xoutput83 net83 VGND VGND VPWR VPWR S4BEG[4] sky130_fd_sc_hd__buf_2
Xoutput94 net94 VGND VGND VPWR VPWR SS4BEG[14] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_2_54 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_315 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_9_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_98 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_10_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_081_ N4END[6] VGND VGND VPWR VPWR net88 sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_11_140 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_11_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_064_ N2END[7] VGND VGND VPWR VPWR net65 sky130_fd_sc_hd__buf_1
XFILLER_11_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_047_ FrameStrobe[15] VGND VGND VPWR VPWR net39 sky130_fd_sc_hd__clkbuf_1
XFILLER_7_266 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_2_Right_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_3 FrameData[12] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput40 net40 VGND VGND VPWR VPWR FrameStrobe_O[16] sky130_fd_sc_hd__buf_2
Xoutput51 net51 VGND VGND VPWR VPWR FrameStrobe_O[8] sky130_fd_sc_hd__buf_2
XFILLER_9_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput5 net5 VGND VGND VPWR VPWR FrameData_O[13] sky130_fd_sc_hd__buf_2
Xoutput62 net62 VGND VGND VPWR VPWR S2BEG[5] sky130_fd_sc_hd__buf_2
Xoutput73 net73 VGND VGND VPWR VPWR S4BEG[0] sky130_fd_sc_hd__buf_2
Xoutput84 net84 VGND VGND VPWR VPWR S4BEG[5] sky130_fd_sc_hd__buf_2
Xoutput95 net95 VGND VGND VPWR VPWR SS4BEG[15] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_2_55 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_327 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_9_114 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_9_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_3_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_080_ N4END[7] VGND VGND VPWR VPWR net87 sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_11_141 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_11_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_063_ N2MID[0] VGND VGND VPWR VPWR net64 sky130_fd_sc_hd__clkbuf_1
XFILLER_2_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_11_285 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_046_ FrameStrobe[14] VGND VGND VPWR VPWR net38 sky130_fd_sc_hd__clkbuf_1
XFILLER_7_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_029_ FrameData[29] VGND VGND VPWR VPWR net22 sky130_fd_sc_hd__clkbuf_2
XANTENNA_4 FrameData[13] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput41 net41 VGND VGND VPWR VPWR FrameStrobe_O[17] sky130_fd_sc_hd__buf_2
Xoutput52 net52 VGND VGND VPWR VPWR FrameStrobe_O[9] sky130_fd_sc_hd__buf_2
XFILLER_9_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xoutput6 net6 VGND VGND VPWR VPWR FrameData_O[14] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_2_56 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput30 net30 VGND VGND VPWR VPWR FrameData_O[7] sky130_fd_sc_hd__buf_2
Xoutput63 net63 VGND VGND VPWR VPWR S2BEG[6] sky130_fd_sc_hd__buf_2
Xoutput85 net85 VGND VGND VPWR VPWR S4BEG[6] sky130_fd_sc_hd__buf_2
Xoutput74 net74 VGND VGND VPWR VPWR S4BEG[10] sky130_fd_sc_hd__buf_2
Xoutput96 net96 VGND VGND VPWR VPWR SS4BEG[1] sky130_fd_sc_hd__buf_2
.ends

