module EF_SRAM (AD_SRAM0,
    AD_SRAM1,
    AD_SRAM2,
    AD_SRAM3,
    AD_SRAM4,
    AD_SRAM5,
    AD_SRAM6,
    AD_SRAM7,
    AD_SRAM8,
    AD_SRAM9,
    BEN_SRAM0,
    BEN_SRAM1,
    BEN_SRAM10,
    BEN_SRAM11,
    BEN_SRAM12,
    BEN_SRAM13,
    BEN_SRAM14,
    BEN_SRAM15,
    BEN_SRAM16,
    BEN_SRAM17,
    BEN_SRAM18,
    BEN_SRAM19,
    BEN_SRAM2,
    BEN_SRAM20,
    BEN_SRAM21,
    BEN_SRAM22,
    BEN_SRAM23,
    BEN_SRAM24,
    BEN_SRAM25,
    BEN_SRAM26,
    BEN_SRAM27,
    BEN_SRAM28,
    BEN_SRAM29,
    BEN_SRAM3,
    BEN_SRAM30,
    BEN_SRAM31,
    BEN_SRAM4,
    BEN_SRAM5,
    BEN_SRAM6,
    BEN_SRAM7,
    BEN_SRAM8,
    BEN_SRAM9,
    CLOCK_SRAM,
    DI_SRAM0,
    DI_SRAM1,
    DI_SRAM10,
    DI_SRAM11,
    DI_SRAM12,
    DI_SRAM13,
    DI_SRAM14,
    DI_SRAM15,
    DI_SRAM16,
    DI_SRAM17,
    DI_SRAM18,
    DI_SRAM19,
    DI_SRAM2,
    DI_SRAM20,
    DI_SRAM21,
    DI_SRAM22,
    DI_SRAM23,
    DI_SRAM24,
    DI_SRAM25,
    DI_SRAM26,
    DI_SRAM27,
    DI_SRAM28,
    DI_SRAM29,
    DI_SRAM3,
    DI_SRAM30,
    DI_SRAM31,
    DI_SRAM4,
    DI_SRAM5,
    DI_SRAM6,
    DI_SRAM7,
    DI_SRAM8,
    DI_SRAM9,
    DO_SRAM0,
    DO_SRAM1,
    DO_SRAM10,
    DO_SRAM11,
    DO_SRAM12,
    DO_SRAM13,
    DO_SRAM14,
    DO_SRAM15,
    DO_SRAM16,
    DO_SRAM17,
    DO_SRAM18,
    DO_SRAM19,
    DO_SRAM2,
    DO_SRAM20,
    DO_SRAM21,
    DO_SRAM22,
    DO_SRAM23,
    DO_SRAM24,
    DO_SRAM25,
    DO_SRAM26,
    DO_SRAM27,
    DO_SRAM28,
    DO_SRAM29,
    DO_SRAM3,
    DO_SRAM30,
    DO_SRAM31,
    DO_SRAM4,
    DO_SRAM5,
    DO_SRAM6,
    DO_SRAM7,
    DO_SRAM8,
    DO_SRAM9,
    EN_SRAM,
    R_WB_SRAM,
    Tile_X0Y0_UserCLKo,
    Tile_X0Y1_UserCLK,
    Tile_X0Y0_E1END,
    Tile_X0Y0_E2END,
    Tile_X0Y0_E2MID,
    Tile_X0Y0_E6END,
    Tile_X0Y0_EE4END,
    Tile_X0Y0_FrameData,
    Tile_X0Y0_FrameData_O,
    Tile_X0Y0_FrameStrobe_O,
    Tile_X0Y0_N1BEG,
    Tile_X0Y0_N2BEG,
    Tile_X0Y0_N2BEGb,
    Tile_X0Y0_N4BEG,
    Tile_X0Y0_S1END,
    Tile_X0Y0_S2END,
    Tile_X0Y0_S2MID,
    Tile_X0Y0_S4END,
    Tile_X0Y0_W1BEG,
    Tile_X0Y0_W2BEG,
    Tile_X0Y0_W2BEGb,
    Tile_X0Y0_W6BEG,
    Tile_X0Y0_WW4BEG,
    Tile_X0Y1_E1END,
    Tile_X0Y1_E2END,
    Tile_X0Y1_E2MID,
    Tile_X0Y1_E6END,
    Tile_X0Y1_EE4END,
    Tile_X0Y1_FrameData,
    Tile_X0Y1_FrameData_O,
    Tile_X0Y1_FrameStrobe,
    Tile_X0Y1_N1END,
    Tile_X0Y1_N2END,
    Tile_X0Y1_N2MID,
    Tile_X0Y1_N4END,
    Tile_X0Y1_S1BEG,
    Tile_X0Y1_S2BEG,
    Tile_X0Y1_S2BEGb,
    Tile_X0Y1_S4BEG,
    Tile_X0Y1_W1BEG,
    Tile_X0Y1_W2BEG,
    Tile_X0Y1_W2BEGb,
    Tile_X0Y1_W6BEG,
    Tile_X0Y1_WW4BEG);
 output AD_SRAM0;
 output AD_SRAM1;
 output AD_SRAM2;
 output AD_SRAM3;
 output AD_SRAM4;
 output AD_SRAM5;
 output AD_SRAM6;
 output AD_SRAM7;
 output AD_SRAM8;
 output AD_SRAM9;
 output BEN_SRAM0;
 output BEN_SRAM1;
 output BEN_SRAM10;
 output BEN_SRAM11;
 output BEN_SRAM12;
 output BEN_SRAM13;
 output BEN_SRAM14;
 output BEN_SRAM15;
 output BEN_SRAM16;
 output BEN_SRAM17;
 output BEN_SRAM18;
 output BEN_SRAM19;
 output BEN_SRAM2;
 output BEN_SRAM20;
 output BEN_SRAM21;
 output BEN_SRAM22;
 output BEN_SRAM23;
 output BEN_SRAM24;
 output BEN_SRAM25;
 output BEN_SRAM26;
 output BEN_SRAM27;
 output BEN_SRAM28;
 output BEN_SRAM29;
 output BEN_SRAM3;
 output BEN_SRAM30;
 output BEN_SRAM31;
 output BEN_SRAM4;
 output BEN_SRAM5;
 output BEN_SRAM6;
 output BEN_SRAM7;
 output BEN_SRAM8;
 output BEN_SRAM9;
 output CLOCK_SRAM;
 output DI_SRAM0;
 output DI_SRAM1;
 output DI_SRAM10;
 output DI_SRAM11;
 output DI_SRAM12;
 output DI_SRAM13;
 output DI_SRAM14;
 output DI_SRAM15;
 output DI_SRAM16;
 output DI_SRAM17;
 output DI_SRAM18;
 output DI_SRAM19;
 output DI_SRAM2;
 output DI_SRAM20;
 output DI_SRAM21;
 output DI_SRAM22;
 output DI_SRAM23;
 output DI_SRAM24;
 output DI_SRAM25;
 output DI_SRAM26;
 output DI_SRAM27;
 output DI_SRAM28;
 output DI_SRAM29;
 output DI_SRAM3;
 output DI_SRAM30;
 output DI_SRAM31;
 output DI_SRAM4;
 output DI_SRAM5;
 output DI_SRAM6;
 output DI_SRAM7;
 output DI_SRAM8;
 output DI_SRAM9;
 input DO_SRAM0;
 input DO_SRAM1;
 input DO_SRAM10;
 input DO_SRAM11;
 input DO_SRAM12;
 input DO_SRAM13;
 input DO_SRAM14;
 input DO_SRAM15;
 input DO_SRAM16;
 input DO_SRAM17;
 input DO_SRAM18;
 input DO_SRAM19;
 input DO_SRAM2;
 input DO_SRAM20;
 input DO_SRAM21;
 input DO_SRAM22;
 input DO_SRAM23;
 input DO_SRAM24;
 input DO_SRAM25;
 input DO_SRAM26;
 input DO_SRAM27;
 input DO_SRAM28;
 input DO_SRAM29;
 input DO_SRAM3;
 input DO_SRAM30;
 input DO_SRAM31;
 input DO_SRAM4;
 input DO_SRAM5;
 input DO_SRAM6;
 input DO_SRAM7;
 input DO_SRAM8;
 input DO_SRAM9;
 output EN_SRAM;
 output R_WB_SRAM;
 output Tile_X0Y0_UserCLKo;
 input Tile_X0Y1_UserCLK;
 input [3:0] Tile_X0Y0_E1END;
 input [7:0] Tile_X0Y0_E2END;
 input [7:0] Tile_X0Y0_E2MID;
 input [11:0] Tile_X0Y0_E6END;
 input [15:0] Tile_X0Y0_EE4END;
 input [31:0] Tile_X0Y0_FrameData;
 output [31:0] Tile_X0Y0_FrameData_O;
 output [19:0] Tile_X0Y0_FrameStrobe_O;
 output [3:0] Tile_X0Y0_N1BEG;
 output [7:0] Tile_X0Y0_N2BEG;
 output [7:0] Tile_X0Y0_N2BEGb;
 output [15:0] Tile_X0Y0_N4BEG;
 input [3:0] Tile_X0Y0_S1END;
 input [7:0] Tile_X0Y0_S2END;
 input [7:0] Tile_X0Y0_S2MID;
 input [15:0] Tile_X0Y0_S4END;
 output [3:0] Tile_X0Y0_W1BEG;
 output [7:0] Tile_X0Y0_W2BEG;
 output [7:0] Tile_X0Y0_W2BEGb;
 output [11:0] Tile_X0Y0_W6BEG;
 output [15:0] Tile_X0Y0_WW4BEG;
 input [3:0] Tile_X0Y1_E1END;
 input [7:0] Tile_X0Y1_E2END;
 input [7:0] Tile_X0Y1_E2MID;
 input [11:0] Tile_X0Y1_E6END;
 input [15:0] Tile_X0Y1_EE4END;
 input [31:0] Tile_X0Y1_FrameData;
 output [31:0] Tile_X0Y1_FrameData_O;
 input [19:0] Tile_X0Y1_FrameStrobe;
 input [3:0] Tile_X0Y1_N1END;
 input [7:0] Tile_X0Y1_N2END;
 input [7:0] Tile_X0Y1_N2MID;
 input [15:0] Tile_X0Y1_N4END;
 output [3:0] Tile_X0Y1_S1BEG;
 output [7:0] Tile_X0Y1_S2BEG;
 output [7:0] Tile_X0Y1_S2BEGb;
 output [15:0] Tile_X0Y1_S4BEG;
 output [3:0] Tile_X0Y1_W1BEG;
 output [7:0] Tile_X0Y1_W2BEG;
 output [7:0] Tile_X0Y1_W2BEGb;
 output [11:0] Tile_X0Y1_W6BEG;
 output [15:0] Tile_X0Y1_WW4BEG;

 wire net248;
 wire net249;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire \Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame0_bit0.Q ;
 wire \Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame0_bit1.Q ;
 wire \Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame0_bit10.Q ;
 wire \Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame0_bit11.Q ;
 wire \Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame0_bit12.Q ;
 wire \Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame0_bit13.Q ;
 wire \Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame0_bit14.Q ;
 wire \Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame0_bit15.Q ;
 wire \Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame0_bit16.Q ;
 wire \Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame0_bit17.Q ;
 wire \Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame0_bit18.Q ;
 wire \Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame0_bit19.Q ;
 wire \Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame0_bit2.Q ;
 wire \Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame0_bit20.Q ;
 wire \Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame0_bit21.Q ;
 wire \Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame0_bit22.Q ;
 wire \Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame0_bit23.Q ;
 wire \Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame0_bit24.Q ;
 wire \Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame0_bit25.Q ;
 wire \Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame0_bit26.Q ;
 wire \Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame0_bit27.Q ;
 wire \Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame0_bit28.Q ;
 wire \Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame0_bit29.Q ;
 wire \Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame0_bit3.Q ;
 wire \Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame0_bit30.Q ;
 wire \Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame0_bit31.Q ;
 wire \Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame0_bit4.Q ;
 wire \Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame0_bit5.Q ;
 wire \Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame0_bit6.Q ;
 wire \Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame0_bit7.Q ;
 wire \Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame0_bit8.Q ;
 wire \Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame0_bit9.Q ;
 wire \Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame1_bit0.Q ;
 wire \Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame1_bit1.Q ;
 wire \Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame1_bit10.Q ;
 wire \Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame1_bit11.Q ;
 wire \Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame1_bit12.Q ;
 wire \Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame1_bit13.Q ;
 wire \Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame1_bit14.Q ;
 wire \Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame1_bit15.Q ;
 wire \Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame1_bit16.Q ;
 wire \Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame1_bit17.Q ;
 wire \Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame1_bit18.Q ;
 wire \Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame1_bit19.Q ;
 wire \Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame1_bit2.Q ;
 wire \Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame1_bit20.Q ;
 wire \Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame1_bit21.Q ;
 wire \Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame1_bit22.Q ;
 wire \Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame1_bit23.Q ;
 wire \Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame1_bit24.Q ;
 wire \Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame1_bit25.Q ;
 wire \Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame1_bit26.Q ;
 wire \Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame1_bit27.Q ;
 wire \Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame1_bit28.Q ;
 wire \Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame1_bit29.Q ;
 wire \Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame1_bit3.Q ;
 wire \Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame1_bit30.Q ;
 wire \Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame1_bit31.Q ;
 wire \Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame1_bit4.Q ;
 wire \Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame1_bit5.Q ;
 wire \Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame1_bit6.Q ;
 wire \Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame1_bit7.Q ;
 wire \Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame1_bit8.Q ;
 wire \Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame1_bit9.Q ;
 wire \Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame2_bit0.Q ;
 wire \Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame2_bit1.Q ;
 wire \Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame2_bit10.Q ;
 wire \Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame2_bit11.Q ;
 wire \Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame2_bit12.Q ;
 wire \Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame2_bit13.Q ;
 wire \Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame2_bit14.Q ;
 wire \Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame2_bit15.Q ;
 wire \Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame2_bit16.Q ;
 wire \Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame2_bit17.Q ;
 wire \Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame2_bit18.Q ;
 wire \Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame2_bit19.Q ;
 wire \Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame2_bit2.Q ;
 wire \Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame2_bit20.Q ;
 wire \Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame2_bit21.Q ;
 wire \Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame2_bit22.Q ;
 wire \Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame2_bit23.Q ;
 wire \Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame2_bit24.Q ;
 wire \Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame2_bit25.Q ;
 wire \Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame2_bit26.Q ;
 wire \Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame2_bit27.Q ;
 wire \Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame2_bit28.Q ;
 wire \Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame2_bit29.Q ;
 wire \Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame2_bit3.Q ;
 wire \Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame2_bit30.Q ;
 wire \Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame2_bit31.Q ;
 wire \Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame2_bit4.Q ;
 wire \Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame2_bit5.Q ;
 wire \Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame2_bit6.Q ;
 wire \Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame2_bit7.Q ;
 wire \Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame2_bit8.Q ;
 wire \Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame2_bit9.Q ;
 wire \Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame3_bit0.Q ;
 wire \Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame3_bit1.Q ;
 wire \Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame3_bit10.Q ;
 wire \Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame3_bit11.Q ;
 wire \Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame3_bit12.Q ;
 wire \Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame3_bit13.Q ;
 wire \Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame3_bit14.Q ;
 wire \Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame3_bit15.Q ;
 wire \Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame3_bit16.Q ;
 wire \Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame3_bit17.Q ;
 wire \Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame3_bit18.Q ;
 wire \Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame3_bit19.Q ;
 wire \Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame3_bit2.Q ;
 wire \Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame3_bit20.Q ;
 wire \Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame3_bit21.Q ;
 wire \Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame3_bit22.Q ;
 wire \Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame3_bit23.Q ;
 wire \Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame3_bit24.Q ;
 wire \Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame3_bit25.Q ;
 wire \Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame3_bit26.Q ;
 wire \Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame3_bit27.Q ;
 wire \Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame3_bit28.Q ;
 wire \Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame3_bit29.Q ;
 wire \Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame3_bit3.Q ;
 wire \Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame3_bit30.Q ;
 wire \Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame3_bit31.Q ;
 wire \Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame3_bit4.Q ;
 wire \Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame3_bit5.Q ;
 wire \Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame3_bit6.Q ;
 wire \Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame3_bit7.Q ;
 wire \Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame3_bit8.Q ;
 wire \Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame3_bit9.Q ;
 wire \Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame4_bit0.Q ;
 wire \Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame4_bit1.Q ;
 wire \Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame4_bit10.Q ;
 wire \Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame4_bit11.Q ;
 wire \Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame4_bit12.Q ;
 wire \Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame4_bit13.Q ;
 wire \Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame4_bit14.Q ;
 wire \Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame4_bit15.Q ;
 wire \Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame4_bit16.Q ;
 wire \Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame4_bit17.Q ;
 wire \Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame4_bit18.Q ;
 wire \Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame4_bit19.Q ;
 wire \Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame4_bit2.Q ;
 wire \Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame4_bit20.Q ;
 wire \Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame4_bit21.Q ;
 wire \Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame4_bit22.Q ;
 wire \Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame4_bit23.Q ;
 wire \Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame4_bit24.Q ;
 wire \Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame4_bit25.Q ;
 wire \Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame4_bit26.Q ;
 wire \Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame4_bit27.Q ;
 wire \Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame4_bit28.Q ;
 wire \Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame4_bit29.Q ;
 wire \Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame4_bit3.Q ;
 wire \Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame4_bit30.Q ;
 wire \Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame4_bit31.Q ;
 wire \Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame4_bit4.Q ;
 wire \Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame4_bit5.Q ;
 wire \Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame4_bit6.Q ;
 wire \Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame4_bit7.Q ;
 wire \Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame4_bit8.Q ;
 wire \Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame4_bit9.Q ;
 wire \Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame5_bit0.Q ;
 wire \Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame5_bit1.Q ;
 wire \Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame5_bit10.Q ;
 wire \Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame5_bit11.Q ;
 wire \Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame5_bit12.Q ;
 wire \Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame5_bit13.Q ;
 wire \Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame5_bit14.Q ;
 wire \Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame5_bit15.Q ;
 wire \Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame5_bit16.Q ;
 wire \Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame5_bit17.Q ;
 wire \Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame5_bit18.Q ;
 wire \Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame5_bit19.Q ;
 wire \Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame5_bit2.Q ;
 wire \Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame5_bit20.Q ;
 wire \Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame5_bit21.Q ;
 wire \Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame5_bit22.Q ;
 wire \Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame5_bit23.Q ;
 wire \Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame5_bit24.Q ;
 wire \Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame5_bit25.Q ;
 wire \Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame5_bit26.Q ;
 wire \Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame5_bit27.Q ;
 wire \Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame5_bit28.Q ;
 wire \Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame5_bit29.Q ;
 wire \Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame5_bit3.Q ;
 wire \Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame5_bit30.Q ;
 wire \Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame5_bit31.Q ;
 wire \Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame5_bit4.Q ;
 wire \Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame5_bit5.Q ;
 wire \Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame5_bit6.Q ;
 wire \Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame5_bit7.Q ;
 wire \Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame5_bit8.Q ;
 wire \Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame5_bit9.Q ;
 wire \Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame6_bit0.Q ;
 wire \Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame6_bit1.Q ;
 wire \Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame6_bit10.Q ;
 wire \Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame6_bit11.Q ;
 wire \Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame6_bit12.Q ;
 wire \Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame6_bit13.Q ;
 wire \Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame6_bit14.Q ;
 wire \Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame6_bit15.Q ;
 wire \Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame6_bit16.Q ;
 wire \Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame6_bit17.Q ;
 wire \Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame6_bit18.Q ;
 wire \Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame6_bit19.Q ;
 wire \Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame6_bit2.Q ;
 wire \Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame6_bit20.Q ;
 wire \Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame6_bit21.Q ;
 wire \Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame6_bit22.Q ;
 wire \Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame6_bit23.Q ;
 wire \Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame6_bit24.Q ;
 wire \Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame6_bit25.Q ;
 wire \Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame6_bit26.Q ;
 wire \Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame6_bit27.Q ;
 wire \Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame6_bit28.Q ;
 wire \Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame6_bit29.Q ;
 wire \Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame6_bit3.Q ;
 wire \Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame6_bit30.Q ;
 wire \Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame6_bit31.Q ;
 wire \Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame6_bit4.Q ;
 wire \Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame6_bit5.Q ;
 wire \Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame6_bit6.Q ;
 wire \Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame6_bit7.Q ;
 wire \Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame6_bit8.Q ;
 wire \Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame6_bit9.Q ;
 wire \Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame7_bit0.Q ;
 wire \Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame7_bit1.Q ;
 wire \Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame7_bit10.Q ;
 wire \Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame7_bit11.Q ;
 wire \Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame7_bit12.Q ;
 wire \Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame7_bit13.Q ;
 wire \Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame7_bit14.Q ;
 wire \Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame7_bit15.Q ;
 wire \Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame7_bit16.Q ;
 wire \Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame7_bit17.Q ;
 wire \Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame7_bit18.Q ;
 wire \Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame7_bit19.Q ;
 wire \Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame7_bit2.Q ;
 wire \Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame7_bit20.Q ;
 wire \Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame7_bit21.Q ;
 wire \Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame7_bit22.Q ;
 wire \Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame7_bit23.Q ;
 wire \Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame7_bit24.Q ;
 wire \Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame7_bit25.Q ;
 wire \Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame7_bit26.Q ;
 wire \Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame7_bit27.Q ;
 wire \Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame7_bit28.Q ;
 wire \Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame7_bit29.Q ;
 wire \Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame7_bit3.Q ;
 wire \Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame7_bit30.Q ;
 wire \Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame7_bit31.Q ;
 wire \Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame7_bit4.Q ;
 wire \Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame7_bit5.Q ;
 wire \Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame7_bit6.Q ;
 wire \Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame7_bit7.Q ;
 wire \Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame7_bit8.Q ;
 wire \Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame7_bit9.Q ;
 wire \Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame8_bit0.Q ;
 wire \Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame8_bit1.Q ;
 wire \Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame8_bit10.Q ;
 wire \Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame8_bit11.Q ;
 wire \Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame8_bit12.Q ;
 wire \Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame8_bit13.Q ;
 wire \Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame8_bit14.Q ;
 wire \Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame8_bit15.Q ;
 wire \Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame8_bit16.Q ;
 wire \Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame8_bit17.Q ;
 wire \Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame8_bit18.Q ;
 wire \Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame8_bit19.Q ;
 wire \Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame8_bit2.Q ;
 wire \Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame8_bit20.Q ;
 wire \Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame8_bit21.Q ;
 wire \Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame8_bit22.Q ;
 wire \Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame8_bit23.Q ;
 wire \Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame8_bit24.Q ;
 wire \Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame8_bit25.Q ;
 wire \Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame8_bit26.Q ;
 wire \Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame8_bit27.Q ;
 wire \Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame8_bit28.Q ;
 wire \Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame8_bit29.Q ;
 wire \Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame8_bit3.Q ;
 wire \Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame8_bit30.Q ;
 wire \Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame8_bit31.Q ;
 wire \Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame8_bit4.Q ;
 wire \Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame8_bit5.Q ;
 wire \Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame8_bit6.Q ;
 wire \Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame8_bit7.Q ;
 wire \Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame8_bit8.Q ;
 wire \Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame8_bit9.Q ;
 wire \Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame9_bit22.Q ;
 wire \Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame9_bit23.Q ;
 wire \Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame9_bit24.Q ;
 wire \Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame9_bit25.Q ;
 wire \Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame9_bit26.Q ;
 wire \Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame9_bit27.Q ;
 wire \Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame9_bit28.Q ;
 wire \Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame9_bit29.Q ;
 wire \Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame9_bit30.Q ;
 wire \Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame9_bit31.Q ;
 wire \Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.J_NS2_BEG0 ;
 wire \Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.J_NS2_BEG1 ;
 wire \Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.J_NS2_BEG2 ;
 wire \Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.J_NS2_BEG3 ;
 wire \Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.J_NS2_BEG4 ;
 wire \Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.J_NS2_BEG5 ;
 wire \Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.J_NS2_BEG6 ;
 wire \Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.J_NS2_BEG7 ;
 wire \Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.J_NS4_BEG0 ;
 wire \Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.J_NS4_BEG1 ;
 wire \Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.J_NS4_BEG10 ;
 wire \Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.J_NS4_BEG11 ;
 wire \Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.J_NS4_BEG12 ;
 wire \Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.J_NS4_BEG13 ;
 wire \Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.J_NS4_BEG14 ;
 wire \Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.J_NS4_BEG15 ;
 wire \Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.J_NS4_BEG2 ;
 wire \Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.J_NS4_BEG3 ;
 wire \Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.J_NS4_BEG4 ;
 wire \Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.J_NS4_BEG5 ;
 wire \Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.J_NS4_BEG6 ;
 wire \Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.J_NS4_BEG7 ;
 wire \Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.J_NS4_BEG8 ;
 wire \Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.J_NS4_BEG9 ;
 wire \Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.N1BEG0 ;
 wire \Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.N1BEG1 ;
 wire \Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.N1BEG2 ;
 wire \Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.N1BEG3 ;
 wire \Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.N1END0 ;
 wire \Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.N1END1 ;
 wire \Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.N1END2 ;
 wire \Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.N1END3 ;
 wire \Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.N2BEG0 ;
 wire \Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.N2BEG1 ;
 wire \Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.N2BEG2 ;
 wire \Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.N2BEG3 ;
 wire \Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.N2BEG4 ;
 wire \Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.N2BEG5 ;
 wire \Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.N2BEG6 ;
 wire \Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.N2BEG7 ;
 wire \Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.N2BEGb0 ;
 wire \Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.N2BEGb1 ;
 wire \Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.N2BEGb2 ;
 wire \Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.N2BEGb3 ;
 wire \Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.N2BEGb4 ;
 wire \Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.N2BEGb5 ;
 wire \Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.N2BEGb6 ;
 wire \Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.N2BEGb7 ;
 wire \Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.N4BEG0 ;
 wire \Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.N4BEG1 ;
 wire \Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.N4BEG2 ;
 wire \Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.N4BEG3 ;
 wire \Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.S2BEG0 ;
 wire \Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.S2BEG1 ;
 wire \Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.S2BEG2 ;
 wire \Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.S2BEG3 ;
 wire \Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.S2BEG4 ;
 wire \Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.S2BEG5 ;
 wire \Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.S2BEG6 ;
 wire \Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.S2BEG7 ;
 wire \Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.S4BEG0 ;
 wire \Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.S4BEG1 ;
 wire \Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.S4BEG2 ;
 wire \Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.S4BEG3 ;
 wire \Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.W1BEG0 ;
 wire \Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.W1BEG1 ;
 wire \Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.W1BEG2 ;
 wire \Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.W1BEG3 ;
 wire \Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.W2BEG0 ;
 wire \Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.W2BEG1 ;
 wire \Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.W2BEG2 ;
 wire \Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.W2BEG3 ;
 wire \Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.W2BEG4 ;
 wire \Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.W2BEG5 ;
 wire \Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.W2BEG6 ;
 wire \Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.W2BEG7 ;
 wire \Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.W2BEGb0 ;
 wire \Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.W2BEGb1 ;
 wire \Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.W2BEGb2 ;
 wire \Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.W2BEGb3 ;
 wire \Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.W2BEGb4 ;
 wire \Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.W2BEGb5 ;
 wire \Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.W2BEGb6 ;
 wire \Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.W2BEGb7 ;
 wire \Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.W6BEG0 ;
 wire \Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.W6BEG1 ;
 wire \Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.W6BEG10 ;
 wire \Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.W6BEG11 ;
 wire \Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.W6BEG2 ;
 wire \Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.W6BEG3 ;
 wire \Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.W6BEG4 ;
 wire \Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.W6BEG5 ;
 wire \Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.W6BEG6 ;
 wire \Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.W6BEG7 ;
 wire \Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.W6BEG8 ;
 wire \Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.W6BEG9 ;
 wire \Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.WW4BEG0 ;
 wire \Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.WW4BEG1 ;
 wire \Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.WW4BEG10 ;
 wire \Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.WW4BEG11 ;
 wire \Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.WW4BEG12 ;
 wire \Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.WW4BEG13 ;
 wire \Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.WW4BEG14 ;
 wire \Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.WW4BEG15 ;
 wire \Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.WW4BEG2 ;
 wire \Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.WW4BEG3 ;
 wire \Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.WW4BEG4 ;
 wire \Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.WW4BEG5 ;
 wire \Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.WW4BEG6 ;
 wire \Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.WW4BEG7 ;
 wire \Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.WW4BEG8 ;
 wire \Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.WW4BEG9 ;
 wire \Tile_X0Y0_EF_SRAM_top.N4BEG_outbuf_10.A ;
 wire \Tile_X0Y0_EF_SRAM_top.N4BEG_outbuf_11.A ;
 wire \Tile_X0Y0_EF_SRAM_top.N4BEG_outbuf_8.A ;
 wire \Tile_X0Y0_EF_SRAM_top.N4BEG_outbuf_9.A ;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net477;
 wire net478;
 wire net479;
 wire net480;
 wire net481;
 wire net482;
 wire net483;
 wire net484;
 wire net485;
 wire net486;
 wire net487;
 wire net488;
 wire net489;
 wire net490;
 wire net491;
 wire net492;
 wire net493;
 wire net494;
 wire net495;
 wire net496;
 wire net497;
 wire net498;
 wire net499;
 wire net500;
 wire net501;
 wire net502;
 wire net503;
 wire net504;
 wire net505;
 wire net506;
 wire net507;
 wire net508;
 wire net509;
 wire net510;
 wire net511;
 wire net512;
 wire net513;
 wire net514;
 wire net515;
 wire net516;
 wire net517;
 wire net518;
 wire net519;
 wire net520;
 wire net521;
 wire net522;
 wire net523;
 wire net524;
 wire net525;
 wire net526;
 wire net527;
 wire net528;
 wire net529;
 wire net530;
 wire net531;
 wire net532;
 wire net533;
 wire net534;
 wire net535;
 wire net536;
 wire net537;
 wire net538;
 wire net539;
 wire net540;
 wire net541;
 wire net542;
 wire net543;
 wire net544;
 wire net545;
 wire net546;
 wire net547;
 wire net548;
 wire net549;
 wire net550;
 wire net551;
 wire net552;
 wire net553;
 wire net554;
 wire net555;
 wire net556;
 wire net557;
 wire net558;
 wire net559;
 wire net560;
 wire net561;
 wire net562;
 wire net563;
 wire net564;
 wire net565;
 wire net566;
 wire net567;
 wire net568;
 wire net569;
 wire net570;
 wire net571;
 wire net572;
 wire net573;
 wire net574;
 wire net575;
 wire net576;
 wire net577;
 wire net578;
 wire \Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame0_bit0.Q ;
 wire \Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame0_bit1.Q ;
 wire \Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame0_bit10.Q ;
 wire \Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame0_bit11.Q ;
 wire \Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame0_bit12.Q ;
 wire \Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame0_bit13.Q ;
 wire \Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame0_bit14.Q ;
 wire \Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame0_bit15.Q ;
 wire \Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame0_bit16.Q ;
 wire \Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame0_bit17.Q ;
 wire \Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame0_bit18.Q ;
 wire \Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame0_bit19.Q ;
 wire \Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame0_bit2.Q ;
 wire \Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame0_bit20.Q ;
 wire \Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame0_bit21.Q ;
 wire \Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame0_bit22.Q ;
 wire \Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame0_bit23.Q ;
 wire \Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame0_bit24.Q ;
 wire \Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame0_bit25.Q ;
 wire \Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame0_bit26.Q ;
 wire \Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame0_bit27.Q ;
 wire \Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame0_bit28.Q ;
 wire \Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame0_bit29.Q ;
 wire \Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame0_bit3.Q ;
 wire \Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame0_bit30.Q ;
 wire \Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame0_bit31.Q ;
 wire \Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame0_bit4.Q ;
 wire \Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame0_bit5.Q ;
 wire \Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame0_bit6.Q ;
 wire \Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame0_bit7.Q ;
 wire \Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame0_bit8.Q ;
 wire \Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame0_bit9.Q ;
 wire \Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame1_bit0.Q ;
 wire \Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame1_bit1.Q ;
 wire \Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame1_bit10.Q ;
 wire \Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame1_bit11.Q ;
 wire \Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame1_bit12.Q ;
 wire \Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame1_bit13.Q ;
 wire \Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame1_bit14.Q ;
 wire \Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame1_bit15.Q ;
 wire \Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame1_bit16.Q ;
 wire \Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame1_bit17.Q ;
 wire \Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame1_bit18.Q ;
 wire \Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame1_bit19.Q ;
 wire \Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame1_bit2.Q ;
 wire \Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame1_bit20.Q ;
 wire \Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame1_bit21.Q ;
 wire \Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame1_bit22.Q ;
 wire \Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame1_bit23.Q ;
 wire \Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame1_bit24.Q ;
 wire \Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame1_bit25.Q ;
 wire \Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame1_bit26.Q ;
 wire \Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame1_bit27.Q ;
 wire \Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame1_bit28.Q ;
 wire \Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame1_bit29.Q ;
 wire \Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame1_bit3.Q ;
 wire \Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame1_bit30.Q ;
 wire \Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame1_bit31.Q ;
 wire \Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame1_bit4.Q ;
 wire \Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame1_bit5.Q ;
 wire \Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame1_bit6.Q ;
 wire \Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame1_bit7.Q ;
 wire \Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame1_bit8.Q ;
 wire \Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame1_bit9.Q ;
 wire \Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame2_bit0.Q ;
 wire \Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame2_bit1.Q ;
 wire \Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame2_bit10.Q ;
 wire \Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame2_bit11.Q ;
 wire \Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame2_bit12.Q ;
 wire \Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame2_bit13.Q ;
 wire \Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame2_bit14.Q ;
 wire \Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame2_bit15.Q ;
 wire \Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame2_bit16.Q ;
 wire \Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame2_bit17.Q ;
 wire \Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame2_bit18.Q ;
 wire \Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame2_bit19.Q ;
 wire \Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame2_bit2.Q ;
 wire \Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame2_bit20.Q ;
 wire \Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame2_bit21.Q ;
 wire \Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame2_bit22.Q ;
 wire \Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame2_bit23.Q ;
 wire \Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame2_bit24.Q ;
 wire \Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame2_bit25.Q ;
 wire \Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame2_bit26.Q ;
 wire \Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame2_bit27.Q ;
 wire \Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame2_bit28.Q ;
 wire \Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame2_bit29.Q ;
 wire \Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame2_bit3.Q ;
 wire \Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame2_bit30.Q ;
 wire \Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame2_bit31.Q ;
 wire \Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame2_bit4.Q ;
 wire \Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame2_bit5.Q ;
 wire \Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame2_bit6.Q ;
 wire \Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame2_bit7.Q ;
 wire \Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame2_bit8.Q ;
 wire \Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame2_bit9.Q ;
 wire \Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame3_bit0.Q ;
 wire \Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame3_bit1.Q ;
 wire \Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame3_bit10.Q ;
 wire \Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame3_bit11.Q ;
 wire \Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame3_bit12.Q ;
 wire \Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame3_bit13.Q ;
 wire \Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame3_bit14.Q ;
 wire \Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame3_bit15.Q ;
 wire \Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame3_bit16.Q ;
 wire \Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame3_bit17.Q ;
 wire \Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame3_bit18.Q ;
 wire \Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame3_bit19.Q ;
 wire \Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame3_bit2.Q ;
 wire \Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame3_bit20.Q ;
 wire \Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame3_bit21.Q ;
 wire \Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame3_bit22.Q ;
 wire \Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame3_bit23.Q ;
 wire \Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame3_bit24.Q ;
 wire \Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame3_bit25.Q ;
 wire \Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame3_bit26.Q ;
 wire \Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame3_bit27.Q ;
 wire \Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame3_bit28.Q ;
 wire \Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame3_bit29.Q ;
 wire \Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame3_bit3.Q ;
 wire \Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame3_bit30.Q ;
 wire \Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame3_bit31.Q ;
 wire \Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame3_bit4.Q ;
 wire \Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame3_bit5.Q ;
 wire \Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame3_bit6.Q ;
 wire \Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame3_bit7.Q ;
 wire \Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame3_bit8.Q ;
 wire \Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame3_bit9.Q ;
 wire \Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame4_bit0.Q ;
 wire \Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame4_bit1.Q ;
 wire \Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame4_bit10.Q ;
 wire \Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame4_bit11.Q ;
 wire \Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame4_bit12.Q ;
 wire \Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame4_bit13.Q ;
 wire \Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame4_bit14.Q ;
 wire \Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame4_bit15.Q ;
 wire \Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame4_bit16.Q ;
 wire \Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame4_bit17.Q ;
 wire \Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame4_bit18.Q ;
 wire \Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame4_bit19.Q ;
 wire \Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame4_bit2.Q ;
 wire \Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame4_bit20.Q ;
 wire \Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame4_bit21.Q ;
 wire \Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame4_bit22.Q ;
 wire \Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame4_bit23.Q ;
 wire \Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame4_bit24.Q ;
 wire \Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame4_bit25.Q ;
 wire \Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame4_bit26.Q ;
 wire \Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame4_bit27.Q ;
 wire \Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame4_bit28.Q ;
 wire \Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame4_bit29.Q ;
 wire \Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame4_bit3.Q ;
 wire \Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame4_bit30.Q ;
 wire \Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame4_bit31.Q ;
 wire \Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame4_bit4.Q ;
 wire \Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame4_bit5.Q ;
 wire \Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame4_bit6.Q ;
 wire \Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame4_bit7.Q ;
 wire \Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame4_bit8.Q ;
 wire \Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame4_bit9.Q ;
 wire \Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame5_bit0.Q ;
 wire \Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame5_bit1.Q ;
 wire \Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame5_bit10.Q ;
 wire \Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame5_bit11.Q ;
 wire \Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame5_bit12.Q ;
 wire \Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame5_bit13.Q ;
 wire \Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame5_bit14.Q ;
 wire \Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame5_bit15.Q ;
 wire \Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame5_bit16.Q ;
 wire \Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame5_bit17.Q ;
 wire \Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame5_bit18.Q ;
 wire \Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame5_bit19.Q ;
 wire \Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame5_bit2.Q ;
 wire \Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame5_bit20.Q ;
 wire \Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame5_bit21.Q ;
 wire \Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame5_bit22.Q ;
 wire \Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame5_bit23.Q ;
 wire \Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame5_bit24.Q ;
 wire \Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame5_bit25.Q ;
 wire \Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame5_bit26.Q ;
 wire \Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame5_bit27.Q ;
 wire \Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame5_bit28.Q ;
 wire \Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame5_bit29.Q ;
 wire \Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame5_bit3.Q ;
 wire \Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame5_bit30.Q ;
 wire \Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame5_bit31.Q ;
 wire \Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame5_bit4.Q ;
 wire \Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame5_bit5.Q ;
 wire \Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame5_bit6.Q ;
 wire \Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame5_bit7.Q ;
 wire \Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame5_bit8.Q ;
 wire \Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame5_bit9.Q ;
 wire \Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame6_bit0.Q ;
 wire \Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame6_bit1.Q ;
 wire \Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame6_bit10.Q ;
 wire \Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame6_bit11.Q ;
 wire \Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame6_bit12.Q ;
 wire \Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame6_bit13.Q ;
 wire \Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame6_bit14.Q ;
 wire \Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame6_bit15.Q ;
 wire \Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame6_bit16.Q ;
 wire \Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame6_bit17.Q ;
 wire \Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame6_bit18.Q ;
 wire \Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame6_bit19.Q ;
 wire \Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame6_bit2.Q ;
 wire \Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame6_bit20.Q ;
 wire \Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame6_bit21.Q ;
 wire \Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame6_bit22.Q ;
 wire \Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame6_bit23.Q ;
 wire \Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame6_bit24.Q ;
 wire \Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame6_bit25.Q ;
 wire \Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame6_bit26.Q ;
 wire \Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame6_bit27.Q ;
 wire \Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame6_bit28.Q ;
 wire \Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame6_bit29.Q ;
 wire \Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame6_bit3.Q ;
 wire \Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame6_bit30.Q ;
 wire \Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame6_bit31.Q ;
 wire \Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame6_bit4.Q ;
 wire \Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame6_bit5.Q ;
 wire \Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame6_bit6.Q ;
 wire \Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame6_bit7.Q ;
 wire \Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame6_bit8.Q ;
 wire \Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame6_bit9.Q ;
 wire \Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame7_bit0.Q ;
 wire \Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame7_bit1.Q ;
 wire \Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame7_bit10.Q ;
 wire \Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame7_bit11.Q ;
 wire \Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame7_bit12.Q ;
 wire \Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame7_bit13.Q ;
 wire \Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame7_bit14.Q ;
 wire \Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame7_bit15.Q ;
 wire \Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame7_bit16.Q ;
 wire \Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame7_bit17.Q ;
 wire \Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame7_bit18.Q ;
 wire \Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame7_bit19.Q ;
 wire \Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame7_bit2.Q ;
 wire \Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame7_bit20.Q ;
 wire \Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame7_bit21.Q ;
 wire \Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame7_bit22.Q ;
 wire \Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame7_bit23.Q ;
 wire \Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame7_bit24.Q ;
 wire \Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame7_bit25.Q ;
 wire \Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame7_bit26.Q ;
 wire \Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame7_bit27.Q ;
 wire \Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame7_bit28.Q ;
 wire \Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame7_bit29.Q ;
 wire \Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame7_bit3.Q ;
 wire \Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame7_bit30.Q ;
 wire \Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame7_bit31.Q ;
 wire \Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame7_bit4.Q ;
 wire \Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame7_bit5.Q ;
 wire \Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame7_bit6.Q ;
 wire \Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame7_bit7.Q ;
 wire \Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame7_bit8.Q ;
 wire \Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame7_bit9.Q ;
 wire \Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame8_bit0.Q ;
 wire \Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame8_bit1.Q ;
 wire \Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame8_bit10.Q ;
 wire \Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame8_bit11.Q ;
 wire \Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame8_bit12.Q ;
 wire \Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame8_bit13.Q ;
 wire \Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame8_bit14.Q ;
 wire \Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame8_bit15.Q ;
 wire \Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame8_bit16.Q ;
 wire \Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame8_bit17.Q ;
 wire \Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame8_bit18.Q ;
 wire \Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame8_bit19.Q ;
 wire \Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame8_bit2.Q ;
 wire \Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame8_bit20.Q ;
 wire \Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame8_bit21.Q ;
 wire \Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame8_bit22.Q ;
 wire \Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame8_bit23.Q ;
 wire \Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame8_bit24.Q ;
 wire \Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame8_bit25.Q ;
 wire \Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame8_bit26.Q ;
 wire \Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame8_bit27.Q ;
 wire \Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame8_bit28.Q ;
 wire \Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame8_bit29.Q ;
 wire \Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame8_bit3.Q ;
 wire \Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame8_bit30.Q ;
 wire \Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame8_bit31.Q ;
 wire \Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame8_bit4.Q ;
 wire \Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame8_bit5.Q ;
 wire \Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame8_bit6.Q ;
 wire \Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame8_bit7.Q ;
 wire \Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame8_bit8.Q ;
 wire \Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame8_bit9.Q ;
 wire \Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame9_bit14.Q ;
 wire \Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame9_bit15.Q ;
 wire \Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame9_bit16.Q ;
 wire \Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame9_bit17.Q ;
 wire \Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame9_bit18.Q ;
 wire \Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame9_bit19.Q ;
 wire \Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame9_bit20.Q ;
 wire \Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame9_bit21.Q ;
 wire \Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame9_bit22.Q ;
 wire \Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame9_bit23.Q ;
 wire \Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame9_bit24.Q ;
 wire \Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame9_bit25.Q ;
 wire \Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame9_bit26.Q ;
 wire \Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame9_bit27.Q ;
 wire \Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame9_bit28.Q ;
 wire \Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame9_bit29.Q ;
 wire \Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame9_bit30.Q ;
 wire \Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame9_bit31.Q ;
 wire \Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.J_NS4_BEG10 ;
 wire \Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.J_NS4_BEG11 ;
 wire \Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.J_NS4_BEG12 ;
 wire \Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.J_NS4_BEG13 ;
 wire \Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.J_NS4_BEG14 ;
 wire \Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.J_NS4_BEG15 ;
 wire \Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.J_NS4_BEG4 ;
 wire \Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.J_NS4_BEG5 ;
 wire \Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.J_NS4_BEG6 ;
 wire \Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.J_NS4_BEG7 ;
 wire \Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.J_NS4_BEG8 ;
 wire \Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.J_NS4_BEG9 ;
 wire \Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.S1BEG0 ;
 wire \Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.S1BEG1 ;
 wire \Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.S1BEG2 ;
 wire \Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.S1BEG3 ;
 wire \Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.S2BEG0 ;
 wire \Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.S2BEG1 ;
 wire \Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.S2BEG2 ;
 wire \Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.S2BEG3 ;
 wire \Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.S2BEG4 ;
 wire \Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.S2BEG5 ;
 wire \Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.S2BEG6 ;
 wire \Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.S2BEG7 ;
 wire \Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.S4BEG0 ;
 wire \Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.S4BEG1 ;
 wire \Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.S4BEG2 ;
 wire \Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.S4BEG3 ;
 wire \Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.W1BEG0 ;
 wire \Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.W1BEG1 ;
 wire \Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.W1BEG2 ;
 wire \Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.W1BEG3 ;
 wire \Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.W2BEG0 ;
 wire \Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.W2BEG1 ;
 wire \Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.W2BEG2 ;
 wire \Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.W2BEG3 ;
 wire \Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.W2BEG4 ;
 wire \Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.W2BEG5 ;
 wire \Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.W2BEG6 ;
 wire \Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.W2BEG7 ;
 wire \Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.W2BEGb0 ;
 wire \Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.W2BEGb1 ;
 wire \Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.W2BEGb2 ;
 wire \Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.W2BEGb3 ;
 wire \Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.W2BEGb4 ;
 wire \Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.W2BEGb5 ;
 wire \Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.W2BEGb6 ;
 wire \Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.W2BEGb7 ;
 wire \Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.W6BEG0 ;
 wire \Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.W6BEG1 ;
 wire \Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.W6BEG10 ;
 wire \Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.W6BEG11 ;
 wire \Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.W6BEG2 ;
 wire \Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.W6BEG3 ;
 wire \Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.W6BEG4 ;
 wire \Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.W6BEG5 ;
 wire \Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.W6BEG6 ;
 wire \Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.W6BEG7 ;
 wire \Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.W6BEG8 ;
 wire \Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.W6BEG9 ;
 wire \Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.WW4BEG0 ;
 wire \Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.WW4BEG1 ;
 wire \Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.WW4BEG10 ;
 wire \Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.WW4BEG11 ;
 wire \Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.WW4BEG12 ;
 wire \Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.WW4BEG13 ;
 wire \Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.WW4BEG14 ;
 wire \Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.WW4BEG15 ;
 wire \Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.WW4BEG2 ;
 wire \Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.WW4BEG3 ;
 wire \Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.WW4BEG4 ;
 wire \Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.WW4BEG5 ;
 wire \Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.WW4BEG6 ;
 wire \Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.WW4BEG7 ;
 wire \Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.WW4BEG8 ;
 wire \Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.WW4BEG9 ;
 wire net579;
 wire net580;
 wire net581;
 wire net582;
 wire net583;
 wire net584;
 wire net585;
 wire net586;
 wire net587;
 wire net588;
 wire net589;
 wire net590;
 wire net591;
 wire net592;
 wire net593;
 wire net594;
 wire net595;
 wire net596;
 wire net597;
 wire net598;
 wire net599;
 wire net600;
 wire net601;
 wire net602;
 wire net603;
 wire net604;
 wire net605;
 wire net606;
 wire net607;
 wire net608;
 wire net609;
 wire net610;
 wire net611;
 wire net612;
 wire net613;
 wire net614;
 wire net615;
 wire net616;
 wire net617;
 wire net618;
 wire net619;
 wire net620;
 wire net621;
 wire net622;
 wire net623;
 wire net624;
 wire net625;
 wire net626;
 wire net627;
 wire net628;
 wire net629;
 wire net630;
 wire net631;
 wire net632;
 wire net633;
 wire net634;
 wire net635;
 wire net636;
 wire net637;
 wire net638;
 wire net639;
 wire net640;
 wire net641;
 wire net642;
 wire net643;
 wire net644;
 wire net645;
 wire net646;
 wire net647;
 wire net648;
 wire net649;
 wire net650;
 wire net651;
 wire net652;
 wire net653;
 wire net654;
 wire net655;
 wire net656;
 wire net657;
 wire net658;
 wire net659;
 wire net660;
 wire net661;
 wire net662;
 wire net663;
 wire net664;
 wire net665;
 wire net666;
 wire net667;
 wire net668;
 wire net669;
 wire net670;
 wire net671;
 wire net672;
 wire net673;
 wire net674;
 wire net675;
 wire net676;
 wire net677;
 wire net678;
 wire net679;
 wire net680;
 wire net681;
 wire net682;
 wire net683;
 wire net684;
 wire net685;
 wire net686;
 wire net687;
 wire net688;
 wire net689;
 wire net690;
 wire net691;
 wire net692;
 wire net693;
 wire net694;
 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire net368;
 wire net369;
 wire net370;
 wire net371;
 wire net372;
 wire net373;
 wire net374;
 wire net375;
 wire net376;
 wire net377;
 wire net378;
 wire net379;
 wire net380;
 wire net381;
 wire net382;
 wire net383;
 wire net384;
 wire net385;
 wire net386;
 wire net387;
 wire net388;
 wire net389;
 wire net390;
 wire net391;
 wire net392;
 wire net393;
 wire net394;
 wire net395;
 wire net396;
 wire net397;
 wire net398;
 wire net399;
 wire net400;
 wire net401;
 wire net402;
 wire net403;
 wire net404;
 wire net405;
 wire net406;
 wire net407;
 wire net408;
 wire net409;
 wire net410;
 wire net411;
 wire net412;
 wire net413;
 wire net414;
 wire net415;
 wire net416;
 wire net417;
 wire net418;
 wire net419;
 wire net420;
 wire net421;
 wire net422;
 wire net423;
 wire net424;
 wire net425;
 wire net426;
 wire net427;
 wire net428;
 wire net429;
 wire net430;
 wire net431;
 wire net432;
 wire net433;
 wire net434;
 wire net435;
 wire net436;
 wire net437;
 wire net438;
 wire net439;
 wire net440;
 wire net441;
 wire net442;
 wire net443;
 wire net444;
 wire net445;
 wire net446;
 wire net447;
 wire net448;
 wire net449;
 wire net450;
 wire net451;
 wire net452;
 wire net453;
 wire net454;
 wire net455;
 wire net456;
 wire net457;
 wire net458;
 wire net459;
 wire net460;
 wire net461;
 wire net462;
 wire net463;
 wire net464;
 wire net465;
 wire net466;
 wire net467;
 wire net468;
 wire net469;
 wire net470;
 wire net471;
 wire net472;
 wire net473;
 wire net474;
 wire net475;
 wire net476;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire clknet_0_Tile_X0Y1_UserCLK;
 wire clknet_1_0__leaf_Tile_X0Y1_UserCLK;
 wire clknet_1_1__leaf_Tile_X0Y1_UserCLK;

 sky130_fd_sc_hd__inv_1 _0221_ (.A(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame0_bit27.Q ),
    .Y(_0000_));
 sky130_fd_sc_hd__inv_1 _0222_ (.A(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame0_bit29.Q ),
    .Y(_0001_));
 sky130_fd_sc_hd__inv_1 _0223_ (.A(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame0_bit31.Q ),
    .Y(_0002_));
 sky130_fd_sc_hd__inv_2 _0224_ (.A(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame2_bit30.Q ),
    .Y(_0003_));
 sky130_fd_sc_hd__inv_2 _0225_ (.A(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame1_bit0.Q ),
    .Y(_0004_));
 sky130_fd_sc_hd__inv_2 _0226_ (.A(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame1_bit2.Q ),
    .Y(_0005_));
 sky130_fd_sc_hd__inv_2 _0227_ (.A(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame1_bit4.Q ),
    .Y(_0006_));
 sky130_fd_sc_hd__inv_2 _0228_ (.A(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame1_bit7.Q ),
    .Y(_0007_));
 sky130_fd_sc_hd__inv_2 _0229_ (.A(net150),
    .Y(_0008_));
 sky130_fd_sc_hd__inv_1 _0230_ (.A(net127),
    .Y(_0009_));
 sky130_fd_sc_hd__inv_2 _0231_ (.A(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame8_bit16.Q ),
    .Y(_0010_));
 sky130_fd_sc_hd__inv_2 _0232_ (.A(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame8_bit19.Q ),
    .Y(_0011_));
 sky130_fd_sc_hd__inv_1 _0233_ (.A(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame8_bit22.Q ),
    .Y(_0012_));
 sky130_fd_sc_hd__inv_2 _0234_ (.A(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame8_bit25.Q ),
    .Y(_0013_));
 sky130_fd_sc_hd__inv_2 _0235_ (.A(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame7_bit20.Q ),
    .Y(_0014_));
 sky130_fd_sc_hd__inv_1 _0236_ (.A(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame7_bit23.Q ),
    .Y(_0015_));
 sky130_fd_sc_hd__inv_1 _0237_ (.A(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame7_bit26.Q ),
    .Y(_0016_));
 sky130_fd_sc_hd__inv_1 _0238_ (.A(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame7_bit29.Q ),
    .Y(_0017_));
 sky130_fd_sc_hd__inv_2 _0239_ (.A(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame0_bit24.Q ),
    .Y(_0018_));
 sky130_fd_sc_hd__inv_1 _0240_ (.A(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame0_bit25.Q ),
    .Y(_0019_));
 sky130_fd_sc_hd__inv_2 _0241_ (.A(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame0_bit26.Q ),
    .Y(_0020_));
 sky130_fd_sc_hd__inv_2 _0242_ (.A(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame0_bit28.Q ),
    .Y(_0021_));
 sky130_fd_sc_hd__inv_2 _0243_ (.A(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame0_bit30.Q ),
    .Y(_0022_));
 sky130_fd_sc_hd__inv_2 _0244_ (.A(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame4_bit22.Q ),
    .Y(_0023_));
 sky130_fd_sc_hd__inv_2 _0245_ (.A(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame4_bit24.Q ),
    .Y(_0024_));
 sky130_fd_sc_hd__inv_2 _0246_ (.A(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame4_bit26.Q ),
    .Y(_0025_));
 sky130_fd_sc_hd__inv_2 _0247_ (.A(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame4_bit28.Q ),
    .Y(_0026_));
 sky130_fd_sc_hd__inv_2 _0248_ (.A(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame4_bit30.Q ),
    .Y(_0027_));
 sky130_fd_sc_hd__inv_1 _0249_ (.A(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame8_bit6.Q ),
    .Y(_0028_));
 sky130_fd_sc_hd__inv_2 _0250_ (.A(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame8_bit7.Q ),
    .Y(_0029_));
 sky130_fd_sc_hd__inv_1 _0251_ (.A(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame8_bit8.Q ),
    .Y(_0030_));
 sky130_fd_sc_hd__inv_1 _0252_ (.A(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame8_bit9.Q ),
    .Y(_0031_));
 sky130_fd_sc_hd__inv_2 _0253_ (.A(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame8_bit10.Q ),
    .Y(_0032_));
 sky130_fd_sc_hd__inv_1 _0254_ (.A(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame8_bit11.Q ),
    .Y(_0033_));
 sky130_fd_sc_hd__inv_1 _0255_ (.A(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame8_bit12.Q ),
    .Y(_0034_));
 sky130_fd_sc_hd__inv_2 _0256_ (.A(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame8_bit13.Q ),
    .Y(_0035_));
 sky130_fd_sc_hd__inv_1 _0257_ (.A(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame8_bit14.Q ),
    .Y(_0036_));
 sky130_fd_sc_hd__inv_1 _0258_ (.A(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame8_bit15.Q ),
    .Y(_0037_));
 sky130_fd_sc_hd__inv_2 _0259_ (.A(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame8_bit16.Q ),
    .Y(_0038_));
 sky130_fd_sc_hd__inv_1 _0260_ (.A(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame8_bit17.Q ),
    .Y(_0039_));
 sky130_fd_sc_hd__inv_1 _0261_ (.A(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame7_bit10.Q ),
    .Y(_0040_));
 sky130_fd_sc_hd__inv_2 _0262_ (.A(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame7_bit11.Q ),
    .Y(_0041_));
 sky130_fd_sc_hd__inv_1 _0263_ (.A(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame7_bit12.Q ),
    .Y(_0042_));
 sky130_fd_sc_hd__inv_1 _0264_ (.A(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame7_bit13.Q ),
    .Y(_0043_));
 sky130_fd_sc_hd__inv_2 _0265_ (.A(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame7_bit14.Q ),
    .Y(_0044_));
 sky130_fd_sc_hd__inv_1 _0266_ (.A(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame7_bit15.Q ),
    .Y(_0045_));
 sky130_fd_sc_hd__inv_1 _0267_ (.A(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame7_bit16.Q ),
    .Y(_0046_));
 sky130_fd_sc_hd__inv_2 _0268_ (.A(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame7_bit17.Q ),
    .Y(_0047_));
 sky130_fd_sc_hd__inv_1 _0269_ (.A(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame7_bit18.Q ),
    .Y(_0048_));
 sky130_fd_sc_hd__inv_1 _0270_ (.A(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame7_bit19.Q ),
    .Y(_0049_));
 sky130_fd_sc_hd__inv_2 _0271_ (.A(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame7_bit20.Q ),
    .Y(_0050_));
 sky130_fd_sc_hd__inv_1 _0272_ (.A(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame7_bit21.Q ),
    .Y(_0051_));
 sky130_fd_sc_hd__inv_2 _0273_ (.A(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame1_bit1.Q ),
    .Y(_0052_));
 sky130_fd_sc_hd__inv_1 _0274_ (.A(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame1_bit4.Q ),
    .Y(_0053_));
 sky130_fd_sc_hd__inv_2 _0275_ (.A(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame1_bit5.Q ),
    .Y(_0054_));
 sky130_fd_sc_hd__mux2_1 _0276_ (.A0(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.N1END1 ),
    .A1(net56),
    .S(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame0_bit26.Q ),
    .X(_0055_));
 sky130_fd_sc_hd__nand2_1 _0277_ (.A(net114),
    .B(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame0_bit27.Q ),
    .Y(_0056_));
 sky130_fd_sc_hd__a2bb2o_1 _0278_ (.A1_N(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame0_bit26.Q ),
    .A2_N(_0056_),
    .B1(_0000_),
    .B2(_0055_),
    .X(_0057_));
 sky130_fd_sc_hd__mux4_2 _0279_ (.A0(net34),
    .A1(net64),
    .A2(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.J_NS4_BEG13 ),
    .A3(_0057_),
    .S0(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame8_bit28.Q ),
    .S1(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame8_bit29.Q ),
    .X(_0058_));
 sky130_fd_sc_hd__o21ba_1 _0280_ (.A1(net221),
    .A2(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame0_bit26.Q ),
    .B1_N(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame0_bit27.Q ),
    .X(_0059_));
 sky130_fd_sc_hd__o21a_1 _0281_ (.A1(net164),
    .A2(_0020_),
    .B1(_0059_),
    .X(_0060_));
 sky130_fd_sc_hd__a31o_1 _0282_ (.A1(_0020_),
    .A2(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame0_bit27.Q ),
    .A3(_0058_),
    .B1(_0060_),
    .X(_0061_));
 sky130_fd_sc_hd__mux4_2 _0283_ (.A0(net142),
    .A1(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.J_NS4_BEG13 ),
    .A2(net168),
    .A3(_0061_),
    .S0(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame9_bit17.Q ),
    .S1(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame9_bit16.Q ),
    .X(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.N1END1 ));
 sky130_fd_sc_hd__mux4_2 _0284_ (.A0(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.N1END1 ),
    .A1(net245),
    .A2(net114),
    .A3(net134),
    .S0(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame0_bit2.Q ),
    .S1(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame0_bit3.Q ),
    .X(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.J_NS4_BEG13 ));
 sky130_fd_sc_hd__mux4_1 _0285_ (.A0(net34),
    .A1(net60),
    .A2(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.J_NS4_BEG13 ),
    .A3(_0057_),
    .S0(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame9_bit24.Q ),
    .S1(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame9_bit25.Q ),
    .X(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.N1BEG1 ));
 sky130_fd_sc_hd__mux2_1 _0286_ (.A0(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.N1END2 ),
    .A1(net57),
    .S(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame0_bit28.Q ),
    .X(_0062_));
 sky130_fd_sc_hd__nand2_1 _0287_ (.A(net115),
    .B(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame0_bit29.Q ),
    .Y(_0063_));
 sky130_fd_sc_hd__a2bb2o_1 _0288_ (.A1_N(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame0_bit28.Q ),
    .A2_N(_0063_),
    .B1(_0001_),
    .B2(_0062_),
    .X(_0064_));
 sky130_fd_sc_hd__mux4_2 _0289_ (.A0(net35),
    .A1(net54),
    .A2(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.J_NS4_BEG14 ),
    .A3(_0064_),
    .S0(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame8_bit30.Q ),
    .S1(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame8_bit31.Q ),
    .X(_0065_));
 sky130_fd_sc_hd__o21ba_1 _0290_ (.A1(net222),
    .A2(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame0_bit28.Q ),
    .B1_N(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame0_bit29.Q ),
    .X(_0066_));
 sky130_fd_sc_hd__o21a_1 _0291_ (.A1(net165),
    .A2(_0021_),
    .B1(_0066_),
    .X(_0067_));
 sky130_fd_sc_hd__a31o_1 _0292_ (.A1(_0021_),
    .A2(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame0_bit29.Q ),
    .A3(_0065_),
    .B1(_0067_),
    .X(_0068_));
 sky130_fd_sc_hd__mux4_2 _0293_ (.A0(net143),
    .A1(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.J_NS4_BEG14 ),
    .A2(net169),
    .A3(_0068_),
    .S0(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame9_bit19.Q ),
    .S1(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame9_bit18.Q ),
    .X(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.N1END2 ));
 sky130_fd_sc_hd__mux4_2 _0294_ (.A0(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.N1END2 ),
    .A1(net246),
    .A2(net115),
    .A3(net135),
    .S0(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame0_bit4.Q ),
    .S1(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame0_bit5.Q ),
    .X(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.J_NS4_BEG14 ));
 sky130_fd_sc_hd__mux4_1 _0295_ (.A0(net35),
    .A1(net61),
    .A2(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.J_NS4_BEG14 ),
    .A3(_0064_),
    .S0(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame9_bit26.Q ),
    .S1(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame9_bit27.Q ),
    .X(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.N1BEG2 ));
 sky130_fd_sc_hd__mux2_1 _0296_ (.A0(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.N1END3 ),
    .A1(net58),
    .S(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame0_bit30.Q ),
    .X(_0069_));
 sky130_fd_sc_hd__nand2_1 _0297_ (.A(net116),
    .B(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame0_bit31.Q ),
    .Y(_0070_));
 sky130_fd_sc_hd__a2bb2o_1 _0298_ (.A1_N(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame0_bit30.Q ),
    .A2_N(_0070_),
    .B1(_0002_),
    .B2(_0069_),
    .X(_0071_));
 sky130_fd_sc_hd__mux4_2 _0299_ (.A0(net36),
    .A1(net55),
    .A2(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.J_NS4_BEG15 ),
    .A3(_0071_),
    .S0(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame7_bit0.Q ),
    .S1(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame7_bit1.Q ),
    .X(_0072_));
 sky130_fd_sc_hd__o21ba_1 _0300_ (.A1(net223),
    .A2(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame0_bit30.Q ),
    .B1_N(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame0_bit31.Q ),
    .X(_0073_));
 sky130_fd_sc_hd__o21a_1 _0301_ (.A1(net166),
    .A2(_0022_),
    .B1(_0073_),
    .X(_0074_));
 sky130_fd_sc_hd__a31o_1 _0302_ (.A1(_0022_),
    .A2(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame0_bit31.Q ),
    .A3(_0072_),
    .B1(_0074_),
    .X(_0075_));
 sky130_fd_sc_hd__mux4_2 _0303_ (.A0(net144),
    .A1(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.J_NS4_BEG15 ),
    .A2(net170),
    .A3(_0075_),
    .S0(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame9_bit21.Q ),
    .S1(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame9_bit20.Q ),
    .X(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.N1END3 ));
 sky130_fd_sc_hd__mux4_2 _0304_ (.A0(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.N1END3 ),
    .A1(net247),
    .A2(net116),
    .A3(net136),
    .S0(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame0_bit6.Q ),
    .S1(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame0_bit7.Q ),
    .X(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.J_NS4_BEG15 ));
 sky130_fd_sc_hd__mux4_1 _0305_ (.A0(net36),
    .A1(net62),
    .A2(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.J_NS4_BEG15 ),
    .A3(_0071_),
    .S0(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame9_bit28.Q ),
    .S1(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame9_bit29.Q ),
    .X(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.N1BEG3 ));
 sky130_fd_sc_hd__mux4_2 _0306_ (.A0(net52),
    .A1(net44),
    .A2(net63),
    .A3(net364),
    .S0(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame7_bit2.Q ),
    .S1(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame7_bit3.Q ),
    .X(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.S2BEG0 ));
 sky130_fd_sc_hd__mux4_1 _0307_ (.A0(net232),
    .A1(net224),
    .A2(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.S2BEG0 ),
    .A3(net125),
    .S0(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame0_bit8.Q ),
    .S1(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame0_bit9.Q ),
    .X(_0076_));
 sky130_fd_sc_hd__mux4_1 _0308_ (.A0(net160),
    .A1(net152),
    .A2(net170),
    .A3(net369),
    .S0(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame9_bit22.Q ),
    .S1(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame9_bit23.Q ),
    .X(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.N2BEGb0 ));
 sky130_fd_sc_hd__mux4_1 _0309_ (.A0(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.N2BEGb0 ),
    .A1(net125),
    .A2(net232),
    .A3(net117),
    .S0(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame0_bit9.Q ),
    .S1(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame0_bit8.Q ),
    .X(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.J_NS2_BEG0 ));
 sky130_fd_sc_hd__mux4_1 _0310_ (.A0(net52),
    .A1(net44),
    .A2(net62),
    .A3(net364),
    .S0(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame9_bit30.Q ),
    .S1(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame9_bit31.Q ),
    .X(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.N2BEG0 ));
 sky130_fd_sc_hd__mux4_2 _0311_ (.A0(net51),
    .A1(net43),
    .A2(net64),
    .A3(net363),
    .S0(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame7_bit4.Q ),
    .S1(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame7_bit5.Q ),
    .X(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.S2BEG1 ));
 sky130_fd_sc_hd__mux4_1 _0312_ (.A0(net233),
    .A1(net225),
    .A2(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.S2BEG1 ),
    .A3(net126),
    .S0(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame0_bit10.Q ),
    .S1(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame0_bit11.Q ),
    .X(_0077_));
 sky130_fd_sc_hd__mux4_1 _0313_ (.A0(net159),
    .A1(net151),
    .A2(net169),
    .A3(net368),
    .S0(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame9_bit24.Q ),
    .S1(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame9_bit25.Q ),
    .X(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.N2BEGb1 ));
 sky130_fd_sc_hd__mux4_1 _0314_ (.A0(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.N2BEGb1 ),
    .A1(net126),
    .A2(net233),
    .A3(net118),
    .S0(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame0_bit11.Q ),
    .S1(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame0_bit10.Q ),
    .X(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.J_NS2_BEG1 ));
 sky130_fd_sc_hd__mux4_1 _0315_ (.A0(net51),
    .A1(net43),
    .A2(net61),
    .A3(net363),
    .S0(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame8_bit0.Q ),
    .S1(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame8_bit1.Q ),
    .X(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.N2BEG1 ));
 sky130_fd_sc_hd__mux4_2 _0316_ (.A0(net50),
    .A1(net42),
    .A2(net54),
    .A3(net362),
    .S0(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame7_bit6.Q ),
    .S1(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame7_bit7.Q ),
    .X(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.S2BEG2 ));
 sky130_fd_sc_hd__mux4_1 _0317_ (.A0(net234),
    .A1(net226),
    .A2(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.S2BEG2 ),
    .A3(net127),
    .S0(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame0_bit12.Q ),
    .S1(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame0_bit13.Q ),
    .X(_0078_));
 sky130_fd_sc_hd__mux4_1 _0318_ (.A0(net158),
    .A1(net150),
    .A2(net168),
    .A3(net367),
    .S0(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame9_bit26.Q ),
    .S1(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame9_bit27.Q ),
    .X(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.N2BEGb2 ));
 sky130_fd_sc_hd__mux4_1 _0319_ (.A0(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.N2BEGb2 ),
    .A1(net127),
    .A2(net234),
    .A3(net119),
    .S0(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame0_bit13.Q ),
    .S1(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame0_bit12.Q ),
    .X(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.J_NS2_BEG2 ));
 sky130_fd_sc_hd__mux4_1 _0320_ (.A0(net50),
    .A1(net42),
    .A2(net60),
    .A3(net362),
    .S0(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame8_bit2.Q ),
    .S1(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame8_bit3.Q ),
    .X(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.N2BEG2 ));
 sky130_fd_sc_hd__mux4_2 _0321_ (.A0(net49),
    .A1(net41),
    .A2(net55),
    .A3(net361),
    .S0(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame7_bit8.Q ),
    .S1(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame7_bit9.Q ),
    .X(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.S2BEG3 ));
 sky130_fd_sc_hd__mux4_1 _0322_ (.A0(net235),
    .A1(net227),
    .A2(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.S2BEG3 ),
    .A3(net128),
    .S0(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame0_bit14.Q ),
    .S1(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame0_bit15.Q ),
    .X(_0079_));
 sky130_fd_sc_hd__mux4_1 _0323_ (.A0(net157),
    .A1(net149),
    .A2(net167),
    .A3(_0079_),
    .S0(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame9_bit28.Q ),
    .S1(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame9_bit29.Q ),
    .X(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.N2BEGb3 ));
 sky130_fd_sc_hd__mux4_2 _0324_ (.A0(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.N2BEGb3 ),
    .A1(net128),
    .A2(net235),
    .A3(net120),
    .S0(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame0_bit15.Q ),
    .S1(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame0_bit14.Q ),
    .X(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.J_NS2_BEG3 ));
 sky130_fd_sc_hd__mux4_1 _0325_ (.A0(net49),
    .A1(net41),
    .A2(net59),
    .A3(net361),
    .S0(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame8_bit4.Q ),
    .S1(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame8_bit5.Q ),
    .X(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.N2BEG3 ));
 sky130_fd_sc_hd__mux4_2 _0326_ (.A0(net33),
    .A1(net40),
    .A2(net48),
    .A3(net360),
    .S0(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame7_bit11.Q ),
    .S1(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame7_bit10.Q ),
    .X(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.S2BEG4 ));
 sky130_fd_sc_hd__mux4_1 _0327_ (.A0(net236),
    .A1(net228),
    .A2(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.S2BEG4 ),
    .A3(net129),
    .S0(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame0_bit16.Q ),
    .S1(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame0_bit17.Q ),
    .X(_0080_));
 sky130_fd_sc_hd__mux4_1 _0328_ (.A0(net156),
    .A1(net148),
    .A2(net166),
    .A3(_0080_),
    .S0(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame9_bit30.Q ),
    .S1(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame9_bit31.Q ),
    .X(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.N2BEGb4 ));
 sky130_fd_sc_hd__mux4_1 _0329_ (.A0(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.N2BEGb4 ),
    .A1(net129),
    .A2(net236),
    .A3(net121),
    .S0(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame0_bit17.Q ),
    .S1(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame0_bit16.Q ),
    .X(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.J_NS2_BEG4 ));
 sky130_fd_sc_hd__mux4_1 _0330_ (.A0(net48),
    .A1(net40),
    .A2(net58),
    .A3(net360),
    .S0(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame8_bit6.Q ),
    .S1(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame8_bit7.Q ),
    .X(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.N2BEG4 ));
 sky130_fd_sc_hd__mux4_1 _0331_ (.A0(net34),
    .A1(net47),
    .A2(net39),
    .A3(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.J_NS2_BEG5 ),
    .S0(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame7_bit12.Q ),
    .S1(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame7_bit13.Q ),
    .X(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.S2BEG5 ));
 sky130_fd_sc_hd__mux4_2 _0332_ (.A0(net237),
    .A1(net229),
    .A2(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.S2BEG5 ),
    .A3(net130),
    .S0(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame0_bit18.Q ),
    .S1(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame0_bit19.Q ),
    .X(_0081_));
 sky130_fd_sc_hd__mux4_1 _0333_ (.A0(net155),
    .A1(net147),
    .A2(net165),
    .A3(_0081_),
    .S0(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame8_bit0.Q ),
    .S1(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame8_bit1.Q ),
    .X(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.N2BEGb5 ));
 sky130_fd_sc_hd__mux4_2 _0334_ (.A0(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.N2BEGb5 ),
    .A1(net130),
    .A2(net237),
    .A3(net122),
    .S0(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame0_bit19.Q ),
    .S1(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame0_bit18.Q ),
    .X(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.J_NS2_BEG5 ));
 sky130_fd_sc_hd__mux4_1 _0335_ (.A0(net47),
    .A1(net39),
    .A2(net57),
    .A3(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.J_NS2_BEG5 ),
    .S0(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame8_bit8.Q ),
    .S1(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame8_bit9.Q ),
    .X(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.N2BEG5 ));
 sky130_fd_sc_hd__mux4_1 _0336_ (.A0(net35),
    .A1(net46),
    .A2(net38),
    .A3(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.J_NS2_BEG6 ),
    .S0(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame7_bit14.Q ),
    .S1(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame7_bit15.Q ),
    .X(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.S2BEG6 ));
 sky130_fd_sc_hd__mux4_2 _0337_ (.A0(net238),
    .A1(net230),
    .A2(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.S2BEG6 ),
    .A3(net131),
    .S0(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame0_bit20.Q ),
    .S1(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame0_bit21.Q ),
    .X(_0082_));
 sky130_fd_sc_hd__mux4_1 _0338_ (.A0(net154),
    .A1(net146),
    .A2(net164),
    .A3(_0082_),
    .S0(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame8_bit2.Q ),
    .S1(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame8_bit3.Q ),
    .X(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.N2BEGb6 ));
 sky130_fd_sc_hd__mux4_2 _0339_ (.A0(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.N2BEGb6 ),
    .A1(net131),
    .A2(net238),
    .A3(net123),
    .S0(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame0_bit21.Q ),
    .S1(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame0_bit20.Q ),
    .X(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.J_NS2_BEG6 ));
 sky130_fd_sc_hd__mux4_1 _0340_ (.A0(net46),
    .A1(net38),
    .A2(net56),
    .A3(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.J_NS2_BEG6 ),
    .S0(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame8_bit10.Q ),
    .S1(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame8_bit11.Q ),
    .X(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.N2BEG6 ));
 sky130_fd_sc_hd__mux4_1 _0341_ (.A0(net36),
    .A1(net45),
    .A2(net37),
    .A3(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.J_NS2_BEG7 ),
    .S0(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame7_bit16.Q ),
    .S1(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame7_bit17.Q ),
    .X(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.S2BEG7 ));
 sky130_fd_sc_hd__mux4_2 _0342_ (.A0(net239),
    .A1(net231),
    .A2(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.S2BEG7 ),
    .A3(net132),
    .S0(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame0_bit22.Q ),
    .S1(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame0_bit23.Q ),
    .X(_0083_));
 sky130_fd_sc_hd__mux4_2 _0343_ (.A0(net153),
    .A1(net145),
    .A2(net161),
    .A3(_0083_),
    .S0(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame8_bit4.Q ),
    .S1(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame8_bit5.Q ),
    .X(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.N2BEGb7 ));
 sky130_fd_sc_hd__mux4_2 _0344_ (.A0(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.N2BEGb7 ),
    .A1(net132),
    .A2(net239),
    .A3(net124),
    .S0(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame0_bit23.Q ),
    .S1(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame0_bit22.Q ),
    .X(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.J_NS2_BEG7 ));
 sky130_fd_sc_hd__mux4_1 _0345_ (.A0(net45),
    .A1(net37),
    .A2(net53),
    .A3(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.J_NS2_BEG7 ),
    .S0(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame8_bit12.Q ),
    .S1(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame8_bit13.Q ),
    .X(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.N2BEG7 ));
 sky130_fd_sc_hd__mux2_1 _0346_ (.A0(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.N1END0 ),
    .A1(net53),
    .S(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame0_bit24.Q ),
    .X(_0084_));
 sky130_fd_sc_hd__and3b_1 _0347_ (.A_N(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame0_bit24.Q ),
    .B(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame0_bit25.Q ),
    .C(net113),
    .X(_0085_));
 sky130_fd_sc_hd__a21o_1 _0348_ (.A1(_0019_),
    .A2(_0084_),
    .B1(_0085_),
    .X(_0086_));
 sky130_fd_sc_hd__mux4_2 _0349_ (.A0(net33),
    .A1(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.J_NS4_BEG12 ),
    .A2(net63),
    .A3(_0086_),
    .S0(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame8_bit27.Q ),
    .S1(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame8_bit26.Q ),
    .X(_0087_));
 sky130_fd_sc_hd__o21ba_1 _0350_ (.A1(net220),
    .A2(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame0_bit24.Q ),
    .B1_N(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame0_bit25.Q ),
    .X(_0088_));
 sky130_fd_sc_hd__o21a_1 _0351_ (.A1(net161),
    .A2(_0018_),
    .B1(_0088_),
    .X(_0089_));
 sky130_fd_sc_hd__a31o_1 _0352_ (.A1(_0018_),
    .A2(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame0_bit25.Q ),
    .A3(_0087_),
    .B1(_0089_),
    .X(_0090_));
 sky130_fd_sc_hd__mux4_2 _0353_ (.A0(net141),
    .A1(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.J_NS4_BEG12 ),
    .A2(net167),
    .A3(_0090_),
    .S0(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame9_bit15.Q ),
    .S1(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame9_bit14.Q ),
    .X(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.N1END0 ));
 sky130_fd_sc_hd__mux4_1 _0354_ (.A0(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.N1END0 ),
    .A1(net11),
    .A2(net113),
    .A3(net17),
    .S0(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame7_bit31.Q ),
    .S1(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame7_bit30.Q ),
    .X(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.W1BEG0 ));
 sky130_fd_sc_hd__mux4_1 _0355_ (.A0(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.N1END1 ),
    .A1(net12),
    .A2(net114),
    .A3(net16),
    .S0(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame6_bit1.Q ),
    .S1(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame6_bit0.Q ),
    .X(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.W1BEG1 ));
 sky130_fd_sc_hd__mux4_1 _0356_ (.A0(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.N1END2 ),
    .A1(net9),
    .A2(net115),
    .A3(net15),
    .S0(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame6_bit3.Q ),
    .S1(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame6_bit2.Q ),
    .X(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.W1BEG2 ));
 sky130_fd_sc_hd__mux4_1 _0357_ (.A0(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.N1END3 ),
    .A1(net10),
    .A2(net116),
    .A3(net14),
    .S0(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame6_bit5.Q ),
    .S1(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame6_bit4.Q ),
    .X(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.W1BEG3 ));
 sky130_fd_sc_hd__mux4_1 _0358_ (.A0(net9),
    .A1(net18),
    .A2(net364),
    .A3(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.J_NS2_BEG7 ),
    .S0(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame6_bit6.Q ),
    .S1(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame6_bit7.Q ),
    .X(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.W2BEG0 ));
 sky130_fd_sc_hd__mux4_1 _0359_ (.A0(net10),
    .A1(net19),
    .A2(net363),
    .A3(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.J_NS2_BEG6 ),
    .S0(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame6_bit8.Q ),
    .S1(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame6_bit9.Q ),
    .X(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.W2BEG1 ));
 sky130_fd_sc_hd__mux4_1 _0360_ (.A0(net11),
    .A1(net20),
    .A2(net362),
    .A3(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.J_NS2_BEG5 ),
    .S0(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame6_bit10.Q ),
    .S1(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame6_bit11.Q ),
    .X(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.W2BEG2 ));
 sky130_fd_sc_hd__mux4_1 _0361_ (.A0(net12),
    .A1(net21),
    .A2(net361),
    .A3(net360),
    .S0(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame6_bit12.Q ),
    .S1(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame6_bit13.Q ),
    .X(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.W2BEG3 ));
 sky130_fd_sc_hd__mux4_1 _0362_ (.A0(net14),
    .A1(net22),
    .A2(net361),
    .A3(net360),
    .S0(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame6_bit14.Q ),
    .S1(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame6_bit15.Q ),
    .X(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.W2BEG4 ));
 sky130_fd_sc_hd__mux4_1 _0363_ (.A0(net15),
    .A1(net23),
    .A2(net362),
    .A3(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.J_NS2_BEG5 ),
    .S0(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame6_bit16.Q ),
    .S1(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame6_bit17.Q ),
    .X(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.W2BEG5 ));
 sky130_fd_sc_hd__mux4_1 _0364_ (.A0(net16),
    .A1(net25),
    .A2(net363),
    .A3(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.J_NS2_BEG6 ),
    .S0(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame6_bit18.Q ),
    .S1(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame6_bit19.Q ),
    .X(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.W2BEG6 ));
 sky130_fd_sc_hd__mux4_1 _0365_ (.A0(net17),
    .A1(net26),
    .A2(net364),
    .A3(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.J_NS2_BEG7 ),
    .S0(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame6_bit20.Q ),
    .S1(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame6_bit21.Q ),
    .X(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.W2BEG7 ));
 sky130_fd_sc_hd__mux4_1 _0366_ (.A0(net9),
    .A1(net18),
    .A2(net364),
    .A3(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.J_NS2_BEG7 ),
    .S0(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame6_bit22.Q ),
    .S1(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame6_bit23.Q ),
    .X(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.W2BEGb0 ));
 sky130_fd_sc_hd__mux4_1 _0367_ (.A0(net10),
    .A1(net19),
    .A2(net363),
    .A3(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.J_NS2_BEG6 ),
    .S0(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame6_bit24.Q ),
    .S1(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame6_bit25.Q ),
    .X(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.W2BEGb1 ));
 sky130_fd_sc_hd__mux4_1 _0368_ (.A0(net11),
    .A1(net20),
    .A2(net362),
    .A3(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.J_NS2_BEG5 ),
    .S0(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame6_bit26.Q ),
    .S1(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame6_bit27.Q ),
    .X(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.W2BEGb2 ));
 sky130_fd_sc_hd__mux4_1 _0369_ (.A0(net12),
    .A1(net21),
    .A2(net361),
    .A3(net360),
    .S0(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame6_bit28.Q ),
    .S1(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame6_bit29.Q ),
    .X(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.W2BEGb3 ));
 sky130_fd_sc_hd__mux4_1 _0370_ (.A0(net14),
    .A1(net22),
    .A2(net361),
    .A3(net360),
    .S0(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame6_bit30.Q ),
    .S1(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame6_bit31.Q ),
    .X(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.W2BEGb4 ));
 sky130_fd_sc_hd__mux4_1 _0371_ (.A0(net15),
    .A1(net23),
    .A2(net362),
    .A3(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.J_NS2_BEG5 ),
    .S0(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame5_bit0.Q ),
    .S1(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame5_bit1.Q ),
    .X(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.W2BEGb5 ));
 sky130_fd_sc_hd__mux4_1 _0372_ (.A0(net16),
    .A1(net25),
    .A2(net363),
    .A3(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.J_NS2_BEG6 ),
    .S0(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame5_bit2.Q ),
    .S1(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame5_bit3.Q ),
    .X(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.W2BEGb6 ));
 sky130_fd_sc_hd__mux4_1 _0373_ (.A0(net17),
    .A1(net26),
    .A2(net364),
    .A3(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.J_NS2_BEG7 ),
    .S0(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame5_bit4.Q ),
    .S1(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame5_bit5.Q ),
    .X(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.W2BEGb7 ));
 sky130_fd_sc_hd__mux4_1 _0374_ (.A0(net9),
    .A1(net22),
    .A2(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.J_NS4_BEG15 ),
    .A3(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.J_NS2_BEG7 ),
    .S0(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame5_bit6.Q ),
    .S1(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame5_bit7.Q ),
    .X(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.WW4BEG0 ));
 sky130_fd_sc_hd__mux4_1 _0375_ (.A0(net10),
    .A1(net23),
    .A2(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.J_NS4_BEG14 ),
    .A3(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.J_NS2_BEG6 ),
    .S0(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame5_bit8.Q ),
    .S1(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame5_bit9.Q ),
    .X(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.WW4BEG1 ));
 sky130_fd_sc_hd__mux4_1 _0376_ (.A0(net11),
    .A1(net25),
    .A2(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.J_NS4_BEG13 ),
    .A3(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.J_NS2_BEG5 ),
    .S0(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame5_bit10.Q ),
    .S1(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame5_bit11.Q ),
    .X(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.WW4BEG2 ));
 sky130_fd_sc_hd__mux4_2 _0377_ (.A0(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.N1END0 ),
    .A1(net244),
    .A2(net113),
    .A3(net133),
    .S0(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame0_bit0.Q ),
    .S1(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame0_bit1.Q ),
    .X(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.J_NS4_BEG12 ));
 sky130_fd_sc_hd__mux4_1 _0378_ (.A0(net12),
    .A1(net26),
    .A2(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.J_NS4_BEG12 ),
    .A3(net360),
    .S0(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame5_bit12.Q ),
    .S1(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame5_bit13.Q ),
    .X(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.WW4BEG3 ));
 sky130_fd_sc_hd__mux4_2 _0379_ (.A0(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.N1END3 ),
    .A1(net247),
    .A2(net116),
    .A3(net136),
    .S0(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame1_bit30.Q ),
    .S1(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame1_bit31.Q ),
    .X(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.J_NS4_BEG11 ));
 sky130_fd_sc_hd__mux4_1 _0380_ (.A0(net14),
    .A1(net18),
    .A2(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.J_NS4_BEG11 ),
    .A3(net361),
    .S0(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame5_bit14.Q ),
    .S1(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame5_bit15.Q ),
    .X(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.WW4BEG4 ));
 sky130_fd_sc_hd__mux4_2 _0381_ (.A0(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.N1END2 ),
    .A1(net246),
    .A2(net115),
    .A3(net135),
    .S0(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame1_bit28.Q ),
    .S1(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame1_bit29.Q ),
    .X(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.J_NS4_BEG10 ));
 sky130_fd_sc_hd__mux4_1 _0382_ (.A0(net15),
    .A1(net19),
    .A2(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.J_NS4_BEG10 ),
    .A3(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.J_NS2_BEG2 ),
    .S0(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame5_bit16.Q ),
    .S1(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame5_bit17.Q ),
    .X(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.WW4BEG5 ));
 sky130_fd_sc_hd__mux4_2 _0383_ (.A0(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.N1END1 ),
    .A1(net245),
    .A2(net114),
    .A3(net134),
    .S0(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame1_bit26.Q ),
    .S1(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame1_bit27.Q ),
    .X(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.J_NS4_BEG9 ));
 sky130_fd_sc_hd__mux4_1 _0384_ (.A0(net16),
    .A1(net20),
    .A2(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.J_NS4_BEG9 ),
    .A3(net363),
    .S0(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame5_bit18.Q ),
    .S1(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame5_bit19.Q ),
    .X(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.WW4BEG6 ));
 sky130_fd_sc_hd__mux4_2 _0385_ (.A0(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.N1END0 ),
    .A1(net244),
    .A2(net113),
    .A3(net133),
    .S0(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame1_bit24.Q ),
    .S1(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame1_bit25.Q ),
    .X(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.J_NS4_BEG8 ));
 sky130_fd_sc_hd__mux4_1 _0386_ (.A0(net17),
    .A1(net21),
    .A2(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.J_NS4_BEG8 ),
    .A3(net364),
    .S0(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame5_bit20.Q ),
    .S1(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame5_bit21.Q ),
    .X(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.WW4BEG7 ));
 sky130_fd_sc_hd__mux4_2 _0387_ (.A0(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.N1END3 ),
    .A1(net247),
    .A2(net116),
    .A3(net136),
    .S0(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame1_bit22.Q ),
    .S1(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame1_bit23.Q ),
    .X(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.J_NS4_BEG7 ));
 sky130_fd_sc_hd__mux4_1 _0388_ (.A0(net14),
    .A1(net18),
    .A2(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.J_NS4_BEG7 ),
    .A3(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.J_NS2_BEG7 ),
    .S0(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame5_bit22.Q ),
    .S1(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame5_bit23.Q ),
    .X(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.WW4BEG8 ));
 sky130_fd_sc_hd__mux4_2 _0389_ (.A0(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.N1END2 ),
    .A1(net246),
    .A2(net115),
    .A3(net135),
    .S0(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame1_bit20.Q ),
    .S1(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame1_bit21.Q ),
    .X(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.J_NS4_BEG6 ));
 sky130_fd_sc_hd__mux4_1 _0390_ (.A0(net15),
    .A1(net19),
    .A2(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.J_NS4_BEG6 ),
    .A3(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.J_NS2_BEG6 ),
    .S0(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame5_bit24.Q ),
    .S1(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame5_bit25.Q ),
    .X(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.WW4BEG9 ));
 sky130_fd_sc_hd__mux4_2 _0391_ (.A0(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.N1END1 ),
    .A1(net245),
    .A2(net114),
    .A3(net134),
    .S0(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame1_bit18.Q ),
    .S1(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame1_bit19.Q ),
    .X(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.J_NS4_BEG5 ));
 sky130_fd_sc_hd__mux4_1 _0392_ (.A0(net16),
    .A1(net20),
    .A2(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.J_NS4_BEG5 ),
    .A3(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.J_NS2_BEG5 ),
    .S0(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame5_bit26.Q ),
    .S1(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame5_bit27.Q ),
    .X(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.WW4BEG10 ));
 sky130_fd_sc_hd__mux4_2 _0393_ (.A0(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.N1END0 ),
    .A1(net244),
    .A2(net113),
    .A3(net133),
    .S0(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame1_bit16.Q ),
    .S1(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame1_bit17.Q ),
    .X(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.J_NS4_BEG4 ));
 sky130_fd_sc_hd__mux4_1 _0394_ (.A0(net17),
    .A1(net21),
    .A2(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.J_NS4_BEG4 ),
    .A3(net360),
    .S0(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame5_bit28.Q ),
    .S1(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame5_bit29.Q ),
    .X(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.WW4BEG11 ));
 sky130_fd_sc_hd__mux4_2 _0395_ (.A0(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.N1END3 ),
    .A1(net247),
    .A2(net116),
    .A3(net136),
    .S0(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame1_bit14.Q ),
    .S1(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame1_bit15.Q ),
    .X(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.J_NS4_BEG3 ));
 sky130_fd_sc_hd__mux4_1 _0396_ (.A0(net9),
    .A1(net22),
    .A2(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.J_NS4_BEG3 ),
    .A3(net361),
    .S0(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame5_bit30.Q ),
    .S1(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame5_bit31.Q ),
    .X(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.WW4BEG12 ));
 sky130_fd_sc_hd__mux4_2 _0397_ (.A0(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.N1END2 ),
    .A1(net246),
    .A2(net115),
    .A3(net135),
    .S0(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame1_bit12.Q ),
    .S1(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame1_bit13.Q ),
    .X(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.J_NS4_BEG2 ));
 sky130_fd_sc_hd__mux4_1 _0398_ (.A0(net10),
    .A1(net23),
    .A2(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.J_NS4_BEG2 ),
    .A3(net362),
    .S0(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame4_bit0.Q ),
    .S1(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame4_bit1.Q ),
    .X(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.WW4BEG13 ));
 sky130_fd_sc_hd__mux4_2 _0399_ (.A0(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.N1END1 ),
    .A1(net245),
    .A2(net114),
    .A3(net134),
    .S0(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame1_bit10.Q ),
    .S1(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame1_bit11.Q ),
    .X(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.J_NS4_BEG1 ));
 sky130_fd_sc_hd__mux4_1 _0400_ (.A0(net11),
    .A1(net25),
    .A2(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.J_NS4_BEG1 ),
    .A3(net363),
    .S0(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame4_bit2.Q ),
    .S1(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame4_bit3.Q ),
    .X(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.WW4BEG14 ));
 sky130_fd_sc_hd__mux4_2 _0401_ (.A0(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.N1END0 ),
    .A1(net244),
    .A2(net113),
    .A3(net133),
    .S0(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame1_bit8.Q ),
    .S1(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame1_bit9.Q ),
    .X(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.J_NS4_BEG0 ));
 sky130_fd_sc_hd__mux4_1 _0402_ (.A0(net12),
    .A1(net26),
    .A2(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.J_NS4_BEG0 ),
    .A3(net364),
    .S0(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame4_bit4.Q ),
    .S1(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame4_bit5.Q ),
    .X(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.WW4BEG15 ));
 sky130_fd_sc_hd__mux4_1 _0403_ (.A0(net244),
    .A1(net133),
    .A2(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.J_NS4_BEG11 ),
    .A3(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.J_NS4_BEG15 ),
    .S0(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame4_bit6.Q ),
    .S1(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame4_bit7.Q ),
    .X(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.W6BEG0 ));
 sky130_fd_sc_hd__mux4_1 _0404_ (.A0(net245),
    .A1(net134),
    .A2(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.J_NS4_BEG10 ),
    .A3(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.J_NS4_BEG14 ),
    .S0(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame4_bit8.Q ),
    .S1(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame4_bit9.Q ),
    .X(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.W6BEG1 ));
 sky130_fd_sc_hd__mux4_1 _0405_ (.A0(net246),
    .A1(net135),
    .A2(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.J_NS4_BEG9 ),
    .A3(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.J_NS4_BEG13 ),
    .S0(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame4_bit10.Q ),
    .S1(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame4_bit11.Q ),
    .X(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.W6BEG2 ));
 sky130_fd_sc_hd__mux4_1 _0406_ (.A0(net247),
    .A1(net136),
    .A2(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.J_NS4_BEG8 ),
    .A3(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.J_NS4_BEG12 ),
    .S0(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame4_bit12.Q ),
    .S1(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame4_bit13.Q ),
    .X(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.W6BEG3 ));
 sky130_fd_sc_hd__mux4_1 _0407_ (.A0(net14),
    .A1(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.J_NS4_BEG11 ),
    .A2(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.J_NS4_BEG7 ),
    .A3(net364),
    .S0(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame4_bit15.Q ),
    .S1(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame4_bit14.Q ),
    .X(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.W6BEG4 ));
 sky130_fd_sc_hd__mux4_1 _0408_ (.A0(net15),
    .A1(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.J_NS4_BEG10 ),
    .A2(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.J_NS4_BEG6 ),
    .A3(net363),
    .S0(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame4_bit17.Q ),
    .S1(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame4_bit16.Q ),
    .X(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.W6BEG5 ));
 sky130_fd_sc_hd__mux4_1 _0409_ (.A0(net16),
    .A1(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.J_NS4_BEG5 ),
    .A2(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.J_NS4_BEG9 ),
    .A3(net362),
    .S0(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame4_bit18.Q ),
    .S1(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame4_bit19.Q ),
    .X(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.W6BEG6 ));
 sky130_fd_sc_hd__mux4_1 _0410_ (.A0(net17),
    .A1(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.J_NS4_BEG4 ),
    .A2(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.J_NS4_BEG8 ),
    .A3(net361),
    .S0(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame4_bit20.Q ),
    .S1(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame4_bit21.Q ),
    .X(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.W6BEG7 ));
 sky130_fd_sc_hd__mux4_1 _0411_ (.A0(net9),
    .A1(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.J_NS4_BEG7 ),
    .A2(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.J_NS4_BEG3 ),
    .A3(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.J_NS2_BEG4 ),
    .S0(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame4_bit23.Q ),
    .S1(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame4_bit22.Q ),
    .X(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.W6BEG8 ));
 sky130_fd_sc_hd__mux4_1 _0412_ (.A0(net10),
    .A1(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.J_NS4_BEG6 ),
    .A2(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.J_NS4_BEG2 ),
    .A3(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.J_NS2_BEG5 ),
    .S0(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame4_bit25.Q ),
    .S1(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame4_bit24.Q ),
    .X(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.W6BEG9 ));
 sky130_fd_sc_hd__mux4_1 _0413_ (.A0(net11),
    .A1(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.J_NS4_BEG5 ),
    .A2(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.J_NS4_BEG1 ),
    .A3(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.J_NS2_BEG6 ),
    .S0(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame4_bit27.Q ),
    .S1(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame4_bit26.Q ),
    .X(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.W6BEG10 ));
 sky130_fd_sc_hd__mux4_1 _0414_ (.A0(net12),
    .A1(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.J_NS4_BEG4 ),
    .A2(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.J_NS4_BEG0 ),
    .A3(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.J_NS2_BEG7 ),
    .S0(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame4_bit29.Q ),
    .S1(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame4_bit28.Q ),
    .X(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.W6BEG11 ));
 sky130_fd_sc_hd__mux4_1 _0415_ (.A0(net65),
    .A1(net79),
    .A2(net53),
    .A3(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.J_NS4_BEG0 ),
    .S0(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame4_bit30.Q ),
    .S1(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame4_bit31.Q ),
    .X(net299));
 sky130_fd_sc_hd__mux4_2 _0416_ (.A0(net72),
    .A1(net80),
    .A2(net56),
    .A3(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.J_NS4_BEG1 ),
    .S0(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame3_bit0.Q ),
    .S1(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame3_bit1.Q ),
    .X(net300));
 sky130_fd_sc_hd__mux4_2 _0417_ (.A0(net73),
    .A1(net66),
    .A2(net57),
    .A3(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.J_NS4_BEG2 ),
    .S0(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame3_bit2.Q ),
    .S1(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame3_bit3.Q ),
    .X(net301));
 sky130_fd_sc_hd__mux4_2 _0418_ (.A0(net74),
    .A1(net67),
    .A2(net58),
    .A3(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.J_NS4_BEG3 ),
    .S0(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame3_bit4.Q ),
    .S1(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame3_bit5.Q ),
    .X(net302));
 sky130_fd_sc_hd__mux4_1 _0419_ (.A0(net75),
    .A1(net68),
    .A2(net59),
    .A3(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.J_NS4_BEG4 ),
    .S0(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame3_bit6.Q ),
    .S1(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame3_bit7.Q ),
    .X(net304));
 sky130_fd_sc_hd__mux4_2 _0420_ (.A0(net76),
    .A1(net69),
    .A2(net60),
    .A3(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.J_NS4_BEG5 ),
    .S0(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame3_bit8.Q ),
    .S1(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame3_bit9.Q ),
    .X(net305));
 sky130_fd_sc_hd__mux4_2 _0421_ (.A0(net77),
    .A1(net70),
    .A2(net61),
    .A3(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.J_NS4_BEG6 ),
    .S0(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame3_bit10.Q ),
    .S1(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame3_bit11.Q ),
    .X(net306));
 sky130_fd_sc_hd__mux4_2 _0422_ (.A0(net78),
    .A1(net71),
    .A2(net62),
    .A3(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.J_NS4_BEG7 ),
    .S0(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame3_bit12.Q ),
    .S1(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame3_bit13.Q ),
    .X(net307));
 sky130_fd_sc_hd__mux4_1 _0423_ (.A0(net65),
    .A1(net79),
    .A2(net63),
    .A3(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.J_NS4_BEG8 ),
    .S0(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame3_bit14.Q ),
    .S1(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame3_bit15.Q ),
    .X(net308));
 sky130_fd_sc_hd__mux4_2 _0424_ (.A0(net72),
    .A1(net80),
    .A2(net64),
    .A3(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.J_NS4_BEG9 ),
    .S0(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame3_bit16.Q ),
    .S1(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame3_bit17.Q ),
    .X(net309));
 sky130_fd_sc_hd__mux4_2 _0425_ (.A0(net73),
    .A1(net66),
    .A2(net54),
    .A3(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.J_NS4_BEG10 ),
    .S0(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame3_bit18.Q ),
    .S1(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame3_bit19.Q ),
    .X(net310));
 sky130_fd_sc_hd__mux4_2 _0426_ (.A0(net74),
    .A1(net67),
    .A2(net55),
    .A3(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.J_NS4_BEG11 ),
    .S0(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame3_bit20.Q ),
    .S1(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame3_bit21.Q ),
    .X(net311));
 sky130_fd_sc_hd__mux4_1 _0427_ (.A0(net33),
    .A1(net75),
    .A2(net68),
    .A3(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.J_NS4_BEG12 ),
    .S0(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame3_bit22.Q ),
    .S1(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame3_bit23.Q ),
    .X(net312));
 sky130_fd_sc_hd__mux4_2 _0428_ (.A0(net34),
    .A1(net76),
    .A2(net69),
    .A3(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.J_NS4_BEG13 ),
    .S0(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame3_bit24.Q ),
    .S1(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame3_bit25.Q ),
    .X(net313));
 sky130_fd_sc_hd__mux4_2 _0429_ (.A0(net35),
    .A1(net77),
    .A2(net70),
    .A3(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.J_NS4_BEG14 ),
    .S0(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame3_bit26.Q ),
    .S1(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame3_bit27.Q ),
    .X(net315));
 sky130_fd_sc_hd__mux4_2 _0430_ (.A0(net36),
    .A1(net78),
    .A2(net71),
    .A3(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.J_NS4_BEG15 ),
    .S0(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame3_bit28.Q ),
    .S1(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame3_bit29.Q ),
    .X(net316));
 sky130_fd_sc_hd__mux4_1 _0431_ (.A0(net65),
    .A1(net79),
    .A2(net53),
    .A3(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.J_NS4_BEG0 ),
    .S0(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame3_bit30.Q ),
    .S1(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame3_bit31.Q ),
    .X(net266));
 sky130_fd_sc_hd__mux4_2 _0432_ (.A0(net72),
    .A1(net80),
    .A2(net56),
    .A3(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.J_NS4_BEG1 ),
    .S0(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame2_bit0.Q ),
    .S1(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame2_bit1.Q ),
    .X(net267));
 sky130_fd_sc_hd__mux4_2 _0433_ (.A0(net73),
    .A1(net66),
    .A2(net57),
    .A3(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.J_NS4_BEG2 ),
    .S0(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame2_bit2.Q ),
    .S1(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame2_bit3.Q ),
    .X(net268));
 sky130_fd_sc_hd__mux4_2 _0434_ (.A0(net74),
    .A1(net67),
    .A2(net58),
    .A3(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.J_NS4_BEG3 ),
    .S0(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame2_bit4.Q ),
    .S1(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame2_bit5.Q ),
    .X(net269));
 sky130_fd_sc_hd__mux4_2 _0435_ (.A0(net75),
    .A1(net68),
    .A2(net59),
    .A3(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.J_NS4_BEG4 ),
    .S0(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame2_bit6.Q ),
    .S1(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame2_bit7.Q ),
    .X(net271));
 sky130_fd_sc_hd__mux4_2 _0436_ (.A0(net76),
    .A1(net69),
    .A2(net60),
    .A3(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.J_NS4_BEG5 ),
    .S0(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame2_bit8.Q ),
    .S1(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame2_bit9.Q ),
    .X(net272));
 sky130_fd_sc_hd__mux4_2 _0437_ (.A0(net77),
    .A1(net70),
    .A2(net61),
    .A3(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.J_NS4_BEG6 ),
    .S0(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame2_bit10.Q ),
    .S1(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame2_bit11.Q ),
    .X(net273));
 sky130_fd_sc_hd__mux4_2 _0438_ (.A0(net78),
    .A1(net71),
    .A2(net62),
    .A3(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.J_NS4_BEG7 ),
    .S0(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame2_bit12.Q ),
    .S1(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame2_bit13.Q ),
    .X(net274));
 sky130_fd_sc_hd__mux4_1 _0439_ (.A0(net65),
    .A1(net79),
    .A2(net63),
    .A3(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.J_NS4_BEG8 ),
    .S0(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame2_bit14.Q ),
    .S1(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame2_bit15.Q ),
    .X(net275));
 sky130_fd_sc_hd__mux4_2 _0440_ (.A0(net72),
    .A1(net80),
    .A2(net64),
    .A3(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.J_NS4_BEG9 ),
    .S0(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame2_bit16.Q ),
    .S1(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame2_bit17.Q ),
    .X(net276));
 sky130_fd_sc_hd__mux4_2 _0441_ (.A0(net73),
    .A1(net66),
    .A2(net54),
    .A3(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.J_NS4_BEG10 ),
    .S0(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame2_bit18.Q ),
    .S1(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame2_bit19.Q ),
    .X(net277));
 sky130_fd_sc_hd__mux4_2 _0442_ (.A0(net74),
    .A1(net67),
    .A2(net55),
    .A3(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.J_NS4_BEG11 ),
    .S0(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame2_bit20.Q ),
    .S1(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame2_bit21.Q ),
    .X(net278));
 sky130_fd_sc_hd__mux4_1 _0443_ (.A0(net33),
    .A1(net75),
    .A2(net68),
    .A3(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.J_NS4_BEG12 ),
    .S0(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame2_bit22.Q ),
    .S1(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame2_bit23.Q ),
    .X(net279));
 sky130_fd_sc_hd__mux4_2 _0444_ (.A0(net34),
    .A1(net76),
    .A2(net69),
    .A3(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.J_NS4_BEG13 ),
    .S0(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame2_bit24.Q ),
    .S1(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame2_bit25.Q ),
    .X(net280));
 sky130_fd_sc_hd__mux4_2 _0445_ (.A0(net35),
    .A1(net77),
    .A2(net70),
    .A3(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.J_NS4_BEG14 ),
    .S0(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame2_bit26.Q ),
    .S1(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame2_bit27.Q ),
    .X(net282));
 sky130_fd_sc_hd__mux4_2 _0446_ (.A0(net36),
    .A1(net78),
    .A2(net71),
    .A3(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.J_NS4_BEG15 ),
    .S0(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame2_bit28.Q ),
    .S1(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame2_bit29.Q ),
    .X(net283));
 sky130_fd_sc_hd__mux2_1 _0447_ (.A0(net45),
    .A1(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.J_NS2_BEG0 ),
    .S(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame2_bit31.Q ),
    .X(_0091_));
 sky130_fd_sc_hd__nand2_1 _0448_ (.A(net37),
    .B(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame2_bit30.Q ),
    .Y(_0092_));
 sky130_fd_sc_hd__a2bb2o_1 _0449_ (.A1_N(_0092_),
    .A2_N(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame2_bit31.Q ),
    .B1(_0003_),
    .B2(_0091_),
    .X(net253));
 sky130_fd_sc_hd__mux2_1 _0450_ (.A0(net46),
    .A1(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.J_NS2_BEG1 ),
    .S(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame1_bit1.Q ),
    .X(_0093_));
 sky130_fd_sc_hd__nand2_1 _0451_ (.A(net38),
    .B(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame1_bit0.Q ),
    .Y(_0094_));
 sky130_fd_sc_hd__a2bb2o_2 _0452_ (.A1_N(_0094_),
    .A2_N(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame1_bit1.Q ),
    .B1(_0004_),
    .B2(_0093_),
    .X(net254));
 sky130_fd_sc_hd__mux2_1 _0453_ (.A0(net47),
    .A1(net362),
    .S(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame1_bit3.Q ),
    .X(_0095_));
 sky130_fd_sc_hd__nand2_1 _0454_ (.A(net39),
    .B(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame1_bit2.Q ),
    .Y(_0096_));
 sky130_fd_sc_hd__a2bb2o_2 _0455_ (.A1_N(_0096_),
    .A2_N(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame1_bit3.Q ),
    .B1(_0005_),
    .B2(_0095_),
    .X(net255));
 sky130_fd_sc_hd__mux2_1 _0456_ (.A0(net48),
    .A1(net361),
    .S(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame1_bit5.Q ),
    .X(_0097_));
 sky130_fd_sc_hd__nand2_1 _0457_ (.A(net40),
    .B(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame1_bit4.Q ),
    .Y(_0098_));
 sky130_fd_sc_hd__a2bb2o_2 _0458_ (.A1_N(_0098_),
    .A2_N(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame1_bit5.Q ),
    .B1(_0006_),
    .B2(_0097_),
    .X(net256));
 sky130_fd_sc_hd__o21ba_1 _0459_ (.A1(net49),
    .A2(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame1_bit7.Q ),
    .B1_N(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame1_bit6.Q ),
    .X(_0099_));
 sky130_fd_sc_hd__o21a_1 _0460_ (.A1(_0007_),
    .A2(net360),
    .B1(_0099_),
    .X(_0100_));
 sky130_fd_sc_hd__a31o_2 _0461_ (.A1(net41),
    .A2(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame1_bit6.Q ),
    .A3(_0007_),
    .B1(_0100_),
    .X(net257));
 sky130_fd_sc_hd__mux4_1 _0462_ (.A0(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.J_NS4_BEG4 ),
    .A1(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.J_NS4_BEG8 ),
    .A2(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.J_NS4_BEG12 ),
    .A3(net364),
    .S0(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame8_bit14.Q ),
    .S1(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame8_bit15.Q ),
    .X(_0101_));
 sky130_fd_sc_hd__nand2b_1 _0463_ (.A_N(net65),
    .B(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame8_bit14.Q ),
    .Y(_0102_));
 sky130_fd_sc_hd__o21ba_1 _0464_ (.A1(net33),
    .A2(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame8_bit14.Q ),
    .B1_N(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame8_bit15.Q ),
    .X(_0103_));
 sky130_fd_sc_hd__mux2_1 _0465_ (.A0(net63),
    .A1(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.J_NS4_BEG0 ),
    .S(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame8_bit14.Q ),
    .X(_0104_));
 sky130_fd_sc_hd__a221o_1 _0466_ (.A1(_0102_),
    .A2(_0103_),
    .B1(_0104_),
    .B2(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame8_bit15.Q ),
    .C1(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame8_bit16.Q ),
    .X(_0105_));
 sky130_fd_sc_hd__o21a_1 _0467_ (.A1(_0010_),
    .A2(_0101_),
    .B1(_0105_),
    .X(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.N4BEG0 ));
 sky130_fd_sc_hd__mux4_1 _0468_ (.A0(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.J_NS4_BEG5 ),
    .A1(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.J_NS4_BEG9 ),
    .A2(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.J_NS4_BEG13 ),
    .A3(net363),
    .S0(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame8_bit17.Q ),
    .S1(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame8_bit18.Q ),
    .X(_0106_));
 sky130_fd_sc_hd__nand2b_1 _0469_ (.A_N(net72),
    .B(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame8_bit17.Q ),
    .Y(_0107_));
 sky130_fd_sc_hd__o21ba_1 _0470_ (.A1(net34),
    .A2(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame8_bit17.Q ),
    .B1_N(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame8_bit18.Q ),
    .X(_0108_));
 sky130_fd_sc_hd__mux2_1 _0471_ (.A0(net64),
    .A1(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.J_NS4_BEG1 ),
    .S(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame8_bit17.Q ),
    .X(_0109_));
 sky130_fd_sc_hd__a221o_1 _0472_ (.A1(_0107_),
    .A2(_0108_),
    .B1(_0109_),
    .B2(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame8_bit18.Q ),
    .C1(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame8_bit19.Q ),
    .X(_0110_));
 sky130_fd_sc_hd__o21a_1 _0473_ (.A1(_0011_),
    .A2(_0106_),
    .B1(_0110_),
    .X(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.N4BEG1 ));
 sky130_fd_sc_hd__mux4_1 _0474_ (.A0(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.J_NS4_BEG6 ),
    .A1(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.J_NS4_BEG10 ),
    .A2(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.J_NS4_BEG14 ),
    .A3(net362),
    .S0(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame8_bit20.Q ),
    .S1(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame8_bit21.Q ),
    .X(_0111_));
 sky130_fd_sc_hd__nand2b_1 _0475_ (.A_N(net73),
    .B(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame8_bit20.Q ),
    .Y(_0112_));
 sky130_fd_sc_hd__o21ba_1 _0476_ (.A1(net35),
    .A2(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame8_bit20.Q ),
    .B1_N(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame8_bit21.Q ),
    .X(_0113_));
 sky130_fd_sc_hd__mux2_1 _0477_ (.A0(net54),
    .A1(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.J_NS4_BEG2 ),
    .S(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame8_bit20.Q ),
    .X(_0114_));
 sky130_fd_sc_hd__a221o_1 _0478_ (.A1(_0112_),
    .A2(_0113_),
    .B1(_0114_),
    .B2(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame8_bit21.Q ),
    .C1(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame8_bit22.Q ),
    .X(_0115_));
 sky130_fd_sc_hd__o21a_1 _0479_ (.A1(_0012_),
    .A2(_0111_),
    .B1(_0115_),
    .X(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.N4BEG2 ));
 sky130_fd_sc_hd__mux4_1 _0480_ (.A0(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.J_NS4_BEG7 ),
    .A1(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.J_NS4_BEG11 ),
    .A2(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.J_NS4_BEG15 ),
    .A3(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.J_NS2_BEG3 ),
    .S0(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame8_bit23.Q ),
    .S1(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame8_bit24.Q ),
    .X(_0116_));
 sky130_fd_sc_hd__nand2b_1 _0481_ (.A_N(net74),
    .B(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame8_bit23.Q ),
    .Y(_0117_));
 sky130_fd_sc_hd__o21ba_1 _0482_ (.A1(net36),
    .A2(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame8_bit23.Q ),
    .B1_N(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame8_bit24.Q ),
    .X(_0118_));
 sky130_fd_sc_hd__mux2_1 _0483_ (.A0(net55),
    .A1(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.J_NS4_BEG3 ),
    .S(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame8_bit23.Q ),
    .X(_0119_));
 sky130_fd_sc_hd__a221o_1 _0484_ (.A1(_0117_),
    .A2(_0118_),
    .B1(_0119_),
    .B2(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame8_bit24.Q ),
    .C1(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame8_bit25.Q ),
    .X(_0120_));
 sky130_fd_sc_hd__o21a_1 _0485_ (.A1(_0013_),
    .A2(_0116_),
    .B1(_0120_),
    .X(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.N4BEG3 ));
 sky130_fd_sc_hd__mux4_1 _0486_ (.A0(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.J_NS4_BEG4 ),
    .A1(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.J_NS4_BEG8 ),
    .A2(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.J_NS4_BEG12 ),
    .A3(net360),
    .S0(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame7_bit18.Q ),
    .S1(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame7_bit19.Q ),
    .X(_0121_));
 sky130_fd_sc_hd__nand2b_1 _0487_ (.A_N(net68),
    .B(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame7_bit18.Q ),
    .Y(_0122_));
 sky130_fd_sc_hd__o21ba_1 _0488_ (.A1(net33),
    .A2(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame7_bit18.Q ),
    .B1_N(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame7_bit19.Q ),
    .X(_0123_));
 sky130_fd_sc_hd__mux2_1 _0489_ (.A0(net59),
    .A1(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.J_NS4_BEG0 ),
    .S(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame7_bit18.Q ),
    .X(_0124_));
 sky130_fd_sc_hd__a221o_1 _0490_ (.A1(_0122_),
    .A2(_0123_),
    .B1(_0124_),
    .B2(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame7_bit19.Q ),
    .C1(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame7_bit20.Q ),
    .X(_0125_));
 sky130_fd_sc_hd__o21a_1 _0491_ (.A1(_0014_),
    .A2(_0121_),
    .B1(_0125_),
    .X(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.S4BEG0 ));
 sky130_fd_sc_hd__mux4_1 _0492_ (.A0(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.J_NS4_BEG5 ),
    .A1(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.J_NS4_BEG9 ),
    .A2(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.J_NS4_BEG13 ),
    .A3(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.J_NS2_BEG5 ),
    .S0(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame7_bit21.Q ),
    .S1(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame7_bit22.Q ),
    .X(_0126_));
 sky130_fd_sc_hd__nand2b_1 _0493_ (.A_N(net69),
    .B(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame7_bit21.Q ),
    .Y(_0127_));
 sky130_fd_sc_hd__o21ba_1 _0494_ (.A1(net34),
    .A2(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame7_bit21.Q ),
    .B1_N(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame7_bit22.Q ),
    .X(_0128_));
 sky130_fd_sc_hd__mux2_1 _0495_ (.A0(net60),
    .A1(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.J_NS4_BEG1 ),
    .S(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame7_bit21.Q ),
    .X(_0129_));
 sky130_fd_sc_hd__a221o_1 _0496_ (.A1(_0127_),
    .A2(_0128_),
    .B1(_0129_),
    .B2(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame7_bit22.Q ),
    .C1(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame7_bit23.Q ),
    .X(_0130_));
 sky130_fd_sc_hd__o21a_1 _0497_ (.A1(_0015_),
    .A2(_0126_),
    .B1(_0130_),
    .X(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.S4BEG1 ));
 sky130_fd_sc_hd__mux4_1 _0498_ (.A0(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.J_NS4_BEG6 ),
    .A1(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.J_NS4_BEG10 ),
    .A2(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.J_NS4_BEG14 ),
    .A3(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.J_NS2_BEG6 ),
    .S0(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame7_bit24.Q ),
    .S1(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame7_bit25.Q ),
    .X(_0131_));
 sky130_fd_sc_hd__nand2b_1 _0499_ (.A_N(net70),
    .B(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame7_bit24.Q ),
    .Y(_0132_));
 sky130_fd_sc_hd__o21ba_1 _0500_ (.A1(net35),
    .A2(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame7_bit24.Q ),
    .B1_N(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame7_bit25.Q ),
    .X(_0133_));
 sky130_fd_sc_hd__mux2_1 _0501_ (.A0(net61),
    .A1(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.J_NS4_BEG2 ),
    .S(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame7_bit24.Q ),
    .X(_0134_));
 sky130_fd_sc_hd__a221o_1 _0502_ (.A1(_0132_),
    .A2(_0133_),
    .B1(_0134_),
    .B2(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame7_bit25.Q ),
    .C1(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame7_bit26.Q ),
    .X(_0135_));
 sky130_fd_sc_hd__o21a_1 _0503_ (.A1(_0016_),
    .A2(_0131_),
    .B1(_0135_),
    .X(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.S4BEG2 ));
 sky130_fd_sc_hd__mux4_1 _0504_ (.A0(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.J_NS4_BEG7 ),
    .A1(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.J_NS4_BEG11 ),
    .A2(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.J_NS4_BEG15 ),
    .A3(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.J_NS2_BEG7 ),
    .S0(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame7_bit27.Q ),
    .S1(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame7_bit28.Q ),
    .X(_0136_));
 sky130_fd_sc_hd__nand2b_1 _0505_ (.A_N(net71),
    .B(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame7_bit27.Q ),
    .Y(_0137_));
 sky130_fd_sc_hd__o21ba_1 _0506_ (.A1(net36),
    .A2(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame7_bit27.Q ),
    .B1_N(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame7_bit28.Q ),
    .X(_0138_));
 sky130_fd_sc_hd__mux2_1 _0507_ (.A0(net62),
    .A1(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.J_NS4_BEG3 ),
    .S(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame7_bit27.Q ),
    .X(_0139_));
 sky130_fd_sc_hd__a221o_1 _0508_ (.A1(_0137_),
    .A2(_0138_),
    .B1(_0139_),
    .B2(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame7_bit28.Q ),
    .C1(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame7_bit29.Q ),
    .X(_0140_));
 sky130_fd_sc_hd__o21a_1 _0509_ (.A1(_0017_),
    .A2(_0136_),
    .B1(_0140_),
    .X(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.S4BEG3 ));
 sky130_fd_sc_hd__mux4_2 _0510_ (.A0(net220),
    .A1(net240),
    .A2(_0087_),
    .A3(net137),
    .S0(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame0_bit0.Q ),
    .S1(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame0_bit1.Q ),
    .X(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.J_NS4_BEG12 ));
 sky130_fd_sc_hd__mux4_2 _0511_ (.A0(net221),
    .A1(net241),
    .A2(_0058_),
    .A3(net138),
    .S0(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame0_bit2.Q ),
    .S1(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame0_bit3.Q ),
    .X(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.J_NS4_BEG13 ));
 sky130_fd_sc_hd__mux4_2 _0512_ (.A0(net222),
    .A1(net242),
    .A2(_0065_),
    .A3(net139),
    .S0(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame0_bit4.Q ),
    .S1(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame0_bit5.Q ),
    .X(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.J_NS4_BEG14 ));
 sky130_fd_sc_hd__mux4_2 _0513_ (.A0(net223),
    .A1(net243),
    .A2(_0072_),
    .A3(net140),
    .S0(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame0_bit6.Q ),
    .S1(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame0_bit7.Q ),
    .X(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.J_NS4_BEG15 ));
 sky130_fd_sc_hd__mux4_1 _0514_ (.A0(net33),
    .A1(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.J_NS4_BEG12 ),
    .A2(net59),
    .A3(_0086_),
    .S0(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame9_bit23.Q ),
    .S1(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame9_bit22.Q ),
    .X(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.N1BEG0 ));
 sky130_fd_sc_hd__mux4_1 _0515_ (.A0(net141),
    .A1(net171),
    .A2(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.J_NS4_BEG12 ),
    .A3(_0090_),
    .S0(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame8_bit18.Q ),
    .S1(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame8_bit19.Q ),
    .X(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.S1BEG0 ));
 sky130_fd_sc_hd__mux4_1 _0516_ (.A0(net142),
    .A1(net172),
    .A2(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.J_NS4_BEG13 ),
    .A3(_0061_),
    .S0(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame8_bit20.Q ),
    .S1(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame8_bit21.Q ),
    .X(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.S1BEG1 ));
 sky130_fd_sc_hd__mux4_1 _0517_ (.A0(net143),
    .A1(net162),
    .A2(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.J_NS4_BEG14 ),
    .A3(_0068_),
    .S0(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame8_bit22.Q ),
    .S1(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame8_bit23.Q ),
    .X(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.S1BEG2 ));
 sky130_fd_sc_hd__mux4_1 _0518_ (.A0(net144),
    .A1(net163),
    .A2(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.J_NS4_BEG15 ),
    .A3(_0075_),
    .S0(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame8_bit24.Q ),
    .S1(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame8_bit25.Q ),
    .X(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.S1BEG3 ));
 sky130_fd_sc_hd__mux4_1 _0519_ (.A0(net160),
    .A1(net152),
    .A2(net171),
    .A3(_0076_),
    .S0(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame8_bit26.Q ),
    .S1(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame8_bit27.Q ),
    .X(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.S2BEG0 ));
 sky130_fd_sc_hd__mux4_1 _0520_ (.A0(net159),
    .A1(net151),
    .A2(net172),
    .A3(_0077_),
    .S0(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame8_bit28.Q ),
    .S1(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame8_bit29.Q ),
    .X(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.S2BEG1 ));
 sky130_fd_sc_hd__mux4_1 _0521_ (.A0(net158),
    .A1(net150),
    .A2(net162),
    .A3(_0078_),
    .S0(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame8_bit30.Q ),
    .S1(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame8_bit31.Q ),
    .X(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.S2BEG2 ));
 sky130_fd_sc_hd__mux4_1 _0522_ (.A0(net157),
    .A1(net149),
    .A2(net163),
    .A3(net366),
    .S0(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame7_bit0.Q ),
    .S1(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame7_bit1.Q ),
    .X(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.S2BEG3 ));
 sky130_fd_sc_hd__mux4_1 _0523_ (.A0(net141),
    .A1(net148),
    .A2(net156),
    .A3(net365),
    .S0(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame7_bit3.Q ),
    .S1(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame7_bit2.Q ),
    .X(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.S2BEG4 ));
 sky130_fd_sc_hd__mux4_1 _0524_ (.A0(net142),
    .A1(net147),
    .A2(net155),
    .A3(_0081_),
    .S0(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame7_bit5.Q ),
    .S1(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame7_bit4.Q ),
    .X(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.S2BEG5 ));
 sky130_fd_sc_hd__mux4_1 _0525_ (.A0(net143),
    .A1(net146),
    .A2(net154),
    .A3(_0082_),
    .S0(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame7_bit7.Q ),
    .S1(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame7_bit6.Q ),
    .X(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.S2BEG6 ));
 sky130_fd_sc_hd__mux4_1 _0526_ (.A0(net144),
    .A1(net145),
    .A2(net153),
    .A3(_0083_),
    .S0(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame7_bit9.Q ),
    .S1(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame7_bit8.Q ),
    .X(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.S2BEG7 ));
 sky130_fd_sc_hd__mux4_1 _0527_ (.A0(net220),
    .A1(net13),
    .A2(_0087_),
    .A3(net30),
    .S0(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame7_bit23.Q ),
    .S1(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame7_bit22.Q ),
    .X(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.W1BEG0 ));
 sky130_fd_sc_hd__mux4_1 _0528_ (.A0(net221),
    .A1(net24),
    .A2(_0058_),
    .A3(net29),
    .S0(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame7_bit25.Q ),
    .S1(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame7_bit24.Q ),
    .X(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.W1BEG1 ));
 sky130_fd_sc_hd__mux4_1 _0529_ (.A0(net222),
    .A1(net1),
    .A2(_0065_),
    .A3(net28),
    .S0(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame7_bit27.Q ),
    .S1(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame7_bit26.Q ),
    .X(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.W1BEG2 ));
 sky130_fd_sc_hd__mux4_1 _0530_ (.A0(net223),
    .A1(net2),
    .A2(_0072_),
    .A3(net27),
    .S0(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame7_bit29.Q ),
    .S1(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame7_bit28.Q ),
    .X(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.W1BEG3 ));
 sky130_fd_sc_hd__mux4_1 _0531_ (.A0(net1),
    .A1(net31),
    .A2(net369),
    .A3(_0083_),
    .S0(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame7_bit30.Q ),
    .S1(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame7_bit31.Q ),
    .X(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.W2BEG0 ));
 sky130_fd_sc_hd__mux4_1 _0532_ (.A0(net2),
    .A1(net32),
    .A2(net368),
    .A3(_0082_),
    .S0(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame6_bit0.Q ),
    .S1(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame6_bit1.Q ),
    .X(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.W2BEG1 ));
 sky130_fd_sc_hd__mux4_1 _0533_ (.A0(net13),
    .A1(net3),
    .A2(net367),
    .A3(_0081_),
    .S0(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame6_bit2.Q ),
    .S1(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame6_bit3.Q ),
    .X(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.W2BEG2 ));
 sky130_fd_sc_hd__mux4_1 _0534_ (.A0(net24),
    .A1(net4),
    .A2(net366),
    .A3(net365),
    .S0(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame6_bit4.Q ),
    .S1(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame6_bit5.Q ),
    .X(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.W2BEG3 ));
 sky130_fd_sc_hd__mux4_1 _0535_ (.A0(net27),
    .A1(net5),
    .A2(net366),
    .A3(net365),
    .S0(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame6_bit6.Q ),
    .S1(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame6_bit7.Q ),
    .X(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.W2BEG4 ));
 sky130_fd_sc_hd__mux4_1 _0536_ (.A0(net28),
    .A1(net6),
    .A2(net367),
    .A3(_0081_),
    .S0(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame6_bit8.Q ),
    .S1(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame6_bit9.Q ),
    .X(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.W2BEG5 ));
 sky130_fd_sc_hd__mux4_1 _0537_ (.A0(net29),
    .A1(net7),
    .A2(net368),
    .A3(_0082_),
    .S0(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame6_bit10.Q ),
    .S1(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame6_bit11.Q ),
    .X(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.W2BEG6 ));
 sky130_fd_sc_hd__mux4_1 _0538_ (.A0(net30),
    .A1(net8),
    .A2(net369),
    .A3(_0083_),
    .S0(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame6_bit12.Q ),
    .S1(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame6_bit13.Q ),
    .X(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.W2BEG7 ));
 sky130_fd_sc_hd__mux4_1 _0539_ (.A0(net1),
    .A1(net31),
    .A2(net369),
    .A3(_0083_),
    .S0(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame6_bit14.Q ),
    .S1(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame6_bit15.Q ),
    .X(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.W2BEGb0 ));
 sky130_fd_sc_hd__mux4_1 _0540_ (.A0(net2),
    .A1(net32),
    .A2(net368),
    .A3(_0082_),
    .S0(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame6_bit16.Q ),
    .S1(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame6_bit17.Q ),
    .X(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.W2BEGb1 ));
 sky130_fd_sc_hd__mux4_1 _0541_ (.A0(net13),
    .A1(net3),
    .A2(net367),
    .A3(_0081_),
    .S0(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame6_bit18.Q ),
    .S1(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame6_bit19.Q ),
    .X(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.W2BEGb2 ));
 sky130_fd_sc_hd__mux4_1 _0542_ (.A0(net24),
    .A1(net4),
    .A2(net366),
    .A3(net365),
    .S0(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame6_bit20.Q ),
    .S1(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame6_bit21.Q ),
    .X(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.W2BEGb3 ));
 sky130_fd_sc_hd__mux4_1 _0543_ (.A0(net27),
    .A1(net5),
    .A2(net366),
    .A3(net365),
    .S0(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame6_bit22.Q ),
    .S1(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame6_bit23.Q ),
    .X(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.W2BEGb4 ));
 sky130_fd_sc_hd__mux4_1 _0544_ (.A0(net28),
    .A1(net6),
    .A2(net367),
    .A3(_0081_),
    .S0(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame6_bit24.Q ),
    .S1(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame6_bit25.Q ),
    .X(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.W2BEGb5 ));
 sky130_fd_sc_hd__mux4_1 _0545_ (.A0(net29),
    .A1(net7),
    .A2(net368),
    .A3(_0082_),
    .S0(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame6_bit26.Q ),
    .S1(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame6_bit27.Q ),
    .X(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.W2BEGb6 ));
 sky130_fd_sc_hd__mux4_1 _0546_ (.A0(net30),
    .A1(net8),
    .A2(net369),
    .A3(_0083_),
    .S0(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame6_bit28.Q ),
    .S1(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame6_bit29.Q ),
    .X(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.W2BEGb7 ));
 sky130_fd_sc_hd__mux4_1 _0547_ (.A0(net1),
    .A1(net5),
    .A2(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.J_NS4_BEG15 ),
    .A3(_0083_),
    .S0(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame6_bit30.Q ),
    .S1(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame6_bit31.Q ),
    .X(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.WW4BEG0 ));
 sky130_fd_sc_hd__mux4_1 _0548_ (.A0(net2),
    .A1(net6),
    .A2(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.J_NS4_BEG14 ),
    .A3(_0082_),
    .S0(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame5_bit0.Q ),
    .S1(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame5_bit1.Q ),
    .X(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.WW4BEG1 ));
 sky130_fd_sc_hd__mux4_1 _0549_ (.A0(net13),
    .A1(net7),
    .A2(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.J_NS4_BEG13 ),
    .A3(_0081_),
    .S0(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame5_bit2.Q ),
    .S1(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame5_bit3.Q ),
    .X(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.WW4BEG2 ));
 sky130_fd_sc_hd__mux4_1 _0550_ (.A0(net24),
    .A1(net8),
    .A2(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.J_NS4_BEG12 ),
    .A3(net365),
    .S0(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame5_bit4.Q ),
    .S1(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame5_bit5.Q ),
    .X(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.WW4BEG3 ));
 sky130_fd_sc_hd__mux4_2 _0551_ (.A0(net223),
    .A1(net243),
    .A2(_0072_),
    .A3(net140),
    .S0(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame1_bit30.Q ),
    .S1(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame1_bit31.Q ),
    .X(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.J_NS4_BEG11 ));
 sky130_fd_sc_hd__mux4_1 _0552_ (.A0(net27),
    .A1(net31),
    .A2(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.J_NS4_BEG11 ),
    .A3(net366),
    .S0(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame5_bit6.Q ),
    .S1(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame5_bit7.Q ),
    .X(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.WW4BEG4 ));
 sky130_fd_sc_hd__mux4_2 _0553_ (.A0(net222),
    .A1(net242),
    .A2(_0065_),
    .A3(net139),
    .S0(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame1_bit28.Q ),
    .S1(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame1_bit29.Q ),
    .X(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.J_NS4_BEG10 ));
 sky130_fd_sc_hd__mux4_1 _0554_ (.A0(net28),
    .A1(net32),
    .A2(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.J_NS4_BEG10 ),
    .A3(net367),
    .S0(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame5_bit8.Q ),
    .S1(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame5_bit9.Q ),
    .X(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.WW4BEG5 ));
 sky130_fd_sc_hd__mux4_2 _0555_ (.A0(net221),
    .A1(net241),
    .A2(_0058_),
    .A3(net138),
    .S0(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame1_bit26.Q ),
    .S1(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame1_bit27.Q ),
    .X(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.J_NS4_BEG9 ));
 sky130_fd_sc_hd__mux4_1 _0556_ (.A0(net29),
    .A1(net3),
    .A2(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.J_NS4_BEG9 ),
    .A3(net368),
    .S0(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame5_bit10.Q ),
    .S1(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame5_bit11.Q ),
    .X(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.WW4BEG6 ));
 sky130_fd_sc_hd__mux4_2 _0557_ (.A0(net220),
    .A1(net240),
    .A2(_0087_),
    .A3(net137),
    .S0(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame1_bit24.Q ),
    .S1(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame1_bit25.Q ),
    .X(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.J_NS4_BEG8 ));
 sky130_fd_sc_hd__mux4_1 _0558_ (.A0(net30),
    .A1(net4),
    .A2(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.J_NS4_BEG8 ),
    .A3(net369),
    .S0(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame5_bit12.Q ),
    .S1(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame5_bit13.Q ),
    .X(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.WW4BEG7 ));
 sky130_fd_sc_hd__mux4_2 _0559_ (.A0(net223),
    .A1(net243),
    .A2(_0072_),
    .A3(net140),
    .S0(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame1_bit22.Q ),
    .S1(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame1_bit23.Q ),
    .X(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.J_NS4_BEG7 ));
 sky130_fd_sc_hd__mux4_1 _0560_ (.A0(net27),
    .A1(net31),
    .A2(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.J_NS4_BEG7 ),
    .A3(_0083_),
    .S0(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame5_bit14.Q ),
    .S1(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame5_bit15.Q ),
    .X(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.WW4BEG8 ));
 sky130_fd_sc_hd__mux4_2 _0561_ (.A0(net222),
    .A1(net242),
    .A2(_0065_),
    .A3(net139),
    .S0(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame1_bit20.Q ),
    .S1(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame1_bit21.Q ),
    .X(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.J_NS4_BEG6 ));
 sky130_fd_sc_hd__mux4_1 _0562_ (.A0(net28),
    .A1(net32),
    .A2(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.J_NS4_BEG6 ),
    .A3(_0082_),
    .S0(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame5_bit16.Q ),
    .S1(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame5_bit17.Q ),
    .X(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.WW4BEG9 ));
 sky130_fd_sc_hd__mux4_2 _0563_ (.A0(net221),
    .A1(net241),
    .A2(_0058_),
    .A3(net138),
    .S0(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame1_bit18.Q ),
    .S1(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame1_bit19.Q ),
    .X(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.J_NS4_BEG5 ));
 sky130_fd_sc_hd__mux4_1 _0564_ (.A0(net29),
    .A1(net3),
    .A2(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.J_NS4_BEG5 ),
    .A3(_0081_),
    .S0(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame5_bit18.Q ),
    .S1(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame5_bit19.Q ),
    .X(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.WW4BEG10 ));
 sky130_fd_sc_hd__mux4_2 _0565_ (.A0(net220),
    .A1(net240),
    .A2(_0087_),
    .A3(net137),
    .S0(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame1_bit16.Q ),
    .S1(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame1_bit17.Q ),
    .X(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.J_NS4_BEG4 ));
 sky130_fd_sc_hd__mux4_1 _0566_ (.A0(net30),
    .A1(net4),
    .A2(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.J_NS4_BEG4 ),
    .A3(net365),
    .S0(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame5_bit20.Q ),
    .S1(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame5_bit21.Q ),
    .X(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.WW4BEG11 ));
 sky130_fd_sc_hd__mux4_2 _0567_ (.A0(net223),
    .A1(net243),
    .A2(_0072_),
    .A3(net140),
    .S0(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame1_bit14.Q ),
    .S1(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame1_bit15.Q ),
    .X(_0141_));
 sky130_fd_sc_hd__mux4_1 _0568_ (.A0(net1),
    .A1(net5),
    .A2(_0141_),
    .A3(net366),
    .S0(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame5_bit22.Q ),
    .S1(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame5_bit23.Q ),
    .X(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.WW4BEG12 ));
 sky130_fd_sc_hd__mux4_2 _0569_ (.A0(net222),
    .A1(net242),
    .A2(_0065_),
    .A3(net139),
    .S0(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame1_bit12.Q ),
    .S1(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame1_bit13.Q ),
    .X(_0142_));
 sky130_fd_sc_hd__mux4_1 _0570_ (.A0(net2),
    .A1(net6),
    .A2(_0142_),
    .A3(net367),
    .S0(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame5_bit24.Q ),
    .S1(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame5_bit25.Q ),
    .X(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.WW4BEG13 ));
 sky130_fd_sc_hd__mux4_2 _0571_ (.A0(net221),
    .A1(net241),
    .A2(_0058_),
    .A3(net138),
    .S0(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame1_bit10.Q ),
    .S1(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame1_bit11.Q ),
    .X(_0143_));
 sky130_fd_sc_hd__mux4_1 _0572_ (.A0(net13),
    .A1(net7),
    .A2(_0143_),
    .A3(net368),
    .S0(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame5_bit26.Q ),
    .S1(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame5_bit27.Q ),
    .X(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.WW4BEG14 ));
 sky130_fd_sc_hd__mux4_2 _0573_ (.A0(net220),
    .A1(net240),
    .A2(_0087_),
    .A3(net137),
    .S0(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame1_bit8.Q ),
    .S1(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame1_bit9.Q ),
    .X(_0144_));
 sky130_fd_sc_hd__mux4_1 _0574_ (.A0(net24),
    .A1(net8),
    .A2(_0144_),
    .A3(net369),
    .S0(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame5_bit28.Q ),
    .S1(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame5_bit29.Q ),
    .X(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.WW4BEG15 ));
 sky130_fd_sc_hd__mux4_1 _0575_ (.A0(net240),
    .A1(net137),
    .A2(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.J_NS4_BEG11 ),
    .A3(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.J_NS4_BEG15 ),
    .S0(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame5_bit30.Q ),
    .S1(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame5_bit31.Q ),
    .X(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.W6BEG0 ));
 sky130_fd_sc_hd__mux4_1 _0576_ (.A0(net241),
    .A1(net138),
    .A2(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.J_NS4_BEG10 ),
    .A3(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.J_NS4_BEG14 ),
    .S0(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame4_bit0.Q ),
    .S1(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame4_bit1.Q ),
    .X(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.W6BEG1 ));
 sky130_fd_sc_hd__mux4_1 _0577_ (.A0(net242),
    .A1(net139),
    .A2(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.J_NS4_BEG9 ),
    .A3(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.J_NS4_BEG13 ),
    .S0(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame4_bit2.Q ),
    .S1(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame4_bit3.Q ),
    .X(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.W6BEG2 ));
 sky130_fd_sc_hd__mux4_1 _0578_ (.A0(net243),
    .A1(net140),
    .A2(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.J_NS4_BEG8 ),
    .A3(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.J_NS4_BEG12 ),
    .S0(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame4_bit4.Q ),
    .S1(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame4_bit5.Q ),
    .X(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.W6BEG3 ));
 sky130_fd_sc_hd__mux4_1 _0579_ (.A0(net27),
    .A1(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.J_NS4_BEG11 ),
    .A2(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.J_NS4_BEG7 ),
    .A3(net369),
    .S0(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame4_bit7.Q ),
    .S1(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame4_bit6.Q ),
    .X(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.W6BEG4 ));
 sky130_fd_sc_hd__mux4_1 _0580_ (.A0(net28),
    .A1(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.J_NS4_BEG10 ),
    .A2(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.J_NS4_BEG6 ),
    .A3(net368),
    .S0(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame4_bit9.Q ),
    .S1(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame4_bit8.Q ),
    .X(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.W6BEG5 ));
 sky130_fd_sc_hd__mux4_1 _0581_ (.A0(net29),
    .A1(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.J_NS4_BEG5 ),
    .A2(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.J_NS4_BEG9 ),
    .A3(net367),
    .S0(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame4_bit10.Q ),
    .S1(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame4_bit11.Q ),
    .X(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.W6BEG6 ));
 sky130_fd_sc_hd__mux4_1 _0582_ (.A0(net30),
    .A1(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.J_NS4_BEG4 ),
    .A2(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.J_NS4_BEG8 ),
    .A3(net366),
    .S0(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame4_bit12.Q ),
    .S1(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame4_bit13.Q ),
    .X(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.W6BEG7 ));
 sky130_fd_sc_hd__mux4_1 _0583_ (.A0(net1),
    .A1(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.J_NS4_BEG7 ),
    .A2(_0141_),
    .A3(net365),
    .S0(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame4_bit15.Q ),
    .S1(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame4_bit14.Q ),
    .X(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.W6BEG8 ));
 sky130_fd_sc_hd__mux4_1 _0584_ (.A0(net2),
    .A1(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.J_NS4_BEG6 ),
    .A2(_0142_),
    .A3(_0081_),
    .S0(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame4_bit17.Q ),
    .S1(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame4_bit16.Q ),
    .X(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.W6BEG9 ));
 sky130_fd_sc_hd__mux4_1 _0585_ (.A0(net13),
    .A1(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.J_NS4_BEG5 ),
    .A2(_0143_),
    .A3(_0082_),
    .S0(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame4_bit19.Q ),
    .S1(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame4_bit18.Q ),
    .X(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.W6BEG10 ));
 sky130_fd_sc_hd__mux4_1 _0586_ (.A0(net24),
    .A1(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.J_NS4_BEG4 ),
    .A2(_0144_),
    .A3(_0083_),
    .S0(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame4_bit21.Q ),
    .S1(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame4_bit20.Q ),
    .X(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.W6BEG11 ));
 sky130_fd_sc_hd__o21ba_1 _0587_ (.A1(net153),
    .A2(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame4_bit22.Q ),
    .B1_N(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame4_bit23.Q ),
    .X(_0145_));
 sky130_fd_sc_hd__o21a_1 _0588_ (.A1(net145),
    .A2(_0023_),
    .B1(_0145_),
    .X(_0146_));
 sky130_fd_sc_hd__a31o_1 _0589_ (.A1(_0023_),
    .A2(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame4_bit23.Q ),
    .A3(net369),
    .B1(_0146_),
    .X(net248));
 sky130_fd_sc_hd__o21ba_1 _0590_ (.A1(net154),
    .A2(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame4_bit24.Q ),
    .B1_N(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame4_bit25.Q ),
    .X(_0147_));
 sky130_fd_sc_hd__o21a_1 _0591_ (.A1(net146),
    .A2(_0024_),
    .B1(_0147_),
    .X(_0148_));
 sky130_fd_sc_hd__a31o_1 _0592_ (.A1(_0024_),
    .A2(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame4_bit25.Q ),
    .A3(net368),
    .B1(_0148_),
    .X(net249));
 sky130_fd_sc_hd__o21ba_1 _0593_ (.A1(net155),
    .A2(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame4_bit26.Q ),
    .B1_N(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame4_bit27.Q ),
    .X(_0149_));
 sky130_fd_sc_hd__o21a_1 _0594_ (.A1(net147),
    .A2(_0025_),
    .B1(_0149_),
    .X(_0150_));
 sky130_fd_sc_hd__a31o_1 _0595_ (.A1(_0025_),
    .A2(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame4_bit27.Q ),
    .A3(net367),
    .B1(_0150_),
    .X(net250));
 sky130_fd_sc_hd__o21ba_1 _0596_ (.A1(net156),
    .A2(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame4_bit28.Q ),
    .B1_N(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame4_bit29.Q ),
    .X(_0151_));
 sky130_fd_sc_hd__o21a_1 _0597_ (.A1(net148),
    .A2(_0026_),
    .B1(_0151_),
    .X(_0152_));
 sky130_fd_sc_hd__a31o_1 _0598_ (.A1(_0026_),
    .A2(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame4_bit29.Q ),
    .A3(net366),
    .B1(_0152_),
    .X(net251));
 sky130_fd_sc_hd__o21ba_1 _0599_ (.A1(net157),
    .A2(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame4_bit30.Q ),
    .B1_N(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame4_bit31.Q ),
    .X(_0153_));
 sky130_fd_sc_hd__o21a_1 _0600_ (.A1(net149),
    .A2(_0027_),
    .B1(_0153_),
    .X(_0154_));
 sky130_fd_sc_hd__a31o_1 _0601_ (.A1(_0027_),
    .A2(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame4_bit31.Q ),
    .A3(net365),
    .B1(_0154_),
    .X(net252));
 sky130_fd_sc_hd__mux4_1 _0602_ (.A0(net173),
    .A1(net187),
    .A2(net161),
    .A3(_0144_),
    .S0(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame3_bit0.Q ),
    .S1(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame3_bit1.Q ),
    .X(net258));
 sky130_fd_sc_hd__mux4_2 _0603_ (.A0(net180),
    .A1(net188),
    .A2(net164),
    .A3(_0143_),
    .S0(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame3_bit2.Q ),
    .S1(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame3_bit3.Q ),
    .X(net259));
 sky130_fd_sc_hd__mux4_2 _0604_ (.A0(net181),
    .A1(net174),
    .A2(net165),
    .A3(_0142_),
    .S0(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame3_bit4.Q ),
    .S1(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame3_bit5.Q ),
    .X(net270));
 sky130_fd_sc_hd__mux4_1 _0605_ (.A0(net182),
    .A1(net175),
    .A2(net166),
    .A3(_0141_),
    .S0(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame3_bit6.Q ),
    .S1(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame3_bit7.Q ),
    .X(net281));
 sky130_fd_sc_hd__mux4_1 _0606_ (.A0(net183),
    .A1(net176),
    .A2(net167),
    .A3(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.J_NS4_BEG4 ),
    .S0(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame3_bit8.Q ),
    .S1(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame3_bit9.Q ),
    .X(net284));
 sky130_fd_sc_hd__mux4_2 _0607_ (.A0(net184),
    .A1(net177),
    .A2(net168),
    .A3(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.J_NS4_BEG5 ),
    .S0(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame3_bit10.Q ),
    .S1(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame3_bit11.Q ),
    .X(net285));
 sky130_fd_sc_hd__mux4_2 _0608_ (.A0(net185),
    .A1(net178),
    .A2(net169),
    .A3(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.J_NS4_BEG6 ),
    .S0(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame3_bit12.Q ),
    .S1(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame3_bit13.Q ),
    .X(net286));
 sky130_fd_sc_hd__mux4_1 _0609_ (.A0(net186),
    .A1(net179),
    .A2(net170),
    .A3(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.J_NS4_BEG7 ),
    .S0(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame3_bit14.Q ),
    .S1(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame3_bit15.Q ),
    .X(net287));
 sky130_fd_sc_hd__mux4_1 _0610_ (.A0(net173),
    .A1(net187),
    .A2(net171),
    .A3(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.J_NS4_BEG8 ),
    .S0(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame3_bit16.Q ),
    .S1(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame3_bit17.Q ),
    .X(net288));
 sky130_fd_sc_hd__mux4_2 _0611_ (.A0(net180),
    .A1(net188),
    .A2(net172),
    .A3(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.J_NS4_BEG9 ),
    .S0(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame3_bit18.Q ),
    .S1(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame3_bit19.Q ),
    .X(net289));
 sky130_fd_sc_hd__mux4_2 _0612_ (.A0(net181),
    .A1(net174),
    .A2(net162),
    .A3(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.J_NS4_BEG10 ),
    .S0(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame3_bit20.Q ),
    .S1(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame3_bit21.Q ),
    .X(net260));
 sky130_fd_sc_hd__mux4_1 _0613_ (.A0(net182),
    .A1(net175),
    .A2(net163),
    .A3(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.J_NS4_BEG11 ),
    .S0(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame3_bit22.Q ),
    .S1(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame3_bit23.Q ),
    .X(net261));
 sky130_fd_sc_hd__mux4_1 _0614_ (.A0(net141),
    .A1(net183),
    .A2(net176),
    .A3(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.J_NS4_BEG12 ),
    .S0(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame3_bit24.Q ),
    .S1(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame3_bit25.Q ),
    .X(net262));
 sky130_fd_sc_hd__mux4_2 _0615_ (.A0(net142),
    .A1(net184),
    .A2(net177),
    .A3(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.J_NS4_BEG13 ),
    .S0(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame3_bit26.Q ),
    .S1(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame3_bit27.Q ),
    .X(net263));
 sky130_fd_sc_hd__mux4_2 _0616_ (.A0(net143),
    .A1(net185),
    .A2(net178),
    .A3(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.J_NS4_BEG14 ),
    .S0(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame3_bit28.Q ),
    .S1(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame3_bit29.Q ),
    .X(net264));
 sky130_fd_sc_hd__mux4_1 _0617_ (.A0(net144),
    .A1(net186),
    .A2(net179),
    .A3(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.J_NS4_BEG15 ),
    .S0(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame3_bit30.Q ),
    .S1(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame3_bit31.Q ),
    .X(net265));
 sky130_fd_sc_hd__mux4_1 _0618_ (.A0(net173),
    .A1(net187),
    .A2(net161),
    .A3(_0144_),
    .S0(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame2_bit0.Q ),
    .S1(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame2_bit1.Q ),
    .X(net291));
 sky130_fd_sc_hd__mux4_2 _0619_ (.A0(net180),
    .A1(net188),
    .A2(net164),
    .A3(_0143_),
    .S0(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame2_bit2.Q ),
    .S1(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame2_bit3.Q ),
    .X(net292));
 sky130_fd_sc_hd__mux4_2 _0620_ (.A0(net181),
    .A1(net174),
    .A2(net165),
    .A3(_0142_),
    .S0(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame2_bit4.Q ),
    .S1(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame2_bit5.Q ),
    .X(net303));
 sky130_fd_sc_hd__mux4_2 _0621_ (.A0(net182),
    .A1(net175),
    .A2(net166),
    .A3(_0141_),
    .S0(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame2_bit6.Q ),
    .S1(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame2_bit7.Q ),
    .X(net314));
 sky130_fd_sc_hd__mux4_1 _0622_ (.A0(net183),
    .A1(net176),
    .A2(net167),
    .A3(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.J_NS4_BEG4 ),
    .S0(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame2_bit8.Q ),
    .S1(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame2_bit9.Q ),
    .X(net317));
 sky130_fd_sc_hd__mux4_2 _0623_ (.A0(net184),
    .A1(net177),
    .A2(net168),
    .A3(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.J_NS4_BEG5 ),
    .S0(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame2_bit10.Q ),
    .S1(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame2_bit11.Q ),
    .X(net318));
 sky130_fd_sc_hd__mux4_2 _0624_ (.A0(net185),
    .A1(net178),
    .A2(net169),
    .A3(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.J_NS4_BEG6 ),
    .S0(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame2_bit12.Q ),
    .S1(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame2_bit13.Q ),
    .X(net319));
 sky130_fd_sc_hd__mux4_2 _0625_ (.A0(net186),
    .A1(net179),
    .A2(net170),
    .A3(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.J_NS4_BEG7 ),
    .S0(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame2_bit14.Q ),
    .S1(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame2_bit15.Q ),
    .X(net320));
 sky130_fd_sc_hd__mux4_1 _0626_ (.A0(net173),
    .A1(net187),
    .A2(net171),
    .A3(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.J_NS4_BEG8 ),
    .S0(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame2_bit16.Q ),
    .S1(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame2_bit17.Q ),
    .X(net321));
 sky130_fd_sc_hd__mux4_2 _0627_ (.A0(net180),
    .A1(net188),
    .A2(net172),
    .A3(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.J_NS4_BEG9 ),
    .S0(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame2_bit18.Q ),
    .S1(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame2_bit19.Q ),
    .X(net322));
 sky130_fd_sc_hd__mux4_2 _0628_ (.A0(net181),
    .A1(net174),
    .A2(net162),
    .A3(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.J_NS4_BEG10 ),
    .S0(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame2_bit20.Q ),
    .S1(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame2_bit21.Q ),
    .X(net293));
 sky130_fd_sc_hd__mux4_2 _0629_ (.A0(net182),
    .A1(net175),
    .A2(net163),
    .A3(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.J_NS4_BEG11 ),
    .S0(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame2_bit22.Q ),
    .S1(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame2_bit23.Q ),
    .X(net294));
 sky130_fd_sc_hd__mux4_1 _0630_ (.A0(net141),
    .A1(net183),
    .A2(net176),
    .A3(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.J_NS4_BEG12 ),
    .S0(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame2_bit24.Q ),
    .S1(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame2_bit25.Q ),
    .X(net295));
 sky130_fd_sc_hd__mux4_2 _0631_ (.A0(net142),
    .A1(net184),
    .A2(net177),
    .A3(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.J_NS4_BEG13 ),
    .S0(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame2_bit26.Q ),
    .S1(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame2_bit27.Q ),
    .X(net296));
 sky130_fd_sc_hd__mux4_2 _0632_ (.A0(net143),
    .A1(net185),
    .A2(net178),
    .A3(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.J_NS4_BEG14 ),
    .S0(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame2_bit28.Q ),
    .S1(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame2_bit29.Q ),
    .X(net297));
 sky130_fd_sc_hd__mux4_2 _0633_ (.A0(net144),
    .A1(net186),
    .A2(net179),
    .A3(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.J_NS4_BEG15 ),
    .S0(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame2_bit30.Q ),
    .S1(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame2_bit31.Q ),
    .X(net298));
 sky130_fd_sc_hd__or2_1 _0634_ (.A(net171),
    .B(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame8_bit6.Q ),
    .X(_0155_));
 sky130_fd_sc_hd__o211a_1 _0635_ (.A1(_0028_),
    .A2(_0144_),
    .B1(_0155_),
    .C1(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame8_bit7.Q ),
    .X(_0156_));
 sky130_fd_sc_hd__mux2_1 _0636_ (.A0(net141),
    .A1(net173),
    .S(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame8_bit6.Q ),
    .X(_0157_));
 sky130_fd_sc_hd__a21o_1 _0637_ (.A1(_0029_),
    .A2(_0157_),
    .B1(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame8_bit8.Q ),
    .X(_0158_));
 sky130_fd_sc_hd__mux4_1 _0638_ (.A0(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.J_NS4_BEG12 ),
    .A1(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.J_NS4_BEG4 ),
    .A2(net369),
    .A3(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.J_NS4_BEG8 ),
    .S0(_0029_),
    .S1(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame8_bit6.Q ),
    .X(_0159_));
 sky130_fd_sc_hd__o22a_1 _0639_ (.A1(_0156_),
    .A2(_0158_),
    .B1(_0159_),
    .B2(_0030_),
    .X(\Tile_X0Y0_EF_SRAM_top.N4BEG_outbuf_8.A ));
 sky130_fd_sc_hd__or2_1 _0640_ (.A(net172),
    .B(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame8_bit9.Q ),
    .X(_0160_));
 sky130_fd_sc_hd__o211a_1 _0641_ (.A1(_0031_),
    .A2(_0143_),
    .B1(_0160_),
    .C1(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame8_bit10.Q ),
    .X(_0161_));
 sky130_fd_sc_hd__mux2_1 _0642_ (.A0(net142),
    .A1(net180),
    .S(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame8_bit9.Q ),
    .X(_0162_));
 sky130_fd_sc_hd__a21o_1 _0643_ (.A1(_0032_),
    .A2(_0162_),
    .B1(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame8_bit11.Q ),
    .X(_0163_));
 sky130_fd_sc_hd__mux4_1 _0644_ (.A0(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.J_NS4_BEG13 ),
    .A1(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.J_NS4_BEG5 ),
    .A2(net368),
    .A3(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.J_NS4_BEG9 ),
    .S0(_0032_),
    .S1(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame8_bit9.Q ),
    .X(_0164_));
 sky130_fd_sc_hd__o22a_1 _0645_ (.A1(_0161_),
    .A2(_0163_),
    .B1(_0164_),
    .B2(_0033_),
    .X(\Tile_X0Y0_EF_SRAM_top.N4BEG_outbuf_9.A ));
 sky130_fd_sc_hd__or2_1 _0646_ (.A(net162),
    .B(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame8_bit12.Q ),
    .X(_0165_));
 sky130_fd_sc_hd__o211a_1 _0647_ (.A1(_0034_),
    .A2(_0142_),
    .B1(_0165_),
    .C1(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame8_bit13.Q ),
    .X(_0166_));
 sky130_fd_sc_hd__mux2_1 _0648_ (.A0(net143),
    .A1(net181),
    .S(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame8_bit12.Q ),
    .X(_0167_));
 sky130_fd_sc_hd__a21o_1 _0649_ (.A1(_0035_),
    .A2(_0167_),
    .B1(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame8_bit14.Q ),
    .X(_0168_));
 sky130_fd_sc_hd__mux4_1 _0650_ (.A0(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.J_NS4_BEG14 ),
    .A1(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.J_NS4_BEG6 ),
    .A2(net367),
    .A3(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.J_NS4_BEG10 ),
    .S0(_0035_),
    .S1(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame8_bit12.Q ),
    .X(_0169_));
 sky130_fd_sc_hd__o22a_1 _0651_ (.A1(_0166_),
    .A2(_0168_),
    .B1(_0169_),
    .B2(_0036_),
    .X(\Tile_X0Y0_EF_SRAM_top.N4BEG_outbuf_10.A ));
 sky130_fd_sc_hd__or2_1 _0652_ (.A(net163),
    .B(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame8_bit15.Q ),
    .X(_0170_));
 sky130_fd_sc_hd__o211a_1 _0653_ (.A1(_0037_),
    .A2(_0141_),
    .B1(_0170_),
    .C1(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame8_bit16.Q ),
    .X(_0171_));
 sky130_fd_sc_hd__mux2_1 _0654_ (.A0(net144),
    .A1(net182),
    .S(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame8_bit15.Q ),
    .X(_0172_));
 sky130_fd_sc_hd__a21o_1 _0655_ (.A1(_0038_),
    .A2(_0172_),
    .B1(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame8_bit17.Q ),
    .X(_0173_));
 sky130_fd_sc_hd__mux4_1 _0656_ (.A0(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.J_NS4_BEG15 ),
    .A1(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.J_NS4_BEG7 ),
    .A2(net366),
    .A3(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.J_NS4_BEG11 ),
    .S0(_0038_),
    .S1(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame8_bit15.Q ),
    .X(_0174_));
 sky130_fd_sc_hd__o22a_1 _0657_ (.A1(_0171_),
    .A2(_0173_),
    .B1(_0174_),
    .B2(_0039_),
    .X(\Tile_X0Y0_EF_SRAM_top.N4BEG_outbuf_11.A ));
 sky130_fd_sc_hd__or2_1 _0658_ (.A(net167),
    .B(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame7_bit10.Q ),
    .X(_0175_));
 sky130_fd_sc_hd__o211a_1 _0659_ (.A1(_0040_),
    .A2(_0144_),
    .B1(_0175_),
    .C1(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame7_bit11.Q ),
    .X(_0176_));
 sky130_fd_sc_hd__mux2_1 _0660_ (.A0(net141),
    .A1(net176),
    .S(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame7_bit10.Q ),
    .X(_0177_));
 sky130_fd_sc_hd__a21o_1 _0661_ (.A1(_0041_),
    .A2(_0177_),
    .B1(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame7_bit12.Q ),
    .X(_0178_));
 sky130_fd_sc_hd__mux4_1 _0662_ (.A0(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.J_NS4_BEG12 ),
    .A1(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.J_NS4_BEG4 ),
    .A2(net365),
    .A3(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.J_NS4_BEG8 ),
    .S0(_0041_),
    .S1(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame7_bit10.Q ),
    .X(_0179_));
 sky130_fd_sc_hd__o22a_1 _0663_ (.A1(_0176_),
    .A2(_0178_),
    .B1(_0179_),
    .B2(_0042_),
    .X(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.S4BEG0 ));
 sky130_fd_sc_hd__or2_1 _0664_ (.A(net168),
    .B(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame7_bit13.Q ),
    .X(_0180_));
 sky130_fd_sc_hd__o211a_1 _0665_ (.A1(_0043_),
    .A2(_0143_),
    .B1(_0180_),
    .C1(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame7_bit14.Q ),
    .X(_0181_));
 sky130_fd_sc_hd__mux2_1 _0666_ (.A0(net142),
    .A1(net177),
    .S(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame7_bit13.Q ),
    .X(_0182_));
 sky130_fd_sc_hd__a21o_1 _0667_ (.A1(_0044_),
    .A2(_0182_),
    .B1(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame7_bit15.Q ),
    .X(_0183_));
 sky130_fd_sc_hd__mux4_1 _0668_ (.A0(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.J_NS4_BEG13 ),
    .A1(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.J_NS4_BEG5 ),
    .A2(_0081_),
    .A3(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.J_NS4_BEG9 ),
    .S0(_0044_),
    .S1(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame7_bit13.Q ),
    .X(_0184_));
 sky130_fd_sc_hd__o22a_1 _0669_ (.A1(_0181_),
    .A2(_0183_),
    .B1(_0184_),
    .B2(_0045_),
    .X(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.S4BEG1 ));
 sky130_fd_sc_hd__or2_1 _0670_ (.A(net169),
    .B(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame7_bit16.Q ),
    .X(_0185_));
 sky130_fd_sc_hd__o211a_1 _0671_ (.A1(_0046_),
    .A2(_0142_),
    .B1(_0185_),
    .C1(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame7_bit17.Q ),
    .X(_0186_));
 sky130_fd_sc_hd__mux2_1 _0672_ (.A0(net143),
    .A1(net178),
    .S(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame7_bit16.Q ),
    .X(_0187_));
 sky130_fd_sc_hd__a21o_1 _0673_ (.A1(_0047_),
    .A2(_0187_),
    .B1(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame7_bit18.Q ),
    .X(_0188_));
 sky130_fd_sc_hd__mux4_1 _0674_ (.A0(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.J_NS4_BEG14 ),
    .A1(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.J_NS4_BEG6 ),
    .A2(_0082_),
    .A3(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.J_NS4_BEG10 ),
    .S0(_0047_),
    .S1(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame7_bit16.Q ),
    .X(_0189_));
 sky130_fd_sc_hd__o22a_1 _0675_ (.A1(_0186_),
    .A2(_0188_),
    .B1(_0189_),
    .B2(_0048_),
    .X(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.S4BEG2 ));
 sky130_fd_sc_hd__or2_1 _0676_ (.A(net170),
    .B(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame7_bit19.Q ),
    .X(_0190_));
 sky130_fd_sc_hd__o211a_1 _0677_ (.A1(_0049_),
    .A2(_0141_),
    .B1(_0190_),
    .C1(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame7_bit20.Q ),
    .X(_0191_));
 sky130_fd_sc_hd__mux2_1 _0678_ (.A0(net144),
    .A1(net179),
    .S(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame7_bit19.Q ),
    .X(_0192_));
 sky130_fd_sc_hd__a21o_1 _0679_ (.A1(_0050_),
    .A2(_0192_),
    .B1(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame7_bit21.Q ),
    .X(_0193_));
 sky130_fd_sc_hd__mux4_1 _0680_ (.A0(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.J_NS4_BEG15 ),
    .A1(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.J_NS4_BEG7 ),
    .A2(_0083_),
    .A3(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.J_NS4_BEG11 ),
    .S0(_0050_),
    .S1(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame7_bit19.Q ),
    .X(_0194_));
 sky130_fd_sc_hd__o22a_1 _0681_ (.A1(_0191_),
    .A2(_0193_),
    .B1(_0194_),
    .B2(_0051_),
    .X(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.S4BEG3 ));
 sky130_fd_sc_hd__or3b_1 _0682_ (.A(net128),
    .B(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame1_bit1.Q ),
    .C_N(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame1_bit2.Q ),
    .X(_0195_));
 sky130_fd_sc_hd__o311a_1 _0683_ (.A1(net149),
    .A2(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame1_bit1.Q ),
    .A3(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame1_bit2.Q ),
    .B1(_0195_),
    .C1(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame1_bit0.Q ),
    .X(_0196_));
 sky130_fd_sc_hd__o31a_1 _0684_ (.A1(_0052_),
    .A2(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame1_bit2.Q ),
    .A3(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.S2BEG0 ),
    .B1(_0196_),
    .X(_0197_));
 sky130_fd_sc_hd__or3_1 _0685_ (.A(net148),
    .B(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame1_bit1.Q ),
    .C(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame1_bit2.Q ),
    .X(_0198_));
 sky130_fd_sc_hd__o21ai_1 _0686_ (.A1(_0008_),
    .A2(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame1_bit2.Q ),
    .B1(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame1_bit1.Q ),
    .Y(_0199_));
 sky130_fd_sc_hd__a21oi_1 _0687_ (.A1(_0009_),
    .A2(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame1_bit2.Q ),
    .B1(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame1_bit0.Q ),
    .Y(_0200_));
 sky130_fd_sc_hd__a31o_1 _0688_ (.A1(_0198_),
    .A2(_0199_),
    .A3(_0200_),
    .B1(_0197_),
    .X(_0201_));
 sky130_fd_sc_hd__mux2_1 _0689_ (.A0(net156),
    .A1(net159),
    .S(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame1_bit0.Q ),
    .X(_0202_));
 sky130_fd_sc_hd__or3b_1 _0690_ (.A(_0202_),
    .B(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame1_bit1.Q ),
    .C_N(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame1_bit2.Q ),
    .X(_0203_));
 sky130_fd_sc_hd__mux2_1 _0691_ (.A0(net238),
    .A1(net226),
    .S(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame1_bit0.Q ),
    .X(_0204_));
 sky130_fd_sc_hd__or3_1 _0692_ (.A(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame1_bit1.Q ),
    .B(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame1_bit2.Q ),
    .C(_0204_),
    .X(_0205_));
 sky130_fd_sc_hd__mux4_1 _0693_ (.A0(net227),
    .A1(net146),
    .A2(net153),
    .A3(net147),
    .S0(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame1_bit2.Q ),
    .S1(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame1_bit0.Q ),
    .X(_0206_));
 sky130_fd_sc_hd__o21ba_1 _0694_ (.A1(_0052_),
    .A2(_0206_),
    .B1_N(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame1_bit3.Q ),
    .X(_0207_));
 sky130_fd_sc_hd__a32o_1 _0695_ (.A1(_0203_),
    .A2(_0205_),
    .A3(_0207_),
    .B1(_0201_),
    .B2(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame1_bit3.Q ),
    .X(net323));
 sky130_fd_sc_hd__or3_1 _0696_ (.A(_0054_),
    .B(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame1_bit6.Q ),
    .C(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.S2BEG0 ),
    .X(_0208_));
 sky130_fd_sc_hd__mux2_1 _0697_ (.A0(net149),
    .A1(net128),
    .S(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame1_bit6.Q ),
    .X(_0209_));
 sky130_fd_sc_hd__o211a_1 _0698_ (.A1(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame1_bit5.Q ),
    .A2(_0209_),
    .B1(_0208_),
    .C1(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame1_bit4.Q ),
    .X(_0210_));
 sky130_fd_sc_hd__nand2_1 _0699_ (.A(net127),
    .B(_0054_),
    .Y(_0211_));
 sky130_fd_sc_hd__nor3_1 _0700_ (.A(net148),
    .B(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame1_bit5.Q ),
    .C(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame1_bit6.Q ),
    .Y(_0212_));
 sky130_fd_sc_hd__a221o_1 _0701_ (.A1(_0008_),
    .A2(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame1_bit5.Q ),
    .B1(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame1_bit6.Q ),
    .B2(_0211_),
    .C1(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame1_bit4.Q ),
    .X(_0213_));
 sky130_fd_sc_hd__or3b_1 _0702_ (.A(net156),
    .B(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame1_bit5.Q ),
    .C_N(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame1_bit6.Q ),
    .X(_0214_));
 sky130_fd_sc_hd__o311a_1 _0703_ (.A1(net238),
    .A2(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame1_bit5.Q ),
    .A3(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame1_bit6.Q ),
    .B1(_0214_),
    .C1(_0053_),
    .X(_0215_));
 sky130_fd_sc_hd__or3b_1 _0704_ (.A(net159),
    .B(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame1_bit5.Q ),
    .C_N(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame1_bit6.Q ),
    .X(_0216_));
 sky130_fd_sc_hd__o311a_1 _0705_ (.A1(net226),
    .A2(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame1_bit5.Q ),
    .A3(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame1_bit6.Q ),
    .B1(_0216_),
    .C1(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame1_bit4.Q ),
    .X(_0217_));
 sky130_fd_sc_hd__mux4_1 _0706_ (.A0(net227),
    .A1(net146),
    .A2(net153),
    .A3(net147),
    .S0(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame1_bit6.Q ),
    .S1(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame1_bit4.Q ),
    .X(_0218_));
 sky130_fd_sc_hd__o22a_1 _0707_ (.A1(_0215_),
    .A2(_0217_),
    .B1(_0218_),
    .B2(_0054_),
    .X(_0219_));
 sky130_fd_sc_hd__o21ai_1 _0708_ (.A1(_0212_),
    .A2(_0213_),
    .B1(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame1_bit7.Q ),
    .Y(_0220_));
 sky130_fd_sc_hd__o22a_1 _0709_ (.A1(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame1_bit7.Q ),
    .A2(_0219_),
    .B1(_0220_),
    .B2(_0210_),
    .X(net324));
 sky130_fd_sc_hd__dlxtp_1 _0710_ (.D(net467),
    .GATE(net446),
    .Q(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame0_bit31.Q ));
 sky130_fd_sc_hd__dlxtp_1 _0711_ (.D(net468),
    .GATE(net446),
    .Q(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame0_bit30.Q ));
 sky130_fd_sc_hd__dlxtp_1 _0712_ (.D(net102),
    .GATE(net447),
    .Q(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame0_bit29.Q ));
 sky130_fd_sc_hd__dlxtp_1 _0713_ (.D(net101),
    .GATE(net447),
    .Q(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame0_bit28.Q ));
 sky130_fd_sc_hd__dlxtp_1 _0714_ (.D(net471),
    .GATE(net446),
    .Q(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame0_bit27.Q ));
 sky130_fd_sc_hd__dlxtp_1 _0715_ (.D(net472),
    .GATE(net446),
    .Q(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame0_bit26.Q ));
 sky130_fd_sc_hd__dlxtp_1 _0716_ (.D(net98),
    .GATE(net448),
    .Q(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame0_bit25.Q ));
 sky130_fd_sc_hd__dlxtp_1 _0717_ (.D(net97),
    .GATE(net448),
    .Q(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame0_bit24.Q ));
 sky130_fd_sc_hd__dlxtp_1 _0718_ (.D(net475),
    .GATE(net445),
    .Q(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame0_bit23.Q ));
 sky130_fd_sc_hd__dlxtp_1 _0719_ (.D(net476),
    .GATE(net445),
    .Q(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame0_bit22.Q ));
 sky130_fd_sc_hd__dlxtp_1 _0720_ (.D(net94),
    .GATE(net447),
    .Q(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame0_bit21.Q ));
 sky130_fd_sc_hd__dlxtp_1 _0721_ (.D(net93),
    .GATE(net447),
    .Q(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame0_bit20.Q ));
 sky130_fd_sc_hd__dlxtp_1 _0722_ (.D(net91),
    .GATE(net447),
    .Q(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame0_bit19.Q ));
 sky130_fd_sc_hd__dlxtp_1 _0723_ (.D(net90),
    .GATE(net447),
    .Q(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame0_bit18.Q ));
 sky130_fd_sc_hd__dlxtp_1 _0724_ (.D(net89),
    .GATE(net444),
    .Q(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame0_bit17.Q ));
 sky130_fd_sc_hd__dlxtp_1 _0725_ (.D(net88),
    .GATE(net444),
    .Q(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame0_bit16.Q ));
 sky130_fd_sc_hd__dlxtp_1 _0726_ (.D(net87),
    .GATE(net444),
    .Q(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame0_bit15.Q ));
 sky130_fd_sc_hd__dlxtp_1 _0727_ (.D(net86),
    .GATE(net444),
    .Q(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame0_bit14.Q ));
 sky130_fd_sc_hd__dlxtp_1 _0728_ (.D(net85),
    .GATE(net444),
    .Q(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame0_bit13.Q ));
 sky130_fd_sc_hd__dlxtp_1 _0729_ (.D(net84),
    .GATE(net444),
    .Q(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame0_bit12.Q ));
 sky130_fd_sc_hd__dlxtp_1 _0730_ (.D(net83),
    .GATE(net444),
    .Q(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame0_bit11.Q ));
 sky130_fd_sc_hd__dlxtp_1 _0731_ (.D(net82),
    .GATE(net444),
    .Q(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame0_bit10.Q ));
 sky130_fd_sc_hd__dlxtp_1 _0732_ (.D(net112),
    .GATE(net444),
    .Q(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame0_bit9.Q ));
 sky130_fd_sc_hd__dlxtp_1 _0733_ (.D(net111),
    .GATE(net444),
    .Q(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame0_bit8.Q ));
 sky130_fd_sc_hd__dlxtp_1 _0734_ (.D(net110),
    .GATE(net446),
    .Q(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame0_bit7.Q ));
 sky130_fd_sc_hd__dlxtp_1 _0735_ (.D(net109),
    .GATE(net446),
    .Q(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame0_bit6.Q ));
 sky130_fd_sc_hd__dlxtp_1 _0736_ (.D(net108),
    .GATE(net446),
    .Q(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame0_bit5.Q ));
 sky130_fd_sc_hd__dlxtp_1 _0737_ (.D(net107),
    .GATE(net446),
    .Q(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame0_bit4.Q ));
 sky130_fd_sc_hd__dlxtp_1 _0738_ (.D(net106),
    .GATE(net446),
    .Q(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame0_bit3.Q ));
 sky130_fd_sc_hd__dlxtp_1 _0739_ (.D(net103),
    .GATE(net446),
    .Q(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame0_bit2.Q ));
 sky130_fd_sc_hd__dlxtp_1 _0740_ (.D(net92),
    .GATE(net445),
    .Q(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame0_bit1.Q ));
 sky130_fd_sc_hd__dlxtp_1 _0741_ (.D(net81),
    .GATE(net445),
    .Q(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame0_bit0.Q ));
 sky130_fd_sc_hd__dlxtp_1 _0742_ (.D(net467),
    .GATE(net438),
    .Q(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame1_bit31.Q ));
 sky130_fd_sc_hd__dlxtp_1 _0743_ (.D(net468),
    .GATE(net438),
    .Q(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame1_bit30.Q ));
 sky130_fd_sc_hd__dlxtp_1 _0744_ (.D(net469),
    .GATE(net437),
    .Q(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame1_bit29.Q ));
 sky130_fd_sc_hd__dlxtp_1 _0745_ (.D(net470),
    .GATE(net437),
    .Q(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame1_bit28.Q ));
 sky130_fd_sc_hd__dlxtp_1 _0746_ (.D(net471),
    .GATE(net436),
    .Q(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame1_bit27.Q ));
 sky130_fd_sc_hd__dlxtp_1 _0747_ (.D(net472),
    .GATE(net436),
    .Q(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame1_bit26.Q ));
 sky130_fd_sc_hd__dlxtp_1 _0748_ (.D(net473),
    .GATE(net438),
    .Q(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame1_bit25.Q ));
 sky130_fd_sc_hd__dlxtp_1 _0749_ (.D(net474),
    .GATE(net438),
    .Q(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame1_bit24.Q ));
 sky130_fd_sc_hd__dlxtp_1 _0750_ (.D(net475),
    .GATE(net438),
    .Q(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame1_bit23.Q ));
 sky130_fd_sc_hd__dlxtp_1 _0751_ (.D(net476),
    .GATE(net438),
    .Q(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame1_bit22.Q ));
 sky130_fd_sc_hd__dlxtp_1 _0752_ (.D(net94),
    .GATE(net439),
    .Q(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame1_bit21.Q ));
 sky130_fd_sc_hd__dlxtp_1 _0753_ (.D(net93),
    .GATE(net437),
    .Q(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame1_bit20.Q ));
 sky130_fd_sc_hd__dlxtp_1 _0754_ (.D(net91),
    .GATE(net437),
    .Q(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame1_bit19.Q ));
 sky130_fd_sc_hd__dlxtp_1 _0755_ (.D(net90),
    .GATE(net437),
    .Q(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame1_bit18.Q ));
 sky130_fd_sc_hd__dlxtp_1 _0756_ (.D(net89),
    .GATE(net438),
    .Q(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame1_bit17.Q ));
 sky130_fd_sc_hd__dlxtp_1 _0757_ (.D(net88),
    .GATE(net438),
    .Q(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame1_bit16.Q ));
 sky130_fd_sc_hd__dlxtp_1 _0758_ (.D(net87),
    .GATE(net439),
    .Q(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame1_bit15.Q ));
 sky130_fd_sc_hd__dlxtp_1 _0759_ (.D(net86),
    .GATE(net437),
    .Q(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame1_bit14.Q ));
 sky130_fd_sc_hd__dlxtp_1 _0760_ (.D(net85),
    .GATE(net439),
    .Q(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame1_bit13.Q ));
 sky130_fd_sc_hd__dlxtp_1 _0761_ (.D(net84),
    .GATE(net439),
    .Q(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame1_bit12.Q ));
 sky130_fd_sc_hd__dlxtp_1 _0762_ (.D(net83),
    .GATE(net437),
    .Q(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame1_bit11.Q ));
 sky130_fd_sc_hd__dlxtp_1 _0763_ (.D(net82),
    .GATE(net437),
    .Q(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame1_bit10.Q ));
 sky130_fd_sc_hd__dlxtp_1 _0764_ (.D(net112),
    .GATE(net438),
    .Q(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame1_bit9.Q ));
 sky130_fd_sc_hd__dlxtp_1 _0765_ (.D(net111),
    .GATE(net438),
    .Q(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame1_bit8.Q ));
 sky130_fd_sc_hd__dlxtp_1 _0766_ (.D(net110),
    .GATE(net436),
    .Q(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame1_bit7.Q ));
 sky130_fd_sc_hd__dlxtp_1 _0767_ (.D(net109),
    .GATE(net436),
    .Q(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame1_bit6.Q ));
 sky130_fd_sc_hd__dlxtp_1 _0768_ (.D(net108),
    .GATE(net436),
    .Q(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame1_bit5.Q ));
 sky130_fd_sc_hd__dlxtp_1 _0769_ (.D(net107),
    .GATE(net436),
    .Q(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame1_bit4.Q ));
 sky130_fd_sc_hd__dlxtp_1 _0770_ (.D(net106),
    .GATE(net436),
    .Q(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame1_bit3.Q ));
 sky130_fd_sc_hd__dlxtp_1 _0771_ (.D(net103),
    .GATE(net436),
    .Q(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame1_bit2.Q ));
 sky130_fd_sc_hd__dlxtp_1 _0772_ (.D(net92),
    .GATE(net436),
    .Q(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame1_bit1.Q ));
 sky130_fd_sc_hd__dlxtp_1 _0773_ (.D(net81),
    .GATE(net436),
    .Q(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame1_bit0.Q ));
 sky130_fd_sc_hd__dlxtp_1 _0774_ (.D(net467),
    .GATE(net427),
    .Q(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame2_bit31.Q ));
 sky130_fd_sc_hd__dlxtp_1 _0775_ (.D(net468),
    .GATE(net427),
    .Q(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame2_bit30.Q ));
 sky130_fd_sc_hd__dlxtp_1 _0776_ (.D(net469),
    .GATE(net430),
    .Q(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame2_bit29.Q ));
 sky130_fd_sc_hd__dlxtp_1 _0777_ (.D(net470),
    .GATE(net430),
    .Q(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame2_bit28.Q ));
 sky130_fd_sc_hd__dlxtp_1 _0778_ (.D(net471),
    .GATE(net429),
    .Q(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame2_bit27.Q ));
 sky130_fd_sc_hd__dlxtp_1 _0779_ (.D(net472),
    .GATE(net427),
    .Q(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame2_bit26.Q ));
 sky130_fd_sc_hd__dlxtp_1 _0780_ (.D(net473),
    .GATE(net427),
    .Q(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame2_bit25.Q ));
 sky130_fd_sc_hd__dlxtp_1 _0781_ (.D(net474),
    .GATE(net427),
    .Q(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame2_bit24.Q ));
 sky130_fd_sc_hd__dlxtp_1 _0782_ (.D(net475),
    .GATE(net430),
    .Q(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame2_bit23.Q ));
 sky130_fd_sc_hd__dlxtp_1 _0783_ (.D(net476),
    .GATE(net430),
    .Q(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame2_bit22.Q ));
 sky130_fd_sc_hd__dlxtp_1 _0784_ (.D(net94),
    .GATE(net427),
    .Q(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame2_bit21.Q ));
 sky130_fd_sc_hd__dlxtp_1 _0785_ (.D(net93),
    .GATE(net427),
    .Q(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame2_bit20.Q ));
 sky130_fd_sc_hd__dlxtp_1 _0786_ (.D(net91),
    .GATE(net428),
    .Q(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame2_bit19.Q ));
 sky130_fd_sc_hd__dlxtp_1 _0787_ (.D(net90),
    .GATE(net429),
    .Q(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame2_bit18.Q ));
 sky130_fd_sc_hd__dlxtp_1 _0788_ (.D(net89),
    .GATE(net428),
    .Q(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame2_bit17.Q ));
 sky130_fd_sc_hd__dlxtp_1 _0789_ (.D(net88),
    .GATE(net428),
    .Q(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame2_bit16.Q ));
 sky130_fd_sc_hd__dlxtp_1 _0790_ (.D(net87),
    .GATE(net430),
    .Q(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame2_bit15.Q ));
 sky130_fd_sc_hd__dlxtp_1 _0791_ (.D(net86),
    .GATE(net430),
    .Q(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame2_bit14.Q ));
 sky130_fd_sc_hd__dlxtp_1 _0792_ (.D(net85),
    .GATE(net430),
    .Q(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame2_bit13.Q ));
 sky130_fd_sc_hd__dlxtp_1 _0793_ (.D(net84),
    .GATE(net430),
    .Q(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame2_bit12.Q ));
 sky130_fd_sc_hd__dlxtp_1 _0794_ (.D(net83),
    .GATE(net429),
    .Q(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame2_bit11.Q ));
 sky130_fd_sc_hd__dlxtp_1 _0795_ (.D(net82),
    .GATE(net427),
    .Q(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame2_bit10.Q ));
 sky130_fd_sc_hd__dlxtp_1 _0796_ (.D(net112),
    .GATE(net428),
    .Q(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame2_bit9.Q ));
 sky130_fd_sc_hd__dlxtp_1 _0797_ (.D(net111),
    .GATE(net428),
    .Q(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame2_bit8.Q ));
 sky130_fd_sc_hd__dlxtp_1 _0798_ (.D(net110),
    .GATE(net430),
    .Q(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame2_bit7.Q ));
 sky130_fd_sc_hd__dlxtp_1 _0799_ (.D(net109),
    .GATE(net430),
    .Q(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame2_bit6.Q ));
 sky130_fd_sc_hd__dlxtp_1 _0800_ (.D(net108),
    .GATE(net427),
    .Q(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame2_bit5.Q ));
 sky130_fd_sc_hd__dlxtp_1 _0801_ (.D(net107),
    .GATE(net427),
    .Q(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame2_bit4.Q ));
 sky130_fd_sc_hd__dlxtp_1 _0802_ (.D(net106),
    .GATE(net428),
    .Q(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame2_bit3.Q ));
 sky130_fd_sc_hd__dlxtp_1 _0803_ (.D(net103),
    .GATE(net428),
    .Q(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame2_bit2.Q ));
 sky130_fd_sc_hd__dlxtp_1 _0804_ (.D(net92),
    .GATE(net428),
    .Q(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame2_bit1.Q ));
 sky130_fd_sc_hd__dlxtp_1 _0805_ (.D(net81),
    .GATE(net428),
    .Q(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame2_bit0.Q ));
 sky130_fd_sc_hd__dlxtp_1 _0806_ (.D(net467),
    .GATE(net420),
    .Q(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame3_bit31.Q ));
 sky130_fd_sc_hd__dlxtp_1 _0807_ (.D(net468),
    .GATE(net420),
    .Q(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame3_bit30.Q ));
 sky130_fd_sc_hd__dlxtp_1 _0808_ (.D(net469),
    .GATE(net423),
    .Q(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame3_bit29.Q ));
 sky130_fd_sc_hd__dlxtp_1 _0809_ (.D(net470),
    .GATE(net423),
    .Q(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame3_bit28.Q ));
 sky130_fd_sc_hd__dlxtp_1 _0810_ (.D(net471),
    .GATE(net422),
    .Q(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame3_bit27.Q ));
 sky130_fd_sc_hd__dlxtp_1 _0811_ (.D(net472),
    .GATE(net422),
    .Q(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame3_bit26.Q ));
 sky130_fd_sc_hd__dlxtp_1 _0812_ (.D(net473),
    .GATE(net422),
    .Q(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame3_bit25.Q ));
 sky130_fd_sc_hd__dlxtp_1 _0813_ (.D(net474),
    .GATE(net422),
    .Q(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame3_bit24.Q ));
 sky130_fd_sc_hd__dlxtp_1 _0814_ (.D(net475),
    .GATE(net420),
    .Q(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame3_bit23.Q ));
 sky130_fd_sc_hd__dlxtp_1 _0815_ (.D(net476),
    .GATE(net420),
    .Q(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame3_bit22.Q ));
 sky130_fd_sc_hd__dlxtp_1 _0816_ (.D(net94),
    .GATE(net422),
    .Q(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame3_bit21.Q ));
 sky130_fd_sc_hd__dlxtp_1 _0817_ (.D(net93),
    .GATE(net422),
    .Q(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame3_bit20.Q ));
 sky130_fd_sc_hd__dlxtp_1 _0818_ (.D(net91),
    .GATE(net423),
    .Q(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame3_bit19.Q ));
 sky130_fd_sc_hd__dlxtp_1 _0819_ (.D(net90),
    .GATE(net421),
    .Q(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame3_bit18.Q ));
 sky130_fd_sc_hd__dlxtp_1 _0820_ (.D(net89),
    .GATE(net421),
    .Q(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame3_bit17.Q ));
 sky130_fd_sc_hd__dlxtp_1 _0821_ (.D(net88),
    .GATE(net421),
    .Q(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame3_bit16.Q ));
 sky130_fd_sc_hd__dlxtp_1 _0822_ (.D(net87),
    .GATE(net420),
    .Q(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame3_bit15.Q ));
 sky130_fd_sc_hd__dlxtp_1 _0823_ (.D(net86),
    .GATE(net420),
    .Q(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame3_bit14.Q ));
 sky130_fd_sc_hd__dlxtp_1 _0824_ (.D(net85),
    .GATE(net420),
    .Q(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame3_bit13.Q ));
 sky130_fd_sc_hd__dlxtp_1 _0825_ (.D(net84),
    .GATE(net420),
    .Q(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame3_bit12.Q ));
 sky130_fd_sc_hd__dlxtp_1 _0826_ (.D(net83),
    .GATE(net422),
    .Q(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame3_bit11.Q ));
 sky130_fd_sc_hd__dlxtp_1 _0827_ (.D(net82),
    .GATE(net422),
    .Q(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame3_bit10.Q ));
 sky130_fd_sc_hd__dlxtp_1 _0828_ (.D(net112),
    .GATE(net421),
    .Q(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame3_bit9.Q ));
 sky130_fd_sc_hd__dlxtp_1 _0829_ (.D(net111),
    .GATE(net421),
    .Q(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame3_bit8.Q ));
 sky130_fd_sc_hd__dlxtp_1 _0830_ (.D(net110),
    .GATE(net420),
    .Q(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame3_bit7.Q ));
 sky130_fd_sc_hd__dlxtp_1 _0831_ (.D(net109),
    .GATE(net420),
    .Q(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame3_bit6.Q ));
 sky130_fd_sc_hd__dlxtp_1 _0832_ (.D(net108),
    .GATE(net422),
    .Q(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame3_bit5.Q ));
 sky130_fd_sc_hd__dlxtp_1 _0833_ (.D(net107),
    .GATE(net422),
    .Q(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame3_bit4.Q ));
 sky130_fd_sc_hd__dlxtp_1 _0834_ (.D(net106),
    .GATE(net421),
    .Q(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame3_bit3.Q ));
 sky130_fd_sc_hd__dlxtp_1 _0835_ (.D(net103),
    .GATE(net421),
    .Q(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame3_bit2.Q ));
 sky130_fd_sc_hd__dlxtp_1 _0836_ (.D(net92),
    .GATE(net421),
    .Q(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame3_bit1.Q ));
 sky130_fd_sc_hd__dlxtp_1 _0837_ (.D(net81),
    .GATE(net421),
    .Q(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame3_bit0.Q ));
 sky130_fd_sc_hd__dlxtp_1 _0838_ (.D(net467),
    .GATE(net414),
    .Q(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame4_bit31.Q ));
 sky130_fd_sc_hd__dlxtp_1 _0839_ (.D(net468),
    .GATE(net414),
    .Q(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame4_bit30.Q ));
 sky130_fd_sc_hd__dlxtp_1 _0840_ (.D(net469),
    .GATE(net415),
    .Q(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame4_bit29.Q ));
 sky130_fd_sc_hd__dlxtp_1 _0841_ (.D(net470),
    .GATE(net415),
    .Q(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame4_bit28.Q ));
 sky130_fd_sc_hd__dlxtp_1 _0842_ (.D(net471),
    .GATE(net411),
    .Q(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame4_bit27.Q ));
 sky130_fd_sc_hd__dlxtp_1 _0843_ (.D(net472),
    .GATE(net411),
    .Q(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame4_bit26.Q ));
 sky130_fd_sc_hd__dlxtp_1 _0844_ (.D(net473),
    .GATE(net411),
    .Q(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame4_bit25.Q ));
 sky130_fd_sc_hd__dlxtp_1 _0845_ (.D(net474),
    .GATE(net411),
    .Q(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame4_bit24.Q ));
 sky130_fd_sc_hd__dlxtp_1 _0846_ (.D(net475),
    .GATE(net412),
    .Q(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame4_bit23.Q ));
 sky130_fd_sc_hd__dlxtp_1 _0847_ (.D(net476),
    .GATE(net412),
    .Q(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame4_bit22.Q ));
 sky130_fd_sc_hd__dlxtp_1 _0848_ (.D(net94),
    .GATE(net415),
    .Q(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame4_bit21.Q ));
 sky130_fd_sc_hd__dlxtp_1 _0849_ (.D(net93),
    .GATE(net415),
    .Q(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame4_bit20.Q ));
 sky130_fd_sc_hd__dlxtp_1 _0850_ (.D(net91),
    .GATE(net411),
    .Q(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame4_bit19.Q ));
 sky130_fd_sc_hd__dlxtp_1 _0851_ (.D(net90),
    .GATE(net411),
    .Q(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame4_bit18.Q ));
 sky130_fd_sc_hd__dlxtp_1 _0852_ (.D(net89),
    .GATE(net412),
    .Q(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame4_bit17.Q ));
 sky130_fd_sc_hd__dlxtp_1 _0853_ (.D(net88),
    .GATE(net412),
    .Q(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame4_bit16.Q ));
 sky130_fd_sc_hd__dlxtp_1 _0854_ (.D(net87),
    .GATE(net415),
    .Q(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame4_bit15.Q ));
 sky130_fd_sc_hd__dlxtp_1 _0855_ (.D(net86),
    .GATE(net415),
    .Q(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame4_bit14.Q ));
 sky130_fd_sc_hd__dlxtp_1 _0856_ (.D(net85),
    .GATE(net414),
    .Q(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame4_bit13.Q ));
 sky130_fd_sc_hd__dlxtp_1 _0857_ (.D(net84),
    .GATE(net414),
    .Q(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame4_bit12.Q ));
 sky130_fd_sc_hd__dlxtp_1 _0858_ (.D(net83),
    .GATE(net413),
    .Q(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame4_bit11.Q ));
 sky130_fd_sc_hd__dlxtp_1 _0859_ (.D(net82),
    .GATE(net413),
    .Q(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame4_bit10.Q ));
 sky130_fd_sc_hd__dlxtp_1 _0860_ (.D(net112),
    .GATE(net413),
    .Q(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame4_bit9.Q ));
 sky130_fd_sc_hd__dlxtp_1 _0861_ (.D(net111),
    .GATE(net413),
    .Q(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame4_bit8.Q ));
 sky130_fd_sc_hd__dlxtp_1 _0862_ (.D(net110),
    .GATE(net415),
    .Q(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame4_bit7.Q ));
 sky130_fd_sc_hd__dlxtp_1 _0863_ (.D(net109),
    .GATE(net415),
    .Q(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame4_bit6.Q ));
 sky130_fd_sc_hd__dlxtp_1 _0864_ (.D(net108),
    .GATE(net415),
    .Q(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame4_bit5.Q ));
 sky130_fd_sc_hd__dlxtp_1 _0865_ (.D(net107),
    .GATE(net415),
    .Q(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame4_bit4.Q ));
 sky130_fd_sc_hd__dlxtp_1 _0866_ (.D(net106),
    .GATE(net411),
    .Q(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame4_bit3.Q ));
 sky130_fd_sc_hd__dlxtp_1 _0867_ (.D(net103),
    .GATE(net411),
    .Q(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame4_bit2.Q ));
 sky130_fd_sc_hd__dlxtp_1 _0868_ (.D(net92),
    .GATE(net411),
    .Q(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame4_bit1.Q ));
 sky130_fd_sc_hd__dlxtp_1 _0869_ (.D(net81),
    .GATE(net411),
    .Q(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame4_bit0.Q ));
 sky130_fd_sc_hd__dlxtp_1 _0870_ (.D(net467),
    .GATE(net403),
    .Q(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame5_bit31.Q ));
 sky130_fd_sc_hd__dlxtp_1 _0871_ (.D(net468),
    .GATE(net402),
    .Q(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame5_bit30.Q ));
 sky130_fd_sc_hd__dlxtp_1 _0872_ (.D(net469),
    .GATE(net402),
    .Q(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame5_bit29.Q ));
 sky130_fd_sc_hd__dlxtp_1 _0873_ (.D(net470),
    .GATE(net402),
    .Q(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame5_bit28.Q ));
 sky130_fd_sc_hd__dlxtp_1 _0874_ (.D(net471),
    .GATE(net402),
    .Q(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame5_bit27.Q ));
 sky130_fd_sc_hd__dlxtp_1 _0875_ (.D(net472),
    .GATE(net402),
    .Q(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame5_bit26.Q ));
 sky130_fd_sc_hd__dlxtp_1 _0876_ (.D(net473),
    .GATE(net404),
    .Q(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame5_bit25.Q ));
 sky130_fd_sc_hd__dlxtp_1 _0877_ (.D(net474),
    .GATE(net404),
    .Q(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame5_bit24.Q ));
 sky130_fd_sc_hd__dlxtp_1 _0878_ (.D(net475),
    .GATE(net402),
    .Q(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame5_bit23.Q ));
 sky130_fd_sc_hd__dlxtp_1 _0879_ (.D(net476),
    .GATE(net402),
    .Q(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame5_bit22.Q ));
 sky130_fd_sc_hd__dlxtp_1 _0880_ (.D(net94),
    .GATE(net403),
    .Q(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame5_bit21.Q ));
 sky130_fd_sc_hd__dlxtp_1 _0881_ (.D(net93),
    .GATE(net403),
    .Q(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame5_bit20.Q ));
 sky130_fd_sc_hd__dlxtp_1 _0882_ (.D(net91),
    .GATE(net402),
    .Q(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame5_bit19.Q ));
 sky130_fd_sc_hd__dlxtp_1 _0883_ (.D(net90),
    .GATE(net402),
    .Q(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame5_bit18.Q ));
 sky130_fd_sc_hd__dlxtp_1 _0884_ (.D(net89),
    .GATE(net404),
    .Q(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame5_bit17.Q ));
 sky130_fd_sc_hd__dlxtp_1 _0885_ (.D(net88),
    .GATE(net404),
    .Q(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame5_bit16.Q ));
 sky130_fd_sc_hd__dlxtp_1 _0886_ (.D(net87),
    .GATE(net403),
    .Q(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame5_bit15.Q ));
 sky130_fd_sc_hd__dlxtp_1 _0887_ (.D(net86),
    .GATE(net403),
    .Q(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame5_bit14.Q ));
 sky130_fd_sc_hd__dlxtp_1 _0888_ (.D(net85),
    .GATE(net405),
    .Q(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame5_bit13.Q ));
 sky130_fd_sc_hd__dlxtp_1 _0889_ (.D(net84),
    .GATE(net405),
    .Q(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame5_bit12.Q ));
 sky130_fd_sc_hd__dlxtp_1 _0890_ (.D(net83),
    .GATE(net402),
    .Q(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame5_bit11.Q ));
 sky130_fd_sc_hd__dlxtp_1 _0891_ (.D(net82),
    .GATE(net404),
    .Q(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame5_bit10.Q ));
 sky130_fd_sc_hd__dlxtp_1 _0892_ (.D(net112),
    .GATE(net404),
    .Q(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame5_bit9.Q ));
 sky130_fd_sc_hd__dlxtp_1 _0893_ (.D(net111),
    .GATE(net404),
    .Q(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame5_bit8.Q ));
 sky130_fd_sc_hd__dlxtp_1 _0894_ (.D(net110),
    .GATE(net405),
    .Q(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame5_bit7.Q ));
 sky130_fd_sc_hd__dlxtp_1 _0895_ (.D(net109),
    .GATE(net405),
    .Q(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame5_bit6.Q ));
 sky130_fd_sc_hd__dlxtp_1 _0896_ (.D(net108),
    .GATE(net405),
    .Q(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame5_bit5.Q ));
 sky130_fd_sc_hd__dlxtp_1 _0897_ (.D(net107),
    .GATE(net405),
    .Q(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame5_bit4.Q ));
 sky130_fd_sc_hd__dlxtp_1 _0898_ (.D(net106),
    .GATE(net405),
    .Q(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame5_bit3.Q ));
 sky130_fd_sc_hd__dlxtp_1 _0899_ (.D(net103),
    .GATE(net405),
    .Q(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame5_bit2.Q ));
 sky130_fd_sc_hd__dlxtp_1 _0900_ (.D(net92),
    .GATE(net405),
    .Q(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame5_bit1.Q ));
 sky130_fd_sc_hd__dlxtp_1 _0901_ (.D(net81),
    .GATE(net405),
    .Q(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame5_bit0.Q ));
 sky130_fd_sc_hd__dlxtp_1 _0902_ (.D(net467),
    .GATE(net397),
    .Q(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame6_bit31.Q ));
 sky130_fd_sc_hd__dlxtp_1 _0903_ (.D(net468),
    .GATE(net396),
    .Q(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame6_bit30.Q ));
 sky130_fd_sc_hd__dlxtp_1 _0904_ (.D(net469),
    .GATE(net396),
    .Q(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame6_bit29.Q ));
 sky130_fd_sc_hd__dlxtp_1 _0905_ (.D(net470),
    .GATE(net396),
    .Q(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame6_bit28.Q ));
 sky130_fd_sc_hd__dlxtp_1 _0906_ (.D(net471),
    .GATE(net396),
    .Q(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame6_bit27.Q ));
 sky130_fd_sc_hd__dlxtp_1 _0907_ (.D(net472),
    .GATE(net396),
    .Q(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame6_bit26.Q ));
 sky130_fd_sc_hd__dlxtp_1 _0908_ (.D(net473),
    .GATE(net396),
    .Q(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame6_bit25.Q ));
 sky130_fd_sc_hd__dlxtp_1 _0909_ (.D(net474),
    .GATE(net396),
    .Q(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame6_bit24.Q ));
 sky130_fd_sc_hd__dlxtp_1 _0910_ (.D(net475),
    .GATE(net394),
    .Q(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame6_bit23.Q ));
 sky130_fd_sc_hd__dlxtp_1 _0911_ (.D(net476),
    .GATE(net394),
    .Q(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame6_bit22.Q ));
 sky130_fd_sc_hd__dlxtp_1 _0912_ (.D(net94),
    .GATE(net396),
    .Q(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame6_bit21.Q ));
 sky130_fd_sc_hd__dlxtp_1 _0913_ (.D(net93),
    .GATE(net395),
    .Q(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame6_bit20.Q ));
 sky130_fd_sc_hd__dlxtp_1 _0914_ (.D(net91),
    .GATE(net396),
    .Q(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame6_bit19.Q ));
 sky130_fd_sc_hd__dlxtp_1 _0915_ (.D(net90),
    .GATE(net396),
    .Q(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame6_bit18.Q ));
 sky130_fd_sc_hd__dlxtp_1 _0916_ (.D(net89),
    .GATE(net394),
    .Q(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame6_bit17.Q ));
 sky130_fd_sc_hd__dlxtp_1 _0917_ (.D(net88),
    .GATE(net394),
    .Q(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame6_bit16.Q ));
 sky130_fd_sc_hd__dlxtp_1 _0918_ (.D(net87),
    .GATE(net395),
    .Q(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame6_bit15.Q ));
 sky130_fd_sc_hd__dlxtp_1 _0919_ (.D(net86),
    .GATE(net395),
    .Q(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame6_bit14.Q ));
 sky130_fd_sc_hd__dlxtp_1 _0920_ (.D(net85),
    .GATE(net394),
    .Q(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame6_bit13.Q ));
 sky130_fd_sc_hd__dlxtp_1 _0921_ (.D(net84),
    .GATE(net394),
    .Q(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame6_bit12.Q ));
 sky130_fd_sc_hd__dlxtp_1 _0922_ (.D(net83),
    .GATE(net394),
    .Q(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame6_bit11.Q ));
 sky130_fd_sc_hd__dlxtp_1 _0923_ (.D(net82),
    .GATE(net394),
    .Q(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame6_bit10.Q ));
 sky130_fd_sc_hd__dlxtp_1 _0924_ (.D(net112),
    .GATE(net395),
    .Q(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame6_bit9.Q ));
 sky130_fd_sc_hd__dlxtp_1 _0925_ (.D(net111),
    .GATE(net394),
    .Q(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame6_bit8.Q ));
 sky130_fd_sc_hd__dlxtp_1 _0926_ (.D(net110),
    .GATE(net394),
    .Q(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame6_bit7.Q ));
 sky130_fd_sc_hd__dlxtp_1 _0927_ (.D(net109),
    .GATE(net395),
    .Q(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame6_bit6.Q ));
 sky130_fd_sc_hd__dlxtp_1 _0928_ (.D(net108),
    .GATE(net397),
    .Q(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame6_bit5.Q ));
 sky130_fd_sc_hd__dlxtp_1 _0929_ (.D(net107),
    .GATE(net397),
    .Q(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame6_bit4.Q ));
 sky130_fd_sc_hd__dlxtp_1 _0930_ (.D(net106),
    .GATE(net397),
    .Q(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame6_bit3.Q ));
 sky130_fd_sc_hd__dlxtp_1 _0931_ (.D(net103),
    .GATE(net397),
    .Q(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame6_bit2.Q ));
 sky130_fd_sc_hd__dlxtp_1 _0932_ (.D(net92),
    .GATE(net395),
    .Q(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame6_bit1.Q ));
 sky130_fd_sc_hd__dlxtp_1 _0933_ (.D(net81),
    .GATE(net395),
    .Q(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame6_bit0.Q ));
 sky130_fd_sc_hd__dlxtp_1 _0934_ (.D(net105),
    .GATE(net388),
    .Q(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame7_bit31.Q ));
 sky130_fd_sc_hd__dlxtp_1 _0935_ (.D(net104),
    .GATE(net388),
    .Q(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame7_bit30.Q ));
 sky130_fd_sc_hd__dlxtp_1 _0936_ (.D(net469),
    .GATE(net388),
    .Q(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame7_bit29.Q ));
 sky130_fd_sc_hd__dlxtp_1 _0937_ (.D(net470),
    .GATE(net388),
    .Q(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame7_bit28.Q ));
 sky130_fd_sc_hd__dlxtp_1 _0938_ (.D(net471),
    .GATE(net388),
    .Q(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame7_bit27.Q ));
 sky130_fd_sc_hd__dlxtp_1 _0939_ (.D(net472),
    .GATE(net387),
    .Q(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame7_bit26.Q ));
 sky130_fd_sc_hd__dlxtp_1 _0940_ (.D(net473),
    .GATE(net387),
    .Q(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame7_bit25.Q ));
 sky130_fd_sc_hd__dlxtp_1 _0941_ (.D(net474),
    .GATE(net387),
    .Q(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame7_bit24.Q ));
 sky130_fd_sc_hd__dlxtp_1 _0942_ (.D(net96),
    .GATE(net385),
    .Q(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame7_bit23.Q ));
 sky130_fd_sc_hd__dlxtp_1 _0943_ (.D(net95),
    .GATE(net386),
    .Q(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame7_bit22.Q ));
 sky130_fd_sc_hd__dlxtp_1 _0944_ (.D(net94),
    .GATE(net386),
    .Q(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame7_bit21.Q ));
 sky130_fd_sc_hd__dlxtp_1 _0945_ (.D(net93),
    .GATE(net388),
    .Q(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame7_bit20.Q ));
 sky130_fd_sc_hd__dlxtp_1 _0946_ (.D(net91),
    .GATE(net388),
    .Q(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame7_bit19.Q ));
 sky130_fd_sc_hd__dlxtp_1 _0947_ (.D(net90),
    .GATE(net388),
    .Q(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame7_bit18.Q ));
 sky130_fd_sc_hd__dlxtp_1 _0948_ (.D(net89),
    .GATE(net385),
    .Q(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame7_bit17.Q ));
 sky130_fd_sc_hd__dlxtp_1 _0949_ (.D(net88),
    .GATE(net385),
    .Q(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame7_bit16.Q ));
 sky130_fd_sc_hd__dlxtp_1 _0950_ (.D(net87),
    .GATE(net385),
    .Q(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame7_bit15.Q ));
 sky130_fd_sc_hd__dlxtp_1 _0951_ (.D(net86),
    .GATE(net386),
    .Q(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame7_bit14.Q ));
 sky130_fd_sc_hd__dlxtp_1 _0952_ (.D(net85),
    .GATE(net386),
    .Q(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame7_bit13.Q ));
 sky130_fd_sc_hd__dlxtp_1 _0953_ (.D(net84),
    .GATE(net386),
    .Q(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame7_bit12.Q ));
 sky130_fd_sc_hd__dlxtp_1 _0954_ (.D(net83),
    .GATE(net385),
    .Q(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame7_bit11.Q ));
 sky130_fd_sc_hd__dlxtp_1 _0955_ (.D(net82),
    .GATE(net385),
    .Q(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame7_bit10.Q ));
 sky130_fd_sc_hd__dlxtp_1 _0956_ (.D(net112),
    .GATE(net385),
    .Q(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame7_bit9.Q ));
 sky130_fd_sc_hd__dlxtp_1 _0957_ (.D(net111),
    .GATE(net385),
    .Q(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame7_bit8.Q ));
 sky130_fd_sc_hd__dlxtp_1 _0958_ (.D(net110),
    .GATE(net386),
    .Q(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame7_bit7.Q ));
 sky130_fd_sc_hd__dlxtp_1 _0959_ (.D(net109),
    .GATE(net386),
    .Q(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame7_bit6.Q ));
 sky130_fd_sc_hd__dlxtp_1 _0960_ (.D(net108),
    .GATE(net386),
    .Q(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame7_bit5.Q ));
 sky130_fd_sc_hd__dlxtp_1 _0961_ (.D(net107),
    .GATE(net386),
    .Q(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame7_bit4.Q ));
 sky130_fd_sc_hd__dlxtp_1 _0962_ (.D(net106),
    .GATE(net385),
    .Q(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame7_bit3.Q ));
 sky130_fd_sc_hd__dlxtp_1 _0963_ (.D(net103),
    .GATE(net385),
    .Q(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame7_bit2.Q ));
 sky130_fd_sc_hd__dlxtp_1 _0964_ (.D(net92),
    .GATE(net387),
    .Q(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame7_bit1.Q ));
 sky130_fd_sc_hd__dlxtp_1 _0965_ (.D(net81),
    .GATE(net387),
    .Q(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame7_bit0.Q ));
 sky130_fd_sc_hd__dlxtp_1 _0966_ (.D(net467),
    .GATE(net379),
    .Q(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame8_bit31.Q ));
 sky130_fd_sc_hd__dlxtp_1 _0967_ (.D(net468),
    .GATE(net379),
    .Q(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame8_bit30.Q ));
 sky130_fd_sc_hd__dlxtp_1 _0968_ (.D(net469),
    .GATE(net377),
    .Q(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame8_bit29.Q ));
 sky130_fd_sc_hd__dlxtp_1 _0969_ (.D(net470),
    .GATE(net377),
    .Q(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame8_bit28.Q ));
 sky130_fd_sc_hd__dlxtp_1 _0970_ (.D(net100),
    .GATE(net380),
    .Q(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame8_bit27.Q ));
 sky130_fd_sc_hd__dlxtp_1 _0971_ (.D(net99),
    .GATE(net380),
    .Q(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame8_bit26.Q ));
 sky130_fd_sc_hd__dlxtp_1 _0972_ (.D(net473),
    .GATE(net379),
    .Q(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame8_bit25.Q ));
 sky130_fd_sc_hd__dlxtp_1 _0973_ (.D(net474),
    .GATE(net380),
    .Q(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame8_bit24.Q ));
 sky130_fd_sc_hd__dlxtp_1 _0974_ (.D(net475),
    .GATE(net380),
    .Q(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame8_bit23.Q ));
 sky130_fd_sc_hd__dlxtp_1 _0975_ (.D(net476),
    .GATE(net378),
    .Q(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame8_bit22.Q ));
 sky130_fd_sc_hd__dlxtp_1 _0976_ (.D(net94),
    .GATE(net378),
    .Q(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame8_bit21.Q ));
 sky130_fd_sc_hd__dlxtp_1 _0977_ (.D(net93),
    .GATE(net378),
    .Q(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame8_bit20.Q ));
 sky130_fd_sc_hd__dlxtp_1 _0978_ (.D(net91),
    .GATE(net378),
    .Q(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame8_bit19.Q ));
 sky130_fd_sc_hd__dlxtp_1 _0979_ (.D(net90),
    .GATE(net378),
    .Q(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame8_bit18.Q ));
 sky130_fd_sc_hd__dlxtp_1 _0980_ (.D(net89),
    .GATE(net378),
    .Q(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame8_bit17.Q ));
 sky130_fd_sc_hd__dlxtp_1 _0981_ (.D(net88),
    .GATE(net380),
    .Q(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame8_bit16.Q ));
 sky130_fd_sc_hd__dlxtp_1 _0982_ (.D(net87),
    .GATE(net380),
    .Q(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame8_bit15.Q ));
 sky130_fd_sc_hd__dlxtp_1 _0983_ (.D(net86),
    .GATE(net380),
    .Q(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame8_bit14.Q ));
 sky130_fd_sc_hd__dlxtp_1 _0984_ (.D(net85),
    .GATE(net377),
    .Q(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame8_bit13.Q ));
 sky130_fd_sc_hd__dlxtp_1 _0985_ (.D(net84),
    .GATE(net377),
    .Q(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame8_bit12.Q ));
 sky130_fd_sc_hd__dlxtp_1 _0986_ (.D(net83),
    .GATE(net378),
    .Q(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame8_bit11.Q ));
 sky130_fd_sc_hd__dlxtp_1 _0987_ (.D(net82),
    .GATE(net378),
    .Q(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame8_bit10.Q ));
 sky130_fd_sc_hd__dlxtp_1 _0988_ (.D(net112),
    .GATE(net378),
    .Q(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame8_bit9.Q ));
 sky130_fd_sc_hd__dlxtp_1 _0989_ (.D(net111),
    .GATE(net378),
    .Q(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame8_bit8.Q ));
 sky130_fd_sc_hd__dlxtp_1 _0990_ (.D(net110),
    .GATE(net380),
    .Q(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame8_bit7.Q ));
 sky130_fd_sc_hd__dlxtp_1 _0991_ (.D(net109),
    .GATE(net380),
    .Q(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame8_bit6.Q ));
 sky130_fd_sc_hd__dlxtp_1 _0992_ (.D(net108),
    .GATE(net377),
    .Q(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame8_bit5.Q ));
 sky130_fd_sc_hd__dlxtp_1 _0993_ (.D(net107),
    .GATE(net377),
    .Q(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame8_bit4.Q ));
 sky130_fd_sc_hd__dlxtp_1 _0994_ (.D(net106),
    .GATE(net377),
    .Q(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame8_bit3.Q ));
 sky130_fd_sc_hd__dlxtp_1 _0995_ (.D(net103),
    .GATE(net377),
    .Q(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame8_bit2.Q ));
 sky130_fd_sc_hd__dlxtp_1 _0996_ (.D(net92),
    .GATE(net377),
    .Q(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame8_bit1.Q ));
 sky130_fd_sc_hd__dlxtp_1 _0997_ (.D(net81),
    .GATE(net377),
    .Q(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame8_bit0.Q ));
 sky130_fd_sc_hd__dlxtp_1 _0998_ (.D(net467),
    .GATE(net372),
    .Q(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame9_bit31.Q ));
 sky130_fd_sc_hd__dlxtp_1 _0999_ (.D(net468),
    .GATE(net372),
    .Q(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame9_bit30.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1000_ (.D(net469),
    .GATE(net219),
    .Q(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame9_bit29.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1001_ (.D(net470),
    .GATE(net372),
    .Q(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame9_bit28.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1002_ (.D(net471),
    .GATE(net372),
    .Q(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame9_bit27.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1003_ (.D(net472),
    .GATE(net372),
    .Q(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame9_bit26.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1004_ (.D(net473),
    .GATE(net372),
    .Q(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame9_bit25.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1005_ (.D(net474),
    .GATE(net372),
    .Q(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame9_bit24.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1006_ (.D(net475),
    .GATE(net372),
    .Q(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame9_bit23.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1007_ (.D(net476),
    .GATE(net372),
    .Q(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_ConfigMem.Inst_frame9_bit22.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1008_ (.D(net449),
    .GATE(net440),
    .Q(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame0_bit31.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1009_ (.D(net450),
    .GATE(net440),
    .Q(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame0_bit30.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1010_ (.D(net208),
    .GATE(net442),
    .Q(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame0_bit29.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1011_ (.D(net207),
    .GATE(net442),
    .Q(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame0_bit28.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1012_ (.D(net206),
    .GATE(net442),
    .Q(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame0_bit27.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1013_ (.D(net205),
    .GATE(net442),
    .Q(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame0_bit26.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1014_ (.D(net204),
    .GATE(net441),
    .Q(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame0_bit25.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1015_ (.D(net203),
    .GATE(net441),
    .Q(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame0_bit24.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1016_ (.D(net457),
    .GATE(net440),
    .Q(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame0_bit23.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1017_ (.D(net458),
    .GATE(net440),
    .Q(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame0_bit22.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1018_ (.D(net459),
    .GATE(net440),
    .Q(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame0_bit21.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1019_ (.D(net460),
    .GATE(net440),
    .Q(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame0_bit20.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1020_ (.D(net461),
    .GATE(net441),
    .Q(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame0_bit19.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1021_ (.D(net462),
    .GATE(net440),
    .Q(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame0_bit18.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1022_ (.D(net463),
    .GATE(net443),
    .Q(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame0_bit17.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1023_ (.D(net464),
    .GATE(net443),
    .Q(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame0_bit16.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1024_ (.D(net465),
    .GATE(net442),
    .Q(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame0_bit15.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1025_ (.D(net466),
    .GATE(net442),
    .Q(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame0_bit14.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1026_ (.D(net193),
    .GATE(net443),
    .Q(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame0_bit13.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1027_ (.D(net192),
    .GATE(net443),
    .Q(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame0_bit12.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1028_ (.D(net191),
    .GATE(net442),
    .Q(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame0_bit11.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1029_ (.D(net190),
    .GATE(net442),
    .Q(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame0_bit10.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1030_ (.D(net218),
    .GATE(net442),
    .Q(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame0_bit9.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1031_ (.D(net217),
    .GATE(net442),
    .Q(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame0_bit8.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1032_ (.D(net216),
    .GATE(net440),
    .Q(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame0_bit7.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1033_ (.D(net215),
    .GATE(net440),
    .Q(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame0_bit6.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1034_ (.D(net214),
    .GATE(net441),
    .Q(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame0_bit5.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1035_ (.D(net213),
    .GATE(net441),
    .Q(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame0_bit4.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1036_ (.D(net212),
    .GATE(net441),
    .Q(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame0_bit3.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1037_ (.D(net209),
    .GATE(net441),
    .Q(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame0_bit2.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1038_ (.D(net198),
    .GATE(net440),
    .Q(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame0_bit1.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1039_ (.D(net189),
    .GATE(net441),
    .Q(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame0_bit0.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1040_ (.D(net449),
    .GATE(net432),
    .Q(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame1_bit31.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1041_ (.D(net450),
    .GATE(net432),
    .Q(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame1_bit30.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1042_ (.D(net451),
    .GATE(net433),
    .Q(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame1_bit29.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1043_ (.D(net452),
    .GATE(net433),
    .Q(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame1_bit28.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1044_ (.D(net453),
    .GATE(net434),
    .Q(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame1_bit27.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1045_ (.D(net454),
    .GATE(net434),
    .Q(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame1_bit26.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1046_ (.D(net455),
    .GATE(net432),
    .Q(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame1_bit25.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1047_ (.D(net456),
    .GATE(net432),
    .Q(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame1_bit24.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1048_ (.D(net457),
    .GATE(net432),
    .Q(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame1_bit23.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1049_ (.D(net458),
    .GATE(net432),
    .Q(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame1_bit22.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1050_ (.D(net459),
    .GATE(net433),
    .Q(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame1_bit21.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1051_ (.D(net460),
    .GATE(net433),
    .Q(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame1_bit20.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1052_ (.D(net461),
    .GATE(net434),
    .Q(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame1_bit19.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1053_ (.D(net462),
    .GATE(net434),
    .Q(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame1_bit18.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1054_ (.D(net463),
    .GATE(net432),
    .Q(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame1_bit17.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1055_ (.D(net464),
    .GATE(net432),
    .Q(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame1_bit16.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1056_ (.D(net465),
    .GATE(net433),
    .Q(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame1_bit15.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1057_ (.D(net466),
    .GATE(net433),
    .Q(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame1_bit14.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1058_ (.D(net193),
    .GATE(net433),
    .Q(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame1_bit13.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1059_ (.D(net192),
    .GATE(net433),
    .Q(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame1_bit12.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1060_ (.D(net191),
    .GATE(net434),
    .Q(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame1_bit11.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1061_ (.D(net190),
    .GATE(net434),
    .Q(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame1_bit10.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1062_ (.D(net218),
    .GATE(net432),
    .Q(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame1_bit9.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1063_ (.D(net217),
    .GATE(net432),
    .Q(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame1_bit8.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1064_ (.D(net216),
    .GATE(net435),
    .Q(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame1_bit7.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1065_ (.D(net215),
    .GATE(net435),
    .Q(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame1_bit6.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1066_ (.D(net214),
    .GATE(net435),
    .Q(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame1_bit5.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1067_ (.D(net213),
    .GATE(net435),
    .Q(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame1_bit4.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1068_ (.D(net212),
    .GATE(net435),
    .Q(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame1_bit3.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1069_ (.D(net209),
    .GATE(net435),
    .Q(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame1_bit2.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1070_ (.D(net198),
    .GATE(net435),
    .Q(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame1_bit1.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1071_ (.D(net189),
    .GATE(net435),
    .Q(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame1_bit0.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1072_ (.D(net449),
    .GATE(net424),
    .Q(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame2_bit31.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1073_ (.D(net450),
    .GATE(net424),
    .Q(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame2_bit30.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1074_ (.D(net451),
    .GATE(net431),
    .Q(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame2_bit29.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1075_ (.D(net452),
    .GATE(net431),
    .Q(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame2_bit28.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1076_ (.D(net453),
    .GATE(net426),
    .Q(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame2_bit27.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1077_ (.D(net454),
    .GATE(net426),
    .Q(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame2_bit26.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1078_ (.D(net455),
    .GATE(net424),
    .Q(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame2_bit25.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1079_ (.D(net456),
    .GATE(net424),
    .Q(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame2_bit24.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1080_ (.D(net457),
    .GATE(net426),
    .Q(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame2_bit23.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1081_ (.D(net458),
    .GATE(net426),
    .Q(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame2_bit22.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1082_ (.D(net459),
    .GATE(net425),
    .Q(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame2_bit21.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1083_ (.D(net460),
    .GATE(net425),
    .Q(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame2_bit20.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1084_ (.D(net197),
    .GATE(net426),
    .Q(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame2_bit19.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1085_ (.D(net196),
    .GATE(net426),
    .Q(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame2_bit18.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1086_ (.D(net463),
    .GATE(net425),
    .Q(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame2_bit17.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1087_ (.D(net464),
    .GATE(net425),
    .Q(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame2_bit16.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1088_ (.D(net465),
    .GATE(net424),
    .Q(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame2_bit15.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1089_ (.D(net466),
    .GATE(net424),
    .Q(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame2_bit14.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1090_ (.D(net193),
    .GATE(net431),
    .Q(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame2_bit13.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1091_ (.D(net192),
    .GATE(net431),
    .Q(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame2_bit12.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1092_ (.D(net191),
    .GATE(net426),
    .Q(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame2_bit11.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1093_ (.D(net190),
    .GATE(net426),
    .Q(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame2_bit10.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1094_ (.D(net218),
    .GATE(net424),
    .Q(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame2_bit9.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1095_ (.D(net217),
    .GATE(net424),
    .Q(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame2_bit8.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1096_ (.D(net216),
    .GATE(net426),
    .Q(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame2_bit7.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1097_ (.D(net215),
    .GATE(net425),
    .Q(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame2_bit6.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1098_ (.D(net214),
    .GATE(net425),
    .Q(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame2_bit5.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1099_ (.D(net213),
    .GATE(net425),
    .Q(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame2_bit4.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1100_ (.D(net212),
    .GATE(net425),
    .Q(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame2_bit3.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1101_ (.D(net209),
    .GATE(net425),
    .Q(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame2_bit2.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1102_ (.D(net198),
    .GATE(net424),
    .Q(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame2_bit1.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1103_ (.D(net189),
    .GATE(net424),
    .Q(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame2_bit0.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1104_ (.D(net449),
    .GATE(net416),
    .Q(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame3_bit31.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1105_ (.D(net450),
    .GATE(net416),
    .Q(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame3_bit30.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1106_ (.D(net451),
    .GATE(net417),
    .Q(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame3_bit29.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1107_ (.D(net452),
    .GATE(net419),
    .Q(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame3_bit28.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1108_ (.D(net453),
    .GATE(net419),
    .Q(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame3_bit27.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1109_ (.D(net454),
    .GATE(net419),
    .Q(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame3_bit26.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1110_ (.D(net455),
    .GATE(net419),
    .Q(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame3_bit25.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1111_ (.D(net456),
    .GATE(net419),
    .Q(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame3_bit24.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1112_ (.D(net202),
    .GATE(net417),
    .Q(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame3_bit23.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1113_ (.D(net201),
    .GATE(net417),
    .Q(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame3_bit22.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1114_ (.D(net200),
    .GATE(net417),
    .Q(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame3_bit21.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1115_ (.D(net199),
    .GATE(net417),
    .Q(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame3_bit20.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1116_ (.D(net461),
    .GATE(net418),
    .Q(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame3_bit19.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1117_ (.D(net462),
    .GATE(net418),
    .Q(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame3_bit18.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1118_ (.D(net463),
    .GATE(net416),
    .Q(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame3_bit17.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1119_ (.D(net464),
    .GATE(net416),
    .Q(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame3_bit16.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1120_ (.D(net465),
    .GATE(net416),
    .Q(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame3_bit15.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1121_ (.D(net466),
    .GATE(net416),
    .Q(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame3_bit14.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1122_ (.D(net193),
    .GATE(net418),
    .Q(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame3_bit13.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1123_ (.D(net192),
    .GATE(net417),
    .Q(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame3_bit12.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1124_ (.D(net191),
    .GATE(net418),
    .Q(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame3_bit11.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1125_ (.D(net190),
    .GATE(net418),
    .Q(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame3_bit10.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1126_ (.D(net218),
    .GATE(net416),
    .Q(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame3_bit9.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1127_ (.D(net217),
    .GATE(net416),
    .Q(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame3_bit8.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1128_ (.D(net216),
    .GATE(net417),
    .Q(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame3_bit7.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1129_ (.D(net215),
    .GATE(net417),
    .Q(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame3_bit6.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1130_ (.D(net214),
    .GATE(net417),
    .Q(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame3_bit5.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1131_ (.D(net213),
    .GATE(net417),
    .Q(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame3_bit4.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1132_ (.D(net212),
    .GATE(net418),
    .Q(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame3_bit3.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1133_ (.D(net209),
    .GATE(net418),
    .Q(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame3_bit2.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1134_ (.D(net198),
    .GATE(net416),
    .Q(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame3_bit1.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1135_ (.D(net189),
    .GATE(net416),
    .Q(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame3_bit0.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1136_ (.D(net211),
    .GATE(net410),
    .Q(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame4_bit31.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1137_ (.D(net210),
    .GATE(net410),
    .Q(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame4_bit30.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1138_ (.D(net451),
    .GATE(net410),
    .Q(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame4_bit29.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1139_ (.D(net452),
    .GATE(net410),
    .Q(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame4_bit28.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1140_ (.D(net453),
    .GATE(net410),
    .Q(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame4_bit27.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1141_ (.D(net454),
    .GATE(net410),
    .Q(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame4_bit26.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1142_ (.D(net455),
    .GATE(net410),
    .Q(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame4_bit25.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1143_ (.D(net456),
    .GATE(net410),
    .Q(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame4_bit24.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1144_ (.D(net457),
    .GATE(net408),
    .Q(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame4_bit23.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1145_ (.D(net458),
    .GATE(net408),
    .Q(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame4_bit22.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1146_ (.D(net459),
    .GATE(net408),
    .Q(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame4_bit21.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1147_ (.D(net460),
    .GATE(net407),
    .Q(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame4_bit20.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1148_ (.D(net461),
    .GATE(net408),
    .Q(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame4_bit19.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1149_ (.D(net462),
    .GATE(net408),
    .Q(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame4_bit18.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1150_ (.D(net463),
    .GATE(net407),
    .Q(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame4_bit17.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1151_ (.D(net464),
    .GATE(net407),
    .Q(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame4_bit16.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1152_ (.D(net465),
    .GATE(net407),
    .Q(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame4_bit15.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1153_ (.D(net466),
    .GATE(net407),
    .Q(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame4_bit14.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1154_ (.D(net193),
    .GATE(net408),
    .Q(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame4_bit13.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1155_ (.D(net192),
    .GATE(net407),
    .Q(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame4_bit12.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1156_ (.D(net191),
    .GATE(net409),
    .Q(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame4_bit11.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1157_ (.D(net190),
    .GATE(net409),
    .Q(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame4_bit10.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1158_ (.D(net218),
    .GATE(net407),
    .Q(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame4_bit9.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1159_ (.D(net217),
    .GATE(net407),
    .Q(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame4_bit8.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1160_ (.D(net216),
    .GATE(net407),
    .Q(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame4_bit7.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1161_ (.D(net215),
    .GATE(net407),
    .Q(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame4_bit6.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1162_ (.D(net214),
    .GATE(net409),
    .Q(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame4_bit5.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1163_ (.D(net213),
    .GATE(net409),
    .Q(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame4_bit4.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1164_ (.D(net212),
    .GATE(net408),
    .Q(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame4_bit3.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1165_ (.D(net209),
    .GATE(net408),
    .Q(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame4_bit2.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1166_ (.D(net198),
    .GATE(net409),
    .Q(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame4_bit1.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1167_ (.D(net189),
    .GATE(net408),
    .Q(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame4_bit0.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1168_ (.D(net449),
    .GATE(net401),
    .Q(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame5_bit31.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1169_ (.D(net450),
    .GATE(net401),
    .Q(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame5_bit30.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1170_ (.D(net451),
    .GATE(net399),
    .Q(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame5_bit29.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1171_ (.D(net452),
    .GATE(net399),
    .Q(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame5_bit28.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1172_ (.D(net453),
    .GATE(net400),
    .Q(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame5_bit27.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1173_ (.D(net454),
    .GATE(net400),
    .Q(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame5_bit26.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1174_ (.D(net455),
    .GATE(net398),
    .Q(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame5_bit25.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1175_ (.D(net456),
    .GATE(net398),
    .Q(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame5_bit24.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1176_ (.D(net457),
    .GATE(net398),
    .Q(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame5_bit23.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1177_ (.D(net458),
    .GATE(net398),
    .Q(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame5_bit22.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1178_ (.D(net459),
    .GATE(net399),
    .Q(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame5_bit21.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1179_ (.D(net460),
    .GATE(net399),
    .Q(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame5_bit20.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1180_ (.D(net461),
    .GATE(net400),
    .Q(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame5_bit19.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1181_ (.D(net462),
    .GATE(net400),
    .Q(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame5_bit18.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1182_ (.D(net463),
    .GATE(net398),
    .Q(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame5_bit17.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1183_ (.D(net464),
    .GATE(net398),
    .Q(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame5_bit16.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1184_ (.D(net465),
    .GATE(net398),
    .Q(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame5_bit15.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1185_ (.D(net466),
    .GATE(net398),
    .Q(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame5_bit14.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1186_ (.D(net193),
    .GATE(net399),
    .Q(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame5_bit13.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1187_ (.D(net192),
    .GATE(net399),
    .Q(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame5_bit12.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1188_ (.D(net191),
    .GATE(net406),
    .Q(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame5_bit11.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1189_ (.D(net190),
    .GATE(net406),
    .Q(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame5_bit10.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1190_ (.D(net218),
    .GATE(net398),
    .Q(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame5_bit9.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1191_ (.D(net217),
    .GATE(net398),
    .Q(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame5_bit8.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1192_ (.D(net216),
    .GATE(net399),
    .Q(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame5_bit7.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1193_ (.D(net215),
    .GATE(net399),
    .Q(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame5_bit6.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1194_ (.D(net214),
    .GATE(net401),
    .Q(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame5_bit5.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1195_ (.D(net213),
    .GATE(net401),
    .Q(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame5_bit4.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1196_ (.D(net212),
    .GATE(net400),
    .Q(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame5_bit3.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1197_ (.D(net209),
    .GATE(net400),
    .Q(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame5_bit2.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1198_ (.D(net198),
    .GATE(net400),
    .Q(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame5_bit1.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1199_ (.D(net189),
    .GATE(net400),
    .Q(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame5_bit0.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1200_ (.D(net449),
    .GATE(net393),
    .Q(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame6_bit31.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1201_ (.D(net450),
    .GATE(net393),
    .Q(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame6_bit30.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1202_ (.D(net451),
    .GATE(net390),
    .Q(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame6_bit29.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1203_ (.D(net452),
    .GATE(net390),
    .Q(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame6_bit28.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1204_ (.D(net453),
    .GATE(net393),
    .Q(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame6_bit27.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1205_ (.D(net454),
    .GATE(net393),
    .Q(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame6_bit26.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1206_ (.D(net455),
    .GATE(net390),
    .Q(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame6_bit25.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1207_ (.D(net456),
    .GATE(net390),
    .Q(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame6_bit24.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1208_ (.D(net457),
    .GATE(net391),
    .Q(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame6_bit23.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1209_ (.D(net458),
    .GATE(net391),
    .Q(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame6_bit22.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1210_ (.D(net459),
    .GATE(net391),
    .Q(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame6_bit21.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1211_ (.D(net460),
    .GATE(net391),
    .Q(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame6_bit20.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1212_ (.D(net461),
    .GATE(net392),
    .Q(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame6_bit19.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1213_ (.D(net462),
    .GATE(net392),
    .Q(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame6_bit18.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1214_ (.D(net463),
    .GATE(net392),
    .Q(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame6_bit17.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1215_ (.D(net464),
    .GATE(net392),
    .Q(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame6_bit16.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1216_ (.D(net465),
    .GATE(net390),
    .Q(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame6_bit15.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1217_ (.D(net466),
    .GATE(net390),
    .Q(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame6_bit14.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1218_ (.D(net193),
    .GATE(net390),
    .Q(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame6_bit13.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1219_ (.D(net192),
    .GATE(net390),
    .Q(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame6_bit12.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1220_ (.D(net191),
    .GATE(net393),
    .Q(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame6_bit11.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1221_ (.D(net190),
    .GATE(net393),
    .Q(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame6_bit10.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1222_ (.D(net218),
    .GATE(net390),
    .Q(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame6_bit9.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1223_ (.D(net217),
    .GATE(net390),
    .Q(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame6_bit8.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1224_ (.D(net216),
    .GATE(net391),
    .Q(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame6_bit7.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1225_ (.D(net215),
    .GATE(net391),
    .Q(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame6_bit6.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1226_ (.D(net214),
    .GATE(net391),
    .Q(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame6_bit5.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1227_ (.D(net213),
    .GATE(net391),
    .Q(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame6_bit4.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1228_ (.D(net212),
    .GATE(net392),
    .Q(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame6_bit3.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1229_ (.D(net209),
    .GATE(net392),
    .Q(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame6_bit2.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1230_ (.D(net198),
    .GATE(net392),
    .Q(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame6_bit1.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1231_ (.D(net189),
    .GATE(net392),
    .Q(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame6_bit0.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1232_ (.D(net449),
    .GATE(net381),
    .Q(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame7_bit31.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1233_ (.D(net450),
    .GATE(net381),
    .Q(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame7_bit30.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1234_ (.D(net451),
    .GATE(net383),
    .Q(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame7_bit29.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1235_ (.D(net452),
    .GATE(net383),
    .Q(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame7_bit28.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1236_ (.D(net453),
    .GATE(net382),
    .Q(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame7_bit27.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1237_ (.D(net454),
    .GATE(net382),
    .Q(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame7_bit26.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1238_ (.D(net455),
    .GATE(net382),
    .Q(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame7_bit25.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1239_ (.D(net456),
    .GATE(net382),
    .Q(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame7_bit24.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1240_ (.D(net457),
    .GATE(net383),
    .Q(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame7_bit23.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1241_ (.D(net458),
    .GATE(net383),
    .Q(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame7_bit22.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1242_ (.D(net459),
    .GATE(net383),
    .Q(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame7_bit21.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1243_ (.D(net460),
    .GATE(net383),
    .Q(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame7_bit20.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1244_ (.D(net461),
    .GATE(net384),
    .Q(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame7_bit19.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1245_ (.D(net462),
    .GATE(net384),
    .Q(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame7_bit18.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1246_ (.D(net463),
    .GATE(net383),
    .Q(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame7_bit17.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1247_ (.D(net464),
    .GATE(net383),
    .Q(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame7_bit16.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1248_ (.D(net195),
    .GATE(net389),
    .Q(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame7_bit15.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1249_ (.D(net194),
    .GATE(net389),
    .Q(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame7_bit14.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1250_ (.D(net193),
    .GATE(net389),
    .Q(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame7_bit13.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1251_ (.D(net192),
    .GATE(net383),
    .Q(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame7_bit12.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1252_ (.D(net191),
    .GATE(net384),
    .Q(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame7_bit11.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1253_ (.D(net190),
    .GATE(net383),
    .Q(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame7_bit10.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1254_ (.D(net218),
    .GATE(net381),
    .Q(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame7_bit9.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1255_ (.D(net217),
    .GATE(net381),
    .Q(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame7_bit8.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1256_ (.D(net216),
    .GATE(net382),
    .Q(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame7_bit7.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1257_ (.D(net215),
    .GATE(net381),
    .Q(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame7_bit6.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1258_ (.D(net214),
    .GATE(net381),
    .Q(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame7_bit5.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1259_ (.D(net213),
    .GATE(net381),
    .Q(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame7_bit4.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1260_ (.D(net212),
    .GATE(net382),
    .Q(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame7_bit3.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1261_ (.D(net209),
    .GATE(net381),
    .Q(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame7_bit2.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1262_ (.D(net198),
    .GATE(net381),
    .Q(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame7_bit1.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1263_ (.D(net189),
    .GATE(net381),
    .Q(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame7_bit0.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1264_ (.D(net449),
    .GATE(net373),
    .Q(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame8_bit31.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1265_ (.D(net450),
    .GATE(net373),
    .Q(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame8_bit30.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1266_ (.D(net451),
    .GATE(net373),
    .Q(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame8_bit29.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1267_ (.D(net452),
    .GATE(net373),
    .Q(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame8_bit28.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1268_ (.D(net453),
    .GATE(net374),
    .Q(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame8_bit27.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1269_ (.D(net454),
    .GATE(net374),
    .Q(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame8_bit26.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1270_ (.D(net455),
    .GATE(net375),
    .Q(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame8_bit25.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1271_ (.D(net456),
    .GATE(net375),
    .Q(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame8_bit24.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1272_ (.D(net457),
    .GATE(net376),
    .Q(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame8_bit23.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1273_ (.D(net458),
    .GATE(net376),
    .Q(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame8_bit22.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1274_ (.D(net459),
    .GATE(net374),
    .Q(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame8_bit21.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1275_ (.D(net460),
    .GATE(net374),
    .Q(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame8_bit20.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1276_ (.D(net461),
    .GATE(net375),
    .Q(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame8_bit19.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1277_ (.D(net462),
    .GATE(net375),
    .Q(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame8_bit18.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1278_ (.D(net463),
    .GATE(net375),
    .Q(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame8_bit17.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1279_ (.D(net464),
    .GATE(net375),
    .Q(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame8_bit16.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1280_ (.D(net465),
    .GATE(net375),
    .Q(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame8_bit15.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1281_ (.D(net466),
    .GATE(net376),
    .Q(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame8_bit14.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1282_ (.D(net193),
    .GATE(net376),
    .Q(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame8_bit13.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1283_ (.D(net192),
    .GATE(net376),
    .Q(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame8_bit12.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1284_ (.D(net191),
    .GATE(net376),
    .Q(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame8_bit11.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1285_ (.D(net190),
    .GATE(net373),
    .Q(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame8_bit10.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1286_ (.D(net218),
    .GATE(net373),
    .Q(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame8_bit9.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1287_ (.D(net217),
    .GATE(net375),
    .Q(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame8_bit8.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1288_ (.D(net216),
    .GATE(net375),
    .Q(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame8_bit7.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1289_ (.D(net215),
    .GATE(net375),
    .Q(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame8_bit6.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1290_ (.D(net214),
    .GATE(net374),
    .Q(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame8_bit5.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1291_ (.D(net213),
    .GATE(net374),
    .Q(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame8_bit4.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1292_ (.D(net212),
    .GATE(net373),
    .Q(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame8_bit3.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1293_ (.D(net209),
    .GATE(net373),
    .Q(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame8_bit2.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1294_ (.D(net198),
    .GATE(net373),
    .Q(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame8_bit1.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1295_ (.D(net189),
    .GATE(net373),
    .Q(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame8_bit0.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1296_ (.D(net449),
    .GATE(net371),
    .Q(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame9_bit31.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1297_ (.D(net450),
    .GATE(net371),
    .Q(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame9_bit30.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1298_ (.D(net451),
    .GATE(net370),
    .Q(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame9_bit29.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1299_ (.D(net452),
    .GATE(net370),
    .Q(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame9_bit28.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1300_ (.D(net453),
    .GATE(net371),
    .Q(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame9_bit27.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1301_ (.D(net454),
    .GATE(net371),
    .Q(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame9_bit26.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1302_ (.D(net455),
    .GATE(net370),
    .Q(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame9_bit25.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1303_ (.D(net456),
    .GATE(net370),
    .Q(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame9_bit24.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1304_ (.D(net457),
    .GATE(net370),
    .Q(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame9_bit23.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1305_ (.D(net458),
    .GATE(net370),
    .Q(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame9_bit22.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1306_ (.D(net459),
    .GATE(net370),
    .Q(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame9_bit21.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1307_ (.D(net460),
    .GATE(net370),
    .Q(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame9_bit20.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1308_ (.D(net461),
    .GATE(net371),
    .Q(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame9_bit19.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1309_ (.D(net462),
    .GATE(net371),
    .Q(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame9_bit18.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1310_ (.D(net463),
    .GATE(net371),
    .Q(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame9_bit17.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1311_ (.D(net464),
    .GATE(net371),
    .Q(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame9_bit16.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1312_ (.D(net465),
    .GATE(net370),
    .Q(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame9_bit15.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1313_ (.D(net466),
    .GATE(net370),
    .Q(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_ConfigMem.Inst_frame9_bit14.Q ));
 sky130_fd_sc_hd__buf_2 _1314_ (.A(clknet_1_0__leaf_Tile_X0Y1_UserCLK),
    .X(net290));
 sky130_fd_sc_hd__buf_1 _1315_ (.A(net81),
    .X(net325));
 sky130_fd_sc_hd__buf_1 _1316_ (.A(net92),
    .X(net336));
 sky130_fd_sc_hd__clkbuf_2 _1317_ (.A(net103),
    .X(net347));
 sky130_fd_sc_hd__clkbuf_2 _1318_ (.A(net106),
    .X(net350));
 sky130_fd_sc_hd__clkbuf_2 _1319_ (.A(net107),
    .X(net351));
 sky130_fd_sc_hd__clkbuf_2 _1320_ (.A(net108),
    .X(net352));
 sky130_fd_sc_hd__buf_1 _1321_ (.A(net109),
    .X(net353));
 sky130_fd_sc_hd__clkbuf_1 _1322_ (.A(net110),
    .X(net354));
 sky130_fd_sc_hd__clkbuf_2 _1323_ (.A(net111),
    .X(net355));
 sky130_fd_sc_hd__clkbuf_2 _1324_ (.A(net112),
    .X(net356));
 sky130_fd_sc_hd__clkbuf_2 _1325_ (.A(net82),
    .X(net326));
 sky130_fd_sc_hd__buf_2 _1326_ (.A(net83),
    .X(net327));
 sky130_fd_sc_hd__buf_1 _1327_ (.A(net84),
    .X(net328));
 sky130_fd_sc_hd__buf_1 _1328_ (.A(net85),
    .X(net329));
 sky130_fd_sc_hd__clkbuf_1 _1329_ (.A(net86),
    .X(net330));
 sky130_fd_sc_hd__buf_1 _1330_ (.A(net87),
    .X(net331));
 sky130_fd_sc_hd__clkbuf_2 _1331_ (.A(net88),
    .X(net332));
 sky130_fd_sc_hd__clkbuf_2 _1332_ (.A(net89),
    .X(net333));
 sky130_fd_sc_hd__clkbuf_2 _1333_ (.A(net90),
    .X(net334));
 sky130_fd_sc_hd__clkbuf_2 _1334_ (.A(net91),
    .X(net335));
 sky130_fd_sc_hd__buf_1 _1335_ (.A(net93),
    .X(net337));
 sky130_fd_sc_hd__clkbuf_2 _1336_ (.A(net94),
    .X(net338));
 sky130_fd_sc_hd__buf_1 _1337_ (.A(net476),
    .X(net339));
 sky130_fd_sc_hd__buf_1 _1338_ (.A(net475),
    .X(net340));
 sky130_fd_sc_hd__clkbuf_2 _1339_ (.A(net474),
    .X(net341));
 sky130_fd_sc_hd__clkbuf_2 _1340_ (.A(net473),
    .X(net342));
 sky130_fd_sc_hd__clkbuf_2 _1341_ (.A(net472),
    .X(net343));
 sky130_fd_sc_hd__clkbuf_2 _1342_ (.A(net471),
    .X(net344));
 sky130_fd_sc_hd__buf_1 _1343_ (.A(net470),
    .X(net345));
 sky130_fd_sc_hd__buf_1 _1344_ (.A(net469),
    .X(net346));
 sky130_fd_sc_hd__buf_1 _1345_ (.A(net468),
    .X(net348));
 sky130_fd_sc_hd__buf_1 _1346_ (.A(net467),
    .X(net349));
 sky130_fd_sc_hd__buf_4 _1347_ (.A(net447),
    .X(net357));
 sky130_fd_sc_hd__clkbuf_2 _1348_ (.A(net437),
    .X(net485));
 sky130_fd_sc_hd__clkbuf_2 _1349_ (.A(net428),
    .X(net486));
 sky130_fd_sc_hd__clkbuf_2 _1350_ (.A(net421),
    .X(net487));
 sky130_fd_sc_hd__clkbuf_2 _1351_ (.A(net414),
    .X(net488));
 sky130_fd_sc_hd__buf_4 _1352_ (.A(net406),
    .X(net489));
 sky130_fd_sc_hd__clkbuf_2 _1353_ (.A(net397),
    .X(net490));
 sky130_fd_sc_hd__clkbuf_1 _1354_ (.A(net387),
    .X(net491));
 sky130_fd_sc_hd__buf_1 _1355_ (.A(net379),
    .X(net492));
 sky130_fd_sc_hd__buf_1 _1356_ (.A(net372),
    .X(net493));
 sky130_fd_sc_hd__clkbuf_1 _1357_ (.A(Tile_X0Y1_FrameStrobe[10]),
    .X(net358));
 sky130_fd_sc_hd__clkbuf_1 _1358_ (.A(Tile_X0Y1_FrameStrobe[11]),
    .X(net359));
 sky130_fd_sc_hd__clkbuf_1 _1359_ (.A(Tile_X0Y1_FrameStrobe[12]),
    .X(net477));
 sky130_fd_sc_hd__clkbuf_1 _1360_ (.A(Tile_X0Y1_FrameStrobe[13]),
    .X(net478));
 sky130_fd_sc_hd__clkbuf_1 _1361_ (.A(Tile_X0Y1_FrameStrobe[14]),
    .X(net479));
 sky130_fd_sc_hd__clkbuf_1 _1362_ (.A(Tile_X0Y1_FrameStrobe[15]),
    .X(net480));
 sky130_fd_sc_hd__clkbuf_1 _1363_ (.A(Tile_X0Y1_FrameStrobe[16]),
    .X(net481));
 sky130_fd_sc_hd__clkbuf_1 _1364_ (.A(Tile_X0Y1_FrameStrobe[17]),
    .X(net482));
 sky130_fd_sc_hd__clkbuf_1 _1365_ (.A(Tile_X0Y1_FrameStrobe[18]),
    .X(net483));
 sky130_fd_sc_hd__clkbuf_1 _1366_ (.A(Tile_X0Y1_FrameStrobe[19]),
    .X(net484));
 sky130_fd_sc_hd__buf_4 _1367_ (.A(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.N1BEG0 ),
    .X(net494));
 sky130_fd_sc_hd__buf_1 _1368_ (.A(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.N1BEG1 ),
    .X(net495));
 sky130_fd_sc_hd__buf_1 _1369_ (.A(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.N1BEG2 ),
    .X(net496));
 sky130_fd_sc_hd__clkbuf_2 _1370_ (.A(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.N1BEG3 ),
    .X(net497));
 sky130_fd_sc_hd__buf_4 _1371_ (.A(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.N2BEG0 ),
    .X(net498));
 sky130_fd_sc_hd__clkbuf_1 _1372_ (.A(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.N2BEG1 ),
    .X(net499));
 sky130_fd_sc_hd__clkbuf_2 _1373_ (.A(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.N2BEG2 ),
    .X(net500));
 sky130_fd_sc_hd__clkbuf_2 _1374_ (.A(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.N2BEG3 ),
    .X(net501));
 sky130_fd_sc_hd__clkbuf_2 _1375_ (.A(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.N2BEG4 ),
    .X(net502));
 sky130_fd_sc_hd__clkbuf_2 _1376_ (.A(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.N2BEG5 ),
    .X(net503));
 sky130_fd_sc_hd__clkbuf_2 _1377_ (.A(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.N2BEG6 ),
    .X(net504));
 sky130_fd_sc_hd__buf_4 _1378_ (.A(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.N2BEG7 ),
    .X(net505));
 sky130_fd_sc_hd__buf_4 _1379_ (.A(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.N2BEGb0 ),
    .X(net506));
 sky130_fd_sc_hd__clkbuf_2 _1380_ (.A(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.N2BEGb1 ),
    .X(net507));
 sky130_fd_sc_hd__clkbuf_2 _1381_ (.A(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.N2BEGb2 ),
    .X(net508));
 sky130_fd_sc_hd__buf_4 _1382_ (.A(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.N2BEGb3 ),
    .X(net509));
 sky130_fd_sc_hd__buf_2 _1383_ (.A(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.N2BEGb4 ),
    .X(net510));
 sky130_fd_sc_hd__clkbuf_2 _1384_ (.A(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.N2BEGb5 ),
    .X(net511));
 sky130_fd_sc_hd__clkbuf_2 _1385_ (.A(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.N2BEGb6 ),
    .X(net512));
 sky130_fd_sc_hd__buf_4 _1386_ (.A(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.N2BEGb7 ),
    .X(net513));
 sky130_fd_sc_hd__buf_4 _1387_ (.A(Tile_X0Y1_N4END[8]),
    .X(net514));
 sky130_fd_sc_hd__buf_4 _1388_ (.A(Tile_X0Y1_N4END[9]),
    .X(net521));
 sky130_fd_sc_hd__buf_4 _1389_ (.A(Tile_X0Y1_N4END[10]),
    .X(net522));
 sky130_fd_sc_hd__buf_4 _1390_ (.A(Tile_X0Y1_N4END[11]),
    .X(net523));
 sky130_fd_sc_hd__buf_4 _1391_ (.A(Tile_X0Y1_N4END[12]),
    .X(net524));
 sky130_fd_sc_hd__buf_4 _1392_ (.A(Tile_X0Y1_N4END[13]),
    .X(net525));
 sky130_fd_sc_hd__buf_4 _1393_ (.A(Tile_X0Y1_N4END[14]),
    .X(net526));
 sky130_fd_sc_hd__buf_4 _1394_ (.A(Tile_X0Y1_N4END[15]),
    .X(net527));
 sky130_fd_sc_hd__buf_4 _1395_ (.A(\Tile_X0Y0_EF_SRAM_top.N4BEG_outbuf_8.A ),
    .X(net528));
 sky130_fd_sc_hd__buf_4 _1396_ (.A(\Tile_X0Y0_EF_SRAM_top.N4BEG_outbuf_9.A ),
    .X(net529));
 sky130_fd_sc_hd__buf_4 _1397_ (.A(\Tile_X0Y0_EF_SRAM_top.N4BEG_outbuf_10.A ),
    .X(net515));
 sky130_fd_sc_hd__buf_4 _1398_ (.A(\Tile_X0Y0_EF_SRAM_top.N4BEG_outbuf_11.A ),
    .X(net516));
 sky130_fd_sc_hd__clkbuf_2 _1399_ (.A(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.N4BEG0 ),
    .X(net517));
 sky130_fd_sc_hd__buf_1 _1400_ (.A(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.N4BEG1 ),
    .X(net518));
 sky130_fd_sc_hd__buf_1 _1401_ (.A(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.N4BEG2 ),
    .X(net519));
 sky130_fd_sc_hd__buf_1 _1402_ (.A(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.N4BEG3 ),
    .X(net520));
 sky130_fd_sc_hd__buf_2 _1403_ (.A(clknet_1_1__leaf_Tile_X0Y1_UserCLK),
    .X(net530));
 sky130_fd_sc_hd__buf_1 _1404_ (.A(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.W1BEG0 ),
    .X(net531));
 sky130_fd_sc_hd__buf_1 _1405_ (.A(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.W1BEG1 ),
    .X(net532));
 sky130_fd_sc_hd__buf_1 _1406_ (.A(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.W1BEG2 ),
    .X(net533));
 sky130_fd_sc_hd__clkbuf_2 _1407_ (.A(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.W1BEG3 ),
    .X(net534));
 sky130_fd_sc_hd__clkbuf_2 _1408_ (.A(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.W2BEG0 ),
    .X(net535));
 sky130_fd_sc_hd__buf_1 _1409_ (.A(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.W2BEG1 ),
    .X(net536));
 sky130_fd_sc_hd__clkbuf_1 _1410_ (.A(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.W2BEG2 ),
    .X(net537));
 sky130_fd_sc_hd__buf_1 _1411_ (.A(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.W2BEG3 ),
    .X(net538));
 sky130_fd_sc_hd__clkbuf_2 _1412_ (.A(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.W2BEG4 ),
    .X(net539));
 sky130_fd_sc_hd__clkbuf_1 _1413_ (.A(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.W2BEG5 ),
    .X(net540));
 sky130_fd_sc_hd__clkbuf_1 _1414_ (.A(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.W2BEG6 ),
    .X(net541));
 sky130_fd_sc_hd__clkbuf_2 _1415_ (.A(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.W2BEG7 ),
    .X(net542));
 sky130_fd_sc_hd__clkbuf_2 _1416_ (.A(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.W2BEGb0 ),
    .X(net543));
 sky130_fd_sc_hd__buf_1 _1417_ (.A(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.W2BEGb1 ),
    .X(net544));
 sky130_fd_sc_hd__clkbuf_1 _1418_ (.A(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.W2BEGb2 ),
    .X(net545));
 sky130_fd_sc_hd__buf_1 _1419_ (.A(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.W2BEGb3 ),
    .X(net546));
 sky130_fd_sc_hd__buf_1 _1420_ (.A(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.W2BEGb4 ),
    .X(net547));
 sky130_fd_sc_hd__buf_1 _1421_ (.A(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.W2BEGb5 ),
    .X(net548));
 sky130_fd_sc_hd__clkbuf_1 _1422_ (.A(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.W2BEGb6 ),
    .X(net549));
 sky130_fd_sc_hd__clkbuf_2 _1423_ (.A(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.W2BEGb7 ),
    .X(net550));
 sky130_fd_sc_hd__buf_1 _1424_ (.A(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.W6BEG0 ),
    .X(net551));
 sky130_fd_sc_hd__buf_1 _1425_ (.A(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.W6BEG1 ),
    .X(net554));
 sky130_fd_sc_hd__clkbuf_1 _1426_ (.A(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.W6BEG2 ),
    .X(net555));
 sky130_fd_sc_hd__buf_1 _1427_ (.A(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.W6BEG3 ),
    .X(net556));
 sky130_fd_sc_hd__clkbuf_2 _1428_ (.A(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.W6BEG4 ),
    .X(net557));
 sky130_fd_sc_hd__buf_1 _1429_ (.A(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.W6BEG5 ),
    .X(net558));
 sky130_fd_sc_hd__clkbuf_1 _1430_ (.A(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.W6BEG6 ),
    .X(net559));
 sky130_fd_sc_hd__buf_1 _1431_ (.A(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.W6BEG7 ),
    .X(net560));
 sky130_fd_sc_hd__buf_1 _1432_ (.A(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.W6BEG8 ),
    .X(net561));
 sky130_fd_sc_hd__clkbuf_1 _1433_ (.A(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.W6BEG9 ),
    .X(net562));
 sky130_fd_sc_hd__clkbuf_1 _1434_ (.A(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.W6BEG10 ),
    .X(net552));
 sky130_fd_sc_hd__clkbuf_2 _1435_ (.A(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.W6BEG11 ),
    .X(net553));
 sky130_fd_sc_hd__clkbuf_2 _1436_ (.A(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.WW4BEG0 ),
    .X(net563));
 sky130_fd_sc_hd__clkbuf_1 _1437_ (.A(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.WW4BEG1 ),
    .X(net570));
 sky130_fd_sc_hd__clkbuf_1 _1438_ (.A(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.WW4BEG2 ),
    .X(net571));
 sky130_fd_sc_hd__clkbuf_2 _1439_ (.A(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.WW4BEG3 ),
    .X(net572));
 sky130_fd_sc_hd__clkbuf_2 _1440_ (.A(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.WW4BEG4 ),
    .X(net573));
 sky130_fd_sc_hd__buf_1 _1441_ (.A(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.WW4BEG5 ),
    .X(net574));
 sky130_fd_sc_hd__clkbuf_1 _1442_ (.A(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.WW4BEG6 ),
    .X(net575));
 sky130_fd_sc_hd__buf_1 _1443_ (.A(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.WW4BEG7 ),
    .X(net576));
 sky130_fd_sc_hd__clkbuf_2 _1444_ (.A(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.WW4BEG8 ),
    .X(net577));
 sky130_fd_sc_hd__buf_1 _1445_ (.A(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.WW4BEG9 ),
    .X(net578));
 sky130_fd_sc_hd__clkbuf_1 _1446_ (.A(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.WW4BEG10 ),
    .X(net564));
 sky130_fd_sc_hd__buf_1 _1447_ (.A(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.WW4BEG11 ),
    .X(net565));
 sky130_fd_sc_hd__clkbuf_2 _1448_ (.A(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.WW4BEG12 ),
    .X(net566));
 sky130_fd_sc_hd__clkbuf_1 _1449_ (.A(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.WW4BEG13 ),
    .X(net567));
 sky130_fd_sc_hd__clkbuf_1 _1450_ (.A(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.WW4BEG14 ),
    .X(net568));
 sky130_fd_sc_hd__clkbuf_2 _1451_ (.A(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.WW4BEG15 ),
    .X(net569));
 sky130_fd_sc_hd__clkbuf_2 _1452_ (.A(net189),
    .X(net579));
 sky130_fd_sc_hd__clkbuf_2 _1453_ (.A(net198),
    .X(net590));
 sky130_fd_sc_hd__buf_4 _1454_ (.A(net209),
    .X(net601));
 sky130_fd_sc_hd__buf_4 _1455_ (.A(net212),
    .X(net604));
 sky130_fd_sc_hd__buf_4 _1456_ (.A(net213),
    .X(net605));
 sky130_fd_sc_hd__buf_4 _1457_ (.A(net214),
    .X(net606));
 sky130_fd_sc_hd__buf_4 _1458_ (.A(net215),
    .X(net607));
 sky130_fd_sc_hd__buf_4 _1459_ (.A(net216),
    .X(net608));
 sky130_fd_sc_hd__buf_4 _1460_ (.A(net217),
    .X(net609));
 sky130_fd_sc_hd__buf_4 _1461_ (.A(net218),
    .X(net610));
 sky130_fd_sc_hd__buf_4 _1462_ (.A(net190),
    .X(net580));
 sky130_fd_sc_hd__buf_4 _1463_ (.A(net191),
    .X(net581));
 sky130_fd_sc_hd__buf_4 _1464_ (.A(net192),
    .X(net582));
 sky130_fd_sc_hd__buf_4 _1465_ (.A(net193),
    .X(net583));
 sky130_fd_sc_hd__buf_4 _1466_ (.A(net466),
    .X(net584));
 sky130_fd_sc_hd__buf_4 _1467_ (.A(net465),
    .X(net585));
 sky130_fd_sc_hd__clkbuf_2 _1468_ (.A(Tile_X0Y1_FrameData[16]),
    .X(net586));
 sky130_fd_sc_hd__buf_4 _1469_ (.A(Tile_X0Y1_FrameData[17]),
    .X(net587));
 sky130_fd_sc_hd__buf_4 _1470_ (.A(net462),
    .X(net588));
 sky130_fd_sc_hd__buf_4 _1471_ (.A(net461),
    .X(net589));
 sky130_fd_sc_hd__buf_4 _1472_ (.A(net460),
    .X(net591));
 sky130_fd_sc_hd__buf_4 _1473_ (.A(net459),
    .X(net592));
 sky130_fd_sc_hd__buf_4 _1474_ (.A(net458),
    .X(net593));
 sky130_fd_sc_hd__buf_4 _1475_ (.A(net457),
    .X(net594));
 sky130_fd_sc_hd__buf_4 _1476_ (.A(net456),
    .X(net595));
 sky130_fd_sc_hd__buf_4 _1477_ (.A(net455),
    .X(net596));
 sky130_fd_sc_hd__buf_4 _1478_ (.A(net454),
    .X(net597));
 sky130_fd_sc_hd__buf_4 _1479_ (.A(net453),
    .X(net598));
 sky130_fd_sc_hd__buf_4 _1480_ (.A(net452),
    .X(net599));
 sky130_fd_sc_hd__buf_4 _1481_ (.A(net451),
    .X(net600));
 sky130_fd_sc_hd__buf_2 _1482_ (.A(net450),
    .X(net602));
 sky130_fd_sc_hd__buf_2 _1483_ (.A(net449),
    .X(net603));
 sky130_fd_sc_hd__clkbuf_2 _1484_ (.A(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.S1BEG0 ),
    .X(net611));
 sky130_fd_sc_hd__clkbuf_2 _1485_ (.A(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.S1BEG1 ),
    .X(net612));
 sky130_fd_sc_hd__buf_1 _1486_ (.A(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.S1BEG2 ),
    .X(net613));
 sky130_fd_sc_hd__buf_1 _1487_ (.A(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.S1BEG3 ),
    .X(net614));
 sky130_fd_sc_hd__clkbuf_2 _1488_ (.A(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.S2BEG0 ),
    .X(net615));
 sky130_fd_sc_hd__clkbuf_2 _1489_ (.A(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.S2BEG1 ),
    .X(net616));
 sky130_fd_sc_hd__clkbuf_2 _1490_ (.A(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.S2BEG2 ),
    .X(net617));
 sky130_fd_sc_hd__clkbuf_2 _1491_ (.A(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.S2BEG3 ),
    .X(net618));
 sky130_fd_sc_hd__clkbuf_2 _1492_ (.A(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.S2BEG4 ),
    .X(net619));
 sky130_fd_sc_hd__clkbuf_2 _1493_ (.A(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.S2BEG5 ),
    .X(net620));
 sky130_fd_sc_hd__clkbuf_2 _1494_ (.A(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.S2BEG6 ),
    .X(net621));
 sky130_fd_sc_hd__buf_1 _1495_ (.A(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.S2BEG7 ),
    .X(net622));
 sky130_fd_sc_hd__clkbuf_2 _1496_ (.A(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.S2BEG0 ),
    .X(net623));
 sky130_fd_sc_hd__buf_4 _1497_ (.A(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.S2BEG1 ),
    .X(net624));
 sky130_fd_sc_hd__clkbuf_2 _1498_ (.A(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.S2BEG2 ),
    .X(net625));
 sky130_fd_sc_hd__clkbuf_2 _1499_ (.A(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.S2BEG3 ),
    .X(net626));
 sky130_fd_sc_hd__clkbuf_2 _1500_ (.A(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.S2BEG4 ),
    .X(net627));
 sky130_fd_sc_hd__buf_2 _1501_ (.A(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.S2BEG5 ),
    .X(net628));
 sky130_fd_sc_hd__clkbuf_2 _1502_ (.A(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.S2BEG6 ),
    .X(net629));
 sky130_fd_sc_hd__clkbuf_2 _1503_ (.A(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.S2BEG7 ),
    .X(net630));
 sky130_fd_sc_hd__buf_4 _1504_ (.A(Tile_X0Y0_S4END[8]),
    .X(net631));
 sky130_fd_sc_hd__buf_4 _1505_ (.A(Tile_X0Y0_S4END[9]),
    .X(net638));
 sky130_fd_sc_hd__buf_4 _1506_ (.A(Tile_X0Y0_S4END[10]),
    .X(net639));
 sky130_fd_sc_hd__buf_4 _1507_ (.A(Tile_X0Y0_S4END[11]),
    .X(net640));
 sky130_fd_sc_hd__buf_4 _1508_ (.A(Tile_X0Y0_S4END[12]),
    .X(net641));
 sky130_fd_sc_hd__buf_4 _1509_ (.A(Tile_X0Y0_S4END[13]),
    .X(net642));
 sky130_fd_sc_hd__buf_4 _1510_ (.A(Tile_X0Y0_S4END[14]),
    .X(net643));
 sky130_fd_sc_hd__buf_4 _1511_ (.A(Tile_X0Y0_S4END[15]),
    .X(net644));
 sky130_fd_sc_hd__buf_4 _1512_ (.A(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.S4BEG0 ),
    .X(net645));
 sky130_fd_sc_hd__buf_4 _1513_ (.A(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.S4BEG1 ),
    .X(net646));
 sky130_fd_sc_hd__buf_4 _1514_ (.A(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.S4BEG2 ),
    .X(net632));
 sky130_fd_sc_hd__buf_4 _1515_ (.A(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.S4BEG3 ),
    .X(net633));
 sky130_fd_sc_hd__buf_1 _1516_ (.A(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.S4BEG0 ),
    .X(net634));
 sky130_fd_sc_hd__buf_4 _1517_ (.A(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.S4BEG1 ),
    .X(net635));
 sky130_fd_sc_hd__buf_1 _1518_ (.A(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.S4BEG2 ),
    .X(net636));
 sky130_fd_sc_hd__buf_1 _1519_ (.A(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.S4BEG3 ),
    .X(net637));
 sky130_fd_sc_hd__clkbuf_2 _1520_ (.A(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.W1BEG0 ),
    .X(net647));
 sky130_fd_sc_hd__clkbuf_1 _1521_ (.A(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.W1BEG1 ),
    .X(net648));
 sky130_fd_sc_hd__buf_1 _1522_ (.A(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.W1BEG2 ),
    .X(net649));
 sky130_fd_sc_hd__clkbuf_2 _1523_ (.A(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.W1BEG3 ),
    .X(net650));
 sky130_fd_sc_hd__clkbuf_2 _1524_ (.A(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.W2BEG0 ),
    .X(net651));
 sky130_fd_sc_hd__buf_1 _1525_ (.A(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.W2BEG1 ),
    .X(net652));
 sky130_fd_sc_hd__buf_1 _1526_ (.A(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.W2BEG2 ),
    .X(net653));
 sky130_fd_sc_hd__buf_1 _1527_ (.A(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.W2BEG3 ),
    .X(net654));
 sky130_fd_sc_hd__buf_1 _1528_ (.A(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.W2BEG4 ),
    .X(net655));
 sky130_fd_sc_hd__buf_1 _1529_ (.A(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.W2BEG5 ),
    .X(net656));
 sky130_fd_sc_hd__buf_1 _1530_ (.A(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.W2BEG6 ),
    .X(net657));
 sky130_fd_sc_hd__buf_1 _1531_ (.A(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.W2BEG7 ),
    .X(net658));
 sky130_fd_sc_hd__buf_1 _1532_ (.A(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.W2BEGb0 ),
    .X(net659));
 sky130_fd_sc_hd__clkbuf_1 _1533_ (.A(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.W2BEGb1 ),
    .X(net660));
 sky130_fd_sc_hd__buf_1 _1534_ (.A(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.W2BEGb2 ),
    .X(net661));
 sky130_fd_sc_hd__buf_1 _1535_ (.A(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.W2BEGb3 ),
    .X(net662));
 sky130_fd_sc_hd__buf_1 _1536_ (.A(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.W2BEGb4 ),
    .X(net663));
 sky130_fd_sc_hd__buf_1 _1537_ (.A(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.W2BEGb5 ),
    .X(net664));
 sky130_fd_sc_hd__buf_1 _1538_ (.A(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.W2BEGb6 ),
    .X(net665));
 sky130_fd_sc_hd__buf_1 _1539_ (.A(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.W2BEGb7 ),
    .X(net666));
 sky130_fd_sc_hd__clkbuf_2 _1540_ (.A(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.W6BEG0 ),
    .X(net667));
 sky130_fd_sc_hd__buf_1 _1541_ (.A(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.W6BEG1 ),
    .X(net670));
 sky130_fd_sc_hd__buf_1 _1542_ (.A(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.W6BEG2 ),
    .X(net671));
 sky130_fd_sc_hd__buf_1 _1543_ (.A(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.W6BEG3 ),
    .X(net672));
 sky130_fd_sc_hd__clkbuf_2 _1544_ (.A(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.W6BEG4 ),
    .X(net673));
 sky130_fd_sc_hd__buf_1 _1545_ (.A(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.W6BEG5 ),
    .X(net674));
 sky130_fd_sc_hd__clkbuf_1 _1546_ (.A(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.W6BEG6 ),
    .X(net675));
 sky130_fd_sc_hd__clkbuf_1 _1547_ (.A(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.W6BEG7 ),
    .X(net676));
 sky130_fd_sc_hd__clkbuf_2 _1548_ (.A(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.W6BEG8 ),
    .X(net677));
 sky130_fd_sc_hd__buf_1 _1549_ (.A(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.W6BEG9 ),
    .X(net678));
 sky130_fd_sc_hd__clkbuf_1 _1550_ (.A(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.W6BEG10 ),
    .X(net668));
 sky130_fd_sc_hd__buf_1 _1551_ (.A(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.W6BEG11 ),
    .X(net669));
 sky130_fd_sc_hd__clkbuf_2 _1552_ (.A(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.WW4BEG0 ),
    .X(net679));
 sky130_fd_sc_hd__buf_1 _1553_ (.A(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.WW4BEG1 ),
    .X(net686));
 sky130_fd_sc_hd__buf_1 _1554_ (.A(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.WW4BEG2 ),
    .X(net687));
 sky130_fd_sc_hd__clkbuf_1 _1555_ (.A(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.WW4BEG3 ),
    .X(net688));
 sky130_fd_sc_hd__buf_1 _1556_ (.A(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.WW4BEG4 ),
    .X(net689));
 sky130_fd_sc_hd__buf_1 _1557_ (.A(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.WW4BEG5 ),
    .X(net690));
 sky130_fd_sc_hd__buf_1 _1558_ (.A(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.WW4BEG6 ),
    .X(net691));
 sky130_fd_sc_hd__buf_1 _1559_ (.A(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.WW4BEG7 ),
    .X(net692));
 sky130_fd_sc_hd__buf_1 _1560_ (.A(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.WW4BEG8 ),
    .X(net693));
 sky130_fd_sc_hd__buf_1 _1561_ (.A(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.WW4BEG9 ),
    .X(net694));
 sky130_fd_sc_hd__clkbuf_1 _1562_ (.A(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.WW4BEG10 ),
    .X(net680));
 sky130_fd_sc_hd__buf_1 _1563_ (.A(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.WW4BEG11 ),
    .X(net681));
 sky130_fd_sc_hd__buf_1 _1564_ (.A(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.WW4BEG12 ),
    .X(net682));
 sky130_fd_sc_hd__buf_1 _1565_ (.A(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.WW4BEG13 ),
    .X(net683));
 sky130_fd_sc_hd__clkbuf_1 _1566_ (.A(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.WW4BEG14 ),
    .X(net684));
 sky130_fd_sc_hd__buf_1 _1567_ (.A(\Tile_X0Y1_EF_SRAM_bot.Inst_EF_SRAM_bot_switch_matrix.WW4BEG15 ),
    .X(net685));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_0_Right_0 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_1_Right_1 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_2_Right_2 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_3_Right_3 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_4_Right_4 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_5_Right_5 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_6_Right_6 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_7_Right_7 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_8_Right_8 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_9_Right_9 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_10_Right_10 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_11_Right_11 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_12_Right_12 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_13_Right_13 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_14_Right_14 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_15_Right_15 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_16_Right_16 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_17_Right_17 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_18_Right_18 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_19_Right_19 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_20_Right_20 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_21_Right_21 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_22_Right_22 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_23_Right_23 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_24_Right_24 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_25_Right_25 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_26_Right_26 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_27_Right_27 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_28_Right_28 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_29_Right_29 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_30_Right_30 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_31_Right_31 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_32_Right_32 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_33_Right_33 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_34_Right_34 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_35_Right_35 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_36_Right_36 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_37_Right_37 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_38_Right_38 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_39_Right_39 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_40_Right_40 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_41_Right_41 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_42_Right_42 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_43_Right_43 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_44_Right_44 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_45_Right_45 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_46_Right_46 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_47_Right_47 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_48_Right_48 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_49_Right_49 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_50_Right_50 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_51_Right_51 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_52_Right_52 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_53_Right_53 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_54_Right_54 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_55_Right_55 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_56_Right_56 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_57_Right_57 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_58_Right_58 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_59_Right_59 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_60_Right_60 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_61_Right_61 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_62_Right_62 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_63_Right_63 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_64_Right_64 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_65_Right_65 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_66_Right_66 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_67_Right_67 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_68_Right_68 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_69_Right_69 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_70_Right_70 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_71_Right_71 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_72_Right_72 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_73_Right_73 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_74_Right_74 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_75_Right_75 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_76_Right_76 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_77_Right_77 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_78_Right_78 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_79_Right_79 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_80_Right_80 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_81_Right_81 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_82_Right_82 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_83_Right_83 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_84_Right_84 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_85_Right_85 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_86_Right_86 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_87_Right_87 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_88_Right_88 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_89_Right_89 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_90_Right_90 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_91_Right_91 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_92_Right_92 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_93_Right_93 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_94_Right_94 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_95_Right_95 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_96_Right_96 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_97_Right_97 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_98_Right_98 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_99_Right_99 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_100_Right_100 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_101_Right_101 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_102_Right_102 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_103_Right_103 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_104_Right_104 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_105_Right_105 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_106_Right_106 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_107_Right_107 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_108_Right_108 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_109_Right_109 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_110_Right_110 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_111_Right_111 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_112_Right_112 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_113_Right_113 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_114_Right_114 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_115_Right_115 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_116_Right_116 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_117_Right_117 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_118_Right_118 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_119_Right_119 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_120_Right_120 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_121_Right_121 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_122_Right_122 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_123_Right_123 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_124_Right_124 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_125_Right_125 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_126_Right_126 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_127_Right_127 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_128_Right_128 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_129_Right_129 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_130_Right_130 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_131_Right_131 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_132_Right_132 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_133_Right_133 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_134_Right_134 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_135_Right_135 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_136_Right_136 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_137_Right_137 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_138_Right_138 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_139_Right_139 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_140_Right_140 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_141_Right_141 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_142_Right_142 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_143_Right_143 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_144_Right_144 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_145_Right_145 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_146_Right_146 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_147_Right_147 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_148_Right_148 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_149_Right_149 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_150_Right_150 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_151_Right_151 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_152_Right_152 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_153_Right_153 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_154_Right_154 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_155_Right_155 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_156_Right_156 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_0_Left_157 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_1_Left_158 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_2_Left_159 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_3_Left_160 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_4_Left_161 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_5_Left_162 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_6_Left_163 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_7_Left_164 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_8_Left_165 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_9_Left_166 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_10_Left_167 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_11_Left_168 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_12_Left_169 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_13_Left_170 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_14_Left_171 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_15_Left_172 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_16_Left_173 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_17_Left_174 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_18_Left_175 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_19_Left_176 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_20_Left_177 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_21_Left_178 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_22_Left_179 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_23_Left_180 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_24_Left_181 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_25_Left_182 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_26_Left_183 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_27_Left_184 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_28_Left_185 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_29_Left_186 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_30_Left_187 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_31_Left_188 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_32_Left_189 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_33_Left_190 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_34_Left_191 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_35_Left_192 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_36_Left_193 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_37_Left_194 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_38_Left_195 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_39_Left_196 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_40_Left_197 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_41_Left_198 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_42_Left_199 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_43_Left_200 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_44_Left_201 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_45_Left_202 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_46_Left_203 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_47_Left_204 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_48_Left_205 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_49_Left_206 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_50_Left_207 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_51_Left_208 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_52_Left_209 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_53_Left_210 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_54_Left_211 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_55_Left_212 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_56_Left_213 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_57_Left_214 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_58_Left_215 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_59_Left_216 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_60_Left_217 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_61_Left_218 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_62_Left_219 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_63_Left_220 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_64_Left_221 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_65_Left_222 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_66_Left_223 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_67_Left_224 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_68_Left_225 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_69_Left_226 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_70_Left_227 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_71_Left_228 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_72_Left_229 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_73_Left_230 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_74_Left_231 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_75_Left_232 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_76_Left_233 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_77_Left_234 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_78_Left_235 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_79_Left_236 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_80_Left_237 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_81_Left_238 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_82_Left_239 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_83_Left_240 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_84_Left_241 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_85_Left_242 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_86_Left_243 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_87_Left_244 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_88_Left_245 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_89_Left_246 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_90_Left_247 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_91_Left_248 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_92_Left_249 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_93_Left_250 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_94_Left_251 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_95_Left_252 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_96_Left_253 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_97_Left_254 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_98_Left_255 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_99_Left_256 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_100_Left_257 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_101_Left_258 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_102_Left_259 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_103_Left_260 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_104_Left_261 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_105_Left_262 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_106_Left_263 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_107_Left_264 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_108_Left_265 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_109_Left_266 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_110_Left_267 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_111_Left_268 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_112_Left_269 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_113_Left_270 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_114_Left_271 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_115_Left_272 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_116_Left_273 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_117_Left_274 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_118_Left_275 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_119_Left_276 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_120_Left_277 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_121_Left_278 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_122_Left_279 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_123_Left_280 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_124_Left_281 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_125_Left_282 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_126_Left_283 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_127_Left_284 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_128_Left_285 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_129_Left_286 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_130_Left_287 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_131_Left_288 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_132_Left_289 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_133_Left_290 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_134_Left_291 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_135_Left_292 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_136_Left_293 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_137_Left_294 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_138_Left_295 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_139_Left_296 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_140_Left_297 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_141_Left_298 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_142_Left_299 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_143_Left_300 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_144_Left_301 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_145_Left_302 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_146_Left_303 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_147_Left_304 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_148_Left_305 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_149_Left_306 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_150_Left_307 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_151_Left_308 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_152_Left_309 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_153_Left_310 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_154_Left_311 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_155_Left_312 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_156_Left_313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_1000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_1001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_1002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_1003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_1004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_1005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_1006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_1007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_1008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_1009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_1010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_1011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_1012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_1013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_1014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_1015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_1016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_1017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_1018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_1019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_1020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_1021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_1022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_1023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_1024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_1025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_1026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_1027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_1028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_1029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_1030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_1031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_1032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_1033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_1034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_1035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_1036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_1037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_1038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_1039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_1040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_1041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_1042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_1043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_1044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_1045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_1046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_1047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_1048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_1049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_1050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_1051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_1052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_1053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_1054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_1055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_1056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_1057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_1058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_1059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_1060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_1061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_1062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_1063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_1064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_1065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_1066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_1067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_1068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_1069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_1070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_1071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_1072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_1073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_1074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_1075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_1076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_1077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_1078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_1079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_1080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_1081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_1082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_1083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_1084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_1085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_1086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_1087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_1088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_1089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_1090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_1091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_1092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_1093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_1094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_1095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_1096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_1097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_1098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_1099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_1100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_1101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_1102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_1103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_1104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_1105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_1106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_1107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_1108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_1109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_1110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_1111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_1112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_1113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_1114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_1115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_1116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_1117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_1118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_1119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_1120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_1121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_1122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_1123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_1124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_1125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_1126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_1127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_1128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_1129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_1130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_1131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_1132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_1133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_1134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_1135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_1136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_1137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_1138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_1139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_1140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_1141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_1142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_1143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_1144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_1145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_1146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_1147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_1148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_1149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_1150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_1151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_1152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_1153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_1154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_1155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_1156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_1157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_1158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_1159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_1160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_1161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_1162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_1163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_1164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_1165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_1166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_1167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_1168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_1169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_1170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_1171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_1172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_1173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_1174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_1175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_1176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_1177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_1178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_1179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_1180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_1181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_1182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_1183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_1184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_1185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_1186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_1187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_1188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_1189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_1190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_1191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_1192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_1193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_1194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_1195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_1196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_1197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_1198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_1199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_1200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_1201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_1202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_1203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_1204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_1205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_1206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_1207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_1208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_1209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_1210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_1211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_1212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_1213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_1214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_1215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_1216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_1217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_1218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_1219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_1220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_1221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_1222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_1223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_1224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_1225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_1226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_1227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_1228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_1229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_1230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_1231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_1232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_1233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_1234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_1235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_1236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_1237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_1238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_1239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_1240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_1241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_1242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_1243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_1244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_1245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_1246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_1247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_1248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_1249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_1250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_1251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_1252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_1253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_1254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_1255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_1256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_1257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_1258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_1259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_1260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_1261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_1262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_1263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_1264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_1265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_1266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_1267 ();
 sky130_fd_sc_hd__buf_2 fanout360 (.A(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.J_NS2_BEG4 ),
    .X(net360));
 sky130_fd_sc_hd__buf_2 fanout361 (.A(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.J_NS2_BEG3 ),
    .X(net361));
 sky130_fd_sc_hd__clkbuf_4 fanout362 (.A(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.J_NS2_BEG2 ),
    .X(net362));
 sky130_fd_sc_hd__buf_2 fanout363 (.A(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.J_NS2_BEG1 ),
    .X(net363));
 sky130_fd_sc_hd__buf_2 fanout364 (.A(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.J_NS2_BEG0 ),
    .X(net364));
 sky130_fd_sc_hd__clkbuf_4 fanout365 (.A(_0080_),
    .X(net365));
 sky130_fd_sc_hd__buf_2 fanout366 (.A(_0079_),
    .X(net366));
 sky130_fd_sc_hd__buf_2 fanout367 (.A(_0078_),
    .X(net367));
 sky130_fd_sc_hd__clkbuf_4 fanout368 (.A(_0077_),
    .X(net368));
 sky130_fd_sc_hd__clkbuf_4 fanout369 (.A(_0076_),
    .X(net369));
 sky130_fd_sc_hd__buf_2 fanout370 (.A(net219),
    .X(net370));
 sky130_fd_sc_hd__clkbuf_2 fanout371 (.A(net219),
    .X(net371));
 sky130_fd_sc_hd__buf_2 fanout372 (.A(net219),
    .X(net372));
 sky130_fd_sc_hd__clkbuf_2 fanout373 (.A(net374),
    .X(net373));
 sky130_fd_sc_hd__clkbuf_2 fanout374 (.A(net376),
    .X(net374));
 sky130_fd_sc_hd__clkbuf_2 fanout375 (.A(net376),
    .X(net375));
 sky130_fd_sc_hd__buf_2 fanout376 (.A(Tile_X0Y1_FrameStrobe[8]),
    .X(net376));
 sky130_fd_sc_hd__clkbuf_4 fanout377 (.A(net379),
    .X(net377));
 sky130_fd_sc_hd__buf_2 fanout378 (.A(net379),
    .X(net378));
 sky130_fd_sc_hd__clkbuf_2 fanout379 (.A(net380),
    .X(net379));
 sky130_fd_sc_hd__buf_2 fanout380 (.A(Tile_X0Y1_FrameStrobe[8]),
    .X(net380));
 sky130_fd_sc_hd__buf_2 fanout381 (.A(net384),
    .X(net381));
 sky130_fd_sc_hd__clkbuf_2 fanout382 (.A(net384),
    .X(net382));
 sky130_fd_sc_hd__clkbuf_2 fanout383 (.A(net384),
    .X(net383));
 sky130_fd_sc_hd__clkbuf_2 fanout384 (.A(net389),
    .X(net384));
 sky130_fd_sc_hd__buf_2 fanout385 (.A(net387),
    .X(net385));
 sky130_fd_sc_hd__buf_2 fanout386 (.A(net387),
    .X(net386));
 sky130_fd_sc_hd__clkbuf_2 fanout387 (.A(net388),
    .X(net387));
 sky130_fd_sc_hd__buf_2 fanout388 (.A(net389),
    .X(net388));
 sky130_fd_sc_hd__clkbuf_2 fanout389 (.A(Tile_X0Y1_FrameStrobe[7]),
    .X(net389));
 sky130_fd_sc_hd__clkbuf_2 fanout390 (.A(net392),
    .X(net390));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout391 (.A(net392),
    .X(net391));
 sky130_fd_sc_hd__buf_2 fanout392 (.A(net393),
    .X(net392));
 sky130_fd_sc_hd__clkbuf_4 fanout393 (.A(Tile_X0Y1_FrameStrobe[6]),
    .X(net393));
 sky130_fd_sc_hd__buf_2 fanout394 (.A(net395),
    .X(net394));
 sky130_fd_sc_hd__buf_2 fanout395 (.A(net397),
    .X(net395));
 sky130_fd_sc_hd__buf_2 fanout396 (.A(net397),
    .X(net396));
 sky130_fd_sc_hd__clkbuf_2 fanout397 (.A(Tile_X0Y1_FrameStrobe[6]),
    .X(net397));
 sky130_fd_sc_hd__clkbuf_2 fanout398 (.A(net400),
    .X(net398));
 sky130_fd_sc_hd__clkbuf_2 fanout399 (.A(net400),
    .X(net399));
 sky130_fd_sc_hd__buf_2 fanout400 (.A(net401),
    .X(net400));
 sky130_fd_sc_hd__clkbuf_2 fanout401 (.A(net406),
    .X(net401));
 sky130_fd_sc_hd__clkbuf_4 fanout402 (.A(net404),
    .X(net402));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout403 (.A(net404),
    .X(net403));
 sky130_fd_sc_hd__buf_2 fanout404 (.A(net406),
    .X(net404));
 sky130_fd_sc_hd__buf_2 fanout405 (.A(net406),
    .X(net405));
 sky130_fd_sc_hd__clkbuf_2 fanout406 (.A(Tile_X0Y1_FrameStrobe[5]),
    .X(net406));
 sky130_fd_sc_hd__clkbuf_2 fanout407 (.A(net408),
    .X(net407));
 sky130_fd_sc_hd__buf_2 fanout408 (.A(net409),
    .X(net408));
 sky130_fd_sc_hd__clkbuf_2 fanout409 (.A(net410),
    .X(net409));
 sky130_fd_sc_hd__buf_2 fanout410 (.A(Tile_X0Y1_FrameStrobe[4]),
    .X(net410));
 sky130_fd_sc_hd__clkbuf_2 fanout411 (.A(net412),
    .X(net411));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout412 (.A(net413),
    .X(net412));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout413 (.A(net414),
    .X(net413));
 sky130_fd_sc_hd__clkbuf_2 fanout414 (.A(Tile_X0Y1_FrameStrobe[4]),
    .X(net414));
 sky130_fd_sc_hd__buf_2 fanout415 (.A(Tile_X0Y1_FrameStrobe[4]),
    .X(net415));
 sky130_fd_sc_hd__clkbuf_2 fanout416 (.A(net419),
    .X(net416));
 sky130_fd_sc_hd__clkbuf_2 fanout417 (.A(net418),
    .X(net417));
 sky130_fd_sc_hd__clkbuf_2 fanout418 (.A(net419),
    .X(net418));
 sky130_fd_sc_hd__buf_2 fanout419 (.A(Tile_X0Y1_FrameStrobe[3]),
    .X(net419));
 sky130_fd_sc_hd__buf_2 fanout420 (.A(net423),
    .X(net420));
 sky130_fd_sc_hd__buf_2 fanout421 (.A(net423),
    .X(net421));
 sky130_fd_sc_hd__clkbuf_2 fanout422 (.A(net423),
    .X(net422));
 sky130_fd_sc_hd__buf_2 fanout423 (.A(Tile_X0Y1_FrameStrobe[3]),
    .X(net423));
 sky130_fd_sc_hd__clkbuf_2 fanout424 (.A(net425),
    .X(net424));
 sky130_fd_sc_hd__buf_2 fanout425 (.A(net426),
    .X(net425));
 sky130_fd_sc_hd__buf_2 fanout426 (.A(net431),
    .X(net426));
 sky130_fd_sc_hd__clkbuf_4 fanout427 (.A(net429),
    .X(net427));
 sky130_fd_sc_hd__buf_2 fanout428 (.A(net429),
    .X(net428));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout429 (.A(net431),
    .X(net429));
 sky130_fd_sc_hd__buf_2 fanout430 (.A(net431),
    .X(net430));
 sky130_fd_sc_hd__clkbuf_4 fanout431 (.A(Tile_X0Y1_FrameStrobe[2]),
    .X(net431));
 sky130_fd_sc_hd__clkbuf_2 fanout432 (.A(net433),
    .X(net432));
 sky130_fd_sc_hd__clkbuf_2 fanout433 (.A(net434),
    .X(net433));
 sky130_fd_sc_hd__clkbuf_2 fanout434 (.A(net435),
    .X(net434));
 sky130_fd_sc_hd__buf_2 fanout435 (.A(Tile_X0Y1_FrameStrobe[1]),
    .X(net435));
 sky130_fd_sc_hd__clkbuf_4 fanout436 (.A(net437),
    .X(net436));
 sky130_fd_sc_hd__clkbuf_2 fanout437 (.A(net439),
    .X(net437));
 sky130_fd_sc_hd__clkbuf_2 fanout438 (.A(Tile_X0Y1_FrameStrobe[1]),
    .X(net438));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout439 (.A(Tile_X0Y1_FrameStrobe[1]),
    .X(net439));
 sky130_fd_sc_hd__buf_2 fanout440 (.A(net443),
    .X(net440));
 sky130_fd_sc_hd__clkbuf_4 fanout441 (.A(net443),
    .X(net441));
 sky130_fd_sc_hd__buf_2 fanout442 (.A(net443),
    .X(net442));
 sky130_fd_sc_hd__clkbuf_2 fanout443 (.A(Tile_X0Y1_FrameStrobe[0]),
    .X(net443));
 sky130_fd_sc_hd__clkbuf_2 fanout444 (.A(net445),
    .X(net444));
 sky130_fd_sc_hd__buf_1 fanout445 (.A(net448),
    .X(net445));
 sky130_fd_sc_hd__buf_2 fanout446 (.A(net448),
    .X(net446));
 sky130_fd_sc_hd__clkbuf_2 fanout447 (.A(net448),
    .X(net447));
 sky130_fd_sc_hd__clkbuf_2 fanout448 (.A(Tile_X0Y1_FrameStrobe[0]),
    .X(net448));
 sky130_fd_sc_hd__buf_4 fanout449 (.A(net211),
    .X(net449));
 sky130_fd_sc_hd__buf_4 fanout450 (.A(net210),
    .X(net450));
 sky130_fd_sc_hd__clkbuf_4 fanout451 (.A(net208),
    .X(net451));
 sky130_fd_sc_hd__clkbuf_4 fanout452 (.A(net207),
    .X(net452));
 sky130_fd_sc_hd__clkbuf_4 fanout453 (.A(net206),
    .X(net453));
 sky130_fd_sc_hd__clkbuf_4 fanout454 (.A(net205),
    .X(net454));
 sky130_fd_sc_hd__buf_4 fanout455 (.A(net204),
    .X(net455));
 sky130_fd_sc_hd__buf_4 fanout456 (.A(net203),
    .X(net456));
 sky130_fd_sc_hd__clkbuf_4 fanout457 (.A(net202),
    .X(net457));
 sky130_fd_sc_hd__clkbuf_4 fanout458 (.A(net201),
    .X(net458));
 sky130_fd_sc_hd__clkbuf_4 fanout459 (.A(net200),
    .X(net459));
 sky130_fd_sc_hd__clkbuf_4 fanout460 (.A(net199),
    .X(net460));
 sky130_fd_sc_hd__clkbuf_4 fanout461 (.A(net197),
    .X(net461));
 sky130_fd_sc_hd__clkbuf_4 fanout462 (.A(net196),
    .X(net462));
 sky130_fd_sc_hd__buf_4 fanout463 (.A(Tile_X0Y1_FrameData[17]),
    .X(net463));
 sky130_fd_sc_hd__buf_4 fanout464 (.A(Tile_X0Y1_FrameData[16]),
    .X(net464));
 sky130_fd_sc_hd__clkbuf_4 fanout465 (.A(net195),
    .X(net465));
 sky130_fd_sc_hd__buf_4 fanout466 (.A(net194),
    .X(net466));
 sky130_fd_sc_hd__buf_2 fanout467 (.A(net105),
    .X(net467));
 sky130_fd_sc_hd__buf_2 fanout468 (.A(net104),
    .X(net468));
 sky130_fd_sc_hd__clkbuf_4 fanout469 (.A(net102),
    .X(net469));
 sky130_fd_sc_hd__clkbuf_4 fanout470 (.A(net101),
    .X(net470));
 sky130_fd_sc_hd__buf_4 fanout471 (.A(net100),
    .X(net471));
 sky130_fd_sc_hd__clkbuf_4 fanout472 (.A(net99),
    .X(net472));
 sky130_fd_sc_hd__clkbuf_4 fanout473 (.A(net98),
    .X(net473));
 sky130_fd_sc_hd__clkbuf_4 fanout474 (.A(net97),
    .X(net474));
 sky130_fd_sc_hd__clkbuf_4 fanout475 (.A(net96),
    .X(net475));
 sky130_fd_sc_hd__clkbuf_4 fanout476 (.A(net95),
    .X(net476));
 sky130_fd_sc_hd__clkbuf_2 input1 (.A(DO_SRAM0),
    .X(net1));
 sky130_fd_sc_hd__clkbuf_2 input2 (.A(DO_SRAM1),
    .X(net2));
 sky130_fd_sc_hd__clkbuf_2 input3 (.A(DO_SRAM10),
    .X(net3));
 sky130_fd_sc_hd__clkbuf_2 input4 (.A(DO_SRAM11),
    .X(net4));
 sky130_fd_sc_hd__dlymetal6s2s_1 input5 (.A(DO_SRAM12),
    .X(net5));
 sky130_fd_sc_hd__clkbuf_2 input6 (.A(DO_SRAM13),
    .X(net6));
 sky130_fd_sc_hd__clkbuf_2 input7 (.A(DO_SRAM14),
    .X(net7));
 sky130_fd_sc_hd__dlymetal6s2s_1 input8 (.A(DO_SRAM15),
    .X(net8));
 sky130_fd_sc_hd__buf_2 input9 (.A(DO_SRAM16),
    .X(net9));
 sky130_fd_sc_hd__clkbuf_4 input10 (.A(DO_SRAM17),
    .X(net10));
 sky130_fd_sc_hd__buf_2 input11 (.A(DO_SRAM18),
    .X(net11));
 sky130_fd_sc_hd__clkbuf_4 input12 (.A(DO_SRAM19),
    .X(net12));
 sky130_fd_sc_hd__clkbuf_2 input13 (.A(DO_SRAM2),
    .X(net13));
 sky130_fd_sc_hd__buf_2 input14 (.A(DO_SRAM20),
    .X(net14));
 sky130_fd_sc_hd__buf_2 input15 (.A(DO_SRAM21),
    .X(net15));
 sky130_fd_sc_hd__clkbuf_4 input16 (.A(DO_SRAM22),
    .X(net16));
 sky130_fd_sc_hd__buf_2 input17 (.A(DO_SRAM23),
    .X(net17));
 sky130_fd_sc_hd__buf_2 input18 (.A(DO_SRAM24),
    .X(net18));
 sky130_fd_sc_hd__clkbuf_2 input19 (.A(DO_SRAM25),
    .X(net19));
 sky130_fd_sc_hd__buf_2 input20 (.A(DO_SRAM26),
    .X(net20));
 sky130_fd_sc_hd__clkbuf_2 input21 (.A(DO_SRAM27),
    .X(net21));
 sky130_fd_sc_hd__buf_2 input22 (.A(DO_SRAM28),
    .X(net22));
 sky130_fd_sc_hd__buf_2 input23 (.A(DO_SRAM29),
    .X(net23));
 sky130_fd_sc_hd__buf_2 input24 (.A(DO_SRAM3),
    .X(net24));
 sky130_fd_sc_hd__buf_2 input25 (.A(DO_SRAM30),
    .X(net25));
 sky130_fd_sc_hd__clkbuf_2 input26 (.A(DO_SRAM31),
    .X(net26));
 sky130_fd_sc_hd__clkbuf_2 input27 (.A(DO_SRAM4),
    .X(net27));
 sky130_fd_sc_hd__clkbuf_2 input28 (.A(DO_SRAM5),
    .X(net28));
 sky130_fd_sc_hd__clkbuf_2 input29 (.A(DO_SRAM6),
    .X(net29));
 sky130_fd_sc_hd__clkbuf_2 input30 (.A(DO_SRAM7),
    .X(net30));
 sky130_fd_sc_hd__dlymetal6s2s_1 input31 (.A(DO_SRAM8),
    .X(net31));
 sky130_fd_sc_hd__clkbuf_2 input32 (.A(DO_SRAM9),
    .X(net32));
 sky130_fd_sc_hd__clkbuf_4 input33 (.A(Tile_X0Y0_E1END[0]),
    .X(net33));
 sky130_fd_sc_hd__buf_2 input34 (.A(Tile_X0Y0_E1END[1]),
    .X(net34));
 sky130_fd_sc_hd__buf_2 input35 (.A(Tile_X0Y0_E1END[2]),
    .X(net35));
 sky130_fd_sc_hd__clkbuf_4 input36 (.A(Tile_X0Y0_E1END[3]),
    .X(net36));
 sky130_fd_sc_hd__clkbuf_2 input37 (.A(Tile_X0Y0_E2END[0]),
    .X(net37));
 sky130_fd_sc_hd__dlymetal6s2s_1 input38 (.A(Tile_X0Y0_E2END[1]),
    .X(net38));
 sky130_fd_sc_hd__dlymetal6s2s_1 input39 (.A(Tile_X0Y0_E2END[2]),
    .X(net39));
 sky130_fd_sc_hd__dlymetal6s2s_1 input40 (.A(Tile_X0Y0_E2END[3]),
    .X(net40));
 sky130_fd_sc_hd__clkbuf_2 input41 (.A(Tile_X0Y0_E2END[4]),
    .X(net41));
 sky130_fd_sc_hd__buf_1 input42 (.A(Tile_X0Y0_E2END[5]),
    .X(net42));
 sky130_fd_sc_hd__buf_1 input43 (.A(Tile_X0Y0_E2END[6]),
    .X(net43));
 sky130_fd_sc_hd__clkbuf_2 input44 (.A(Tile_X0Y0_E2END[7]),
    .X(net44));
 sky130_fd_sc_hd__clkbuf_2 input45 (.A(Tile_X0Y0_E2MID[0]),
    .X(net45));
 sky130_fd_sc_hd__dlymetal6s2s_1 input46 (.A(Tile_X0Y0_E2MID[1]),
    .X(net46));
 sky130_fd_sc_hd__buf_1 input47 (.A(Tile_X0Y0_E2MID[2]),
    .X(net47));
 sky130_fd_sc_hd__dlymetal6s2s_1 input48 (.A(Tile_X0Y0_E2MID[3]),
    .X(net48));
 sky130_fd_sc_hd__clkbuf_2 input49 (.A(Tile_X0Y0_E2MID[4]),
    .X(net49));
 sky130_fd_sc_hd__buf_1 input50 (.A(Tile_X0Y0_E2MID[5]),
    .X(net50));
 sky130_fd_sc_hd__buf_1 input51 (.A(Tile_X0Y0_E2MID[6]),
    .X(net51));
 sky130_fd_sc_hd__clkbuf_2 input52 (.A(Tile_X0Y0_E2MID[7]),
    .X(net52));
 sky130_fd_sc_hd__buf_2 input53 (.A(Tile_X0Y0_E6END[0]),
    .X(net53));
 sky130_fd_sc_hd__clkbuf_2 input54 (.A(Tile_X0Y0_E6END[10]),
    .X(net54));
 sky130_fd_sc_hd__clkbuf_2 input55 (.A(Tile_X0Y0_E6END[11]),
    .X(net55));
 sky130_fd_sc_hd__clkbuf_2 input56 (.A(Tile_X0Y0_E6END[1]),
    .X(net56));
 sky130_fd_sc_hd__clkbuf_2 input57 (.A(Tile_X0Y0_E6END[2]),
    .X(net57));
 sky130_fd_sc_hd__clkbuf_2 input58 (.A(Tile_X0Y0_E6END[3]),
    .X(net58));
 sky130_fd_sc_hd__buf_2 input59 (.A(Tile_X0Y0_E6END[4]),
    .X(net59));
 sky130_fd_sc_hd__clkbuf_2 input60 (.A(Tile_X0Y0_E6END[5]),
    .X(net60));
 sky130_fd_sc_hd__clkbuf_2 input61 (.A(Tile_X0Y0_E6END[6]),
    .X(net61));
 sky130_fd_sc_hd__buf_2 input62 (.A(Tile_X0Y0_E6END[7]),
    .X(net62));
 sky130_fd_sc_hd__buf_2 input63 (.A(Tile_X0Y0_E6END[8]),
    .X(net63));
 sky130_fd_sc_hd__dlymetal6s2s_1 input64 (.A(Tile_X0Y0_E6END[9]),
    .X(net64));
 sky130_fd_sc_hd__buf_2 input65 (.A(Tile_X0Y0_EE4END[0]),
    .X(net65));
 sky130_fd_sc_hd__buf_1 input66 (.A(Tile_X0Y0_EE4END[10]),
    .X(net66));
 sky130_fd_sc_hd__clkbuf_2 input67 (.A(Tile_X0Y0_EE4END[11]),
    .X(net67));
 sky130_fd_sc_hd__buf_2 input68 (.A(Tile_X0Y0_EE4END[12]),
    .X(net68));
 sky130_fd_sc_hd__buf_1 input69 (.A(Tile_X0Y0_EE4END[13]),
    .X(net69));
 sky130_fd_sc_hd__dlymetal6s2s_1 input70 (.A(Tile_X0Y0_EE4END[14]),
    .X(net70));
 sky130_fd_sc_hd__clkbuf_2 input71 (.A(Tile_X0Y0_EE4END[15]),
    .X(net71));
 sky130_fd_sc_hd__buf_1 input72 (.A(Tile_X0Y0_EE4END[1]),
    .X(net72));
 sky130_fd_sc_hd__buf_1 input73 (.A(Tile_X0Y0_EE4END[2]),
    .X(net73));
 sky130_fd_sc_hd__clkbuf_2 input74 (.A(Tile_X0Y0_EE4END[3]),
    .X(net74));
 sky130_fd_sc_hd__clkbuf_2 input75 (.A(Tile_X0Y0_EE4END[4]),
    .X(net75));
 sky130_fd_sc_hd__buf_1 input76 (.A(Tile_X0Y0_EE4END[5]),
    .X(net76));
 sky130_fd_sc_hd__dlymetal6s2s_1 input77 (.A(Tile_X0Y0_EE4END[6]),
    .X(net77));
 sky130_fd_sc_hd__clkbuf_2 input78 (.A(Tile_X0Y0_EE4END[7]),
    .X(net78));
 sky130_fd_sc_hd__clkbuf_2 input79 (.A(Tile_X0Y0_EE4END[8]),
    .X(net79));
 sky130_fd_sc_hd__buf_1 input80 (.A(Tile_X0Y0_EE4END[9]),
    .X(net80));
 sky130_fd_sc_hd__clkbuf_4 input81 (.A(Tile_X0Y0_FrameData[0]),
    .X(net81));
 sky130_fd_sc_hd__clkbuf_4 input82 (.A(Tile_X0Y0_FrameData[10]),
    .X(net82));
 sky130_fd_sc_hd__clkbuf_4 input83 (.A(Tile_X0Y0_FrameData[11]),
    .X(net83));
 sky130_fd_sc_hd__buf_4 input84 (.A(Tile_X0Y0_FrameData[12]),
    .X(net84));
 sky130_fd_sc_hd__buf_4 input85 (.A(Tile_X0Y0_FrameData[13]),
    .X(net85));
 sky130_fd_sc_hd__buf_4 input86 (.A(Tile_X0Y0_FrameData[14]),
    .X(net86));
 sky130_fd_sc_hd__buf_4 input87 (.A(Tile_X0Y0_FrameData[15]),
    .X(net87));
 sky130_fd_sc_hd__buf_4 input88 (.A(Tile_X0Y0_FrameData[16]),
    .X(net88));
 sky130_fd_sc_hd__buf_4 input89 (.A(Tile_X0Y0_FrameData[17]),
    .X(net89));
 sky130_fd_sc_hd__clkbuf_4 input90 (.A(Tile_X0Y0_FrameData[18]),
    .X(net90));
 sky130_fd_sc_hd__clkbuf_4 input91 (.A(Tile_X0Y0_FrameData[19]),
    .X(net91));
 sky130_fd_sc_hd__clkbuf_4 input92 (.A(Tile_X0Y0_FrameData[1]),
    .X(net92));
 sky130_fd_sc_hd__buf_4 input93 (.A(Tile_X0Y0_FrameData[20]),
    .X(net93));
 sky130_fd_sc_hd__buf_4 input94 (.A(Tile_X0Y0_FrameData[21]),
    .X(net94));
 sky130_fd_sc_hd__buf_1 input95 (.A(Tile_X0Y0_FrameData[22]),
    .X(net95));
 sky130_fd_sc_hd__dlymetal6s2s_1 input96 (.A(Tile_X0Y0_FrameData[23]),
    .X(net96));
 sky130_fd_sc_hd__clkbuf_2 input97 (.A(Tile_X0Y0_FrameData[24]),
    .X(net97));
 sky130_fd_sc_hd__clkbuf_2 input98 (.A(Tile_X0Y0_FrameData[25]),
    .X(net98));
 sky130_fd_sc_hd__clkbuf_2 input99 (.A(Tile_X0Y0_FrameData[26]),
    .X(net99));
 sky130_fd_sc_hd__clkbuf_2 input100 (.A(Tile_X0Y0_FrameData[27]),
    .X(net100));
 sky130_fd_sc_hd__clkbuf_2 input101 (.A(Tile_X0Y0_FrameData[28]),
    .X(net101));
 sky130_fd_sc_hd__clkbuf_2 input102 (.A(Tile_X0Y0_FrameData[29]),
    .X(net102));
 sky130_fd_sc_hd__clkbuf_4 input103 (.A(Tile_X0Y0_FrameData[2]),
    .X(net103));
 sky130_fd_sc_hd__clkbuf_2 input104 (.A(Tile_X0Y0_FrameData[30]),
    .X(net104));
 sky130_fd_sc_hd__clkbuf_2 input105 (.A(Tile_X0Y0_FrameData[31]),
    .X(net105));
 sky130_fd_sc_hd__clkbuf_4 input106 (.A(Tile_X0Y0_FrameData[3]),
    .X(net106));
 sky130_fd_sc_hd__clkbuf_4 input107 (.A(Tile_X0Y0_FrameData[4]),
    .X(net107));
 sky130_fd_sc_hd__clkbuf_4 input108 (.A(Tile_X0Y0_FrameData[5]),
    .X(net108));
 sky130_fd_sc_hd__clkbuf_4 input109 (.A(Tile_X0Y0_FrameData[6]),
    .X(net109));
 sky130_fd_sc_hd__clkbuf_4 input110 (.A(Tile_X0Y0_FrameData[7]),
    .X(net110));
 sky130_fd_sc_hd__buf_4 input111 (.A(Tile_X0Y0_FrameData[8]),
    .X(net111));
 sky130_fd_sc_hd__buf_4 input112 (.A(Tile_X0Y0_FrameData[9]),
    .X(net112));
 sky130_fd_sc_hd__buf_2 input113 (.A(Tile_X0Y0_S1END[0]),
    .X(net113));
 sky130_fd_sc_hd__buf_2 input114 (.A(Tile_X0Y0_S1END[1]),
    .X(net114));
 sky130_fd_sc_hd__clkbuf_2 input115 (.A(Tile_X0Y0_S1END[2]),
    .X(net115));
 sky130_fd_sc_hd__clkbuf_2 input116 (.A(Tile_X0Y0_S1END[3]),
    .X(net116));
 sky130_fd_sc_hd__clkbuf_2 input117 (.A(Tile_X0Y0_S2END[0]),
    .X(net117));
 sky130_fd_sc_hd__clkbuf_2 input118 (.A(Tile_X0Y0_S2END[1]),
    .X(net118));
 sky130_fd_sc_hd__clkbuf_2 input119 (.A(Tile_X0Y0_S2END[2]),
    .X(net119));
 sky130_fd_sc_hd__clkbuf_2 input120 (.A(Tile_X0Y0_S2END[3]),
    .X(net120));
 sky130_fd_sc_hd__dlymetal6s2s_1 input121 (.A(Tile_X0Y0_S2END[4]),
    .X(net121));
 sky130_fd_sc_hd__clkbuf_2 input122 (.A(Tile_X0Y0_S2END[5]),
    .X(net122));
 sky130_fd_sc_hd__clkbuf_2 input123 (.A(Tile_X0Y0_S2END[6]),
    .X(net123));
 sky130_fd_sc_hd__clkbuf_2 input124 (.A(Tile_X0Y0_S2END[7]),
    .X(net124));
 sky130_fd_sc_hd__clkbuf_2 input125 (.A(Tile_X0Y0_S2MID[0]),
    .X(net125));
 sky130_fd_sc_hd__clkbuf_2 input126 (.A(Tile_X0Y0_S2MID[1]),
    .X(net126));
 sky130_fd_sc_hd__buf_2 input127 (.A(Tile_X0Y0_S2MID[2]),
    .X(net127));
 sky130_fd_sc_hd__buf_2 input128 (.A(Tile_X0Y0_S2MID[3]),
    .X(net128));
 sky130_fd_sc_hd__clkbuf_2 input129 (.A(Tile_X0Y0_S2MID[4]),
    .X(net129));
 sky130_fd_sc_hd__clkbuf_2 input130 (.A(Tile_X0Y0_S2MID[5]),
    .X(net130));
 sky130_fd_sc_hd__clkbuf_2 input131 (.A(Tile_X0Y0_S2MID[6]),
    .X(net131));
 sky130_fd_sc_hd__clkbuf_2 input132 (.A(Tile_X0Y0_S2MID[7]),
    .X(net132));
 sky130_fd_sc_hd__clkbuf_2 input133 (.A(Tile_X0Y0_S4END[0]),
    .X(net133));
 sky130_fd_sc_hd__buf_2 input134 (.A(Tile_X0Y0_S4END[1]),
    .X(net134));
 sky130_fd_sc_hd__clkbuf_2 input135 (.A(Tile_X0Y0_S4END[2]),
    .X(net135));
 sky130_fd_sc_hd__clkbuf_2 input136 (.A(Tile_X0Y0_S4END[3]),
    .X(net136));
 sky130_fd_sc_hd__clkbuf_4 input137 (.A(Tile_X0Y0_S4END[4]),
    .X(net137));
 sky130_fd_sc_hd__clkbuf_4 input138 (.A(Tile_X0Y0_S4END[5]),
    .X(net138));
 sky130_fd_sc_hd__clkbuf_4 input139 (.A(Tile_X0Y0_S4END[6]),
    .X(net139));
 sky130_fd_sc_hd__clkbuf_4 input140 (.A(Tile_X0Y0_S4END[7]),
    .X(net140));
 sky130_fd_sc_hd__buf_2 input141 (.A(Tile_X0Y1_E1END[0]),
    .X(net141));
 sky130_fd_sc_hd__buf_2 input142 (.A(Tile_X0Y1_E1END[1]),
    .X(net142));
 sky130_fd_sc_hd__clkbuf_2 input143 (.A(Tile_X0Y1_E1END[2]),
    .X(net143));
 sky130_fd_sc_hd__buf_2 input144 (.A(Tile_X0Y1_E1END[3]),
    .X(net144));
 sky130_fd_sc_hd__dlymetal6s2s_1 input145 (.A(Tile_X0Y1_E2END[0]),
    .X(net145));
 sky130_fd_sc_hd__clkbuf_2 input146 (.A(Tile_X0Y1_E2END[1]),
    .X(net146));
 sky130_fd_sc_hd__clkbuf_2 input147 (.A(Tile_X0Y1_E2END[2]),
    .X(net147));
 sky130_fd_sc_hd__clkbuf_2 input148 (.A(Tile_X0Y1_E2END[3]),
    .X(net148));
 sky130_fd_sc_hd__buf_2 input149 (.A(Tile_X0Y1_E2END[4]),
    .X(net149));
 sky130_fd_sc_hd__clkbuf_2 input150 (.A(Tile_X0Y1_E2END[5]),
    .X(net150));
 sky130_fd_sc_hd__buf_1 input151 (.A(Tile_X0Y1_E2END[6]),
    .X(net151));
 sky130_fd_sc_hd__clkbuf_2 input152 (.A(Tile_X0Y1_E2END[7]),
    .X(net152));
 sky130_fd_sc_hd__clkbuf_2 input153 (.A(Tile_X0Y1_E2MID[0]),
    .X(net153));
 sky130_fd_sc_hd__clkbuf_2 input154 (.A(Tile_X0Y1_E2MID[1]),
    .X(net154));
 sky130_fd_sc_hd__dlymetal6s2s_1 input155 (.A(Tile_X0Y1_E2MID[2]),
    .X(net155));
 sky130_fd_sc_hd__clkbuf_2 input156 (.A(Tile_X0Y1_E2MID[3]),
    .X(net156));
 sky130_fd_sc_hd__clkbuf_2 input157 (.A(Tile_X0Y1_E2MID[4]),
    .X(net157));
 sky130_fd_sc_hd__dlymetal6s2s_1 input158 (.A(Tile_X0Y1_E2MID[5]),
    .X(net158));
 sky130_fd_sc_hd__clkbuf_2 input159 (.A(Tile_X0Y1_E2MID[6]),
    .X(net159));
 sky130_fd_sc_hd__clkbuf_2 input160 (.A(Tile_X0Y1_E2MID[7]),
    .X(net160));
 sky130_fd_sc_hd__clkbuf_2 input161 (.A(Tile_X0Y1_E6END[0]),
    .X(net161));
 sky130_fd_sc_hd__clkbuf_2 input162 (.A(Tile_X0Y1_E6END[10]),
    .X(net162));
 sky130_fd_sc_hd__clkbuf_2 input163 (.A(Tile_X0Y1_E6END[11]),
    .X(net163));
 sky130_fd_sc_hd__buf_1 input164 (.A(Tile_X0Y1_E6END[1]),
    .X(net164));
 sky130_fd_sc_hd__buf_1 input165 (.A(Tile_X0Y1_E6END[2]),
    .X(net165));
 sky130_fd_sc_hd__clkbuf_2 input166 (.A(Tile_X0Y1_E6END[3]),
    .X(net166));
 sky130_fd_sc_hd__clkbuf_2 input167 (.A(Tile_X0Y1_E6END[4]),
    .X(net167));
 sky130_fd_sc_hd__clkbuf_2 input168 (.A(Tile_X0Y1_E6END[5]),
    .X(net168));
 sky130_fd_sc_hd__clkbuf_2 input169 (.A(Tile_X0Y1_E6END[6]),
    .X(net169));
 sky130_fd_sc_hd__buf_2 input170 (.A(Tile_X0Y1_E6END[7]),
    .X(net170));
 sky130_fd_sc_hd__clkbuf_2 input171 (.A(Tile_X0Y1_E6END[8]),
    .X(net171));
 sky130_fd_sc_hd__dlymetal6s2s_1 input172 (.A(Tile_X0Y1_E6END[9]),
    .X(net172));
 sky130_fd_sc_hd__clkbuf_2 input173 (.A(Tile_X0Y1_EE4END[0]),
    .X(net173));
 sky130_fd_sc_hd__buf_1 input174 (.A(Tile_X0Y1_EE4END[10]),
    .X(net174));
 sky130_fd_sc_hd__dlymetal6s2s_1 input175 (.A(Tile_X0Y1_EE4END[11]),
    .X(net175));
 sky130_fd_sc_hd__clkbuf_2 input176 (.A(Tile_X0Y1_EE4END[12]),
    .X(net176));
 sky130_fd_sc_hd__dlymetal6s2s_1 input177 (.A(Tile_X0Y1_EE4END[13]),
    .X(net177));
 sky130_fd_sc_hd__dlymetal6s2s_1 input178 (.A(Tile_X0Y1_EE4END[14]),
    .X(net178));
 sky130_fd_sc_hd__clkbuf_2 input179 (.A(Tile_X0Y1_EE4END[15]),
    .X(net179));
 sky130_fd_sc_hd__dlymetal6s2s_1 input180 (.A(Tile_X0Y1_EE4END[1]),
    .X(net180));
 sky130_fd_sc_hd__dlymetal6s2s_1 input181 (.A(Tile_X0Y1_EE4END[2]),
    .X(net181));
 sky130_fd_sc_hd__clkbuf_2 input182 (.A(Tile_X0Y1_EE4END[3]),
    .X(net182));
 sky130_fd_sc_hd__clkbuf_2 input183 (.A(Tile_X0Y1_EE4END[4]),
    .X(net183));
 sky130_fd_sc_hd__buf_1 input184 (.A(Tile_X0Y1_EE4END[5]),
    .X(net184));
 sky130_fd_sc_hd__buf_1 input185 (.A(Tile_X0Y1_EE4END[6]),
    .X(net185));
 sky130_fd_sc_hd__clkbuf_2 input186 (.A(Tile_X0Y1_EE4END[7]),
    .X(net186));
 sky130_fd_sc_hd__clkbuf_2 input187 (.A(Tile_X0Y1_EE4END[8]),
    .X(net187));
 sky130_fd_sc_hd__buf_1 input188 (.A(Tile_X0Y1_EE4END[9]),
    .X(net188));
 sky130_fd_sc_hd__buf_4 input189 (.A(Tile_X0Y1_FrameData[0]),
    .X(net189));
 sky130_fd_sc_hd__clkbuf_4 input190 (.A(Tile_X0Y1_FrameData[10]),
    .X(net190));
 sky130_fd_sc_hd__clkbuf_4 input191 (.A(Tile_X0Y1_FrameData[11]),
    .X(net191));
 sky130_fd_sc_hd__clkbuf_4 input192 (.A(Tile_X0Y1_FrameData[12]),
    .X(net192));
 sky130_fd_sc_hd__clkbuf_4 input193 (.A(Tile_X0Y1_FrameData[13]),
    .X(net193));
 sky130_fd_sc_hd__buf_1 input194 (.A(Tile_X0Y1_FrameData[14]),
    .X(net194));
 sky130_fd_sc_hd__buf_1 input195 (.A(Tile_X0Y1_FrameData[15]),
    .X(net195));
 sky130_fd_sc_hd__clkbuf_1 input196 (.A(Tile_X0Y1_FrameData[18]),
    .X(net196));
 sky130_fd_sc_hd__clkbuf_1 input197 (.A(Tile_X0Y1_FrameData[19]),
    .X(net197));
 sky130_fd_sc_hd__buf_4 input198 (.A(Tile_X0Y1_FrameData[1]),
    .X(net198));
 sky130_fd_sc_hd__buf_1 input199 (.A(Tile_X0Y1_FrameData[20]),
    .X(net199));
 sky130_fd_sc_hd__buf_1 input200 (.A(Tile_X0Y1_FrameData[21]),
    .X(net200));
 sky130_fd_sc_hd__dlymetal6s2s_1 input201 (.A(Tile_X0Y1_FrameData[22]),
    .X(net201));
 sky130_fd_sc_hd__dlymetal6s2s_1 input202 (.A(Tile_X0Y1_FrameData[23]),
    .X(net202));
 sky130_fd_sc_hd__clkbuf_2 input203 (.A(Tile_X0Y1_FrameData[24]),
    .X(net203));
 sky130_fd_sc_hd__clkbuf_2 input204 (.A(Tile_X0Y1_FrameData[25]),
    .X(net204));
 sky130_fd_sc_hd__buf_1 input205 (.A(Tile_X0Y1_FrameData[26]),
    .X(net205));
 sky130_fd_sc_hd__buf_1 input206 (.A(Tile_X0Y1_FrameData[27]),
    .X(net206));
 sky130_fd_sc_hd__buf_1 input207 (.A(Tile_X0Y1_FrameData[28]),
    .X(net207));
 sky130_fd_sc_hd__buf_1 input208 (.A(Tile_X0Y1_FrameData[29]),
    .X(net208));
 sky130_fd_sc_hd__buf_2 input209 (.A(Tile_X0Y1_FrameData[2]),
    .X(net209));
 sky130_fd_sc_hd__buf_1 input210 (.A(Tile_X0Y1_FrameData[30]),
    .X(net210));
 sky130_fd_sc_hd__buf_1 input211 (.A(Tile_X0Y1_FrameData[31]),
    .X(net211));
 sky130_fd_sc_hd__clkbuf_4 input212 (.A(Tile_X0Y1_FrameData[3]),
    .X(net212));
 sky130_fd_sc_hd__clkbuf_4 input213 (.A(Tile_X0Y1_FrameData[4]),
    .X(net213));
 sky130_fd_sc_hd__clkbuf_4 input214 (.A(Tile_X0Y1_FrameData[5]),
    .X(net214));
 sky130_fd_sc_hd__clkbuf_4 input215 (.A(Tile_X0Y1_FrameData[6]),
    .X(net215));
 sky130_fd_sc_hd__clkbuf_4 input216 (.A(Tile_X0Y1_FrameData[7]),
    .X(net216));
 sky130_fd_sc_hd__buf_4 input217 (.A(Tile_X0Y1_FrameData[8]),
    .X(net217));
 sky130_fd_sc_hd__buf_4 input218 (.A(Tile_X0Y1_FrameData[9]),
    .X(net218));
 sky130_fd_sc_hd__clkbuf_4 input219 (.A(Tile_X0Y1_FrameStrobe[9]),
    .X(net219));
 sky130_fd_sc_hd__buf_2 input220 (.A(Tile_X0Y1_N1END[0]),
    .X(net220));
 sky130_fd_sc_hd__clkbuf_2 input221 (.A(Tile_X0Y1_N1END[1]),
    .X(net221));
 sky130_fd_sc_hd__buf_2 input222 (.A(Tile_X0Y1_N1END[2]),
    .X(net222));
 sky130_fd_sc_hd__buf_2 input223 (.A(Tile_X0Y1_N1END[3]),
    .X(net223));
 sky130_fd_sc_hd__clkbuf_2 input224 (.A(Tile_X0Y1_N2END[0]),
    .X(net224));
 sky130_fd_sc_hd__clkbuf_2 input225 (.A(Tile_X0Y1_N2END[1]),
    .X(net225));
 sky130_fd_sc_hd__clkbuf_2 input226 (.A(Tile_X0Y1_N2END[2]),
    .X(net226));
 sky130_fd_sc_hd__clkbuf_2 input227 (.A(Tile_X0Y1_N2END[3]),
    .X(net227));
 sky130_fd_sc_hd__clkbuf_2 input228 (.A(Tile_X0Y1_N2END[4]),
    .X(net228));
 sky130_fd_sc_hd__clkbuf_2 input229 (.A(Tile_X0Y1_N2END[5]),
    .X(net229));
 sky130_fd_sc_hd__clkbuf_2 input230 (.A(Tile_X0Y1_N2END[6]),
    .X(net230));
 sky130_fd_sc_hd__clkbuf_2 input231 (.A(Tile_X0Y1_N2END[7]),
    .X(net231));
 sky130_fd_sc_hd__buf_2 input232 (.A(Tile_X0Y1_N2MID[0]),
    .X(net232));
 sky130_fd_sc_hd__clkbuf_2 input233 (.A(Tile_X0Y1_N2MID[1]),
    .X(net233));
 sky130_fd_sc_hd__clkbuf_2 input234 (.A(Tile_X0Y1_N2MID[2]),
    .X(net234));
 sky130_fd_sc_hd__clkbuf_2 input235 (.A(Tile_X0Y1_N2MID[3]),
    .X(net235));
 sky130_fd_sc_hd__clkbuf_2 input236 (.A(Tile_X0Y1_N2MID[4]),
    .X(net236));
 sky130_fd_sc_hd__clkbuf_2 input237 (.A(Tile_X0Y1_N2MID[5]),
    .X(net237));
 sky130_fd_sc_hd__buf_2 input238 (.A(Tile_X0Y1_N2MID[6]),
    .X(net238));
 sky130_fd_sc_hd__buf_2 input239 (.A(Tile_X0Y1_N2MID[7]),
    .X(net239));
 sky130_fd_sc_hd__clkbuf_2 input240 (.A(Tile_X0Y1_N4END[0]),
    .X(net240));
 sky130_fd_sc_hd__clkbuf_2 input241 (.A(Tile_X0Y1_N4END[1]),
    .X(net241));
 sky130_fd_sc_hd__clkbuf_2 input242 (.A(Tile_X0Y1_N4END[2]),
    .X(net242));
 sky130_fd_sc_hd__clkbuf_2 input243 (.A(Tile_X0Y1_N4END[3]),
    .X(net243));
 sky130_fd_sc_hd__clkbuf_4 input244 (.A(Tile_X0Y1_N4END[4]),
    .X(net244));
 sky130_fd_sc_hd__buf_2 input245 (.A(Tile_X0Y1_N4END[5]),
    .X(net245));
 sky130_fd_sc_hd__buf_2 input246 (.A(Tile_X0Y1_N4END[6]),
    .X(net246));
 sky130_fd_sc_hd__clkbuf_4 input247 (.A(Tile_X0Y1_N4END[7]),
    .X(net247));
 sky130_fd_sc_hd__buf_2 output248 (.A(net248),
    .X(AD_SRAM0));
 sky130_fd_sc_hd__buf_2 output249 (.A(net249),
    .X(AD_SRAM1));
 sky130_fd_sc_hd__buf_2 output250 (.A(net250),
    .X(AD_SRAM2));
 sky130_fd_sc_hd__buf_2 output251 (.A(net251),
    .X(AD_SRAM3));
 sky130_fd_sc_hd__buf_2 output252 (.A(net252),
    .X(AD_SRAM4));
 sky130_fd_sc_hd__buf_2 output253 (.A(net253),
    .X(AD_SRAM5));
 sky130_fd_sc_hd__buf_2 output254 (.A(net254),
    .X(AD_SRAM6));
 sky130_fd_sc_hd__buf_2 output255 (.A(net255),
    .X(AD_SRAM7));
 sky130_fd_sc_hd__buf_2 output256 (.A(net256),
    .X(AD_SRAM8));
 sky130_fd_sc_hd__buf_2 output257 (.A(net257),
    .X(AD_SRAM9));
 sky130_fd_sc_hd__buf_2 output258 (.A(net258),
    .X(BEN_SRAM0));
 sky130_fd_sc_hd__buf_2 output259 (.A(net259),
    .X(BEN_SRAM1));
 sky130_fd_sc_hd__buf_2 output260 (.A(net260),
    .X(BEN_SRAM10));
 sky130_fd_sc_hd__buf_2 output261 (.A(net261),
    .X(BEN_SRAM11));
 sky130_fd_sc_hd__buf_2 output262 (.A(net262),
    .X(BEN_SRAM12));
 sky130_fd_sc_hd__buf_2 output263 (.A(net263),
    .X(BEN_SRAM13));
 sky130_fd_sc_hd__buf_2 output264 (.A(net264),
    .X(BEN_SRAM14));
 sky130_fd_sc_hd__buf_2 output265 (.A(net265),
    .X(BEN_SRAM15));
 sky130_fd_sc_hd__buf_2 output266 (.A(net266),
    .X(BEN_SRAM16));
 sky130_fd_sc_hd__buf_2 output267 (.A(net267),
    .X(BEN_SRAM17));
 sky130_fd_sc_hd__buf_2 output268 (.A(net268),
    .X(BEN_SRAM18));
 sky130_fd_sc_hd__buf_2 output269 (.A(net269),
    .X(BEN_SRAM19));
 sky130_fd_sc_hd__buf_2 output270 (.A(net270),
    .X(BEN_SRAM2));
 sky130_fd_sc_hd__buf_2 output271 (.A(net271),
    .X(BEN_SRAM20));
 sky130_fd_sc_hd__buf_2 output272 (.A(net272),
    .X(BEN_SRAM21));
 sky130_fd_sc_hd__buf_2 output273 (.A(net273),
    .X(BEN_SRAM22));
 sky130_fd_sc_hd__buf_2 output274 (.A(net274),
    .X(BEN_SRAM23));
 sky130_fd_sc_hd__buf_2 output275 (.A(net275),
    .X(BEN_SRAM24));
 sky130_fd_sc_hd__buf_2 output276 (.A(net276),
    .X(BEN_SRAM25));
 sky130_fd_sc_hd__buf_2 output277 (.A(net277),
    .X(BEN_SRAM26));
 sky130_fd_sc_hd__buf_2 output278 (.A(net278),
    .X(BEN_SRAM27));
 sky130_fd_sc_hd__buf_2 output279 (.A(net279),
    .X(BEN_SRAM28));
 sky130_fd_sc_hd__buf_2 output280 (.A(net280),
    .X(BEN_SRAM29));
 sky130_fd_sc_hd__buf_2 output281 (.A(net281),
    .X(BEN_SRAM3));
 sky130_fd_sc_hd__buf_2 output282 (.A(net282),
    .X(BEN_SRAM30));
 sky130_fd_sc_hd__buf_2 output283 (.A(net283),
    .X(BEN_SRAM31));
 sky130_fd_sc_hd__buf_2 output284 (.A(net284),
    .X(BEN_SRAM4));
 sky130_fd_sc_hd__buf_2 output285 (.A(net285),
    .X(BEN_SRAM5));
 sky130_fd_sc_hd__buf_2 output286 (.A(net286),
    .X(BEN_SRAM6));
 sky130_fd_sc_hd__buf_2 output287 (.A(net287),
    .X(BEN_SRAM7));
 sky130_fd_sc_hd__buf_2 output288 (.A(net288),
    .X(BEN_SRAM8));
 sky130_fd_sc_hd__buf_2 output289 (.A(net289),
    .X(BEN_SRAM9));
 sky130_fd_sc_hd__buf_1 output290 (.A(net290),
    .X(CLOCK_SRAM));
 sky130_fd_sc_hd__buf_2 output291 (.A(net291),
    .X(DI_SRAM0));
 sky130_fd_sc_hd__buf_2 output292 (.A(net292),
    .X(DI_SRAM1));
 sky130_fd_sc_hd__buf_2 output293 (.A(net293),
    .X(DI_SRAM10));
 sky130_fd_sc_hd__buf_2 output294 (.A(net294),
    .X(DI_SRAM11));
 sky130_fd_sc_hd__buf_2 output295 (.A(net295),
    .X(DI_SRAM12));
 sky130_fd_sc_hd__buf_2 output296 (.A(net296),
    .X(DI_SRAM13));
 sky130_fd_sc_hd__buf_2 output297 (.A(net297),
    .X(DI_SRAM14));
 sky130_fd_sc_hd__buf_2 output298 (.A(net298),
    .X(DI_SRAM15));
 sky130_fd_sc_hd__buf_2 output299 (.A(net299),
    .X(DI_SRAM16));
 sky130_fd_sc_hd__buf_2 output300 (.A(net300),
    .X(DI_SRAM17));
 sky130_fd_sc_hd__buf_2 output301 (.A(net301),
    .X(DI_SRAM18));
 sky130_fd_sc_hd__buf_2 output302 (.A(net302),
    .X(DI_SRAM19));
 sky130_fd_sc_hd__buf_2 output303 (.A(net303),
    .X(DI_SRAM2));
 sky130_fd_sc_hd__buf_2 output304 (.A(net304),
    .X(DI_SRAM20));
 sky130_fd_sc_hd__buf_2 output305 (.A(net305),
    .X(DI_SRAM21));
 sky130_fd_sc_hd__buf_2 output306 (.A(net306),
    .X(DI_SRAM22));
 sky130_fd_sc_hd__buf_2 output307 (.A(net307),
    .X(DI_SRAM23));
 sky130_fd_sc_hd__buf_2 output308 (.A(net308),
    .X(DI_SRAM24));
 sky130_fd_sc_hd__buf_2 output309 (.A(net309),
    .X(DI_SRAM25));
 sky130_fd_sc_hd__buf_2 output310 (.A(net310),
    .X(DI_SRAM26));
 sky130_fd_sc_hd__buf_2 output311 (.A(net311),
    .X(DI_SRAM27));
 sky130_fd_sc_hd__buf_2 output312 (.A(net312),
    .X(DI_SRAM28));
 sky130_fd_sc_hd__buf_2 output313 (.A(net313),
    .X(DI_SRAM29));
 sky130_fd_sc_hd__buf_2 output314 (.A(net314),
    .X(DI_SRAM3));
 sky130_fd_sc_hd__buf_2 output315 (.A(net315),
    .X(DI_SRAM30));
 sky130_fd_sc_hd__buf_2 output316 (.A(net316),
    .X(DI_SRAM31));
 sky130_fd_sc_hd__buf_2 output317 (.A(net317),
    .X(DI_SRAM4));
 sky130_fd_sc_hd__buf_2 output318 (.A(net318),
    .X(DI_SRAM5));
 sky130_fd_sc_hd__buf_2 output319 (.A(net319),
    .X(DI_SRAM6));
 sky130_fd_sc_hd__buf_2 output320 (.A(net320),
    .X(DI_SRAM7));
 sky130_fd_sc_hd__buf_2 output321 (.A(net321),
    .X(DI_SRAM8));
 sky130_fd_sc_hd__buf_2 output322 (.A(net322),
    .X(DI_SRAM9));
 sky130_fd_sc_hd__buf_2 output323 (.A(net323),
    .X(EN_SRAM));
 sky130_fd_sc_hd__buf_2 output324 (.A(net324),
    .X(R_WB_SRAM));
 sky130_fd_sc_hd__buf_2 output325 (.A(net325),
    .X(Tile_X0Y0_FrameData_O[0]));
 sky130_fd_sc_hd__buf_2 output326 (.A(net326),
    .X(Tile_X0Y0_FrameData_O[10]));
 sky130_fd_sc_hd__buf_2 output327 (.A(net327),
    .X(Tile_X0Y0_FrameData_O[11]));
 sky130_fd_sc_hd__buf_2 output328 (.A(net328),
    .X(Tile_X0Y0_FrameData_O[12]));
 sky130_fd_sc_hd__buf_2 output329 (.A(net329),
    .X(Tile_X0Y0_FrameData_O[13]));
 sky130_fd_sc_hd__buf_2 output330 (.A(net330),
    .X(Tile_X0Y0_FrameData_O[14]));
 sky130_fd_sc_hd__buf_2 output331 (.A(net331),
    .X(Tile_X0Y0_FrameData_O[15]));
 sky130_fd_sc_hd__buf_2 output332 (.A(net332),
    .X(Tile_X0Y0_FrameData_O[16]));
 sky130_fd_sc_hd__buf_2 output333 (.A(net333),
    .X(Tile_X0Y0_FrameData_O[17]));
 sky130_fd_sc_hd__buf_2 output334 (.A(net334),
    .X(Tile_X0Y0_FrameData_O[18]));
 sky130_fd_sc_hd__buf_2 output335 (.A(net335),
    .X(Tile_X0Y0_FrameData_O[19]));
 sky130_fd_sc_hd__buf_2 output336 (.A(net336),
    .X(Tile_X0Y0_FrameData_O[1]));
 sky130_fd_sc_hd__buf_2 output337 (.A(net337),
    .X(Tile_X0Y0_FrameData_O[20]));
 sky130_fd_sc_hd__buf_2 output338 (.A(net338),
    .X(Tile_X0Y0_FrameData_O[21]));
 sky130_fd_sc_hd__buf_2 output339 (.A(net339),
    .X(Tile_X0Y0_FrameData_O[22]));
 sky130_fd_sc_hd__buf_2 output340 (.A(net340),
    .X(Tile_X0Y0_FrameData_O[23]));
 sky130_fd_sc_hd__buf_2 output341 (.A(net341),
    .X(Tile_X0Y0_FrameData_O[24]));
 sky130_fd_sc_hd__buf_2 output342 (.A(net342),
    .X(Tile_X0Y0_FrameData_O[25]));
 sky130_fd_sc_hd__buf_2 output343 (.A(net343),
    .X(Tile_X0Y0_FrameData_O[26]));
 sky130_fd_sc_hd__buf_2 output344 (.A(net344),
    .X(Tile_X0Y0_FrameData_O[27]));
 sky130_fd_sc_hd__buf_2 output345 (.A(net345),
    .X(Tile_X0Y0_FrameData_O[28]));
 sky130_fd_sc_hd__buf_2 output346 (.A(net346),
    .X(Tile_X0Y0_FrameData_O[29]));
 sky130_fd_sc_hd__buf_2 output347 (.A(net347),
    .X(Tile_X0Y0_FrameData_O[2]));
 sky130_fd_sc_hd__buf_2 output348 (.A(net348),
    .X(Tile_X0Y0_FrameData_O[30]));
 sky130_fd_sc_hd__buf_2 output349 (.A(net349),
    .X(Tile_X0Y0_FrameData_O[31]));
 sky130_fd_sc_hd__buf_2 output350 (.A(net350),
    .X(Tile_X0Y0_FrameData_O[3]));
 sky130_fd_sc_hd__buf_2 output351 (.A(net351),
    .X(Tile_X0Y0_FrameData_O[4]));
 sky130_fd_sc_hd__buf_2 output352 (.A(net352),
    .X(Tile_X0Y0_FrameData_O[5]));
 sky130_fd_sc_hd__buf_2 output353 (.A(net353),
    .X(Tile_X0Y0_FrameData_O[6]));
 sky130_fd_sc_hd__buf_2 output354 (.A(net354),
    .X(Tile_X0Y0_FrameData_O[7]));
 sky130_fd_sc_hd__buf_2 output355 (.A(net355),
    .X(Tile_X0Y0_FrameData_O[8]));
 sky130_fd_sc_hd__buf_2 output356 (.A(net356),
    .X(Tile_X0Y0_FrameData_O[9]));
 sky130_fd_sc_hd__buf_2 output357 (.A(net357),
    .X(Tile_X0Y0_FrameStrobe_O[0]));
 sky130_fd_sc_hd__buf_2 output358 (.A(net358),
    .X(Tile_X0Y0_FrameStrobe_O[10]));
 sky130_fd_sc_hd__buf_2 output359 (.A(net359),
    .X(Tile_X0Y0_FrameStrobe_O[11]));
 sky130_fd_sc_hd__buf_2 output360 (.A(net477),
    .X(Tile_X0Y0_FrameStrobe_O[12]));
 sky130_fd_sc_hd__buf_2 output361 (.A(net478),
    .X(Tile_X0Y0_FrameStrobe_O[13]));
 sky130_fd_sc_hd__buf_2 output362 (.A(net479),
    .X(Tile_X0Y0_FrameStrobe_O[14]));
 sky130_fd_sc_hd__buf_2 output363 (.A(net480),
    .X(Tile_X0Y0_FrameStrobe_O[15]));
 sky130_fd_sc_hd__buf_2 output364 (.A(net481),
    .X(Tile_X0Y0_FrameStrobe_O[16]));
 sky130_fd_sc_hd__buf_2 output365 (.A(net482),
    .X(Tile_X0Y0_FrameStrobe_O[17]));
 sky130_fd_sc_hd__buf_2 output366 (.A(net483),
    .X(Tile_X0Y0_FrameStrobe_O[18]));
 sky130_fd_sc_hd__buf_2 output367 (.A(net484),
    .X(Tile_X0Y0_FrameStrobe_O[19]));
 sky130_fd_sc_hd__buf_2 output368 (.A(net485),
    .X(Tile_X0Y0_FrameStrobe_O[1]));
 sky130_fd_sc_hd__buf_2 output369 (.A(net486),
    .X(Tile_X0Y0_FrameStrobe_O[2]));
 sky130_fd_sc_hd__buf_2 output370 (.A(net487),
    .X(Tile_X0Y0_FrameStrobe_O[3]));
 sky130_fd_sc_hd__buf_2 output371 (.A(net488),
    .X(Tile_X0Y0_FrameStrobe_O[4]));
 sky130_fd_sc_hd__buf_2 output372 (.A(net489),
    .X(Tile_X0Y0_FrameStrobe_O[5]));
 sky130_fd_sc_hd__buf_2 output373 (.A(net490),
    .X(Tile_X0Y0_FrameStrobe_O[6]));
 sky130_fd_sc_hd__buf_2 output374 (.A(net491),
    .X(Tile_X0Y0_FrameStrobe_O[7]));
 sky130_fd_sc_hd__buf_2 output375 (.A(net492),
    .X(Tile_X0Y0_FrameStrobe_O[8]));
 sky130_fd_sc_hd__buf_2 output376 (.A(net493),
    .X(Tile_X0Y0_FrameStrobe_O[9]));
 sky130_fd_sc_hd__buf_2 output377 (.A(net494),
    .X(Tile_X0Y0_N1BEG[0]));
 sky130_fd_sc_hd__buf_2 output378 (.A(net495),
    .X(Tile_X0Y0_N1BEG[1]));
 sky130_fd_sc_hd__buf_2 output379 (.A(net496),
    .X(Tile_X0Y0_N1BEG[2]));
 sky130_fd_sc_hd__buf_2 output380 (.A(net497),
    .X(Tile_X0Y0_N1BEG[3]));
 sky130_fd_sc_hd__buf_2 output381 (.A(net498),
    .X(Tile_X0Y0_N2BEG[0]));
 sky130_fd_sc_hd__buf_2 output382 (.A(net499),
    .X(Tile_X0Y0_N2BEG[1]));
 sky130_fd_sc_hd__buf_2 output383 (.A(net500),
    .X(Tile_X0Y0_N2BEG[2]));
 sky130_fd_sc_hd__buf_2 output384 (.A(net501),
    .X(Tile_X0Y0_N2BEG[3]));
 sky130_fd_sc_hd__buf_2 output385 (.A(net502),
    .X(Tile_X0Y0_N2BEG[4]));
 sky130_fd_sc_hd__buf_2 output386 (.A(net503),
    .X(Tile_X0Y0_N2BEG[5]));
 sky130_fd_sc_hd__buf_2 output387 (.A(net504),
    .X(Tile_X0Y0_N2BEG[6]));
 sky130_fd_sc_hd__buf_2 output388 (.A(net505),
    .X(Tile_X0Y0_N2BEG[7]));
 sky130_fd_sc_hd__buf_2 output389 (.A(net506),
    .X(Tile_X0Y0_N2BEGb[0]));
 sky130_fd_sc_hd__buf_2 output390 (.A(net507),
    .X(Tile_X0Y0_N2BEGb[1]));
 sky130_fd_sc_hd__buf_2 output391 (.A(net508),
    .X(Tile_X0Y0_N2BEGb[2]));
 sky130_fd_sc_hd__buf_2 output392 (.A(net509),
    .X(Tile_X0Y0_N2BEGb[3]));
 sky130_fd_sc_hd__buf_2 output393 (.A(net510),
    .X(Tile_X0Y0_N2BEGb[4]));
 sky130_fd_sc_hd__buf_2 output394 (.A(net511),
    .X(Tile_X0Y0_N2BEGb[5]));
 sky130_fd_sc_hd__buf_2 output395 (.A(net512),
    .X(Tile_X0Y0_N2BEGb[6]));
 sky130_fd_sc_hd__buf_2 output396 (.A(net513),
    .X(Tile_X0Y0_N2BEGb[7]));
 sky130_fd_sc_hd__buf_2 output397 (.A(net514),
    .X(Tile_X0Y0_N4BEG[0]));
 sky130_fd_sc_hd__buf_2 output398 (.A(net515),
    .X(Tile_X0Y0_N4BEG[10]));
 sky130_fd_sc_hd__buf_2 output399 (.A(net516),
    .X(Tile_X0Y0_N4BEG[11]));
 sky130_fd_sc_hd__buf_2 output400 (.A(net517),
    .X(Tile_X0Y0_N4BEG[12]));
 sky130_fd_sc_hd__buf_2 output401 (.A(net518),
    .X(Tile_X0Y0_N4BEG[13]));
 sky130_fd_sc_hd__buf_2 output402 (.A(net519),
    .X(Tile_X0Y0_N4BEG[14]));
 sky130_fd_sc_hd__buf_2 output403 (.A(net520),
    .X(Tile_X0Y0_N4BEG[15]));
 sky130_fd_sc_hd__buf_2 output404 (.A(net521),
    .X(Tile_X0Y0_N4BEG[1]));
 sky130_fd_sc_hd__buf_2 output405 (.A(net522),
    .X(Tile_X0Y0_N4BEG[2]));
 sky130_fd_sc_hd__buf_2 output406 (.A(net523),
    .X(Tile_X0Y0_N4BEG[3]));
 sky130_fd_sc_hd__buf_2 output407 (.A(net524),
    .X(Tile_X0Y0_N4BEG[4]));
 sky130_fd_sc_hd__buf_2 output408 (.A(net525),
    .X(Tile_X0Y0_N4BEG[5]));
 sky130_fd_sc_hd__buf_2 output409 (.A(net526),
    .X(Tile_X0Y0_N4BEG[6]));
 sky130_fd_sc_hd__buf_2 output410 (.A(net527),
    .X(Tile_X0Y0_N4BEG[7]));
 sky130_fd_sc_hd__buf_2 output411 (.A(net528),
    .X(Tile_X0Y0_N4BEG[8]));
 sky130_fd_sc_hd__buf_2 output412 (.A(net529),
    .X(Tile_X0Y0_N4BEG[9]));
 sky130_fd_sc_hd__buf_1 output413 (.A(net530),
    .X(Tile_X0Y0_UserCLKo));
 sky130_fd_sc_hd__buf_2 output414 (.A(net531),
    .X(Tile_X0Y0_W1BEG[0]));
 sky130_fd_sc_hd__buf_2 output415 (.A(net532),
    .X(Tile_X0Y0_W1BEG[1]));
 sky130_fd_sc_hd__buf_2 output416 (.A(net533),
    .X(Tile_X0Y0_W1BEG[2]));
 sky130_fd_sc_hd__buf_2 output417 (.A(net534),
    .X(Tile_X0Y0_W1BEG[3]));
 sky130_fd_sc_hd__buf_2 output418 (.A(net535),
    .X(Tile_X0Y0_W2BEG[0]));
 sky130_fd_sc_hd__buf_2 output419 (.A(net536),
    .X(Tile_X0Y0_W2BEG[1]));
 sky130_fd_sc_hd__buf_2 output420 (.A(net537),
    .X(Tile_X0Y0_W2BEG[2]));
 sky130_fd_sc_hd__buf_2 output421 (.A(net538),
    .X(Tile_X0Y0_W2BEG[3]));
 sky130_fd_sc_hd__buf_2 output422 (.A(net539),
    .X(Tile_X0Y0_W2BEG[4]));
 sky130_fd_sc_hd__buf_2 output423 (.A(net540),
    .X(Tile_X0Y0_W2BEG[5]));
 sky130_fd_sc_hd__buf_2 output424 (.A(net541),
    .X(Tile_X0Y0_W2BEG[6]));
 sky130_fd_sc_hd__buf_2 output425 (.A(net542),
    .X(Tile_X0Y0_W2BEG[7]));
 sky130_fd_sc_hd__buf_2 output426 (.A(net543),
    .X(Tile_X0Y0_W2BEGb[0]));
 sky130_fd_sc_hd__buf_2 output427 (.A(net544),
    .X(Tile_X0Y0_W2BEGb[1]));
 sky130_fd_sc_hd__buf_2 output428 (.A(net545),
    .X(Tile_X0Y0_W2BEGb[2]));
 sky130_fd_sc_hd__buf_2 output429 (.A(net546),
    .X(Tile_X0Y0_W2BEGb[3]));
 sky130_fd_sc_hd__buf_2 output430 (.A(net547),
    .X(Tile_X0Y0_W2BEGb[4]));
 sky130_fd_sc_hd__buf_2 output431 (.A(net548),
    .X(Tile_X0Y0_W2BEGb[5]));
 sky130_fd_sc_hd__buf_2 output432 (.A(net549),
    .X(Tile_X0Y0_W2BEGb[6]));
 sky130_fd_sc_hd__buf_2 output433 (.A(net550),
    .X(Tile_X0Y0_W2BEGb[7]));
 sky130_fd_sc_hd__buf_2 output434 (.A(net551),
    .X(Tile_X0Y0_W6BEG[0]));
 sky130_fd_sc_hd__buf_2 output435 (.A(net552),
    .X(Tile_X0Y0_W6BEG[10]));
 sky130_fd_sc_hd__buf_2 output436 (.A(net553),
    .X(Tile_X0Y0_W6BEG[11]));
 sky130_fd_sc_hd__buf_2 output437 (.A(net554),
    .X(Tile_X0Y0_W6BEG[1]));
 sky130_fd_sc_hd__buf_2 output438 (.A(net555),
    .X(Tile_X0Y0_W6BEG[2]));
 sky130_fd_sc_hd__buf_2 output439 (.A(net556),
    .X(Tile_X0Y0_W6BEG[3]));
 sky130_fd_sc_hd__buf_2 output440 (.A(net557),
    .X(Tile_X0Y0_W6BEG[4]));
 sky130_fd_sc_hd__buf_2 output441 (.A(net558),
    .X(Tile_X0Y0_W6BEG[5]));
 sky130_fd_sc_hd__buf_2 output442 (.A(net559),
    .X(Tile_X0Y0_W6BEG[6]));
 sky130_fd_sc_hd__buf_2 output443 (.A(net560),
    .X(Tile_X0Y0_W6BEG[7]));
 sky130_fd_sc_hd__buf_2 output444 (.A(net561),
    .X(Tile_X0Y0_W6BEG[8]));
 sky130_fd_sc_hd__buf_2 output445 (.A(net562),
    .X(Tile_X0Y0_W6BEG[9]));
 sky130_fd_sc_hd__buf_2 output446 (.A(net563),
    .X(Tile_X0Y0_WW4BEG[0]));
 sky130_fd_sc_hd__buf_2 output447 (.A(net564),
    .X(Tile_X0Y0_WW4BEG[10]));
 sky130_fd_sc_hd__buf_2 output448 (.A(net565),
    .X(Tile_X0Y0_WW4BEG[11]));
 sky130_fd_sc_hd__buf_2 output449 (.A(net566),
    .X(Tile_X0Y0_WW4BEG[12]));
 sky130_fd_sc_hd__buf_2 output450 (.A(net567),
    .X(Tile_X0Y0_WW4BEG[13]));
 sky130_fd_sc_hd__buf_2 output451 (.A(net568),
    .X(Tile_X0Y0_WW4BEG[14]));
 sky130_fd_sc_hd__buf_2 output452 (.A(net569),
    .X(Tile_X0Y0_WW4BEG[15]));
 sky130_fd_sc_hd__buf_2 output453 (.A(net570),
    .X(Tile_X0Y0_WW4BEG[1]));
 sky130_fd_sc_hd__buf_2 output454 (.A(net571),
    .X(Tile_X0Y0_WW4BEG[2]));
 sky130_fd_sc_hd__buf_2 output455 (.A(net572),
    .X(Tile_X0Y0_WW4BEG[3]));
 sky130_fd_sc_hd__buf_2 output456 (.A(net573),
    .X(Tile_X0Y0_WW4BEG[4]));
 sky130_fd_sc_hd__buf_2 output457 (.A(net574),
    .X(Tile_X0Y0_WW4BEG[5]));
 sky130_fd_sc_hd__buf_2 output458 (.A(net575),
    .X(Tile_X0Y0_WW4BEG[6]));
 sky130_fd_sc_hd__buf_2 output459 (.A(net576),
    .X(Tile_X0Y0_WW4BEG[7]));
 sky130_fd_sc_hd__buf_2 output460 (.A(net577),
    .X(Tile_X0Y0_WW4BEG[8]));
 sky130_fd_sc_hd__buf_2 output461 (.A(net578),
    .X(Tile_X0Y0_WW4BEG[9]));
 sky130_fd_sc_hd__buf_2 output462 (.A(net579),
    .X(Tile_X0Y1_FrameData_O[0]));
 sky130_fd_sc_hd__buf_2 output463 (.A(net580),
    .X(Tile_X0Y1_FrameData_O[10]));
 sky130_fd_sc_hd__buf_2 output464 (.A(net581),
    .X(Tile_X0Y1_FrameData_O[11]));
 sky130_fd_sc_hd__buf_2 output465 (.A(net582),
    .X(Tile_X0Y1_FrameData_O[12]));
 sky130_fd_sc_hd__buf_2 output466 (.A(net583),
    .X(Tile_X0Y1_FrameData_O[13]));
 sky130_fd_sc_hd__buf_2 output467 (.A(net584),
    .X(Tile_X0Y1_FrameData_O[14]));
 sky130_fd_sc_hd__buf_2 output468 (.A(net585),
    .X(Tile_X0Y1_FrameData_O[15]));
 sky130_fd_sc_hd__buf_2 output469 (.A(net586),
    .X(Tile_X0Y1_FrameData_O[16]));
 sky130_fd_sc_hd__buf_2 output470 (.A(net587),
    .X(Tile_X0Y1_FrameData_O[17]));
 sky130_fd_sc_hd__buf_2 output471 (.A(net588),
    .X(Tile_X0Y1_FrameData_O[18]));
 sky130_fd_sc_hd__buf_2 output472 (.A(net589),
    .X(Tile_X0Y1_FrameData_O[19]));
 sky130_fd_sc_hd__buf_2 output473 (.A(net590),
    .X(Tile_X0Y1_FrameData_O[1]));
 sky130_fd_sc_hd__buf_2 output474 (.A(net591),
    .X(Tile_X0Y1_FrameData_O[20]));
 sky130_fd_sc_hd__buf_2 output475 (.A(net592),
    .X(Tile_X0Y1_FrameData_O[21]));
 sky130_fd_sc_hd__buf_2 output476 (.A(net593),
    .X(Tile_X0Y1_FrameData_O[22]));
 sky130_fd_sc_hd__buf_2 output477 (.A(net594),
    .X(Tile_X0Y1_FrameData_O[23]));
 sky130_fd_sc_hd__buf_2 output478 (.A(net595),
    .X(Tile_X0Y1_FrameData_O[24]));
 sky130_fd_sc_hd__buf_2 output479 (.A(net596),
    .X(Tile_X0Y1_FrameData_O[25]));
 sky130_fd_sc_hd__buf_2 output480 (.A(net597),
    .X(Tile_X0Y1_FrameData_O[26]));
 sky130_fd_sc_hd__buf_2 output481 (.A(net598),
    .X(Tile_X0Y1_FrameData_O[27]));
 sky130_fd_sc_hd__buf_2 output482 (.A(net599),
    .X(Tile_X0Y1_FrameData_O[28]));
 sky130_fd_sc_hd__buf_2 output483 (.A(net600),
    .X(Tile_X0Y1_FrameData_O[29]));
 sky130_fd_sc_hd__buf_2 output484 (.A(net601),
    .X(Tile_X0Y1_FrameData_O[2]));
 sky130_fd_sc_hd__buf_2 output485 (.A(net602),
    .X(Tile_X0Y1_FrameData_O[30]));
 sky130_fd_sc_hd__buf_2 output486 (.A(net603),
    .X(Tile_X0Y1_FrameData_O[31]));
 sky130_fd_sc_hd__buf_2 output487 (.A(net604),
    .X(Tile_X0Y1_FrameData_O[3]));
 sky130_fd_sc_hd__buf_2 output488 (.A(net605),
    .X(Tile_X0Y1_FrameData_O[4]));
 sky130_fd_sc_hd__buf_2 output489 (.A(net606),
    .X(Tile_X0Y1_FrameData_O[5]));
 sky130_fd_sc_hd__buf_2 output490 (.A(net607),
    .X(Tile_X0Y1_FrameData_O[6]));
 sky130_fd_sc_hd__buf_2 output491 (.A(net608),
    .X(Tile_X0Y1_FrameData_O[7]));
 sky130_fd_sc_hd__buf_2 output492 (.A(net609),
    .X(Tile_X0Y1_FrameData_O[8]));
 sky130_fd_sc_hd__buf_2 output493 (.A(net610),
    .X(Tile_X0Y1_FrameData_O[9]));
 sky130_fd_sc_hd__buf_2 output494 (.A(net611),
    .X(Tile_X0Y1_S1BEG[0]));
 sky130_fd_sc_hd__buf_2 output495 (.A(net612),
    .X(Tile_X0Y1_S1BEG[1]));
 sky130_fd_sc_hd__buf_2 output496 (.A(net613),
    .X(Tile_X0Y1_S1BEG[2]));
 sky130_fd_sc_hd__buf_2 output497 (.A(net614),
    .X(Tile_X0Y1_S1BEG[3]));
 sky130_fd_sc_hd__buf_2 output498 (.A(net615),
    .X(Tile_X0Y1_S2BEG[0]));
 sky130_fd_sc_hd__buf_2 output499 (.A(net616),
    .X(Tile_X0Y1_S2BEG[1]));
 sky130_fd_sc_hd__buf_2 output500 (.A(net617),
    .X(Tile_X0Y1_S2BEG[2]));
 sky130_fd_sc_hd__buf_2 output501 (.A(net618),
    .X(Tile_X0Y1_S2BEG[3]));
 sky130_fd_sc_hd__buf_2 output502 (.A(net619),
    .X(Tile_X0Y1_S2BEG[4]));
 sky130_fd_sc_hd__buf_2 output503 (.A(net620),
    .X(Tile_X0Y1_S2BEG[5]));
 sky130_fd_sc_hd__buf_2 output504 (.A(net621),
    .X(Tile_X0Y1_S2BEG[6]));
 sky130_fd_sc_hd__buf_2 output505 (.A(net622),
    .X(Tile_X0Y1_S2BEG[7]));
 sky130_fd_sc_hd__buf_2 output506 (.A(net623),
    .X(Tile_X0Y1_S2BEGb[0]));
 sky130_fd_sc_hd__buf_2 output507 (.A(net624),
    .X(Tile_X0Y1_S2BEGb[1]));
 sky130_fd_sc_hd__buf_2 output508 (.A(net625),
    .X(Tile_X0Y1_S2BEGb[2]));
 sky130_fd_sc_hd__buf_2 output509 (.A(net626),
    .X(Tile_X0Y1_S2BEGb[3]));
 sky130_fd_sc_hd__buf_2 output510 (.A(net627),
    .X(Tile_X0Y1_S2BEGb[4]));
 sky130_fd_sc_hd__buf_2 output511 (.A(net628),
    .X(Tile_X0Y1_S2BEGb[5]));
 sky130_fd_sc_hd__buf_2 output512 (.A(net629),
    .X(Tile_X0Y1_S2BEGb[6]));
 sky130_fd_sc_hd__buf_2 output513 (.A(net630),
    .X(Tile_X0Y1_S2BEGb[7]));
 sky130_fd_sc_hd__buf_2 output514 (.A(net631),
    .X(Tile_X0Y1_S4BEG[0]));
 sky130_fd_sc_hd__buf_2 output515 (.A(net632),
    .X(Tile_X0Y1_S4BEG[10]));
 sky130_fd_sc_hd__buf_2 output516 (.A(net633),
    .X(Tile_X0Y1_S4BEG[11]));
 sky130_fd_sc_hd__buf_2 output517 (.A(net634),
    .X(Tile_X0Y1_S4BEG[12]));
 sky130_fd_sc_hd__buf_2 output518 (.A(net635),
    .X(Tile_X0Y1_S4BEG[13]));
 sky130_fd_sc_hd__buf_2 output519 (.A(net636),
    .X(Tile_X0Y1_S4BEG[14]));
 sky130_fd_sc_hd__buf_2 output520 (.A(net637),
    .X(Tile_X0Y1_S4BEG[15]));
 sky130_fd_sc_hd__buf_2 output521 (.A(net638),
    .X(Tile_X0Y1_S4BEG[1]));
 sky130_fd_sc_hd__buf_2 output522 (.A(net639),
    .X(Tile_X0Y1_S4BEG[2]));
 sky130_fd_sc_hd__buf_2 output523 (.A(net640),
    .X(Tile_X0Y1_S4BEG[3]));
 sky130_fd_sc_hd__buf_2 output524 (.A(net641),
    .X(Tile_X0Y1_S4BEG[4]));
 sky130_fd_sc_hd__buf_2 output525 (.A(net642),
    .X(Tile_X0Y1_S4BEG[5]));
 sky130_fd_sc_hd__buf_2 output526 (.A(net643),
    .X(Tile_X0Y1_S4BEG[6]));
 sky130_fd_sc_hd__buf_2 output527 (.A(net644),
    .X(Tile_X0Y1_S4BEG[7]));
 sky130_fd_sc_hd__buf_2 output528 (.A(net645),
    .X(Tile_X0Y1_S4BEG[8]));
 sky130_fd_sc_hd__buf_2 output529 (.A(net646),
    .X(Tile_X0Y1_S4BEG[9]));
 sky130_fd_sc_hd__buf_2 output530 (.A(net647),
    .X(Tile_X0Y1_W1BEG[0]));
 sky130_fd_sc_hd__buf_2 output531 (.A(net648),
    .X(Tile_X0Y1_W1BEG[1]));
 sky130_fd_sc_hd__buf_2 output532 (.A(net649),
    .X(Tile_X0Y1_W1BEG[2]));
 sky130_fd_sc_hd__buf_2 output533 (.A(net650),
    .X(Tile_X0Y1_W1BEG[3]));
 sky130_fd_sc_hd__buf_2 output534 (.A(net651),
    .X(Tile_X0Y1_W2BEG[0]));
 sky130_fd_sc_hd__buf_2 output535 (.A(net652),
    .X(Tile_X0Y1_W2BEG[1]));
 sky130_fd_sc_hd__buf_2 output536 (.A(net653),
    .X(Tile_X0Y1_W2BEG[2]));
 sky130_fd_sc_hd__buf_2 output537 (.A(net654),
    .X(Tile_X0Y1_W2BEG[3]));
 sky130_fd_sc_hd__buf_2 output538 (.A(net655),
    .X(Tile_X0Y1_W2BEG[4]));
 sky130_fd_sc_hd__buf_2 output539 (.A(net656),
    .X(Tile_X0Y1_W2BEG[5]));
 sky130_fd_sc_hd__buf_2 output540 (.A(net657),
    .X(Tile_X0Y1_W2BEG[6]));
 sky130_fd_sc_hd__buf_2 output541 (.A(net658),
    .X(Tile_X0Y1_W2BEG[7]));
 sky130_fd_sc_hd__buf_2 output542 (.A(net659),
    .X(Tile_X0Y1_W2BEGb[0]));
 sky130_fd_sc_hd__buf_2 output543 (.A(net660),
    .X(Tile_X0Y1_W2BEGb[1]));
 sky130_fd_sc_hd__buf_2 output544 (.A(net661),
    .X(Tile_X0Y1_W2BEGb[2]));
 sky130_fd_sc_hd__buf_2 output545 (.A(net662),
    .X(Tile_X0Y1_W2BEGb[3]));
 sky130_fd_sc_hd__buf_2 output546 (.A(net663),
    .X(Tile_X0Y1_W2BEGb[4]));
 sky130_fd_sc_hd__buf_2 output547 (.A(net664),
    .X(Tile_X0Y1_W2BEGb[5]));
 sky130_fd_sc_hd__buf_2 output548 (.A(net665),
    .X(Tile_X0Y1_W2BEGb[6]));
 sky130_fd_sc_hd__buf_2 output549 (.A(net666),
    .X(Tile_X0Y1_W2BEGb[7]));
 sky130_fd_sc_hd__buf_2 output550 (.A(net667),
    .X(Tile_X0Y1_W6BEG[0]));
 sky130_fd_sc_hd__buf_2 output551 (.A(net668),
    .X(Tile_X0Y1_W6BEG[10]));
 sky130_fd_sc_hd__buf_2 output552 (.A(net669),
    .X(Tile_X0Y1_W6BEG[11]));
 sky130_fd_sc_hd__buf_2 output553 (.A(net670),
    .X(Tile_X0Y1_W6BEG[1]));
 sky130_fd_sc_hd__buf_2 output554 (.A(net671),
    .X(Tile_X0Y1_W6BEG[2]));
 sky130_fd_sc_hd__buf_2 output555 (.A(net672),
    .X(Tile_X0Y1_W6BEG[3]));
 sky130_fd_sc_hd__buf_2 output556 (.A(net673),
    .X(Tile_X0Y1_W6BEG[4]));
 sky130_fd_sc_hd__buf_2 output557 (.A(net674),
    .X(Tile_X0Y1_W6BEG[5]));
 sky130_fd_sc_hd__buf_2 output558 (.A(net675),
    .X(Tile_X0Y1_W6BEG[6]));
 sky130_fd_sc_hd__buf_2 output559 (.A(net676),
    .X(Tile_X0Y1_W6BEG[7]));
 sky130_fd_sc_hd__buf_2 output560 (.A(net677),
    .X(Tile_X0Y1_W6BEG[8]));
 sky130_fd_sc_hd__buf_2 output561 (.A(net678),
    .X(Tile_X0Y1_W6BEG[9]));
 sky130_fd_sc_hd__buf_2 output562 (.A(net679),
    .X(Tile_X0Y1_WW4BEG[0]));
 sky130_fd_sc_hd__buf_2 output563 (.A(net680),
    .X(Tile_X0Y1_WW4BEG[10]));
 sky130_fd_sc_hd__buf_2 output564 (.A(net681),
    .X(Tile_X0Y1_WW4BEG[11]));
 sky130_fd_sc_hd__buf_2 output565 (.A(net682),
    .X(Tile_X0Y1_WW4BEG[12]));
 sky130_fd_sc_hd__buf_2 output566 (.A(net683),
    .X(Tile_X0Y1_WW4BEG[13]));
 sky130_fd_sc_hd__buf_2 output567 (.A(net684),
    .X(Tile_X0Y1_WW4BEG[14]));
 sky130_fd_sc_hd__buf_2 output568 (.A(net685),
    .X(Tile_X0Y1_WW4BEG[15]));
 sky130_fd_sc_hd__buf_2 output569 (.A(net686),
    .X(Tile_X0Y1_WW4BEG[1]));
 sky130_fd_sc_hd__buf_2 output570 (.A(net687),
    .X(Tile_X0Y1_WW4BEG[2]));
 sky130_fd_sc_hd__buf_2 output571 (.A(net688),
    .X(Tile_X0Y1_WW4BEG[3]));
 sky130_fd_sc_hd__buf_2 output572 (.A(net689),
    .X(Tile_X0Y1_WW4BEG[4]));
 sky130_fd_sc_hd__buf_2 output573 (.A(net690),
    .X(Tile_X0Y1_WW4BEG[5]));
 sky130_fd_sc_hd__buf_2 output574 (.A(net691),
    .X(Tile_X0Y1_WW4BEG[6]));
 sky130_fd_sc_hd__buf_2 output575 (.A(net692),
    .X(Tile_X0Y1_WW4BEG[7]));
 sky130_fd_sc_hd__buf_2 output576 (.A(net693),
    .X(Tile_X0Y1_WW4BEG[8]));
 sky130_fd_sc_hd__buf_2 output577 (.A(net694),
    .X(Tile_X0Y1_WW4BEG[9]));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_Tile_X0Y1_UserCLK (.A(Tile_X0Y1_UserCLK),
    .X(clknet_0_Tile_X0Y1_UserCLK));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_Tile_X0Y1_UserCLK (.A(clknet_0_Tile_X0Y1_UserCLK),
    .X(clknet_1_0__leaf_Tile_X0Y1_UserCLK));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_Tile_X0Y1_UserCLK (.A(clknet_0_Tile_X0Y1_UserCLK),
    .X(clknet_1_1__leaf_Tile_X0Y1_UserCLK));
 sky130_fd_sc_hd__diode_2 ANTENNA_1 (.DIODE(net256));
 sky130_fd_sc_hd__diode_2 ANTENNA_2 (.DIODE(net267));
 sky130_fd_sc_hd__diode_2 ANTENNA_3 (.DIODE(net268));
 sky130_fd_sc_hd__diode_2 ANTENNA_4 (.DIODE(net269));
 sky130_fd_sc_hd__diode_2 ANTENNA_5 (.DIODE(net272));
 sky130_fd_sc_hd__diode_2 ANTENNA_6 (.DIODE(net273));
 sky130_fd_sc_hd__diode_2 ANTENNA_7 (.DIODE(net276));
 sky130_fd_sc_hd__diode_2 ANTENNA_8 (.DIODE(net277));
 sky130_fd_sc_hd__diode_2 ANTENNA_9 (.DIODE(net278));
 sky130_fd_sc_hd__diode_2 ANTENNA_10 (.DIODE(net300));
 sky130_fd_sc_hd__diode_2 ANTENNA_11 (.DIODE(net301));
 sky130_fd_sc_hd__diode_2 ANTENNA_12 (.DIODE(net310));
 sky130_fd_sc_hd__diode_2 ANTENNA_13 (.DIODE(net323));
 sky130_fd_sc_hd__diode_2 ANTENNA_14 (.DIODE(\Tile_X0Y0_EF_SRAM_top.Inst_EF_SRAM_top_switch_matrix.S2BEG1 ));
 sky130_fd_sc_hd__diode_2 ANTENNA_15 (.DIODE(net326));
 sky130_fd_sc_hd__diode_2 ANTENNA_16 (.DIODE(net327));
 sky130_fd_sc_hd__diode_2 ANTENNA_17 (.DIODE(net333));
 sky130_fd_sc_hd__diode_2 ANTENNA_18 (.DIODE(net335));
 sky130_fd_sc_hd__diode_2 ANTENNA_19 (.DIODE(net338));
 sky130_fd_sc_hd__diode_2 ANTENNA_20 (.DIODE(net350));
 sky130_fd_sc_hd__diode_2 ANTENNA_21 (.DIODE(net356));
 sky130_fd_sc_hd__diode_2 ANTENNA_22 (.DIODE(net489));
 sky130_fd_sc_hd__diode_2 ANTENNA_23 (.DIODE(net498));
 sky130_fd_sc_hd__diode_2 ANTENNA_24 (.DIODE(net505));
 sky130_fd_sc_hd__diode_2 ANTENNA_25 (.DIODE(net506));
 sky130_fd_sc_hd__diode_2 ANTENNA_26 (.DIODE(net509));
 sky130_fd_sc_hd__diode_2 ANTENNA_27 (.DIODE(net514));
 sky130_fd_sc_hd__diode_2 ANTENNA_28 (.DIODE(net514));
 sky130_fd_sc_hd__diode_2 ANTENNA_29 (.DIODE(net514));
 sky130_fd_sc_hd__diode_2 ANTENNA_30 (.DIODE(net514));
 sky130_fd_sc_hd__diode_2 ANTENNA_31 (.DIODE(net514));
 sky130_fd_sc_hd__diode_2 ANTENNA_32 (.DIODE(net514));
 sky130_fd_sc_hd__diode_2 ANTENNA_33 (.DIODE(net514));
 sky130_fd_sc_hd__diode_2 ANTENNA_34 (.DIODE(net514));
 sky130_fd_sc_hd__diode_2 ANTENNA_35 (.DIODE(net514));
 sky130_fd_sc_hd__diode_2 ANTENNA_36 (.DIODE(net514));
 sky130_fd_sc_hd__diode_2 ANTENNA_37 (.DIODE(net515));
 sky130_fd_sc_hd__diode_2 ANTENNA_38 (.DIODE(net515));
 sky130_fd_sc_hd__diode_2 ANTENNA_39 (.DIODE(net515));
 sky130_fd_sc_hd__diode_2 ANTENNA_40 (.DIODE(net515));
 sky130_fd_sc_hd__diode_2 ANTENNA_41 (.DIODE(net517));
 sky130_fd_sc_hd__diode_2 ANTENNA_42 (.DIODE(net521));
 sky130_fd_sc_hd__diode_2 ANTENNA_43 (.DIODE(net521));
 sky130_fd_sc_hd__diode_2 ANTENNA_44 (.DIODE(net521));
 sky130_fd_sc_hd__diode_2 ANTENNA_45 (.DIODE(net521));
 sky130_fd_sc_hd__diode_2 ANTENNA_46 (.DIODE(net521));
 sky130_fd_sc_hd__diode_2 ANTENNA_47 (.DIODE(net521));
 sky130_fd_sc_hd__diode_2 ANTENNA_48 (.DIODE(net522));
 sky130_fd_sc_hd__diode_2 ANTENNA_49 (.DIODE(net523));
 sky130_fd_sc_hd__diode_2 ANTENNA_50 (.DIODE(net523));
 sky130_fd_sc_hd__diode_2 ANTENNA_51 (.DIODE(net523));
 sky130_fd_sc_hd__diode_2 ANTENNA_52 (.DIODE(net523));
 sky130_fd_sc_hd__diode_2 ANTENNA_53 (.DIODE(net523));
 sky130_fd_sc_hd__diode_2 ANTENNA_54 (.DIODE(net523));
 sky130_fd_sc_hd__diode_2 ANTENNA_55 (.DIODE(net523));
 sky130_fd_sc_hd__diode_2 ANTENNA_56 (.DIODE(net523));
 sky130_fd_sc_hd__diode_2 ANTENNA_57 (.DIODE(net523));
 sky130_fd_sc_hd__diode_2 ANTENNA_58 (.DIODE(net523));
 sky130_fd_sc_hd__diode_2 ANTENNA_59 (.DIODE(net525));
 sky130_fd_sc_hd__diode_2 ANTENNA_60 (.DIODE(net525));
 sky130_fd_sc_hd__diode_2 ANTENNA_61 (.DIODE(net525));
 sky130_fd_sc_hd__diode_2 ANTENNA_62 (.DIODE(net525));
 sky130_fd_sc_hd__diode_2 ANTENNA_63 (.DIODE(net525));
 sky130_fd_sc_hd__diode_2 ANTENNA_64 (.DIODE(net525));
 sky130_fd_sc_hd__diode_2 ANTENNA_65 (.DIODE(net526));
 sky130_fd_sc_hd__diode_2 ANTENNA_66 (.DIODE(net526));
 sky130_fd_sc_hd__diode_2 ANTENNA_67 (.DIODE(net526));
 sky130_fd_sc_hd__diode_2 ANTENNA_68 (.DIODE(net526));
 sky130_fd_sc_hd__diode_2 ANTENNA_69 (.DIODE(net526));
 sky130_fd_sc_hd__diode_2 ANTENNA_70 (.DIODE(net526));
 sky130_fd_sc_hd__diode_2 ANTENNA_71 (.DIODE(net526));
 sky130_fd_sc_hd__diode_2 ANTENNA_72 (.DIODE(net527));
 sky130_fd_sc_hd__diode_2 ANTENNA_73 (.DIODE(net527));
 sky130_fd_sc_hd__diode_2 ANTENNA_74 (.DIODE(net527));
 sky130_fd_sc_hd__diode_2 ANTENNA_75 (.DIODE(net527));
 sky130_fd_sc_hd__diode_2 ANTENNA_76 (.DIODE(net528));
 sky130_fd_sc_hd__diode_2 ANTENNA_77 (.DIODE(net535));
 sky130_fd_sc_hd__diode_2 ANTENNA_78 (.DIODE(net539));
 sky130_fd_sc_hd__diode_2 ANTENNA_79 (.DIODE(net547));
 sky130_fd_sc_hd__diode_2 ANTENNA_80 (.DIODE(Tile_X0Y1_FrameData[17]));
 sky130_fd_sc_hd__diode_2 ANTENNA_81 (.DIODE(Tile_X0Y1_FrameData[17]));
 sky130_fd_sc_hd__diode_2 ANTENNA_82 (.DIODE(Tile_X0Y1_FrameData[17]));
 sky130_fd_sc_hd__diode_2 ANTENNA_83 (.DIODE(Tile_X0Y1_FrameData[17]));
 sky130_fd_sc_hd__diode_2 ANTENNA_84 (.DIODE(net581));
 sky130_fd_sc_hd__diode_2 ANTENNA_85 (.DIODE(net583));
 sky130_fd_sc_hd__diode_2 ANTENNA_86 (.DIODE(net588));
 sky130_fd_sc_hd__diode_2 ANTENNA_87 (.DIODE(net592));
 sky130_fd_sc_hd__diode_2 ANTENNA_88 (.DIODE(net593));
 sky130_fd_sc_hd__diode_2 ANTENNA_89 (.DIODE(net593));
 sky130_fd_sc_hd__diode_2 ANTENNA_90 (.DIODE(net596));
 sky130_fd_sc_hd__diode_2 ANTENNA_91 (.DIODE(net597));
 sky130_fd_sc_hd__diode_2 ANTENNA_92 (.DIODE(net598));
 sky130_fd_sc_hd__diode_2 ANTENNA_93 (.DIODE(net599));
 sky130_fd_sc_hd__diode_2 ANTENNA_94 (.DIODE(net601));
 sky130_fd_sc_hd__diode_2 ANTENNA_95 (.DIODE(net606));
 sky130_fd_sc_hd__diode_2 ANTENNA_96 (.DIODE(Tile_X0Y1_FrameStrobe[10]));
 sky130_fd_sc_hd__diode_2 ANTENNA_97 (.DIODE(Tile_X0Y1_FrameStrobe[11]));
 sky130_fd_sc_hd__diode_2 ANTENNA_98 (.DIODE(Tile_X0Y1_FrameStrobe[12]));
 sky130_fd_sc_hd__diode_2 ANTENNA_99 (.DIODE(Tile_X0Y1_FrameStrobe[14]));
 sky130_fd_sc_hd__diode_2 ANTENNA_100 (.DIODE(Tile_X0Y1_FrameStrobe[15]));
 sky130_fd_sc_hd__diode_2 ANTENNA_101 (.DIODE(Tile_X0Y1_FrameStrobe[16]));
 sky130_fd_sc_hd__diode_2 ANTENNA_102 (.DIODE(Tile_X0Y1_FrameStrobe[17]));
 sky130_fd_sc_hd__diode_2 ANTENNA_103 (.DIODE(Tile_X0Y1_FrameStrobe[18]));
 sky130_fd_sc_hd__diode_2 ANTENNA_104 (.DIODE(Tile_X0Y1_FrameStrobe[18]));
 sky130_fd_sc_hd__diode_2 ANTENNA_105 (.DIODE(Tile_X0Y1_FrameStrobe[18]));
 sky130_fd_sc_hd__diode_2 ANTENNA_106 (.DIODE(Tile_X0Y1_FrameStrobe[18]));
 sky130_fd_sc_hd__diode_2 ANTENNA_107 (.DIODE(Tile_X0Y1_FrameStrobe[18]));
 sky130_fd_sc_hd__diode_2 ANTENNA_108 (.DIODE(Tile_X0Y1_FrameStrobe[18]));
 sky130_fd_sc_hd__diode_2 ANTENNA_109 (.DIODE(Tile_X0Y1_FrameStrobe[18]));
 sky130_fd_sc_hd__diode_2 ANTENNA_110 (.DIODE(Tile_X0Y1_FrameStrobe[18]));
 sky130_fd_sc_hd__diode_2 ANTENNA_111 (.DIODE(Tile_X0Y1_FrameStrobe[19]));
 sky130_fd_sc_hd__diode_2 ANTENNA_112 (.DIODE(Tile_X0Y1_FrameStrobe[19]));
 sky130_fd_sc_hd__diode_2 ANTENNA_113 (.DIODE(Tile_X0Y1_FrameStrobe[19]));
 sky130_fd_sc_hd__diode_2 ANTENNA_114 (.DIODE(Tile_X0Y1_FrameStrobe[19]));
 sky130_fd_sc_hd__diode_2 ANTENNA_115 (.DIODE(Tile_X0Y1_FrameStrobe[2]));
 sky130_fd_sc_hd__diode_2 ANTENNA_116 (.DIODE(Tile_X0Y1_FrameStrobe[4]));
 sky130_fd_sc_hd__diode_2 ANTENNA_117 (.DIODE(Tile_X0Y1_FrameStrobe[5]));
 sky130_fd_sc_hd__diode_2 ANTENNA_118 (.DIODE(Tile_X0Y1_FrameStrobe[6]));
 sky130_fd_sc_hd__diode_2 ANTENNA_119 (.DIODE(Tile_X0Y1_FrameStrobe[6]));
 sky130_fd_sc_hd__diode_2 ANTENNA_120 (.DIODE(Tile_X0Y1_FrameStrobe[7]));
 sky130_fd_sc_hd__diode_2 ANTENNA_121 (.DIODE(Tile_X0Y1_FrameStrobe[8]));
 sky130_fd_sc_hd__diode_2 ANTENNA_122 (.DIODE(Tile_X0Y1_FrameStrobe[8]));
 sky130_fd_sc_hd__diode_2 ANTENNA_123 (.DIODE(net615));
 sky130_fd_sc_hd__diode_2 ANTENNA_124 (.DIODE(net628));
 sky130_fd_sc_hd__diode_2 ANTENNA_125 (.DIODE(net635));
 sky130_fd_sc_hd__diode_2 ANTENNA_126 (.DIODE(net639));
 sky130_fd_sc_hd__diode_2 ANTENNA_127 (.DIODE(net640));
 sky130_fd_sc_hd__diode_2 ANTENNA_128 (.DIODE(net640));
 sky130_fd_sc_hd__diode_2 ANTENNA_129 (.DIODE(net642));
 sky130_fd_sc_hd__diode_2 ANTENNA_130 (.DIODE(net642));
 sky130_fd_sc_hd__diode_2 ANTENNA_131 (.DIODE(net642));
 sky130_fd_sc_hd__diode_2 ANTENNA_132 (.DIODE(net642));
 sky130_fd_sc_hd__diode_2 ANTENNA_133 (.DIODE(net642));
 sky130_fd_sc_hd__diode_2 ANTENNA_134 (.DIODE(net642));
 sky130_fd_sc_hd__diode_2 ANTENNA_135 (.DIODE(net642));
 sky130_fd_sc_hd__diode_2 ANTENNA_136 (.DIODE(net642));
 sky130_fd_sc_hd__diode_2 ANTENNA_137 (.DIODE(net642));
 sky130_fd_sc_hd__diode_2 ANTENNA_138 (.DIODE(net643));
 sky130_fd_sc_hd__diode_2 ANTENNA_139 (.DIODE(net643));
 sky130_fd_sc_hd__diode_2 ANTENNA_140 (.DIODE(net643));
 sky130_fd_sc_hd__diode_2 ANTENNA_141 (.DIODE(net646));
 sky130_fd_sc_hd__diode_2 ANTENNA_142 (.DIODE(net646));
 sky130_fd_sc_hd__diode_2 ANTENNA_143 (.DIODE(net646));
 sky130_fd_sc_hd__diode_2 ANTENNA_144 (.DIODE(net646));
 sky130_fd_sc_hd__diode_2 ANTENNA_145 (.DIODE(net646));
 sky130_fd_sc_hd__diode_2 ANTENNA_146 (.DIODE(net646));
 sky130_fd_sc_hd__diode_2 ANTENNA_147 (.DIODE(net646));
 sky130_fd_sc_hd__diode_2 ANTENNA_148 (.DIODE(net11));
 sky130_fd_sc_hd__diode_2 ANTENNA_149 (.DIODE(net21));
 sky130_fd_sc_hd__diode_2 ANTENNA_150 (.DIODE(net44));
 sky130_fd_sc_hd__diode_2 ANTENNA_151 (.DIODE(net44));
 sky130_fd_sc_hd__diode_2 ANTENNA_152 (.DIODE(net52));
 sky130_fd_sc_hd__diode_2 ANTENNA_153 (.DIODE(net52));
 sky130_fd_sc_hd__diode_2 ANTENNA_154 (.DIODE(net118));
 sky130_fd_sc_hd__diode_2 ANTENNA_155 (.DIODE(net118));
 sky130_fd_sc_hd__diode_2 ANTENNA_156 (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 ANTENNA_157 (.DIODE(net152));
 sky130_fd_sc_hd__diode_2 ANTENNA_158 (.DIODE(net152));
 sky130_fd_sc_hd__diode_2 ANTENNA_159 (.DIODE(net225));
 sky130_fd_sc_hd__diode_2 ANTENNA_160 (.DIODE(net524));
 sky130_fd_sc_hd__diode_2 ANTENNA_161 (.DIODE(net524));
 sky130_fd_sc_hd__diode_2 ANTENNA_162 (.DIODE(net524));
 sky130_fd_sc_hd__diode_2 ANTENNA_163 (.DIODE(net524));
 sky130_fd_sc_hd__diode_2 ANTENNA_164 (.DIODE(net524));
 sky130_fd_sc_hd__diode_2 ANTENNA_165 (.DIODE(net611));
 sky130_fd_sc_hd__diode_2 ANTENNA_166 (.DIODE(net631));
 sky130_fd_sc_hd__diode_2 ANTENNA_167 (.DIODE(net631));
 sky130_fd_sc_hd__diode_2 ANTENNA_168 (.DIODE(net644));
 sky130_fd_sc_hd__diode_2 ANTENNA_169 (.DIODE(net692));
 sky130_fd_sc_hd__diode_2 ANTENNA_170 (.DIODE(net25));
 sky130_fd_sc_hd__diode_2 ANTENNA_171 (.DIODE(net25));
 sky130_fd_sc_hd__diode_2 ANTENNA_172 (.DIODE(net25));
 sky130_fd_sc_hd__diode_2 ANTENNA_173 (.DIODE(net25));
 sky130_fd_sc_hd__diode_2 ANTENNA_174 (.DIODE(net45));
 sky130_fd_sc_hd__diode_2 ANTENNA_175 (.DIODE(net45));
 sky130_fd_sc_hd__diode_2 ANTENNA_176 (.DIODE(net45));
 sky130_fd_sc_hd__diode_2 ANTENNA_177 (.DIODE(net511));
 sky130_ef_sc_hd__decap_12 FILLER_0_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_213 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_229 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_287 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_33 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_38 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_50 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_86 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_92 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_104 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_137 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_158 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_162 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_181 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_203 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_227 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_245 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_109 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_213 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_227 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_231 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_321 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_30 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_42 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_52 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_227 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_231 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_239 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_227 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_235 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_321 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_123 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_135 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_147 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_227 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_235 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_239 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_153 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_165 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_173 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_188 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_227 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_321 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_35 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_203 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_227 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_256 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_268 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_37 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_159 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_193 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_203 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_211 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_227 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_259 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_271 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_283 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_321 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_119 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_131 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_143 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_189 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_213 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_220 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_247 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_139 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_157 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_321 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_137 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_193 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_213 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_153 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_188 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_219 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_231 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_321 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_150 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_167 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_179 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_246 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_321 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_64 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_147 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_193 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_220 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_229 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_287 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_290 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_308 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_109 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_202 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_282 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_321 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_214 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_229 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_242 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_254 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_65 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_81 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_100 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_121 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_226 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_230 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_256 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_268 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_280 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_321 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_89 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_241 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_121 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_168 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_265 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_321 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_150 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_99 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_110 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_144 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_156 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_174 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_321 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_155 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_205 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_221 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_235 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_260 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_61 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_98 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_124 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_138 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_147 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_155 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_246 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_260 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_321 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_23 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_52 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_101 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_193 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_201 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_216 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_229 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_254 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_311 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_11 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_25 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_195 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_224 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_248 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_321 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_23 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_36 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_72 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_84 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_151 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_158 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_170 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_194 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_223 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_231 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_246 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_286 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_321 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_78 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_90 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_156 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_35 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_59 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_119 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_139 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_150 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_154 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_188 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_203 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_234 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_238 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_274 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_321 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_35 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_39 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_71 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_75 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_200 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_249 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_262 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_301 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_313 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_50 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_58 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_71 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_83 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_127 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_161 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_288 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_300 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_321 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_13 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_72 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_80 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_17 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_35 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_88 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_118 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_157 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_321 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_39 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_146 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_238 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_262 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_13 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_121 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_129 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_159 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_176 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_188 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_205 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_329 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_78 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_90 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_110 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_121 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_160 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_215 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_264 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_301 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_313 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_44 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_129 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_159 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_232 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_244 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_248 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_282 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_22 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_71 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_79 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_95 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_99 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_146 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_191 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_203 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_327 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_44 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_56 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_62 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_161 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_200 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_208 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_238 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_246 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_272 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_17 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_52 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_119 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_131 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_146 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_220 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_279 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_311 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_323 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_153 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_195 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_203 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_234 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_18 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_30 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_101 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_117 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_148 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_160 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_216 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_274 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_300 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_312 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_320 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_16 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_72 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_232 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_244 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_259 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_284 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_28 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_52 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_78 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_90 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_110 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_137 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_155 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_189 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_202 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_212 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_249 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_171 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_175 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_190 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_248 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_259 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_285 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_43 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_73 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_104 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_134 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_146 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_154 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_200 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_212 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_231 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_14 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_63 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_67 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_82 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_159 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_171 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_192 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_265 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_285 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_38 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_50 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_198 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_210 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_234 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_314 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_80 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_206 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_218 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_224 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_321 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_13 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_28 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_52 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_87 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_17 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_284 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_237 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_327 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_112 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_138 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_147 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_160 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_287 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_329 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_64 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_76 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_88 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_133 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_162 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_175 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_188 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_200 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_208 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_222 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_263 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_284 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_308 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_320 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_47 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_112 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_76 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_88 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_108 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_129 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_241 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_317 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_71 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_105 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_117 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_178 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_190 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_33 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_65 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_86 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_143 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_199 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_223 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_314 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_88 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_148 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_160 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_221 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_261 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_6 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_144 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_184 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_196 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_263 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_267 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_314 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_58 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_66 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_80 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_91 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_103 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_115 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_161 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_174 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_221 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_261 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_300 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_12 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_54 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_79 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_91 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_249 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_267 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_317 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_61 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_73 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_165 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_183 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_200 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_214 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_248 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_267 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_275 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_290 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_13 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_25 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_37 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_52 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_84 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_96 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_164 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_201 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_237 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_14 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_73 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_78 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_66_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_112 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_66_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_171 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_224 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_266 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_290 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_22 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_34 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_90 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_134 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_146 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_243 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_258 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_9 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_22 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_65 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_103 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_190 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_212 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_224 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_36 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_48 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_88 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_100 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_119 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_139 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_152 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_198 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_241 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_254 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_11 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_105 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_117 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_159 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_171 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_185 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_227 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_290 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_43 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_89 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_110 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_121 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_193 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_211 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_311 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_327 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_37 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_64 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_103 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_139 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_147 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_234 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_246 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_329 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_71 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_75 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_88 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_94 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_145 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_202 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_222 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_238 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_250 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_262 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_270 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_66 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_78 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_116 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_127 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_187 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_199 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_317 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_174 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_275 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_287 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_77 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_109 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_163 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_166 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_173 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_243 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_255 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_317 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_115 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_174 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_215 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_234 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_79_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_94 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_133 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_157 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_160 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_185 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_249 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_263 ();
 sky130_fd_sc_hd__decap_3 FILLER_79_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_317 ();
 sky130_fd_sc_hd__decap_3 FILLER_79_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_58 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_70 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_157 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_162 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_168 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_176 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_195 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_251 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_290 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_35 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_59 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_95 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_135 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_147 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_159 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_200 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_290 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_327 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_33 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_73 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_80 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_147 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_159 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_171 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_178 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_184 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_188 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_227 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_240 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_269 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_290 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_78 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_90 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_240 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_252 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_260 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_317 ();
 sky130_fd_sc_hd__decap_3 FILLER_83_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_84_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_91 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_104 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_116 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_128 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_156 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_161 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_173 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_84_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_229 ();
 sky130_fd_sc_hd__decap_3 FILLER_84_235 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_244 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_259 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_284 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_329 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_85_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_37 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_54 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_73 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_95 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_107 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_126 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_150 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_162 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_198 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_222 ();
 sky130_fd_sc_hd__decap_3 FILLER_85_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_262 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_317 ();
 sky130_fd_sc_hd__decap_3 FILLER_85_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_36 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_42 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_83 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_116 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_138 ();
 sky130_fd_sc_hd__decap_3 FILLER_86_159 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_164 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_172 ();
 sky130_fd_sc_hd__decap_3 FILLER_86_185 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_261 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_273 ();
 sky130_fd_sc_hd__decap_3 FILLER_86_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_81 ();
 sky130_fd_sc_hd__decap_3 FILLER_87_95 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_122 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_148 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_166 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_189 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_203 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_239 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_279 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_308 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_320 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_88_7 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_88_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_35 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_59 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_71 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_118 ();
 sky130_fd_sc_hd__decap_8 FILLER_88_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_160 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_178 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_190 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_203 ();
 sky130_fd_sc_hd__decap_3 FILLER_88_215 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_88_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_88_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_89_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_89_137 ();
 sky130_fd_sc_hd__decap_3 FILLER_89_161 ();
 sky130_fd_sc_hd__decap_3 FILLER_89_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_184 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_196 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_200 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_222 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_243 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_255 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_267 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_314 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_59 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_71 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_153 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_90_193 ();
 sky130_fd_sc_hd__decap_3 FILLER_90_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_231 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_275 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_329 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_38 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_50 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_111 ();
 sky130_fd_sc_hd__decap_3 FILLER_91_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_161 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_191 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_249 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_254 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_262 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_317 ();
 sky130_fd_sc_hd__decap_3 FILLER_91_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_92_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_92_35 ();
 sky130_fd_sc_hd__decap_3 FILLER_92_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_67 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_71 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_92_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_117 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_92_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_161 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_260 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_272 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_284 ();
 sky130_fd_sc_hd__decap_8 FILLER_92_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_92_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_24 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_93_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_140 ();
 sky130_fd_sc_hd__decap_3 FILLER_93_148 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_267 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_317 ();
 sky130_fd_sc_hd__decap_3 FILLER_93_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_61 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_109 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_162 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_192 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_213 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_94_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_94_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_94_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_94_314 ();
 sky130_fd_sc_hd__decap_3 FILLER_94_322 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_95_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_90 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_129 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_142 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_150 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_95_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_177 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_297 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_318 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_324 ();
 sky130_fd_sc_hd__decap_3 FILLER_95_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_59 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_71 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_109 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_127 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_162 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_174 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_227 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_234 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_265 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_285 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_97_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_81 ();
 sky130_fd_sc_hd__decap_3 FILLER_97_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_137 ();
 sky130_fd_sc_hd__decap_3 FILLER_97_149 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_293 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_305 ();
 sky130_fd_sc_hd__decap_3 FILLER_97_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_98_7 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_160 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_174 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_221 ();
 sky130_fd_sc_hd__decap_3 FILLER_98_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_250 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_259 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_272 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_284 ();
 sky130_fd_sc_hd__decap_3 FILLER_98_292 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_52 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_67 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_91 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_95 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_99 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_124 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_148 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_160 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_179 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_187 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_201 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_99_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_99_241 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_284 ();
 sky130_fd_sc_hd__decap_3 FILLER_99_296 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_320 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_71 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_114 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_119 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_183 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_282 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_338 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_148 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_160 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_213 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_284 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_296 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_320 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_54 ();
 sky130_fd_sc_hd__decap_8 FILLER_102_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_102_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_124 ();
 sky130_fd_sc_hd__decap_8 FILLER_102_159 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_102_221 ();
 sky130_fd_sc_hd__decap_3 FILLER_102_229 ();
 sky130_fd_sc_hd__decap_8 FILLER_102_244 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_321 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_11 ();
 sky130_fd_sc_hd__decap_3 FILLER_103_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_75 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_87 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_117 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_130 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_103_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_249 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_103_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_293 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_317 ();
 sky130_fd_sc_hd__decap_3 FILLER_103_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_37 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_82 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_91 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_104 ();
 sky130_fd_sc_hd__decap_3 FILLER_104_112 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_161 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_173 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_104_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_277 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_23 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_35 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_105_81 ();
 sky130_fd_sc_hd__decap_3 FILLER_105_89 ();
 sky130_fd_sc_hd__decap_8 FILLER_105_104 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_105_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_105_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_105_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_293 ();
 sky130_fd_sc_hd__decap_8 FILLER_105_320 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_35 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_66 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_78 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_101 ();
 sky130_fd_sc_hd__decap_8 FILLER_106_132 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_202 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_214 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_226 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_283 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_106_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_52 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_132 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_144 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_156 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_107_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_107_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_248 ();
 sky130_fd_sc_hd__decap_8 FILLER_107_260 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_314 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_7 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_32 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_56 ();
 sky130_fd_sc_hd__decap_3 FILLER_108_68 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_83 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_106 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_136 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_154 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_108_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_108_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_338 ();
 sky130_fd_sc_hd__decap_3 FILLER_109_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_30 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_109_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_84 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_90 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_94 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_106 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_132 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_109_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_196 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_200 ();
 sky130_fd_sc_hd__decap_8 FILLER_109_216 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_243 ();
 sky130_fd_sc_hd__decap_8 FILLER_109_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_109_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_109_317 ();
 sky130_fd_sc_hd__decap_3 FILLER_109_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_110_7 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_33 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_80 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_123 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_192 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_230 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_110_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_40 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_60 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_72 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_96 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_102 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_149 ();
 sky130_fd_sc_hd__decap_8 FILLER_111_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_111_165 ();
 sky130_fd_sc_hd__decap_3 FILLER_111_181 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_196 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_202 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_314 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_112_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_56 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_72 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_91 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_116 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_128 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_157 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_112_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_217 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_258 ();
 sky130_fd_sc_hd__decap_3 FILLER_112_270 ();
 sky130_fd_sc_hd__decap_3 FILLER_112_297 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_112_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_43 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_113_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_150 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_162 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_258 ();
 sky130_fd_sc_hd__decap_8 FILLER_113_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_113_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_114_17 ();
 sky130_fd_sc_hd__decap_3 FILLER_114_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_109 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_148 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_160 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_172 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_184 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_114_265 ();
 sky130_fd_sc_hd__decap_8 FILLER_114_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_114_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_16 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_28 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_52 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_81 ();
 sky130_fd_sc_hd__decap_3 FILLER_115_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_115_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_150 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_162 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_249 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_115_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_37 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_49 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_61 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_116_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_159 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_16 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_117_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_98 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_157 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_162 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_185 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_204 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_216 ();
 sky130_fd_sc_hd__decap_3 FILLER_117_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_252 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_317 ();
 sky130_fd_sc_hd__decap_3 FILLER_117_325 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_54 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_60 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_106 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_118 ();
 sky130_fd_sc_hd__decap_8 FILLER_118_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_161 ();
 sky130_fd_sc_hd__decap_3 FILLER_118_175 ();
 sky130_fd_sc_hd__decap_8 FILLER_118_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_229 ();
 sky130_fd_sc_hd__decap_8 FILLER_118_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_118_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_287 ();
 sky130_fd_sc_hd__decap_8 FILLER_118_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_7 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_98 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_125 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_143 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_175 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_191 ();
 sky130_fd_sc_hd__decap_8 FILLER_119_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_119_266 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_306 ();
 sky130_fd_sc_hd__decap_8 FILLER_119_318 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_7 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_21 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_34 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_54 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_66 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_120_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_120_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_120_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_120_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_175 ();
 sky130_fd_sc_hd__decap_8 FILLER_120_188 ();
 sky130_fd_sc_hd__decap_8 FILLER_120_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_120_205 ();
 sky130_fd_sc_hd__decap_3 FILLER_120_220 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_226 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_230 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_287 ();
 sky130_fd_sc_hd__decap_8 FILLER_120_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_20 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_24 ();
 sky130_fd_sc_hd__decap_8 FILLER_121_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_121_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_81 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_132 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_144 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_156 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_175 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_184 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_196 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_220 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_245 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_266 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_306 ();
 sky130_fd_sc_hd__decap_8 FILLER_121_318 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_14 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_43 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_67 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_83 ();
 sky130_fd_sc_hd__decap_3 FILLER_122_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_100 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_136 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_154 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_161 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_173 ();
 sky130_fd_sc_hd__decap_8 FILLER_122_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_122_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_13 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_37 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_87 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_156 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_59 ();
 sky130_fd_sc_hd__decap_3 FILLER_124_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_124_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_124_161 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_168 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_321 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_16 ();
 sky130_fd_sc_hd__decap_8 FILLER_125_28 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_36 ();
 sky130_fd_sc_hd__decap_8 FILLER_125_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_65 ();
 sky130_fd_sc_hd__decap_3 FILLER_125_84 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_119 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_147 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_167 ();
 sky130_fd_sc_hd__decap_3 FILLER_125_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_245 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_257 ();
 sky130_fd_sc_hd__decap_8 FILLER_125_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_125_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_126_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_37 ();
 sky130_fd_sc_hd__decap_8 FILLER_126_56 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_64 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_82 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_103 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_115 ();
 sky130_fd_sc_hd__decap_3 FILLER_126_127 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_138 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_126_150 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_158 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_217 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_229 ();
 sky130_fd_sc_hd__decap_8 FILLER_126_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_126_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_280 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_292 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_321 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_9 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_21 ();
 sky130_fd_sc_hd__decap_8 FILLER_127_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_127_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_127_83 ();
 sky130_fd_sc_hd__decap_3 FILLER_127_91 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_106 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_127_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_183 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_257 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_59 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_71 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_159 ();
 sky130_fd_sc_hd__decap_3 FILLER_128_163 ();
 sky130_fd_sc_hd__decap_8 FILLER_128_170 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_195 ();
 sky130_fd_sc_hd__decap_3 FILLER_128_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_221 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_321 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_16 ();
 sky130_fd_sc_hd__decap_8 FILLER_129_28 ();
 sky130_fd_sc_hd__decap_8 FILLER_129_48 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_243 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_256 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_260 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_121 ();
 sky130_fd_sc_hd__decap_8 FILLER_130_132 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_221 ();
 sky130_fd_sc_hd__decap_3 FILLER_130_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_321 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_131_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_73 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_86 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_98 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_110 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_117 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_131_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_237 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_71 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_88 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_100 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_112 ();
 sky130_fd_sc_hd__decap_8 FILLER_132_155 ();
 sky130_fd_sc_hd__decap_3 FILLER_132_163 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_178 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_190 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_132_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_132_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_267 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_321 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_23 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_35 ();
 sky130_fd_sc_hd__decap_3 FILLER_133_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_96 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_150 ();
 sky130_fd_sc_hd__decap_8 FILLER_133_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_191 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_203 ();
 sky130_fd_sc_hd__decap_8 FILLER_133_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_134_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_134_104 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_119 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_130 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_144 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_168 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_213 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_226 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_277 ();
 sky130_fd_sc_hd__decap_3 FILLER_134_289 ();
 sky130_fd_sc_hd__decap_8 FILLER_134_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_321 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_17 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_135_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_135_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_135_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_180 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_192 ();
 sky130_fd_sc_hd__decap_8 FILLER_135_204 ();
 sky130_fd_sc_hd__decap_3 FILLER_135_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_240 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_252 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_13 ();
 sky130_fd_sc_hd__decap_3 FILLER_136_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_58 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_70 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_136_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_321 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_87 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_125 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_184 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_198 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_255 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_138_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_118 ();
 sky130_fd_sc_hd__decap_8 FILLER_138_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_159 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_246 ();
 sky130_fd_sc_hd__decap_8 FILLER_138_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_269 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_138_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_321 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_333 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_30 ();
 sky130_fd_sc_hd__decap_3 FILLER_139_42 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_87 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_145 ();
 sky130_fd_sc_hd__decap_8 FILLER_139_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_139_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_223 ();
 sky130_fd_sc_hd__decap_3 FILLER_139_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_242 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_254 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_58 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_82 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_91 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_165 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_140_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_218 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_230 ();
 sky130_fd_sc_hd__decap_8 FILLER_140_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_321 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_141_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_143 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_142_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_105 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_119 ();
 sky130_fd_sc_hd__decap_8 FILLER_142_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_321 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_321 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_12 ();
 sky130_fd_sc_hd__decap_8 FILLER_146_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_146_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_96 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_102 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_114 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_147 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_159 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_171 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_321 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_96 ();
 sky130_fd_sc_hd__decap_8 FILLER_147_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_13 ();
 sky130_fd_sc_hd__decap_3 FILLER_148_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_148_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_96 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_102 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_114 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_148_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_321 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_149_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_96 ();
 sky130_fd_sc_hd__decap_8 FILLER_149_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_149_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_83 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_91 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_96 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_102 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_106 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_112 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_115 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_150_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_321 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_151_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_151_81 ();
 sky130_fd_sc_hd__decap_3 FILLER_151_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_96 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_102 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_106 ();
 sky130_fd_sc_hd__decap_3 FILLER_151_117 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_122 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_146 ();
 sky130_fd_sc_hd__decap_8 FILLER_151_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_151_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_240 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_252 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_255 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_152_11 ();
 sky130_fd_sc_hd__decap_3 FILLER_152_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_83 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_91 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_96 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_106 ();
 sky130_fd_sc_hd__decap_3 FILLER_152_110 ();
 sky130_fd_sc_hd__decap_3 FILLER_152_117 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_122 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_244 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_248 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_256 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_260 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_284 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_321 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_34 ();
 sky130_fd_sc_hd__decap_8 FILLER_153_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_91 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_96 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_110 ();
 sky130_fd_sc_hd__decap_3 FILLER_153_117 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_122 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_146 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_158 ();
 sky130_fd_sc_hd__decap_3 FILLER_153_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_176 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_188 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_200 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_212 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_229 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_245 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_83 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_98 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_106 ();
 sky130_fd_sc_hd__decap_3 FILLER_154_110 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_119 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_122 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_257 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_269 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_154_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_321 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_33 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_38 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_50 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_67 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_86 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_98 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_134 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_143 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_158 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_162 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_201 ();
 sky130_fd_sc_hd__decap_8 FILLER_155_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_231 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_240 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_252 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_270 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_155_287 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_303 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_311 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_156_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_23 ();
 sky130_fd_sc_hd__decap_3 FILLER_156_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_156_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_156_117 ();
 sky130_fd_sc_hd__decap_3 FILLER_156_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_182 ();
 sky130_fd_sc_hd__decap_3 FILLER_156_211 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_231 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_156_277 ();
 sky130_fd_sc_hd__decap_3 FILLER_156_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_156_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_337 ();
endmodule
