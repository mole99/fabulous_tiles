magic
tech ihp-sg13g2
magscale 1 2
timestamp 1743692326
<< metal1 >>
rect 1152 9848 45216 9872
rect 1152 9808 3688 9848
rect 3728 9808 3770 9848
rect 3810 9808 3852 9848
rect 3892 9808 3934 9848
rect 3974 9808 4016 9848
rect 4056 9808 18808 9848
rect 18848 9808 18890 9848
rect 18930 9808 18972 9848
rect 19012 9808 19054 9848
rect 19094 9808 19136 9848
rect 19176 9808 33928 9848
rect 33968 9808 34010 9848
rect 34050 9808 34092 9848
rect 34132 9808 34174 9848
rect 34214 9808 34256 9848
rect 34296 9808 45216 9848
rect 1152 9784 45216 9808
rect 3387 9680 3429 9689
rect 3387 9640 3388 9680
rect 3428 9640 3429 9680
rect 3387 9631 3429 9640
rect 8187 9680 8229 9689
rect 8187 9640 8188 9680
rect 8228 9640 8229 9680
rect 8187 9631 8229 9640
rect 9915 9680 9957 9689
rect 9915 9640 9916 9680
rect 9956 9640 9957 9680
rect 9915 9631 9957 9640
rect 11547 9680 11589 9689
rect 11547 9640 11548 9680
rect 11588 9640 11589 9680
rect 11547 9631 11589 9640
rect 12315 9680 12357 9689
rect 12315 9640 12316 9680
rect 12356 9640 12357 9680
rect 12315 9631 12357 9640
rect 14523 9680 14565 9689
rect 14523 9640 14524 9680
rect 14564 9640 14565 9680
rect 14523 9631 14565 9640
rect 15675 9680 15717 9689
rect 15675 9640 15676 9680
rect 15716 9640 15717 9680
rect 15675 9631 15717 9640
rect 18075 9680 18117 9689
rect 18075 9640 18076 9680
rect 18116 9640 18117 9680
rect 18075 9631 18117 9640
rect 22011 9680 22053 9689
rect 22011 9640 22012 9680
rect 22052 9640 22053 9680
rect 22011 9631 22053 9640
rect 28443 9680 28485 9689
rect 28443 9640 28444 9680
rect 28484 9640 28485 9680
rect 28443 9631 28485 9640
rect 29211 9680 29253 9689
rect 29211 9640 29212 9680
rect 29252 9640 29253 9680
rect 29211 9631 29253 9640
rect 32283 9680 32325 9689
rect 32283 9640 32284 9680
rect 32324 9640 32325 9680
rect 32283 9631 32325 9640
rect 36891 9680 36933 9689
rect 36891 9640 36892 9680
rect 36932 9640 36933 9680
rect 36891 9631 36933 9640
rect 37275 9680 37317 9689
rect 37275 9640 37276 9680
rect 37316 9640 37317 9680
rect 37275 9631 37317 9640
rect 38811 9680 38853 9689
rect 38811 9640 38812 9680
rect 38852 9640 38853 9680
rect 38811 9631 38853 9640
rect 39195 9680 39237 9689
rect 39195 9640 39196 9680
rect 39236 9640 39237 9680
rect 39195 9631 39237 9640
rect 43227 9680 43269 9689
rect 43227 9640 43228 9680
rect 43268 9640 43269 9680
rect 43227 9631 43269 9640
rect 44379 9680 44421 9689
rect 44379 9640 44380 9680
rect 44420 9640 44421 9680
rect 44379 9631 44421 9640
rect 8331 9596 8373 9605
rect 8331 9556 8332 9596
rect 8372 9556 8373 9596
rect 8331 9547 8373 9556
rect 9531 9596 9573 9605
rect 9531 9556 9532 9596
rect 9572 9556 9573 9596
rect 9531 9547 9573 9556
rect 10059 9596 10101 9605
rect 10059 9556 10060 9596
rect 10100 9556 10101 9596
rect 10059 9547 10101 9556
rect 11931 9596 11973 9605
rect 11931 9556 11932 9596
rect 11972 9556 11973 9596
rect 11931 9547 11973 9556
rect 20139 9596 20181 9605
rect 20139 9556 20140 9596
rect 20180 9556 20181 9596
rect 20139 9547 20181 9556
rect 22107 9596 22149 9605
rect 22107 9556 22108 9596
rect 22148 9556 22149 9596
rect 22107 9547 22149 9556
rect 25227 9596 25269 9605
rect 25227 9556 25228 9596
rect 25268 9556 25269 9596
rect 25227 9547 25269 9556
rect 27531 9596 27573 9605
rect 27531 9556 27532 9596
rect 27572 9556 27573 9596
rect 27531 9547 27573 9556
rect 31803 9596 31845 9605
rect 31803 9556 31804 9596
rect 31844 9556 31845 9596
rect 31803 9547 31845 9556
rect 34299 9596 34341 9605
rect 34299 9556 34300 9596
rect 34340 9556 34341 9596
rect 34299 9547 34341 9556
rect 35595 9596 35637 9605
rect 35595 9556 35596 9596
rect 35636 9556 35637 9596
rect 35595 9547 35637 9556
rect 36123 9596 36165 9605
rect 36123 9556 36124 9596
rect 36164 9556 36165 9596
rect 36123 9547 36165 9556
rect 36507 9596 36549 9605
rect 36507 9556 36508 9596
rect 36548 9556 36549 9596
rect 36507 9547 36549 9556
rect 1227 9512 1269 9521
rect 1227 9472 1228 9512
rect 1268 9472 1269 9512
rect 1227 9463 1269 9472
rect 1611 9512 1653 9521
rect 1611 9472 1612 9512
rect 1652 9472 1653 9512
rect 1611 9463 1653 9472
rect 1995 9512 2037 9521
rect 1995 9472 1996 9512
rect 2036 9472 2037 9512
rect 1995 9463 2037 9472
rect 2379 9512 2421 9521
rect 2379 9472 2380 9512
rect 2420 9472 2421 9512
rect 2379 9463 2421 9472
rect 2763 9512 2805 9521
rect 2763 9472 2764 9512
rect 2804 9472 2805 9512
rect 2763 9463 2805 9472
rect 3147 9512 3189 9521
rect 3147 9472 3148 9512
rect 3188 9472 3189 9512
rect 3147 9463 3189 9472
rect 7947 9512 7989 9521
rect 7947 9472 7948 9512
rect 7988 9472 7989 9512
rect 7947 9463 7989 9472
rect 9291 9512 9333 9521
rect 9291 9472 9292 9512
rect 9332 9472 9333 9512
rect 9291 9463 9333 9472
rect 9675 9512 9717 9521
rect 9675 9472 9676 9512
rect 9716 9472 9717 9512
rect 9675 9463 9717 9472
rect 11307 9512 11349 9521
rect 11307 9472 11308 9512
rect 11348 9472 11349 9512
rect 11307 9463 11349 9472
rect 11691 9512 11733 9521
rect 11691 9472 11692 9512
rect 11732 9472 11733 9512
rect 11691 9463 11733 9472
rect 12075 9512 12117 9521
rect 12075 9472 12076 9512
rect 12116 9472 12117 9512
rect 12075 9463 12117 9472
rect 14283 9512 14325 9521
rect 14283 9472 14284 9512
rect 14324 9472 14325 9512
rect 14283 9463 14325 9472
rect 14667 9512 14709 9521
rect 14667 9472 14668 9512
rect 14708 9472 14709 9512
rect 14667 9463 14709 9472
rect 15051 9512 15093 9521
rect 15051 9472 15052 9512
rect 15092 9472 15093 9512
rect 15051 9463 15093 9472
rect 15435 9512 15477 9521
rect 15435 9472 15436 9512
rect 15476 9472 15477 9512
rect 15435 9463 15477 9472
rect 15819 9512 15861 9521
rect 15819 9472 15820 9512
rect 15860 9472 15861 9512
rect 15819 9463 15861 9472
rect 17835 9512 17877 9521
rect 17835 9472 17836 9512
rect 17876 9472 17877 9512
rect 17835 9463 17877 9472
rect 18795 9512 18837 9521
rect 18795 9472 18796 9512
rect 18836 9472 18837 9512
rect 18795 9463 18837 9472
rect 18987 9512 19029 9521
rect 18987 9472 18988 9512
rect 19028 9472 19029 9512
rect 18987 9463 19029 9472
rect 20619 9512 20661 9521
rect 20619 9472 20620 9512
rect 20660 9472 20661 9512
rect 20619 9463 20661 9472
rect 21195 9512 21237 9521
rect 21195 9472 21196 9512
rect 21236 9472 21237 9512
rect 21195 9463 21237 9472
rect 21339 9512 21381 9521
rect 21339 9472 21340 9512
rect 21380 9472 21381 9512
rect 21339 9463 21381 9472
rect 21579 9512 21621 9521
rect 21579 9472 21580 9512
rect 21620 9472 21621 9512
rect 21579 9463 21621 9472
rect 21771 9512 21813 9521
rect 21771 9472 21772 9512
rect 21812 9472 21813 9512
rect 21771 9463 21813 9472
rect 22347 9512 22389 9521
rect 22347 9472 22348 9512
rect 22388 9472 22389 9512
rect 22347 9463 22389 9472
rect 22731 9512 22773 9521
rect 22731 9472 22732 9512
rect 22772 9472 22773 9512
rect 22731 9463 22773 9472
rect 23115 9512 23157 9521
rect 23115 9472 23116 9512
rect 23156 9472 23157 9512
rect 23115 9463 23157 9472
rect 23307 9512 23349 9521
rect 23307 9472 23308 9512
rect 23348 9472 23349 9512
rect 23307 9463 23349 9472
rect 23883 9512 23925 9521
rect 23883 9472 23884 9512
rect 23924 9472 23925 9512
rect 23883 9463 23925 9472
rect 24267 9512 24309 9521
rect 24267 9472 24268 9512
rect 24308 9472 24309 9512
rect 24267 9463 24309 9472
rect 25611 9512 25653 9521
rect 25611 9472 25612 9512
rect 25652 9472 25653 9512
rect 25611 9463 25653 9472
rect 25803 9512 25845 9521
rect 25803 9472 25804 9512
rect 25844 9472 25845 9512
rect 25803 9463 25845 9472
rect 26187 9512 26229 9521
rect 26187 9472 26188 9512
rect 26228 9472 26229 9512
rect 26187 9463 26229 9472
rect 27915 9512 27957 9521
rect 27915 9472 27916 9512
rect 27956 9472 27957 9512
rect 27915 9463 27957 9472
rect 28299 9512 28341 9521
rect 28299 9472 28300 9512
rect 28340 9472 28341 9512
rect 28299 9463 28341 9472
rect 28683 9512 28725 9521
rect 28683 9472 28684 9512
rect 28724 9472 28725 9512
rect 28683 9463 28725 9472
rect 29067 9512 29109 9521
rect 29067 9472 29068 9512
rect 29108 9472 29109 9512
rect 29067 9463 29109 9472
rect 29451 9512 29493 9521
rect 29451 9472 29452 9512
rect 29492 9472 29493 9512
rect 29451 9463 29493 9472
rect 29835 9512 29877 9521
rect 29835 9472 29836 9512
rect 29876 9472 29877 9512
rect 29835 9463 29877 9472
rect 30027 9512 30069 9521
rect 30027 9472 30028 9512
rect 30068 9472 30069 9512
rect 30027 9463 30069 9472
rect 30603 9512 30645 9521
rect 30603 9472 30604 9512
rect 30644 9472 30645 9512
rect 30603 9463 30645 9472
rect 30987 9512 31029 9521
rect 30987 9472 30988 9512
rect 31028 9472 31029 9512
rect 30987 9463 31029 9472
rect 31371 9512 31413 9521
rect 31371 9472 31372 9512
rect 31412 9472 31413 9512
rect 31371 9463 31413 9472
rect 31563 9512 31605 9521
rect 31563 9472 31564 9512
rect 31604 9472 31605 9512
rect 31563 9463 31605 9472
rect 32139 9512 32181 9521
rect 32139 9472 32140 9512
rect 32180 9472 32181 9512
rect 32139 9463 32181 9472
rect 32523 9512 32565 9521
rect 32523 9472 32524 9512
rect 32564 9472 32565 9512
rect 32523 9463 32565 9472
rect 34539 9512 34581 9521
rect 34539 9472 34540 9512
rect 34580 9472 34581 9512
rect 34539 9463 34581 9472
rect 35979 9512 36021 9521
rect 35979 9472 35980 9512
rect 36020 9472 36021 9512
rect 35979 9463 36021 9472
rect 36363 9512 36405 9521
rect 36363 9472 36364 9512
rect 36404 9472 36405 9512
rect 36363 9463 36405 9472
rect 36747 9512 36789 9521
rect 36747 9472 36748 9512
rect 36788 9472 36789 9512
rect 36747 9463 36789 9472
rect 37131 9512 37173 9521
rect 37131 9472 37132 9512
rect 37172 9472 37173 9512
rect 37131 9463 37173 9472
rect 37515 9512 37557 9521
rect 37515 9472 37516 9512
rect 37556 9472 37557 9512
rect 37515 9463 37557 9472
rect 37899 9512 37941 9521
rect 37899 9472 37900 9512
rect 37940 9472 37941 9512
rect 37899 9463 37941 9472
rect 38283 9512 38325 9521
rect 38283 9472 38284 9512
rect 38324 9472 38325 9512
rect 38283 9463 38325 9472
rect 38667 9512 38709 9521
rect 38667 9472 38668 9512
rect 38708 9472 38709 9512
rect 38667 9463 38709 9472
rect 39051 9512 39093 9521
rect 39051 9472 39052 9512
rect 39092 9472 39093 9512
rect 39051 9463 39093 9472
rect 39435 9512 39477 9521
rect 39435 9472 39436 9512
rect 39476 9472 39477 9512
rect 39435 9463 39477 9472
rect 39819 9512 39861 9521
rect 39819 9472 39820 9512
rect 39860 9472 39861 9512
rect 39819 9463 39861 9472
rect 41019 9512 41061 9521
rect 41019 9472 41020 9512
rect 41060 9472 41061 9512
rect 41019 9463 41061 9472
rect 41259 9512 41301 9521
rect 41259 9472 41260 9512
rect 41300 9472 41301 9512
rect 41259 9463 41301 9472
rect 42603 9512 42645 9521
rect 42603 9472 42604 9512
rect 42644 9472 42645 9512
rect 42603 9463 42645 9472
rect 42987 9512 43029 9521
rect 42987 9472 42988 9512
rect 43028 9472 43029 9512
rect 42987 9463 43029 9472
rect 43467 9512 43509 9521
rect 43467 9472 43468 9512
rect 43508 9472 43509 9512
rect 43467 9463 43509 9472
rect 43755 9512 43797 9521
rect 43755 9472 43756 9512
rect 43796 9472 43797 9512
rect 43755 9463 43797 9472
rect 44139 9512 44181 9521
rect 44139 9472 44140 9512
rect 44180 9472 44181 9512
rect 44139 9463 44181 9472
rect 44523 9512 44565 9521
rect 44523 9472 44524 9512
rect 44564 9472 44565 9512
rect 44523 9463 44565 9472
rect 45099 9512 45141 9521
rect 45099 9472 45100 9512
rect 45140 9472 45141 9512
rect 45099 9463 45141 9472
rect 6315 9428 6357 9437
rect 6315 9388 6316 9428
rect 6356 9388 6357 9428
rect 6315 9379 6357 9388
rect 7555 9428 7613 9429
rect 9003 9428 9045 9437
rect 10731 9428 10773 9437
rect 7555 9388 7564 9428
rect 7604 9388 7613 9428
rect 7555 9387 7613 9388
rect 8715 9419 8757 9428
rect 8715 9379 8716 9419
rect 8756 9379 8757 9419
rect 9003 9388 9004 9428
rect 9044 9388 9045 9428
rect 9003 9379 9045 9388
rect 10443 9419 10485 9428
rect 10443 9379 10444 9419
rect 10484 9379 10485 9419
rect 10731 9388 10732 9428
rect 10772 9388 10773 9428
rect 10731 9379 10773 9388
rect 12643 9428 12701 9429
rect 12643 9388 12652 9428
rect 12692 9388 12701 9428
rect 12643 9387 12701 9388
rect 13899 9428 13941 9437
rect 13899 9388 13900 9428
rect 13940 9388 13941 9428
rect 13899 9379 13941 9388
rect 16203 9428 16245 9437
rect 16203 9388 16204 9428
rect 16244 9388 16245 9428
rect 16203 9379 16245 9388
rect 17443 9428 17501 9429
rect 17443 9388 17452 9428
rect 17492 9388 17501 9428
rect 17443 9387 17501 9388
rect 19467 9428 19509 9437
rect 19467 9388 19468 9428
rect 19508 9388 19509 9428
rect 19467 9379 19509 9388
rect 19738 9428 19796 9429
rect 19738 9388 19747 9428
rect 19787 9388 19796 9428
rect 19738 9387 19796 9388
rect 24555 9428 24597 9437
rect 24555 9388 24556 9428
rect 24596 9388 24597 9428
rect 24555 9379 24597 9388
rect 24826 9428 24884 9429
rect 24826 9388 24835 9428
rect 24875 9388 24884 9428
rect 24826 9387 24884 9388
rect 26859 9428 26901 9437
rect 26859 9388 26860 9428
rect 26900 9388 26901 9428
rect 26859 9379 26901 9388
rect 27106 9428 27164 9429
rect 27106 9388 27115 9428
rect 27155 9388 27164 9428
rect 27106 9387 27164 9388
rect 27226 9428 27284 9429
rect 27226 9388 27235 9428
rect 27275 9388 27284 9428
rect 27226 9387 27284 9388
rect 32715 9428 32757 9437
rect 32715 9388 32716 9428
rect 32756 9388 32757 9428
rect 32715 9379 32757 9388
rect 33955 9428 34013 9429
rect 33955 9388 33964 9428
rect 34004 9388 34013 9428
rect 33955 9387 34013 9388
rect 34923 9428 34965 9437
rect 34923 9388 34924 9428
rect 34964 9388 34965 9428
rect 34923 9379 34965 9388
rect 35194 9428 35252 9429
rect 35194 9388 35203 9428
rect 35243 9388 35252 9428
rect 35194 9387 35252 9388
rect 8715 9370 8757 9379
rect 10443 9370 10485 9379
rect 8619 9344 8661 9353
rect 8619 9304 8620 9344
rect 8660 9304 8661 9344
rect 8619 9295 8661 9304
rect 10347 9344 10389 9353
rect 10347 9304 10348 9344
rect 10388 9304 10389 9344
rect 10347 9295 10389 9304
rect 12459 9344 12501 9353
rect 12459 9304 12460 9344
rect 12500 9304 12501 9344
rect 12459 9295 12501 9304
rect 14907 9344 14949 9353
rect 14907 9304 14908 9344
rect 14948 9304 14949 9344
rect 14907 9295 14949 9304
rect 19851 9344 19893 9353
rect 19851 9304 19852 9344
rect 19892 9304 19893 9344
rect 19851 9295 19893 9304
rect 20859 9344 20901 9353
rect 20859 9304 20860 9344
rect 20900 9304 20901 9344
rect 20859 9295 20901 9304
rect 23547 9344 23589 9353
rect 23547 9304 23548 9344
rect 23588 9304 23589 9344
rect 23547 9295 23589 9304
rect 24939 9344 24981 9353
rect 24939 9304 24940 9344
rect 24980 9304 24981 9344
rect 24939 9295 24981 9304
rect 29595 9344 29637 9353
rect 29595 9304 29596 9344
rect 29636 9304 29637 9344
rect 29595 9295 29637 9304
rect 30267 9344 30309 9353
rect 30267 9304 30268 9344
rect 30308 9304 30309 9344
rect 30267 9295 30309 9304
rect 35307 9344 35349 9353
rect 35307 9304 35308 9344
rect 35348 9304 35349 9344
rect 35307 9295 35349 9304
rect 39579 9344 39621 9353
rect 39579 9304 39580 9344
rect 39620 9304 39621 9344
rect 39579 9295 39621 9304
rect 44763 9344 44805 9353
rect 44763 9304 44764 9344
rect 44804 9304 44805 9344
rect 44763 9295 44805 9304
rect 1467 9260 1509 9269
rect 1467 9220 1468 9260
rect 1508 9220 1509 9260
rect 1467 9211 1509 9220
rect 1851 9260 1893 9269
rect 1851 9220 1852 9260
rect 1892 9220 1893 9260
rect 1851 9211 1893 9220
rect 2235 9260 2277 9269
rect 2235 9220 2236 9260
rect 2276 9220 2277 9260
rect 2235 9211 2277 9220
rect 2619 9260 2661 9269
rect 2619 9220 2620 9260
rect 2660 9220 2661 9260
rect 2619 9211 2661 9220
rect 3003 9260 3045 9269
rect 3003 9220 3004 9260
rect 3044 9220 3045 9260
rect 3003 9211 3045 9220
rect 7755 9260 7797 9269
rect 7755 9220 7756 9260
rect 7796 9220 7797 9260
rect 7755 9211 7797 9220
rect 15291 9260 15333 9269
rect 15291 9220 15292 9260
rect 15332 9220 15333 9260
rect 15291 9211 15333 9220
rect 16059 9260 16101 9269
rect 16059 9220 16060 9260
rect 16100 9220 16101 9260
rect 16059 9211 16101 9220
rect 17643 9260 17685 9269
rect 17643 9220 17644 9260
rect 17684 9220 17685 9260
rect 17643 9211 17685 9220
rect 18411 9260 18453 9269
rect 18411 9220 18412 9260
rect 18452 9220 18453 9260
rect 18411 9211 18453 9220
rect 18555 9260 18597 9269
rect 18555 9220 18556 9260
rect 18596 9220 18597 9260
rect 18555 9211 18597 9220
rect 19227 9260 19269 9269
rect 19227 9220 19228 9260
rect 19268 9220 19269 9260
rect 19227 9211 19269 9220
rect 20955 9260 20997 9269
rect 20955 9220 20956 9260
rect 20996 9220 20997 9260
rect 20955 9211 20997 9220
rect 22491 9260 22533 9269
rect 22491 9220 22492 9260
rect 22532 9220 22533 9260
rect 22491 9211 22533 9220
rect 22875 9260 22917 9269
rect 22875 9220 22876 9260
rect 22916 9220 22917 9260
rect 22875 9211 22917 9220
rect 23643 9260 23685 9269
rect 23643 9220 23644 9260
rect 23684 9220 23685 9260
rect 23643 9211 23685 9220
rect 24027 9260 24069 9269
rect 24027 9220 24028 9260
rect 24068 9220 24069 9260
rect 24027 9211 24069 9220
rect 25371 9260 25413 9269
rect 25371 9220 25372 9260
rect 25412 9220 25413 9260
rect 25371 9211 25413 9220
rect 26043 9260 26085 9269
rect 26043 9220 26044 9260
rect 26084 9220 26085 9260
rect 26043 9211 26085 9220
rect 26427 9260 26469 9269
rect 26427 9220 26428 9260
rect 26468 9220 26469 9260
rect 26427 9211 26469 9220
rect 27675 9260 27717 9269
rect 27675 9220 27676 9260
rect 27716 9220 27717 9260
rect 27675 9211 27717 9220
rect 28059 9260 28101 9269
rect 28059 9220 28060 9260
rect 28100 9220 28101 9260
rect 28059 9211 28101 9220
rect 28827 9260 28869 9269
rect 28827 9220 28828 9260
rect 28868 9220 28869 9260
rect 28827 9211 28869 9220
rect 30363 9260 30405 9269
rect 30363 9220 30364 9260
rect 30404 9220 30405 9260
rect 30363 9211 30405 9220
rect 30747 9260 30789 9269
rect 30747 9220 30748 9260
rect 30788 9220 30789 9260
rect 30747 9211 30789 9220
rect 31131 9260 31173 9269
rect 31131 9220 31132 9260
rect 31172 9220 31173 9260
rect 31131 9211 31173 9220
rect 31899 9260 31941 9269
rect 31899 9220 31900 9260
rect 31940 9220 31941 9260
rect 31899 9211 31941 9220
rect 34155 9260 34197 9269
rect 34155 9220 34156 9260
rect 34196 9220 34197 9260
rect 34155 9211 34197 9220
rect 35739 9260 35781 9269
rect 35739 9220 35740 9260
rect 35780 9220 35781 9260
rect 35739 9211 35781 9220
rect 37659 9260 37701 9269
rect 37659 9220 37660 9260
rect 37700 9220 37701 9260
rect 37659 9211 37701 9220
rect 38043 9260 38085 9269
rect 38043 9220 38044 9260
rect 38084 9220 38085 9260
rect 38043 9211 38085 9220
rect 38427 9260 38469 9269
rect 38427 9220 38428 9260
rect 38468 9220 38469 9260
rect 38427 9211 38469 9220
rect 40186 9260 40244 9261
rect 40186 9220 40195 9260
rect 40235 9220 40244 9260
rect 40186 9219 40244 9220
rect 40474 9260 40532 9261
rect 40474 9220 40483 9260
rect 40523 9220 40532 9260
rect 40474 9219 40532 9220
rect 40762 9260 40820 9261
rect 40762 9220 40771 9260
rect 40811 9220 40820 9260
rect 40762 9219 40820 9220
rect 41434 9260 41492 9261
rect 41434 9220 41443 9260
rect 41483 9220 41492 9260
rect 41434 9219 41492 9220
rect 41722 9260 41780 9261
rect 41722 9220 41731 9260
rect 41771 9220 41780 9260
rect 41722 9219 41780 9220
rect 42010 9260 42068 9261
rect 42010 9220 42019 9260
rect 42059 9220 42068 9260
rect 42010 9219 42068 9220
rect 42298 9260 42356 9261
rect 42298 9220 42307 9260
rect 42347 9220 42356 9260
rect 42298 9219 42356 9220
rect 42843 9260 42885 9269
rect 42843 9220 42844 9260
rect 42884 9220 42885 9260
rect 42843 9211 42885 9220
rect 43450 9260 43508 9261
rect 43450 9220 43459 9260
rect 43499 9220 43508 9260
rect 43450 9219 43508 9220
rect 43995 9260 44037 9269
rect 43995 9220 43996 9260
rect 44036 9220 44037 9260
rect 43995 9211 44037 9220
rect 44859 9260 44901 9269
rect 44859 9220 44860 9260
rect 44900 9220 44901 9260
rect 44859 9211 44901 9220
rect 1152 9092 45216 9116
rect 1152 9052 4928 9092
rect 4968 9052 5010 9092
rect 5050 9052 5092 9092
rect 5132 9052 5174 9092
rect 5214 9052 5256 9092
rect 5296 9052 20048 9092
rect 20088 9052 20130 9092
rect 20170 9052 20212 9092
rect 20252 9052 20294 9092
rect 20334 9052 20376 9092
rect 20416 9052 35168 9092
rect 35208 9052 35250 9092
rect 35290 9052 35332 9092
rect 35372 9052 35414 9092
rect 35454 9052 35496 9092
rect 35536 9052 45216 9092
rect 1152 9028 45216 9052
rect 1467 8924 1509 8933
rect 1467 8884 1468 8924
rect 1508 8884 1509 8924
rect 1467 8875 1509 8884
rect 2619 8924 2661 8933
rect 2619 8884 2620 8924
rect 2660 8884 2661 8924
rect 2619 8875 2661 8884
rect 8235 8924 8277 8933
rect 8235 8884 8236 8924
rect 8276 8884 8277 8924
rect 8235 8875 8277 8884
rect 10731 8924 10773 8933
rect 10731 8884 10732 8924
rect 10772 8884 10773 8924
rect 10731 8875 10773 8884
rect 13563 8924 13605 8933
rect 13563 8884 13564 8924
rect 13604 8884 13605 8924
rect 13563 8875 13605 8884
rect 13947 8924 13989 8933
rect 13947 8884 13948 8924
rect 13988 8884 13989 8924
rect 13947 8875 13989 8884
rect 15531 8924 15573 8933
rect 15531 8884 15532 8924
rect 15572 8884 15573 8924
rect 15531 8875 15573 8884
rect 16155 8924 16197 8933
rect 16155 8884 16156 8924
rect 16196 8884 16197 8924
rect 16155 8875 16197 8884
rect 17739 8924 17781 8933
rect 17739 8884 17740 8924
rect 17780 8884 17781 8924
rect 17739 8875 17781 8884
rect 22635 8924 22677 8933
rect 22635 8884 22636 8924
rect 22676 8884 22677 8924
rect 22635 8875 22677 8884
rect 26283 8924 26325 8933
rect 26283 8884 26284 8924
rect 26324 8884 26325 8924
rect 26283 8875 26325 8884
rect 32667 8924 32709 8933
rect 32667 8884 32668 8924
rect 32708 8884 32709 8924
rect 32667 8875 32709 8884
rect 35259 8924 35301 8933
rect 35259 8884 35260 8924
rect 35300 8884 35301 8924
rect 35259 8875 35301 8884
rect 35979 8924 36021 8933
rect 35979 8884 35980 8924
rect 36020 8884 36021 8924
rect 35979 8875 36021 8884
rect 38331 8924 38373 8933
rect 38331 8884 38332 8924
rect 38372 8884 38373 8924
rect 38331 8875 38373 8884
rect 40923 8924 40965 8933
rect 40923 8884 40924 8924
rect 40964 8884 40965 8924
rect 40923 8875 40965 8884
rect 41355 8924 41397 8933
rect 41355 8884 41356 8924
rect 41396 8884 41397 8924
rect 41355 8875 41397 8884
rect 41722 8924 41780 8925
rect 41722 8884 41731 8924
rect 41771 8884 41780 8924
rect 41722 8883 41780 8884
rect 42795 8924 42837 8933
rect 42795 8884 42796 8924
rect 42836 8884 42837 8924
rect 42795 8875 42837 8884
rect 43707 8924 43749 8933
rect 43707 8884 43708 8924
rect 43748 8884 43749 8924
rect 43707 8875 43749 8884
rect 44379 8924 44421 8933
rect 44379 8884 44380 8924
rect 44420 8884 44421 8924
rect 44379 8875 44421 8884
rect 5835 8840 5877 8849
rect 5835 8800 5836 8840
rect 5876 8800 5877 8840
rect 5835 8791 5877 8800
rect 11211 8840 11253 8849
rect 11211 8800 11212 8840
rect 11252 8800 11253 8840
rect 11211 8791 11253 8800
rect 13179 8840 13221 8849
rect 13179 8800 13180 8840
rect 13220 8800 13221 8840
rect 13179 8791 13221 8800
rect 18267 8840 18309 8849
rect 18267 8800 18268 8840
rect 18308 8800 18309 8840
rect 18267 8791 18309 8800
rect 27243 8840 27285 8849
rect 27243 8800 27244 8840
rect 27284 8800 27285 8840
rect 27243 8791 27285 8800
rect 28347 8840 28389 8849
rect 28347 8800 28348 8840
rect 28388 8800 28389 8840
rect 28347 8791 28389 8800
rect 30699 8840 30741 8849
rect 30699 8800 30700 8840
rect 30740 8800 30741 8840
rect 30699 8791 30741 8800
rect 32571 8840 32613 8849
rect 32571 8800 32572 8840
rect 32612 8800 32613 8840
rect 32571 8791 32613 8800
rect 33675 8840 33717 8849
rect 33675 8800 33676 8840
rect 33716 8800 33717 8840
rect 33675 8791 33717 8800
rect 34827 8840 34869 8849
rect 34827 8800 34828 8840
rect 34868 8800 34869 8840
rect 34827 8791 34869 8800
rect 35163 8840 35205 8849
rect 35163 8800 35164 8840
rect 35204 8800 35205 8840
rect 35163 8791 35205 8800
rect 39387 8840 39429 8849
rect 39387 8800 39388 8840
rect 39428 8800 39429 8840
rect 39387 8791 39429 8800
rect 43323 8840 43365 8849
rect 43323 8800 43324 8840
rect 43364 8800 43365 8840
rect 43323 8791 43365 8800
rect 4395 8756 4437 8765
rect 6795 8756 6837 8765
rect 8986 8756 9044 8757
rect 4395 8716 4396 8756
rect 4436 8716 4437 8756
rect 4395 8707 4437 8716
rect 5643 8747 5685 8756
rect 5643 8707 5644 8747
rect 5684 8707 5685 8747
rect 6795 8716 6796 8756
rect 6836 8716 6837 8756
rect 6795 8707 6837 8716
rect 8043 8747 8085 8756
rect 8043 8707 8044 8747
rect 8084 8707 8085 8747
rect 8986 8716 8995 8756
rect 9035 8716 9044 8756
rect 8986 8715 9044 8716
rect 9099 8756 9141 8765
rect 9099 8716 9100 8756
rect 9140 8716 9141 8756
rect 9099 8707 9141 8716
rect 9483 8756 9525 8765
rect 12651 8756 12693 8765
rect 9483 8716 9484 8756
rect 9524 8716 9525 8756
rect 9483 8707 9525 8716
rect 10059 8747 10101 8756
rect 10059 8707 10060 8747
rect 10100 8707 10101 8747
rect 5643 8698 5685 8707
rect 8043 8698 8085 8707
rect 10059 8698 10101 8707
rect 10539 8747 10581 8756
rect 10539 8707 10540 8747
rect 10580 8707 10581 8747
rect 10539 8698 10581 8707
rect 11403 8747 11445 8756
rect 11403 8707 11404 8747
rect 11444 8707 11445 8747
rect 12651 8716 12652 8756
rect 12692 8716 12693 8756
rect 12651 8707 12693 8716
rect 14091 8756 14133 8765
rect 16299 8756 16341 8765
rect 18861 8756 18903 8765
rect 14091 8716 14092 8756
rect 14132 8716 14133 8756
rect 14091 8707 14133 8716
rect 15339 8747 15381 8756
rect 15339 8707 15340 8747
rect 15380 8707 15381 8747
rect 16299 8716 16300 8756
rect 16340 8716 16341 8756
rect 16299 8707 16341 8716
rect 17547 8747 17589 8756
rect 17547 8707 17548 8747
rect 17588 8707 17589 8747
rect 18861 8716 18862 8756
rect 18902 8716 18903 8756
rect 18861 8707 18903 8716
rect 18987 8756 19029 8765
rect 18987 8716 18988 8756
rect 19028 8716 19029 8756
rect 18987 8707 19029 8716
rect 19371 8756 19413 8765
rect 19371 8716 19372 8756
rect 19412 8716 19413 8756
rect 19371 8707 19413 8716
rect 19934 8756 19992 8757
rect 20890 8756 20948 8757
rect 19934 8716 19943 8756
rect 19983 8716 19992 8756
rect 19934 8715 19992 8716
rect 20427 8747 20469 8756
rect 20427 8707 20428 8747
rect 20468 8707 20469 8747
rect 20890 8716 20899 8756
rect 20939 8716 20948 8756
rect 20890 8715 20948 8716
rect 21003 8756 21045 8765
rect 21003 8716 21004 8756
rect 21044 8716 21045 8756
rect 21003 8707 21045 8716
rect 21387 8756 21429 8765
rect 22827 8756 22869 8765
rect 21387 8716 21388 8756
rect 21428 8716 21429 8756
rect 21387 8707 21429 8716
rect 21963 8747 22005 8756
rect 21963 8707 21964 8747
rect 22004 8707 22005 8747
rect 11403 8698 11445 8707
rect 15339 8698 15381 8707
rect 17547 8698 17589 8707
rect 20427 8698 20469 8707
rect 21963 8698 22005 8707
rect 22443 8747 22485 8756
rect 22443 8707 22444 8747
rect 22484 8707 22485 8747
rect 22827 8716 22828 8756
rect 22868 8716 22869 8756
rect 22827 8707 22869 8716
rect 24538 8756 24596 8757
rect 24538 8716 24547 8756
rect 24587 8716 24596 8756
rect 24538 8715 24596 8716
rect 24651 8756 24693 8765
rect 24651 8716 24652 8756
rect 24692 8716 24693 8756
rect 24071 8714 24129 8715
rect 22443 8698 22485 8707
rect 1227 8672 1269 8681
rect 1227 8632 1228 8672
rect 1268 8632 1269 8672
rect 1227 8623 1269 8632
rect 1611 8672 1653 8681
rect 1611 8632 1612 8672
rect 1652 8632 1653 8672
rect 1611 8623 1653 8632
rect 1995 8672 2037 8681
rect 1995 8632 1996 8672
rect 2036 8632 2037 8672
rect 1995 8623 2037 8632
rect 2235 8672 2277 8681
rect 2235 8632 2236 8672
rect 2276 8632 2277 8672
rect 2235 8623 2277 8632
rect 2379 8672 2421 8681
rect 2379 8632 2380 8672
rect 2420 8632 2421 8672
rect 2379 8623 2421 8632
rect 8523 8672 8565 8681
rect 8523 8632 8524 8672
rect 8564 8632 8565 8672
rect 8523 8623 8565 8632
rect 8763 8672 8805 8681
rect 8763 8632 8764 8672
rect 8804 8632 8805 8672
rect 8763 8623 8805 8632
rect 9579 8672 9621 8681
rect 9579 8632 9580 8672
rect 9620 8632 9621 8672
rect 9579 8623 9621 8632
rect 12939 8672 12981 8681
rect 12939 8632 12940 8672
rect 12980 8632 12981 8672
rect 12939 8623 12981 8632
rect 13323 8672 13365 8681
rect 13323 8632 13324 8672
rect 13364 8632 13365 8672
rect 13323 8623 13365 8632
rect 13707 8672 13749 8681
rect 13707 8632 13708 8672
rect 13748 8632 13749 8672
rect 13707 8623 13749 8632
rect 15915 8672 15957 8681
rect 15915 8632 15916 8672
rect 15956 8632 15957 8672
rect 15915 8623 15957 8632
rect 18027 8672 18069 8681
rect 18027 8632 18028 8672
rect 18068 8632 18069 8672
rect 18027 8623 18069 8632
rect 18411 8672 18453 8681
rect 18411 8632 18412 8672
rect 18452 8632 18453 8672
rect 18411 8623 18453 8632
rect 18651 8672 18693 8681
rect 18651 8632 18652 8672
rect 18692 8632 18693 8672
rect 18651 8623 18693 8632
rect 19467 8672 19509 8681
rect 19467 8632 19468 8672
rect 19508 8632 19509 8672
rect 19467 8623 19509 8632
rect 20650 8672 20708 8673
rect 20650 8632 20659 8672
rect 20699 8632 20708 8672
rect 20650 8631 20708 8632
rect 21483 8672 21525 8681
rect 24071 8674 24080 8714
rect 24120 8674 24129 8714
rect 24651 8707 24693 8716
rect 25035 8756 25077 8765
rect 26859 8756 26901 8765
rect 25035 8716 25036 8756
rect 25076 8716 25077 8756
rect 25035 8707 25077 8716
rect 25611 8747 25653 8756
rect 25611 8707 25612 8747
rect 25652 8707 25653 8747
rect 25611 8698 25653 8707
rect 26091 8747 26133 8756
rect 26091 8707 26092 8747
rect 26132 8707 26133 8747
rect 26859 8716 26860 8756
rect 26900 8716 26901 8756
rect 26859 8707 26901 8716
rect 27130 8756 27188 8757
rect 30507 8756 30549 8765
rect 32139 8756 32181 8765
rect 27130 8716 27139 8756
rect 27179 8716 27188 8756
rect 27130 8715 27188 8716
rect 29259 8747 29301 8756
rect 29259 8707 29260 8747
rect 29300 8707 29301 8747
rect 30507 8716 30508 8756
rect 30548 8716 30549 8756
rect 30507 8707 30549 8716
rect 30891 8747 30933 8756
rect 30891 8707 30892 8747
rect 30932 8707 30933 8747
rect 32139 8716 32140 8756
rect 32180 8716 32181 8756
rect 32139 8707 32181 8716
rect 33291 8756 33333 8765
rect 33291 8716 33292 8756
rect 33332 8716 33333 8756
rect 33291 8707 33333 8716
rect 33562 8756 33620 8757
rect 33562 8716 33571 8756
rect 33611 8716 33620 8756
rect 33562 8715 33620 8716
rect 34443 8756 34485 8765
rect 34443 8716 34444 8756
rect 34484 8716 34485 8756
rect 34443 8707 34485 8716
rect 34714 8756 34772 8757
rect 37419 8756 37461 8765
rect 34714 8716 34723 8756
rect 34763 8716 34772 8756
rect 34714 8715 34772 8716
rect 36171 8747 36213 8756
rect 36171 8707 36172 8747
rect 36212 8707 36213 8747
rect 37419 8716 37420 8756
rect 37460 8716 37461 8756
rect 37419 8707 37461 8716
rect 42891 8756 42933 8765
rect 42891 8716 42892 8756
rect 42932 8716 42933 8756
rect 42891 8707 42933 8716
rect 44715 8756 44757 8765
rect 44715 8716 44716 8756
rect 44756 8716 44757 8756
rect 44715 8707 44757 8716
rect 26091 8698 26133 8707
rect 29259 8698 29301 8707
rect 30891 8698 30933 8707
rect 36171 8698 36213 8707
rect 24071 8673 24129 8674
rect 21483 8632 21484 8672
rect 21524 8632 21525 8672
rect 21483 8623 21525 8632
rect 25131 8672 25173 8681
rect 25131 8632 25132 8672
rect 25172 8632 25173 8672
rect 25131 8623 25173 8632
rect 27675 8672 27717 8681
rect 27675 8632 27676 8672
rect 27716 8632 27717 8672
rect 27675 8623 27717 8632
rect 27915 8672 27957 8681
rect 27915 8632 27916 8672
rect 27956 8632 27957 8672
rect 27915 8623 27957 8632
rect 28107 8672 28149 8681
rect 28107 8632 28108 8672
rect 28148 8632 28149 8672
rect 28107 8623 28149 8632
rect 28683 8672 28725 8681
rect 28683 8632 28684 8672
rect 28724 8632 28725 8672
rect 28683 8623 28725 8632
rect 29050 8672 29108 8673
rect 29050 8632 29059 8672
rect 29099 8632 29108 8672
rect 29050 8631 29108 8632
rect 32331 8672 32373 8681
rect 32331 8632 32332 8672
rect 32372 8632 32373 8672
rect 32331 8623 32373 8632
rect 32907 8672 32949 8681
rect 32907 8632 32908 8672
rect 32948 8632 32949 8672
rect 32907 8623 32949 8632
rect 35499 8672 35541 8681
rect 35499 8632 35500 8672
rect 35540 8632 35541 8672
rect 35499 8623 35541 8632
rect 37563 8672 37605 8681
rect 37563 8632 37564 8672
rect 37604 8632 37605 8672
rect 37563 8623 37605 8632
rect 37803 8672 37845 8681
rect 37803 8632 37804 8672
rect 37844 8632 37845 8672
rect 37803 8623 37845 8632
rect 37947 8672 37989 8681
rect 37947 8632 37948 8672
rect 37988 8632 37989 8672
rect 37947 8623 37989 8632
rect 38187 8672 38229 8681
rect 38187 8632 38188 8672
rect 38228 8632 38229 8672
rect 38187 8623 38229 8632
rect 38571 8672 38613 8681
rect 38571 8632 38572 8672
rect 38612 8632 38613 8672
rect 38571 8623 38613 8632
rect 38715 8672 38757 8681
rect 38715 8632 38716 8672
rect 38756 8632 38757 8672
rect 38715 8623 38757 8632
rect 38955 8672 38997 8681
rect 38955 8632 38956 8672
rect 38996 8632 38997 8672
rect 38955 8623 38997 8632
rect 39147 8672 39189 8681
rect 39147 8632 39148 8672
rect 39188 8632 39189 8672
rect 39147 8623 39189 8632
rect 39531 8672 39573 8681
rect 39531 8632 39532 8672
rect 39572 8632 39573 8672
rect 39531 8623 39573 8632
rect 39867 8672 39909 8681
rect 39867 8632 39868 8672
rect 39908 8632 39909 8672
rect 39867 8623 39909 8632
rect 40107 8672 40149 8681
rect 40107 8632 40108 8672
rect 40148 8632 40149 8672
rect 40107 8623 40149 8632
rect 40491 8672 40533 8681
rect 40491 8632 40492 8672
rect 40532 8632 40533 8672
rect 40491 8623 40533 8632
rect 40779 8672 40821 8681
rect 40779 8632 40780 8672
rect 40820 8632 40821 8672
rect 40779 8623 40821 8632
rect 41163 8672 41205 8681
rect 41163 8632 41164 8672
rect 41204 8632 41205 8672
rect 41163 8623 41205 8632
rect 42027 8672 42069 8681
rect 42027 8632 42028 8672
rect 42068 8632 42069 8672
rect 42027 8623 42069 8632
rect 42315 8672 42357 8681
rect 42315 8632 42316 8672
rect 42356 8632 42357 8672
rect 42315 8623 42357 8632
rect 42603 8672 42645 8681
rect 42603 8632 42604 8672
rect 42644 8632 42645 8672
rect 42603 8623 42645 8632
rect 43083 8672 43125 8681
rect 43083 8632 43084 8672
rect 43124 8632 43125 8672
rect 43083 8623 43125 8632
rect 43467 8672 43509 8681
rect 43467 8632 43468 8672
rect 43508 8632 43509 8672
rect 43467 8623 43509 8632
rect 43947 8672 43989 8681
rect 43947 8632 43948 8672
rect 43988 8632 43989 8672
rect 43947 8623 43989 8632
rect 44139 8672 44181 8681
rect 44139 8632 44140 8672
rect 44180 8632 44181 8672
rect 44139 8623 44181 8632
rect 44907 8672 44949 8681
rect 44907 8632 44908 8672
rect 44948 8632 44949 8672
rect 44907 8623 44949 8632
rect 28443 8588 28485 8597
rect 28443 8548 28444 8588
rect 28484 8548 28485 8588
rect 28443 8539 28485 8548
rect 39771 8588 39813 8597
rect 39771 8548 39772 8588
rect 39812 8548 39813 8588
rect 39771 8539 39813 8548
rect 1851 8504 1893 8513
rect 1851 8464 1852 8504
rect 1892 8464 1893 8504
rect 1851 8455 1893 8464
rect 24267 8504 24309 8513
rect 24267 8464 24268 8504
rect 24308 8464 24309 8504
rect 24267 8455 24309 8464
rect 27531 8504 27573 8513
rect 27531 8464 27532 8504
rect 27572 8464 27573 8504
rect 27531 8455 27573 8464
rect 33963 8504 34005 8513
rect 33963 8464 33964 8504
rect 34004 8464 34005 8504
rect 33963 8455 34005 8464
rect 45147 8504 45189 8513
rect 45147 8464 45148 8504
rect 45188 8464 45189 8504
rect 45147 8455 45189 8464
rect 1152 8336 45216 8360
rect 1152 8296 3688 8336
rect 3728 8296 3770 8336
rect 3810 8296 3852 8336
rect 3892 8296 3934 8336
rect 3974 8296 4016 8336
rect 4056 8296 18808 8336
rect 18848 8296 18890 8336
rect 18930 8296 18972 8336
rect 19012 8296 19054 8336
rect 19094 8296 19136 8336
rect 19176 8296 33928 8336
rect 33968 8296 34010 8336
rect 34050 8296 34092 8336
rect 34132 8296 34174 8336
rect 34214 8296 34256 8336
rect 34296 8296 45216 8336
rect 1152 8272 45216 8296
rect 4347 8168 4389 8177
rect 4347 8128 4348 8168
rect 4388 8128 4389 8168
rect 4347 8119 4389 8128
rect 10251 8168 10293 8177
rect 10251 8128 10252 8168
rect 10292 8128 10293 8168
rect 10251 8119 10293 8128
rect 11835 8168 11877 8177
rect 11835 8128 11836 8168
rect 11876 8128 11877 8168
rect 11835 8119 11877 8128
rect 16443 8168 16485 8177
rect 16443 8128 16444 8168
rect 16484 8128 16485 8168
rect 16443 8119 16485 8128
rect 25899 8168 25941 8177
rect 25899 8128 25900 8168
rect 25940 8128 25941 8168
rect 25899 8119 25941 8128
rect 30651 8168 30693 8177
rect 30651 8128 30652 8168
rect 30692 8128 30693 8168
rect 30651 8119 30693 8128
rect 32811 8168 32853 8177
rect 32811 8128 32812 8168
rect 32852 8128 32853 8168
rect 32811 8119 32853 8128
rect 39387 8168 39429 8177
rect 39387 8128 39388 8168
rect 39428 8128 39429 8168
rect 39387 8119 39429 8128
rect 44379 8168 44421 8177
rect 44379 8128 44380 8168
rect 44420 8128 44421 8168
rect 44379 8119 44421 8128
rect 12219 8084 12261 8093
rect 12219 8044 12220 8084
rect 12260 8044 12261 8084
rect 12219 8035 12261 8044
rect 20043 8084 20085 8093
rect 20043 8044 20044 8084
rect 20084 8044 20085 8084
rect 20043 8035 20085 8044
rect 22827 8084 22869 8093
rect 22827 8044 22828 8084
rect 22868 8044 22869 8084
rect 22827 8035 22869 8044
rect 30555 8084 30597 8093
rect 30555 8044 30556 8084
rect 30596 8044 30597 8084
rect 30555 8035 30597 8044
rect 36507 8084 36549 8093
rect 36507 8044 36508 8084
rect 36548 8044 36549 8084
rect 36507 8035 36549 8044
rect 1227 8000 1269 8009
rect 1227 7960 1228 8000
rect 1268 7960 1269 8000
rect 1227 7951 1269 7960
rect 1611 8000 1653 8009
rect 1611 7960 1612 8000
rect 1652 7960 1653 8000
rect 1611 7951 1653 7960
rect 4107 8000 4149 8009
rect 4107 7960 4108 8000
rect 4148 7960 4149 8000
rect 4107 7951 4149 7960
rect 9483 8000 9525 8009
rect 9483 7960 9484 8000
rect 9524 7960 9525 8000
rect 9483 7951 9525 7960
rect 9723 8000 9765 8009
rect 9723 7960 9724 8000
rect 9764 7960 9765 8000
rect 9723 7951 9765 7960
rect 9867 8000 9909 8009
rect 9867 7960 9868 8000
rect 9908 7960 9909 8000
rect 9867 7951 9909 7960
rect 11211 8000 11253 8009
rect 11211 7960 11212 8000
rect 11252 7960 11253 8000
rect 11211 7951 11253 7960
rect 11595 8000 11637 8009
rect 11595 7960 11596 8000
rect 11636 7960 11637 8000
rect 11595 7951 11637 7960
rect 11979 8000 12021 8009
rect 11979 7960 11980 8000
rect 12020 7960 12021 8000
rect 11979 7951 12021 7960
rect 12346 8000 12404 8001
rect 12346 7960 12355 8000
rect 12395 7960 12404 8000
rect 12346 7959 12404 7960
rect 16203 8000 16245 8009
rect 16203 7960 16204 8000
rect 16244 7960 16245 8000
rect 16203 7951 16245 7960
rect 16587 8000 16629 8009
rect 16587 7960 16588 8000
rect 16628 7960 16629 8000
rect 16587 7951 16629 7960
rect 16971 8000 17013 8009
rect 16971 7960 16972 8000
rect 17012 7960 17013 8000
rect 16971 7951 17013 7960
rect 17211 8000 17253 8009
rect 17211 7960 17212 8000
rect 17252 7960 17253 8000
rect 17211 7951 17253 7960
rect 20715 8000 20757 8009
rect 20715 7960 20716 8000
rect 20756 7960 20757 8000
rect 20715 7951 20757 7960
rect 21099 8000 21141 8009
rect 21099 7960 21100 8000
rect 21140 7960 21141 8000
rect 21099 7951 21141 7960
rect 21483 8000 21525 8009
rect 21483 7960 21484 8000
rect 21524 7960 21525 8000
rect 21483 7951 21525 7960
rect 21675 8000 21717 8009
rect 21675 7960 21676 8000
rect 21716 7960 21717 8000
rect 21675 7951 21717 7960
rect 22971 8000 23013 8009
rect 22971 7960 22972 8000
rect 23012 7960 23013 8000
rect 22971 7951 23013 7960
rect 23211 8000 23253 8009
rect 23211 7960 23212 8000
rect 23252 7960 23253 8000
rect 23211 7951 23253 7960
rect 23355 8000 23397 8009
rect 23355 7960 23356 8000
rect 23396 7960 23397 8000
rect 23355 7951 23397 7960
rect 23595 8000 23637 8009
rect 23595 7960 23596 8000
rect 23636 7960 23637 8000
rect 23595 7951 23637 7960
rect 28491 8000 28533 8009
rect 28491 7960 28492 8000
rect 28532 7960 28533 8000
rect 28491 7951 28533 7960
rect 30123 8000 30165 8009
rect 30123 7960 30124 8000
rect 30164 7960 30165 8000
rect 30123 7951 30165 7960
rect 30315 8000 30357 8009
rect 30315 7960 30316 8000
rect 30356 7960 30357 8000
rect 30315 7951 30357 7960
rect 30891 8000 30933 8009
rect 30891 7960 30892 8000
rect 30932 7960 30933 8000
rect 30891 7951 30933 7960
rect 34635 8000 34677 8009
rect 34635 7960 34636 8000
rect 34676 7960 34677 8000
rect 34635 7951 34677 7960
rect 36123 8000 36165 8009
rect 36123 7960 36124 8000
rect 36164 7960 36165 8000
rect 36123 7951 36165 7960
rect 36363 8000 36405 8009
rect 36363 7960 36364 8000
rect 36404 7960 36405 8000
rect 36363 7951 36405 7960
rect 36747 8000 36789 8009
rect 36747 7960 36748 8000
rect 36788 7960 36789 8000
rect 36747 7951 36789 7960
rect 37131 8000 37173 8009
rect 37131 7960 37132 8000
rect 37172 7960 37173 8000
rect 37131 7951 37173 7960
rect 39627 8000 39669 8009
rect 39627 7960 39628 8000
rect 39668 7960 39669 8000
rect 39627 7951 39669 7960
rect 41451 8000 41493 8009
rect 41451 7960 41452 8000
rect 41492 7960 41493 8000
rect 41451 7951 41493 7960
rect 42123 8000 42165 8009
rect 42123 7960 42124 8000
rect 42164 7960 42165 8000
rect 42123 7951 42165 7960
rect 44139 8000 44181 8009
rect 44139 7960 44140 8000
rect 44180 7960 44181 8000
rect 44139 7951 44181 7960
rect 44523 8000 44565 8009
rect 44523 7960 44524 8000
rect 44564 7960 44565 8000
rect 44523 7951 44565 7960
rect 44907 8000 44949 8009
rect 44907 7960 44908 8000
rect 44948 7960 44949 8000
rect 44907 7951 44949 7960
rect 4491 7916 4533 7925
rect 4491 7876 4492 7916
rect 4532 7876 4533 7916
rect 4491 7867 4533 7876
rect 5731 7916 5789 7917
rect 5731 7876 5740 7916
rect 5780 7876 5789 7916
rect 5731 7875 5789 7876
rect 7563 7916 7605 7925
rect 7563 7876 7564 7916
rect 7604 7876 7605 7916
rect 7563 7867 7605 7876
rect 8803 7916 8861 7917
rect 10923 7916 10965 7925
rect 8803 7876 8812 7916
rect 8852 7876 8861 7916
rect 8803 7875 8861 7876
rect 10635 7907 10677 7916
rect 10635 7867 10636 7907
rect 10676 7867 10677 7907
rect 10923 7876 10924 7916
rect 10964 7876 10965 7916
rect 10923 7867 10965 7876
rect 12547 7916 12605 7917
rect 12547 7876 12556 7916
rect 12596 7876 12605 7916
rect 12547 7875 12605 7876
rect 13803 7916 13845 7925
rect 13803 7876 13804 7916
rect 13844 7876 13845 7916
rect 13803 7867 13845 7876
rect 14283 7916 14325 7925
rect 14283 7876 14284 7916
rect 14324 7876 14325 7916
rect 14283 7867 14325 7876
rect 15523 7916 15581 7917
rect 15523 7876 15532 7916
rect 15572 7876 15581 7916
rect 15523 7875 15581 7876
rect 17355 7916 17397 7925
rect 17355 7876 17356 7916
rect 17396 7876 17397 7916
rect 17355 7867 17397 7876
rect 18595 7916 18653 7917
rect 18595 7876 18604 7916
rect 18644 7876 18653 7916
rect 18595 7875 18653 7876
rect 19371 7916 19413 7925
rect 19371 7876 19372 7916
rect 19412 7876 19413 7916
rect 19371 7867 19413 7876
rect 19642 7916 19700 7917
rect 19642 7876 19651 7916
rect 19691 7876 19700 7916
rect 19642 7875 19700 7876
rect 22155 7916 22197 7925
rect 22155 7876 22156 7916
rect 22196 7876 22197 7916
rect 22155 7867 22197 7876
rect 22426 7916 22484 7917
rect 22426 7876 22435 7916
rect 22475 7876 22484 7916
rect 22426 7875 22484 7876
rect 24459 7916 24501 7925
rect 24459 7876 24460 7916
rect 24500 7876 24501 7916
rect 24459 7867 24501 7876
rect 25699 7916 25757 7917
rect 25699 7876 25708 7916
rect 25748 7876 25757 7916
rect 25699 7875 25757 7876
rect 26283 7916 26325 7925
rect 26283 7876 26284 7916
rect 26324 7876 26325 7916
rect 26283 7867 26325 7876
rect 27523 7916 27581 7917
rect 27523 7876 27532 7916
rect 27572 7876 27581 7916
rect 27523 7875 27581 7876
rect 27994 7916 28052 7917
rect 27994 7876 28003 7916
rect 28043 7876 28052 7916
rect 27994 7875 28052 7876
rect 28107 7916 28149 7925
rect 28107 7876 28108 7916
rect 28148 7876 28149 7916
rect 28107 7867 28149 7876
rect 28587 7916 28629 7925
rect 28587 7876 28588 7916
rect 28628 7876 28629 7916
rect 28587 7867 28629 7876
rect 29059 7916 29117 7917
rect 29059 7876 29068 7916
rect 29108 7876 29117 7916
rect 29059 7875 29117 7876
rect 29547 7916 29605 7917
rect 29547 7876 29556 7916
rect 29596 7876 29605 7916
rect 29547 7875 29605 7876
rect 31371 7916 31413 7925
rect 31371 7876 31372 7916
rect 31412 7876 31413 7916
rect 31371 7867 31413 7876
rect 32611 7916 32669 7917
rect 32611 7876 32620 7916
rect 32660 7876 32669 7916
rect 32611 7875 32669 7876
rect 33003 7916 33045 7925
rect 33003 7876 33004 7916
rect 33044 7876 33045 7916
rect 33003 7867 33045 7876
rect 34243 7916 34301 7917
rect 34243 7876 34252 7916
rect 34292 7876 34301 7916
rect 34243 7875 34301 7876
rect 35307 7916 35349 7925
rect 35307 7876 35308 7916
rect 35348 7876 35349 7916
rect 35307 7867 35349 7876
rect 35578 7916 35636 7917
rect 35578 7876 35587 7916
rect 35627 7876 35636 7916
rect 35578 7875 35636 7876
rect 36027 7916 36069 7925
rect 36027 7876 36028 7916
rect 36068 7876 36069 7916
rect 36027 7867 36069 7876
rect 37515 7916 37557 7925
rect 37515 7876 37516 7916
rect 37556 7876 37557 7916
rect 37515 7867 37557 7876
rect 38755 7916 38813 7917
rect 38755 7876 38764 7916
rect 38804 7876 38813 7916
rect 38755 7875 38813 7876
rect 10635 7858 10677 7867
rect 10539 7832 10581 7841
rect 10539 7792 10540 7832
rect 10580 7792 10581 7832
rect 10539 7783 10581 7792
rect 16827 7832 16869 7841
rect 16827 7792 16828 7832
rect 16868 7792 16869 7832
rect 16827 7783 16869 7792
rect 18795 7832 18837 7841
rect 18795 7792 18796 7832
rect 18836 7792 18837 7832
rect 18795 7783 18837 7792
rect 19739 7832 19781 7841
rect 19739 7792 19740 7832
rect 19780 7792 19781 7832
rect 19739 7783 19781 7792
rect 21243 7832 21285 7841
rect 21243 7792 21244 7832
rect 21284 7792 21285 7832
rect 21243 7783 21285 7792
rect 22539 7832 22581 7841
rect 22539 7792 22540 7832
rect 22580 7792 22581 7832
rect 22539 7783 22581 7792
rect 27723 7832 27765 7841
rect 27723 7792 27724 7832
rect 27764 7792 27765 7832
rect 27723 7783 27765 7792
rect 34875 7832 34917 7841
rect 34875 7792 34876 7832
rect 34916 7792 34917 7832
rect 34875 7783 34917 7792
rect 35691 7832 35733 7841
rect 35691 7792 35692 7832
rect 35732 7792 35733 7832
rect 35691 7783 35733 7792
rect 36891 7832 36933 7841
rect 36891 7792 36892 7832
rect 36932 7792 36933 7832
rect 36891 7783 36933 7792
rect 41835 7832 41877 7841
rect 41835 7792 41836 7832
rect 41876 7792 41877 7832
rect 41835 7783 41877 7792
rect 42411 7832 42453 7841
rect 42411 7792 42412 7832
rect 42452 7792 42453 7832
rect 42411 7783 42453 7792
rect 42699 7832 42741 7841
rect 42699 7792 42700 7832
rect 42740 7792 42741 7832
rect 42699 7783 42741 7792
rect 42987 7832 43029 7841
rect 42987 7792 42988 7832
rect 43028 7792 43029 7832
rect 42987 7783 43029 7792
rect 43275 7832 43317 7841
rect 43275 7792 43276 7832
rect 43316 7792 43317 7832
rect 43275 7783 43317 7792
rect 1467 7748 1509 7757
rect 1467 7708 1468 7748
rect 1508 7708 1509 7748
rect 1467 7699 1509 7708
rect 1851 7748 1893 7757
rect 1851 7708 1852 7748
rect 1892 7708 1893 7748
rect 1851 7699 1893 7708
rect 5931 7748 5973 7757
rect 5931 7708 5932 7748
rect 5972 7708 5973 7748
rect 5931 7699 5973 7708
rect 9003 7748 9045 7757
rect 9003 7708 9004 7748
rect 9044 7708 9045 7748
rect 9003 7699 9045 7708
rect 10107 7748 10149 7757
rect 10107 7708 10108 7748
rect 10148 7708 10149 7748
rect 10107 7699 10149 7708
rect 11451 7748 11493 7757
rect 11451 7708 11452 7748
rect 11492 7708 11493 7748
rect 11451 7699 11493 7708
rect 15723 7748 15765 7757
rect 15723 7708 15724 7748
rect 15764 7708 15765 7748
rect 15723 7699 15765 7708
rect 20475 7748 20517 7757
rect 20475 7708 20476 7748
rect 20516 7708 20517 7748
rect 20475 7699 20517 7708
rect 20859 7748 20901 7757
rect 20859 7708 20860 7748
rect 20900 7708 20901 7748
rect 20859 7699 20901 7708
rect 21915 7748 21957 7757
rect 21915 7708 21916 7748
rect 21956 7708 21957 7748
rect 21915 7699 21957 7708
rect 29739 7748 29781 7757
rect 29739 7708 29740 7748
rect 29780 7708 29781 7748
rect 29739 7699 29781 7708
rect 29883 7748 29925 7757
rect 29883 7708 29884 7748
rect 29924 7708 29925 7748
rect 29883 7699 29925 7708
rect 34443 7748 34485 7757
rect 34443 7708 34444 7748
rect 34484 7708 34485 7748
rect 34443 7699 34485 7708
rect 38955 7748 38997 7757
rect 38955 7708 38956 7748
rect 38996 7708 38997 7748
rect 38955 7699 38997 7708
rect 40954 7748 41012 7749
rect 40954 7708 40963 7748
rect 41003 7708 41012 7748
rect 40954 7707 41012 7708
rect 41211 7748 41253 7757
rect 41211 7708 41212 7748
rect 41252 7708 41253 7748
rect 41211 7699 41253 7708
rect 42202 7748 42260 7749
rect 42202 7708 42211 7748
rect 42251 7708 42260 7748
rect 42202 7707 42260 7708
rect 43642 7748 43700 7749
rect 43642 7708 43651 7748
rect 43691 7708 43700 7748
rect 43642 7707 43700 7708
rect 43834 7748 43892 7749
rect 43834 7708 43843 7748
rect 43883 7708 43892 7748
rect 43834 7707 43892 7708
rect 44763 7748 44805 7757
rect 44763 7708 44764 7748
rect 44804 7708 44805 7748
rect 44763 7699 44805 7708
rect 45147 7748 45189 7757
rect 45147 7708 45148 7748
rect 45188 7708 45189 7748
rect 45147 7699 45189 7708
rect 1152 7580 45216 7604
rect 1152 7540 4928 7580
rect 4968 7540 5010 7580
rect 5050 7540 5092 7580
rect 5132 7540 5174 7580
rect 5214 7540 5256 7580
rect 5296 7540 20048 7580
rect 20088 7540 20130 7580
rect 20170 7540 20212 7580
rect 20252 7540 20294 7580
rect 20334 7540 20376 7580
rect 20416 7540 35168 7580
rect 35208 7540 35250 7580
rect 35290 7540 35332 7580
rect 35372 7540 35414 7580
rect 35454 7540 35496 7580
rect 35536 7540 45216 7580
rect 1152 7516 45216 7540
rect 10107 7412 10149 7421
rect 10107 7372 10108 7412
rect 10148 7372 10149 7412
rect 10107 7363 10149 7372
rect 29355 7412 29397 7421
rect 29355 7372 29356 7412
rect 29396 7372 29397 7412
rect 29355 7363 29397 7372
rect 33339 7412 33381 7421
rect 33339 7372 33340 7412
rect 33380 7372 33381 7412
rect 33339 7363 33381 7372
rect 33723 7412 33765 7421
rect 33723 7372 33724 7412
rect 33764 7372 33765 7412
rect 33723 7363 33765 7372
rect 41818 7412 41876 7413
rect 41818 7372 41827 7412
rect 41867 7372 41876 7412
rect 41818 7371 41876 7372
rect 42490 7412 42548 7413
rect 42490 7372 42499 7412
rect 42539 7372 42548 7412
rect 42490 7371 42548 7372
rect 42778 7412 42836 7413
rect 42778 7372 42787 7412
rect 42827 7372 42836 7412
rect 42778 7371 42836 7372
rect 9771 7328 9813 7337
rect 9771 7288 9772 7328
rect 9812 7288 9813 7328
rect 9771 7279 9813 7288
rect 11019 7328 11061 7337
rect 11019 7288 11020 7328
rect 11060 7288 11061 7328
rect 11019 7279 11061 7288
rect 21675 7328 21717 7337
rect 21675 7288 21676 7328
rect 21716 7288 21717 7328
rect 21675 7279 21717 7288
rect 32955 7328 32997 7337
rect 32955 7288 32956 7328
rect 32996 7288 32997 7328
rect 32955 7279 32997 7288
rect 9387 7244 9429 7253
rect 9387 7204 9388 7244
rect 9428 7204 9429 7244
rect 9387 7195 9429 7204
rect 9658 7244 9716 7245
rect 9658 7204 9667 7244
rect 9707 7204 9716 7244
rect 9658 7203 9716 7204
rect 10635 7244 10677 7253
rect 10635 7204 10636 7244
rect 10676 7204 10677 7244
rect 10635 7195 10677 7204
rect 10906 7244 10964 7245
rect 10906 7204 10915 7244
rect 10955 7204 10964 7244
rect 10906 7203 10964 7204
rect 17067 7244 17109 7253
rect 21291 7244 21333 7253
rect 17067 7204 17068 7244
rect 17108 7204 17109 7244
rect 17067 7195 17109 7204
rect 18315 7235 18357 7244
rect 18315 7195 18316 7235
rect 18356 7195 18357 7235
rect 21291 7204 21292 7244
rect 21332 7204 21333 7244
rect 21291 7195 21333 7204
rect 21562 7244 21620 7245
rect 21562 7204 21571 7244
rect 21611 7204 21620 7244
rect 21562 7203 21620 7204
rect 23019 7244 23061 7253
rect 23019 7204 23020 7244
rect 23060 7204 23061 7244
rect 23019 7195 23061 7204
rect 23266 7244 23324 7245
rect 23266 7204 23275 7244
rect 23315 7204 23324 7244
rect 23266 7203 23324 7204
rect 23386 7244 23444 7245
rect 23386 7204 23395 7244
rect 23435 7204 23444 7244
rect 23386 7203 23444 7204
rect 27915 7244 27957 7253
rect 30699 7244 30741 7253
rect 34426 7244 34484 7245
rect 27915 7204 27916 7244
rect 27956 7204 27957 7244
rect 27915 7195 27957 7204
rect 29163 7235 29205 7244
rect 29163 7195 29164 7235
rect 29204 7195 29205 7235
rect 30699 7204 30700 7244
rect 30740 7204 30741 7244
rect 30699 7195 30741 7204
rect 31947 7235 31989 7244
rect 31947 7195 31948 7235
rect 31988 7195 31989 7235
rect 34426 7204 34435 7244
rect 34475 7204 34484 7244
rect 34426 7203 34484 7204
rect 34539 7244 34581 7253
rect 34539 7204 34540 7244
rect 34580 7204 34581 7244
rect 34539 7195 34581 7204
rect 34923 7244 34965 7253
rect 39435 7244 39477 7253
rect 34923 7204 34924 7244
rect 34964 7204 34965 7244
rect 34923 7195 34965 7204
rect 35499 7235 35541 7244
rect 35499 7195 35500 7235
rect 35540 7195 35541 7235
rect 18315 7186 18357 7195
rect 29163 7186 29205 7195
rect 31947 7186 31989 7195
rect 35499 7186 35541 7195
rect 35979 7235 36021 7244
rect 35979 7195 35980 7235
rect 36020 7195 36021 7235
rect 39435 7204 39436 7244
rect 39476 7204 39477 7244
rect 39435 7195 39477 7204
rect 40683 7235 40725 7244
rect 40683 7195 40684 7235
rect 40724 7195 40725 7235
rect 35979 7186 36021 7195
rect 40683 7186 40725 7195
rect 1227 7160 1269 7169
rect 1227 7120 1228 7160
rect 1268 7120 1269 7160
rect 1227 7111 1269 7120
rect 1611 7160 1653 7169
rect 1611 7120 1612 7160
rect 1652 7120 1653 7160
rect 1611 7111 1653 7120
rect 1851 7160 1893 7169
rect 1851 7120 1852 7160
rect 1892 7120 1893 7160
rect 1851 7111 1893 7120
rect 3531 7160 3573 7169
rect 3531 7120 3532 7160
rect 3572 7120 3573 7160
rect 3531 7111 3573 7120
rect 6315 7160 6357 7169
rect 6315 7120 6316 7160
rect 6356 7120 6357 7160
rect 6315 7111 6357 7120
rect 6555 7160 6597 7169
rect 6555 7120 6556 7160
rect 6596 7120 6597 7160
rect 6555 7111 6597 7120
rect 8139 7160 8181 7169
rect 8139 7120 8140 7160
rect 8180 7120 8181 7160
rect 8139 7111 8181 7120
rect 8523 7160 8565 7169
rect 8523 7120 8524 7160
rect 8564 7120 8565 7160
rect 8523 7111 8565 7120
rect 8907 7160 8949 7169
rect 8907 7120 8908 7160
rect 8948 7120 8949 7160
rect 8907 7111 8949 7120
rect 9147 7160 9189 7169
rect 9147 7120 9148 7160
rect 9188 7120 9189 7160
rect 9147 7111 9189 7120
rect 11691 7160 11733 7169
rect 11691 7120 11692 7160
rect 11732 7120 11733 7160
rect 11691 7111 11733 7120
rect 12075 7160 12117 7169
rect 12075 7120 12076 7160
rect 12116 7120 12117 7160
rect 12075 7111 12117 7120
rect 12459 7160 12501 7169
rect 12459 7120 12460 7160
rect 12500 7120 12501 7160
rect 12459 7111 12501 7120
rect 12843 7160 12885 7169
rect 12843 7120 12844 7160
rect 12884 7120 12885 7160
rect 12843 7111 12885 7120
rect 13227 7160 13269 7169
rect 13227 7120 13228 7160
rect 13268 7120 13269 7160
rect 13227 7111 13269 7120
rect 13467 7160 13509 7169
rect 13467 7120 13468 7160
rect 13508 7120 13509 7160
rect 13467 7111 13509 7120
rect 13611 7160 13653 7169
rect 13611 7120 13612 7160
rect 13652 7120 13653 7160
rect 13611 7111 13653 7120
rect 13995 7160 14037 7169
rect 13995 7120 13996 7160
rect 14036 7120 14037 7160
rect 13995 7111 14037 7120
rect 14379 7160 14421 7169
rect 14379 7120 14380 7160
rect 14420 7120 14421 7160
rect 14379 7111 14421 7120
rect 14763 7160 14805 7169
rect 14763 7120 14764 7160
rect 14804 7120 14805 7160
rect 14763 7111 14805 7120
rect 15003 7160 15045 7169
rect 15003 7120 15004 7160
rect 15044 7120 15045 7160
rect 15003 7111 15045 7120
rect 15147 7160 15189 7169
rect 15147 7120 15148 7160
rect 15188 7120 15189 7160
rect 15147 7111 15189 7120
rect 15531 7160 15573 7169
rect 15531 7120 15532 7160
rect 15572 7120 15573 7160
rect 15531 7111 15573 7120
rect 15915 7160 15957 7169
rect 15915 7120 15916 7160
rect 15956 7120 15957 7160
rect 15915 7111 15957 7120
rect 16299 7160 16341 7169
rect 16299 7120 16300 7160
rect 16340 7120 16341 7160
rect 16299 7111 16341 7120
rect 16683 7160 16725 7169
rect 16683 7120 16684 7160
rect 16724 7120 16725 7160
rect 16683 7111 16725 7120
rect 18891 7160 18933 7169
rect 18891 7120 18892 7160
rect 18932 7120 18933 7160
rect 18891 7111 18933 7120
rect 19275 7160 19317 7169
rect 19275 7120 19276 7160
rect 19316 7120 19317 7160
rect 19275 7111 19317 7120
rect 19659 7160 19701 7169
rect 19659 7120 19660 7160
rect 19700 7120 19701 7160
rect 19659 7111 19701 7120
rect 19899 7160 19941 7169
rect 19899 7120 19900 7160
rect 19940 7120 19941 7160
rect 19899 7111 19941 7120
rect 20235 7160 20277 7169
rect 20235 7120 20236 7160
rect 20276 7120 20277 7160
rect 20235 7111 20277 7120
rect 20619 7160 20661 7169
rect 20619 7120 20620 7160
rect 20660 7120 20661 7160
rect 20619 7111 20661 7120
rect 20763 7160 20805 7169
rect 20763 7120 20764 7160
rect 20804 7120 20805 7160
rect 20763 7111 20805 7120
rect 21003 7160 21045 7169
rect 21003 7120 21004 7160
rect 21044 7120 21045 7160
rect 21003 7111 21045 7120
rect 22347 7160 22389 7169
rect 22347 7120 22348 7160
rect 22388 7120 22389 7160
rect 22347 7111 22389 7120
rect 22539 7160 22581 7169
rect 22539 7120 22540 7160
rect 22580 7120 22581 7160
rect 22539 7111 22581 7120
rect 23979 7160 24021 7169
rect 23979 7120 23980 7160
rect 24020 7120 24021 7160
rect 23979 7111 24021 7120
rect 25131 7160 25173 7169
rect 25131 7120 25132 7160
rect 25172 7120 25173 7160
rect 25131 7111 25173 7120
rect 25707 7160 25749 7169
rect 25707 7120 25708 7160
rect 25748 7120 25749 7160
rect 25707 7111 25749 7120
rect 26091 7160 26133 7169
rect 26091 7120 26092 7160
rect 26132 7120 26133 7160
rect 26091 7111 26133 7120
rect 27051 7160 27093 7169
rect 27051 7120 27052 7160
rect 27092 7120 27093 7160
rect 27051 7111 27093 7120
rect 27723 7160 27765 7169
rect 27723 7120 27724 7160
rect 27764 7120 27765 7160
rect 27723 7111 27765 7120
rect 29499 7160 29541 7169
rect 29499 7120 29500 7160
rect 29540 7120 29541 7160
rect 29499 7111 29541 7120
rect 30123 7160 30165 7169
rect 30123 7120 30124 7160
rect 30164 7120 30165 7160
rect 30123 7111 30165 7120
rect 30315 7160 30357 7169
rect 30315 7120 30316 7160
rect 30356 7120 30357 7160
rect 30315 7111 30357 7120
rect 32523 7160 32565 7169
rect 32523 7120 32524 7160
rect 32564 7120 32565 7160
rect 32523 7111 32565 7120
rect 32715 7160 32757 7169
rect 32715 7120 32716 7160
rect 32756 7120 32757 7160
rect 32715 7111 32757 7120
rect 33099 7160 33141 7169
rect 33099 7120 33100 7160
rect 33140 7120 33141 7160
rect 33099 7111 33141 7120
rect 33483 7160 33525 7169
rect 33483 7120 33484 7160
rect 33524 7120 33525 7160
rect 33483 7111 33525 7120
rect 34059 7160 34101 7169
rect 34059 7120 34060 7160
rect 34100 7120 34101 7160
rect 34059 7111 34101 7120
rect 35019 7160 35061 7169
rect 35019 7120 35020 7160
rect 35060 7120 35061 7160
rect 35019 7111 35061 7120
rect 36555 7160 36597 7169
rect 36555 7120 36556 7160
rect 36596 7120 36597 7160
rect 36555 7111 36597 7120
rect 36939 7160 36981 7169
rect 36939 7120 36940 7160
rect 36980 7120 36981 7160
rect 36939 7111 36981 7120
rect 37323 7160 37365 7169
rect 37323 7120 37324 7160
rect 37364 7120 37365 7160
rect 37323 7111 37365 7120
rect 37707 7160 37749 7169
rect 37707 7120 37708 7160
rect 37748 7120 37749 7160
rect 37707 7111 37749 7120
rect 42219 7160 42261 7169
rect 42219 7120 42220 7160
rect 42260 7120 42261 7160
rect 42219 7111 42261 7120
rect 43179 7160 43221 7169
rect 43179 7120 43180 7160
rect 43220 7120 43221 7160
rect 43179 7111 43221 7120
rect 43467 7160 43509 7169
rect 43467 7120 43468 7160
rect 43508 7120 43509 7160
rect 43467 7111 43509 7120
rect 43755 7160 43797 7169
rect 43755 7120 43756 7160
rect 43796 7120 43797 7160
rect 43755 7111 43797 7120
rect 44043 7160 44085 7169
rect 44043 7120 44044 7160
rect 44084 7120 44085 7160
rect 44043 7111 44085 7120
rect 44331 7160 44373 7169
rect 44331 7120 44332 7160
rect 44372 7120 44373 7160
rect 44331 7111 44373 7120
rect 44523 7160 44565 7169
rect 44523 7120 44524 7160
rect 44564 7120 44565 7160
rect 44523 7111 44565 7120
rect 44907 7160 44949 7169
rect 44907 7120 44908 7160
rect 44948 7120 44949 7160
rect 44907 7111 44949 7120
rect 12315 7076 12357 7085
rect 12315 7036 12316 7076
rect 12356 7036 12357 7076
rect 12315 7027 12357 7036
rect 14235 7076 14277 7085
rect 14235 7036 14236 7076
rect 14276 7036 14277 7076
rect 14235 7027 14277 7036
rect 15771 7076 15813 7085
rect 15771 7036 15772 7076
rect 15812 7036 15813 7076
rect 15771 7027 15813 7036
rect 16539 7076 16581 7085
rect 16539 7036 16540 7076
rect 16580 7036 16581 7076
rect 16539 7027 16581 7036
rect 19515 7076 19557 7085
rect 19515 7036 19516 7076
rect 19556 7036 19557 7076
rect 19515 7027 19557 7036
rect 21963 7076 22005 7085
rect 21963 7036 21964 7076
rect 22004 7036 22005 7076
rect 21963 7027 22005 7036
rect 27483 7076 27525 7085
rect 27483 7036 27484 7076
rect 27524 7036 27525 7076
rect 27483 7027 27525 7036
rect 29787 7076 29829 7085
rect 29787 7036 29788 7076
rect 29828 7036 29829 7076
rect 29787 7027 29829 7036
rect 32139 7076 32181 7085
rect 32139 7036 32140 7076
rect 32180 7036 32181 7076
rect 32139 7027 32181 7036
rect 44763 7076 44805 7085
rect 44763 7036 44764 7076
rect 44804 7036 44805 7076
rect 44763 7027 44805 7036
rect 1467 6992 1509 7001
rect 1467 6952 1468 6992
rect 1508 6952 1509 6992
rect 1467 6943 1509 6952
rect 3771 6992 3813 7001
rect 3771 6952 3772 6992
rect 3812 6952 3813 6992
rect 3771 6943 3813 6952
rect 8379 6992 8421 7001
rect 8379 6952 8380 6992
rect 8420 6952 8421 6992
rect 8379 6943 8421 6952
rect 8763 6992 8805 7001
rect 8763 6952 8764 6992
rect 8804 6952 8805 6992
rect 8763 6943 8805 6952
rect 11307 6992 11349 7001
rect 11307 6952 11308 6992
rect 11348 6952 11349 6992
rect 11307 6943 11349 6952
rect 11931 6992 11973 7001
rect 11931 6952 11932 6992
rect 11972 6952 11973 6992
rect 11931 6943 11973 6952
rect 12699 6992 12741 7001
rect 12699 6952 12700 6992
rect 12740 6952 12741 6992
rect 12699 6943 12741 6952
rect 13083 6992 13125 7001
rect 13083 6952 13084 6992
rect 13124 6952 13125 6992
rect 13083 6943 13125 6952
rect 13851 6992 13893 7001
rect 13851 6952 13852 6992
rect 13892 6952 13893 6992
rect 13851 6943 13893 6952
rect 14619 6992 14661 7001
rect 14619 6952 14620 6992
rect 14660 6952 14661 6992
rect 14619 6943 14661 6952
rect 15387 6992 15429 7001
rect 15387 6952 15388 6992
rect 15428 6952 15429 6992
rect 15387 6943 15429 6952
rect 16155 6992 16197 7001
rect 16155 6952 16156 6992
rect 16196 6952 16197 6992
rect 16155 6943 16197 6952
rect 16923 6992 16965 7001
rect 16923 6952 16924 6992
rect 16964 6952 16965 6992
rect 16923 6943 16965 6952
rect 18507 6992 18549 7001
rect 18507 6952 18508 6992
rect 18548 6952 18549 6992
rect 18507 6943 18549 6952
rect 19131 6992 19173 7001
rect 19131 6952 19132 6992
rect 19172 6952 19173 6992
rect 19131 6943 19173 6952
rect 19995 6992 20037 7001
rect 19995 6952 19996 6992
rect 20036 6952 20037 6992
rect 19995 6943 20037 6952
rect 20379 6992 20421 7001
rect 20379 6952 20380 6992
rect 20420 6952 20421 6992
rect 20379 6943 20421 6952
rect 22107 6992 22149 7001
rect 22107 6952 22108 6992
rect 22148 6952 22149 6992
rect 22107 6943 22149 6952
rect 22779 6992 22821 7001
rect 22779 6952 22780 6992
rect 22820 6952 22821 6992
rect 22779 6943 22821 6952
rect 23691 6992 23733 7001
rect 23691 6952 23692 6992
rect 23732 6952 23733 6992
rect 23691 6943 23733 6952
rect 24219 6992 24261 7001
rect 24219 6952 24220 6992
rect 24260 6952 24261 6992
rect 24219 6943 24261 6952
rect 25371 6992 25413 7001
rect 25371 6952 25372 6992
rect 25412 6952 25413 6992
rect 25371 6943 25413 6952
rect 25947 6992 25989 7001
rect 25947 6952 25948 6992
rect 25988 6952 25989 6992
rect 25947 6943 25989 6952
rect 26331 6992 26373 7001
rect 26331 6952 26332 6992
rect 26372 6952 26373 6992
rect 26331 6943 26373 6952
rect 27291 6992 27333 7001
rect 27291 6952 27292 6992
rect 27332 6952 27333 6992
rect 27291 6943 27333 6952
rect 29883 6992 29925 7001
rect 29883 6952 29884 6992
rect 29924 6952 29925 6992
rect 29883 6943 29925 6952
rect 30555 6992 30597 7001
rect 30555 6952 30556 6992
rect 30596 6952 30597 6992
rect 30555 6943 30597 6952
rect 32283 6992 32325 7001
rect 32283 6952 32284 6992
rect 32324 6952 32325 6992
rect 32283 6943 32325 6952
rect 33819 6992 33861 7001
rect 33819 6952 33820 6992
rect 33860 6952 33861 6992
rect 33819 6943 33861 6952
rect 36202 6992 36260 6993
rect 36202 6952 36211 6992
rect 36251 6952 36260 6992
rect 36202 6951 36260 6952
rect 36315 6992 36357 7001
rect 36315 6952 36316 6992
rect 36356 6952 36357 6992
rect 36315 6943 36357 6952
rect 36699 6992 36741 7001
rect 36699 6952 36700 6992
rect 36740 6952 36741 6992
rect 36699 6943 36741 6952
rect 37083 6992 37125 7001
rect 37083 6952 37084 6992
rect 37124 6952 37125 6992
rect 37083 6943 37125 6952
rect 37467 6992 37509 7001
rect 37467 6952 37468 6992
rect 37508 6952 37509 6992
rect 37467 6943 37509 6952
rect 40875 6992 40917 7001
rect 40875 6952 40876 6992
rect 40916 6952 40917 6992
rect 40875 6943 40917 6952
rect 41979 6992 42021 7001
rect 41979 6952 41980 6992
rect 42020 6952 42021 6992
rect 41979 6943 42021 6952
rect 45147 6992 45189 7001
rect 45147 6952 45148 6992
rect 45188 6952 45189 6992
rect 45147 6943 45189 6952
rect 1152 6824 45216 6848
rect 1152 6784 3688 6824
rect 3728 6784 3770 6824
rect 3810 6784 3852 6824
rect 3892 6784 3934 6824
rect 3974 6784 4016 6824
rect 4056 6784 18808 6824
rect 18848 6784 18890 6824
rect 18930 6784 18972 6824
rect 19012 6784 19054 6824
rect 19094 6784 19136 6824
rect 19176 6784 33928 6824
rect 33968 6784 34010 6824
rect 34050 6784 34092 6824
rect 34132 6784 34174 6824
rect 34214 6784 34256 6824
rect 34296 6784 45216 6824
rect 1152 6760 45216 6784
rect 10107 6656 10149 6665
rect 10107 6616 10108 6656
rect 10148 6616 10149 6656
rect 10107 6607 10149 6616
rect 12507 6656 12549 6665
rect 12507 6616 12508 6656
rect 12548 6616 12549 6656
rect 12507 6607 12549 6616
rect 12891 6656 12933 6665
rect 12891 6616 12892 6656
rect 12932 6616 12933 6656
rect 12891 6607 12933 6616
rect 13275 6656 13317 6665
rect 13275 6616 13276 6656
rect 13316 6616 13317 6656
rect 13275 6607 13317 6616
rect 15291 6656 15333 6665
rect 15291 6616 15292 6656
rect 15332 6616 15333 6656
rect 15291 6607 15333 6616
rect 17403 6656 17445 6665
rect 17403 6616 17404 6656
rect 17444 6616 17445 6656
rect 17403 6607 17445 6616
rect 17787 6656 17829 6665
rect 17787 6616 17788 6656
rect 17828 6616 17829 6656
rect 17787 6607 17829 6616
rect 18459 6656 18501 6665
rect 18459 6616 18460 6656
rect 18500 6616 18501 6656
rect 18459 6607 18501 6616
rect 20043 6656 20085 6665
rect 20043 6616 20044 6656
rect 20084 6616 20085 6656
rect 20043 6607 20085 6616
rect 22155 6656 22197 6665
rect 22155 6616 22156 6656
rect 22196 6616 22197 6656
rect 22155 6607 22197 6616
rect 36747 6656 36789 6665
rect 36747 6616 36748 6656
rect 36788 6616 36789 6656
rect 36747 6607 36789 6616
rect 41835 6656 41877 6665
rect 41835 6616 41836 6656
rect 41876 6616 41877 6656
rect 41835 6607 41877 6616
rect 43995 6656 44037 6665
rect 43995 6616 43996 6656
rect 44036 6616 44037 6656
rect 43995 6607 44037 6616
rect 27963 6572 28005 6581
rect 27963 6532 27964 6572
rect 28004 6532 28005 6572
rect 27963 6523 28005 6532
rect 34347 6572 34389 6581
rect 34347 6532 34348 6572
rect 34388 6532 34389 6572
rect 34347 6523 34389 6532
rect 35307 6572 35349 6581
rect 35307 6532 35308 6572
rect 35348 6532 35349 6572
rect 35307 6523 35349 6532
rect 36555 6572 36597 6581
rect 36555 6532 36556 6572
rect 36596 6532 36597 6572
rect 36555 6523 36597 6532
rect 42795 6572 42837 6581
rect 42795 6532 42796 6572
rect 42836 6532 42837 6572
rect 42795 6523 42837 6532
rect 1227 6488 1269 6497
rect 1227 6448 1228 6488
rect 1268 6448 1269 6488
rect 1227 6439 1269 6448
rect 1611 6488 1653 6497
rect 1611 6448 1612 6488
rect 1652 6448 1653 6488
rect 1611 6439 1653 6448
rect 6219 6488 6261 6497
rect 6219 6448 6220 6488
rect 6260 6448 6261 6488
rect 6219 6439 6261 6448
rect 7642 6488 7700 6489
rect 7642 6448 7651 6488
rect 7691 6448 7700 6488
rect 7642 6447 7700 6448
rect 9483 6488 9525 6497
rect 9483 6448 9484 6488
rect 9524 6448 9525 6488
rect 9483 6439 9525 6448
rect 9867 6488 9909 6497
rect 9867 6448 9868 6488
rect 9908 6448 9909 6488
rect 9867 6439 9909 6448
rect 10827 6488 10869 6497
rect 10827 6448 10828 6488
rect 10868 6448 10869 6488
rect 10827 6439 10869 6448
rect 12267 6488 12309 6497
rect 12267 6448 12268 6488
rect 12308 6448 12309 6488
rect 12267 6439 12309 6448
rect 12651 6488 12693 6497
rect 12651 6448 12652 6488
rect 12692 6448 12693 6488
rect 12651 6439 12693 6448
rect 13035 6488 13077 6497
rect 13035 6448 13036 6488
rect 13076 6448 13077 6488
rect 13035 6439 13077 6448
rect 15531 6488 15573 6497
rect 15531 6448 15532 6488
rect 15572 6448 15573 6488
rect 15531 6439 15573 6448
rect 17643 6488 17685 6497
rect 17643 6448 17644 6488
rect 17684 6448 17685 6488
rect 17643 6439 17685 6448
rect 18027 6488 18069 6497
rect 18027 6448 18028 6488
rect 18068 6448 18069 6488
rect 18027 6439 18069 6448
rect 18219 6488 18261 6497
rect 18219 6448 18220 6488
rect 18260 6448 18261 6488
rect 18219 6439 18261 6448
rect 20235 6488 20277 6497
rect 20235 6448 20236 6488
rect 20276 6448 20277 6488
rect 20235 6439 20277 6448
rect 20475 6488 20517 6497
rect 20475 6448 20476 6488
rect 20516 6448 20517 6488
rect 20475 6439 20517 6448
rect 22923 6488 22965 6497
rect 22923 6448 22924 6488
rect 22964 6448 22965 6488
rect 22923 6439 22965 6448
rect 24555 6488 24597 6497
rect 24555 6448 24556 6488
rect 24596 6448 24597 6488
rect 24555 6439 24597 6448
rect 27147 6488 27189 6497
rect 27147 6448 27148 6488
rect 27188 6448 27189 6488
rect 27147 6439 27189 6448
rect 28203 6488 28245 6497
rect 28203 6448 28204 6488
rect 28244 6448 28245 6488
rect 28203 6439 28245 6448
rect 39531 6488 39573 6497
rect 39531 6448 39532 6488
rect 39572 6448 39573 6488
rect 39531 6439 39573 6448
rect 43179 6488 43221 6497
rect 43179 6448 43180 6488
rect 43220 6448 43221 6488
rect 43179 6439 43221 6448
rect 44235 6488 44277 6497
rect 44235 6448 44236 6488
rect 44276 6448 44277 6488
rect 44235 6439 44277 6448
rect 44523 6488 44565 6497
rect 44523 6448 44524 6488
rect 44564 6448 44565 6488
rect 44523 6439 44565 6448
rect 44907 6488 44949 6497
rect 44907 6448 44908 6488
rect 44948 6448 44949 6488
rect 44907 6439 44949 6448
rect 3723 6404 3765 6413
rect 3723 6364 3724 6404
rect 3764 6364 3765 6404
rect 3723 6355 3765 6364
rect 4963 6404 5021 6405
rect 4963 6364 4972 6404
rect 5012 6364 5021 6404
rect 4963 6363 5021 6364
rect 5722 6404 5780 6405
rect 5722 6364 5731 6404
rect 5771 6364 5780 6404
rect 5722 6363 5780 6364
rect 5835 6404 5877 6413
rect 5835 6364 5836 6404
rect 5876 6364 5877 6404
rect 5835 6355 5877 6364
rect 6315 6404 6357 6413
rect 6315 6364 6316 6404
rect 6356 6364 6357 6404
rect 6315 6355 6357 6364
rect 6787 6404 6845 6405
rect 6787 6364 6796 6404
rect 6836 6364 6845 6404
rect 6787 6363 6845 6364
rect 7306 6404 7364 6405
rect 7306 6364 7315 6404
rect 7355 6364 7364 6404
rect 7306 6363 7364 6364
rect 7843 6404 7901 6405
rect 7843 6364 7852 6404
rect 7892 6364 7901 6404
rect 7843 6363 7901 6364
rect 9099 6404 9141 6413
rect 9099 6364 9100 6404
rect 9140 6364 9141 6404
rect 9099 6355 9141 6364
rect 10317 6403 10359 6412
rect 10317 6363 10318 6403
rect 10358 6363 10359 6403
rect 10317 6354 10359 6363
rect 10443 6404 10485 6413
rect 10443 6364 10444 6404
rect 10484 6364 10485 6404
rect 10443 6355 10485 6364
rect 10923 6404 10965 6413
rect 10923 6364 10924 6404
rect 10964 6364 10965 6404
rect 10923 6355 10965 6364
rect 11395 6404 11453 6405
rect 11395 6364 11404 6404
rect 11444 6364 11453 6404
rect 11395 6363 11453 6364
rect 11914 6404 11972 6405
rect 11914 6364 11923 6404
rect 11963 6364 11972 6404
rect 11914 6363 11972 6364
rect 13603 6404 13661 6405
rect 13603 6364 13612 6404
rect 13652 6364 13661 6404
rect 13603 6363 13661 6364
rect 14859 6404 14901 6413
rect 14859 6364 14860 6404
rect 14900 6364 14901 6404
rect 14859 6355 14901 6364
rect 16003 6404 16061 6405
rect 16003 6364 16012 6404
rect 16052 6364 16061 6404
rect 16003 6363 16061 6364
rect 17259 6404 17301 6413
rect 17259 6364 17260 6404
rect 17300 6364 17301 6404
rect 17259 6355 17301 6364
rect 18603 6404 18645 6413
rect 18603 6364 18604 6404
rect 18644 6364 18645 6404
rect 18603 6355 18645 6364
rect 19843 6404 19901 6405
rect 19843 6364 19852 6404
rect 19892 6364 19901 6404
rect 19843 6363 19901 6364
rect 20715 6404 20757 6413
rect 20715 6364 20716 6404
rect 20756 6364 20757 6404
rect 20715 6355 20757 6364
rect 21963 6404 22021 6405
rect 21963 6364 21972 6404
rect 22012 6364 22021 6404
rect 21963 6363 22021 6364
rect 22426 6404 22484 6405
rect 22426 6364 22435 6404
rect 22475 6364 22484 6404
rect 22426 6363 22484 6364
rect 22539 6404 22581 6413
rect 22539 6364 22540 6404
rect 22580 6364 22581 6404
rect 22539 6355 22581 6364
rect 23019 6404 23061 6413
rect 23019 6364 23020 6404
rect 23060 6364 23061 6404
rect 23019 6355 23061 6364
rect 23491 6404 23549 6405
rect 23491 6364 23500 6404
rect 23540 6364 23549 6404
rect 23491 6363 23549 6364
rect 24010 6404 24068 6405
rect 24010 6364 24019 6404
rect 24059 6364 24068 6404
rect 24010 6363 24068 6364
rect 25219 6404 25277 6405
rect 25219 6364 25228 6404
rect 25268 6364 25277 6404
rect 25219 6363 25277 6364
rect 26475 6404 26517 6413
rect 26475 6364 26476 6404
rect 26516 6364 26517 6404
rect 26475 6355 26517 6364
rect 28675 6404 28733 6405
rect 28675 6364 28684 6404
rect 28724 6364 28733 6404
rect 28675 6363 28733 6364
rect 29931 6404 29973 6413
rect 29931 6364 29932 6404
rect 29972 6364 29973 6404
rect 29931 6355 29973 6364
rect 30315 6404 30357 6413
rect 30315 6364 30316 6404
rect 30356 6364 30357 6404
rect 30315 6355 30357 6364
rect 31555 6404 31613 6405
rect 31555 6364 31564 6404
rect 31604 6364 31613 6404
rect 31555 6363 31613 6364
rect 31947 6404 31989 6413
rect 31947 6364 31948 6404
rect 31988 6364 31989 6404
rect 31947 6355 31989 6364
rect 33187 6404 33245 6405
rect 33187 6364 33196 6404
rect 33236 6364 33245 6404
rect 33187 6363 33245 6364
rect 33675 6404 33717 6413
rect 33675 6364 33676 6404
rect 33716 6364 33717 6404
rect 33675 6355 33717 6364
rect 33946 6404 34004 6405
rect 33946 6364 33955 6404
rect 33995 6364 34004 6404
rect 33946 6363 34004 6364
rect 34635 6404 34677 6413
rect 34635 6364 34636 6404
rect 34676 6364 34677 6404
rect 34635 6355 34677 6364
rect 34906 6404 34964 6405
rect 34906 6364 34915 6404
rect 34955 6364 34964 6404
rect 34906 6363 34964 6364
rect 35883 6404 35925 6413
rect 35883 6364 35884 6404
rect 35924 6364 35925 6404
rect 35883 6355 35925 6364
rect 36130 6404 36188 6405
rect 36130 6364 36139 6404
rect 36179 6364 36188 6404
rect 36130 6363 36188 6364
rect 36250 6404 36308 6405
rect 36250 6364 36259 6404
rect 36299 6364 36308 6404
rect 36250 6363 36308 6364
rect 36931 6404 36989 6405
rect 36931 6364 36940 6404
rect 36980 6364 36989 6404
rect 36931 6363 36989 6364
rect 38187 6404 38229 6413
rect 38187 6364 38188 6404
rect 38228 6364 38229 6404
rect 38187 6355 38229 6364
rect 39021 6404 39063 6413
rect 39021 6364 39022 6404
rect 39062 6364 39063 6404
rect 39021 6355 39063 6364
rect 39147 6404 39189 6413
rect 39147 6364 39148 6404
rect 39188 6364 39189 6404
rect 39147 6355 39189 6364
rect 39627 6404 39669 6413
rect 39627 6364 39628 6404
rect 39668 6364 39669 6404
rect 39627 6355 39669 6364
rect 40099 6404 40157 6405
rect 40099 6364 40108 6404
rect 40148 6364 40157 6404
rect 40099 6363 40157 6364
rect 40587 6404 40645 6405
rect 40587 6364 40596 6404
rect 40636 6364 40645 6404
rect 40587 6363 40645 6364
rect 41163 6404 41205 6413
rect 41163 6364 41164 6404
rect 41204 6364 41205 6404
rect 41163 6355 41205 6364
rect 41434 6404 41492 6405
rect 41434 6364 41443 6404
rect 41483 6364 41492 6404
rect 41434 6363 41492 6364
rect 42123 6404 42165 6413
rect 42123 6364 42124 6404
rect 42164 6364 42165 6404
rect 42123 6355 42165 6364
rect 42394 6404 42452 6405
rect 42394 6364 42403 6404
rect 42443 6364 42452 6404
rect 42394 6363 42452 6364
rect 24315 6320 24357 6329
rect 24315 6280 24316 6320
rect 24356 6280 24357 6320
rect 24315 6271 24357 6280
rect 25035 6320 25077 6329
rect 25035 6280 25036 6320
rect 25076 6280 25077 6320
rect 25035 6271 25077 6280
rect 28491 6320 28533 6329
rect 28491 6280 28492 6320
rect 28532 6280 28533 6320
rect 28491 6271 28533 6280
rect 34059 6320 34101 6329
rect 34059 6280 34060 6320
rect 34100 6280 34101 6320
rect 34059 6271 34101 6280
rect 35019 6320 35061 6329
rect 35019 6280 35020 6320
rect 35060 6280 35061 6320
rect 35019 6271 35061 6280
rect 41547 6320 41589 6329
rect 41547 6280 41548 6320
rect 41588 6280 41589 6320
rect 41547 6271 41589 6280
rect 42507 6320 42549 6329
rect 42507 6280 42508 6320
rect 42548 6280 42549 6320
rect 42507 6271 42549 6280
rect 45147 6320 45189 6329
rect 45147 6280 45148 6320
rect 45188 6280 45189 6320
rect 45147 6271 45189 6280
rect 1467 6236 1509 6245
rect 1467 6196 1468 6236
rect 1508 6196 1509 6236
rect 1467 6187 1509 6196
rect 1851 6236 1893 6245
rect 1851 6196 1852 6236
rect 1892 6196 1893 6236
rect 1851 6187 1893 6196
rect 5163 6236 5205 6245
rect 5163 6196 5164 6236
rect 5204 6196 5205 6236
rect 5163 6187 5205 6196
rect 7467 6236 7509 6245
rect 7467 6196 7468 6236
rect 7508 6196 7509 6236
rect 7467 6187 7509 6196
rect 9723 6236 9765 6245
rect 9723 6196 9724 6236
rect 9764 6196 9765 6236
rect 9723 6187 9765 6196
rect 12075 6236 12117 6245
rect 12075 6196 12076 6236
rect 12116 6196 12117 6236
rect 12075 6187 12117 6196
rect 13419 6236 13461 6245
rect 13419 6196 13420 6236
rect 13460 6196 13461 6236
rect 13419 6187 13461 6196
rect 15819 6236 15861 6245
rect 15819 6196 15820 6236
rect 15860 6196 15861 6236
rect 15819 6187 15861 6196
rect 24171 6236 24213 6245
rect 24171 6196 24172 6236
rect 24212 6196 24213 6236
rect 24171 6187 24213 6196
rect 27387 6236 27429 6245
rect 27387 6196 27388 6236
rect 27428 6196 27429 6236
rect 27387 6187 27429 6196
rect 31755 6236 31797 6245
rect 31755 6196 31756 6236
rect 31796 6196 31797 6236
rect 31755 6187 31797 6196
rect 33387 6236 33429 6245
rect 33387 6196 33388 6236
rect 33428 6196 33429 6236
rect 33387 6187 33429 6196
rect 40779 6236 40821 6245
rect 40779 6196 40780 6236
rect 40820 6196 40821 6236
rect 40779 6187 40821 6196
rect 42939 6236 42981 6245
rect 42939 6196 42940 6236
rect 42980 6196 42981 6236
rect 42939 6187 42981 6196
rect 43546 6236 43604 6237
rect 43546 6196 43555 6236
rect 43595 6196 43604 6236
rect 43546 6195 43604 6196
rect 43834 6236 43892 6237
rect 43834 6196 43843 6236
rect 43883 6196 43892 6236
rect 43834 6195 43892 6196
rect 44763 6236 44805 6245
rect 44763 6196 44764 6236
rect 44804 6196 44805 6236
rect 44763 6187 44805 6196
rect 1152 6068 45216 6092
rect 1152 6028 4928 6068
rect 4968 6028 5010 6068
rect 5050 6028 5092 6068
rect 5132 6028 5174 6068
rect 5214 6028 5256 6068
rect 5296 6028 20048 6068
rect 20088 6028 20130 6068
rect 20170 6028 20212 6068
rect 20252 6028 20294 6068
rect 20334 6028 20376 6068
rect 20416 6028 35168 6068
rect 35208 6028 35250 6068
rect 35290 6028 35332 6068
rect 35372 6028 35414 6068
rect 35454 6028 35496 6068
rect 35536 6028 45216 6068
rect 1152 6004 45216 6028
rect 32475 5900 32517 5909
rect 32475 5860 32476 5900
rect 32516 5860 32517 5900
rect 32475 5851 32517 5860
rect 41931 5900 41973 5909
rect 41931 5860 41932 5900
rect 41972 5860 41973 5900
rect 41931 5851 41973 5860
rect 43162 5900 43220 5901
rect 43162 5860 43171 5900
rect 43211 5860 43220 5900
rect 43162 5859 43220 5860
rect 43450 5900 43508 5901
rect 43450 5860 43459 5900
rect 43499 5860 43508 5900
rect 43450 5859 43508 5860
rect 44235 5900 44277 5909
rect 44235 5860 44236 5900
rect 44276 5860 44277 5900
rect 44235 5851 44277 5860
rect 6027 5816 6069 5825
rect 6027 5776 6028 5816
rect 6068 5776 6069 5816
rect 6027 5767 6069 5776
rect 8811 5816 8853 5825
rect 8811 5776 8812 5816
rect 8852 5776 8853 5816
rect 8811 5767 8853 5776
rect 11115 5816 11157 5825
rect 11115 5776 11116 5816
rect 11156 5776 11157 5816
rect 11115 5767 11157 5776
rect 11835 5816 11877 5825
rect 11835 5776 11836 5816
rect 11876 5776 11877 5816
rect 11835 5767 11877 5776
rect 23691 5816 23733 5825
rect 23691 5776 23692 5816
rect 23732 5776 23733 5816
rect 23691 5767 23733 5776
rect 3531 5732 3573 5741
rect 5643 5732 5685 5741
rect 3531 5692 3532 5732
rect 3572 5692 3573 5732
rect 3531 5683 3573 5692
rect 4783 5723 4825 5732
rect 4783 5683 4784 5723
rect 4824 5683 4825 5723
rect 5643 5692 5644 5732
rect 5684 5692 5685 5732
rect 5643 5683 5685 5692
rect 5914 5732 5972 5733
rect 5914 5692 5923 5732
rect 5963 5692 5972 5732
rect 5914 5691 5972 5692
rect 8932 5732 8990 5733
rect 8932 5692 8941 5732
rect 8981 5692 8990 5732
rect 8932 5691 8990 5692
rect 9195 5732 9237 5741
rect 9195 5692 9196 5732
rect 9236 5692 9237 5732
rect 9195 5683 9237 5692
rect 10731 5732 10773 5741
rect 10731 5692 10732 5732
rect 10772 5692 10773 5732
rect 10731 5683 10773 5692
rect 11002 5732 11060 5733
rect 14723 5732 14765 5741
rect 17163 5732 17205 5741
rect 11002 5692 11011 5732
rect 11051 5692 11060 5732
rect 11002 5691 11060 5692
rect 13515 5723 13557 5732
rect 13515 5683 13516 5723
rect 13556 5683 13557 5723
rect 14723 5692 14724 5732
rect 14764 5692 14765 5732
rect 14723 5683 14765 5692
rect 15915 5723 15957 5732
rect 15915 5683 15916 5723
rect 15956 5683 15957 5723
rect 17163 5692 17164 5732
rect 17204 5692 17205 5732
rect 17163 5683 17205 5692
rect 18027 5732 18069 5741
rect 20043 5732 20085 5741
rect 23307 5732 23349 5741
rect 18027 5692 18028 5732
rect 18068 5692 18069 5732
rect 18027 5683 18069 5692
rect 19275 5723 19317 5732
rect 19275 5683 19276 5723
rect 19316 5683 19317 5723
rect 20043 5692 20044 5732
rect 20084 5692 20085 5732
rect 20043 5683 20085 5692
rect 21291 5723 21333 5732
rect 21291 5683 21292 5723
rect 21332 5683 21333 5723
rect 23307 5692 23308 5732
rect 23348 5692 23349 5732
rect 23307 5683 23349 5692
rect 23578 5732 23636 5733
rect 27147 5732 27189 5741
rect 23578 5692 23587 5732
rect 23627 5692 23636 5732
rect 23578 5691 23636 5692
rect 25899 5723 25941 5732
rect 25899 5683 25900 5723
rect 25940 5683 25941 5723
rect 27147 5692 27148 5732
rect 27188 5692 27189 5732
rect 27147 5683 27189 5692
rect 27627 5732 27669 5741
rect 30507 5732 30549 5741
rect 33370 5732 33428 5733
rect 27627 5692 27628 5732
rect 27668 5692 27669 5732
rect 27627 5683 27669 5692
rect 28875 5723 28917 5732
rect 28875 5683 28876 5723
rect 28916 5683 28917 5723
rect 30507 5692 30508 5732
rect 30548 5692 30549 5732
rect 30507 5683 30549 5692
rect 31755 5723 31797 5732
rect 31755 5683 31756 5723
rect 31796 5683 31797 5723
rect 33370 5692 33379 5732
rect 33419 5692 33428 5732
rect 33370 5691 33428 5692
rect 33483 5732 33525 5741
rect 35146 5732 35204 5733
rect 33483 5692 33484 5732
rect 33524 5692 33525 5732
rect 33483 5683 33525 5692
rect 34443 5723 34485 5732
rect 34443 5683 34444 5723
rect 34484 5683 34485 5723
rect 4783 5674 4825 5683
rect 13515 5674 13557 5683
rect 15915 5674 15957 5683
rect 19275 5674 19317 5683
rect 21291 5674 21333 5683
rect 25899 5674 25941 5683
rect 28875 5674 28917 5683
rect 31755 5674 31797 5683
rect 34443 5674 34485 5683
rect 34923 5723 34965 5732
rect 34923 5683 34924 5723
rect 34964 5683 34965 5723
rect 35146 5692 35155 5732
rect 35195 5692 35204 5732
rect 35146 5691 35204 5692
rect 38571 5732 38613 5741
rect 40491 5732 40533 5741
rect 38571 5692 38572 5732
rect 38612 5692 38613 5732
rect 38571 5683 38613 5692
rect 39819 5723 39861 5732
rect 39819 5683 39820 5723
rect 39860 5683 39861 5723
rect 40491 5692 40492 5732
rect 40532 5692 40533 5732
rect 40491 5683 40533 5692
rect 41739 5723 41781 5732
rect 41739 5683 41740 5723
rect 41780 5683 41781 5723
rect 34923 5674 34965 5683
rect 39819 5674 39861 5683
rect 41739 5674 41781 5683
rect 1227 5648 1269 5657
rect 1227 5608 1228 5648
rect 1268 5608 1269 5648
rect 1227 5599 1269 5608
rect 1611 5648 1653 5657
rect 1611 5608 1612 5648
rect 1652 5608 1653 5648
rect 1611 5599 1653 5608
rect 1995 5648 2037 5657
rect 1995 5608 1996 5648
rect 2036 5608 2037 5648
rect 1995 5599 2037 5608
rect 6507 5648 6549 5657
rect 6507 5608 6508 5648
rect 6548 5608 6549 5648
rect 6507 5599 6549 5608
rect 10251 5648 10293 5657
rect 10251 5608 10252 5648
rect 10292 5608 10293 5648
rect 10251 5599 10293 5608
rect 11595 5648 11637 5657
rect 11595 5608 11596 5648
rect 11636 5608 11637 5648
rect 11595 5599 11637 5608
rect 11979 5648 12021 5657
rect 11979 5608 11980 5648
rect 12020 5608 12021 5648
rect 11979 5599 12021 5608
rect 12411 5648 12453 5657
rect 12411 5608 12412 5648
rect 12452 5608 12453 5648
rect 12411 5599 12453 5608
rect 12651 5648 12693 5657
rect 12651 5608 12652 5648
rect 12692 5608 12693 5648
rect 12651 5599 12693 5608
rect 12843 5648 12885 5657
rect 12843 5608 12844 5648
rect 12884 5608 12885 5648
rect 12843 5599 12885 5608
rect 13306 5648 13364 5649
rect 13306 5608 13315 5648
rect 13355 5608 13364 5648
rect 13306 5607 13364 5608
rect 14955 5648 14997 5657
rect 14955 5608 14956 5648
rect 14996 5608 14997 5648
rect 14955 5599 14997 5608
rect 15531 5648 15573 5657
rect 15531 5608 15532 5648
rect 15572 5608 15573 5648
rect 15531 5599 15573 5608
rect 22107 5648 22149 5657
rect 22107 5608 22108 5648
rect 22148 5608 22149 5648
rect 22107 5599 22149 5608
rect 22347 5648 22389 5657
rect 22347 5608 22348 5648
rect 22388 5608 22389 5648
rect 22347 5599 22389 5608
rect 24363 5648 24405 5657
rect 24363 5608 24364 5648
rect 24404 5608 24405 5648
rect 24363 5599 24405 5608
rect 25323 5648 25365 5657
rect 25323 5608 25324 5648
rect 25364 5608 25365 5648
rect 25323 5599 25365 5608
rect 25690 5648 25748 5649
rect 25690 5608 25699 5648
rect 25739 5608 25748 5648
rect 25690 5607 25748 5608
rect 29451 5648 29493 5657
rect 29451 5608 29452 5648
rect 29492 5608 29493 5648
rect 29451 5599 29493 5608
rect 29835 5648 29877 5657
rect 29835 5608 29836 5648
rect 29876 5608 29877 5648
rect 29835 5599 29877 5608
rect 32331 5648 32373 5657
rect 32331 5608 32332 5648
rect 32372 5608 32373 5648
rect 32331 5599 32373 5608
rect 32715 5648 32757 5657
rect 32715 5608 32716 5648
rect 32756 5608 32757 5648
rect 32715 5599 32757 5608
rect 33099 5648 33141 5657
rect 33099 5608 33100 5648
rect 33140 5608 33141 5648
rect 33099 5599 33141 5608
rect 33871 5648 33913 5657
rect 33871 5608 33872 5648
rect 33912 5608 33913 5648
rect 33871 5599 33913 5608
rect 33994 5648 34052 5649
rect 33994 5608 34003 5648
rect 34043 5608 34052 5648
rect 33994 5607 34052 5608
rect 35259 5648 35301 5657
rect 35259 5608 35260 5648
rect 35300 5608 35301 5648
rect 35259 5599 35301 5608
rect 35499 5648 35541 5657
rect 35499 5608 35500 5648
rect 35540 5608 35541 5648
rect 35499 5599 35541 5608
rect 35883 5648 35925 5657
rect 35883 5608 35884 5648
rect 35924 5608 35925 5648
rect 35883 5599 35925 5608
rect 36267 5648 36309 5657
rect 36267 5608 36268 5648
rect 36308 5608 36309 5648
rect 36267 5599 36309 5608
rect 37179 5648 37221 5657
rect 37179 5608 37180 5648
rect 37220 5608 37221 5648
rect 37179 5599 37221 5608
rect 37419 5648 37461 5657
rect 37419 5608 37420 5648
rect 37460 5608 37461 5648
rect 37419 5599 37461 5608
rect 37995 5648 38037 5657
rect 37995 5608 37996 5648
rect 38036 5608 38037 5648
rect 37995 5599 38037 5608
rect 42891 5648 42933 5657
rect 42891 5608 42892 5648
rect 42932 5608 42933 5648
rect 42891 5599 42933 5608
rect 43179 5648 43221 5657
rect 43179 5608 43180 5648
rect 43220 5608 43221 5648
rect 43179 5599 43221 5608
rect 43755 5648 43797 5657
rect 43755 5608 43756 5648
rect 43796 5608 43797 5648
rect 43755 5599 43797 5608
rect 44331 5648 44373 5657
rect 44331 5608 44332 5648
rect 44372 5608 44373 5648
rect 44331 5599 44373 5608
rect 44523 5648 44565 5657
rect 44523 5608 44524 5648
rect 44564 5608 44565 5648
rect 44523 5599 44565 5608
rect 44907 5648 44949 5657
rect 44907 5608 44908 5648
rect 44948 5608 44949 5648
rect 44907 5599 44949 5608
rect 45147 5648 45189 5657
rect 45147 5608 45148 5648
rect 45188 5608 45189 5648
rect 45147 5599 45189 5608
rect 2235 5564 2277 5573
rect 2235 5524 2236 5564
rect 2276 5524 2277 5564
rect 2235 5515 2277 5524
rect 6315 5564 6357 5573
rect 6315 5524 6316 5564
rect 6356 5524 6357 5564
rect 6315 5515 6357 5524
rect 11403 5564 11445 5573
rect 11403 5524 11404 5564
rect 11444 5524 11445 5564
rect 11403 5515 11445 5524
rect 15195 5564 15237 5573
rect 15195 5524 15196 5564
rect 15236 5524 15237 5564
rect 15195 5515 15237 5524
rect 19467 5564 19509 5573
rect 19467 5524 19468 5564
rect 19508 5524 19509 5564
rect 19467 5515 19509 5524
rect 21483 5564 21525 5573
rect 21483 5524 21484 5564
rect 21524 5524 21525 5564
rect 21483 5515 21525 5524
rect 24123 5564 24165 5573
rect 24123 5524 24124 5564
rect 24164 5524 24165 5564
rect 24123 5515 24165 5524
rect 25563 5564 25605 5573
rect 25563 5524 25564 5564
rect 25604 5524 25605 5564
rect 25563 5515 25605 5524
rect 29067 5564 29109 5573
rect 29067 5524 29068 5564
rect 29108 5524 29109 5564
rect 29067 5515 29109 5524
rect 31947 5564 31989 5573
rect 31947 5524 31948 5564
rect 31988 5524 31989 5564
rect 31947 5515 31989 5524
rect 32091 5564 32133 5573
rect 32091 5524 32092 5564
rect 32132 5524 32133 5564
rect 32091 5515 32133 5524
rect 1467 5480 1509 5489
rect 1467 5440 1468 5480
rect 1508 5440 1509 5480
rect 1467 5431 1509 5440
rect 1851 5480 1893 5489
rect 1851 5440 1852 5480
rect 1892 5440 1893 5480
rect 1851 5431 1893 5440
rect 4971 5480 5013 5489
rect 4971 5440 4972 5480
rect 5012 5440 5013 5480
rect 4971 5431 5013 5440
rect 6747 5480 6789 5489
rect 6747 5440 6748 5480
rect 6788 5440 6789 5480
rect 6747 5431 6789 5440
rect 8523 5480 8565 5489
rect 8523 5440 8524 5480
rect 8564 5440 8565 5480
rect 8523 5431 8565 5440
rect 10491 5480 10533 5489
rect 10491 5440 10492 5480
rect 10532 5440 10533 5480
rect 10491 5431 10533 5440
rect 12219 5480 12261 5489
rect 12219 5440 12220 5480
rect 12260 5440 12261 5480
rect 12219 5431 12261 5440
rect 13083 5480 13125 5489
rect 13083 5440 13084 5480
rect 13124 5440 13125 5480
rect 13083 5431 13125 5440
rect 15291 5480 15333 5489
rect 15291 5440 15292 5480
rect 15332 5440 15333 5480
rect 15291 5431 15333 5440
rect 15723 5480 15765 5489
rect 15723 5440 15724 5480
rect 15764 5440 15765 5480
rect 15723 5431 15765 5440
rect 23979 5480 24021 5489
rect 23979 5440 23980 5480
rect 24020 5440 24021 5480
rect 23979 5431 24021 5440
rect 29211 5480 29253 5489
rect 29211 5440 29212 5480
rect 29252 5440 29253 5480
rect 29211 5431 29253 5440
rect 30075 5480 30117 5489
rect 30075 5440 30076 5480
rect 30116 5440 30117 5480
rect 30075 5431 30117 5440
rect 32859 5480 32901 5489
rect 32859 5440 32860 5480
rect 32900 5440 32901 5480
rect 32859 5431 32901 5440
rect 35643 5480 35685 5489
rect 35643 5440 35644 5480
rect 35684 5440 35685 5480
rect 35643 5431 35685 5440
rect 36027 5480 36069 5489
rect 36027 5440 36028 5480
rect 36068 5440 36069 5480
rect 36027 5431 36069 5440
rect 38235 5480 38277 5489
rect 38235 5440 38236 5480
rect 38276 5440 38277 5480
rect 38235 5431 38277 5440
rect 40011 5480 40053 5489
rect 40011 5440 40012 5480
rect 40052 5440 40053 5480
rect 40011 5431 40053 5440
rect 44763 5480 44805 5489
rect 44763 5440 44764 5480
rect 44804 5440 44805 5480
rect 44763 5431 44805 5440
rect 1152 5312 45216 5336
rect 1152 5272 3688 5312
rect 3728 5272 3770 5312
rect 3810 5272 3852 5312
rect 3892 5272 3934 5312
rect 3974 5272 4016 5312
rect 4056 5272 18808 5312
rect 18848 5272 18890 5312
rect 18930 5272 18972 5312
rect 19012 5272 19054 5312
rect 19094 5272 19136 5312
rect 19176 5272 33928 5312
rect 33968 5272 34010 5312
rect 34050 5272 34092 5312
rect 34132 5272 34174 5312
rect 34214 5272 34256 5312
rect 34296 5272 45216 5312
rect 1152 5248 45216 5272
rect 6123 5144 6165 5153
rect 6123 5104 6124 5144
rect 6164 5104 6165 5144
rect 6123 5095 6165 5104
rect 11451 5144 11493 5153
rect 11451 5104 11452 5144
rect 11492 5104 11493 5144
rect 11451 5095 11493 5104
rect 12363 5144 12405 5153
rect 12363 5104 12364 5144
rect 12404 5104 12405 5144
rect 12363 5095 12405 5104
rect 14235 5144 14277 5153
rect 14235 5104 14236 5144
rect 14276 5104 14277 5144
rect 14235 5095 14277 5104
rect 36363 5144 36405 5153
rect 36363 5104 36364 5144
rect 36404 5104 36405 5144
rect 36363 5095 36405 5104
rect 7083 5060 7125 5069
rect 7083 5020 7084 5060
rect 7124 5020 7125 5060
rect 7083 5011 7125 5020
rect 14619 5060 14661 5069
rect 14619 5020 14620 5060
rect 14660 5020 14661 5060
rect 14619 5011 14661 5020
rect 33771 5060 33813 5069
rect 33771 5020 33772 5060
rect 33812 5020 33813 5060
rect 33771 5011 33813 5020
rect 39195 5060 39237 5069
rect 39195 5020 39196 5060
rect 39236 5020 39237 5060
rect 39195 5011 39237 5020
rect 41451 5060 41493 5069
rect 41451 5020 41452 5060
rect 41492 5020 41493 5060
rect 41451 5011 41493 5020
rect 1227 4976 1269 4985
rect 1227 4936 1228 4976
rect 1268 4936 1269 4976
rect 1227 4927 1269 4936
rect 1611 4976 1653 4985
rect 1611 4936 1612 4976
rect 1652 4936 1653 4976
rect 1611 4927 1653 4936
rect 9771 4976 9813 4985
rect 9771 4936 9772 4976
rect 9812 4936 9813 4976
rect 9771 4927 9813 4936
rect 11691 4976 11733 4985
rect 11691 4936 11692 4976
rect 11732 4936 11733 4976
rect 11691 4927 11733 4936
rect 11883 4976 11925 4985
rect 11883 4936 11884 4976
rect 11924 4936 11925 4976
rect 11883 4927 11925 4936
rect 14475 4976 14517 4985
rect 14475 4936 14476 4976
rect 14516 4936 14517 4976
rect 14475 4927 14517 4936
rect 14859 4976 14901 4985
rect 14859 4936 14860 4976
rect 14900 4936 14901 4976
rect 14859 4927 14901 4936
rect 19755 4976 19797 4985
rect 19755 4936 19756 4976
rect 19796 4936 19797 4976
rect 19755 4927 19797 4936
rect 20091 4976 20133 4985
rect 20091 4936 20092 4976
rect 20132 4936 20133 4976
rect 20091 4927 20133 4936
rect 20331 4976 20373 4985
rect 20331 4936 20332 4976
rect 20372 4936 20373 4976
rect 20331 4927 20373 4936
rect 25995 4976 26037 4985
rect 25995 4936 25996 4976
rect 26036 4936 26037 4976
rect 25995 4927 26037 4936
rect 29163 4976 29205 4985
rect 29163 4936 29164 4976
rect 29204 4936 29205 4976
rect 29163 4927 29205 4936
rect 34155 4976 34197 4985
rect 34155 4936 34156 4976
rect 34196 4936 34197 4976
rect 34155 4927 34197 4936
rect 38955 4976 38997 4985
rect 38955 4936 38956 4976
rect 38996 4936 38997 4976
rect 38955 4927 38997 4936
rect 40299 4976 40341 4985
rect 40299 4936 40300 4976
rect 40340 4936 40341 4976
rect 40299 4927 40341 4936
rect 44091 4976 44133 4985
rect 44091 4936 44092 4976
rect 44132 4936 44133 4976
rect 44091 4927 44133 4936
rect 44331 4976 44373 4985
rect 44331 4936 44332 4976
rect 44372 4936 44373 4976
rect 44331 4927 44373 4936
rect 44523 4976 44565 4985
rect 44523 4936 44524 4976
rect 44564 4936 44565 4976
rect 44523 4927 44565 4936
rect 44907 4976 44949 4985
rect 44907 4936 44908 4976
rect 44948 4936 44949 4976
rect 44907 4927 44949 4936
rect 45147 4976 45189 4985
rect 45147 4936 45148 4976
rect 45188 4936 45189 4976
rect 45147 4927 45189 4936
rect 5451 4892 5493 4901
rect 5451 4852 5452 4892
rect 5492 4852 5493 4892
rect 5451 4843 5493 4852
rect 5722 4892 5780 4893
rect 5722 4852 5731 4892
rect 5771 4852 5780 4892
rect 5722 4851 5780 4852
rect 6411 4892 6453 4901
rect 6411 4852 6412 4892
rect 6452 4852 6453 4892
rect 6411 4843 6453 4852
rect 6682 4892 6740 4893
rect 6682 4852 6691 4892
rect 6731 4852 6740 4892
rect 6682 4851 6740 4852
rect 7563 4892 7605 4901
rect 7563 4852 7564 4892
rect 7604 4852 7605 4892
rect 7563 4843 7605 4852
rect 8803 4892 8861 4893
rect 8803 4852 8812 4892
rect 8852 4852 8861 4892
rect 8803 4851 8861 4852
rect 9274 4892 9332 4893
rect 9274 4852 9283 4892
rect 9323 4852 9332 4892
rect 9274 4851 9332 4852
rect 9387 4892 9429 4901
rect 9387 4852 9388 4892
rect 9428 4852 9429 4892
rect 9387 4843 9429 4852
rect 9867 4892 9909 4901
rect 9867 4852 9868 4892
rect 9908 4852 9909 4892
rect 9867 4843 9909 4852
rect 10339 4892 10397 4893
rect 10339 4852 10348 4892
rect 10388 4852 10397 4892
rect 10339 4851 10397 4852
rect 10858 4892 10916 4893
rect 10858 4852 10867 4892
rect 10907 4852 10916 4892
rect 10858 4851 10916 4852
rect 12547 4892 12605 4893
rect 12547 4852 12556 4892
rect 12596 4852 12605 4892
rect 12547 4851 12605 4852
rect 13803 4892 13845 4901
rect 13803 4852 13804 4892
rect 13844 4852 13845 4892
rect 13803 4843 13845 4852
rect 15235 4892 15293 4893
rect 15235 4852 15244 4892
rect 15284 4852 15293 4892
rect 15235 4851 15293 4852
rect 16491 4892 16533 4901
rect 16491 4852 16492 4892
rect 16532 4852 16533 4892
rect 16491 4843 16533 4852
rect 17067 4892 17109 4901
rect 17067 4852 17068 4892
rect 17108 4852 17109 4892
rect 17067 4843 17109 4852
rect 18307 4892 18365 4893
rect 18307 4852 18316 4892
rect 18356 4852 18365 4892
rect 18307 4851 18365 4852
rect 21099 4892 21141 4901
rect 21099 4852 21100 4892
rect 21140 4852 21141 4892
rect 21099 4843 21141 4852
rect 22347 4892 22405 4893
rect 22347 4852 22356 4892
rect 22396 4852 22405 4892
rect 22347 4851 22405 4852
rect 22923 4892 22965 4901
rect 22923 4852 22924 4892
rect 22964 4852 22965 4892
rect 22923 4843 22965 4852
rect 24163 4892 24221 4893
rect 24163 4852 24172 4892
rect 24212 4852 24221 4892
rect 24163 4851 24221 4852
rect 33099 4892 33141 4901
rect 33099 4852 33100 4892
rect 33140 4852 33141 4892
rect 33099 4843 33141 4852
rect 33370 4892 33428 4893
rect 33370 4852 33379 4892
rect 33419 4852 33428 4892
rect 33370 4851 33428 4852
rect 34923 4892 34965 4901
rect 34923 4852 34924 4892
rect 34964 4852 34965 4892
rect 34923 4843 34965 4852
rect 36163 4892 36221 4893
rect 36163 4852 36172 4892
rect 36212 4852 36221 4892
rect 36163 4851 36221 4852
rect 37323 4892 37365 4901
rect 37323 4852 37324 4892
rect 37364 4852 37365 4892
rect 37323 4843 37365 4852
rect 38563 4892 38621 4893
rect 38563 4852 38572 4892
rect 38612 4852 38621 4892
rect 38563 4851 38621 4852
rect 40779 4892 40821 4901
rect 40779 4852 40780 4892
rect 40820 4852 40821 4892
rect 40779 4843 40821 4852
rect 41050 4892 41108 4893
rect 41050 4852 41059 4892
rect 41099 4852 41108 4892
rect 41050 4851 41108 4852
rect 1467 4808 1509 4817
rect 1467 4768 1468 4808
rect 1508 4768 1509 4808
rect 1467 4759 1509 4768
rect 5835 4808 5877 4817
rect 5835 4768 5836 4808
rect 5876 4768 5877 4808
rect 5835 4759 5877 4768
rect 6795 4808 6837 4817
rect 6795 4768 6796 4808
rect 6836 4768 6837 4808
rect 6795 4759 6837 4768
rect 9003 4808 9045 4817
rect 9003 4768 9004 4808
rect 9044 4768 9045 4808
rect 9003 4759 9045 4768
rect 14235 4808 14277 4817
rect 14235 4768 14236 4808
rect 14276 4768 14277 4808
rect 14235 4759 14277 4768
rect 19995 4808 20037 4817
rect 19995 4768 19996 4808
rect 20036 4768 20037 4808
rect 19995 4759 20037 4768
rect 29403 4808 29445 4817
rect 29403 4768 29404 4808
rect 29444 4768 29445 4808
rect 29403 4759 29445 4768
rect 33483 4808 33525 4817
rect 33483 4768 33484 4808
rect 33524 4768 33525 4808
rect 33483 4759 33525 4768
rect 33915 4808 33957 4817
rect 33915 4768 33916 4808
rect 33956 4768 33957 4808
rect 33915 4759 33957 4768
rect 41163 4808 41205 4817
rect 41163 4768 41164 4808
rect 41204 4768 41205 4808
rect 41163 4759 41205 4768
rect 1851 4724 1893 4733
rect 1851 4684 1852 4724
rect 1892 4684 1893 4724
rect 1851 4675 1893 4684
rect 11019 4724 11061 4733
rect 11019 4684 11020 4724
rect 11060 4684 11061 4724
rect 11019 4675 11061 4684
rect 12123 4724 12165 4733
rect 12123 4684 12124 4724
rect 12164 4684 12165 4724
rect 12123 4675 12165 4684
rect 15051 4724 15093 4733
rect 15051 4684 15052 4724
rect 15092 4684 15093 4724
rect 15051 4675 15093 4684
rect 18507 4724 18549 4733
rect 18507 4684 18508 4724
rect 18548 4684 18549 4724
rect 18507 4675 18549 4684
rect 22539 4724 22581 4733
rect 22539 4684 22540 4724
rect 22580 4684 22581 4724
rect 22539 4675 22581 4684
rect 24363 4724 24405 4733
rect 24363 4684 24364 4724
rect 24404 4684 24405 4724
rect 24363 4675 24405 4684
rect 26235 4724 26277 4733
rect 26235 4684 26236 4724
rect 26276 4684 26277 4724
rect 26235 4675 26277 4684
rect 38763 4724 38805 4733
rect 38763 4684 38764 4724
rect 38804 4684 38805 4724
rect 38763 4675 38805 4684
rect 40539 4724 40581 4733
rect 40539 4684 40540 4724
rect 40580 4684 40581 4724
rect 40539 4675 40581 4684
rect 42970 4724 43028 4725
rect 42970 4684 42979 4724
rect 43019 4684 43028 4724
rect 42970 4683 43028 4684
rect 43258 4724 43316 4725
rect 43258 4684 43267 4724
rect 43307 4684 43316 4724
rect 43258 4683 43316 4684
rect 43834 4724 43892 4725
rect 43834 4684 43843 4724
rect 43883 4684 43892 4724
rect 43834 4683 43892 4684
rect 44763 4724 44805 4733
rect 44763 4684 44764 4724
rect 44804 4684 44805 4724
rect 44763 4675 44805 4684
rect 1152 4556 45216 4580
rect 1152 4516 4928 4556
rect 4968 4516 5010 4556
rect 5050 4516 5092 4556
rect 5132 4516 5174 4556
rect 5214 4516 5256 4556
rect 5296 4516 20048 4556
rect 20088 4516 20130 4556
rect 20170 4516 20212 4556
rect 20252 4516 20294 4556
rect 20334 4516 20376 4556
rect 20416 4516 35168 4556
rect 35208 4516 35250 4556
rect 35290 4516 35332 4556
rect 35372 4516 35414 4556
rect 35454 4516 35496 4556
rect 35536 4516 45216 4556
rect 1152 4492 45216 4516
rect 24027 4388 24069 4397
rect 24027 4348 24028 4388
rect 24068 4348 24069 4388
rect 24027 4339 24069 4348
rect 42202 4388 42260 4389
rect 42202 4348 42211 4388
rect 42251 4348 42260 4388
rect 42202 4347 42260 4348
rect 42490 4388 42548 4389
rect 42490 4348 42499 4388
rect 42539 4348 42548 4388
rect 42490 4347 42548 4348
rect 42778 4388 42836 4389
rect 42778 4348 42787 4388
rect 42827 4348 42836 4388
rect 42778 4347 42836 4348
rect 43546 4388 43604 4389
rect 43546 4348 43555 4388
rect 43595 4348 43604 4388
rect 43546 4347 43604 4348
rect 44218 4388 44276 4389
rect 44218 4348 44227 4388
rect 44267 4348 44276 4388
rect 44218 4347 44276 4348
rect 6219 4304 6261 4313
rect 6219 4264 6220 4304
rect 6260 4264 6261 4304
rect 6219 4255 6261 4264
rect 8842 4304 8900 4305
rect 8842 4264 8851 4304
rect 8891 4264 8900 4304
rect 8842 4263 8900 4264
rect 9243 4304 9285 4313
rect 9243 4264 9244 4304
rect 9284 4264 9285 4304
rect 9243 4255 9285 4264
rect 9867 4304 9909 4313
rect 9867 4264 9868 4304
rect 9908 4264 9909 4304
rect 9867 4255 9909 4264
rect 11259 4304 11301 4313
rect 11259 4264 11260 4304
rect 11300 4264 11301 4304
rect 11259 4255 11301 4264
rect 13707 4304 13749 4313
rect 13707 4264 13708 4304
rect 13748 4264 13749 4304
rect 13707 4255 13749 4264
rect 15243 4304 15285 4313
rect 15243 4264 15244 4304
rect 15284 4264 15285 4304
rect 15243 4255 15285 4264
rect 18507 4304 18549 4313
rect 18507 4264 18508 4304
rect 18548 4264 18549 4304
rect 18507 4255 18549 4264
rect 22347 4304 22389 4313
rect 22347 4264 22348 4304
rect 22388 4264 22389 4304
rect 22347 4255 22389 4264
rect 31179 4304 31221 4313
rect 31179 4264 31180 4304
rect 31220 4264 31221 4304
rect 31179 4255 31221 4264
rect 39339 4304 39381 4313
rect 39339 4264 39340 4304
rect 39380 4264 39381 4304
rect 39339 4255 39381 4264
rect 43851 4304 43893 4313
rect 43851 4264 43852 4304
rect 43892 4264 43893 4304
rect 43851 4255 43893 4264
rect 45147 4304 45189 4313
rect 45147 4264 45148 4304
rect 45188 4264 45189 4304
rect 45147 4255 45189 4264
rect 4779 4220 4821 4229
rect 7066 4220 7124 4221
rect 4779 4180 4780 4220
rect 4820 4180 4821 4220
rect 4779 4171 4821 4180
rect 6027 4211 6069 4220
rect 6027 4171 6028 4211
rect 6068 4171 6069 4211
rect 7066 4180 7075 4220
rect 7115 4180 7124 4220
rect 7066 4179 7124 4180
rect 7179 4220 7221 4229
rect 7179 4180 7180 4220
rect 7220 4180 7221 4220
rect 7179 4171 7221 4180
rect 7563 4220 7605 4229
rect 9483 4220 9525 4229
rect 7563 4180 7564 4220
rect 7604 4180 7605 4220
rect 7563 4171 7605 4180
rect 8139 4211 8181 4220
rect 8139 4171 8140 4211
rect 8180 4171 8181 4211
rect 6027 4162 6069 4171
rect 8139 4162 8181 4171
rect 8619 4211 8661 4220
rect 8619 4171 8620 4211
rect 8660 4171 8661 4211
rect 9483 4180 9484 4220
rect 9524 4180 9525 4220
rect 9483 4171 9525 4180
rect 9754 4220 9812 4221
rect 9754 4180 9763 4220
rect 9803 4180 9812 4220
rect 9754 4179 9812 4180
rect 12267 4220 12309 4229
rect 15364 4220 15422 4221
rect 12267 4180 12268 4220
rect 12308 4180 12309 4220
rect 12267 4171 12309 4180
rect 13515 4211 13557 4220
rect 13515 4171 13516 4211
rect 13556 4171 13557 4211
rect 15364 4180 15373 4220
rect 15413 4180 15422 4220
rect 15364 4179 15422 4180
rect 15627 4220 15669 4229
rect 15627 4180 15628 4220
rect 15668 4180 15669 4220
rect 15627 4171 15669 4180
rect 16875 4220 16917 4229
rect 19947 4220 19989 4229
rect 16875 4180 16876 4220
rect 16916 4180 16917 4220
rect 16875 4171 16917 4180
rect 18123 4211 18165 4220
rect 18123 4171 18124 4211
rect 18164 4171 18165 4211
rect 8619 4162 8661 4171
rect 13515 4162 13557 4171
rect 18123 4162 18165 4171
rect 18699 4211 18741 4220
rect 18699 4171 18700 4211
rect 18740 4171 18741 4211
rect 19947 4180 19948 4220
rect 19988 4180 19989 4220
rect 19947 4171 19989 4180
rect 20907 4220 20949 4229
rect 25611 4220 25653 4229
rect 27243 4220 27285 4229
rect 20907 4180 20908 4220
rect 20948 4180 20949 4220
rect 20907 4171 20949 4180
rect 22155 4211 22197 4220
rect 22155 4171 22156 4211
rect 22196 4171 22197 4211
rect 18699 4162 18741 4171
rect 22155 4162 22197 4171
rect 24363 4211 24405 4220
rect 24363 4171 24364 4211
rect 24404 4171 24405 4211
rect 25611 4180 25612 4220
rect 25652 4180 25653 4220
rect 25611 4171 25653 4180
rect 25995 4211 26037 4220
rect 25995 4171 25996 4211
rect 26036 4171 26037 4211
rect 27243 4180 27244 4220
rect 27284 4180 27285 4220
rect 27243 4171 27285 4180
rect 27627 4220 27669 4229
rect 29739 4220 29781 4229
rect 32602 4220 32660 4221
rect 27627 4180 27628 4220
rect 27668 4180 27669 4220
rect 27627 4171 27669 4180
rect 28875 4211 28917 4220
rect 28875 4171 28876 4211
rect 28916 4171 28917 4211
rect 29739 4180 29740 4220
rect 29780 4180 29781 4220
rect 29739 4171 29781 4180
rect 30987 4211 31029 4220
rect 30987 4171 30988 4211
rect 31028 4171 31029 4211
rect 32602 4180 32611 4220
rect 32651 4180 32660 4220
rect 32602 4179 32660 4180
rect 32715 4220 32757 4229
rect 32715 4180 32716 4220
rect 32756 4180 32757 4220
rect 32715 4171 32757 4180
rect 33092 4220 33134 4229
rect 37227 4220 37269 4229
rect 38907 4220 38949 4229
rect 33092 4180 33093 4220
rect 33133 4180 33134 4220
rect 33092 4171 33134 4180
rect 33675 4211 33717 4220
rect 33675 4171 33676 4211
rect 33716 4171 33717 4211
rect 24363 4162 24405 4171
rect 25995 4162 26037 4171
rect 28875 4162 28917 4171
rect 30987 4162 31029 4171
rect 33675 4162 33717 4171
rect 34155 4211 34197 4220
rect 34155 4171 34156 4211
rect 34196 4171 34197 4211
rect 37227 4180 37228 4220
rect 37268 4180 37269 4220
rect 37227 4171 37269 4180
rect 38475 4211 38517 4220
rect 38475 4171 38476 4211
rect 38516 4171 38517 4211
rect 38907 4180 38908 4220
rect 38948 4180 38949 4220
rect 38907 4171 38949 4180
rect 39226 4220 39284 4221
rect 41643 4220 41685 4229
rect 39226 4180 39235 4220
rect 39275 4180 39284 4220
rect 39226 4179 39284 4180
rect 40395 4211 40437 4220
rect 40395 4171 40396 4211
rect 40436 4171 40437 4211
rect 41643 4180 41644 4220
rect 41684 4180 41685 4220
rect 41643 4171 41685 4180
rect 43467 4220 43509 4229
rect 43467 4180 43468 4220
rect 43508 4180 43509 4220
rect 43467 4171 43509 4180
rect 34155 4162 34197 4171
rect 38475 4162 38517 4171
rect 40395 4162 40437 4171
rect 1227 4136 1269 4145
rect 1227 4096 1228 4136
rect 1268 4096 1269 4136
rect 1227 4087 1269 4096
rect 1467 4136 1509 4145
rect 1467 4096 1468 4136
rect 1508 4096 1509 4136
rect 1467 4087 1509 4096
rect 1611 4136 1653 4145
rect 1611 4096 1612 4136
rect 1652 4096 1653 4136
rect 1611 4087 1653 4096
rect 4107 4136 4149 4145
rect 4107 4096 4108 4136
rect 4148 4096 4149 4136
rect 4107 4087 4149 4096
rect 6411 4136 6453 4145
rect 6411 4096 6412 4136
rect 6452 4096 6453 4136
rect 6411 4087 6453 4096
rect 7659 4136 7701 4145
rect 7659 4096 7660 4136
rect 7700 4096 7701 4136
rect 7659 4087 7701 4096
rect 9003 4136 9045 4145
rect 9003 4096 9004 4136
rect 9044 4096 9045 4136
rect 9003 4087 9045 4096
rect 10203 4136 10245 4145
rect 10203 4096 10204 4136
rect 10244 4096 10245 4136
rect 10203 4087 10245 4096
rect 10347 4136 10389 4145
rect 10347 4096 10348 4136
rect 10388 4096 10389 4136
rect 10347 4087 10389 4096
rect 11019 4136 11061 4145
rect 11019 4096 11020 4136
rect 11060 4096 11061 4136
rect 11019 4087 11061 4096
rect 13947 4136 13989 4145
rect 13947 4096 13948 4136
rect 13988 4096 13989 4136
rect 13947 4087 13989 4096
rect 14187 4136 14229 4145
rect 14187 4096 14188 4136
rect 14228 4096 14229 4136
rect 14187 4087 14229 4096
rect 20139 4136 20181 4145
rect 20139 4096 20140 4136
rect 20180 4096 20181 4136
rect 20139 4087 20181 4096
rect 20523 4136 20565 4145
rect 20523 4096 20524 4136
rect 20564 4096 20565 4136
rect 20523 4087 20565 4096
rect 23787 4136 23829 4145
rect 23787 4096 23788 4136
rect 23828 4096 23829 4136
rect 23787 4087 23829 4096
rect 29451 4136 29493 4145
rect 29451 4096 29452 4136
rect 29492 4096 29493 4136
rect 29451 4087 29493 4096
rect 33195 4136 33237 4145
rect 33195 4096 33196 4136
rect 33236 4096 33237 4136
rect 33195 4087 33237 4096
rect 34731 4136 34773 4145
rect 34731 4096 34732 4136
rect 34772 4096 34773 4136
rect 34731 4087 34773 4096
rect 34923 4136 34965 4145
rect 34923 4096 34924 4136
rect 34964 4096 34965 4136
rect 34923 4087 34965 4096
rect 35979 4136 36021 4145
rect 35979 4096 35980 4136
rect 36020 4096 36021 4136
rect 35979 4087 36021 4096
rect 39771 4136 39813 4145
rect 39771 4096 39772 4136
rect 39812 4096 39813 4136
rect 39771 4087 39813 4096
rect 40011 4136 40053 4145
rect 40011 4096 40012 4136
rect 40052 4096 40053 4136
rect 40011 4087 40053 4096
rect 42027 4136 42069 4145
rect 42027 4096 42028 4136
rect 42068 4096 42069 4136
rect 42027 4087 42069 4096
rect 43179 4136 43221 4145
rect 43179 4096 43180 4136
rect 43220 4096 43221 4136
rect 43179 4087 43221 4096
rect 44523 4136 44565 4145
rect 44523 4096 44524 4136
rect 44564 4096 44565 4136
rect 44523 4087 44565 4096
rect 44907 4136 44949 4145
rect 44907 4096 44908 4136
rect 44948 4096 44949 4136
rect 44907 4087 44949 4096
rect 1851 4052 1893 4061
rect 1851 4012 1852 4052
rect 1892 4012 1893 4052
rect 1851 4003 1893 4012
rect 18315 4052 18357 4061
rect 18315 4012 18316 4052
rect 18356 4012 18357 4052
rect 18315 4003 18357 4012
rect 20379 4052 20421 4061
rect 20379 4012 20380 4052
rect 20420 4012 20421 4052
rect 20379 4003 20421 4012
rect 20763 4052 20805 4061
rect 20763 4012 20764 4052
rect 20804 4012 20805 4052
rect 20763 4003 20805 4012
rect 24171 4052 24213 4061
rect 24171 4012 24172 4052
rect 24212 4012 24213 4052
rect 24171 4003 24213 4012
rect 34491 4052 34533 4061
rect 34491 4012 34492 4052
rect 34532 4012 34533 4052
rect 34491 4003 34533 4012
rect 38667 4052 38709 4061
rect 38667 4012 38668 4052
rect 38708 4012 38709 4052
rect 38667 4003 38709 4012
rect 39627 4052 39669 4061
rect 39627 4012 39628 4052
rect 39668 4012 39669 4052
rect 39627 4003 39669 4012
rect 44763 4052 44805 4061
rect 44763 4012 44764 4052
rect 44804 4012 44805 4052
rect 44763 4003 44805 4012
rect 4347 3968 4389 3977
rect 4347 3928 4348 3968
rect 4388 3928 4389 3968
rect 4347 3919 4389 3928
rect 6651 3968 6693 3977
rect 6651 3928 6652 3968
rect 6692 3928 6693 3968
rect 6651 3919 6693 3928
rect 10587 3968 10629 3977
rect 10587 3928 10588 3968
rect 10628 3928 10629 3968
rect 10587 3919 10629 3928
rect 14955 3968 14997 3977
rect 14955 3928 14956 3968
rect 14996 3928 14997 3968
rect 14955 3919 14997 3928
rect 25803 3968 25845 3977
rect 25803 3928 25804 3968
rect 25844 3928 25845 3968
rect 25803 3919 25845 3928
rect 29067 3968 29109 3977
rect 29067 3928 29068 3968
rect 29108 3928 29109 3968
rect 29067 3919 29109 3928
rect 29211 3968 29253 3977
rect 29211 3928 29212 3968
rect 29252 3928 29253 3968
rect 29211 3919 29253 3928
rect 34378 3968 34436 3969
rect 34378 3928 34387 3968
rect 34427 3928 34436 3968
rect 34378 3927 34436 3928
rect 35163 3968 35205 3977
rect 35163 3928 35164 3968
rect 35204 3928 35205 3968
rect 35163 3919 35205 3928
rect 36219 3968 36261 3977
rect 36219 3928 36220 3968
rect 36260 3928 36261 3968
rect 36219 3919 36261 3928
rect 40203 3968 40245 3977
rect 40203 3928 40204 3968
rect 40244 3928 40245 3968
rect 40203 3919 40245 3928
rect 41787 3968 41829 3977
rect 41787 3928 41788 3968
rect 41828 3928 41829 3968
rect 41787 3919 41829 3928
rect 1152 3800 45216 3824
rect 1152 3760 3688 3800
rect 3728 3760 3770 3800
rect 3810 3760 3852 3800
rect 3892 3760 3934 3800
rect 3974 3760 4016 3800
rect 4056 3760 18808 3800
rect 18848 3760 18890 3800
rect 18930 3760 18972 3800
rect 19012 3760 19054 3800
rect 19094 3760 19136 3800
rect 19176 3760 33928 3800
rect 33968 3760 34010 3800
rect 34050 3760 34092 3800
rect 34132 3760 34174 3800
rect 34214 3760 34256 3800
rect 34296 3760 45216 3800
rect 1152 3736 45216 3760
rect 14619 3632 14661 3641
rect 14619 3592 14620 3632
rect 14660 3592 14661 3632
rect 14619 3583 14661 3592
rect 43995 3632 44037 3641
rect 43995 3592 43996 3632
rect 44036 3592 44037 3632
rect 43995 3583 44037 3592
rect 45147 3632 45189 3641
rect 45147 3592 45148 3632
rect 45188 3592 45189 3632
rect 45147 3583 45189 3592
rect 1467 3548 1509 3557
rect 1467 3508 1468 3548
rect 1508 3508 1509 3548
rect 1467 3499 1509 3508
rect 1851 3548 1893 3557
rect 1851 3508 1852 3548
rect 1892 3508 1893 3548
rect 1851 3499 1893 3508
rect 5355 3548 5397 3557
rect 5355 3508 5356 3548
rect 5396 3508 5397 3548
rect 5355 3499 5397 3508
rect 8139 3548 8181 3557
rect 8139 3508 8140 3548
rect 8180 3508 8181 3548
rect 8139 3499 8181 3508
rect 8571 3548 8613 3557
rect 8571 3508 8572 3548
rect 8612 3508 8613 3548
rect 8571 3499 8613 3508
rect 13803 3548 13845 3557
rect 13803 3508 13804 3548
rect 13844 3508 13845 3548
rect 13803 3499 13845 3508
rect 14235 3548 14277 3557
rect 14235 3508 14236 3548
rect 14276 3508 14277 3548
rect 14235 3499 14277 3508
rect 18987 3548 19029 3557
rect 18987 3508 18988 3548
rect 19028 3508 19029 3548
rect 18987 3499 19029 3508
rect 24651 3548 24693 3557
rect 24651 3508 24652 3548
rect 24692 3508 24693 3548
rect 24651 3499 24693 3508
rect 29547 3548 29589 3557
rect 29547 3508 29548 3548
rect 29588 3508 29589 3548
rect 29547 3499 29589 3508
rect 31947 3548 31989 3557
rect 31947 3508 31948 3548
rect 31988 3508 31989 3548
rect 31947 3499 31989 3508
rect 33483 3548 33525 3557
rect 33483 3508 33484 3548
rect 33524 3508 33525 3548
rect 33483 3499 33525 3508
rect 1227 3464 1269 3473
rect 1227 3424 1228 3464
rect 1268 3424 1269 3464
rect 1227 3415 1269 3424
rect 1611 3464 1653 3473
rect 1611 3424 1612 3464
rect 1652 3424 1653 3464
rect 1611 3415 1653 3424
rect 8331 3464 8373 3473
rect 8331 3424 8332 3464
rect 8372 3424 8373 3464
rect 8331 3415 8373 3424
rect 8715 3464 8757 3473
rect 8715 3424 8716 3464
rect 8756 3424 8757 3464
rect 8715 3415 8757 3424
rect 13995 3464 14037 3473
rect 13995 3424 13996 3464
rect 14036 3424 14037 3464
rect 13995 3415 14037 3424
rect 14859 3464 14901 3473
rect 14859 3424 14860 3464
rect 14900 3424 14901 3464
rect 14859 3415 14901 3424
rect 15627 3464 15669 3473
rect 15627 3424 15628 3464
rect 15668 3424 15669 3464
rect 15627 3415 15669 3424
rect 18027 3464 18069 3473
rect 18027 3424 18028 3464
rect 18068 3424 18069 3464
rect 16683 3413 16725 3422
rect 18027 3415 18069 3424
rect 19371 3464 19413 3473
rect 19371 3424 19372 3464
rect 19412 3424 19413 3464
rect 19371 3415 19413 3424
rect 21003 3464 21045 3473
rect 21003 3424 21004 3464
rect 21044 3424 21045 3464
rect 21003 3415 21045 3424
rect 24795 3464 24837 3473
rect 24795 3424 24796 3464
rect 24836 3424 24837 3464
rect 24795 3415 24837 3424
rect 25035 3464 25077 3473
rect 25035 3424 25036 3464
rect 25076 3424 25077 3464
rect 25035 3415 25077 3424
rect 25707 3464 25749 3473
rect 25707 3424 25708 3464
rect 25748 3424 25749 3464
rect 25707 3415 25749 3424
rect 29787 3464 29829 3473
rect 29787 3424 29788 3464
rect 29828 3424 29829 3464
rect 29787 3415 29829 3424
rect 30027 3464 30069 3473
rect 30027 3424 30028 3464
rect 30068 3424 30069 3464
rect 30027 3415 30069 3424
rect 33867 3464 33909 3473
rect 33867 3424 33868 3464
rect 33908 3424 33909 3464
rect 33867 3415 33909 3424
rect 38571 3464 38613 3473
rect 38571 3424 38572 3464
rect 38612 3424 38613 3464
rect 38571 3415 38613 3424
rect 44235 3464 44277 3473
rect 44235 3424 44236 3464
rect 44276 3424 44277 3464
rect 44235 3415 44277 3424
rect 44619 3464 44661 3473
rect 44619 3424 44620 3464
rect 44660 3424 44661 3464
rect 44619 3415 44661 3424
rect 44907 3464 44949 3473
rect 44907 3424 44908 3464
rect 44948 3424 44949 3464
rect 44907 3415 44949 3424
rect 3915 3380 3957 3389
rect 3915 3340 3916 3380
rect 3956 3340 3957 3380
rect 3915 3331 3957 3340
rect 5155 3380 5213 3381
rect 5155 3340 5164 3380
rect 5204 3340 5213 3380
rect 5155 3339 5213 3340
rect 7467 3380 7509 3389
rect 7467 3340 7468 3380
rect 7508 3340 7509 3380
rect 7467 3331 7509 3340
rect 7738 3380 7796 3381
rect 7738 3340 7747 3380
rect 7787 3340 7796 3380
rect 7738 3339 7796 3340
rect 11403 3380 11445 3389
rect 11403 3340 11404 3380
rect 11444 3340 11445 3380
rect 11403 3331 11445 3340
rect 12643 3380 12701 3381
rect 12643 3340 12652 3380
rect 12692 3340 12701 3380
rect 12643 3339 12701 3340
rect 13131 3380 13173 3389
rect 13131 3340 13132 3380
rect 13172 3340 13173 3380
rect 13131 3331 13173 3340
rect 13402 3380 13460 3381
rect 13402 3340 13411 3380
rect 13451 3340 13460 3380
rect 13402 3339 13460 3340
rect 15130 3380 15188 3381
rect 15130 3340 15139 3380
rect 15179 3340 15188 3380
rect 15130 3339 15188 3340
rect 15243 3380 15285 3389
rect 15243 3340 15244 3380
rect 15284 3340 15285 3380
rect 15243 3331 15285 3340
rect 15723 3380 15765 3389
rect 15723 3340 15724 3380
rect 15764 3340 15765 3380
rect 15723 3331 15765 3340
rect 16195 3380 16253 3381
rect 16195 3340 16204 3380
rect 16244 3340 16253 3380
rect 16683 3373 16684 3413
rect 16724 3373 16725 3413
rect 16683 3364 16725 3373
rect 18315 3380 18357 3389
rect 16195 3339 16253 3340
rect 18315 3340 18316 3380
rect 18356 3340 18357 3380
rect 18315 3331 18357 3340
rect 18586 3380 18644 3381
rect 18586 3340 18595 3380
rect 18635 3340 18644 3380
rect 18586 3339 18644 3340
rect 23979 3380 24021 3389
rect 23979 3340 23980 3380
rect 24020 3340 24021 3380
rect 23979 3331 24021 3340
rect 24250 3380 24308 3381
rect 24250 3340 24259 3380
rect 24299 3340 24308 3380
rect 24250 3339 24308 3340
rect 26379 3380 26421 3389
rect 26379 3340 26380 3380
rect 26420 3340 26421 3380
rect 26379 3331 26421 3340
rect 27619 3380 27677 3381
rect 27619 3340 27628 3380
rect 27668 3340 27677 3380
rect 27619 3339 27677 3340
rect 28875 3380 28917 3389
rect 28875 3340 28876 3380
rect 28916 3340 28917 3380
rect 28875 3331 28917 3340
rect 29146 3380 29204 3381
rect 29146 3340 29155 3380
rect 29195 3340 29204 3380
rect 29146 3339 29204 3340
rect 30507 3380 30549 3389
rect 30507 3340 30508 3380
rect 30548 3340 30549 3380
rect 30507 3331 30549 3340
rect 31747 3380 31805 3381
rect 31747 3340 31756 3380
rect 31796 3340 31805 3380
rect 31747 3339 31805 3340
rect 32811 3380 32853 3389
rect 32811 3340 32812 3380
rect 32852 3340 32853 3380
rect 32811 3331 32853 3340
rect 33082 3380 33140 3381
rect 33082 3340 33091 3380
rect 33131 3340 33140 3380
rect 33082 3339 33140 3340
rect 36171 3380 36213 3389
rect 36171 3340 36172 3380
rect 36212 3340 36213 3380
rect 36171 3331 36213 3340
rect 37415 3380 37473 3381
rect 37415 3340 37424 3380
rect 37464 3340 37473 3380
rect 37415 3339 37473 3340
rect 38074 3380 38132 3381
rect 38074 3340 38083 3380
rect 38123 3340 38132 3380
rect 38074 3339 38132 3340
rect 38187 3380 38229 3389
rect 38187 3340 38188 3380
rect 38228 3340 38229 3380
rect 38187 3331 38229 3340
rect 38667 3380 38709 3389
rect 38667 3340 38668 3380
rect 38708 3340 38709 3380
rect 38667 3331 38709 3340
rect 39139 3380 39197 3381
rect 39139 3340 39148 3380
rect 39188 3340 39197 3380
rect 39139 3339 39197 3340
rect 39658 3380 39716 3381
rect 39658 3340 39667 3380
rect 39707 3340 39716 3380
rect 39658 3339 39716 3340
rect 41355 3380 41397 3389
rect 41355 3340 41356 3380
rect 41396 3340 41397 3380
rect 41355 3331 41397 3340
rect 43755 3380 43797 3389
rect 43755 3340 43756 3380
rect 43796 3340 43797 3380
rect 43755 3331 43797 3340
rect 7851 3296 7893 3305
rect 7851 3256 7852 3296
rect 7892 3256 7893 3296
rect 7851 3247 7893 3256
rect 12843 3296 12885 3305
rect 12843 3256 12844 3296
rect 12884 3256 12885 3296
rect 12843 3247 12885 3256
rect 13515 3296 13557 3305
rect 13515 3256 13516 3296
rect 13556 3256 13557 3296
rect 13515 3247 13557 3256
rect 18699 3296 18741 3305
rect 18699 3256 18700 3296
rect 18740 3256 18741 3296
rect 18699 3247 18741 3256
rect 19131 3296 19173 3305
rect 19131 3256 19132 3296
rect 19172 3256 19173 3296
rect 19131 3247 19173 3256
rect 24363 3296 24405 3305
rect 24363 3256 24364 3296
rect 24404 3256 24405 3296
rect 24363 3247 24405 3256
rect 29259 3296 29301 3305
rect 29259 3256 29260 3296
rect 29300 3256 29301 3296
rect 29259 3247 29301 3256
rect 33179 3296 33221 3305
rect 33179 3256 33180 3296
rect 33220 3256 33221 3296
rect 33179 3247 33221 3256
rect 33627 3296 33669 3305
rect 33627 3256 33628 3296
rect 33668 3256 33669 3296
rect 33627 3247 33669 3256
rect 37611 3296 37653 3305
rect 37611 3256 37612 3296
rect 37652 3256 37653 3296
rect 37611 3247 37653 3256
rect 44379 3296 44421 3305
rect 44379 3256 44380 3296
rect 44420 3256 44421 3296
rect 44379 3247 44421 3256
rect 8955 3212 8997 3221
rect 8955 3172 8956 3212
rect 8996 3172 8997 3212
rect 8955 3163 8997 3172
rect 16875 3212 16917 3221
rect 16875 3172 16876 3212
rect 16916 3172 16917 3212
rect 16875 3163 16917 3172
rect 17787 3212 17829 3221
rect 17787 3172 17788 3212
rect 17828 3172 17829 3212
rect 17787 3163 17829 3172
rect 21243 3212 21285 3221
rect 21243 3172 21244 3212
rect 21284 3172 21285 3212
rect 21243 3163 21285 3172
rect 25467 3212 25509 3221
rect 25467 3172 25468 3212
rect 25508 3172 25509 3212
rect 25467 3163 25509 3172
rect 27819 3212 27861 3221
rect 27819 3172 27820 3212
rect 27860 3172 27861 3212
rect 27819 3163 27861 3172
rect 39819 3212 39861 3221
rect 39819 3172 39820 3212
rect 39860 3172 39861 3212
rect 39819 3163 39861 3172
rect 41626 3212 41684 3213
rect 41626 3172 41635 3212
rect 41675 3172 41684 3212
rect 41626 3171 41684 3172
rect 41914 3212 41972 3213
rect 41914 3172 41923 3212
rect 41963 3172 41972 3212
rect 41914 3171 41972 3172
rect 42202 3212 42260 3213
rect 42202 3172 42211 3212
rect 42251 3172 42260 3212
rect 42202 3171 42260 3172
rect 42490 3212 42548 3213
rect 42490 3172 42499 3212
rect 42539 3172 42548 3212
rect 42490 3171 42548 3172
rect 42778 3212 42836 3213
rect 42778 3172 42787 3212
rect 42827 3172 42836 3212
rect 42778 3171 42836 3172
rect 43066 3212 43124 3213
rect 43066 3172 43075 3212
rect 43115 3172 43124 3212
rect 43066 3171 43124 3172
rect 43354 3212 43412 3213
rect 43354 3172 43363 3212
rect 43403 3172 43412 3212
rect 43354 3171 43412 3172
rect 1152 3044 45216 3068
rect 1152 3004 4928 3044
rect 4968 3004 5010 3044
rect 5050 3004 5092 3044
rect 5132 3004 5174 3044
rect 5214 3004 5256 3044
rect 5296 3004 20048 3044
rect 20088 3004 20130 3044
rect 20170 3004 20212 3044
rect 20252 3004 20294 3044
rect 20334 3004 20376 3044
rect 20416 3004 35168 3044
rect 35208 3004 35250 3044
rect 35290 3004 35332 3044
rect 35372 3004 35414 3044
rect 35454 3004 35496 3044
rect 35536 3004 45216 3044
rect 1152 2980 45216 3004
rect 5595 2876 5637 2885
rect 5595 2836 5596 2876
rect 5636 2836 5637 2876
rect 5595 2827 5637 2836
rect 7179 2876 7221 2885
rect 7179 2836 7180 2876
rect 7220 2836 7221 2876
rect 7179 2827 7221 2836
rect 9003 2876 9045 2885
rect 9003 2836 9004 2876
rect 9044 2836 9045 2876
rect 9003 2827 9045 2836
rect 9627 2876 9669 2885
rect 9627 2836 9628 2876
rect 9668 2836 9669 2876
rect 9627 2827 9669 2836
rect 11211 2876 11253 2885
rect 11211 2836 11212 2876
rect 11252 2836 11253 2876
rect 11211 2827 11253 2836
rect 15435 2876 15477 2885
rect 15435 2836 15436 2876
rect 15476 2836 15477 2876
rect 15435 2827 15477 2836
rect 20907 2876 20949 2885
rect 20907 2836 20908 2876
rect 20948 2836 20949 2876
rect 20907 2827 20949 2836
rect 24843 2876 24885 2885
rect 24843 2836 24844 2876
rect 24884 2836 24885 2876
rect 24843 2827 24885 2836
rect 27531 2876 27573 2885
rect 27531 2836 27532 2876
rect 27572 2836 27573 2876
rect 27531 2827 27573 2836
rect 30027 2876 30069 2885
rect 30027 2836 30028 2876
rect 30068 2836 30069 2876
rect 30027 2827 30069 2836
rect 34059 2876 34101 2885
rect 34059 2836 34060 2876
rect 34100 2836 34101 2876
rect 34059 2827 34101 2836
rect 40762 2876 40820 2877
rect 40762 2836 40771 2876
rect 40811 2836 40820 2876
rect 40762 2835 40820 2836
rect 41050 2876 41108 2877
rect 41050 2836 41059 2876
rect 41099 2836 41108 2876
rect 41050 2835 41108 2836
rect 41307 2876 41349 2885
rect 41307 2836 41308 2876
rect 41348 2836 41349 2876
rect 41307 2827 41349 2836
rect 41691 2876 41733 2885
rect 41691 2836 41692 2876
rect 41732 2836 41733 2876
rect 41691 2827 41733 2836
rect 42459 2876 42501 2885
rect 42459 2836 42460 2876
rect 42500 2836 42501 2876
rect 42459 2827 42501 2836
rect 43066 2876 43124 2877
rect 43066 2836 43075 2876
rect 43115 2836 43124 2876
rect 43066 2835 43124 2836
rect 45147 2876 45189 2885
rect 45147 2836 45148 2876
rect 45188 2836 45189 2876
rect 45147 2827 45189 2836
rect 1467 2792 1509 2801
rect 1467 2752 1468 2792
rect 1508 2752 1509 2792
rect 1467 2743 1509 2752
rect 18603 2792 18645 2801
rect 18603 2752 18604 2792
rect 18644 2752 18645 2792
rect 18603 2743 18645 2752
rect 22635 2792 22677 2801
rect 22635 2752 22636 2792
rect 22676 2752 22677 2792
rect 22635 2743 22677 2752
rect 24987 2792 25029 2801
rect 24987 2752 24988 2792
rect 25028 2752 25029 2792
rect 24987 2743 25029 2752
rect 30555 2792 30597 2801
rect 30555 2752 30556 2792
rect 30596 2752 30597 2792
rect 30555 2743 30597 2752
rect 30987 2792 31029 2801
rect 30987 2752 30988 2792
rect 31028 2752 31029 2792
rect 30987 2743 31029 2752
rect 35739 2792 35781 2801
rect 35739 2752 35740 2792
rect 35780 2752 35781 2792
rect 35739 2743 35781 2752
rect 38091 2792 38133 2801
rect 38091 2752 38092 2792
rect 38132 2752 38133 2792
rect 38091 2743 38133 2752
rect 38763 2792 38805 2801
rect 38763 2752 38764 2792
rect 38804 2752 38805 2792
rect 38763 2743 38805 2752
rect 44763 2792 44805 2801
rect 44763 2752 44764 2792
rect 44804 2752 44805 2792
rect 44763 2743 44805 2752
rect 5739 2708 5781 2717
rect 7563 2708 7605 2717
rect 9771 2708 9813 2717
rect 11403 2708 11445 2717
rect 13323 2708 13365 2717
rect 5739 2668 5740 2708
rect 5780 2668 5781 2708
rect 5739 2659 5781 2668
rect 6987 2699 7029 2708
rect 6987 2659 6988 2699
rect 7028 2659 7029 2699
rect 7563 2668 7564 2708
rect 7604 2668 7605 2708
rect 7563 2659 7605 2668
rect 8811 2699 8853 2708
rect 8811 2659 8812 2699
rect 8852 2659 8853 2699
rect 9771 2668 9772 2708
rect 9812 2668 9813 2708
rect 9771 2659 9813 2668
rect 11019 2699 11061 2708
rect 11019 2659 11020 2699
rect 11060 2659 11061 2699
rect 11403 2668 11404 2708
rect 11444 2668 11445 2708
rect 11403 2659 11445 2668
rect 12651 2699 12693 2708
rect 12651 2659 12652 2699
rect 12692 2659 12693 2699
rect 13323 2668 13324 2708
rect 13364 2668 13365 2708
rect 13323 2659 13365 2668
rect 13444 2708 13502 2709
rect 13444 2668 13453 2708
rect 13493 2668 13502 2708
rect 13444 2667 13502 2668
rect 13707 2708 13749 2717
rect 13707 2668 13708 2708
rect 13748 2668 13749 2708
rect 13707 2659 13749 2668
rect 13995 2708 14037 2717
rect 15706 2708 15764 2709
rect 13995 2668 13996 2708
rect 14036 2668 14037 2708
rect 13995 2659 14037 2668
rect 15243 2699 15285 2708
rect 15243 2659 15244 2699
rect 15284 2659 15285 2699
rect 15706 2668 15715 2708
rect 15755 2668 15764 2708
rect 15706 2667 15764 2668
rect 15819 2708 15861 2717
rect 15819 2668 15820 2708
rect 15860 2668 15861 2708
rect 15819 2659 15861 2668
rect 16203 2708 16245 2717
rect 18219 2708 18261 2717
rect 16203 2668 16204 2708
rect 16244 2668 16245 2708
rect 16203 2659 16245 2668
rect 16779 2699 16821 2708
rect 16779 2659 16780 2699
rect 16820 2659 16821 2699
rect 6987 2650 7029 2659
rect 8811 2650 8853 2659
rect 11019 2650 11061 2659
rect 12651 2650 12693 2659
rect 15243 2650 15285 2659
rect 16779 2650 16821 2659
rect 17259 2699 17301 2708
rect 17259 2659 17260 2699
rect 17300 2659 17301 2699
rect 18219 2668 18220 2708
rect 18260 2668 18261 2708
rect 18219 2659 18261 2668
rect 18490 2708 18548 2709
rect 18490 2668 18499 2708
rect 18539 2668 18548 2708
rect 18490 2667 18548 2668
rect 19162 2708 19220 2709
rect 19162 2668 19171 2708
rect 19211 2668 19220 2708
rect 19162 2667 19220 2668
rect 19275 2708 19317 2717
rect 19275 2668 19276 2708
rect 19316 2668 19317 2708
rect 19275 2659 19317 2668
rect 19659 2708 19701 2717
rect 21195 2708 21237 2717
rect 23098 2708 23156 2709
rect 19659 2668 19660 2708
rect 19700 2668 19701 2708
rect 19659 2659 19701 2668
rect 20235 2699 20277 2708
rect 20235 2659 20236 2699
rect 20276 2659 20277 2699
rect 17259 2650 17301 2659
rect 20235 2650 20277 2659
rect 20715 2699 20757 2708
rect 20715 2659 20716 2699
rect 20756 2659 20757 2699
rect 21195 2668 21196 2708
rect 21236 2668 21237 2708
rect 21195 2659 21237 2668
rect 22443 2699 22485 2708
rect 22443 2659 22444 2699
rect 22484 2659 22485 2699
rect 23098 2668 23107 2708
rect 23147 2668 23156 2708
rect 23098 2667 23156 2668
rect 23211 2708 23253 2717
rect 23211 2668 23212 2708
rect 23252 2668 23253 2708
rect 23211 2659 23253 2668
rect 23595 2708 23637 2717
rect 25323 2708 25365 2717
rect 23595 2668 23596 2708
rect 23636 2668 23637 2708
rect 23595 2659 23637 2668
rect 24171 2699 24213 2708
rect 24171 2659 24172 2699
rect 24212 2659 24213 2699
rect 20715 2650 20757 2659
rect 22443 2650 22485 2659
rect 24171 2650 24213 2659
rect 24651 2699 24693 2708
rect 24651 2659 24652 2699
rect 24692 2659 24693 2699
rect 25323 2668 25324 2708
rect 25364 2668 25365 2708
rect 25323 2659 25365 2668
rect 25444 2708 25502 2709
rect 25444 2668 25453 2708
rect 25493 2668 25502 2708
rect 25444 2667 25502 2668
rect 25707 2708 25749 2717
rect 25707 2668 25708 2708
rect 25748 2668 25749 2708
rect 25707 2659 25749 2668
rect 26091 2708 26133 2717
rect 28282 2708 28340 2709
rect 26091 2668 26092 2708
rect 26132 2668 26133 2708
rect 26091 2659 26133 2668
rect 27339 2699 27381 2708
rect 27339 2659 27340 2699
rect 27380 2659 27381 2699
rect 28282 2668 28291 2708
rect 28331 2668 28340 2708
rect 28282 2667 28340 2668
rect 28395 2708 28437 2717
rect 28395 2668 28396 2708
rect 28436 2668 28437 2708
rect 28395 2659 28437 2668
rect 28779 2708 28821 2717
rect 32427 2708 32469 2717
rect 28779 2668 28780 2708
rect 28820 2668 28821 2708
rect 28779 2659 28821 2668
rect 29355 2699 29397 2708
rect 29355 2659 29356 2699
rect 29396 2659 29397 2699
rect 24651 2650 24693 2659
rect 27339 2650 27381 2659
rect 29355 2650 29397 2659
rect 29835 2699 29877 2708
rect 29835 2659 29836 2699
rect 29876 2659 29877 2699
rect 29835 2650 29877 2659
rect 31179 2699 31221 2708
rect 31179 2659 31180 2699
rect 31220 2659 31221 2699
rect 32427 2668 32428 2708
rect 32468 2668 32469 2708
rect 32427 2659 32469 2668
rect 32619 2708 32661 2717
rect 34923 2708 34965 2717
rect 32619 2668 32620 2708
rect 32660 2668 32661 2708
rect 32619 2659 32661 2668
rect 33867 2699 33909 2708
rect 33867 2659 33868 2699
rect 33908 2659 33909 2699
rect 34923 2668 34924 2708
rect 34964 2668 34965 2708
rect 34923 2659 34965 2668
rect 35170 2708 35228 2709
rect 35170 2668 35179 2708
rect 35219 2668 35228 2708
rect 35170 2667 35228 2668
rect 35290 2708 35348 2709
rect 35290 2668 35299 2708
rect 35339 2668 35348 2708
rect 35290 2667 35348 2668
rect 36651 2708 36693 2717
rect 38379 2708 38421 2717
rect 36651 2668 36652 2708
rect 36692 2668 36693 2708
rect 36651 2659 36693 2668
rect 37899 2699 37941 2708
rect 37899 2659 37900 2699
rect 37940 2659 37941 2699
rect 38379 2668 38380 2708
rect 38420 2668 38421 2708
rect 38379 2659 38421 2668
rect 38650 2708 38708 2709
rect 38650 2668 38659 2708
rect 38699 2668 38708 2708
rect 38650 2667 38708 2668
rect 31179 2650 31221 2659
rect 33867 2650 33909 2659
rect 37899 2650 37941 2659
rect 1227 2624 1269 2633
rect 1227 2584 1228 2624
rect 1268 2584 1269 2624
rect 1227 2575 1269 2584
rect 1611 2624 1653 2633
rect 1611 2584 1612 2624
rect 1652 2584 1653 2624
rect 1611 2575 1653 2584
rect 1995 2624 2037 2633
rect 1995 2584 1996 2624
rect 2036 2584 2037 2624
rect 1995 2575 2037 2584
rect 5355 2624 5397 2633
rect 5355 2584 5356 2624
rect 5396 2584 5397 2624
rect 5355 2575 5397 2584
rect 9387 2624 9429 2633
rect 9387 2584 9388 2624
rect 9428 2584 9429 2624
rect 9387 2575 9429 2584
rect 16299 2624 16341 2633
rect 16299 2584 16300 2624
rect 16340 2584 16341 2624
rect 16299 2575 16341 2584
rect 17739 2624 17781 2633
rect 17739 2584 17740 2624
rect 17780 2584 17781 2624
rect 17739 2575 17781 2584
rect 19755 2624 19797 2633
rect 19755 2584 19756 2624
rect 19796 2584 19797 2624
rect 19755 2575 19797 2584
rect 23691 2624 23733 2633
rect 23691 2584 23692 2624
rect 23732 2584 23733 2624
rect 23691 2575 23733 2584
rect 27915 2624 27957 2633
rect 27915 2584 27916 2624
rect 27956 2584 27957 2624
rect 27915 2575 27957 2584
rect 28875 2624 28917 2633
rect 28875 2584 28876 2624
rect 28916 2584 28917 2624
rect 28875 2575 28917 2584
rect 30411 2624 30453 2633
rect 30411 2584 30412 2624
rect 30452 2584 30453 2624
rect 30411 2575 30453 2584
rect 30795 2624 30837 2633
rect 30795 2584 30796 2624
rect 30836 2584 30837 2624
rect 30795 2575 30837 2584
rect 35979 2624 36021 2633
rect 35979 2584 35980 2624
rect 36020 2584 36021 2624
rect 35979 2575 36021 2584
rect 36267 2624 36309 2633
rect 36267 2584 36268 2624
rect 36308 2584 36309 2624
rect 36267 2575 36309 2584
rect 39099 2624 39141 2633
rect 39099 2584 39100 2624
rect 39140 2584 39141 2624
rect 39099 2575 39141 2584
rect 39435 2624 39477 2633
rect 39435 2584 39436 2624
rect 39476 2584 39477 2624
rect 39435 2575 39477 2584
rect 41547 2624 41589 2633
rect 41547 2584 41548 2624
rect 41588 2584 41589 2624
rect 41547 2575 41589 2584
rect 41931 2624 41973 2633
rect 41931 2584 41932 2624
rect 41972 2584 41973 2624
rect 41931 2575 41973 2584
rect 42075 2624 42117 2633
rect 42075 2584 42076 2624
rect 42116 2584 42117 2624
rect 42075 2575 42117 2584
rect 42315 2624 42357 2633
rect 42315 2584 42316 2624
rect 42356 2584 42357 2624
rect 42315 2575 42357 2584
rect 42699 2624 42741 2633
rect 42699 2584 42700 2624
rect 42740 2584 42741 2624
rect 42699 2575 42741 2584
rect 43083 2624 43125 2633
rect 43083 2584 43084 2624
rect 43124 2584 43125 2624
rect 43083 2575 43125 2584
rect 43371 2624 43413 2633
rect 43371 2584 43372 2624
rect 43412 2584 43413 2624
rect 43371 2575 43413 2584
rect 43755 2624 43797 2633
rect 43755 2584 43756 2624
rect 43796 2584 43797 2624
rect 43755 2575 43797 2584
rect 44331 2624 44373 2633
rect 44331 2584 44332 2624
rect 44372 2584 44373 2624
rect 44331 2575 44373 2584
rect 44523 2624 44565 2633
rect 44523 2584 44524 2624
rect 44564 2584 44565 2624
rect 44523 2575 44565 2584
rect 44907 2624 44949 2633
rect 44907 2584 44908 2624
rect 44948 2584 44949 2624
rect 44907 2575 44949 2584
rect 2235 2540 2277 2549
rect 2235 2500 2236 2540
rect 2276 2500 2277 2540
rect 2235 2491 2277 2500
rect 27675 2540 27717 2549
rect 27675 2500 27676 2540
rect 27716 2500 27717 2540
rect 27675 2491 27717 2500
rect 35595 2540 35637 2549
rect 35595 2500 35596 2540
rect 35636 2500 35637 2540
rect 35595 2491 35637 2500
rect 43995 2540 44037 2549
rect 43995 2500 43996 2540
rect 44036 2500 44037 2540
rect 43995 2491 44037 2500
rect 1851 2456 1893 2465
rect 1851 2416 1852 2456
rect 1892 2416 1893 2456
rect 1851 2407 1893 2416
rect 12843 2456 12885 2465
rect 12843 2416 12844 2456
rect 12884 2416 12885 2456
rect 12843 2407 12885 2416
rect 13035 2456 13077 2465
rect 13035 2416 13036 2456
rect 13076 2416 13077 2456
rect 13035 2407 13077 2416
rect 17482 2456 17540 2457
rect 17482 2416 17491 2456
rect 17531 2416 17540 2456
rect 17482 2415 17540 2416
rect 17979 2456 18021 2465
rect 17979 2416 17980 2456
rect 18020 2416 18021 2456
rect 17979 2407 18021 2416
rect 18891 2456 18933 2465
rect 18891 2416 18892 2456
rect 18932 2416 18933 2456
rect 18891 2407 18933 2416
rect 30171 2456 30213 2465
rect 30171 2416 30172 2456
rect 30212 2416 30213 2456
rect 30171 2407 30213 2416
rect 36507 2456 36549 2465
rect 36507 2416 36508 2456
rect 36548 2416 36549 2456
rect 36507 2407 36549 2416
rect 39195 2456 39237 2465
rect 39195 2416 39196 2456
rect 39236 2416 39237 2456
rect 39195 2407 39237 2416
rect 43611 2456 43653 2465
rect 43611 2416 43612 2456
rect 43652 2416 43653 2456
rect 43611 2407 43653 2416
rect 44091 2456 44133 2465
rect 44091 2416 44092 2456
rect 44132 2416 44133 2456
rect 44091 2407 44133 2416
rect 1152 2288 45216 2312
rect 1152 2248 3688 2288
rect 3728 2248 3770 2288
rect 3810 2248 3852 2288
rect 3892 2248 3934 2288
rect 3974 2248 4016 2288
rect 4056 2248 18808 2288
rect 18848 2248 18890 2288
rect 18930 2248 18972 2288
rect 19012 2248 19054 2288
rect 19094 2248 19136 2288
rect 19176 2248 33928 2288
rect 33968 2248 34010 2288
rect 34050 2248 34092 2288
rect 34132 2248 34174 2288
rect 34214 2248 34256 2288
rect 34296 2248 45216 2288
rect 1152 2224 45216 2248
rect 1851 2120 1893 2129
rect 1851 2080 1852 2120
rect 1892 2080 1893 2120
rect 1851 2071 1893 2080
rect 2619 2120 2661 2129
rect 2619 2080 2620 2120
rect 2660 2080 2661 2120
rect 2619 2071 2661 2080
rect 4251 2120 4293 2129
rect 4251 2080 4252 2120
rect 4292 2080 4293 2120
rect 4251 2071 4293 2080
rect 5979 2120 6021 2129
rect 5979 2080 5980 2120
rect 6020 2080 6021 2120
rect 5979 2071 6021 2080
rect 8763 2120 8805 2129
rect 8763 2080 8764 2120
rect 8804 2080 8805 2120
rect 8763 2071 8805 2080
rect 9147 2120 9189 2129
rect 9147 2080 9148 2120
rect 9188 2080 9189 2120
rect 9147 2071 9189 2080
rect 10731 2120 10773 2129
rect 10731 2080 10732 2120
rect 10772 2080 10773 2120
rect 10731 2071 10773 2080
rect 13947 2120 13989 2129
rect 13947 2080 13948 2120
rect 13988 2080 13989 2120
rect 13947 2071 13989 2080
rect 16539 2120 16581 2129
rect 16539 2080 16540 2120
rect 16580 2080 16581 2120
rect 16539 2071 16581 2080
rect 16971 2120 17013 2129
rect 16971 2080 16972 2120
rect 17012 2080 17013 2120
rect 16971 2071 17013 2080
rect 20619 2120 20661 2129
rect 20619 2080 20620 2120
rect 20660 2080 20661 2120
rect 20619 2071 20661 2080
rect 34251 2120 34293 2129
rect 34251 2080 34252 2120
rect 34292 2080 34293 2120
rect 34251 2071 34293 2080
rect 35163 2120 35205 2129
rect 35163 2080 35164 2120
rect 35204 2080 35205 2120
rect 35163 2071 35205 2080
rect 36987 2120 37029 2129
rect 36987 2080 36988 2120
rect 37028 2080 37029 2120
rect 36987 2071 37029 2080
rect 39003 2120 39045 2129
rect 39003 2080 39004 2120
rect 39044 2080 39045 2120
rect 39003 2071 39045 2080
rect 40443 2120 40485 2129
rect 40443 2080 40444 2120
rect 40484 2080 40485 2120
rect 40443 2071 40485 2080
rect 41883 2120 41925 2129
rect 41883 2080 41884 2120
rect 41924 2080 41925 2120
rect 41883 2071 41925 2080
rect 42843 2120 42885 2129
rect 42843 2080 42844 2120
rect 42884 2080 42885 2120
rect 42843 2071 42885 2080
rect 3483 2036 3525 2045
rect 3483 1996 3484 2036
rect 3524 1996 3525 2036
rect 3483 1987 3525 1996
rect 4827 2036 4869 2045
rect 4827 1996 4828 2036
rect 4868 1996 4869 2036
rect 4827 1987 4869 1996
rect 12219 2036 12261 2045
rect 12219 1996 12220 2036
rect 12260 1996 12261 2036
rect 12219 1987 12261 1996
rect 13803 2036 13845 2045
rect 13803 1996 13804 2036
rect 13844 1996 13845 2036
rect 13803 1987 13845 1996
rect 14619 2036 14661 2045
rect 14619 1996 14620 2036
rect 14660 1996 14661 2036
rect 14619 1987 14661 1996
rect 24651 2036 24693 2045
rect 24651 1996 24652 2036
rect 24692 1996 24693 2036
rect 24651 1987 24693 1996
rect 25179 2036 25221 2045
rect 25179 1996 25180 2036
rect 25220 1996 25221 2036
rect 25179 1987 25221 1996
rect 28683 2036 28725 2045
rect 28683 1996 28684 2036
rect 28724 1996 28725 2036
rect 28683 1987 28725 1996
rect 31611 2036 31653 2045
rect 31611 1996 31612 2036
rect 31652 1996 31653 2036
rect 31611 1987 31653 1996
rect 45147 2036 45189 2045
rect 45147 1996 45148 2036
rect 45188 1996 45189 2036
rect 45147 1987 45189 1996
rect 1227 1952 1269 1961
rect 1227 1912 1228 1952
rect 1268 1912 1269 1952
rect 1227 1903 1269 1912
rect 1611 1952 1653 1961
rect 1611 1912 1612 1952
rect 1652 1912 1653 1952
rect 1611 1903 1653 1912
rect 1995 1952 2037 1961
rect 1995 1912 1996 1952
rect 2036 1912 2037 1952
rect 1995 1903 2037 1912
rect 2379 1952 2421 1961
rect 2379 1912 2380 1952
rect 2420 1912 2421 1952
rect 2379 1903 2421 1912
rect 3243 1952 3285 1961
rect 3243 1912 3244 1952
rect 3284 1912 3285 1952
rect 3243 1903 3285 1912
rect 4011 1952 4053 1961
rect 4011 1912 4012 1952
rect 4052 1912 4053 1952
rect 4011 1903 4053 1912
rect 4587 1952 4629 1961
rect 4587 1912 4588 1952
rect 4628 1912 4629 1952
rect 4587 1903 4629 1912
rect 4971 1952 5013 1961
rect 4971 1912 4972 1952
rect 5012 1912 5013 1952
rect 4971 1903 5013 1912
rect 5211 1952 5253 1961
rect 5211 1912 5212 1952
rect 5252 1912 5253 1952
rect 5211 1903 5253 1912
rect 5386 1952 5444 1953
rect 5386 1912 5395 1952
rect 5435 1912 5444 1952
rect 5386 1911 5444 1912
rect 5739 1952 5781 1961
rect 5739 1912 5740 1952
rect 5780 1912 5781 1952
rect 5739 1903 5781 1912
rect 6123 1952 6165 1961
rect 6123 1912 6124 1952
rect 6164 1912 6165 1952
rect 6123 1903 6165 1912
rect 6507 1952 6549 1961
rect 6507 1912 6508 1952
rect 6548 1912 6549 1952
rect 6507 1903 6549 1912
rect 8523 1952 8565 1961
rect 8523 1912 8524 1952
rect 8564 1912 8565 1952
rect 8523 1903 8565 1912
rect 8907 1952 8949 1961
rect 8907 1912 8908 1952
rect 8948 1912 8949 1952
rect 8907 1903 8949 1912
rect 10923 1952 10965 1961
rect 10923 1912 10924 1952
rect 10964 1912 10965 1952
rect 10923 1903 10965 1912
rect 11499 1952 11541 1961
rect 11499 1912 11500 1952
rect 11540 1912 11541 1952
rect 11499 1903 11541 1912
rect 11883 1952 11925 1961
rect 11883 1912 11884 1952
rect 11924 1912 11925 1952
rect 11883 1903 11925 1912
rect 12459 1952 12501 1961
rect 12459 1912 12460 1952
rect 12500 1912 12501 1952
rect 12459 1903 12501 1912
rect 12603 1952 12645 1961
rect 12603 1912 12604 1952
rect 12644 1912 12645 1952
rect 12603 1903 12645 1912
rect 12843 1952 12885 1961
rect 12843 1912 12844 1952
rect 12884 1912 12885 1952
rect 12843 1903 12885 1912
rect 14187 1952 14229 1961
rect 14187 1912 14188 1952
rect 14228 1912 14229 1952
rect 14187 1903 14229 1912
rect 14379 1952 14421 1961
rect 14379 1912 14380 1952
rect 14420 1912 14421 1952
rect 14379 1903 14421 1912
rect 14763 1952 14805 1961
rect 14763 1912 14764 1952
rect 14804 1912 14805 1952
rect 14763 1903 14805 1912
rect 15003 1952 15045 1961
rect 15003 1912 15004 1952
rect 15044 1912 15045 1952
rect 15003 1903 15045 1912
rect 15627 1952 15669 1961
rect 15627 1912 15628 1952
rect 15668 1912 15669 1952
rect 15627 1903 15669 1912
rect 15819 1952 15861 1961
rect 15819 1912 15820 1952
rect 15860 1912 15861 1952
rect 15819 1903 15861 1912
rect 16203 1952 16245 1961
rect 16203 1912 16204 1952
rect 16244 1912 16245 1952
rect 16203 1903 16245 1912
rect 16779 1952 16821 1961
rect 16779 1912 16780 1952
rect 16820 1912 16821 1952
rect 16779 1903 16821 1912
rect 18603 1952 18645 1961
rect 18603 1912 18604 1952
rect 18644 1912 18645 1952
rect 18603 1903 18645 1912
rect 18987 1952 19029 1961
rect 18987 1912 18988 1952
rect 19028 1912 19029 1952
rect 18987 1903 19029 1912
rect 19563 1952 19605 1961
rect 19563 1912 19564 1952
rect 19604 1912 19605 1952
rect 19563 1903 19605 1912
rect 19851 1952 19893 1961
rect 19851 1912 19852 1952
rect 19892 1912 19893 1952
rect 19851 1903 19893 1912
rect 20235 1952 20277 1961
rect 20235 1912 20236 1952
rect 20276 1912 20277 1952
rect 20235 1903 20277 1912
rect 22635 1952 22677 1961
rect 22635 1912 22636 1952
rect 22676 1912 22677 1952
rect 22635 1903 22677 1912
rect 23242 1952 23300 1953
rect 23242 1912 23251 1952
rect 23291 1912 23300 1952
rect 23242 1911 23300 1912
rect 23499 1952 23541 1961
rect 23499 1912 23500 1952
rect 23540 1912 23541 1952
rect 23499 1903 23541 1912
rect 24795 1952 24837 1961
rect 24795 1912 24796 1952
rect 24836 1912 24837 1952
rect 24795 1903 24837 1912
rect 25035 1952 25077 1961
rect 25035 1912 25036 1952
rect 25076 1912 25077 1952
rect 25035 1903 25077 1912
rect 25419 1952 25461 1961
rect 25419 1912 25420 1952
rect 25460 1912 25461 1952
rect 25419 1903 25461 1912
rect 25803 1952 25845 1961
rect 25803 1912 25804 1952
rect 25844 1912 25845 1952
rect 25803 1903 25845 1912
rect 30027 1952 30069 1961
rect 30027 1912 30028 1952
rect 30068 1912 30069 1952
rect 30027 1903 30069 1912
rect 31371 1952 31413 1961
rect 31371 1912 31372 1952
rect 31412 1912 31413 1952
rect 31371 1903 31413 1912
rect 31851 1952 31893 1961
rect 31851 1912 31852 1952
rect 31892 1912 31893 1952
rect 31851 1903 31893 1912
rect 32091 1952 32133 1961
rect 32091 1912 32092 1952
rect 32132 1912 32133 1952
rect 32091 1903 32133 1912
rect 34923 1952 34965 1961
rect 34923 1912 34924 1952
rect 34964 1912 34965 1952
rect 34923 1903 34965 1912
rect 36747 1952 36789 1961
rect 36747 1912 36748 1952
rect 36788 1912 36789 1952
rect 36747 1903 36789 1912
rect 39243 1952 39285 1961
rect 39243 1912 39244 1952
rect 39284 1912 39285 1952
rect 39243 1903 39285 1912
rect 40299 1952 40341 1961
rect 40299 1912 40300 1952
rect 40340 1912 40341 1952
rect 40299 1903 40341 1912
rect 40683 1952 40725 1961
rect 40683 1912 40684 1952
rect 40724 1912 40725 1952
rect 40683 1903 40725 1912
rect 42123 1952 42165 1961
rect 42123 1912 42124 1952
rect 42164 1912 42165 1952
rect 42123 1903 42165 1912
rect 42603 1952 42645 1961
rect 42603 1912 42604 1952
rect 42644 1912 42645 1952
rect 42603 1903 42645 1912
rect 42987 1952 43029 1961
rect 42987 1912 42988 1952
rect 43028 1912 43029 1952
rect 42987 1903 43029 1912
rect 43371 1952 43413 1961
rect 43371 1912 43372 1952
rect 43412 1912 43413 1952
rect 43371 1903 43413 1912
rect 43755 1952 43797 1961
rect 43755 1912 43756 1952
rect 43796 1912 43797 1952
rect 43755 1903 43797 1912
rect 44091 1952 44133 1961
rect 44091 1912 44092 1952
rect 44132 1912 44133 1952
rect 44091 1903 44133 1912
rect 44331 1952 44373 1961
rect 44331 1912 44332 1952
rect 44372 1912 44373 1952
rect 44331 1903 44373 1912
rect 44715 1952 44757 1961
rect 44715 1912 44716 1952
rect 44756 1912 44757 1952
rect 44715 1903 44757 1912
rect 44907 1952 44949 1961
rect 44907 1912 44908 1952
rect 44948 1912 44949 1952
rect 44907 1903 44949 1912
rect 6891 1868 6933 1877
rect 6891 1828 6892 1868
rect 6932 1828 6933 1868
rect 6891 1819 6933 1828
rect 8131 1868 8189 1869
rect 8131 1828 8140 1868
rect 8180 1828 8189 1868
rect 8131 1827 8189 1828
rect 9291 1868 9333 1877
rect 9291 1828 9292 1868
rect 9332 1828 9333 1868
rect 9291 1819 9333 1828
rect 10531 1868 10589 1869
rect 10531 1828 10540 1868
rect 10580 1828 10589 1868
rect 10531 1827 10589 1828
rect 13131 1868 13173 1877
rect 13131 1828 13132 1868
rect 13172 1828 13173 1868
rect 13131 1819 13173 1828
rect 13402 1868 13460 1869
rect 13402 1828 13411 1868
rect 13451 1828 13460 1868
rect 13402 1827 13460 1828
rect 17155 1868 17213 1869
rect 17155 1828 17164 1868
rect 17204 1828 17213 1868
rect 17155 1827 17213 1828
rect 18411 1868 18453 1877
rect 18411 1828 18412 1868
rect 18452 1828 18453 1868
rect 18411 1819 18453 1828
rect 20803 1868 20861 1869
rect 20803 1828 20812 1868
rect 20852 1828 20861 1868
rect 20803 1827 20861 1828
rect 22059 1868 22101 1877
rect 22059 1828 22060 1868
rect 22100 1828 22101 1868
rect 22059 1819 22101 1828
rect 23979 1868 24021 1877
rect 23979 1828 23980 1868
rect 24020 1828 24021 1868
rect 23979 1819 24021 1828
rect 24226 1868 24284 1869
rect 24226 1828 24235 1868
rect 24275 1828 24284 1868
rect 24226 1827 24284 1828
rect 24346 1868 24404 1869
rect 24346 1828 24355 1868
rect 24395 1828 24404 1868
rect 24346 1827 24404 1828
rect 25995 1868 26037 1877
rect 25995 1828 25996 1868
rect 26036 1828 26037 1868
rect 25995 1819 26037 1828
rect 27235 1868 27293 1869
rect 27235 1828 27244 1868
rect 27284 1828 27293 1868
rect 27235 1827 27293 1828
rect 28011 1868 28053 1877
rect 28011 1828 28012 1868
rect 28052 1828 28053 1868
rect 28011 1819 28053 1828
rect 28282 1868 28340 1869
rect 28282 1828 28291 1868
rect 28331 1828 28340 1868
rect 28282 1827 28340 1828
rect 28971 1868 29013 1877
rect 28971 1828 28972 1868
rect 29012 1828 29013 1868
rect 28971 1819 29013 1828
rect 29242 1868 29300 1869
rect 29242 1828 29251 1868
rect 29291 1828 29300 1868
rect 29242 1827 29300 1828
rect 29691 1868 29733 1877
rect 29691 1828 29692 1868
rect 29732 1828 29733 1868
rect 29691 1819 29733 1828
rect 32811 1868 32853 1877
rect 32811 1828 32812 1868
rect 32852 1828 32853 1868
rect 32811 1819 32853 1828
rect 34051 1868 34109 1869
rect 34051 1828 34060 1868
rect 34100 1828 34109 1868
rect 34051 1827 34109 1828
rect 1467 1784 1509 1793
rect 1467 1744 1468 1784
rect 1508 1744 1509 1784
rect 1467 1735 1509 1744
rect 11739 1784 11781 1793
rect 11739 1744 11740 1784
rect 11780 1744 11781 1784
rect 11739 1735 11781 1744
rect 12123 1784 12165 1793
rect 12123 1744 12124 1784
rect 12164 1744 12165 1784
rect 12123 1735 12165 1744
rect 13515 1784 13557 1793
rect 13515 1744 13516 1784
rect 13556 1744 13557 1784
rect 13515 1735 13557 1744
rect 16443 1784 16485 1793
rect 16443 1744 16444 1784
rect 16484 1744 16485 1784
rect 16443 1735 16485 1744
rect 19227 1784 19269 1793
rect 19227 1744 19228 1784
rect 19268 1744 19269 1784
rect 19227 1735 19269 1744
rect 25563 1784 25605 1793
rect 25563 1744 25564 1784
rect 25604 1744 25605 1784
rect 25563 1735 25605 1744
rect 27435 1784 27477 1793
rect 27435 1744 27436 1784
rect 27476 1744 27477 1784
rect 27435 1735 27477 1744
rect 28395 1784 28437 1793
rect 28395 1744 28396 1784
rect 28436 1744 28437 1784
rect 28395 1735 28437 1744
rect 29355 1784 29397 1793
rect 29355 1744 29356 1784
rect 29396 1744 29397 1784
rect 29355 1735 29397 1744
rect 42411 1784 42453 1793
rect 42411 1744 42412 1784
rect 42452 1744 42453 1784
rect 42411 1735 42453 1744
rect 43995 1784 44037 1793
rect 43995 1744 43996 1784
rect 44036 1744 44037 1784
rect 43995 1735 44037 1744
rect 2235 1700 2277 1709
rect 2235 1660 2236 1700
rect 2276 1660 2277 1700
rect 2235 1651 2277 1660
rect 5595 1700 5637 1709
rect 5595 1660 5596 1700
rect 5636 1660 5637 1700
rect 5595 1651 5637 1660
rect 6363 1700 6405 1709
rect 6363 1660 6364 1700
rect 6404 1660 6405 1700
rect 6363 1651 6405 1660
rect 6747 1700 6789 1709
rect 6747 1660 6748 1700
rect 6788 1660 6789 1700
rect 6747 1651 6789 1660
rect 8331 1700 8373 1709
rect 8331 1660 8332 1700
rect 8372 1660 8373 1700
rect 8331 1651 8373 1660
rect 11163 1700 11205 1709
rect 11163 1660 11164 1700
rect 11204 1660 11205 1700
rect 11163 1651 11205 1660
rect 15387 1700 15429 1709
rect 15387 1660 15388 1700
rect 15428 1660 15429 1700
rect 15387 1651 15429 1660
rect 16059 1700 16101 1709
rect 16059 1660 16060 1700
rect 16100 1660 16101 1700
rect 16059 1651 16101 1660
rect 18843 1700 18885 1709
rect 18843 1660 18844 1700
rect 18884 1660 18885 1700
rect 18843 1651 18885 1660
rect 19323 1700 19365 1709
rect 19323 1660 19324 1700
rect 19364 1660 19365 1700
rect 19323 1651 19365 1660
rect 20091 1700 20133 1709
rect 20091 1660 20092 1700
rect 20132 1660 20133 1700
rect 20091 1651 20133 1660
rect 20475 1700 20517 1709
rect 20475 1660 20476 1700
rect 20516 1660 20517 1700
rect 20475 1651 20517 1660
rect 22395 1700 22437 1709
rect 22395 1660 22396 1700
rect 22436 1660 22437 1700
rect 22395 1651 22437 1660
rect 23067 1700 23109 1709
rect 23067 1660 23068 1700
rect 23108 1660 23109 1700
rect 23067 1651 23109 1660
rect 23739 1700 23781 1709
rect 23739 1660 23740 1700
rect 23780 1660 23781 1700
rect 23739 1651 23781 1660
rect 29787 1700 29829 1709
rect 29787 1660 29788 1700
rect 29828 1660 29829 1700
rect 29787 1651 29829 1660
rect 40282 1700 40340 1701
rect 40282 1660 40291 1700
rect 40331 1660 40340 1700
rect 40282 1659 40340 1660
rect 41067 1700 41109 1709
rect 41067 1660 41068 1700
rect 41108 1660 41109 1700
rect 41067 1651 41109 1660
rect 41355 1700 41397 1709
rect 41355 1660 41356 1700
rect 41396 1660 41397 1700
rect 41355 1651 41397 1660
rect 41643 1700 41685 1709
rect 41643 1660 41644 1700
rect 41684 1660 41685 1700
rect 41643 1651 41685 1660
rect 42315 1700 42357 1709
rect 42315 1660 42316 1700
rect 42356 1660 42357 1700
rect 42315 1651 42357 1660
rect 43227 1700 43269 1709
rect 43227 1660 43228 1700
rect 43268 1660 43269 1700
rect 43227 1651 43269 1660
rect 43611 1700 43653 1709
rect 43611 1660 43612 1700
rect 43652 1660 43653 1700
rect 43611 1651 43653 1660
rect 1152 1532 45216 1556
rect 1152 1492 4928 1532
rect 4968 1492 5010 1532
rect 5050 1492 5092 1532
rect 5132 1492 5174 1532
rect 5214 1492 5256 1532
rect 5296 1492 20048 1532
rect 20088 1492 20130 1532
rect 20170 1492 20212 1532
rect 20252 1492 20294 1532
rect 20334 1492 20376 1532
rect 20416 1492 35168 1532
rect 35208 1492 35250 1532
rect 35290 1492 35332 1532
rect 35372 1492 35414 1532
rect 35454 1492 35496 1532
rect 35536 1492 45216 1532
rect 1152 1468 45216 1492
<< via1 >>
rect 3688 9808 3728 9848
rect 3770 9808 3810 9848
rect 3852 9808 3892 9848
rect 3934 9808 3974 9848
rect 4016 9808 4056 9848
rect 18808 9808 18848 9848
rect 18890 9808 18930 9848
rect 18972 9808 19012 9848
rect 19054 9808 19094 9848
rect 19136 9808 19176 9848
rect 33928 9808 33968 9848
rect 34010 9808 34050 9848
rect 34092 9808 34132 9848
rect 34174 9808 34214 9848
rect 34256 9808 34296 9848
rect 3388 9640 3428 9680
rect 8188 9640 8228 9680
rect 9916 9640 9956 9680
rect 11548 9640 11588 9680
rect 12316 9640 12356 9680
rect 14524 9640 14564 9680
rect 15676 9640 15716 9680
rect 18076 9640 18116 9680
rect 22012 9640 22052 9680
rect 28444 9640 28484 9680
rect 29212 9640 29252 9680
rect 32284 9640 32324 9680
rect 36892 9640 36932 9680
rect 37276 9640 37316 9680
rect 38812 9640 38852 9680
rect 39196 9640 39236 9680
rect 43228 9640 43268 9680
rect 44380 9640 44420 9680
rect 8332 9556 8372 9596
rect 9532 9556 9572 9596
rect 10060 9556 10100 9596
rect 11932 9556 11972 9596
rect 20140 9556 20180 9596
rect 22108 9556 22148 9596
rect 25228 9556 25268 9596
rect 27532 9556 27572 9596
rect 31804 9556 31844 9596
rect 34300 9556 34340 9596
rect 35596 9556 35636 9596
rect 36124 9556 36164 9596
rect 36508 9556 36548 9596
rect 1228 9472 1268 9512
rect 1612 9472 1652 9512
rect 1996 9472 2036 9512
rect 2380 9472 2420 9512
rect 2764 9472 2804 9512
rect 3148 9472 3188 9512
rect 7948 9472 7988 9512
rect 9292 9472 9332 9512
rect 9676 9472 9716 9512
rect 11308 9472 11348 9512
rect 11692 9472 11732 9512
rect 12076 9472 12116 9512
rect 14284 9472 14324 9512
rect 14668 9472 14708 9512
rect 15052 9472 15092 9512
rect 15436 9472 15476 9512
rect 15820 9472 15860 9512
rect 17836 9472 17876 9512
rect 18796 9472 18836 9512
rect 18988 9472 19028 9512
rect 20620 9472 20660 9512
rect 21196 9472 21236 9512
rect 21340 9472 21380 9512
rect 21580 9472 21620 9512
rect 21772 9472 21812 9512
rect 22348 9472 22388 9512
rect 22732 9472 22772 9512
rect 23116 9472 23156 9512
rect 23308 9472 23348 9512
rect 23884 9472 23924 9512
rect 24268 9472 24308 9512
rect 25612 9472 25652 9512
rect 25804 9472 25844 9512
rect 26188 9472 26228 9512
rect 27916 9472 27956 9512
rect 28300 9472 28340 9512
rect 28684 9472 28724 9512
rect 29068 9472 29108 9512
rect 29452 9472 29492 9512
rect 29836 9472 29876 9512
rect 30028 9472 30068 9512
rect 30604 9472 30644 9512
rect 30988 9472 31028 9512
rect 31372 9472 31412 9512
rect 31564 9472 31604 9512
rect 32140 9472 32180 9512
rect 32524 9472 32564 9512
rect 34540 9472 34580 9512
rect 35980 9472 36020 9512
rect 36364 9472 36404 9512
rect 36748 9472 36788 9512
rect 37132 9472 37172 9512
rect 37516 9472 37556 9512
rect 37900 9472 37940 9512
rect 38284 9472 38324 9512
rect 38668 9472 38708 9512
rect 39052 9472 39092 9512
rect 39436 9472 39476 9512
rect 39820 9472 39860 9512
rect 41020 9472 41060 9512
rect 41260 9472 41300 9512
rect 42604 9472 42644 9512
rect 42988 9472 43028 9512
rect 43468 9472 43508 9512
rect 43756 9472 43796 9512
rect 44140 9472 44180 9512
rect 44524 9472 44564 9512
rect 45100 9472 45140 9512
rect 6316 9388 6356 9428
rect 7564 9388 7604 9428
rect 8716 9379 8756 9419
rect 9004 9388 9044 9428
rect 10444 9379 10484 9419
rect 10732 9388 10772 9428
rect 12652 9388 12692 9428
rect 13900 9388 13940 9428
rect 16204 9388 16244 9428
rect 17452 9388 17492 9428
rect 19468 9388 19508 9428
rect 19747 9388 19787 9428
rect 24556 9388 24596 9428
rect 24835 9388 24875 9428
rect 26860 9388 26900 9428
rect 27115 9388 27155 9428
rect 27235 9388 27275 9428
rect 32716 9388 32756 9428
rect 33964 9388 34004 9428
rect 34924 9388 34964 9428
rect 35203 9388 35243 9428
rect 8620 9304 8660 9344
rect 10348 9304 10388 9344
rect 12460 9304 12500 9344
rect 14908 9304 14948 9344
rect 19852 9304 19892 9344
rect 20860 9304 20900 9344
rect 23548 9304 23588 9344
rect 24940 9304 24980 9344
rect 29596 9304 29636 9344
rect 30268 9304 30308 9344
rect 35308 9304 35348 9344
rect 39580 9304 39620 9344
rect 44764 9304 44804 9344
rect 1468 9220 1508 9260
rect 1852 9220 1892 9260
rect 2236 9220 2276 9260
rect 2620 9220 2660 9260
rect 3004 9220 3044 9260
rect 7756 9220 7796 9260
rect 15292 9220 15332 9260
rect 16060 9220 16100 9260
rect 17644 9220 17684 9260
rect 18412 9220 18452 9260
rect 18556 9220 18596 9260
rect 19228 9220 19268 9260
rect 20956 9220 20996 9260
rect 22492 9220 22532 9260
rect 22876 9220 22916 9260
rect 23644 9220 23684 9260
rect 24028 9220 24068 9260
rect 25372 9220 25412 9260
rect 26044 9220 26084 9260
rect 26428 9220 26468 9260
rect 27676 9220 27716 9260
rect 28060 9220 28100 9260
rect 28828 9220 28868 9260
rect 30364 9220 30404 9260
rect 30748 9220 30788 9260
rect 31132 9220 31172 9260
rect 31900 9220 31940 9260
rect 34156 9220 34196 9260
rect 35740 9220 35780 9260
rect 37660 9220 37700 9260
rect 38044 9220 38084 9260
rect 38428 9220 38468 9260
rect 40195 9220 40235 9260
rect 40483 9220 40523 9260
rect 40771 9220 40811 9260
rect 41443 9220 41483 9260
rect 41731 9220 41771 9260
rect 42019 9220 42059 9260
rect 42307 9220 42347 9260
rect 42844 9220 42884 9260
rect 43459 9220 43499 9260
rect 43996 9220 44036 9260
rect 44860 9220 44900 9260
rect 4928 9052 4968 9092
rect 5010 9052 5050 9092
rect 5092 9052 5132 9092
rect 5174 9052 5214 9092
rect 5256 9052 5296 9092
rect 20048 9052 20088 9092
rect 20130 9052 20170 9092
rect 20212 9052 20252 9092
rect 20294 9052 20334 9092
rect 20376 9052 20416 9092
rect 35168 9052 35208 9092
rect 35250 9052 35290 9092
rect 35332 9052 35372 9092
rect 35414 9052 35454 9092
rect 35496 9052 35536 9092
rect 1468 8884 1508 8924
rect 2620 8884 2660 8924
rect 8236 8884 8276 8924
rect 10732 8884 10772 8924
rect 13564 8884 13604 8924
rect 13948 8884 13988 8924
rect 15532 8884 15572 8924
rect 16156 8884 16196 8924
rect 17740 8884 17780 8924
rect 22636 8884 22676 8924
rect 26284 8884 26324 8924
rect 32668 8884 32708 8924
rect 35260 8884 35300 8924
rect 35980 8884 36020 8924
rect 38332 8884 38372 8924
rect 40924 8884 40964 8924
rect 41356 8884 41396 8924
rect 41731 8884 41771 8924
rect 42796 8884 42836 8924
rect 43708 8884 43748 8924
rect 44380 8884 44420 8924
rect 5836 8800 5876 8840
rect 11212 8800 11252 8840
rect 13180 8800 13220 8840
rect 18268 8800 18308 8840
rect 27244 8800 27284 8840
rect 28348 8800 28388 8840
rect 30700 8800 30740 8840
rect 32572 8800 32612 8840
rect 33676 8800 33716 8840
rect 34828 8800 34868 8840
rect 35164 8800 35204 8840
rect 39388 8800 39428 8840
rect 43324 8800 43364 8840
rect 4396 8716 4436 8756
rect 5644 8707 5684 8747
rect 6796 8716 6836 8756
rect 8044 8707 8084 8747
rect 8995 8716 9035 8756
rect 9100 8716 9140 8756
rect 9484 8716 9524 8756
rect 10060 8707 10100 8747
rect 10540 8707 10580 8747
rect 11404 8707 11444 8747
rect 12652 8716 12692 8756
rect 14092 8716 14132 8756
rect 15340 8707 15380 8747
rect 16300 8716 16340 8756
rect 17548 8707 17588 8747
rect 18862 8716 18902 8756
rect 18988 8716 19028 8756
rect 19372 8716 19412 8756
rect 19943 8716 19983 8756
rect 20428 8707 20468 8747
rect 20899 8716 20939 8756
rect 21004 8716 21044 8756
rect 21388 8716 21428 8756
rect 21964 8707 22004 8747
rect 22444 8707 22484 8747
rect 22828 8716 22868 8756
rect 24547 8716 24587 8756
rect 24652 8716 24692 8756
rect 1228 8632 1268 8672
rect 1612 8632 1652 8672
rect 1996 8632 2036 8672
rect 2236 8632 2276 8672
rect 2380 8632 2420 8672
rect 8524 8632 8564 8672
rect 8764 8632 8804 8672
rect 9580 8632 9620 8672
rect 12940 8632 12980 8672
rect 13324 8632 13364 8672
rect 13708 8632 13748 8672
rect 15916 8632 15956 8672
rect 18028 8632 18068 8672
rect 18412 8632 18452 8672
rect 18652 8632 18692 8672
rect 19468 8632 19508 8672
rect 20659 8632 20699 8672
rect 24080 8674 24120 8714
rect 25036 8716 25076 8756
rect 25612 8707 25652 8747
rect 26092 8707 26132 8747
rect 26860 8716 26900 8756
rect 27139 8716 27179 8756
rect 29260 8707 29300 8747
rect 30508 8716 30548 8756
rect 30892 8707 30932 8747
rect 32140 8716 32180 8756
rect 33292 8716 33332 8756
rect 33571 8716 33611 8756
rect 34444 8716 34484 8756
rect 34723 8716 34763 8756
rect 36172 8707 36212 8747
rect 37420 8716 37460 8756
rect 42892 8716 42932 8756
rect 44716 8716 44756 8756
rect 21484 8632 21524 8672
rect 25132 8632 25172 8672
rect 27676 8632 27716 8672
rect 27916 8632 27956 8672
rect 28108 8632 28148 8672
rect 28684 8632 28724 8672
rect 29059 8632 29099 8672
rect 32332 8632 32372 8672
rect 32908 8632 32948 8672
rect 35500 8632 35540 8672
rect 37564 8632 37604 8672
rect 37804 8632 37844 8672
rect 37948 8632 37988 8672
rect 38188 8632 38228 8672
rect 38572 8632 38612 8672
rect 38716 8632 38756 8672
rect 38956 8632 38996 8672
rect 39148 8632 39188 8672
rect 39532 8632 39572 8672
rect 39868 8632 39908 8672
rect 40108 8632 40148 8672
rect 40492 8632 40532 8672
rect 40780 8632 40820 8672
rect 41164 8632 41204 8672
rect 42028 8632 42068 8672
rect 42316 8632 42356 8672
rect 42604 8632 42644 8672
rect 43084 8632 43124 8672
rect 43468 8632 43508 8672
rect 43948 8632 43988 8672
rect 44140 8632 44180 8672
rect 44908 8632 44948 8672
rect 28444 8548 28484 8588
rect 39772 8548 39812 8588
rect 1852 8464 1892 8504
rect 24268 8464 24308 8504
rect 27532 8464 27572 8504
rect 33964 8464 34004 8504
rect 45148 8464 45188 8504
rect 3688 8296 3728 8336
rect 3770 8296 3810 8336
rect 3852 8296 3892 8336
rect 3934 8296 3974 8336
rect 4016 8296 4056 8336
rect 18808 8296 18848 8336
rect 18890 8296 18930 8336
rect 18972 8296 19012 8336
rect 19054 8296 19094 8336
rect 19136 8296 19176 8336
rect 33928 8296 33968 8336
rect 34010 8296 34050 8336
rect 34092 8296 34132 8336
rect 34174 8296 34214 8336
rect 34256 8296 34296 8336
rect 4348 8128 4388 8168
rect 10252 8128 10292 8168
rect 11836 8128 11876 8168
rect 16444 8128 16484 8168
rect 25900 8128 25940 8168
rect 30652 8128 30692 8168
rect 32812 8128 32852 8168
rect 39388 8128 39428 8168
rect 44380 8128 44420 8168
rect 12220 8044 12260 8084
rect 20044 8044 20084 8084
rect 22828 8044 22868 8084
rect 30556 8044 30596 8084
rect 36508 8044 36548 8084
rect 1228 7960 1268 8000
rect 1612 7960 1652 8000
rect 4108 7960 4148 8000
rect 9484 7960 9524 8000
rect 9724 7960 9764 8000
rect 9868 7960 9908 8000
rect 11212 7960 11252 8000
rect 11596 7960 11636 8000
rect 11980 7960 12020 8000
rect 12355 7960 12395 8000
rect 16204 7960 16244 8000
rect 16588 7960 16628 8000
rect 16972 7960 17012 8000
rect 17212 7960 17252 8000
rect 20716 7960 20756 8000
rect 21100 7960 21140 8000
rect 21484 7960 21524 8000
rect 21676 7960 21716 8000
rect 22972 7960 23012 8000
rect 23212 7960 23252 8000
rect 23356 7960 23396 8000
rect 23596 7960 23636 8000
rect 28492 7960 28532 8000
rect 30124 7960 30164 8000
rect 30316 7960 30356 8000
rect 30892 7960 30932 8000
rect 34636 7960 34676 8000
rect 36124 7960 36164 8000
rect 36364 7960 36404 8000
rect 36748 7960 36788 8000
rect 37132 7960 37172 8000
rect 39628 7960 39668 8000
rect 41452 7960 41492 8000
rect 42124 7960 42164 8000
rect 44140 7960 44180 8000
rect 44524 7960 44564 8000
rect 44908 7960 44948 8000
rect 4492 7876 4532 7916
rect 5740 7876 5780 7916
rect 7564 7876 7604 7916
rect 8812 7876 8852 7916
rect 10636 7867 10676 7907
rect 10924 7876 10964 7916
rect 12556 7876 12596 7916
rect 13804 7876 13844 7916
rect 14284 7876 14324 7916
rect 15532 7876 15572 7916
rect 17356 7876 17396 7916
rect 18604 7876 18644 7916
rect 19372 7876 19412 7916
rect 19651 7876 19691 7916
rect 22156 7876 22196 7916
rect 22435 7876 22475 7916
rect 24460 7876 24500 7916
rect 25708 7876 25748 7916
rect 26284 7876 26324 7916
rect 27532 7876 27572 7916
rect 28003 7876 28043 7916
rect 28108 7876 28148 7916
rect 28588 7876 28628 7916
rect 29068 7876 29108 7916
rect 29556 7876 29596 7916
rect 31372 7876 31412 7916
rect 32620 7876 32660 7916
rect 33004 7876 33044 7916
rect 34252 7876 34292 7916
rect 35308 7876 35348 7916
rect 35587 7876 35627 7916
rect 36028 7876 36068 7916
rect 37516 7876 37556 7916
rect 38764 7876 38804 7916
rect 10540 7792 10580 7832
rect 16828 7792 16868 7832
rect 18796 7792 18836 7832
rect 19740 7792 19780 7832
rect 21244 7792 21284 7832
rect 22540 7792 22580 7832
rect 27724 7792 27764 7832
rect 34876 7792 34916 7832
rect 35692 7792 35732 7832
rect 36892 7792 36932 7832
rect 41836 7792 41876 7832
rect 42412 7792 42452 7832
rect 42700 7792 42740 7832
rect 42988 7792 43028 7832
rect 43276 7792 43316 7832
rect 1468 7708 1508 7748
rect 1852 7708 1892 7748
rect 5932 7708 5972 7748
rect 9004 7708 9044 7748
rect 10108 7708 10148 7748
rect 11452 7708 11492 7748
rect 15724 7708 15764 7748
rect 20476 7708 20516 7748
rect 20860 7708 20900 7748
rect 21916 7708 21956 7748
rect 29740 7708 29780 7748
rect 29884 7708 29924 7748
rect 34444 7708 34484 7748
rect 38956 7708 38996 7748
rect 40963 7708 41003 7748
rect 41212 7708 41252 7748
rect 42211 7708 42251 7748
rect 43651 7708 43691 7748
rect 43843 7708 43883 7748
rect 44764 7708 44804 7748
rect 45148 7708 45188 7748
rect 4928 7540 4968 7580
rect 5010 7540 5050 7580
rect 5092 7540 5132 7580
rect 5174 7540 5214 7580
rect 5256 7540 5296 7580
rect 20048 7540 20088 7580
rect 20130 7540 20170 7580
rect 20212 7540 20252 7580
rect 20294 7540 20334 7580
rect 20376 7540 20416 7580
rect 35168 7540 35208 7580
rect 35250 7540 35290 7580
rect 35332 7540 35372 7580
rect 35414 7540 35454 7580
rect 35496 7540 35536 7580
rect 10108 7372 10148 7412
rect 29356 7372 29396 7412
rect 33340 7372 33380 7412
rect 33724 7372 33764 7412
rect 41827 7372 41867 7412
rect 42499 7372 42539 7412
rect 42787 7372 42827 7412
rect 9772 7288 9812 7328
rect 11020 7288 11060 7328
rect 21676 7288 21716 7328
rect 32956 7288 32996 7328
rect 9388 7204 9428 7244
rect 9667 7204 9707 7244
rect 10636 7204 10676 7244
rect 10915 7204 10955 7244
rect 17068 7204 17108 7244
rect 18316 7195 18356 7235
rect 21292 7204 21332 7244
rect 21571 7204 21611 7244
rect 23020 7204 23060 7244
rect 23275 7204 23315 7244
rect 23395 7204 23435 7244
rect 27916 7204 27956 7244
rect 29164 7195 29204 7235
rect 30700 7204 30740 7244
rect 31948 7195 31988 7235
rect 34435 7204 34475 7244
rect 34540 7204 34580 7244
rect 34924 7204 34964 7244
rect 35500 7195 35540 7235
rect 35980 7195 36020 7235
rect 39436 7204 39476 7244
rect 40684 7195 40724 7235
rect 1228 7120 1268 7160
rect 1612 7120 1652 7160
rect 1852 7120 1892 7160
rect 3532 7120 3572 7160
rect 6316 7120 6356 7160
rect 6556 7120 6596 7160
rect 8140 7120 8180 7160
rect 8524 7120 8564 7160
rect 8908 7120 8948 7160
rect 9148 7120 9188 7160
rect 11692 7120 11732 7160
rect 12076 7120 12116 7160
rect 12460 7120 12500 7160
rect 12844 7120 12884 7160
rect 13228 7120 13268 7160
rect 13468 7120 13508 7160
rect 13612 7120 13652 7160
rect 13996 7120 14036 7160
rect 14380 7120 14420 7160
rect 14764 7120 14804 7160
rect 15004 7120 15044 7160
rect 15148 7120 15188 7160
rect 15532 7120 15572 7160
rect 15916 7120 15956 7160
rect 16300 7120 16340 7160
rect 16684 7120 16724 7160
rect 18892 7120 18932 7160
rect 19276 7120 19316 7160
rect 19660 7120 19700 7160
rect 19900 7120 19940 7160
rect 20236 7120 20276 7160
rect 20620 7120 20660 7160
rect 20764 7120 20804 7160
rect 21004 7120 21044 7160
rect 22348 7120 22388 7160
rect 22540 7120 22580 7160
rect 23980 7120 24020 7160
rect 25132 7120 25172 7160
rect 25708 7120 25748 7160
rect 26092 7120 26132 7160
rect 27052 7120 27092 7160
rect 27724 7120 27764 7160
rect 29500 7120 29540 7160
rect 30124 7120 30164 7160
rect 30316 7120 30356 7160
rect 32524 7120 32564 7160
rect 32716 7120 32756 7160
rect 33100 7120 33140 7160
rect 33484 7120 33524 7160
rect 34060 7120 34100 7160
rect 35020 7120 35060 7160
rect 36556 7120 36596 7160
rect 36940 7120 36980 7160
rect 37324 7120 37364 7160
rect 37708 7120 37748 7160
rect 42220 7120 42260 7160
rect 43180 7120 43220 7160
rect 43468 7120 43508 7160
rect 43756 7120 43796 7160
rect 44044 7120 44084 7160
rect 44332 7120 44372 7160
rect 44524 7120 44564 7160
rect 44908 7120 44948 7160
rect 12316 7036 12356 7076
rect 14236 7036 14276 7076
rect 15772 7036 15812 7076
rect 16540 7036 16580 7076
rect 19516 7036 19556 7076
rect 21964 7036 22004 7076
rect 27484 7036 27524 7076
rect 29788 7036 29828 7076
rect 32140 7036 32180 7076
rect 44764 7036 44804 7076
rect 1468 6952 1508 6992
rect 3772 6952 3812 6992
rect 8380 6952 8420 6992
rect 8764 6952 8804 6992
rect 11308 6952 11348 6992
rect 11932 6952 11972 6992
rect 12700 6952 12740 6992
rect 13084 6952 13124 6992
rect 13852 6952 13892 6992
rect 14620 6952 14660 6992
rect 15388 6952 15428 6992
rect 16156 6952 16196 6992
rect 16924 6952 16964 6992
rect 18508 6952 18548 6992
rect 19132 6952 19172 6992
rect 19996 6952 20036 6992
rect 20380 6952 20420 6992
rect 22108 6952 22148 6992
rect 22780 6952 22820 6992
rect 23692 6952 23732 6992
rect 24220 6952 24260 6992
rect 25372 6952 25412 6992
rect 25948 6952 25988 6992
rect 26332 6952 26372 6992
rect 27292 6952 27332 6992
rect 29884 6952 29924 6992
rect 30556 6952 30596 6992
rect 32284 6952 32324 6992
rect 33820 6952 33860 6992
rect 36211 6952 36251 6992
rect 36316 6952 36356 6992
rect 36700 6952 36740 6992
rect 37084 6952 37124 6992
rect 37468 6952 37508 6992
rect 40876 6952 40916 6992
rect 41980 6952 42020 6992
rect 45148 6952 45188 6992
rect 3688 6784 3728 6824
rect 3770 6784 3810 6824
rect 3852 6784 3892 6824
rect 3934 6784 3974 6824
rect 4016 6784 4056 6824
rect 18808 6784 18848 6824
rect 18890 6784 18930 6824
rect 18972 6784 19012 6824
rect 19054 6784 19094 6824
rect 19136 6784 19176 6824
rect 33928 6784 33968 6824
rect 34010 6784 34050 6824
rect 34092 6784 34132 6824
rect 34174 6784 34214 6824
rect 34256 6784 34296 6824
rect 10108 6616 10148 6656
rect 12508 6616 12548 6656
rect 12892 6616 12932 6656
rect 13276 6616 13316 6656
rect 15292 6616 15332 6656
rect 17404 6616 17444 6656
rect 17788 6616 17828 6656
rect 18460 6616 18500 6656
rect 20044 6616 20084 6656
rect 22156 6616 22196 6656
rect 36748 6616 36788 6656
rect 41836 6616 41876 6656
rect 43996 6616 44036 6656
rect 27964 6532 28004 6572
rect 34348 6532 34388 6572
rect 35308 6532 35348 6572
rect 36556 6532 36596 6572
rect 42796 6532 42836 6572
rect 1228 6448 1268 6488
rect 1612 6448 1652 6488
rect 6220 6448 6260 6488
rect 7651 6448 7691 6488
rect 9484 6448 9524 6488
rect 9868 6448 9908 6488
rect 10828 6448 10868 6488
rect 12268 6448 12308 6488
rect 12652 6448 12692 6488
rect 13036 6448 13076 6488
rect 15532 6448 15572 6488
rect 17644 6448 17684 6488
rect 18028 6448 18068 6488
rect 18220 6448 18260 6488
rect 20236 6448 20276 6488
rect 20476 6448 20516 6488
rect 22924 6448 22964 6488
rect 24556 6448 24596 6488
rect 27148 6448 27188 6488
rect 28204 6448 28244 6488
rect 39532 6448 39572 6488
rect 43180 6448 43220 6488
rect 44236 6448 44276 6488
rect 44524 6448 44564 6488
rect 44908 6448 44948 6488
rect 3724 6364 3764 6404
rect 4972 6364 5012 6404
rect 5731 6364 5771 6404
rect 5836 6364 5876 6404
rect 6316 6364 6356 6404
rect 6796 6364 6836 6404
rect 7315 6364 7355 6404
rect 7852 6364 7892 6404
rect 9100 6364 9140 6404
rect 10318 6363 10358 6403
rect 10444 6364 10484 6404
rect 10924 6364 10964 6404
rect 11404 6364 11444 6404
rect 11923 6364 11963 6404
rect 13612 6364 13652 6404
rect 14860 6364 14900 6404
rect 16012 6364 16052 6404
rect 17260 6364 17300 6404
rect 18604 6364 18644 6404
rect 19852 6364 19892 6404
rect 20716 6364 20756 6404
rect 21972 6364 22012 6404
rect 22435 6364 22475 6404
rect 22540 6364 22580 6404
rect 23020 6364 23060 6404
rect 23500 6364 23540 6404
rect 24019 6364 24059 6404
rect 25228 6364 25268 6404
rect 26476 6364 26516 6404
rect 28684 6364 28724 6404
rect 29932 6364 29972 6404
rect 30316 6364 30356 6404
rect 31564 6364 31604 6404
rect 31948 6364 31988 6404
rect 33196 6364 33236 6404
rect 33676 6364 33716 6404
rect 33955 6364 33995 6404
rect 34636 6364 34676 6404
rect 34915 6364 34955 6404
rect 35884 6364 35924 6404
rect 36139 6364 36179 6404
rect 36259 6364 36299 6404
rect 36940 6364 36980 6404
rect 38188 6364 38228 6404
rect 39022 6364 39062 6404
rect 39148 6364 39188 6404
rect 39628 6364 39668 6404
rect 40108 6364 40148 6404
rect 40596 6364 40636 6404
rect 41164 6364 41204 6404
rect 41443 6364 41483 6404
rect 42124 6364 42164 6404
rect 42403 6364 42443 6404
rect 24316 6280 24356 6320
rect 25036 6280 25076 6320
rect 28492 6280 28532 6320
rect 34060 6280 34100 6320
rect 35020 6280 35060 6320
rect 41548 6280 41588 6320
rect 42508 6280 42548 6320
rect 45148 6280 45188 6320
rect 1468 6196 1508 6236
rect 1852 6196 1892 6236
rect 5164 6196 5204 6236
rect 7468 6196 7508 6236
rect 9724 6196 9764 6236
rect 12076 6196 12116 6236
rect 13420 6196 13460 6236
rect 15820 6196 15860 6236
rect 24172 6196 24212 6236
rect 27388 6196 27428 6236
rect 31756 6196 31796 6236
rect 33388 6196 33428 6236
rect 40780 6196 40820 6236
rect 42940 6196 42980 6236
rect 43555 6196 43595 6236
rect 43843 6196 43883 6236
rect 44764 6196 44804 6236
rect 4928 6028 4968 6068
rect 5010 6028 5050 6068
rect 5092 6028 5132 6068
rect 5174 6028 5214 6068
rect 5256 6028 5296 6068
rect 20048 6028 20088 6068
rect 20130 6028 20170 6068
rect 20212 6028 20252 6068
rect 20294 6028 20334 6068
rect 20376 6028 20416 6068
rect 35168 6028 35208 6068
rect 35250 6028 35290 6068
rect 35332 6028 35372 6068
rect 35414 6028 35454 6068
rect 35496 6028 35536 6068
rect 32476 5860 32516 5900
rect 41932 5860 41972 5900
rect 43171 5860 43211 5900
rect 43459 5860 43499 5900
rect 44236 5860 44276 5900
rect 6028 5776 6068 5816
rect 8812 5776 8852 5816
rect 11116 5776 11156 5816
rect 11836 5776 11876 5816
rect 23692 5776 23732 5816
rect 3532 5692 3572 5732
rect 4784 5683 4824 5723
rect 5644 5692 5684 5732
rect 5923 5692 5963 5732
rect 8941 5692 8981 5732
rect 9196 5692 9236 5732
rect 10732 5692 10772 5732
rect 11011 5692 11051 5732
rect 13516 5683 13556 5723
rect 14724 5692 14764 5732
rect 15916 5683 15956 5723
rect 17164 5692 17204 5732
rect 18028 5692 18068 5732
rect 19276 5683 19316 5723
rect 20044 5692 20084 5732
rect 21292 5683 21332 5723
rect 23308 5692 23348 5732
rect 23587 5692 23627 5732
rect 25900 5683 25940 5723
rect 27148 5692 27188 5732
rect 27628 5692 27668 5732
rect 28876 5683 28916 5723
rect 30508 5692 30548 5732
rect 31756 5683 31796 5723
rect 33379 5692 33419 5732
rect 33484 5692 33524 5732
rect 34444 5683 34484 5723
rect 34924 5683 34964 5723
rect 35155 5692 35195 5732
rect 38572 5692 38612 5732
rect 39820 5683 39860 5723
rect 40492 5692 40532 5732
rect 41740 5683 41780 5723
rect 1228 5608 1268 5648
rect 1612 5608 1652 5648
rect 1996 5608 2036 5648
rect 6508 5608 6548 5648
rect 10252 5608 10292 5648
rect 11596 5608 11636 5648
rect 11980 5608 12020 5648
rect 12412 5608 12452 5648
rect 12652 5608 12692 5648
rect 12844 5608 12884 5648
rect 13315 5608 13355 5648
rect 14956 5608 14996 5648
rect 15532 5608 15572 5648
rect 22108 5608 22148 5648
rect 22348 5608 22388 5648
rect 24364 5608 24404 5648
rect 25324 5608 25364 5648
rect 25699 5608 25739 5648
rect 29452 5608 29492 5648
rect 29836 5608 29876 5648
rect 32332 5608 32372 5648
rect 32716 5608 32756 5648
rect 33100 5608 33140 5648
rect 33872 5608 33912 5648
rect 34003 5608 34043 5648
rect 35260 5608 35300 5648
rect 35500 5608 35540 5648
rect 35884 5608 35924 5648
rect 36268 5608 36308 5648
rect 37180 5608 37220 5648
rect 37420 5608 37460 5648
rect 37996 5608 38036 5648
rect 42892 5608 42932 5648
rect 43180 5608 43220 5648
rect 43756 5608 43796 5648
rect 44332 5608 44372 5648
rect 44524 5608 44564 5648
rect 44908 5608 44948 5648
rect 45148 5608 45188 5648
rect 2236 5524 2276 5564
rect 6316 5524 6356 5564
rect 11404 5524 11444 5564
rect 15196 5524 15236 5564
rect 19468 5524 19508 5564
rect 21484 5524 21524 5564
rect 24124 5524 24164 5564
rect 25564 5524 25604 5564
rect 29068 5524 29108 5564
rect 31948 5524 31988 5564
rect 32092 5524 32132 5564
rect 1468 5440 1508 5480
rect 1852 5440 1892 5480
rect 4972 5440 5012 5480
rect 6748 5440 6788 5480
rect 8524 5440 8564 5480
rect 10492 5440 10532 5480
rect 12220 5440 12260 5480
rect 13084 5440 13124 5480
rect 15292 5440 15332 5480
rect 15724 5440 15764 5480
rect 23980 5440 24020 5480
rect 29212 5440 29252 5480
rect 30076 5440 30116 5480
rect 32860 5440 32900 5480
rect 35644 5440 35684 5480
rect 36028 5440 36068 5480
rect 38236 5440 38276 5480
rect 40012 5440 40052 5480
rect 44764 5440 44804 5480
rect 3688 5272 3728 5312
rect 3770 5272 3810 5312
rect 3852 5272 3892 5312
rect 3934 5272 3974 5312
rect 4016 5272 4056 5312
rect 18808 5272 18848 5312
rect 18890 5272 18930 5312
rect 18972 5272 19012 5312
rect 19054 5272 19094 5312
rect 19136 5272 19176 5312
rect 33928 5272 33968 5312
rect 34010 5272 34050 5312
rect 34092 5272 34132 5312
rect 34174 5272 34214 5312
rect 34256 5272 34296 5312
rect 6124 5104 6164 5144
rect 11452 5104 11492 5144
rect 12364 5104 12404 5144
rect 14236 5104 14276 5144
rect 36364 5104 36404 5144
rect 7084 5020 7124 5060
rect 14620 5020 14660 5060
rect 33772 5020 33812 5060
rect 39196 5020 39236 5060
rect 41452 5020 41492 5060
rect 1228 4936 1268 4976
rect 1612 4936 1652 4976
rect 9772 4936 9812 4976
rect 11692 4936 11732 4976
rect 11884 4936 11924 4976
rect 14476 4936 14516 4976
rect 14860 4936 14900 4976
rect 19756 4936 19796 4976
rect 20092 4936 20132 4976
rect 20332 4936 20372 4976
rect 25996 4936 26036 4976
rect 29164 4936 29204 4976
rect 34156 4936 34196 4976
rect 38956 4936 38996 4976
rect 40300 4936 40340 4976
rect 44092 4936 44132 4976
rect 44332 4936 44372 4976
rect 44524 4936 44564 4976
rect 44908 4936 44948 4976
rect 45148 4936 45188 4976
rect 5452 4852 5492 4892
rect 5731 4852 5771 4892
rect 6412 4852 6452 4892
rect 6691 4852 6731 4892
rect 7564 4852 7604 4892
rect 8812 4852 8852 4892
rect 9283 4852 9323 4892
rect 9388 4852 9428 4892
rect 9868 4852 9908 4892
rect 10348 4852 10388 4892
rect 10867 4852 10907 4892
rect 12556 4852 12596 4892
rect 13804 4852 13844 4892
rect 15244 4852 15284 4892
rect 16492 4852 16532 4892
rect 17068 4852 17108 4892
rect 18316 4852 18356 4892
rect 21100 4852 21140 4892
rect 22356 4852 22396 4892
rect 22924 4852 22964 4892
rect 24172 4852 24212 4892
rect 33100 4852 33140 4892
rect 33379 4852 33419 4892
rect 34924 4852 34964 4892
rect 36172 4852 36212 4892
rect 37324 4852 37364 4892
rect 38572 4852 38612 4892
rect 40780 4852 40820 4892
rect 41059 4852 41099 4892
rect 1468 4768 1508 4808
rect 5836 4768 5876 4808
rect 6796 4768 6836 4808
rect 9004 4768 9044 4808
rect 14236 4768 14276 4808
rect 19996 4768 20036 4808
rect 29404 4768 29444 4808
rect 33484 4768 33524 4808
rect 33916 4768 33956 4808
rect 41164 4768 41204 4808
rect 1852 4684 1892 4724
rect 11020 4684 11060 4724
rect 12124 4684 12164 4724
rect 15052 4684 15092 4724
rect 18508 4684 18548 4724
rect 22540 4684 22580 4724
rect 24364 4684 24404 4724
rect 26236 4684 26276 4724
rect 38764 4684 38804 4724
rect 40540 4684 40580 4724
rect 42979 4684 43019 4724
rect 43267 4684 43307 4724
rect 43843 4684 43883 4724
rect 44764 4684 44804 4724
rect 4928 4516 4968 4556
rect 5010 4516 5050 4556
rect 5092 4516 5132 4556
rect 5174 4516 5214 4556
rect 5256 4516 5296 4556
rect 20048 4516 20088 4556
rect 20130 4516 20170 4556
rect 20212 4516 20252 4556
rect 20294 4516 20334 4556
rect 20376 4516 20416 4556
rect 35168 4516 35208 4556
rect 35250 4516 35290 4556
rect 35332 4516 35372 4556
rect 35414 4516 35454 4556
rect 35496 4516 35536 4556
rect 24028 4348 24068 4388
rect 42211 4348 42251 4388
rect 42499 4348 42539 4388
rect 42787 4348 42827 4388
rect 43555 4348 43595 4388
rect 44227 4348 44267 4388
rect 6220 4264 6260 4304
rect 8851 4264 8891 4304
rect 9244 4264 9284 4304
rect 9868 4264 9908 4304
rect 11260 4264 11300 4304
rect 13708 4264 13748 4304
rect 15244 4264 15284 4304
rect 18508 4264 18548 4304
rect 22348 4264 22388 4304
rect 31180 4264 31220 4304
rect 39340 4264 39380 4304
rect 43852 4264 43892 4304
rect 45148 4264 45188 4304
rect 4780 4180 4820 4220
rect 6028 4171 6068 4211
rect 7075 4180 7115 4220
rect 7180 4180 7220 4220
rect 7564 4180 7604 4220
rect 8140 4171 8180 4211
rect 8620 4171 8660 4211
rect 9484 4180 9524 4220
rect 9763 4180 9803 4220
rect 12268 4180 12308 4220
rect 13516 4171 13556 4211
rect 15373 4180 15413 4220
rect 15628 4180 15668 4220
rect 16876 4180 16916 4220
rect 18124 4171 18164 4211
rect 18700 4171 18740 4211
rect 19948 4180 19988 4220
rect 20908 4180 20948 4220
rect 22156 4171 22196 4211
rect 24364 4171 24404 4211
rect 25612 4180 25652 4220
rect 25996 4171 26036 4211
rect 27244 4180 27284 4220
rect 27628 4180 27668 4220
rect 28876 4171 28916 4211
rect 29740 4180 29780 4220
rect 30988 4171 31028 4211
rect 32611 4180 32651 4220
rect 32716 4180 32756 4220
rect 33093 4180 33133 4220
rect 33676 4171 33716 4211
rect 34156 4171 34196 4211
rect 37228 4180 37268 4220
rect 38476 4171 38516 4211
rect 38908 4180 38948 4220
rect 39235 4180 39275 4220
rect 40396 4171 40436 4211
rect 41644 4180 41684 4220
rect 43468 4180 43508 4220
rect 1228 4096 1268 4136
rect 1468 4096 1508 4136
rect 1612 4096 1652 4136
rect 4108 4096 4148 4136
rect 6412 4096 6452 4136
rect 7660 4096 7700 4136
rect 9004 4096 9044 4136
rect 10204 4096 10244 4136
rect 10348 4096 10388 4136
rect 11020 4096 11060 4136
rect 13948 4096 13988 4136
rect 14188 4096 14228 4136
rect 20140 4096 20180 4136
rect 20524 4096 20564 4136
rect 23788 4096 23828 4136
rect 29452 4096 29492 4136
rect 33196 4096 33236 4136
rect 34732 4096 34772 4136
rect 34924 4096 34964 4136
rect 35980 4096 36020 4136
rect 39772 4096 39812 4136
rect 40012 4096 40052 4136
rect 42028 4096 42068 4136
rect 43180 4096 43220 4136
rect 44524 4096 44564 4136
rect 44908 4096 44948 4136
rect 1852 4012 1892 4052
rect 18316 4012 18356 4052
rect 20380 4012 20420 4052
rect 20764 4012 20804 4052
rect 24172 4012 24212 4052
rect 34492 4012 34532 4052
rect 38668 4012 38708 4052
rect 39628 4012 39668 4052
rect 44764 4012 44804 4052
rect 4348 3928 4388 3968
rect 6652 3928 6692 3968
rect 10588 3928 10628 3968
rect 14956 3928 14996 3968
rect 25804 3928 25844 3968
rect 29068 3928 29108 3968
rect 29212 3928 29252 3968
rect 34387 3928 34427 3968
rect 35164 3928 35204 3968
rect 36220 3928 36260 3968
rect 40204 3928 40244 3968
rect 41788 3928 41828 3968
rect 3688 3760 3728 3800
rect 3770 3760 3810 3800
rect 3852 3760 3892 3800
rect 3934 3760 3974 3800
rect 4016 3760 4056 3800
rect 18808 3760 18848 3800
rect 18890 3760 18930 3800
rect 18972 3760 19012 3800
rect 19054 3760 19094 3800
rect 19136 3760 19176 3800
rect 33928 3760 33968 3800
rect 34010 3760 34050 3800
rect 34092 3760 34132 3800
rect 34174 3760 34214 3800
rect 34256 3760 34296 3800
rect 14620 3592 14660 3632
rect 43996 3592 44036 3632
rect 45148 3592 45188 3632
rect 1468 3508 1508 3548
rect 1852 3508 1892 3548
rect 5356 3508 5396 3548
rect 8140 3508 8180 3548
rect 8572 3508 8612 3548
rect 13804 3508 13844 3548
rect 14236 3508 14276 3548
rect 18988 3508 19028 3548
rect 24652 3508 24692 3548
rect 29548 3508 29588 3548
rect 31948 3508 31988 3548
rect 33484 3508 33524 3548
rect 1228 3424 1268 3464
rect 1612 3424 1652 3464
rect 8332 3424 8372 3464
rect 8716 3424 8756 3464
rect 13996 3424 14036 3464
rect 14860 3424 14900 3464
rect 15628 3424 15668 3464
rect 18028 3424 18068 3464
rect 19372 3424 19412 3464
rect 21004 3424 21044 3464
rect 24796 3424 24836 3464
rect 25036 3424 25076 3464
rect 25708 3424 25748 3464
rect 29788 3424 29828 3464
rect 30028 3424 30068 3464
rect 33868 3424 33908 3464
rect 38572 3424 38612 3464
rect 44236 3424 44276 3464
rect 44620 3424 44660 3464
rect 44908 3424 44948 3464
rect 3916 3340 3956 3380
rect 5164 3340 5204 3380
rect 7468 3340 7508 3380
rect 7747 3340 7787 3380
rect 11404 3340 11444 3380
rect 12652 3340 12692 3380
rect 13132 3340 13172 3380
rect 13411 3340 13451 3380
rect 15139 3340 15179 3380
rect 15244 3340 15284 3380
rect 15724 3340 15764 3380
rect 16204 3340 16244 3380
rect 16684 3373 16724 3413
rect 18316 3340 18356 3380
rect 18595 3340 18635 3380
rect 23980 3340 24020 3380
rect 24259 3340 24299 3380
rect 26380 3340 26420 3380
rect 27628 3340 27668 3380
rect 28876 3340 28916 3380
rect 29155 3340 29195 3380
rect 30508 3340 30548 3380
rect 31756 3340 31796 3380
rect 32812 3340 32852 3380
rect 33091 3340 33131 3380
rect 36172 3340 36212 3380
rect 37424 3340 37464 3380
rect 38083 3340 38123 3380
rect 38188 3340 38228 3380
rect 38668 3340 38708 3380
rect 39148 3340 39188 3380
rect 39667 3340 39707 3380
rect 41356 3340 41396 3380
rect 43756 3340 43796 3380
rect 7852 3256 7892 3296
rect 12844 3256 12884 3296
rect 13516 3256 13556 3296
rect 18700 3256 18740 3296
rect 19132 3256 19172 3296
rect 24364 3256 24404 3296
rect 29260 3256 29300 3296
rect 33180 3256 33220 3296
rect 33628 3256 33668 3296
rect 37612 3256 37652 3296
rect 44380 3256 44420 3296
rect 8956 3172 8996 3212
rect 16876 3172 16916 3212
rect 17788 3172 17828 3212
rect 21244 3172 21284 3212
rect 25468 3172 25508 3212
rect 27820 3172 27860 3212
rect 39820 3172 39860 3212
rect 41635 3172 41675 3212
rect 41923 3172 41963 3212
rect 42211 3172 42251 3212
rect 42499 3172 42539 3212
rect 42787 3172 42827 3212
rect 43075 3172 43115 3212
rect 43363 3172 43403 3212
rect 4928 3004 4968 3044
rect 5010 3004 5050 3044
rect 5092 3004 5132 3044
rect 5174 3004 5214 3044
rect 5256 3004 5296 3044
rect 20048 3004 20088 3044
rect 20130 3004 20170 3044
rect 20212 3004 20252 3044
rect 20294 3004 20334 3044
rect 20376 3004 20416 3044
rect 35168 3004 35208 3044
rect 35250 3004 35290 3044
rect 35332 3004 35372 3044
rect 35414 3004 35454 3044
rect 35496 3004 35536 3044
rect 5596 2836 5636 2876
rect 7180 2836 7220 2876
rect 9004 2836 9044 2876
rect 9628 2836 9668 2876
rect 11212 2836 11252 2876
rect 15436 2836 15476 2876
rect 20908 2836 20948 2876
rect 24844 2836 24884 2876
rect 27532 2836 27572 2876
rect 30028 2836 30068 2876
rect 34060 2836 34100 2876
rect 40771 2836 40811 2876
rect 41059 2836 41099 2876
rect 41308 2836 41348 2876
rect 41692 2836 41732 2876
rect 42460 2836 42500 2876
rect 43075 2836 43115 2876
rect 45148 2836 45188 2876
rect 1468 2752 1508 2792
rect 18604 2752 18644 2792
rect 22636 2752 22676 2792
rect 24988 2752 25028 2792
rect 30556 2752 30596 2792
rect 30988 2752 31028 2792
rect 35740 2752 35780 2792
rect 38092 2752 38132 2792
rect 38764 2752 38804 2792
rect 44764 2752 44804 2792
rect 5740 2668 5780 2708
rect 6988 2659 7028 2699
rect 7564 2668 7604 2708
rect 8812 2659 8852 2699
rect 9772 2668 9812 2708
rect 11020 2659 11060 2699
rect 11404 2668 11444 2708
rect 12652 2659 12692 2699
rect 13324 2668 13364 2708
rect 13453 2668 13493 2708
rect 13708 2668 13748 2708
rect 13996 2668 14036 2708
rect 15244 2659 15284 2699
rect 15715 2668 15755 2708
rect 15820 2668 15860 2708
rect 16204 2668 16244 2708
rect 16780 2659 16820 2699
rect 17260 2659 17300 2699
rect 18220 2668 18260 2708
rect 18499 2668 18539 2708
rect 19171 2668 19211 2708
rect 19276 2668 19316 2708
rect 19660 2668 19700 2708
rect 20236 2659 20276 2699
rect 20716 2659 20756 2699
rect 21196 2668 21236 2708
rect 22444 2659 22484 2699
rect 23107 2668 23147 2708
rect 23212 2668 23252 2708
rect 23596 2668 23636 2708
rect 24172 2659 24212 2699
rect 24652 2659 24692 2699
rect 25324 2668 25364 2708
rect 25453 2668 25493 2708
rect 25708 2668 25748 2708
rect 26092 2668 26132 2708
rect 27340 2659 27380 2699
rect 28291 2668 28331 2708
rect 28396 2668 28436 2708
rect 28780 2668 28820 2708
rect 29356 2659 29396 2699
rect 29836 2659 29876 2699
rect 31180 2659 31220 2699
rect 32428 2668 32468 2708
rect 32620 2668 32660 2708
rect 33868 2659 33908 2699
rect 34924 2668 34964 2708
rect 35179 2668 35219 2708
rect 35299 2668 35339 2708
rect 36652 2668 36692 2708
rect 37900 2659 37940 2699
rect 38380 2668 38420 2708
rect 38659 2668 38699 2708
rect 1228 2584 1268 2624
rect 1612 2584 1652 2624
rect 1996 2584 2036 2624
rect 5356 2584 5396 2624
rect 9388 2584 9428 2624
rect 16300 2584 16340 2624
rect 17740 2584 17780 2624
rect 19756 2584 19796 2624
rect 23692 2584 23732 2624
rect 27916 2584 27956 2624
rect 28876 2584 28916 2624
rect 30412 2584 30452 2624
rect 30796 2584 30836 2624
rect 35980 2584 36020 2624
rect 36268 2584 36308 2624
rect 39100 2584 39140 2624
rect 39436 2584 39476 2624
rect 41548 2584 41588 2624
rect 41932 2584 41972 2624
rect 42076 2584 42116 2624
rect 42316 2584 42356 2624
rect 42700 2584 42740 2624
rect 43084 2584 43124 2624
rect 43372 2584 43412 2624
rect 43756 2584 43796 2624
rect 44332 2584 44372 2624
rect 44524 2584 44564 2624
rect 44908 2584 44948 2624
rect 2236 2500 2276 2540
rect 27676 2500 27716 2540
rect 35596 2500 35636 2540
rect 43996 2500 44036 2540
rect 1852 2416 1892 2456
rect 12844 2416 12884 2456
rect 13036 2416 13076 2456
rect 17491 2416 17531 2456
rect 17980 2416 18020 2456
rect 18892 2416 18932 2456
rect 30172 2416 30212 2456
rect 36508 2416 36548 2456
rect 39196 2416 39236 2456
rect 43612 2416 43652 2456
rect 44092 2416 44132 2456
rect 3688 2248 3728 2288
rect 3770 2248 3810 2288
rect 3852 2248 3892 2288
rect 3934 2248 3974 2288
rect 4016 2248 4056 2288
rect 18808 2248 18848 2288
rect 18890 2248 18930 2288
rect 18972 2248 19012 2288
rect 19054 2248 19094 2288
rect 19136 2248 19176 2288
rect 33928 2248 33968 2288
rect 34010 2248 34050 2288
rect 34092 2248 34132 2288
rect 34174 2248 34214 2288
rect 34256 2248 34296 2288
rect 1852 2080 1892 2120
rect 2620 2080 2660 2120
rect 4252 2080 4292 2120
rect 5980 2080 6020 2120
rect 8764 2080 8804 2120
rect 9148 2080 9188 2120
rect 10732 2080 10772 2120
rect 13948 2080 13988 2120
rect 16540 2080 16580 2120
rect 16972 2080 17012 2120
rect 20620 2080 20660 2120
rect 34252 2080 34292 2120
rect 35164 2080 35204 2120
rect 36988 2080 37028 2120
rect 39004 2080 39044 2120
rect 40444 2080 40484 2120
rect 41884 2080 41924 2120
rect 42844 2080 42884 2120
rect 3484 1996 3524 2036
rect 4828 1996 4868 2036
rect 12220 1996 12260 2036
rect 13804 1996 13844 2036
rect 14620 1996 14660 2036
rect 24652 1996 24692 2036
rect 25180 1996 25220 2036
rect 28684 1996 28724 2036
rect 31612 1996 31652 2036
rect 45148 1996 45188 2036
rect 1228 1912 1268 1952
rect 1612 1912 1652 1952
rect 1996 1912 2036 1952
rect 2380 1912 2420 1952
rect 3244 1912 3284 1952
rect 4012 1912 4052 1952
rect 4588 1912 4628 1952
rect 4972 1912 5012 1952
rect 5212 1912 5252 1952
rect 5395 1912 5435 1952
rect 5740 1912 5780 1952
rect 6124 1912 6164 1952
rect 6508 1912 6548 1952
rect 8524 1912 8564 1952
rect 8908 1912 8948 1952
rect 10924 1912 10964 1952
rect 11500 1912 11540 1952
rect 11884 1912 11924 1952
rect 12460 1912 12500 1952
rect 12604 1912 12644 1952
rect 12844 1912 12884 1952
rect 14188 1912 14228 1952
rect 14380 1912 14420 1952
rect 14764 1912 14804 1952
rect 15004 1912 15044 1952
rect 15628 1912 15668 1952
rect 15820 1912 15860 1952
rect 16204 1912 16244 1952
rect 16780 1912 16820 1952
rect 18604 1912 18644 1952
rect 18988 1912 19028 1952
rect 19564 1912 19604 1952
rect 19852 1912 19892 1952
rect 20236 1912 20276 1952
rect 22636 1912 22676 1952
rect 23251 1912 23291 1952
rect 23500 1912 23540 1952
rect 24796 1912 24836 1952
rect 25036 1912 25076 1952
rect 25420 1912 25460 1952
rect 25804 1912 25844 1952
rect 30028 1912 30068 1952
rect 31372 1912 31412 1952
rect 31852 1912 31892 1952
rect 32092 1912 32132 1952
rect 34924 1912 34964 1952
rect 36748 1912 36788 1952
rect 39244 1912 39284 1952
rect 40300 1912 40340 1952
rect 40684 1912 40724 1952
rect 42124 1912 42164 1952
rect 42604 1912 42644 1952
rect 42988 1912 43028 1952
rect 43372 1912 43412 1952
rect 43756 1912 43796 1952
rect 44092 1912 44132 1952
rect 44332 1912 44372 1952
rect 44716 1912 44756 1952
rect 44908 1912 44948 1952
rect 6892 1828 6932 1868
rect 8140 1828 8180 1868
rect 9292 1828 9332 1868
rect 10540 1828 10580 1868
rect 13132 1828 13172 1868
rect 13411 1828 13451 1868
rect 17164 1828 17204 1868
rect 18412 1828 18452 1868
rect 20812 1828 20852 1868
rect 22060 1828 22100 1868
rect 23980 1828 24020 1868
rect 24235 1828 24275 1868
rect 24355 1828 24395 1868
rect 25996 1828 26036 1868
rect 27244 1828 27284 1868
rect 28012 1828 28052 1868
rect 28291 1828 28331 1868
rect 28972 1828 29012 1868
rect 29251 1828 29291 1868
rect 29692 1828 29732 1868
rect 32812 1828 32852 1868
rect 34060 1828 34100 1868
rect 1468 1744 1508 1784
rect 11740 1744 11780 1784
rect 12124 1744 12164 1784
rect 13516 1744 13556 1784
rect 16444 1744 16484 1784
rect 19228 1744 19268 1784
rect 25564 1744 25604 1784
rect 27436 1744 27476 1784
rect 28396 1744 28436 1784
rect 29356 1744 29396 1784
rect 42412 1744 42452 1784
rect 43996 1744 44036 1784
rect 2236 1660 2276 1700
rect 5596 1660 5636 1700
rect 6364 1660 6404 1700
rect 6748 1660 6788 1700
rect 8332 1660 8372 1700
rect 11164 1660 11204 1700
rect 15388 1660 15428 1700
rect 16060 1660 16100 1700
rect 18844 1660 18884 1700
rect 19324 1660 19364 1700
rect 20092 1660 20132 1700
rect 20476 1660 20516 1700
rect 22396 1660 22436 1700
rect 23068 1660 23108 1700
rect 23740 1660 23780 1700
rect 29788 1660 29828 1700
rect 40291 1660 40331 1700
rect 41068 1660 41108 1700
rect 41356 1660 41396 1700
rect 41644 1660 41684 1700
rect 42316 1660 42356 1700
rect 43228 1660 43268 1700
rect 43612 1660 43652 1700
rect 4928 1492 4968 1532
rect 5010 1492 5050 1532
rect 5092 1492 5132 1532
rect 5174 1492 5214 1532
rect 5256 1492 5296 1532
rect 20048 1492 20088 1532
rect 20130 1492 20170 1532
rect 20212 1492 20252 1532
rect 20294 1492 20334 1532
rect 20376 1492 20416 1532
rect 35168 1492 35208 1532
rect 35250 1492 35290 1532
rect 35332 1492 35372 1532
rect 35414 1492 35454 1532
rect 35496 1492 35536 1532
<< metal2 >>
rect 19939 11068 19948 11108
rect 19988 11068 21196 11108
rect 21236 11068 21245 11108
rect 0 11024 90 11044
rect 46278 11024 46368 11044
rect 0 10984 1324 11024
rect 1364 10984 1373 11024
rect 44707 10984 44716 11024
rect 44756 10984 46368 11024
rect 0 10964 90 10984
rect 46278 10964 46368 10984
rect 18403 10900 18412 10940
rect 18452 10900 21004 10940
rect 21044 10900 21053 10940
rect 28675 10732 28684 10772
rect 28724 10732 32332 10772
rect 32372 10732 32381 10772
rect 0 10688 90 10708
rect 46278 10688 46368 10708
rect 0 10648 1132 10688
rect 1172 10648 1181 10688
rect 44227 10648 44236 10688
rect 44276 10648 46368 10688
rect 0 10628 90 10648
rect 46278 10628 46368 10648
rect 0 10352 90 10372
rect 46278 10352 46368 10372
rect 0 10312 1420 10352
rect 1460 10312 1469 10352
rect 34435 10312 34444 10352
rect 34484 10312 39148 10352
rect 39188 10312 39197 10352
rect 43267 10312 43276 10352
rect 43316 10312 46368 10352
rect 0 10292 90 10312
rect 46278 10292 46368 10312
rect 30595 10228 30604 10268
rect 30644 10228 34924 10268
rect 34964 10228 34973 10268
rect 12940 10144 17644 10184
rect 17684 10144 17693 10184
rect 18211 10144 18220 10184
rect 18260 10144 18836 10184
rect 12940 10100 12980 10144
rect 18796 10100 18836 10144
rect 21580 10144 22868 10184
rect 21580 10100 21620 10144
rect 22828 10100 22868 10144
rect 23020 10144 23404 10184
rect 23444 10144 23453 10184
rect 24556 10144 28724 10184
rect 23020 10100 23060 10144
rect 24556 10100 24596 10144
rect 28684 10100 28724 10144
rect 3427 10060 3436 10100
rect 3476 10060 12980 10100
rect 13036 10060 15820 10100
rect 15860 10060 15869 10100
rect 16291 10060 16300 10100
rect 16340 10060 18604 10100
rect 18644 10060 18653 10100
rect 18796 10060 21004 10100
rect 21044 10060 21053 10100
rect 21475 10060 21484 10100
rect 21524 10060 21620 10100
rect 21667 10060 21676 10100
rect 21716 10060 22732 10100
rect 22772 10060 22781 10100
rect 22828 10060 23060 10100
rect 23116 10060 24596 10100
rect 24643 10060 24652 10100
rect 24692 10060 25804 10100
rect 25844 10060 25853 10100
rect 28684 10060 29548 10100
rect 29588 10060 29597 10100
rect 31747 10060 31756 10100
rect 31796 10060 36460 10100
rect 36500 10060 36509 10100
rect 36643 10060 36652 10100
rect 36692 10060 41452 10100
rect 41492 10060 41501 10100
rect 0 10016 90 10036
rect 13036 10016 13076 10060
rect 23116 10016 23156 10060
rect 46278 10016 46368 10036
rect 0 9976 1268 10016
rect 2275 9976 2284 10016
rect 2324 9976 12652 10016
rect 12692 9976 12701 10016
rect 12835 9976 12844 10016
rect 12884 9976 13076 10016
rect 13411 9976 13420 10016
rect 13460 9976 23156 10016
rect 23203 9976 23212 10016
rect 23252 9976 33140 10016
rect 33859 9976 33868 10016
rect 33908 9976 37900 10016
rect 37940 9976 37949 10016
rect 38659 9976 38668 10016
rect 38708 9976 42220 10016
rect 42260 9976 42269 10016
rect 44419 9976 44428 10016
rect 44468 9976 46368 10016
rect 0 9956 90 9976
rect 1228 9848 1268 9976
rect 33100 9932 33140 9976
rect 46278 9956 46368 9976
rect 1315 9892 1324 9932
rect 1364 9892 2900 9932
rect 8227 9892 8236 9932
rect 8276 9892 11788 9932
rect 11828 9892 11837 9932
rect 12067 9892 12076 9932
rect 12116 9892 15052 9932
rect 15092 9892 15101 9932
rect 15244 9892 21292 9932
rect 21332 9892 21341 9932
rect 29635 9892 29644 9932
rect 29684 9892 31468 9932
rect 31508 9892 31517 9932
rect 33100 9892 33772 9932
rect 33812 9892 33821 9932
rect 38179 9892 38188 9932
rect 38228 9892 41068 9932
rect 41108 9892 41117 9932
rect 41539 9892 41548 9932
rect 41588 9892 45140 9932
rect 1228 9808 2420 9848
rect 0 9680 90 9700
rect 0 9640 2036 9680
rect 0 9620 90 9640
rect 1411 9556 1420 9596
rect 1460 9556 1748 9596
rect 1097 9472 1228 9512
rect 1268 9472 1277 9512
rect 1603 9472 1612 9512
rect 1652 9472 1661 9512
rect 0 9344 90 9364
rect 1612 9344 1652 9472
rect 1708 9428 1748 9556
rect 1996 9512 2036 9640
rect 2380 9512 2420 9808
rect 2860 9512 2900 9892
rect 3679 9808 3688 9848
rect 3728 9808 3770 9848
rect 3810 9808 3852 9848
rect 3892 9808 3934 9848
rect 3974 9808 4016 9848
rect 4056 9808 4065 9848
rect 5644 9808 10924 9848
rect 10964 9808 10973 9848
rect 11020 9808 13324 9848
rect 13364 9808 13373 9848
rect 3379 9640 3388 9680
rect 3428 9640 3436 9680
rect 3476 9640 3559 9680
rect 1987 9472 1996 9512
rect 2036 9472 2045 9512
rect 2371 9472 2380 9512
rect 2420 9472 2429 9512
rect 2755 9472 2764 9512
rect 2804 9472 2813 9512
rect 2860 9472 3148 9512
rect 3188 9472 3197 9512
rect 2764 9428 2804 9472
rect 1708 9388 2804 9428
rect 5644 9344 5684 9808
rect 11020 9764 11060 9808
rect 15244 9764 15284 9892
rect 15811 9808 15820 9848
rect 15860 9808 18220 9848
rect 18260 9808 18269 9848
rect 18799 9808 18808 9848
rect 18848 9808 18890 9848
rect 18930 9808 18972 9848
rect 19012 9808 19054 9848
rect 19094 9808 19136 9848
rect 19176 9808 19185 9848
rect 19267 9808 19276 9848
rect 19316 9808 20044 9848
rect 20084 9808 20093 9848
rect 22252 9808 23116 9848
rect 23156 9808 23165 9848
rect 28579 9808 28588 9848
rect 28628 9808 33388 9848
rect 33428 9808 33437 9848
rect 33919 9808 33928 9848
rect 33968 9808 34010 9848
rect 34050 9808 34092 9848
rect 34132 9808 34174 9848
rect 34214 9808 34256 9848
rect 34296 9808 34305 9848
rect 39043 9808 39052 9848
rect 39092 9808 44140 9848
rect 44180 9808 44189 9848
rect 6211 9724 6220 9764
rect 6260 9724 9964 9764
rect 10004 9724 10013 9764
rect 10060 9724 11060 9764
rect 11116 9724 15284 9764
rect 15340 9724 17548 9764
rect 17588 9724 17597 9764
rect 17644 9724 19372 9764
rect 19412 9724 19421 9764
rect 10060 9680 10100 9724
rect 11116 9680 11156 9724
rect 15340 9680 15380 9724
rect 17644 9680 17684 9724
rect 8105 9640 8188 9680
rect 8228 9640 8236 9680
rect 8276 9640 8285 9680
rect 9907 9640 9916 9680
rect 9956 9640 10100 9680
rect 10243 9640 10252 9680
rect 10292 9640 11156 9680
rect 11539 9640 11548 9680
rect 11588 9640 12076 9680
rect 12116 9640 12125 9680
rect 12307 9640 12316 9680
rect 12356 9640 12844 9680
rect 12884 9640 12893 9680
rect 14515 9640 14524 9680
rect 14564 9640 15380 9680
rect 15427 9640 15436 9680
rect 15476 9640 15485 9680
rect 15667 9640 15676 9680
rect 15716 9640 17684 9680
rect 18067 9640 18076 9680
rect 18116 9640 20620 9680
rect 20660 9640 20669 9680
rect 21100 9640 21580 9680
rect 21620 9640 21629 9680
rect 21929 9640 22012 9680
rect 22052 9640 22060 9680
rect 22100 9640 22109 9680
rect 15436 9596 15476 9640
rect 7660 9556 8084 9596
rect 8131 9556 8140 9596
rect 8180 9556 8332 9596
rect 8372 9556 8381 9596
rect 8428 9556 9428 9596
rect 9523 9556 9532 9596
rect 9572 9556 9812 9596
rect 9929 9556 10060 9596
rect 10100 9556 10109 9596
rect 11923 9556 11932 9596
rect 11972 9556 15476 9596
rect 16492 9556 18124 9596
rect 18164 9556 18173 9596
rect 18796 9556 19948 9596
rect 19988 9556 19997 9596
rect 20131 9556 20140 9596
rect 20180 9556 20716 9596
rect 20756 9556 20765 9596
rect 7660 9512 7700 9556
rect 8044 9512 8084 9556
rect 8428 9512 8468 9556
rect 9388 9512 9428 9556
rect 9772 9512 9812 9556
rect 5731 9472 5740 9512
rect 5780 9472 7700 9512
rect 7817 9472 7948 9512
rect 7988 9472 7997 9512
rect 8044 9472 8468 9512
rect 8620 9472 8812 9512
rect 8852 9472 8861 9512
rect 9161 9472 9292 9512
rect 9332 9472 9341 9512
rect 9388 9472 9620 9512
rect 9667 9472 9676 9512
rect 9716 9472 9725 9512
rect 9772 9472 11252 9512
rect 11299 9472 11308 9512
rect 11348 9472 11479 9512
rect 11683 9472 11692 9512
rect 11732 9472 11884 9512
rect 11924 9472 11933 9512
rect 12067 9472 12076 9512
rect 12116 9472 12268 9512
rect 12308 9472 12317 9512
rect 13411 9472 13420 9512
rect 13460 9472 14284 9512
rect 14324 9472 14333 9512
rect 14659 9472 14668 9512
rect 14708 9472 14764 9512
rect 14804 9472 14839 9512
rect 15043 9472 15052 9512
rect 15092 9472 15101 9512
rect 15305 9472 15436 9512
rect 15476 9472 15485 9512
rect 15689 9472 15820 9512
rect 15860 9472 15869 9512
rect 15916 9472 16204 9512
rect 16244 9472 16253 9512
rect 7564 9428 7604 9472
rect 8620 9428 8660 9472
rect 5827 9388 5836 9428
rect 5876 9388 6316 9428
rect 6356 9388 6365 9428
rect 7564 9379 7604 9388
rect 7660 9388 8660 9428
rect 8716 9419 8756 9428
rect 0 9304 1652 9344
rect 1708 9304 5684 9344
rect 0 9284 90 9304
rect 1708 9260 1748 9304
rect 1459 9220 1468 9260
rect 1508 9220 1748 9260
rect 1843 9220 1852 9260
rect 1892 9220 1901 9260
rect 2227 9220 2236 9260
rect 2276 9220 2516 9260
rect 2611 9220 2620 9260
rect 2660 9220 2860 9260
rect 2900 9220 2909 9260
rect 2995 9220 3004 9260
rect 3044 9220 4204 9260
rect 4244 9220 4253 9260
rect 1852 9092 1892 9220
rect 2476 9176 2516 9220
rect 7660 9176 7700 9388
rect 8873 9388 9004 9428
rect 9044 9388 9053 9428
rect 8716 9344 8756 9379
rect 9580 9344 9620 9472
rect 9676 9428 9716 9472
rect 11212 9428 11252 9472
rect 12652 9428 12692 9437
rect 15052 9428 15092 9472
rect 15916 9428 15956 9472
rect 9676 9388 10252 9428
rect 10292 9388 10301 9428
rect 10444 9419 10676 9428
rect 10484 9388 10676 9419
rect 10723 9388 10732 9428
rect 10772 9388 10781 9428
rect 11212 9388 12596 9428
rect 12643 9388 12652 9428
rect 12692 9388 12823 9428
rect 13891 9388 13900 9428
rect 13940 9388 13949 9428
rect 14275 9388 14284 9428
rect 14324 9388 15092 9428
rect 15139 9388 15148 9428
rect 15188 9388 15956 9428
rect 16099 9388 16108 9428
rect 16148 9388 16204 9428
rect 16244 9388 16279 9428
rect 10444 9370 10484 9379
rect 10636 9344 10676 9388
rect 10732 9344 10772 9388
rect 8489 9304 8620 9344
rect 8660 9304 8669 9344
rect 8716 9304 9484 9344
rect 9524 9304 9533 9344
rect 9580 9304 9964 9344
rect 10004 9304 10013 9344
rect 10217 9304 10348 9344
rect 10388 9304 10397 9344
rect 10627 9304 10636 9344
rect 10676 9304 10685 9344
rect 10732 9304 12460 9344
rect 12500 9304 12509 9344
rect 12556 9260 12596 9388
rect 12652 9379 12692 9388
rect 13900 9344 13940 9388
rect 16492 9344 16532 9556
rect 18796 9512 18836 9556
rect 21100 9512 21140 9640
rect 21196 9556 21676 9596
rect 21716 9556 21725 9596
rect 21859 9556 21868 9596
rect 21908 9556 22108 9596
rect 22148 9556 22157 9596
rect 21196 9512 21236 9556
rect 22252 9512 22292 9808
rect 22924 9724 23308 9764
rect 23348 9724 23357 9764
rect 27043 9724 27052 9764
rect 27092 9724 30260 9764
rect 32131 9724 32140 9764
rect 32180 9724 35780 9764
rect 22924 9596 22964 9724
rect 30220 9680 30260 9724
rect 35740 9680 35780 9724
rect 22348 9556 22964 9596
rect 23020 9640 23500 9680
rect 23540 9640 23549 9680
rect 24739 9640 24748 9680
rect 24788 9640 25132 9680
rect 25172 9640 28444 9680
rect 28484 9640 28493 9680
rect 29059 9640 29068 9680
rect 29108 9640 29212 9680
rect 29252 9640 29261 9680
rect 30220 9640 32284 9680
rect 32324 9640 32333 9680
rect 33475 9640 33484 9680
rect 33524 9640 34444 9680
rect 34484 9640 34493 9680
rect 35740 9640 36892 9680
rect 36932 9640 36941 9680
rect 37219 9640 37228 9680
rect 37268 9640 37276 9680
rect 37316 9640 37399 9680
rect 38755 9640 38764 9680
rect 38804 9640 38812 9680
rect 38852 9640 38935 9680
rect 39139 9640 39148 9680
rect 39188 9640 39196 9680
rect 39236 9640 39319 9680
rect 43219 9640 43228 9680
rect 43268 9640 43276 9680
rect 43316 9640 43399 9680
rect 44297 9640 44380 9680
rect 44420 9640 44428 9680
rect 44468 9640 44477 9680
rect 22348 9512 22388 9556
rect 23020 9512 23060 9640
rect 23116 9556 23692 9596
rect 23732 9556 23741 9596
rect 23884 9556 24076 9596
rect 24116 9556 24125 9596
rect 24835 9556 24844 9596
rect 24884 9556 25028 9596
rect 25219 9556 25228 9596
rect 25268 9556 26612 9596
rect 27523 9556 27532 9596
rect 27572 9556 30644 9596
rect 30691 9556 30700 9596
rect 30740 9556 31412 9596
rect 31459 9556 31468 9596
rect 31508 9556 31604 9596
rect 31651 9556 31660 9596
rect 31700 9556 31709 9596
rect 31795 9556 31804 9596
rect 31844 9556 33140 9596
rect 33763 9556 33772 9596
rect 33812 9556 34300 9596
rect 34340 9556 34349 9596
rect 35465 9556 35596 9596
rect 35636 9556 35645 9596
rect 35971 9556 35980 9596
rect 36020 9556 36067 9596
rect 36115 9556 36124 9596
rect 36164 9556 36172 9596
rect 36212 9556 36295 9596
rect 36451 9556 36460 9596
rect 36500 9556 36508 9596
rect 36548 9556 36631 9596
rect 36748 9556 38996 9596
rect 39331 9556 39340 9596
rect 39380 9556 44564 9596
rect 23116 9512 23156 9556
rect 23884 9512 23924 9556
rect 17539 9472 17548 9512
rect 17588 9472 17836 9512
rect 17876 9472 17885 9512
rect 18787 9472 18796 9512
rect 18836 9472 18845 9512
rect 18979 9472 18988 9512
rect 19028 9472 20140 9512
rect 20180 9472 20189 9512
rect 20611 9472 20620 9512
rect 20660 9472 21140 9512
rect 21187 9472 21196 9512
rect 21236 9472 21245 9512
rect 21292 9472 21340 9512
rect 21380 9472 21389 9512
rect 21571 9472 21580 9512
rect 21620 9472 21629 9512
rect 21763 9472 21772 9512
rect 21812 9472 22292 9512
rect 22339 9472 22348 9512
rect 22388 9472 22397 9512
rect 22723 9472 22732 9512
rect 22772 9472 23060 9512
rect 23107 9472 23116 9512
rect 23156 9472 23165 9512
rect 23299 9472 23308 9512
rect 23348 9472 23357 9512
rect 23875 9472 23884 9512
rect 23924 9472 23933 9512
rect 24137 9472 24268 9512
rect 24308 9472 24317 9512
rect 17452 9428 17492 9437
rect 21292 9428 21332 9472
rect 21580 9428 21620 9472
rect 23308 9428 23348 9472
rect 24988 9428 25028 9556
rect 26572 9512 26612 9556
rect 30604 9512 30644 9556
rect 31372 9512 31412 9556
rect 31564 9512 31604 9556
rect 31660 9512 31700 9556
rect 33100 9512 33140 9556
rect 35980 9512 36020 9556
rect 36748 9512 36788 9556
rect 25219 9472 25228 9512
rect 25268 9472 25612 9512
rect 25652 9472 25661 9512
rect 25795 9472 25804 9512
rect 25844 9472 25975 9512
rect 26179 9472 26188 9512
rect 26228 9472 26237 9512
rect 26572 9472 27916 9512
rect 27956 9472 27965 9512
rect 28169 9472 28300 9512
rect 28340 9472 28349 9512
rect 28553 9472 28684 9512
rect 28724 9472 28733 9512
rect 28867 9472 28876 9512
rect 28916 9472 29068 9512
rect 29108 9472 29117 9512
rect 29321 9472 29452 9512
rect 29492 9472 29501 9512
rect 29705 9472 29836 9512
rect 29876 9472 29885 9512
rect 30019 9472 30028 9512
rect 30068 9472 30077 9512
rect 30595 9472 30604 9512
rect 30644 9472 30653 9512
rect 30979 9472 30988 9512
rect 31028 9472 31037 9512
rect 31363 9472 31372 9512
rect 31412 9472 31421 9512
rect 31555 9472 31564 9512
rect 31604 9472 31613 9512
rect 31660 9472 32140 9512
rect 32180 9472 32189 9512
rect 32323 9472 32332 9512
rect 32372 9472 32524 9512
rect 32564 9472 32573 9512
rect 32707 9472 32716 9512
rect 32756 9472 33044 9512
rect 33100 9472 33868 9512
rect 33908 9472 33917 9512
rect 34409 9472 34540 9512
rect 34580 9472 34589 9512
rect 34924 9472 35924 9512
rect 35971 9472 35980 9512
rect 36020 9472 36029 9512
rect 36355 9472 36364 9512
rect 36404 9472 36413 9512
rect 36739 9472 36748 9512
rect 36788 9472 36797 9512
rect 37123 9472 37132 9512
rect 37172 9472 37228 9512
rect 37268 9472 37303 9512
rect 37507 9472 37516 9512
rect 37556 9472 37565 9512
rect 37699 9472 37708 9512
rect 37748 9472 37900 9512
rect 37940 9472 37949 9512
rect 38275 9472 38284 9512
rect 38324 9472 38333 9512
rect 38537 9472 38668 9512
rect 38708 9472 38717 9512
rect 26188 9428 26228 9472
rect 30028 9428 30068 9472
rect 30988 9428 31028 9472
rect 33004 9428 33044 9472
rect 33964 9428 34004 9437
rect 34924 9428 34964 9472
rect 35884 9428 35924 9472
rect 36364 9428 36404 9472
rect 37516 9428 37556 9472
rect 38284 9428 38324 9472
rect 38956 9428 38996 9556
rect 44524 9512 44564 9556
rect 45100 9512 45140 9892
rect 46278 9680 46368 9700
rect 45187 9640 45196 9680
rect 45236 9640 46368 9680
rect 46278 9620 46368 9640
rect 39043 9472 39052 9512
rect 39092 9472 39223 9512
rect 39427 9472 39436 9512
rect 39476 9472 39764 9512
rect 39811 9472 39820 9512
rect 39860 9472 41020 9512
rect 41060 9472 41069 9512
rect 41251 9472 41260 9512
rect 41300 9472 42316 9512
rect 42356 9472 42365 9512
rect 42473 9472 42604 9512
rect 42644 9472 42653 9512
rect 42979 9472 42988 9512
rect 43028 9472 43037 9512
rect 43459 9472 43468 9512
rect 43508 9472 43756 9512
rect 43796 9472 43805 9512
rect 44131 9472 44140 9512
rect 44180 9472 44189 9512
rect 44515 9472 44524 9512
rect 44564 9472 44573 9512
rect 45091 9472 45100 9512
rect 45140 9472 45149 9512
rect 17492 9388 17836 9428
rect 17876 9388 17885 9428
rect 18787 9388 18796 9428
rect 18836 9388 19468 9428
rect 19508 9388 19517 9428
rect 19738 9388 19747 9428
rect 19787 9388 19796 9428
rect 19843 9388 19852 9428
rect 19892 9388 20908 9428
rect 20948 9388 20957 9428
rect 21283 9388 21292 9428
rect 21332 9388 21341 9428
rect 21580 9388 22924 9428
rect 22964 9388 22973 9428
rect 23308 9388 23884 9428
rect 23924 9388 23933 9428
rect 24425 9388 24556 9428
rect 24596 9388 24605 9428
rect 24739 9388 24748 9428
rect 24788 9388 24835 9428
rect 24875 9388 24919 9428
rect 24988 9388 26228 9428
rect 26851 9388 26860 9428
rect 26900 9388 26909 9428
rect 26993 9388 27052 9428
rect 27092 9388 27115 9428
rect 27155 9388 27173 9428
rect 27226 9388 27235 9428
rect 27275 9388 27436 9428
rect 27476 9388 27485 9428
rect 27619 9388 27628 9428
rect 27668 9388 30068 9428
rect 30115 9388 30124 9428
rect 30164 9388 31028 9428
rect 32419 9388 32428 9428
rect 32468 9388 32716 9428
rect 32756 9388 32812 9428
rect 32852 9388 32916 9428
rect 33004 9388 33964 9428
rect 34915 9388 34924 9428
rect 34964 9388 34973 9428
rect 35194 9388 35203 9428
rect 35243 9388 35252 9428
rect 35884 9388 35980 9428
rect 36020 9388 36029 9428
rect 36364 9388 37420 9428
rect 37460 9388 37469 9428
rect 37516 9388 38188 9428
rect 38228 9388 38237 9428
rect 38284 9388 38900 9428
rect 38956 9388 39628 9428
rect 39668 9388 39677 9428
rect 17452 9379 17492 9388
rect 13900 9304 14188 9344
rect 14228 9304 14237 9344
rect 14899 9304 14908 9344
rect 14948 9304 16532 9344
rect 17548 9304 19372 9344
rect 19412 9304 19421 9344
rect 17548 9260 17588 9304
rect 19756 9260 19796 9388
rect 19852 9344 19892 9388
rect 26860 9344 26900 9388
rect 33964 9379 34004 9388
rect 35212 9344 35252 9388
rect 19843 9304 19852 9344
rect 19892 9304 19968 9344
rect 20851 9304 20860 9344
rect 20900 9304 22444 9344
rect 22484 9304 22493 9344
rect 23539 9304 23548 9344
rect 23588 9304 24308 9344
rect 24809 9304 24940 9344
rect 24980 9304 24989 9344
rect 26860 9304 29068 9344
rect 29108 9304 29117 9344
rect 29539 9304 29548 9344
rect 29588 9304 29596 9344
rect 29636 9304 29719 9344
rect 30108 9304 30220 9344
rect 30260 9304 30268 9344
rect 30308 9304 33140 9344
rect 7747 9220 7756 9260
rect 7796 9220 7805 9260
rect 8035 9220 8044 9260
rect 8084 9220 10444 9260
rect 10484 9220 10493 9260
rect 12556 9220 13132 9260
rect 13172 9220 13181 9260
rect 15283 9220 15292 9260
rect 15332 9220 15572 9260
rect 16051 9220 16060 9260
rect 16100 9220 17588 9260
rect 17635 9220 17644 9260
rect 17684 9220 18124 9260
rect 18164 9220 18173 9260
rect 18281 9220 18412 9260
rect 18452 9220 18461 9260
rect 18547 9220 18556 9260
rect 18596 9220 18604 9260
rect 18644 9220 18727 9260
rect 19097 9220 19180 9260
rect 19220 9220 19228 9260
rect 19268 9220 19277 9260
rect 19747 9220 19756 9260
rect 19796 9220 19805 9260
rect 20035 9220 20044 9260
rect 20084 9220 20900 9260
rect 20947 9220 20956 9260
rect 20996 9220 21292 9260
rect 21332 9220 21341 9260
rect 22339 9220 22348 9260
rect 22388 9220 22492 9260
rect 22532 9220 22541 9260
rect 22627 9220 22636 9260
rect 22676 9220 22876 9260
rect 22916 9220 22925 9260
rect 23561 9220 23644 9260
rect 23684 9220 23692 9260
rect 23732 9220 23741 9260
rect 23875 9220 23884 9260
rect 23924 9220 24028 9260
rect 24068 9220 24077 9260
rect 2476 9136 7700 9176
rect 7756 9092 7796 9220
rect 15532 9176 15572 9220
rect 9571 9136 9580 9176
rect 9620 9136 10636 9176
rect 10676 9136 10685 9176
rect 13795 9136 13804 9176
rect 13844 9136 15148 9176
rect 15188 9136 15197 9176
rect 15532 9136 18508 9176
rect 18548 9136 18557 9176
rect 19948 9136 20620 9176
rect 20660 9136 20669 9176
rect 19948 9092 19988 9136
rect 20860 9092 20900 9220
rect 24268 9176 24308 9304
rect 33100 9260 33140 9304
rect 34060 9304 35252 9344
rect 35299 9304 35308 9344
rect 35348 9304 35479 9344
rect 35596 9304 38764 9344
rect 38804 9304 38813 9344
rect 34060 9260 34100 9304
rect 35596 9260 35636 9304
rect 38860 9260 38900 9388
rect 39724 9344 39764 9472
rect 42988 9428 43028 9472
rect 41347 9388 41356 9428
rect 41396 9388 43028 9428
rect 44140 9344 44180 9472
rect 38947 9304 38956 9344
rect 38996 9304 39580 9344
rect 39620 9304 39629 9344
rect 39724 9304 42028 9344
rect 42068 9304 42077 9344
rect 42403 9304 42412 9344
rect 42452 9304 44180 9344
rect 44236 9388 45188 9428
rect 44236 9260 44276 9388
rect 45148 9344 45188 9388
rect 46278 9344 46368 9364
rect 44755 9304 44764 9344
rect 44804 9304 45004 9344
rect 45044 9304 45053 9344
rect 45148 9304 46368 9344
rect 46278 9284 46368 9304
rect 24451 9220 24460 9260
rect 24500 9220 25372 9260
rect 25412 9220 25421 9260
rect 25516 9220 25900 9260
rect 25940 9220 25949 9260
rect 26035 9220 26044 9260
rect 26084 9220 26092 9260
rect 26132 9220 26215 9260
rect 26275 9220 26284 9260
rect 26324 9220 26428 9260
rect 26468 9220 26477 9260
rect 27331 9220 27340 9260
rect 27380 9220 27676 9260
rect 27716 9220 27725 9260
rect 27811 9220 27820 9260
rect 27860 9220 28060 9260
rect 28100 9220 28109 9260
rect 28697 9220 28780 9260
rect 28820 9220 28828 9260
rect 28868 9220 28877 9260
rect 30233 9220 30316 9260
rect 30356 9220 30364 9260
rect 30404 9220 30413 9260
rect 30595 9220 30604 9260
rect 30644 9220 30748 9260
rect 30788 9220 30797 9260
rect 31123 9220 31132 9260
rect 31172 9220 31276 9260
rect 31316 9220 31325 9260
rect 31891 9220 31900 9260
rect 31940 9220 32044 9260
rect 32084 9220 32093 9260
rect 33100 9220 34100 9260
rect 34147 9220 34156 9260
rect 34196 9220 34327 9260
rect 34819 9220 34828 9260
rect 34868 9220 35636 9260
rect 35731 9220 35740 9260
rect 35780 9220 35884 9260
rect 35924 9220 35933 9260
rect 37507 9220 37516 9260
rect 37556 9220 37660 9260
rect 37700 9220 37709 9260
rect 37795 9220 37804 9260
rect 37844 9220 38044 9260
rect 38084 9220 38093 9260
rect 38179 9220 38188 9260
rect 38228 9220 38428 9260
rect 38468 9220 38477 9260
rect 38860 9220 40052 9260
rect 40186 9220 40195 9260
rect 40244 9220 40483 9260
rect 40523 9220 40771 9260
rect 40811 9220 41443 9260
rect 41483 9220 41731 9260
rect 41780 9220 42019 9260
rect 42059 9220 42307 9260
rect 42347 9220 42356 9260
rect 42835 9220 42844 9260
rect 42884 9220 43028 9260
rect 43075 9220 43084 9260
rect 43124 9220 43459 9260
rect 43499 9220 43508 9260
rect 43987 9220 43996 9260
rect 44036 9220 44276 9260
rect 44323 9220 44332 9260
rect 44372 9220 44860 9260
rect 44900 9220 44909 9260
rect 25516 9176 25556 9220
rect 40012 9176 40052 9220
rect 42316 9176 42356 9220
rect 21571 9136 21580 9176
rect 21620 9136 21868 9176
rect 21908 9136 21917 9176
rect 24268 9136 25556 9176
rect 27148 9136 34388 9176
rect 34435 9136 34444 9176
rect 34484 9136 36884 9176
rect 36931 9136 36940 9176
rect 36980 9136 39188 9176
rect 40012 9136 40492 9176
rect 40532 9136 40541 9176
rect 42316 9136 42892 9176
rect 42932 9136 42941 9176
rect 27148 9092 27188 9136
rect 34348 9092 34388 9136
rect 36844 9092 36884 9136
rect 1852 9052 4108 9092
rect 4148 9052 4157 9092
rect 4919 9052 4928 9092
rect 4968 9052 5010 9092
rect 5050 9052 5092 9092
rect 5132 9052 5174 9092
rect 5214 9052 5256 9092
rect 5296 9052 5305 9092
rect 7756 9052 18892 9092
rect 18932 9052 18941 9092
rect 19555 9052 19564 9092
rect 19604 9052 19988 9092
rect 20039 9052 20048 9092
rect 20088 9052 20130 9092
rect 20170 9052 20212 9092
rect 20252 9052 20294 9092
rect 20334 9052 20376 9092
rect 20416 9052 20425 9092
rect 20860 9052 27188 9092
rect 28387 9052 28396 9092
rect 28436 9052 33196 9092
rect 33236 9052 33245 9092
rect 34348 9052 34828 9092
rect 34868 9052 34877 9092
rect 35159 9052 35168 9092
rect 35208 9052 35250 9092
rect 35290 9052 35332 9092
rect 35372 9052 35414 9092
rect 35454 9052 35496 9092
rect 35536 9052 35545 9092
rect 36844 9052 37996 9092
rect 38036 9052 38045 9092
rect 0 9008 90 9028
rect 0 8968 1228 9008
rect 1268 8968 1277 9008
rect 1468 8968 12844 9008
rect 12884 8968 12893 9008
rect 12940 8968 15436 9008
rect 15476 8968 15485 9008
rect 15532 8968 20468 9008
rect 0 8948 90 8968
rect 1468 8924 1508 8968
rect 12940 8924 12980 8968
rect 15532 8924 15572 8968
rect 20428 8924 20468 8968
rect 20620 8968 22388 9008
rect 22435 8968 22444 9008
rect 22484 8968 24172 9008
rect 24212 8968 24221 9008
rect 26179 8968 26188 9008
rect 26228 8968 28108 9008
rect 28148 8968 28157 9008
rect 28579 8968 28588 9008
rect 28628 8968 32852 9008
rect 32995 8968 33004 9008
rect 33044 8968 38516 9008
rect 20620 8924 20660 8968
rect 1459 8884 1468 8924
rect 1508 8884 1517 8924
rect 2611 8884 2620 8924
rect 2660 8884 8044 8924
rect 8084 8884 8093 8924
rect 8227 8884 8236 8924
rect 8276 8884 9004 8924
rect 9044 8884 9053 8924
rect 10601 8884 10732 8924
rect 10772 8884 10781 8924
rect 10924 8884 12980 8924
rect 13555 8884 13564 8924
rect 13604 8884 13804 8924
rect 13844 8884 13853 8924
rect 13939 8884 13948 8924
rect 13988 8884 15476 8924
rect 15523 8884 15532 8924
rect 15572 8884 15581 8924
rect 16147 8884 16156 8924
rect 16196 8884 16300 8924
rect 16340 8884 16349 8924
rect 17731 8884 17740 8924
rect 17780 8884 18796 8924
rect 18836 8884 18845 8924
rect 19276 8884 20332 8924
rect 20372 8884 20381 8924
rect 20428 8884 20660 8924
rect 10924 8840 10964 8884
rect 1123 8800 1132 8840
rect 1172 8800 2420 8840
rect 4099 8800 4108 8840
rect 4148 8800 5780 8840
rect 5827 8800 5836 8840
rect 5876 8800 8468 8840
rect 8515 8800 8524 8840
rect 8564 8800 10252 8840
rect 10292 8800 10301 8840
rect 10444 8800 10964 8840
rect 11203 8800 11212 8840
rect 11252 8800 11261 8840
rect 13171 8800 13180 8840
rect 13220 8800 15148 8840
rect 15188 8800 15197 8840
rect 1036 8716 2036 8756
rect 2275 8716 2284 8756
rect 2324 8716 2333 8756
rect 0 8672 90 8692
rect 1036 8672 1076 8716
rect 1996 8672 2036 8716
rect 2284 8672 2324 8716
rect 2380 8672 2420 8800
rect 5740 8756 5780 8800
rect 8428 8756 8468 8800
rect 3523 8716 3532 8756
rect 3572 8716 4396 8756
rect 4436 8716 4445 8756
rect 5513 8716 5644 8756
rect 5684 8716 5693 8756
rect 5740 8716 6796 8756
rect 6836 8716 6845 8756
rect 8044 8747 8084 8756
rect 5644 8698 5684 8707
rect 8428 8716 8995 8756
rect 9035 8716 9044 8756
rect 9091 8716 9100 8756
rect 9140 8716 9196 8756
rect 9236 8716 9271 8756
rect 9353 8716 9484 8756
rect 9524 8716 9533 8756
rect 10025 8747 10156 8756
rect 10025 8716 10060 8747
rect 8044 8672 8084 8707
rect 10100 8716 10156 8747
rect 10196 8716 10205 8756
rect 10060 8698 10100 8707
rect 10444 8672 10484 8800
rect 11212 8756 11252 8800
rect 15436 8756 15476 8884
rect 15724 8800 16588 8840
rect 16628 8800 16637 8840
rect 17548 8800 18028 8840
rect 18068 8800 18077 8840
rect 18259 8800 18268 8840
rect 18308 8800 19180 8840
rect 19220 8800 19229 8840
rect 15724 8756 15764 8800
rect 10540 8747 11252 8756
rect 10580 8716 11252 8747
rect 11369 8747 11500 8756
rect 11369 8716 11404 8747
rect 10540 8698 10580 8707
rect 11444 8716 11500 8747
rect 11540 8716 11549 8756
rect 11971 8716 11980 8756
rect 12020 8736 12500 8756
rect 12643 8736 12652 8756
rect 12020 8716 12652 8736
rect 12692 8716 12701 8756
rect 12931 8716 12940 8756
rect 12980 8716 14092 8756
rect 14132 8716 14188 8756
rect 14228 8716 14292 8756
rect 15209 8716 15340 8756
rect 15380 8716 15389 8756
rect 15436 8716 15764 8756
rect 15811 8716 15820 8756
rect 15860 8716 16108 8756
rect 16148 8716 16300 8756
rect 16340 8716 16349 8756
rect 17548 8747 17588 8800
rect 11404 8698 11444 8707
rect 12460 8696 12692 8716
rect 15340 8698 15380 8707
rect 17548 8698 17588 8707
rect 18028 8716 18604 8756
rect 18644 8716 18653 8756
rect 18731 8716 18796 8756
rect 18836 8716 18862 8756
rect 18902 8716 18911 8756
rect 18979 8716 18988 8756
rect 19028 8716 19159 8756
rect 18028 8672 18068 8716
rect 19276 8672 19316 8884
rect 22348 8840 22388 8968
rect 32812 8924 32852 8968
rect 38476 8924 38516 8968
rect 39148 8924 39188 9136
rect 39235 9052 39244 9092
rect 39284 9052 40300 9092
rect 40340 9052 40349 9092
rect 42988 9008 43028 9220
rect 46278 9008 46368 9028
rect 40771 8968 40780 9008
rect 40820 8968 42836 9008
rect 42988 8968 46368 9008
rect 41356 8924 41396 8968
rect 42796 8924 42836 8968
rect 46278 8948 46368 8968
rect 22627 8884 22636 8924
rect 22676 8884 23212 8924
rect 23252 8884 23261 8924
rect 24835 8884 24844 8924
rect 24884 8884 26284 8924
rect 26324 8884 26333 8924
rect 26467 8884 26476 8924
rect 26516 8884 32668 8924
rect 32708 8884 32717 8924
rect 32812 8884 34004 8924
rect 34627 8884 34636 8924
rect 34676 8884 35060 8924
rect 35251 8884 35260 8924
rect 35300 8884 35692 8924
rect 35732 8884 35741 8924
rect 35849 8884 35980 8924
rect 36020 8884 36029 8924
rect 36163 8884 36172 8924
rect 36212 8884 38332 8924
rect 38372 8884 38381 8924
rect 38476 8884 39092 8924
rect 39148 8884 40924 8924
rect 40964 8884 40973 8924
rect 41347 8884 41356 8924
rect 41396 8884 41405 8924
rect 41609 8884 41731 8924
rect 41780 8884 41789 8924
rect 42787 8884 42796 8924
rect 42836 8884 42845 8924
rect 43699 8884 43708 8924
rect 43748 8884 44236 8924
rect 44276 8884 44285 8924
rect 44371 8884 44380 8924
rect 44420 8884 45196 8924
rect 45236 8884 45245 8924
rect 19372 8800 22060 8840
rect 22100 8800 22109 8840
rect 22348 8800 22964 8840
rect 19372 8756 19412 8800
rect 22924 8756 22964 8800
rect 26764 8800 27188 8840
rect 27235 8800 27244 8840
rect 27284 8800 27415 8840
rect 28265 8800 28348 8840
rect 28388 8800 28396 8840
rect 28436 8800 28445 8840
rect 28588 8800 30700 8840
rect 30740 8800 30749 8840
rect 30883 8800 30892 8840
rect 30932 8800 32276 8840
rect 32563 8800 32572 8840
rect 32612 8800 33044 8840
rect 33475 8800 33484 8840
rect 33524 8800 33676 8840
rect 33716 8800 33868 8840
rect 33908 8800 33917 8840
rect 26764 8756 26804 8800
rect 27148 8756 27188 8800
rect 28588 8756 28628 8800
rect 32236 8756 32276 8800
rect 19363 8716 19372 8756
rect 19412 8716 19421 8756
rect 19747 8716 19756 8756
rect 19796 8716 19943 8756
rect 19983 8716 20332 8756
rect 20372 8716 20381 8756
rect 20428 8747 20468 8756
rect 20890 8716 20899 8756
rect 20939 8716 20948 8756
rect 20995 8716 21004 8756
rect 21044 8716 21100 8756
rect 21140 8716 21175 8756
rect 21379 8716 21388 8756
rect 21428 8716 21437 8756
rect 21964 8747 22100 8756
rect 0 8632 1076 8672
rect 1123 8632 1132 8672
rect 1172 8632 1228 8672
rect 1268 8632 1303 8672
rect 1603 8632 1612 8672
rect 1652 8632 1661 8672
rect 1987 8632 1996 8672
rect 2036 8632 2045 8672
rect 2227 8632 2236 8672
rect 2276 8632 2324 8672
rect 2371 8632 2380 8672
rect 2420 8632 2429 8672
rect 8044 8632 8468 8672
rect 8515 8632 8524 8672
rect 8564 8632 8695 8672
rect 8755 8632 8764 8672
rect 8804 8632 9524 8672
rect 9571 8632 9580 8672
rect 9620 8632 9751 8672
rect 10156 8632 10484 8672
rect 11875 8632 11884 8672
rect 11924 8632 12268 8672
rect 12308 8632 12317 8672
rect 12931 8632 12940 8672
rect 12980 8632 13132 8672
rect 13172 8632 13181 8672
rect 13315 8632 13324 8672
rect 13364 8632 13373 8672
rect 13699 8632 13708 8672
rect 13748 8632 13804 8672
rect 13844 8632 13879 8672
rect 14755 8632 14764 8672
rect 14804 8632 15148 8672
rect 15188 8632 15197 8672
rect 15785 8632 15916 8672
rect 15956 8632 15965 8672
rect 18019 8632 18028 8672
rect 18068 8632 18077 8672
rect 18281 8632 18316 8672
rect 18356 8632 18412 8672
rect 18452 8632 18461 8672
rect 18643 8632 18652 8672
rect 18692 8632 19316 8672
rect 19459 8632 19468 8672
rect 19508 8632 20236 8672
rect 20276 8632 20285 8672
rect 0 8612 90 8632
rect 0 8336 90 8356
rect 1612 8336 1652 8632
rect 8428 8588 8468 8632
rect 9484 8588 9524 8632
rect 10156 8588 10196 8632
rect 13324 8588 13364 8632
rect 8428 8548 8620 8588
rect 8660 8548 8669 8588
rect 9484 8548 10196 8588
rect 13219 8548 13228 8588
rect 13268 8548 13364 8588
rect 1843 8464 1852 8504
rect 1892 8464 13900 8504
rect 13940 8464 13949 8504
rect 14371 8464 14380 8504
rect 14420 8464 15820 8504
rect 15860 8464 15869 8504
rect 17251 8464 17260 8504
rect 17300 8464 19276 8504
rect 19316 8464 19325 8504
rect 20428 8420 20468 8707
rect 20908 8672 20948 8716
rect 21388 8672 21428 8716
rect 22004 8716 22100 8747
rect 22313 8716 22348 8756
rect 22388 8747 22484 8756
rect 22388 8716 22444 8747
rect 21964 8698 22004 8707
rect 22060 8672 22100 8716
rect 22697 8716 22828 8756
rect 22868 8716 22877 8756
rect 22924 8716 23788 8756
rect 23828 8716 23837 8756
rect 24080 8714 24120 8723
rect 22444 8698 22484 8707
rect 24076 8674 24080 8714
rect 20515 8632 20524 8672
rect 20564 8632 20659 8672
rect 20699 8632 20708 8672
rect 20899 8632 20908 8672
rect 20948 8632 20995 8672
rect 21187 8632 21196 8672
rect 21236 8632 21428 8672
rect 21475 8632 21484 8672
rect 21524 8632 21676 8672
rect 21716 8632 21725 8672
rect 22051 8632 22060 8672
rect 22100 8632 22109 8672
rect 24076 8665 24120 8674
rect 24172 8716 24547 8756
rect 24587 8716 24596 8756
rect 24643 8716 24652 8756
rect 24692 8716 24823 8756
rect 25027 8716 25036 8756
rect 25076 8716 25502 8756
rect 25603 8716 25612 8756
rect 25652 8716 25783 8756
rect 25961 8716 26092 8756
rect 26132 8716 26141 8756
rect 26188 8716 26804 8756
rect 26851 8716 26860 8756
rect 26900 8716 26909 8756
rect 27130 8716 27139 8756
rect 27179 8716 27188 8756
rect 27244 8716 28628 8756
rect 29225 8747 29356 8756
rect 29225 8716 29260 8747
rect 24076 8588 24116 8665
rect 24067 8548 24076 8588
rect 24116 8548 24125 8588
rect 24172 8504 24212 8716
rect 25036 8672 25076 8716
rect 25462 8672 25502 8716
rect 25612 8698 25652 8707
rect 26092 8698 26132 8707
rect 24355 8632 24364 8672
rect 24404 8632 25076 8672
rect 25123 8632 25132 8672
rect 25172 8632 25303 8672
rect 25462 8632 25556 8672
rect 25516 8588 25556 8632
rect 26188 8588 26228 8716
rect 26860 8672 26900 8716
rect 27244 8672 27284 8716
rect 29300 8716 29356 8747
rect 29396 8716 29405 8756
rect 30403 8716 30412 8756
rect 30452 8716 30508 8756
rect 30548 8716 30583 8756
rect 30892 8747 31468 8756
rect 29260 8698 29300 8707
rect 30932 8716 31468 8747
rect 31508 8716 31517 8756
rect 32009 8716 32140 8756
rect 32180 8716 32189 8756
rect 32236 8716 32948 8756
rect 30892 8698 30932 8707
rect 32908 8672 32948 8716
rect 33004 8672 33044 8800
rect 33161 8716 33292 8756
rect 33332 8716 33341 8756
rect 33449 8716 33571 8756
rect 33620 8716 33629 8756
rect 33964 8672 34004 8884
rect 34051 8800 34060 8840
rect 34100 8800 34540 8840
rect 34580 8800 34828 8840
rect 34868 8800 34877 8840
rect 35020 8756 35060 8884
rect 35155 8800 35164 8840
rect 35204 8800 38996 8840
rect 34147 8716 34156 8756
rect 34196 8716 34444 8756
rect 34484 8716 34493 8756
rect 34714 8716 34723 8756
rect 34763 8716 34772 8756
rect 35020 8716 35980 8756
rect 36020 8716 36029 8756
rect 36172 8747 36212 8756
rect 34732 8672 34772 8716
rect 37411 8716 37420 8756
rect 37460 8716 37516 8756
rect 37556 8716 37591 8756
rect 37891 8716 37900 8756
rect 37940 8716 37949 8756
rect 38572 8716 38860 8756
rect 38900 8716 38909 8756
rect 36172 8672 36212 8707
rect 37900 8672 37940 8716
rect 38572 8672 38612 8716
rect 38956 8672 38996 8800
rect 39052 8756 39092 8884
rect 39379 8800 39388 8840
rect 39428 8800 41260 8840
rect 41300 8800 41309 8840
rect 43315 8800 43324 8840
rect 43364 8800 45044 8840
rect 39052 8716 39572 8756
rect 39619 8716 39628 8756
rect 39668 8716 39677 8756
rect 40003 8716 40012 8756
rect 40052 8716 41204 8756
rect 42883 8716 42892 8756
rect 42932 8716 44716 8756
rect 44756 8716 44765 8756
rect 39532 8672 39572 8716
rect 39628 8672 39668 8716
rect 41164 8672 41204 8716
rect 44716 8672 44756 8716
rect 45004 8672 45044 8800
rect 46278 8672 46368 8692
rect 26860 8632 27284 8672
rect 27427 8632 27436 8672
rect 27476 8632 27676 8672
rect 27716 8632 27725 8672
rect 27811 8632 27820 8672
rect 27860 8632 27916 8672
rect 27956 8632 27991 8672
rect 28099 8632 28108 8672
rect 28148 8632 28279 8672
rect 28553 8632 28684 8672
rect 28724 8632 28733 8672
rect 28937 8632 29059 8672
rect 29108 8632 29117 8672
rect 30979 8632 30988 8672
rect 31028 8632 32332 8672
rect 32372 8632 32381 8672
rect 32899 8632 32908 8672
rect 32948 8632 32957 8672
rect 33004 8632 33196 8672
rect 33236 8632 33245 8672
rect 33379 8632 33388 8672
rect 33428 8632 33908 8672
rect 33964 8632 34772 8672
rect 34915 8632 34924 8672
rect 34964 8632 35500 8672
rect 35540 8632 35549 8672
rect 35779 8632 35788 8672
rect 35828 8632 36212 8672
rect 36268 8632 37564 8672
rect 37604 8632 37613 8672
rect 37673 8632 37804 8672
rect 37844 8632 37853 8672
rect 37900 8632 37948 8672
rect 37988 8632 37997 8672
rect 38179 8632 38188 8672
rect 38228 8632 38516 8672
rect 38563 8632 38572 8672
rect 38612 8632 38621 8672
rect 38707 8632 38716 8672
rect 38756 8632 38764 8672
rect 38804 8632 38887 8672
rect 38947 8632 38956 8672
rect 38996 8632 39005 8672
rect 39139 8632 39148 8672
rect 39188 8632 39319 8672
rect 39523 8632 39532 8672
rect 39572 8632 39581 8672
rect 39628 8632 39868 8672
rect 39908 8632 39917 8672
rect 40099 8632 40108 8672
rect 40148 8632 40157 8672
rect 40387 8632 40396 8672
rect 40436 8632 40492 8672
rect 40532 8632 40567 8672
rect 40649 8632 40780 8672
rect 40820 8632 40829 8672
rect 41155 8632 41164 8672
rect 41204 8632 41213 8672
rect 42019 8632 42028 8672
rect 42068 8632 42316 8672
rect 42356 8632 42604 8672
rect 42644 8632 42653 8672
rect 42953 8632 43084 8672
rect 43124 8632 43133 8672
rect 43337 8632 43468 8672
rect 43508 8632 43517 8672
rect 43939 8632 43948 8672
rect 43988 8632 44140 8672
rect 44180 8632 44189 8672
rect 44716 8632 44908 8672
rect 44948 8632 44957 8672
rect 45004 8632 46368 8672
rect 33868 8588 33908 8632
rect 36268 8588 36308 8632
rect 24451 8548 24460 8588
rect 24500 8548 24596 8588
rect 25516 8548 26228 8588
rect 26284 8548 28444 8588
rect 28484 8548 28493 8588
rect 28963 8548 28972 8588
rect 29012 8548 29740 8588
rect 29780 8548 29789 8588
rect 29923 8548 29932 8588
rect 29972 8548 33004 8588
rect 33044 8548 33053 8588
rect 33868 8548 36308 8588
rect 24556 8504 24596 8548
rect 26284 8504 26324 8548
rect 38476 8504 38516 8632
rect 40108 8588 40148 8632
rect 38851 8548 38860 8588
rect 38900 8548 39772 8588
rect 39812 8548 40148 8588
rect 40492 8588 40532 8632
rect 42028 8588 42068 8632
rect 40492 8548 41740 8588
rect 41780 8548 42068 8588
rect 42604 8588 42644 8632
rect 43948 8588 43988 8632
rect 46278 8612 46368 8632
rect 42604 8548 43988 8588
rect 23779 8464 23788 8504
rect 23828 8464 24212 8504
rect 24259 8464 24268 8504
rect 24308 8464 24439 8504
rect 24556 8464 26324 8504
rect 27401 8464 27532 8504
rect 27572 8464 27581 8504
rect 28579 8464 28588 8504
rect 28628 8464 30220 8504
rect 30260 8464 30269 8504
rect 33955 8464 33964 8504
rect 34004 8464 35980 8504
rect 36020 8464 36029 8504
rect 36172 8464 38380 8504
rect 38420 8464 38429 8504
rect 38476 8464 41164 8504
rect 41204 8464 41213 8504
rect 45139 8464 45148 8504
rect 45188 8464 45772 8504
rect 45812 8464 45821 8504
rect 36172 8420 36212 8464
rect 8620 8380 10100 8420
rect 11011 8380 11020 8420
rect 11060 8380 19268 8420
rect 19939 8380 19948 8420
rect 19988 8380 20332 8420
rect 20372 8380 20381 8420
rect 20428 8380 20620 8420
rect 20660 8380 20669 8420
rect 22723 8380 22732 8420
rect 22772 8380 30260 8420
rect 32899 8380 32908 8420
rect 32948 8380 34868 8420
rect 34915 8380 34924 8420
rect 34964 8380 36212 8420
rect 36259 8380 36268 8420
rect 36308 8380 43220 8420
rect 0 8296 1652 8336
rect 3679 8296 3688 8336
rect 3728 8296 3770 8336
rect 3810 8296 3852 8336
rect 3892 8296 3934 8336
rect 3974 8296 4016 8336
rect 4056 8296 4065 8336
rect 0 8276 90 8296
rect 8620 8168 8660 8380
rect 10060 8252 10100 8380
rect 19228 8336 19268 8380
rect 14563 8296 14572 8336
rect 14612 8296 18604 8336
rect 18644 8296 18653 8336
rect 18799 8296 18808 8336
rect 18848 8296 18890 8336
rect 18930 8296 18972 8336
rect 19012 8296 19054 8336
rect 19094 8296 19136 8336
rect 19176 8296 19185 8336
rect 19228 8296 28780 8336
rect 28820 8296 28829 8336
rect 10060 8212 29932 8252
rect 29972 8212 29981 8252
rect 30220 8168 30260 8380
rect 34828 8336 34868 8380
rect 32515 8296 32524 8336
rect 32564 8296 33140 8336
rect 33919 8296 33928 8336
rect 33968 8296 34010 8336
rect 34050 8296 34092 8336
rect 34132 8296 34174 8336
rect 34214 8296 34256 8336
rect 34296 8296 34305 8336
rect 34828 8296 35060 8336
rect 35203 8296 35212 8336
rect 35252 8296 40204 8336
rect 40244 8296 40253 8336
rect 33100 8252 33140 8296
rect 30787 8212 30796 8252
rect 30836 8212 32716 8252
rect 32756 8212 32765 8252
rect 33100 8212 34732 8252
rect 34772 8212 34781 8252
rect 34828 8212 34924 8252
rect 34964 8212 34973 8252
rect 34828 8168 34868 8212
rect 4339 8128 4348 8168
rect 4388 8128 8660 8168
rect 10121 8128 10252 8168
rect 10292 8128 10301 8168
rect 11827 8128 11836 8168
rect 11876 8128 13612 8168
rect 13652 8128 13661 8168
rect 16435 8128 16444 8168
rect 16484 8128 17932 8168
rect 17972 8128 17981 8168
rect 19084 8128 22388 8168
rect 22435 8128 22444 8168
rect 22484 8128 25708 8168
rect 25748 8128 25757 8168
rect 25891 8128 25900 8168
rect 25940 8128 26092 8168
rect 26132 8128 26141 8168
rect 26284 8128 28148 8168
rect 28195 8128 28204 8168
rect 28244 8128 30164 8168
rect 30220 8128 30652 8168
rect 30692 8128 30701 8168
rect 32803 8128 32812 8168
rect 32852 8128 33292 8168
rect 33332 8128 33341 8168
rect 33772 8128 34868 8168
rect 652 8044 1132 8084
rect 1172 8044 1181 8084
rect 7171 8044 7180 8084
rect 7220 8044 9908 8084
rect 9955 8044 9964 8084
rect 10004 8044 10636 8084
rect 10676 8044 10685 8084
rect 10732 8044 11788 8084
rect 11828 8044 11837 8084
rect 12211 8044 12220 8084
rect 12260 8044 14092 8084
rect 14132 8044 14141 8084
rect 14188 8044 16628 8084
rect 0 8000 90 8020
rect 652 8000 692 8044
rect 9868 8000 9908 8044
rect 10732 8000 10772 8044
rect 14188 8000 14228 8044
rect 16588 8000 16628 8044
rect 16972 8044 17260 8084
rect 17300 8044 17309 8084
rect 16972 8000 17012 8044
rect 19084 8000 19124 8128
rect 20035 8044 20044 8084
rect 20084 8044 20524 8084
rect 20564 8044 20573 8084
rect 20716 8044 21388 8084
rect 21428 8044 21437 8084
rect 21484 8044 22156 8084
rect 22196 8044 22205 8084
rect 20716 8000 20756 8044
rect 21484 8000 21524 8044
rect 22348 8000 22388 8128
rect 22819 8044 22828 8084
rect 22868 8044 23636 8084
rect 23596 8000 23636 8044
rect 23692 8044 26188 8084
rect 26228 8044 26237 8084
rect 0 7960 692 8000
rect 1097 7960 1228 8000
rect 1268 7960 1277 8000
rect 1603 7960 1612 8000
rect 1652 7960 1661 8000
rect 3977 7960 4108 8000
rect 4148 7960 4157 8000
rect 9353 7960 9484 8000
rect 9524 7960 9533 8000
rect 9715 7960 9724 8000
rect 9764 7960 9812 8000
rect 9859 7960 9868 8000
rect 9908 7960 9917 8000
rect 10060 7960 10772 8000
rect 10819 7960 10828 8000
rect 10868 7960 11116 8000
rect 11156 7960 11212 8000
rect 11252 7960 11261 8000
rect 11465 7960 11500 8000
rect 11540 7960 11596 8000
rect 11636 7960 11645 8000
rect 11849 7960 11980 8000
rect 12020 7960 12029 8000
rect 12346 7960 12355 8000
rect 12395 7960 12404 8000
rect 13603 7960 13612 8000
rect 13652 7960 14228 8000
rect 16195 7960 16204 8000
rect 16244 7960 16300 8000
rect 16340 7960 16375 8000
rect 16579 7960 16588 8000
rect 16628 7960 16637 8000
rect 16963 7960 16972 8000
rect 17012 7960 17021 8000
rect 17203 7960 17212 8000
rect 17252 7960 17452 8000
rect 17492 7960 17501 8000
rect 18787 7960 18796 8000
rect 18836 7960 19124 8000
rect 19747 7960 19756 8000
rect 19796 7960 19805 8000
rect 20707 7960 20716 8000
rect 20756 7960 20765 8000
rect 21091 7960 21100 8000
rect 21140 7960 21149 8000
rect 21475 7960 21484 8000
rect 21524 7960 21533 8000
rect 21667 7960 21676 8000
rect 21716 7960 22252 8000
rect 22292 7960 22301 8000
rect 22348 7960 22972 8000
rect 23012 7960 23021 8000
rect 23081 7960 23212 8000
rect 23252 7960 23261 8000
rect 23347 7960 23356 8000
rect 23396 7960 23404 8000
rect 23444 7960 23527 8000
rect 23587 7960 23596 8000
rect 23636 7960 23645 8000
rect 0 7940 90 7960
rect 1612 7832 1652 7960
rect 4108 7916 4148 7960
rect 5740 7916 5780 7925
rect 8812 7916 8852 7925
rect 4108 7876 4492 7916
rect 4532 7876 4541 7916
rect 5609 7876 5740 7916
rect 5780 7876 5789 7916
rect 6787 7876 6796 7916
rect 6836 7876 7564 7916
rect 7604 7876 7613 7916
rect 9772 7916 9812 7960
rect 10060 7916 10100 7960
rect 12364 7916 12404 7960
rect 12556 7916 12596 7925
rect 15532 7916 15572 7925
rect 18604 7916 18644 7925
rect 19756 7916 19796 7960
rect 21100 7916 21140 7960
rect 23692 7916 23732 8044
rect 26284 8000 26324 8128
rect 28108 8084 28148 8128
rect 26371 8044 26380 8084
rect 26420 8044 27668 8084
rect 28099 8044 28108 8084
rect 28148 8044 28157 8084
rect 25708 7960 26324 8000
rect 27628 8000 27668 8044
rect 30124 8000 30164 8128
rect 33772 8084 33812 8128
rect 35020 8084 35060 8296
rect 35107 8212 35116 8252
rect 35156 8212 40396 8252
rect 40436 8212 40445 8252
rect 35971 8128 35980 8168
rect 36020 8128 37172 8168
rect 37411 8128 37420 8168
rect 37460 8128 39388 8168
rect 39428 8128 39437 8168
rect 30211 8044 30220 8084
rect 30260 8044 30269 8084
rect 30547 8044 30556 8084
rect 30596 8044 33812 8084
rect 33868 8044 34676 8084
rect 34723 8044 34732 8084
rect 34772 8044 34781 8084
rect 35020 8044 36508 8084
rect 36548 8044 36557 8084
rect 30220 8000 30260 8044
rect 33868 8000 33908 8044
rect 34636 8000 34676 8044
rect 34732 8000 34772 8044
rect 37132 8000 37172 8128
rect 37315 8044 37324 8084
rect 37364 8044 39148 8084
rect 39188 8044 39197 8084
rect 27628 7960 28492 8000
rect 28532 7960 28541 8000
rect 30115 7960 30124 8000
rect 30164 7960 30173 8000
rect 30220 7960 30316 8000
rect 30356 7960 30365 8000
rect 30883 7960 30892 8000
rect 30932 7960 30941 8000
rect 32707 7960 32716 8000
rect 32756 7960 33908 8000
rect 34627 7960 34636 8000
rect 34676 7960 34685 8000
rect 34732 7960 36124 8000
rect 36164 7960 36173 8000
rect 36233 7960 36364 8000
rect 36404 7960 36413 8000
rect 36617 7960 36748 8000
rect 36788 7960 36797 8000
rect 37123 7960 37132 8000
rect 37172 7960 37181 8000
rect 25708 7916 25748 7960
rect 27532 7916 27572 7925
rect 29068 7916 29108 7925
rect 30892 7916 30932 7960
rect 32620 7916 32660 7925
rect 34252 7916 34292 7925
rect 37564 7916 37604 8044
rect 43180 8000 43220 8380
rect 46278 8336 46368 8356
rect 44995 8296 45004 8336
rect 45044 8296 46368 8336
rect 46278 8276 46368 8296
rect 44371 8128 44380 8168
rect 44420 8128 44716 8168
rect 44756 8128 44765 8168
rect 46278 8000 46368 8020
rect 39619 7960 39628 8000
rect 39668 7960 39677 8000
rect 40675 7960 40684 8000
rect 40724 7960 41452 8000
rect 41492 7960 41501 8000
rect 41731 7960 41740 8000
rect 41780 7960 42124 8000
rect 42164 7960 42173 8000
rect 43180 7960 44140 8000
rect 44180 7960 44189 8000
rect 44323 7960 44332 8000
rect 44372 7960 44524 8000
rect 44564 7960 44573 8000
rect 44899 7960 44908 8000
rect 44948 7960 44957 8000
rect 45763 7960 45772 8000
rect 45812 7960 46368 8000
rect 38764 7916 38804 7925
rect 39628 7916 39668 7960
rect 44908 7916 44948 7960
rect 46278 7940 46368 7960
rect 9772 7876 10100 7916
rect 10505 7876 10636 7916
rect 10676 7876 10685 7916
rect 10915 7876 10924 7916
rect 10964 7876 12404 7916
rect 12521 7876 12556 7916
rect 12596 7876 12652 7916
rect 12692 7876 12701 7916
rect 13027 7876 13036 7916
rect 13076 7876 13804 7916
rect 13844 7876 13853 7916
rect 14249 7876 14284 7916
rect 14324 7876 14380 7916
rect 14420 7876 14429 7916
rect 15331 7876 15340 7916
rect 15380 7876 15532 7916
rect 15572 7876 15820 7916
rect 15860 7876 15869 7916
rect 17059 7876 17068 7916
rect 17108 7876 17356 7916
rect 17396 7876 17405 7916
rect 18019 7876 18028 7916
rect 18068 7876 18604 7916
rect 19363 7876 19372 7916
rect 19412 7876 19421 7916
rect 19642 7876 19651 7916
rect 19691 7876 19796 7916
rect 19939 7876 19948 7916
rect 19988 7876 19997 7916
rect 20131 7876 20140 7916
rect 20180 7876 20428 7916
rect 20468 7876 20477 7916
rect 21100 7876 21772 7916
rect 21812 7876 21821 7916
rect 22147 7876 22156 7916
rect 22196 7876 22205 7916
rect 22426 7876 22435 7916
rect 22475 7876 23732 7916
rect 23779 7876 23788 7916
rect 23828 7876 24460 7916
rect 24500 7876 24509 7916
rect 25795 7876 25804 7916
rect 25844 7876 26284 7916
rect 26324 7876 26333 7916
rect 5740 7867 5780 7876
rect 844 7792 1652 7832
rect 8812 7832 8852 7876
rect 12556 7867 12596 7876
rect 10636 7858 10676 7867
rect 13804 7832 13844 7876
rect 15532 7867 15572 7876
rect 18604 7867 18644 7876
rect 19372 7832 19412 7876
rect 19948 7832 19988 7876
rect 22156 7832 22196 7876
rect 25708 7832 25748 7876
rect 27532 7832 27572 7876
rect 27724 7876 28003 7916
rect 28043 7876 28052 7916
rect 28099 7876 28108 7916
rect 28148 7876 28157 7916
rect 28457 7876 28588 7916
rect 28628 7876 28637 7916
rect 29347 7876 29356 7916
rect 29396 7876 29556 7916
rect 29596 7876 29605 7916
rect 29731 7876 29740 7916
rect 29780 7876 30932 7916
rect 31241 7876 31372 7916
rect 31412 7876 32140 7916
rect 32180 7876 32189 7916
rect 32803 7876 32812 7916
rect 32852 7876 33004 7916
rect 33044 7876 33053 7916
rect 34147 7876 34156 7916
rect 34196 7876 34252 7916
rect 34292 7876 34327 7916
rect 34915 7876 34924 7916
rect 34964 7876 35308 7916
rect 35348 7876 35357 7916
rect 35572 7876 35587 7916
rect 35627 7876 35636 7916
rect 36019 7876 36028 7916
rect 36068 7876 37460 7916
rect 37507 7876 37516 7916
rect 37556 7876 37604 7916
rect 38659 7876 38668 7916
rect 38708 7876 38764 7916
rect 38804 7876 39820 7916
rect 39860 7876 39869 7916
rect 41251 7876 41260 7916
rect 41300 7876 44948 7916
rect 27724 7832 27764 7876
rect 8812 7792 10004 7832
rect 10339 7792 10348 7832
rect 10388 7792 10540 7832
rect 10580 7792 10589 7832
rect 11116 7792 12172 7832
rect 12212 7792 12221 7832
rect 13804 7792 14572 7832
rect 14612 7792 14621 7832
rect 16819 7792 16828 7832
rect 16868 7792 18220 7832
rect 18260 7792 18269 7832
rect 18787 7792 18796 7832
rect 18836 7792 19412 7832
rect 19459 7792 19468 7832
rect 19508 7792 19740 7832
rect 19780 7792 19789 7832
rect 19948 7792 21244 7832
rect 21284 7792 21293 7832
rect 21667 7792 21676 7832
rect 21716 7792 22196 7832
rect 22243 7792 22252 7832
rect 22292 7792 22540 7832
rect 22580 7792 22828 7832
rect 22868 7792 22877 7832
rect 24163 7792 24172 7832
rect 24212 7792 25748 7832
rect 25987 7792 25996 7832
rect 26036 7792 27340 7832
rect 27380 7792 27572 7832
rect 27715 7792 27724 7832
rect 27764 7792 27773 7832
rect 0 7664 90 7684
rect 844 7664 884 7792
rect 1459 7708 1468 7748
rect 1508 7708 1708 7748
rect 1748 7708 1757 7748
rect 1843 7708 1852 7748
rect 1892 7708 2860 7748
rect 2900 7708 2909 7748
rect 5801 7708 5932 7748
rect 5972 7708 5981 7748
rect 8995 7708 9004 7748
rect 9044 7708 9053 7748
rect 0 7624 884 7664
rect 0 7604 90 7624
rect 4919 7540 4928 7580
rect 4968 7540 5010 7580
rect 5050 7540 5092 7580
rect 5132 7540 5174 7580
rect 5214 7540 5256 7580
rect 5296 7540 5305 7580
rect 0 7328 90 7348
rect 0 7288 1228 7328
rect 1268 7288 1277 7328
rect 0 7268 90 7288
rect 9004 7244 9044 7708
rect 9964 7664 10004 7792
rect 11116 7748 11156 7792
rect 28108 7748 28148 7876
rect 29068 7832 29108 7876
rect 32620 7832 32660 7876
rect 34252 7867 34292 7876
rect 35572 7832 35612 7876
rect 37420 7832 37460 7876
rect 38764 7867 38804 7876
rect 29068 7792 31124 7832
rect 31651 7792 31660 7832
rect 31700 7792 32660 7832
rect 33283 7792 33292 7832
rect 33332 7792 33716 7832
rect 31084 7748 31124 7792
rect 33676 7748 33716 7792
rect 34348 7792 34580 7832
rect 34867 7792 34876 7832
rect 34916 7792 35612 7832
rect 35657 7792 35692 7832
rect 35732 7792 35788 7832
rect 35828 7792 35837 7832
rect 35971 7792 35980 7832
rect 36020 7792 36892 7832
rect 36932 7792 36941 7832
rect 37420 7792 37708 7832
rect 37748 7792 37757 7832
rect 40972 7792 41836 7832
rect 41876 7792 42412 7832
rect 42452 7792 42700 7832
rect 42740 7792 42988 7832
rect 43028 7792 43276 7832
rect 43316 7792 43325 7832
rect 34348 7748 34388 7792
rect 10099 7708 10108 7748
rect 10148 7708 11156 7748
rect 11443 7708 11452 7748
rect 11492 7708 15052 7748
rect 15092 7708 15101 7748
rect 15331 7708 15340 7748
rect 15380 7708 15724 7748
rect 15764 7708 15773 7748
rect 19843 7708 19852 7748
rect 19892 7708 20476 7748
rect 20516 7708 20525 7748
rect 20851 7708 20860 7748
rect 20900 7708 21100 7748
rect 21140 7708 21149 7748
rect 21907 7708 21916 7748
rect 21956 7708 22444 7748
rect 22484 7708 22493 7748
rect 24643 7708 24652 7748
rect 24692 7708 28148 7748
rect 28387 7708 28396 7748
rect 28436 7708 29740 7748
rect 29780 7708 29789 7748
rect 29875 7708 29884 7748
rect 29924 7708 29932 7748
rect 29972 7708 30055 7748
rect 31084 7708 33580 7748
rect 33620 7708 33629 7748
rect 33676 7708 34388 7748
rect 34435 7708 34444 7748
rect 34484 7708 34493 7748
rect 9964 7624 11500 7664
rect 11540 7624 11549 7664
rect 12163 7624 12172 7664
rect 12212 7624 19756 7664
rect 19796 7624 19805 7664
rect 19900 7624 34252 7664
rect 34292 7624 34301 7664
rect 9091 7540 9100 7580
rect 9140 7540 14764 7580
rect 14804 7540 14813 7580
rect 15523 7540 15532 7580
rect 15572 7540 19700 7580
rect 19660 7496 19700 7540
rect 19900 7496 19940 7624
rect 20039 7540 20048 7580
rect 20088 7540 20130 7580
rect 20170 7540 20212 7580
rect 20252 7540 20294 7580
rect 20334 7540 20376 7580
rect 20416 7540 20425 7580
rect 27619 7540 27628 7580
rect 27668 7540 28396 7580
rect 28436 7540 28445 7580
rect 29059 7540 29068 7580
rect 29108 7540 34156 7580
rect 34196 7540 34205 7580
rect 10540 7456 11156 7496
rect 15043 7456 15052 7496
rect 15092 7456 19604 7496
rect 19660 7456 19940 7496
rect 20044 7456 29492 7496
rect 9667 7372 9676 7412
rect 9716 7372 10108 7412
rect 10148 7372 10157 7412
rect 10540 7328 10580 7456
rect 11116 7328 11156 7456
rect 19564 7412 19604 7456
rect 20044 7412 20084 7456
rect 29452 7412 29492 7456
rect 9641 7288 9772 7328
rect 9812 7288 10580 7328
rect 10636 7288 10732 7328
rect 10772 7288 10781 7328
rect 11011 7288 11020 7328
rect 11060 7288 11156 7328
rect 11836 7372 18796 7412
rect 18836 7372 18845 7412
rect 19564 7372 20084 7412
rect 20140 7372 21716 7412
rect 22435 7372 22444 7412
rect 22484 7372 28052 7412
rect 29225 7372 29356 7412
rect 29396 7372 29405 7412
rect 29452 7372 33100 7412
rect 33140 7372 33149 7412
rect 33331 7372 33340 7412
rect 33380 7372 33580 7412
rect 33620 7372 33629 7412
rect 33715 7372 33724 7412
rect 33764 7372 33964 7412
rect 34004 7372 34013 7412
rect 10636 7244 10676 7288
rect 9004 7204 9388 7244
rect 9428 7204 9437 7244
rect 9658 7204 9667 7244
rect 9707 7204 10444 7244
rect 10484 7204 10493 7244
rect 10627 7204 10636 7244
rect 10676 7204 10685 7244
rect 10889 7204 10915 7244
rect 10955 7204 11020 7244
rect 11060 7204 11069 7244
rect 67 7120 76 7160
rect 116 7120 1228 7160
rect 1268 7120 1277 7160
rect 1603 7120 1612 7160
rect 1652 7120 1661 7160
rect 1843 7120 1852 7160
rect 1892 7120 3532 7160
rect 3572 7120 3581 7160
rect 6185 7120 6316 7160
rect 6356 7120 6365 7160
rect 6547 7120 6556 7160
rect 6596 7120 7180 7160
rect 7220 7120 7229 7160
rect 8009 7120 8140 7160
rect 8180 7120 8189 7160
rect 8515 7120 8524 7160
rect 8564 7120 8573 7160
rect 8777 7120 8908 7160
rect 8948 7120 8957 7160
rect 9139 7120 9148 7160
rect 9188 7120 10732 7160
rect 10772 7120 10781 7160
rect 11561 7120 11692 7160
rect 11732 7120 11741 7160
rect 1612 7076 1652 7120
rect 172 7036 1652 7076
rect 8524 7076 8564 7120
rect 11836 7076 11876 7372
rect 20140 7328 20180 7372
rect 21676 7328 21716 7372
rect 28012 7328 28052 7372
rect 13891 7288 13900 7328
rect 13940 7288 18892 7328
rect 18932 7288 18941 7328
rect 19459 7288 19468 7328
rect 19508 7288 20180 7328
rect 21667 7288 21676 7328
rect 21716 7288 21725 7328
rect 21955 7288 21964 7328
rect 22004 7288 22580 7328
rect 23011 7288 23020 7328
rect 23060 7288 23069 7328
rect 23212 7288 23596 7328
rect 23636 7288 23645 7328
rect 25603 7288 25612 7328
rect 25652 7288 27724 7328
rect 27764 7288 27773 7328
rect 28012 7288 31084 7328
rect 31124 7288 31133 7328
rect 31843 7288 31852 7328
rect 31892 7288 32276 7328
rect 32947 7288 32956 7328
rect 32996 7288 34348 7328
rect 34388 7288 34397 7328
rect 12460 7204 12940 7244
rect 12980 7204 12989 7244
rect 13516 7204 14476 7244
rect 14516 7204 14525 7244
rect 15052 7204 15380 7244
rect 12460 7160 12500 7204
rect 13516 7160 13556 7204
rect 15052 7160 15092 7204
rect 11945 7120 11980 7160
rect 12020 7120 12076 7160
rect 12116 7120 12125 7160
rect 12451 7120 12460 7160
rect 12500 7120 12509 7160
rect 12713 7120 12844 7160
rect 12884 7120 12893 7160
rect 13027 7120 13036 7160
rect 13076 7120 13228 7160
rect 13268 7120 13277 7160
rect 13459 7120 13468 7160
rect 13508 7120 13556 7160
rect 13603 7120 13612 7160
rect 13652 7120 13661 7160
rect 13865 7120 13900 7160
rect 13940 7120 13996 7160
rect 14036 7120 14045 7160
rect 14249 7120 14380 7160
rect 14420 7120 14429 7160
rect 14563 7120 14572 7160
rect 14612 7120 14764 7160
rect 14804 7120 14813 7160
rect 14995 7120 15004 7160
rect 15044 7120 15092 7160
rect 15139 7120 15148 7160
rect 15188 7120 15284 7160
rect 13612 7076 13652 7120
rect 8524 7036 11876 7076
rect 12307 7036 12316 7076
rect 12356 7036 13516 7076
rect 13556 7036 13565 7076
rect 13612 7036 14092 7076
rect 14132 7036 14141 7076
rect 14227 7036 14236 7076
rect 14276 7036 14860 7076
rect 14900 7036 14909 7076
rect 0 6992 90 7012
rect 0 6952 76 6992
rect 116 6952 125 6992
rect 0 6932 90 6952
rect 0 6656 90 6676
rect 172 6656 212 7036
rect 1459 6952 1468 6992
rect 1508 6952 1748 6992
rect 3763 6952 3772 6992
rect 3812 6952 4300 6992
rect 4340 6952 4349 6992
rect 8371 6952 8380 6992
rect 8420 6952 8660 6992
rect 8755 6952 8764 6992
rect 8804 6952 10540 6992
rect 10580 6952 10589 6992
rect 10723 6952 10732 6992
rect 10772 6952 11116 6992
rect 11156 6952 11165 6992
rect 11299 6952 11308 6992
rect 11348 6952 11788 6992
rect 11828 6952 11837 6992
rect 11923 6952 11932 6992
rect 11972 6952 12404 6992
rect 12691 6952 12700 6992
rect 12740 6952 12940 6992
rect 12980 6952 12989 6992
rect 13075 6952 13084 6992
rect 13124 6952 13708 6992
rect 13748 6952 13757 6992
rect 13843 6952 13852 6992
rect 13892 6952 14380 6992
rect 14420 6952 14429 6992
rect 14611 6952 14620 6992
rect 14660 6952 14764 6992
rect 14804 6952 14813 6992
rect 1708 6908 1748 6952
rect 8620 6908 8660 6952
rect 12364 6908 12404 6952
rect 1708 6868 8564 6908
rect 8620 6868 9964 6908
rect 10004 6868 10013 6908
rect 12364 6868 12748 6908
rect 12788 6868 12797 6908
rect 8524 6824 8564 6868
rect 3679 6784 3688 6824
rect 3728 6784 3770 6824
rect 3810 6784 3852 6824
rect 3892 6784 3934 6824
rect 3974 6784 4016 6824
rect 4056 6784 4065 6824
rect 8524 6784 11212 6824
rect 11252 6784 11261 6824
rect 12892 6784 13324 6824
rect 13364 6784 13373 6824
rect 0 6616 212 6656
rect 4972 6700 12748 6740
rect 12788 6700 12797 6740
rect 0 6596 90 6616
rect 67 6448 76 6488
rect 116 6448 1228 6488
rect 1268 6448 1277 6488
rect 1603 6448 1612 6488
rect 1652 6448 1661 6488
rect 1612 6404 1652 6448
rect 4972 6404 5012 6700
rect 12892 6656 12932 6784
rect 15244 6740 15284 7120
rect 15340 7076 15380 7204
rect 16204 7204 16492 7244
rect 16532 7204 16541 7244
rect 16684 7204 17068 7244
rect 17108 7204 17117 7244
rect 17443 7204 17452 7244
rect 17492 7235 18356 7244
rect 17492 7204 18316 7235
rect 15523 7120 15532 7160
rect 15572 7120 15703 7160
rect 15907 7120 15916 7160
rect 15956 7120 16108 7160
rect 16148 7120 16157 7160
rect 16204 7076 16244 7204
rect 16684 7160 16724 7204
rect 18403 7204 18412 7244
rect 18452 7204 19316 7244
rect 18316 7186 18356 7195
rect 19276 7160 19316 7204
rect 19372 7204 20084 7244
rect 20515 7204 20524 7244
rect 20564 7204 20573 7244
rect 21161 7204 21292 7244
rect 21332 7204 21341 7244
rect 21449 7204 21571 7244
rect 21620 7204 22156 7244
rect 22196 7204 22205 7244
rect 16291 7120 16300 7160
rect 16340 7120 16471 7160
rect 16675 7120 16684 7160
rect 16724 7120 16855 7160
rect 18883 7120 18892 7160
rect 18932 7120 19063 7160
rect 19267 7120 19276 7160
rect 19316 7120 19325 7160
rect 19372 7076 19412 7204
rect 20044 7160 20084 7204
rect 20524 7160 20564 7204
rect 22540 7160 22580 7288
rect 23020 7244 23060 7288
rect 23212 7244 23252 7288
rect 32236 7244 32276 7288
rect 34444 7244 34484 7708
rect 34540 7664 34580 7792
rect 35572 7748 35612 7792
rect 40972 7748 41012 7792
rect 35572 7708 36076 7748
rect 36116 7708 36125 7748
rect 38825 7708 38956 7748
rect 38996 7708 39005 7748
rect 39235 7708 39244 7748
rect 39284 7708 40780 7748
rect 40820 7708 40963 7748
rect 41003 7708 41012 7748
rect 41068 7708 41212 7748
rect 41252 7708 41261 7748
rect 42202 7708 42211 7748
rect 42251 7708 43651 7748
rect 43691 7708 43843 7748
rect 43883 7708 43892 7748
rect 44755 7708 44764 7748
rect 44804 7708 44813 7748
rect 45139 7708 45148 7748
rect 45188 7708 45772 7748
rect 45812 7708 45821 7748
rect 41068 7664 41108 7708
rect 34540 7624 41108 7664
rect 35159 7540 35168 7580
rect 35208 7540 35250 7580
rect 35290 7540 35332 7580
rect 35372 7540 35414 7580
rect 35454 7540 35496 7580
rect 35536 7540 35545 7580
rect 36739 7540 36748 7580
rect 36788 7540 40972 7580
rect 41012 7540 41021 7580
rect 42220 7412 42260 7708
rect 44764 7664 44804 7708
rect 46278 7664 46368 7684
rect 44764 7624 46368 7664
rect 46278 7604 46368 7624
rect 36355 7372 36364 7412
rect 36404 7372 41452 7412
rect 41492 7372 41501 7412
rect 41705 7372 41827 7412
rect 41876 7372 41885 7412
rect 42220 7372 42499 7412
rect 42539 7372 42787 7412
rect 42827 7372 42836 7412
rect 46278 7328 46368 7348
rect 34540 7288 34828 7328
rect 34868 7288 34877 7328
rect 35500 7288 36076 7328
rect 36116 7288 36125 7328
rect 37891 7288 37900 7328
rect 37940 7288 39916 7328
rect 39956 7288 39965 7328
rect 45763 7288 45772 7328
rect 45812 7288 46368 7328
rect 34540 7244 34580 7288
rect 23011 7204 23020 7244
rect 23060 7204 23107 7244
rect 23212 7204 23275 7244
rect 23315 7204 23324 7244
rect 23386 7204 23395 7244
rect 23435 7204 23444 7244
rect 27139 7204 27148 7244
rect 27188 7223 27860 7244
rect 27907 7223 27916 7244
rect 27188 7204 27916 7223
rect 27956 7204 27965 7244
rect 29059 7204 29068 7244
rect 29108 7235 29239 7244
rect 29108 7204 29164 7235
rect 23404 7160 23444 7204
rect 27820 7183 27956 7204
rect 29204 7204 29239 7235
rect 29452 7204 29548 7244
rect 29588 7204 30700 7244
rect 30740 7204 30749 7244
rect 31651 7204 31660 7244
rect 31700 7235 32140 7244
rect 31700 7204 31948 7235
rect 29164 7186 29204 7195
rect 29452 7160 29492 7204
rect 31988 7204 32140 7235
rect 32180 7204 32189 7244
rect 32236 7204 33140 7244
rect 33667 7204 33676 7244
rect 33716 7204 34196 7244
rect 34426 7204 34435 7244
rect 34475 7204 34484 7244
rect 34531 7204 34540 7244
rect 34580 7204 34589 7244
rect 34636 7204 34924 7244
rect 34964 7204 34973 7244
rect 35500 7235 35540 7288
rect 46278 7268 46368 7288
rect 31948 7186 31988 7195
rect 33100 7160 33140 7204
rect 34156 7160 34196 7204
rect 19529 7120 19660 7160
rect 19700 7120 19709 7160
rect 19817 7120 19900 7160
rect 19940 7120 19948 7160
rect 19988 7120 19997 7160
rect 20044 7120 20180 7160
rect 20227 7120 20236 7160
rect 20276 7120 20564 7160
rect 20611 7120 20620 7160
rect 20660 7120 20669 7160
rect 20755 7120 20764 7160
rect 20804 7120 20812 7160
rect 20852 7120 20935 7160
rect 20995 7120 21004 7160
rect 21044 7120 21964 7160
rect 22004 7120 22013 7160
rect 22339 7120 22348 7160
rect 22388 7120 22397 7160
rect 22531 7120 22540 7160
rect 22580 7120 22589 7160
rect 22819 7120 22828 7160
rect 22868 7120 23444 7160
rect 23779 7120 23788 7160
rect 23828 7120 23980 7160
rect 24020 7120 24029 7160
rect 25001 7120 25036 7160
rect 25076 7120 25132 7160
rect 25172 7120 25181 7160
rect 25315 7120 25324 7160
rect 25364 7120 25708 7160
rect 25748 7120 25757 7160
rect 26083 7120 26092 7160
rect 26132 7120 26141 7160
rect 26921 7120 26956 7160
rect 26996 7120 27052 7160
rect 27092 7120 27101 7160
rect 27523 7120 27532 7160
rect 27572 7120 27724 7160
rect 27764 7120 27773 7160
rect 29452 7120 29500 7160
rect 29540 7120 29549 7160
rect 29635 7120 29644 7160
rect 29684 7120 30124 7160
rect 30164 7120 30173 7160
rect 30281 7120 30316 7160
rect 30356 7120 30412 7160
rect 30452 7120 30461 7160
rect 32044 7120 32524 7160
rect 32564 7120 32573 7160
rect 32707 7120 32716 7160
rect 32756 7120 32887 7160
rect 33091 7120 33100 7160
rect 33140 7120 33149 7160
rect 33475 7120 33484 7160
rect 33524 7120 33533 7160
rect 33929 7120 34060 7160
rect 34100 7120 34109 7160
rect 34156 7120 34540 7160
rect 34580 7120 34589 7160
rect 20140 7076 20180 7120
rect 20620 7076 20660 7120
rect 22348 7076 22388 7120
rect 26092 7076 26132 7120
rect 32044 7076 32084 7120
rect 33484 7076 33524 7120
rect 34636 7076 34676 7204
rect 35849 7204 35980 7244
rect 36020 7204 36029 7244
rect 36460 7204 37076 7244
rect 39305 7204 39436 7244
rect 39476 7204 39485 7244
rect 40553 7204 40684 7244
rect 40724 7204 40733 7244
rect 35500 7186 35540 7195
rect 35980 7186 36020 7195
rect 34723 7120 34732 7160
rect 34772 7120 35020 7160
rect 35060 7120 35069 7160
rect 36460 7076 36500 7204
rect 37036 7160 37076 7204
rect 40684 7186 40724 7195
rect 36547 7120 36556 7160
rect 36596 7120 36605 7160
rect 36809 7120 36940 7160
rect 36980 7120 36989 7160
rect 37036 7120 37324 7160
rect 37364 7120 37373 7160
rect 37577 7120 37708 7160
rect 37748 7120 37757 7160
rect 42211 7120 42220 7160
rect 42260 7120 42269 7160
rect 43171 7120 43180 7160
rect 43220 7120 43276 7160
rect 43316 7120 43468 7160
rect 43508 7120 43756 7160
rect 43796 7120 43852 7160
rect 43892 7120 44044 7160
rect 44084 7120 44332 7160
rect 44372 7120 44524 7160
rect 44564 7120 44573 7160
rect 44777 7120 44908 7160
rect 44948 7120 44957 7160
rect 15340 7036 15572 7076
rect 15763 7036 15772 7076
rect 15812 7036 16244 7076
rect 16531 7036 16540 7076
rect 16580 7036 17164 7076
rect 17204 7036 17213 7076
rect 18988 7036 19412 7076
rect 19507 7036 19516 7076
rect 19556 7036 19852 7076
rect 19892 7036 19901 7076
rect 20140 7036 20564 7076
rect 20620 7036 20716 7076
rect 20756 7036 20765 7076
rect 21955 7036 21964 7076
rect 22004 7036 22388 7076
rect 23203 7036 23212 7076
rect 23252 7036 25132 7076
rect 25172 7036 25181 7076
rect 25411 7036 25420 7076
rect 25460 7036 26132 7076
rect 27331 7036 27340 7076
rect 27380 7036 27484 7076
rect 27524 7036 27533 7076
rect 29657 7036 29740 7076
rect 29780 7036 29788 7076
rect 29828 7036 29837 7076
rect 30019 7036 30028 7076
rect 30068 7036 32084 7076
rect 32131 7036 32140 7076
rect 32180 7036 32620 7076
rect 32660 7036 32669 7076
rect 32803 7036 32812 7076
rect 32852 7036 33524 7076
rect 33859 7036 33868 7076
rect 33908 7036 34676 7076
rect 35587 7036 35596 7076
rect 35636 7036 36500 7076
rect 36556 7076 36596 7120
rect 42220 7076 42260 7120
rect 36556 7036 38092 7076
rect 38132 7036 38141 7076
rect 41836 7036 42260 7076
rect 44755 7036 44764 7076
rect 44804 7036 46156 7076
rect 46196 7036 46205 7076
rect 15532 6992 15572 7036
rect 18988 6992 19028 7036
rect 20524 6992 20564 7036
rect 15379 6952 15388 6992
rect 15428 6952 15476 6992
rect 15532 6952 16012 6992
rect 16052 6952 16061 6992
rect 16147 6952 16156 6992
rect 16196 6952 16780 6992
rect 16820 6952 16829 6992
rect 16915 6952 16924 6992
rect 16964 6952 17068 6992
rect 17108 6952 17117 6992
rect 18499 6952 18508 6992
rect 18548 6952 19028 6992
rect 19123 6952 19132 6992
rect 19172 6952 19180 6992
rect 19220 6952 19303 6992
rect 19987 6952 19996 6992
rect 20036 6952 20140 6992
rect 20180 6952 20189 6992
rect 20371 6952 20380 6992
rect 20420 6952 20468 6992
rect 20524 6952 20908 6992
rect 20948 6952 20957 6992
rect 21571 6952 21580 6992
rect 21620 6952 22108 6992
rect 22148 6952 22157 6992
rect 22771 6952 22780 6992
rect 22820 6952 23404 6992
rect 23444 6952 23453 6992
rect 23561 6952 23692 6992
rect 23732 6952 23741 6992
rect 24211 6952 24220 6992
rect 24260 6952 24364 6992
rect 24404 6952 24413 6992
rect 25363 6952 25372 6992
rect 25412 6952 25844 6992
rect 25891 6952 25900 6992
rect 25940 6952 25948 6992
rect 25988 6952 26071 6992
rect 26323 6952 26332 6992
rect 26372 6952 27052 6992
rect 27092 6952 27101 6992
rect 27283 6952 27292 6992
rect 27332 6952 29644 6992
rect 29684 6952 29693 6992
rect 29875 6952 29884 6992
rect 29924 6952 29933 6992
rect 30547 6952 30556 6992
rect 30596 6952 31852 6992
rect 31892 6952 31901 6992
rect 32227 6952 32236 6992
rect 32276 6952 32284 6992
rect 32324 6952 32407 6992
rect 32995 6952 33004 6992
rect 33044 6952 33820 6992
rect 33860 6952 33869 6992
rect 34540 6952 36211 6992
rect 36251 6952 36260 6992
rect 36307 6952 36316 6992
rect 36356 6952 36404 6992
rect 15436 6824 15476 6952
rect 20428 6908 20468 6952
rect 25804 6908 25844 6952
rect 29884 6908 29924 6952
rect 34540 6908 34580 6952
rect 36364 6908 36404 6952
rect 20428 6868 21004 6908
rect 21044 6868 21053 6908
rect 25804 6868 26572 6908
rect 26612 6868 26621 6908
rect 26755 6868 26764 6908
rect 26804 6868 29924 6908
rect 30019 6868 30028 6908
rect 30068 6868 32716 6908
rect 32756 6868 32765 6908
rect 33571 6868 33580 6908
rect 33620 6868 34580 6908
rect 34627 6868 34636 6908
rect 34676 6868 36404 6908
rect 36460 6952 36700 6992
rect 36740 6952 36749 6992
rect 36835 6952 36844 6992
rect 36884 6952 37084 6992
rect 37124 6952 37133 6992
rect 37315 6952 37324 6992
rect 37364 6952 37468 6992
rect 37508 6952 37517 6992
rect 40867 6952 40876 6992
rect 40916 6952 41260 6992
rect 41300 6952 41309 6992
rect 36460 6824 36500 6952
rect 15436 6784 16396 6824
rect 16436 6784 16445 6824
rect 18799 6784 18808 6824
rect 18848 6784 18890 6824
rect 18930 6784 18972 6824
rect 19012 6784 19054 6824
rect 19094 6784 19136 6824
rect 19176 6784 19185 6824
rect 26659 6784 26668 6824
rect 26708 6784 29740 6824
rect 29780 6784 29789 6824
rect 33919 6784 33928 6824
rect 33968 6784 34010 6824
rect 34050 6784 34092 6824
rect 34132 6784 34174 6824
rect 34214 6784 34256 6824
rect 34296 6784 34305 6824
rect 34435 6784 34444 6824
rect 34484 6784 36500 6824
rect 13276 6700 13516 6740
rect 13556 6700 13565 6740
rect 14371 6700 14380 6740
rect 14420 6700 14668 6740
rect 14708 6700 14717 6740
rect 15244 6700 15916 6740
rect 15956 6700 15965 6740
rect 16483 6700 16492 6740
rect 16532 6700 22636 6740
rect 22676 6700 22685 6740
rect 29827 6700 29836 6740
rect 29876 6700 32716 6740
rect 32756 6700 32765 6740
rect 13276 6656 13316 6700
rect 41836 6656 41876 7036
rect 46278 6992 46368 7012
rect 41923 6952 41932 6992
rect 41972 6952 41980 6992
rect 42020 6952 42103 6992
rect 45139 6952 45148 6992
rect 45188 6952 46368 6992
rect 46278 6932 46368 6952
rect 46278 6656 46368 6676
rect 10099 6616 10108 6656
rect 10148 6616 11116 6656
rect 11156 6616 11165 6656
rect 12425 6616 12508 6656
rect 12548 6616 12556 6656
rect 12596 6616 12605 6656
rect 12883 6616 12892 6656
rect 12932 6616 12941 6656
rect 13267 6616 13276 6656
rect 13316 6616 13325 6656
rect 15235 6616 15244 6656
rect 15284 6616 15292 6656
rect 15332 6616 15415 6656
rect 17347 6616 17356 6656
rect 17396 6616 17404 6656
rect 17444 6616 17527 6656
rect 17731 6616 17740 6656
rect 17780 6616 17788 6656
rect 17828 6616 17911 6656
rect 18451 6616 18460 6656
rect 18500 6616 18700 6656
rect 18740 6616 18749 6656
rect 20035 6616 20044 6656
rect 20084 6616 20620 6656
rect 20660 6616 20669 6656
rect 22147 6616 22156 6656
rect 22196 6616 22924 6656
rect 22964 6616 22973 6656
rect 23203 6616 23212 6656
rect 23252 6616 26668 6656
rect 26708 6616 26717 6656
rect 27043 6616 27052 6656
rect 27092 6616 32812 6656
rect 32852 6616 32861 6656
rect 33955 6616 33964 6656
rect 34004 6616 34828 6656
rect 34868 6616 34877 6656
rect 35971 6616 35980 6656
rect 36020 6616 36748 6656
rect 36788 6616 36797 6656
rect 37027 6616 37036 6656
rect 37076 6616 40244 6656
rect 41827 6616 41836 6656
rect 41876 6616 41885 6656
rect 42019 6616 42028 6656
rect 42068 6616 43996 6656
rect 44036 6616 44045 6656
rect 46243 6616 46252 6656
rect 46292 6616 46368 6656
rect 40204 6572 40244 6616
rect 46278 6596 46368 6616
rect 5731 6532 5740 6572
rect 5780 6532 7892 6572
rect 10147 6532 10156 6572
rect 10196 6532 12172 6572
rect 12212 6532 12221 6572
rect 13036 6532 14324 6572
rect 5740 6448 5932 6488
rect 5972 6448 5981 6488
rect 6089 6448 6220 6488
rect 6260 6448 6269 6488
rect 7642 6448 7651 6488
rect 7691 6448 7700 6488
rect 5740 6404 5780 6448
rect 6796 6404 6836 6413
rect 7660 6404 7700 6448
rect 172 6364 1652 6404
rect 3523 6364 3532 6404
rect 3572 6364 3724 6404
rect 3764 6364 3773 6404
rect 5722 6364 5731 6404
rect 5771 6364 5780 6404
rect 5827 6364 5836 6404
rect 5876 6364 6164 6404
rect 6281 6364 6316 6404
rect 6356 6364 6412 6404
rect 6452 6364 6461 6404
rect 6665 6364 6796 6404
rect 6836 6364 6845 6404
rect 7306 6364 7315 6404
rect 7355 6364 7700 6404
rect 7852 6404 7892 6532
rect 9475 6448 9484 6488
rect 9524 6448 9676 6488
rect 9716 6448 9725 6488
rect 9859 6448 9868 6488
rect 9908 6448 10252 6488
rect 10292 6448 10301 6488
rect 10444 6404 10484 6532
rect 13036 6488 13076 6532
rect 10819 6448 10828 6488
rect 10868 6448 11020 6488
rect 11060 6448 11069 6488
rect 12137 6448 12268 6488
rect 12308 6448 12317 6488
rect 12521 6448 12556 6488
rect 12596 6448 12652 6488
rect 12692 6448 12701 6488
rect 13027 6448 13036 6488
rect 13076 6448 13085 6488
rect 11404 6404 11444 6413
rect 8803 6364 8812 6404
rect 8852 6364 9100 6404
rect 9140 6364 9388 6404
rect 9428 6364 9437 6404
rect 10060 6364 10156 6404
rect 10196 6364 10205 6404
rect 0 6320 90 6340
rect 0 6280 76 6320
rect 116 6280 125 6320
rect 0 6260 90 6280
rect 0 5984 90 6004
rect 172 5984 212 6364
rect 4972 6355 5012 6364
rect 1459 6196 1468 6236
rect 1508 6196 1556 6236
rect 1843 6196 1852 6236
rect 1892 6196 2900 6236
rect 5155 6196 5164 6236
rect 5204 6196 5644 6236
rect 5684 6196 5693 6236
rect 0 5944 212 5984
rect 0 5924 90 5944
rect 1516 5900 1556 6196
rect 2860 5984 2900 6196
rect 6124 6152 6164 6364
rect 6796 6355 6836 6364
rect 7852 6355 7892 6364
rect 10060 6320 10100 6364
rect 10252 6363 10318 6403
rect 10358 6363 10367 6403
rect 10435 6364 10444 6404
rect 10484 6364 10493 6404
rect 10627 6364 10636 6404
rect 10676 6364 10924 6404
rect 10964 6364 10973 6404
rect 11369 6364 11404 6404
rect 11444 6364 11500 6404
rect 11540 6364 11549 6404
rect 11914 6364 11923 6404
rect 11963 6364 12652 6404
rect 12692 6364 12701 6404
rect 10252 6320 10292 6363
rect 11404 6320 11444 6364
rect 13036 6320 13076 6448
rect 9187 6280 9196 6320
rect 9236 6280 10100 6320
rect 10243 6280 10252 6320
rect 10292 6280 10301 6320
rect 10435 6280 10444 6320
rect 10484 6280 11444 6320
rect 11980 6280 13076 6320
rect 13612 6404 13652 6413
rect 14284 6404 14324 6532
rect 18220 6532 23020 6572
rect 23060 6532 23069 6572
rect 23404 6532 24268 6572
rect 24308 6532 27964 6572
rect 28004 6532 28013 6572
rect 28099 6532 28108 6572
rect 28148 6532 28724 6572
rect 28867 6532 28876 6572
rect 28916 6532 32620 6572
rect 32660 6532 32669 6572
rect 34217 6532 34348 6572
rect 34388 6532 34397 6572
rect 35299 6532 35308 6572
rect 35348 6532 35596 6572
rect 35636 6532 35645 6572
rect 35779 6532 35788 6572
rect 35828 6532 36308 6572
rect 36547 6532 36556 6572
rect 36596 6532 37420 6572
rect 37460 6532 37469 6572
rect 40204 6532 42412 6572
rect 42452 6532 42461 6572
rect 42787 6532 42796 6572
rect 42836 6532 43220 6572
rect 18220 6488 18260 6532
rect 23404 6488 23444 6532
rect 14371 6448 14380 6488
rect 14420 6448 15532 6488
rect 15572 6448 15581 6488
rect 17513 6448 17644 6488
rect 17684 6448 17693 6488
rect 17897 6448 18028 6488
rect 18068 6448 18077 6488
rect 18211 6448 18220 6488
rect 18260 6448 18269 6488
rect 19939 6448 19948 6488
rect 19988 6448 20236 6488
rect 20276 6448 20285 6488
rect 20467 6448 20476 6488
rect 20516 6448 21772 6488
rect 21812 6448 21821 6488
rect 22147 6448 22156 6488
rect 22196 6448 22924 6488
rect 22964 6448 22973 6488
rect 23020 6448 23444 6488
rect 24425 6448 24556 6488
rect 24596 6448 24605 6488
rect 25315 6448 25324 6488
rect 25364 6448 26516 6488
rect 27017 6448 27148 6488
rect 27188 6448 27197 6488
rect 27907 6448 27916 6488
rect 27956 6448 28204 6488
rect 28244 6448 28253 6488
rect 16012 6404 16052 6413
rect 19852 6404 19892 6413
rect 20476 6404 20516 6448
rect 23020 6404 23060 6448
rect 23500 6404 23540 6413
rect 25228 6404 25268 6413
rect 26476 6404 26516 6448
rect 28684 6404 28724 6532
rect 28771 6448 28780 6488
rect 28820 6448 31468 6488
rect 31508 6448 31517 6488
rect 31564 6404 31604 6413
rect 33196 6404 33236 6413
rect 36268 6404 36308 6532
rect 43180 6488 43220 6532
rect 44044 6532 44948 6572
rect 39523 6448 39532 6488
rect 39572 6448 39581 6488
rect 40300 6448 41492 6488
rect 43171 6448 43180 6488
rect 43220 6448 43229 6488
rect 36940 6404 36980 6413
rect 14284 6364 14668 6404
rect 14708 6364 14860 6404
rect 14900 6364 14909 6404
rect 15043 6364 15052 6404
rect 15092 6364 16012 6404
rect 16052 6364 16061 6404
rect 17129 6364 17260 6404
rect 17300 6364 17309 6404
rect 18115 6364 18124 6404
rect 18164 6364 18604 6404
rect 18644 6364 18653 6404
rect 19171 6364 19180 6404
rect 19220 6364 19852 6404
rect 19892 6364 20516 6404
rect 20585 6364 20716 6404
rect 20756 6364 20765 6404
rect 21929 6364 21972 6404
rect 22012 6364 22060 6404
rect 22100 6364 22109 6404
rect 22243 6364 22252 6404
rect 22292 6364 22435 6404
rect 22475 6364 22484 6404
rect 22531 6364 22540 6404
rect 22580 6364 22711 6404
rect 23011 6364 23020 6404
rect 23060 6364 23069 6404
rect 23465 6364 23500 6404
rect 23540 6364 23596 6404
rect 23636 6364 23645 6404
rect 24010 6364 24019 6404
rect 24059 6364 25076 6404
rect 13612 6320 13652 6364
rect 16012 6355 16052 6364
rect 19852 6355 19892 6364
rect 23500 6355 23540 6364
rect 25036 6320 25076 6364
rect 25268 6364 25900 6404
rect 25940 6364 25949 6404
rect 26467 6364 26476 6404
rect 26516 6364 26525 6404
rect 28963 6364 28972 6404
rect 29012 6364 29548 6404
rect 29588 6364 29932 6404
rect 29972 6364 30316 6404
rect 30356 6364 30420 6404
rect 31363 6364 31372 6404
rect 31412 6364 31564 6404
rect 31939 6364 31948 6404
rect 31988 6364 32044 6404
rect 32084 6364 32119 6404
rect 32227 6364 32236 6404
rect 32276 6364 33196 6404
rect 25228 6355 25268 6364
rect 28684 6320 28724 6364
rect 31564 6355 31604 6364
rect 33196 6355 33236 6364
rect 33292 6364 33676 6404
rect 33716 6364 33725 6404
rect 33772 6364 33955 6404
rect 33995 6364 34004 6404
rect 34156 6364 34636 6404
rect 34676 6364 34685 6404
rect 34819 6364 34828 6404
rect 34868 6364 34915 6404
rect 34955 6364 34999 6404
rect 35849 6364 35884 6404
rect 35924 6364 35980 6404
rect 36020 6364 36029 6404
rect 36076 6364 36139 6404
rect 36179 6364 36188 6404
rect 36250 6364 36259 6404
rect 36299 6364 36308 6404
rect 36739 6364 36748 6404
rect 36788 6364 36940 6404
rect 38057 6364 38188 6404
rect 38228 6364 38237 6404
rect 38891 6364 38956 6404
rect 38996 6364 39022 6404
rect 39062 6364 39071 6404
rect 39139 6364 39148 6404
rect 39188 6364 39197 6404
rect 13612 6280 13653 6320
rect 13891 6280 13900 6320
rect 13940 6280 15956 6320
rect 16099 6280 16108 6320
rect 16148 6280 19468 6320
rect 19508 6280 19517 6320
rect 20428 6280 23060 6320
rect 11980 6236 12020 6280
rect 7337 6196 7468 6236
rect 7508 6196 7517 6236
rect 9715 6196 9724 6236
rect 9764 6196 10004 6236
rect 11107 6196 11116 6236
rect 11156 6196 12020 6236
rect 12067 6196 12076 6236
rect 12116 6196 12268 6236
rect 12308 6196 12317 6236
rect 13324 6196 13420 6236
rect 13460 6196 13469 6236
rect 9964 6152 10004 6196
rect 13324 6152 13364 6196
rect 13613 6152 13653 6280
rect 15916 6236 15956 6280
rect 20428 6236 20468 6280
rect 23020 6236 23060 6280
rect 23596 6280 24316 6320
rect 24356 6280 24365 6320
rect 25027 6280 25036 6320
rect 25076 6280 25085 6320
rect 27331 6280 27340 6320
rect 27380 6280 28492 6320
rect 28532 6280 28541 6320
rect 28675 6280 28684 6320
rect 28724 6280 28800 6320
rect 31660 6280 33004 6320
rect 33044 6280 33053 6320
rect 23596 6236 23636 6280
rect 13987 6196 13996 6236
rect 14036 6196 15820 6236
rect 15860 6196 15869 6236
rect 15916 6196 20468 6236
rect 20515 6196 20524 6236
rect 20564 6196 22252 6236
rect 22292 6196 22301 6236
rect 23020 6196 23636 6236
rect 24163 6196 24172 6236
rect 24212 6196 25900 6236
rect 25940 6196 25949 6236
rect 27379 6196 27388 6236
rect 27428 6196 28300 6236
rect 28340 6196 28349 6236
rect 31660 6152 31700 6280
rect 33292 6236 33332 6364
rect 33772 6320 33812 6364
rect 33667 6280 33676 6320
rect 33716 6280 33812 6320
rect 33929 6280 34060 6320
rect 34100 6280 34109 6320
rect 34156 6236 34196 6364
rect 34627 6280 34636 6320
rect 34676 6280 35020 6320
rect 35060 6280 35788 6320
rect 35828 6280 35837 6320
rect 31747 6196 31756 6236
rect 31796 6196 33332 6236
rect 33379 6196 33388 6236
rect 33428 6196 34196 6236
rect 36076 6236 36116 6364
rect 36940 6355 36980 6364
rect 39148 6320 39188 6364
rect 37891 6280 37900 6320
rect 37940 6280 39188 6320
rect 39532 6236 39572 6448
rect 40108 6404 40148 6413
rect 40300 6404 40340 6448
rect 41452 6404 41492 6448
rect 39619 6364 39628 6404
rect 39668 6364 39799 6404
rect 39977 6364 40108 6404
rect 40148 6364 40340 6404
rect 40579 6364 40588 6404
rect 40636 6364 40759 6404
rect 41129 6364 41164 6404
rect 41204 6364 41260 6404
rect 41300 6364 41309 6404
rect 41434 6364 41443 6404
rect 41483 6364 41492 6404
rect 41993 6364 42124 6404
rect 42164 6364 42173 6404
rect 42281 6364 42403 6404
rect 42452 6364 42461 6404
rect 40108 6355 40148 6364
rect 40867 6280 40876 6320
rect 40916 6280 41548 6320
rect 41588 6280 42508 6320
rect 42548 6280 42557 6320
rect 36076 6196 39572 6236
rect 40387 6196 40396 6236
rect 40436 6196 40780 6236
rect 40820 6196 40829 6236
rect 41731 6196 41740 6236
rect 41780 6196 42940 6236
rect 42980 6196 42989 6236
rect 43546 6196 43555 6236
rect 43595 6196 43843 6236
rect 43892 6196 43901 6236
rect 36076 6152 36116 6196
rect 6124 6112 9196 6152
rect 9236 6112 9245 6152
rect 9964 6112 13268 6152
rect 13315 6112 13324 6152
rect 13364 6112 13373 6152
rect 13613 6112 15820 6152
rect 15860 6112 15869 6152
rect 16003 6112 16012 6152
rect 16052 6112 19180 6152
rect 19220 6112 19229 6152
rect 19651 6112 19660 6152
rect 19700 6112 23212 6152
rect 23252 6112 23261 6152
rect 23587 6112 23596 6152
rect 23636 6112 31700 6152
rect 31747 6112 31756 6152
rect 31796 6112 36116 6152
rect 39619 6112 39628 6152
rect 39668 6112 42412 6152
rect 42452 6112 42461 6152
rect 13228 6068 13268 6112
rect 44044 6068 44084 6532
rect 44908 6488 44948 6532
rect 44227 6448 44236 6488
rect 44276 6448 44285 6488
rect 44393 6448 44428 6488
rect 44468 6448 44524 6488
rect 44564 6448 44573 6488
rect 44899 6448 44908 6488
rect 44948 6448 44957 6488
rect 4919 6028 4928 6068
rect 4968 6028 5010 6068
rect 5050 6028 5092 6068
rect 5132 6028 5174 6068
rect 5214 6028 5256 6068
rect 5296 6028 5305 6068
rect 13228 6028 18412 6068
rect 18452 6028 18461 6068
rect 20039 6028 20048 6068
rect 20088 6028 20130 6068
rect 20170 6028 20212 6068
rect 20252 6028 20294 6068
rect 20334 6028 20376 6068
rect 20416 6028 20425 6068
rect 20716 6028 26764 6068
rect 26804 6028 26813 6068
rect 28972 6028 35060 6068
rect 35159 6028 35168 6068
rect 35208 6028 35250 6068
rect 35290 6028 35332 6068
rect 35372 6028 35414 6068
rect 35454 6028 35496 6068
rect 35536 6028 35545 6068
rect 36355 6028 36364 6068
rect 36404 6028 44084 6068
rect 20716 5984 20756 6028
rect 2860 5944 12748 5984
rect 12788 5944 12797 5984
rect 13891 5944 13900 5984
rect 13940 5944 20756 5984
rect 20803 5944 20812 5984
rect 20852 5944 28876 5984
rect 28916 5944 28925 5984
rect 28972 5900 29012 6028
rect 35020 5984 35060 6028
rect 44236 5984 44276 6448
rect 46278 6320 46368 6340
rect 45139 6280 45148 6320
rect 45188 6280 46368 6320
rect 46278 6260 46368 6280
rect 44755 6196 44764 6236
rect 44804 6196 44813 6236
rect 44764 6152 44804 6196
rect 44764 6112 46252 6152
rect 46292 6112 46301 6152
rect 46278 5984 46368 6004
rect 31555 5944 31564 5984
rect 31604 5944 32516 5984
rect 35020 5944 41932 5984
rect 41972 5944 41981 5984
rect 44236 5944 44372 5984
rect 46243 5944 46252 5984
rect 46292 5944 46368 5984
rect 32476 5900 32516 5944
rect 1516 5860 12940 5900
rect 12980 5860 12989 5900
rect 13987 5860 13996 5900
rect 14036 5860 22924 5900
rect 22964 5860 22973 5900
rect 23107 5860 23116 5900
rect 23156 5860 29012 5900
rect 29635 5860 29644 5900
rect 29684 5860 31988 5900
rect 32467 5860 32476 5900
rect 32516 5860 32525 5900
rect 41923 5860 41932 5900
rect 41972 5860 42124 5900
rect 42164 5860 42173 5900
rect 43162 5860 43171 5900
rect 43211 5860 43459 5900
rect 43499 5860 44236 5900
rect 44276 5860 44285 5900
rect 31948 5816 31988 5860
rect 44332 5816 44372 5944
rect 46278 5924 46368 5944
rect 5923 5776 5932 5816
rect 5972 5776 6028 5816
rect 6068 5776 8756 5816
rect 8803 5776 8812 5816
rect 8852 5776 9676 5816
rect 9716 5776 9725 5816
rect 10339 5776 10348 5816
rect 10388 5776 11116 5816
rect 11156 5776 11165 5816
rect 11827 5776 11836 5816
rect 11876 5776 13036 5816
rect 13076 5776 13085 5816
rect 15820 5776 16492 5816
rect 16532 5776 17204 5816
rect 19267 5776 19276 5816
rect 19316 5776 21332 5816
rect 21571 5776 21580 5816
rect 21620 5776 22732 5816
rect 22772 5776 22781 5816
rect 23212 5776 23692 5816
rect 23732 5776 23741 5816
rect 31660 5776 31892 5816
rect 31948 5776 39628 5816
rect 39668 5776 39677 5816
rect 40771 5776 40780 5816
rect 40820 5776 44372 5816
rect 3401 5692 3532 5732
rect 3572 5692 3581 5732
rect 4771 5692 4780 5732
rect 4820 5723 4951 5732
rect 4824 5692 4951 5723
rect 5513 5692 5644 5732
rect 5684 5692 5693 5732
rect 5914 5692 5923 5732
rect 5963 5692 6220 5732
rect 6260 5692 6269 5732
rect 4784 5674 4824 5683
rect 0 5648 90 5668
rect 8716 5648 8756 5776
rect 15820 5732 15860 5776
rect 17164 5732 17204 5776
rect 21292 5732 21332 5776
rect 8932 5692 8941 5732
rect 8981 5692 9004 5732
rect 9044 5692 9121 5732
rect 9187 5692 9196 5732
rect 9236 5692 10676 5732
rect 10723 5692 10732 5732
rect 10772 5692 10781 5732
rect 10889 5692 11011 5732
rect 11060 5692 11069 5732
rect 13516 5723 13556 5732
rect 0 5608 1228 5648
rect 1268 5608 1277 5648
rect 1603 5608 1612 5648
rect 1652 5608 1661 5648
rect 1865 5608 1996 5648
rect 2036 5608 2045 5648
rect 6412 5608 6508 5648
rect 6548 5608 6557 5648
rect 8716 5608 9772 5648
rect 9812 5608 9821 5648
rect 10051 5608 10060 5648
rect 10100 5608 10252 5648
rect 10292 5608 10301 5648
rect 0 5588 90 5608
rect 1612 5564 1652 5608
rect 172 5524 1652 5564
rect 2227 5524 2236 5564
rect 2276 5524 4684 5564
rect 4724 5524 4733 5564
rect 4876 5524 5836 5564
rect 5876 5524 5885 5564
rect 6185 5524 6316 5564
rect 6356 5524 6365 5564
rect 0 5312 90 5332
rect 172 5312 212 5524
rect 4876 5480 4916 5524
rect 6412 5480 6452 5608
rect 1459 5440 1468 5480
rect 1508 5440 1517 5480
rect 1843 5440 1852 5480
rect 1892 5440 4916 5480
rect 4963 5440 4972 5480
rect 5012 5440 5452 5480
rect 5492 5440 5501 5480
rect 6124 5440 6452 5480
rect 6739 5440 6748 5480
rect 6788 5440 8332 5480
rect 8372 5440 8381 5480
rect 8515 5440 8524 5480
rect 8564 5440 9004 5480
rect 9044 5440 9053 5480
rect 10409 5440 10492 5480
rect 10532 5440 10540 5480
rect 10580 5440 10589 5480
rect 1468 5396 1508 5440
rect 1468 5356 6028 5396
rect 6068 5356 6077 5396
rect 0 5272 212 5312
rect 3679 5272 3688 5312
rect 3728 5272 3770 5312
rect 3810 5272 3852 5312
rect 3892 5272 3934 5312
rect 3974 5272 4016 5312
rect 4056 5272 4065 5312
rect 0 5252 90 5272
rect 6124 5144 6164 5440
rect 10636 5312 10676 5692
rect 10732 5396 10772 5692
rect 14659 5692 14668 5732
rect 14708 5692 14724 5732
rect 14764 5692 14839 5732
rect 14956 5692 15860 5732
rect 15907 5692 15916 5732
rect 15956 5692 16087 5732
rect 17155 5692 17164 5732
rect 17204 5692 18028 5732
rect 18068 5692 18077 5732
rect 19276 5723 19316 5732
rect 11587 5608 11596 5648
rect 11636 5608 11645 5648
rect 11779 5608 11788 5648
rect 11828 5608 11980 5648
rect 12020 5608 12029 5648
rect 12355 5608 12364 5648
rect 12404 5608 12412 5648
rect 12452 5608 12535 5648
rect 12643 5608 12652 5648
rect 12692 5608 12701 5648
rect 12835 5608 12844 5648
rect 12884 5608 12980 5648
rect 13123 5608 13132 5648
rect 13172 5608 13315 5648
rect 13355 5608 13364 5648
rect 11596 5564 11636 5608
rect 11395 5524 11404 5564
rect 11444 5524 11636 5564
rect 12652 5564 12692 5608
rect 12940 5564 12980 5608
rect 13516 5564 13556 5683
rect 14956 5648 14996 5692
rect 15916 5674 15956 5683
rect 19913 5692 20044 5732
rect 20084 5692 20716 5732
rect 20756 5692 21004 5732
rect 21044 5692 21053 5732
rect 21292 5723 21388 5732
rect 19276 5648 19316 5683
rect 21332 5692 21388 5723
rect 21428 5692 21492 5732
rect 22252 5692 22540 5732
rect 22580 5692 22589 5732
rect 21292 5674 21332 5683
rect 22252 5648 22292 5692
rect 23212 5648 23252 5776
rect 31660 5732 31700 5776
rect 31852 5732 31892 5776
rect 23299 5692 23308 5732
rect 23348 5692 23404 5732
rect 23444 5692 23479 5732
rect 23578 5692 23587 5732
rect 23627 5692 24268 5732
rect 24308 5692 24317 5732
rect 25900 5723 25940 5732
rect 25987 5692 25996 5732
rect 26036 5692 27148 5732
rect 27188 5692 27197 5732
rect 27497 5692 27532 5732
rect 27572 5692 27628 5732
rect 27668 5692 27677 5732
rect 28876 5723 28916 5732
rect 14179 5608 14188 5648
rect 14228 5608 14956 5648
rect 14996 5608 15005 5648
rect 15052 5608 15532 5648
rect 15572 5608 15764 5648
rect 19276 5608 19948 5648
rect 19988 5608 19997 5648
rect 21948 5608 22060 5648
rect 22100 5608 22108 5648
rect 22148 5608 22292 5648
rect 22339 5608 22348 5648
rect 22388 5608 22444 5648
rect 22484 5608 22519 5648
rect 23011 5608 23020 5648
rect 23060 5608 23252 5648
rect 23683 5608 23692 5648
rect 23732 5608 24364 5648
rect 24404 5608 24413 5648
rect 25123 5608 25132 5648
rect 25172 5608 25324 5648
rect 25364 5608 25373 5648
rect 25577 5608 25699 5648
rect 25748 5608 25757 5648
rect 15052 5564 15092 5608
rect 15724 5564 15764 5608
rect 12652 5524 12748 5564
rect 12788 5524 12797 5564
rect 12931 5524 12940 5564
rect 12980 5524 12989 5564
rect 13516 5524 14668 5564
rect 14708 5524 15092 5564
rect 15187 5524 15196 5564
rect 15236 5524 15628 5564
rect 15668 5524 15677 5564
rect 15724 5524 18932 5564
rect 19459 5524 19468 5564
rect 19508 5524 20524 5564
rect 20564 5524 20573 5564
rect 21283 5524 21292 5564
rect 21332 5524 21484 5564
rect 21524 5524 21533 5564
rect 18892 5480 18932 5524
rect 22348 5480 22388 5608
rect 23020 5524 24124 5564
rect 24164 5524 24173 5564
rect 25481 5524 25564 5564
rect 25604 5524 25612 5564
rect 25652 5524 25661 5564
rect 23020 5480 23060 5524
rect 12211 5440 12220 5480
rect 12260 5440 12652 5480
rect 12692 5440 12701 5480
rect 13075 5440 13084 5480
rect 13124 5440 15148 5480
rect 15188 5440 15197 5480
rect 15283 5440 15292 5480
rect 15332 5440 15436 5480
rect 15476 5440 15485 5480
rect 15715 5440 15724 5480
rect 15764 5440 15773 5480
rect 15907 5440 15916 5480
rect 15956 5440 17836 5480
rect 17876 5440 18836 5480
rect 18892 5440 22388 5480
rect 22444 5440 23060 5480
rect 23971 5440 23980 5480
rect 24020 5440 24556 5480
rect 24596 5440 24605 5480
rect 15724 5396 15764 5440
rect 10732 5356 15764 5396
rect 18796 5396 18836 5440
rect 18796 5356 22252 5396
rect 22292 5356 22301 5396
rect 22444 5312 22484 5440
rect 25900 5396 25940 5683
rect 29251 5692 29260 5732
rect 29300 5692 30508 5732
rect 30548 5692 30557 5732
rect 31084 5692 31700 5732
rect 31756 5723 31796 5732
rect 28876 5648 28916 5683
rect 29836 5648 29876 5692
rect 26179 5608 26188 5648
rect 26228 5608 28876 5648
rect 28916 5608 28925 5648
rect 29321 5608 29452 5648
rect 29492 5608 29501 5648
rect 29827 5608 29836 5648
rect 29876 5608 29885 5648
rect 31084 5564 31124 5692
rect 31852 5692 33379 5732
rect 33419 5692 33428 5732
rect 33475 5692 33484 5732
rect 33524 5692 33676 5732
rect 33716 5692 33964 5732
rect 34004 5692 34013 5732
rect 34444 5723 34636 5732
rect 31756 5648 31796 5683
rect 34484 5692 34636 5723
rect 34676 5692 34685 5732
rect 34819 5692 34828 5732
rect 34868 5723 34999 5732
rect 34868 5692 34924 5723
rect 34444 5674 34484 5683
rect 29059 5524 29068 5564
rect 29108 5524 31124 5564
rect 31372 5608 31796 5648
rect 32323 5608 32332 5648
rect 32372 5608 32381 5648
rect 32707 5608 32716 5648
rect 32756 5608 32908 5648
rect 32948 5608 32957 5648
rect 33091 5608 33100 5648
rect 33140 5608 33196 5648
rect 33236 5608 33271 5648
rect 33741 5608 33868 5648
rect 33912 5608 33921 5648
rect 33964 5608 34003 5648
rect 34043 5608 34060 5648
rect 34100 5608 34212 5648
rect 31372 5480 31412 5608
rect 32332 5564 32372 5608
rect 33964 5564 34004 5608
rect 31747 5524 31756 5564
rect 31796 5524 31948 5564
rect 31988 5524 31997 5564
rect 32044 5524 32092 5564
rect 32132 5524 32141 5564
rect 32332 5524 33004 5564
rect 33044 5524 33053 5564
rect 33475 5524 33484 5564
rect 33524 5524 34004 5564
rect 28963 5440 28972 5480
rect 29012 5440 29212 5480
rect 29252 5440 29261 5480
rect 30067 5440 30076 5480
rect 30116 5440 30220 5480
rect 30260 5440 30269 5480
rect 30556 5440 31412 5480
rect 30556 5396 30596 5440
rect 32044 5396 32084 5524
rect 32803 5440 32812 5480
rect 32852 5440 32860 5480
rect 32900 5440 32983 5480
rect 33859 5440 33868 5480
rect 33908 5440 34444 5480
rect 34484 5440 34493 5480
rect 34636 5396 34676 5692
rect 34964 5692 34999 5723
rect 35146 5692 35155 5732
rect 35195 5692 36308 5732
rect 38563 5692 38572 5732
rect 38612 5692 38956 5732
rect 38996 5692 39436 5732
rect 39476 5692 39485 5732
rect 39689 5692 39820 5732
rect 39860 5692 39869 5732
rect 40291 5692 40300 5732
rect 40340 5692 40492 5732
rect 40532 5692 40541 5732
rect 40675 5692 40684 5732
rect 40724 5723 41780 5732
rect 40724 5692 41740 5723
rect 34924 5674 34964 5683
rect 36268 5648 36308 5692
rect 39820 5674 39860 5683
rect 41740 5674 41780 5683
rect 46278 5648 46368 5668
rect 35011 5608 35020 5648
rect 35060 5608 35260 5648
rect 35300 5608 35309 5648
rect 35465 5608 35500 5648
rect 35540 5608 35596 5648
rect 35636 5608 35645 5648
rect 35875 5608 35884 5648
rect 35924 5608 35933 5648
rect 36259 5608 36268 5648
rect 36308 5608 36317 5648
rect 36451 5608 36460 5648
rect 36500 5608 37180 5648
rect 37220 5608 37229 5648
rect 37289 5608 37420 5648
rect 37460 5608 37469 5648
rect 37865 5608 37996 5648
rect 38036 5608 38860 5648
rect 38900 5608 38909 5648
rect 42857 5608 42892 5648
rect 42932 5608 42988 5648
rect 43028 5608 43180 5648
rect 43220 5608 43229 5648
rect 43721 5608 43756 5648
rect 43796 5608 43852 5648
rect 43892 5608 43901 5648
rect 44323 5608 44332 5648
rect 44372 5608 44524 5648
rect 44564 5608 44573 5648
rect 44899 5608 44908 5648
rect 44948 5608 44957 5648
rect 45139 5608 45148 5648
rect 45188 5608 46368 5648
rect 35884 5564 35924 5608
rect 44908 5564 44948 5608
rect 46278 5588 46368 5608
rect 35788 5524 35924 5564
rect 36163 5524 36172 5564
rect 36212 5524 42412 5564
rect 42452 5524 42461 5564
rect 43180 5524 44948 5564
rect 35107 5440 35116 5480
rect 35156 5440 35644 5480
rect 35684 5440 35693 5480
rect 23020 5356 29396 5396
rect 30115 5356 30124 5396
rect 30164 5356 30596 5396
rect 31171 5356 31180 5396
rect 31220 5356 32084 5396
rect 32707 5356 32716 5396
rect 32756 5356 34676 5396
rect 35788 5396 35828 5524
rect 35897 5440 35980 5480
rect 36020 5440 36028 5480
rect 36068 5440 36077 5480
rect 38227 5440 38236 5480
rect 38276 5440 38572 5480
rect 38612 5440 38621 5480
rect 40003 5440 40012 5480
rect 40052 5440 40588 5480
rect 40628 5440 40637 5480
rect 35788 5356 42508 5396
rect 42548 5356 42557 5396
rect 23020 5312 23060 5356
rect 10636 5272 12404 5312
rect 12643 5272 12652 5312
rect 12692 5272 15532 5312
rect 15572 5272 15581 5312
rect 17347 5272 17356 5312
rect 17396 5272 18124 5312
rect 18164 5272 18173 5312
rect 18799 5272 18808 5312
rect 18848 5272 18890 5312
rect 18930 5272 18972 5312
rect 19012 5272 19054 5312
rect 19094 5272 19136 5312
rect 19176 5272 19185 5312
rect 19267 5272 19276 5312
rect 19316 5272 22484 5312
rect 22531 5272 22540 5312
rect 22580 5272 23060 5312
rect 23788 5272 27532 5312
rect 27572 5272 27581 5312
rect 12364 5144 12404 5272
rect 23788 5228 23828 5272
rect 29356 5228 29396 5356
rect 31939 5272 31948 5312
rect 31988 5272 32812 5312
rect 32852 5272 32861 5312
rect 33919 5272 33928 5312
rect 33968 5272 34010 5312
rect 34050 5272 34092 5312
rect 34132 5272 34174 5312
rect 34214 5272 34256 5312
rect 34296 5272 34305 5312
rect 35020 5272 41644 5312
rect 41684 5272 41693 5312
rect 12460 5188 14188 5228
rect 14228 5188 14237 5228
rect 14755 5188 14764 5228
rect 14804 5188 23828 5228
rect 28876 5188 29260 5228
rect 29300 5188 29309 5228
rect 29356 5188 31660 5228
rect 31700 5188 31709 5228
rect 6115 5104 6124 5144
rect 6164 5104 6173 5144
rect 8515 5104 8524 5144
rect 8564 5104 8716 5144
rect 8756 5104 8765 5144
rect 11395 5104 11404 5144
rect 11444 5104 11452 5144
rect 11492 5104 11575 5144
rect 12355 5104 12364 5144
rect 12404 5104 12413 5144
rect 12460 5060 12500 5188
rect 28876 5144 28916 5188
rect 35020 5144 35060 5272
rect 43180 5228 43220 5524
rect 44755 5440 44764 5480
rect 44804 5440 46252 5480
rect 46292 5440 46301 5480
rect 46278 5312 46368 5332
rect 46243 5272 46252 5312
rect 46292 5272 46368 5312
rect 46278 5252 46368 5272
rect 35107 5188 35116 5228
rect 35156 5188 43220 5228
rect 12739 5104 12748 5144
rect 12788 5104 14236 5144
rect 14276 5104 14285 5144
rect 14380 5104 23596 5144
rect 23636 5104 23645 5144
rect 24076 5104 28916 5144
rect 28963 5104 28972 5144
rect 29012 5104 31372 5144
rect 31412 5104 31421 5144
rect 33187 5104 33196 5144
rect 33236 5104 35060 5144
rect 36067 5104 36076 5144
rect 36116 5104 36364 5144
rect 36404 5104 36413 5144
rect 36547 5104 36556 5144
rect 36596 5104 44564 5144
rect 1036 5020 1996 5060
rect 2036 5020 2045 5060
rect 6403 5020 6412 5060
rect 6452 5020 7084 5060
rect 7124 5020 7133 5060
rect 7564 5020 12500 5060
rect 12556 5020 14188 5060
rect 14228 5020 14237 5060
rect 0 4976 90 4996
rect 1036 4976 1076 5020
rect 0 4936 1076 4976
rect 1219 4936 1228 4976
rect 1268 4936 1277 4976
rect 1481 4936 1612 4976
rect 1652 4936 1661 4976
rect 0 4916 90 4936
rect 1228 4808 1268 4936
rect 7564 4892 7604 5020
rect 9187 4936 9196 4976
rect 9236 4936 9428 4976
rect 9667 4936 9676 4976
rect 9716 4936 9772 4976
rect 9812 4936 9847 4976
rect 11561 4936 11692 4976
rect 11732 4936 11741 4976
rect 11875 4936 11884 4976
rect 11924 4936 12055 4976
rect 8812 4892 8852 4901
rect 9388 4892 9428 4936
rect 10348 4892 10388 4901
rect 12556 4892 12596 5020
rect 14380 4976 14420 5104
rect 14476 5020 14620 5060
rect 14660 5020 14668 5060
rect 14708 5020 14791 5060
rect 14956 5020 17356 5060
rect 17396 5020 17405 5060
rect 17548 5020 18412 5060
rect 18452 5020 18461 5060
rect 20332 5020 23980 5060
rect 24020 5020 24029 5060
rect 14476 4976 14516 5020
rect 12643 4936 12652 4976
rect 12692 4936 14420 4976
rect 14467 4936 14476 4976
rect 14516 4936 14525 4976
rect 14729 4936 14764 4976
rect 14804 4936 14860 4976
rect 14900 4936 14909 4976
rect 14956 4892 14996 5020
rect 5321 4852 5452 4892
rect 5492 4852 5501 4892
rect 5609 4852 5731 4892
rect 5780 4852 5789 4892
rect 6307 4852 6316 4892
rect 6356 4852 6412 4892
rect 6452 4852 6487 4892
rect 6682 4852 6691 4892
rect 6740 4852 6871 4892
rect 7433 4852 7564 4892
rect 7604 4852 7613 4892
rect 8611 4852 8620 4892
rect 8660 4852 8812 4892
rect 8812 4843 8852 4852
rect 9004 4852 9283 4892
rect 9323 4852 9332 4892
rect 9379 4852 9388 4892
rect 9428 4852 9437 4892
rect 9737 4852 9772 4892
rect 9812 4852 9868 4892
rect 9908 4852 9917 4892
rect 9964 4852 10348 4892
rect 10858 4852 10867 4892
rect 10907 4852 11212 4892
rect 11252 4852 11261 4892
rect 11587 4852 11596 4892
rect 11636 4852 12460 4892
rect 12500 4852 12509 4892
rect 13769 4852 13804 4892
rect 13844 4852 13900 4892
rect 13940 4852 13949 4892
rect 14092 4852 14996 4892
rect 15244 4892 15284 4901
rect 17548 4892 17588 5020
rect 20332 4976 20372 5020
rect 19747 4936 19756 4976
rect 19796 4936 19948 4976
rect 19988 4936 20092 4976
rect 20132 4936 20148 4976
rect 20323 4936 20332 4976
rect 20372 4936 20381 4976
rect 20428 4936 23692 4976
rect 23732 4936 23741 4976
rect 15284 4852 15532 4892
rect 15572 4852 15581 4892
rect 16361 4852 16492 4892
rect 16532 4852 16541 4892
rect 17059 4852 17068 4892
rect 17108 4852 17260 4892
rect 17300 4852 17588 4892
rect 18316 4892 18356 4901
rect 20428 4892 20468 4936
rect 18356 4852 20468 4892
rect 20515 4852 20524 4892
rect 20564 4852 21100 4892
rect 21140 4852 21149 4892
rect 22313 4852 22356 4892
rect 22396 4852 22444 4892
rect 22484 4852 22493 4892
rect 22627 4852 22636 4892
rect 22676 4852 22924 4892
rect 22964 4852 23788 4892
rect 23828 4852 23837 4892
rect 9004 4808 9044 4852
rect 9964 4808 10004 4852
rect 10348 4843 10388 4852
rect 12556 4843 12596 4852
rect 14092 4808 14132 4852
rect 15244 4843 15284 4852
rect 18316 4808 18356 4852
rect 24076 4808 24116 5104
rect 24163 5020 24172 5060
rect 24212 5020 33100 5060
rect 33140 5020 33149 5060
rect 33763 5020 33772 5060
rect 33812 5020 34732 5060
rect 34772 5020 34781 5060
rect 37324 5020 38996 5060
rect 39187 5020 39196 5060
rect 39236 5020 41204 5060
rect 41443 5020 41452 5060
rect 41492 5020 42028 5060
rect 42068 5020 42077 5060
rect 43747 5020 43756 5060
rect 43796 5020 44372 5060
rect 24259 4936 24268 4976
rect 24308 4936 25748 4976
rect 25865 4936 25996 4976
rect 26036 4936 26045 4976
rect 27043 4936 27052 4976
rect 27092 4936 28972 4976
rect 29012 4936 29021 4976
rect 29155 4936 29164 4976
rect 29204 4936 29213 4976
rect 29731 4936 29740 4976
rect 29780 4936 32524 4976
rect 32564 4936 34100 4976
rect 34147 4936 34156 4976
rect 34196 4936 34348 4976
rect 34388 4936 34397 4976
rect 24172 4892 24212 4901
rect 25708 4892 25748 4936
rect 29164 4892 29204 4936
rect 24212 4852 24556 4892
rect 24596 4852 24605 4892
rect 25708 4852 27148 4892
rect 27188 4852 27197 4892
rect 28579 4852 28588 4892
rect 28628 4852 29164 4892
rect 29204 4852 29213 4892
rect 32611 4852 32620 4892
rect 32660 4852 33100 4892
rect 33140 4852 33149 4892
rect 33283 4852 33292 4892
rect 33332 4852 33379 4892
rect 33419 4852 33868 4892
rect 33908 4852 33917 4892
rect 24172 4843 24212 4852
rect 27148 4808 27188 4852
rect 34060 4808 34100 4936
rect 36172 4892 36212 4901
rect 37324 4892 37364 5020
rect 38956 4976 38996 5020
rect 38825 4936 38956 4976
rect 38996 4936 39005 4976
rect 40169 4936 40300 4976
rect 40340 4936 40349 4976
rect 40579 4936 40588 4976
rect 40628 4936 41108 4976
rect 38572 4892 38612 4901
rect 41068 4892 41108 4936
rect 34793 4852 34924 4892
rect 34964 4852 34973 4892
rect 37315 4852 37324 4892
rect 37364 4852 37373 4892
rect 38441 4852 38572 4892
rect 38612 4852 38621 4892
rect 39427 4852 39436 4892
rect 39476 4852 40780 4892
rect 40820 4852 40829 4892
rect 41050 4852 41059 4892
rect 41099 4852 41108 4892
rect 41164 4892 41204 5020
rect 44332 4976 44372 5020
rect 44524 4976 44564 5104
rect 46278 4976 46368 4996
rect 41251 4936 41260 4976
rect 41300 4936 44092 4976
rect 44132 4936 44141 4976
rect 44323 4936 44332 4976
rect 44372 4936 44381 4976
rect 44515 4936 44524 4976
rect 44564 4936 44573 4976
rect 44899 4936 44908 4976
rect 44948 4936 44957 4976
rect 45139 4936 45148 4976
rect 45188 4936 46368 4976
rect 44908 4892 44948 4936
rect 46278 4916 46368 4936
rect 41164 4852 44236 4892
rect 44276 4852 44285 4892
rect 44524 4852 44948 4892
rect 36172 4808 36212 4852
rect 67 4768 76 4808
rect 116 4768 1268 4808
rect 1459 4768 1468 4808
rect 1508 4768 4396 4808
rect 4436 4768 4445 4808
rect 5827 4768 5836 4808
rect 5876 4768 6796 4808
rect 6836 4768 8524 4808
rect 8564 4768 8573 4808
rect 8995 4768 9004 4808
rect 9044 4768 9053 4808
rect 9955 4768 9964 4808
rect 10004 4768 10013 4808
rect 10444 4768 12404 4808
rect 10444 4724 10484 4768
rect 12364 4724 12404 4768
rect 12940 4768 14132 4808
rect 14227 4768 14236 4808
rect 14276 4768 15188 4808
rect 15811 4768 15820 4808
rect 15860 4768 18356 4808
rect 18403 4768 18412 4808
rect 18452 4768 18644 4808
rect 18691 4768 18700 4808
rect 18740 4768 19996 4808
rect 20036 4768 21580 4808
rect 21620 4768 21629 4808
rect 22444 4768 24116 4808
rect 24259 4768 24268 4808
rect 24308 4768 27052 4808
rect 27092 4768 27101 4808
rect 27148 4768 29404 4808
rect 29444 4768 29453 4808
rect 33187 4768 33196 4808
rect 33236 4768 33484 4808
rect 33524 4768 33533 4808
rect 33667 4768 33676 4808
rect 33716 4768 33916 4808
rect 33956 4768 33965 4808
rect 34060 4768 37996 4808
rect 38036 4768 38045 4808
rect 12940 4724 12980 4768
rect 15148 4724 15188 4768
rect 18604 4724 18644 4768
rect 22444 4724 22484 4768
rect 38572 4724 38612 4852
rect 40867 4768 40876 4808
rect 40916 4768 41164 4808
rect 41204 4768 41213 4808
rect 41260 4768 44084 4808
rect 1843 4684 1852 4724
rect 1892 4684 5684 4724
rect 6019 4684 6028 4724
rect 6068 4684 10484 4724
rect 10889 4684 11020 4724
rect 11060 4684 11069 4724
rect 12115 4684 12124 4724
rect 12164 4684 12172 4724
rect 12212 4684 12295 4724
rect 12364 4684 12980 4724
rect 13315 4684 13324 4724
rect 13364 4684 13612 4724
rect 13652 4684 13661 4724
rect 15043 4684 15052 4724
rect 15092 4684 15101 4724
rect 15148 4684 16724 4724
rect 18211 4684 18220 4724
rect 18260 4684 18508 4724
rect 18548 4684 18557 4724
rect 18604 4684 22484 4724
rect 22531 4684 22540 4724
rect 22580 4684 23060 4724
rect 24067 4684 24076 4724
rect 24116 4684 24364 4724
rect 24404 4684 24413 4724
rect 26227 4684 26236 4724
rect 26276 4684 29068 4724
rect 29108 4684 29117 4724
rect 29251 4684 29260 4724
rect 29300 4684 29452 4724
rect 29492 4684 30124 4724
rect 30164 4684 38612 4724
rect 38755 4684 38764 4724
rect 38804 4684 38935 4724
rect 40531 4684 40540 4724
rect 40580 4684 41068 4724
rect 41108 4684 41117 4724
rect 0 4640 90 4660
rect 0 4600 76 4640
rect 116 4600 125 4640
rect 0 4580 90 4600
rect 5644 4556 5684 4684
rect 15052 4640 15092 4684
rect 16684 4640 16724 4684
rect 23020 4640 23060 4684
rect 41260 4640 41300 4768
rect 42857 4684 42979 4724
rect 43028 4684 43267 4724
rect 43307 4684 43316 4724
rect 43721 4684 43843 4724
rect 43892 4684 43901 4724
rect 8035 4600 8044 4640
rect 8084 4600 9100 4640
rect 9140 4600 9149 4640
rect 9475 4600 9484 4640
rect 9524 4600 15092 4640
rect 15235 4600 15244 4640
rect 15284 4600 15820 4640
rect 15860 4600 15869 4640
rect 16684 4600 22924 4640
rect 22964 4600 22973 4640
rect 23020 4600 31660 4640
rect 31700 4600 31709 4640
rect 35683 4600 35692 4640
rect 35732 4600 41300 4640
rect 44044 4640 44084 4768
rect 44524 4640 44564 4852
rect 44755 4684 44764 4724
rect 44804 4684 44813 4724
rect 44044 4600 44564 4640
rect 44764 4640 44804 4684
rect 46278 4640 46368 4660
rect 44764 4600 46368 4640
rect 46278 4580 46368 4600
rect 4919 4516 4928 4556
rect 4968 4516 5010 4556
rect 5050 4516 5092 4556
rect 5132 4516 5174 4556
rect 5214 4516 5256 4556
rect 5296 4516 5305 4556
rect 5644 4516 17260 4556
rect 17300 4516 17309 4556
rect 20039 4516 20048 4556
rect 20088 4516 20130 4556
rect 20170 4516 20212 4556
rect 20252 4516 20294 4556
rect 20334 4516 20376 4556
rect 20416 4516 20425 4556
rect 23971 4516 23980 4556
rect 24020 4516 28492 4556
rect 28532 4516 28541 4556
rect 35159 4516 35168 4556
rect 35208 4516 35250 4556
rect 35290 4516 35332 4556
rect 35372 4516 35414 4556
rect 35454 4516 35496 4556
rect 35536 4516 35545 4556
rect 38179 4516 38188 4556
rect 38228 4516 43756 4556
rect 43796 4516 43805 4556
rect 8611 4432 8620 4472
rect 8660 4432 9964 4472
rect 10004 4432 10013 4472
rect 10531 4432 10540 4472
rect 10580 4432 14476 4472
rect 14516 4432 14525 4472
rect 15139 4432 15148 4472
rect 15188 4432 32908 4472
rect 32948 4432 32957 4472
rect 39907 4432 39916 4472
rect 39956 4432 42260 4472
rect 42220 4388 42260 4432
rect 8323 4348 8332 4388
rect 8372 4348 13324 4388
rect 13364 4348 13373 4388
rect 15811 4348 15820 4388
rect 15860 4348 21332 4388
rect 21379 4348 21388 4388
rect 21428 4348 23788 4388
rect 23828 4348 23837 4388
rect 24019 4348 24028 4388
rect 24068 4348 24172 4388
rect 24212 4348 24221 4388
rect 24355 4348 24364 4388
rect 24404 4348 32236 4388
rect 32276 4348 32285 4388
rect 33283 4348 33292 4388
rect 33332 4348 40588 4388
rect 40628 4348 40637 4388
rect 42202 4348 42211 4388
rect 42251 4348 42499 4388
rect 42539 4348 42787 4388
rect 42827 4348 42836 4388
rect 43546 4348 43555 4388
rect 43595 4348 44227 4388
rect 44267 4348 44276 4388
rect 0 4304 90 4324
rect 0 4264 1612 4304
rect 1652 4264 1661 4304
rect 2860 4264 6164 4304
rect 6211 4264 6220 4304
rect 6260 4264 7124 4304
rect 0 4244 90 4264
rect 2860 4220 2900 4264
rect 6124 4220 6164 4264
rect 7084 4220 7124 4264
rect 7180 4264 7948 4304
rect 7988 4264 7997 4304
rect 8140 4264 8756 4304
rect 8842 4264 8851 4304
rect 8891 4264 8908 4304
rect 8948 4264 9031 4304
rect 9161 4264 9244 4304
rect 9284 4264 9292 4304
rect 9332 4264 9341 4304
rect 9667 4264 9676 4304
rect 9716 4264 9868 4304
rect 9908 4264 9917 4304
rect 11251 4264 11260 4304
rect 11300 4264 11692 4304
rect 11732 4264 11741 4304
rect 13699 4264 13708 4304
rect 13748 4264 14668 4304
rect 14708 4264 14717 4304
rect 15139 4264 15148 4304
rect 15188 4264 15244 4304
rect 15284 4264 15319 4304
rect 18377 4264 18412 4304
rect 18452 4264 18508 4304
rect 18548 4264 18557 4304
rect 20899 4264 20908 4304
rect 20948 4264 20957 4304
rect 7180 4220 7220 4264
rect 1516 4180 2900 4220
rect 4771 4180 4780 4220
rect 4820 4180 4829 4220
rect 5897 4180 6028 4220
rect 6068 4180 6077 4220
rect 6124 4180 6892 4220
rect 6932 4180 6941 4220
rect 7066 4180 7075 4220
rect 7115 4180 7124 4220
rect 7171 4180 7180 4220
rect 7220 4180 7229 4220
rect 7555 4180 7564 4220
rect 7604 4180 8044 4220
rect 8084 4180 8093 4220
rect 8140 4211 8180 4264
rect 8716 4220 8756 4264
rect 20908 4220 20948 4264
rect 21292 4220 21332 4348
rect 46278 4304 46368 4324
rect 22217 4264 22348 4304
rect 22388 4264 22397 4304
rect 23491 4264 23500 4304
rect 23540 4264 31124 4304
rect 31171 4264 31180 4304
rect 31220 4264 32620 4304
rect 32660 4264 32669 4304
rect 33091 4264 33100 4304
rect 33140 4264 34924 4304
rect 34964 4264 34973 4304
rect 38755 4264 38764 4304
rect 38804 4264 38900 4304
rect 38947 4264 38956 4304
rect 38996 4264 39044 4304
rect 39139 4264 39148 4304
rect 39188 4264 39340 4304
rect 39380 4264 39389 4304
rect 40291 4264 40300 4304
rect 40340 4264 41684 4304
rect 43721 4264 43852 4304
rect 43892 4264 43901 4304
rect 45139 4264 45148 4304
rect 45188 4264 46368 4304
rect 29740 4220 29780 4264
rect 1516 4136 1556 4180
rect 4780 4136 4820 4180
rect 6028 4162 6068 4171
rect 8489 4180 8620 4220
rect 8660 4180 8669 4220
rect 8716 4180 9428 4220
rect 9475 4180 9484 4220
rect 9524 4180 9655 4220
rect 9754 4180 9763 4220
rect 9803 4180 10060 4220
rect 10100 4180 10109 4220
rect 11971 4180 11980 4220
rect 12020 4180 12268 4220
rect 12308 4180 12317 4220
rect 13123 4180 13132 4220
rect 13172 4211 13708 4220
rect 13172 4180 13516 4211
rect 8140 4162 8180 4171
rect 8620 4162 8660 4171
rect 9388 4136 9428 4180
rect 9772 4136 9812 4180
rect 13556 4180 13708 4211
rect 13748 4180 13757 4220
rect 15364 4180 15373 4220
rect 15413 4180 15436 4220
rect 15476 4180 15553 4220
rect 15619 4180 15628 4220
rect 15668 4180 15799 4220
rect 16867 4180 16876 4220
rect 16916 4180 16925 4220
rect 17923 4180 17932 4220
rect 17972 4211 18164 4220
rect 17972 4180 18124 4211
rect 13516 4162 13556 4171
rect 13708 4136 13748 4180
rect 67 4096 76 4136
rect 116 4096 1228 4136
rect 1268 4096 1277 4136
rect 1459 4096 1468 4136
rect 1508 4096 1556 4136
rect 1603 4096 1612 4136
rect 1652 4096 1661 4136
rect 3977 4096 4108 4136
rect 4148 4096 4820 4136
rect 6281 4096 6412 4136
rect 6452 4096 6461 4136
rect 7529 4096 7660 4136
rect 7700 4096 7709 4136
rect 8873 4096 9004 4136
rect 9044 4096 9053 4136
rect 9388 4096 9812 4136
rect 10195 4096 10204 4136
rect 10244 4096 10348 4136
rect 10388 4096 10397 4136
rect 10889 4096 11020 4136
rect 11060 4096 11069 4136
rect 13708 4096 13948 4136
rect 13988 4096 13997 4136
rect 14179 4096 14188 4136
rect 14228 4096 15820 4136
rect 15860 4096 15869 4136
rect 0 3968 90 3988
rect 0 3928 76 3968
rect 116 3928 125 3968
rect 0 3908 90 3928
rect 0 3632 90 3652
rect 1612 3632 1652 4096
rect 16876 4052 16916 4180
rect 18124 4162 18164 4171
rect 18700 4211 18740 4220
rect 18787 4180 18796 4220
rect 18836 4180 19948 4220
rect 19988 4180 20852 4220
rect 20899 4180 20908 4220
rect 20948 4180 20995 4220
rect 21292 4211 24940 4220
rect 21292 4180 22156 4211
rect 18700 4136 18740 4171
rect 20812 4136 20852 4180
rect 22196 4180 24364 4211
rect 22156 4162 22196 4171
rect 24404 4180 24940 4211
rect 24980 4180 24989 4220
rect 25123 4180 25132 4220
rect 25172 4180 25324 4220
rect 25364 4180 25612 4220
rect 25652 4180 25661 4220
rect 25900 4211 26900 4220
rect 25900 4180 25996 4211
rect 24364 4162 24404 4171
rect 25900 4136 25940 4180
rect 26036 4180 26900 4211
rect 27113 4180 27244 4220
rect 27284 4180 27628 4220
rect 27668 4180 27677 4220
rect 28745 4180 28876 4220
rect 28916 4180 28925 4220
rect 29731 4180 29740 4220
rect 29780 4180 29789 4220
rect 30988 4211 31028 4220
rect 25996 4162 26036 4171
rect 18700 4096 19948 4136
rect 19988 4096 20140 4136
rect 20180 4096 20189 4136
rect 20419 4096 20428 4136
rect 20468 4096 20524 4136
rect 20564 4096 20599 4136
rect 20812 4096 22060 4136
rect 22100 4096 22109 4136
rect 22243 4096 22252 4136
rect 22292 4096 23500 4136
rect 23540 4096 23549 4136
rect 23657 4096 23692 4136
rect 23732 4096 23788 4136
rect 23828 4096 23837 4136
rect 23884 4096 24308 4136
rect 24547 4096 24556 4136
rect 24596 4096 25940 4136
rect 26860 4136 26900 4180
rect 28876 4162 28916 4171
rect 30988 4136 31028 4171
rect 26860 4096 28588 4136
rect 28628 4096 28637 4136
rect 29155 4096 29164 4136
rect 29204 4096 29452 4136
rect 29492 4096 31028 4136
rect 31084 4136 31124 4264
rect 31939 4180 31948 4220
rect 31988 4180 32611 4220
rect 32651 4180 32660 4220
rect 32707 4180 32716 4220
rect 32756 4180 32812 4220
rect 32852 4180 32887 4220
rect 33084 4180 33093 4220
rect 33133 4180 33292 4220
rect 33332 4180 33341 4220
rect 33676 4211 33868 4220
rect 33716 4180 33868 4211
rect 33908 4180 33917 4220
rect 34156 4211 34348 4220
rect 33676 4162 33716 4171
rect 34196 4180 34348 4211
rect 34388 4180 34397 4220
rect 34156 4162 34196 4171
rect 34924 4136 34964 4264
rect 38860 4220 38900 4264
rect 39004 4220 39044 4264
rect 41644 4220 41684 4264
rect 46278 4244 46368 4264
rect 37123 4180 37132 4220
rect 37172 4180 37228 4220
rect 37268 4180 37303 4220
rect 37987 4180 37996 4220
rect 38036 4211 38516 4220
rect 38036 4180 38476 4211
rect 38860 4180 38908 4220
rect 38948 4180 38957 4220
rect 39004 4180 39235 4220
rect 39275 4180 39284 4220
rect 39331 4180 39340 4220
rect 39380 4211 40436 4220
rect 39380 4180 40396 4211
rect 38476 4162 38516 4171
rect 41635 4180 41644 4220
rect 41684 4180 41693 4220
rect 42979 4180 42988 4220
rect 43028 4180 43468 4220
rect 43508 4180 43517 4220
rect 40396 4162 40436 4171
rect 31084 4096 33004 4136
rect 33044 4096 33053 4136
rect 33187 4096 33196 4136
rect 33236 4096 33388 4136
rect 33428 4096 33437 4136
rect 34601 4096 34732 4136
rect 34772 4096 34781 4136
rect 34915 4096 34924 4136
rect 34964 4096 34973 4136
rect 35971 4096 35980 4136
rect 36020 4096 36172 4136
rect 36212 4096 37516 4136
rect 37556 4096 37565 4136
rect 39523 4096 39532 4136
rect 39572 4096 39772 4136
rect 39812 4096 39821 4136
rect 40003 4096 40012 4136
rect 40052 4096 40061 4136
rect 41897 4096 42028 4136
rect 42068 4096 42077 4136
rect 43049 4096 43084 4136
rect 43124 4096 43180 4136
rect 43220 4096 43284 4136
rect 44393 4096 44524 4136
rect 44564 4096 44573 4136
rect 44777 4096 44908 4136
rect 44948 4096 44957 4136
rect 23884 4052 23924 4096
rect 24268 4052 24308 4096
rect 40012 4052 40052 4096
rect 1843 4012 1852 4052
rect 1892 4012 13364 4052
rect 13603 4012 13612 4052
rect 13652 4012 16684 4052
rect 16724 4012 16916 4052
rect 18307 4012 18316 4052
rect 18356 4012 19276 4052
rect 19316 4012 19325 4052
rect 20131 4012 20140 4052
rect 20180 4012 20380 4052
rect 20420 4012 20524 4052
rect 20564 4012 20580 4052
rect 20755 4012 20764 4052
rect 20804 4012 22484 4052
rect 23107 4012 23116 4052
rect 23156 4012 23924 4052
rect 23971 4012 23980 4052
rect 24020 4012 24172 4052
rect 24212 4012 24221 4052
rect 24268 4012 34492 4052
rect 34532 4012 34541 4052
rect 34627 4012 34636 4052
rect 34676 4012 38476 4052
rect 38516 4012 38525 4052
rect 38659 4012 38668 4052
rect 38708 4012 39436 4052
rect 39476 4012 39485 4052
rect 39619 4012 39628 4052
rect 39668 4012 40052 4052
rect 44755 4012 44764 4052
rect 44804 4012 45620 4052
rect 13324 3968 13364 4012
rect 22444 3968 22484 4012
rect 45580 3968 45620 4012
rect 46278 3968 46368 3988
rect 4339 3928 4348 3968
rect 4388 3928 6548 3968
rect 6643 3928 6652 3968
rect 6692 3928 9812 3968
rect 10579 3928 10588 3968
rect 10628 3928 13228 3968
rect 13268 3928 13277 3968
rect 13324 3928 14708 3968
rect 14825 3928 14860 3968
rect 14900 3928 14956 3968
rect 14996 3928 15005 3968
rect 15619 3928 15628 3968
rect 15668 3928 17452 3968
rect 17492 3928 17501 3968
rect 18316 3928 20428 3968
rect 20468 3928 20908 3968
rect 20948 3928 20957 3968
rect 22444 3928 23060 3968
rect 25673 3928 25708 3968
rect 25748 3928 25804 3968
rect 25844 3928 25853 3968
rect 28937 3928 28972 3968
rect 29012 3928 29068 3968
rect 29108 3928 29117 3968
rect 29203 3928 29212 3968
rect 29252 3928 29740 3968
rect 29780 3928 29789 3968
rect 30211 3928 30220 3968
rect 30260 3928 32140 3968
rect 32180 3928 32189 3968
rect 32515 3928 32524 3968
rect 32564 3928 34387 3968
rect 34427 3928 34436 3968
rect 35155 3928 35164 3968
rect 35204 3928 35596 3968
rect 35636 3928 35645 3968
rect 36211 3928 36220 3968
rect 36260 3928 39628 3968
rect 39668 3928 39677 3968
rect 40073 3928 40204 3968
rect 40244 3928 40253 3968
rect 41657 3928 41740 3968
rect 41780 3928 41788 3968
rect 41828 3928 41837 3968
rect 45580 3928 46368 3968
rect 3679 3760 3688 3800
rect 3728 3760 3770 3800
rect 3810 3760 3852 3800
rect 3892 3760 3934 3800
rect 3974 3760 4016 3800
rect 4056 3760 4065 3800
rect 6508 3716 6548 3928
rect 9772 3884 9812 3928
rect 14668 3884 14708 3928
rect 18316 3884 18356 3928
rect 23020 3884 23060 3928
rect 46278 3908 46368 3928
rect 7843 3844 7852 3884
rect 7892 3844 9676 3884
rect 9716 3844 9725 3884
rect 9772 3844 14380 3884
rect 14420 3844 14429 3884
rect 14668 3844 18356 3884
rect 18403 3844 18412 3884
rect 18452 3844 18604 3884
rect 18644 3844 18653 3884
rect 18700 3844 22636 3884
rect 22676 3844 22685 3884
rect 23020 3844 31852 3884
rect 31892 3844 31901 3884
rect 32323 3844 32332 3884
rect 32372 3844 44948 3884
rect 18700 3800 18740 3844
rect 6883 3760 6892 3800
rect 6932 3760 11116 3800
rect 11156 3760 11165 3800
rect 14092 3760 18740 3800
rect 18799 3760 18808 3800
rect 18848 3760 18890 3800
rect 18930 3760 18972 3800
rect 19012 3760 19054 3800
rect 19094 3760 19136 3800
rect 19176 3760 19185 3800
rect 19459 3760 19468 3800
rect 19508 3760 32524 3800
rect 32564 3760 32573 3800
rect 33919 3760 33928 3800
rect 33968 3760 34010 3800
rect 34050 3760 34092 3800
rect 34132 3760 34174 3800
rect 34214 3760 34256 3800
rect 34296 3760 34305 3800
rect 35395 3760 35404 3800
rect 35444 3760 44428 3800
rect 44468 3760 44477 3800
rect 6508 3676 13708 3716
rect 13748 3676 13757 3716
rect 14092 3632 14132 3760
rect 14179 3676 14188 3716
rect 14228 3676 29260 3716
rect 29300 3676 29309 3716
rect 29356 3676 30604 3716
rect 30644 3676 30653 3716
rect 36931 3676 36940 3716
rect 36980 3676 44276 3716
rect 29356 3632 29396 3676
rect 0 3592 1652 3632
rect 2860 3592 14132 3632
rect 14563 3592 14572 3632
rect 14612 3592 14620 3632
rect 14660 3592 14743 3632
rect 15427 3592 15436 3632
rect 15476 3592 15628 3632
rect 15668 3592 18796 3632
rect 18836 3592 18845 3632
rect 18892 3592 24844 3632
rect 24884 3592 24893 3632
rect 25123 3592 25132 3632
rect 25172 3592 29396 3632
rect 29635 3592 29644 3632
rect 29684 3592 40684 3632
rect 40724 3592 40733 3632
rect 42211 3592 42220 3632
rect 42260 3592 43996 3632
rect 44036 3592 44045 3632
rect 0 3572 90 3592
rect 2860 3548 2900 3592
rect 1459 3508 1468 3548
rect 1508 3508 1748 3548
rect 1843 3508 1852 3548
rect 1892 3508 2900 3548
rect 5347 3508 5356 3548
rect 5396 3508 6316 3548
rect 6356 3508 6365 3548
rect 8131 3508 8140 3548
rect 8180 3508 8189 3548
rect 8563 3508 8572 3548
rect 8612 3508 12460 3548
rect 12500 3508 12509 3548
rect 12556 3508 13612 3548
rect 13652 3508 13661 3548
rect 13795 3508 13804 3548
rect 13844 3508 14036 3548
rect 14153 3508 14236 3548
rect 14276 3508 14284 3548
rect 14324 3508 14333 3548
rect 15004 3508 15724 3548
rect 15764 3508 15773 3548
rect 16684 3508 18604 3548
rect 18644 3508 18653 3548
rect 67 3424 76 3464
rect 116 3424 1228 3464
rect 1268 3424 1277 3464
rect 1603 3424 1612 3464
rect 1652 3424 1661 3464
rect 0 3296 90 3316
rect 0 3256 76 3296
rect 116 3256 125 3296
rect 0 3236 90 3256
rect 1612 3128 1652 3424
rect 1708 3212 1748 3508
rect 8140 3464 8180 3508
rect 12556 3464 12596 3508
rect 13996 3464 14036 3508
rect 8140 3424 8332 3464
rect 8372 3424 8381 3464
rect 8515 3424 8524 3464
rect 8564 3424 8716 3464
rect 8756 3424 8765 3464
rect 8812 3424 12596 3464
rect 12931 3424 12940 3464
rect 12980 3424 13516 3464
rect 13556 3424 13565 3464
rect 13987 3424 13996 3464
rect 14036 3424 14045 3464
rect 14729 3424 14860 3464
rect 14900 3424 14909 3464
rect 5164 3380 5204 3389
rect 3523 3340 3532 3380
rect 3572 3340 3916 3380
rect 3956 3340 4108 3380
rect 4148 3340 4157 3380
rect 4771 3340 4780 3380
rect 4820 3340 5164 3380
rect 5204 3340 6988 3380
rect 7028 3340 7037 3380
rect 7337 3340 7468 3380
rect 7508 3340 7517 3380
rect 7651 3340 7660 3380
rect 7700 3340 7747 3380
rect 7787 3340 7831 3380
rect 5164 3331 5204 3340
rect 7721 3256 7852 3296
rect 7892 3256 7901 3296
rect 8812 3212 8852 3424
rect 12652 3380 12692 3389
rect 11395 3340 11404 3380
rect 11444 3340 11980 3380
rect 12020 3340 12029 3380
rect 12556 3340 12652 3380
rect 12556 3296 12596 3340
rect 12652 3331 12692 3340
rect 12844 3340 13132 3380
rect 13172 3340 13181 3380
rect 13289 3340 13411 3380
rect 13460 3340 13469 3380
rect 12844 3296 12884 3340
rect 9283 3256 9292 3296
rect 9332 3256 12364 3296
rect 12404 3256 12413 3296
rect 12547 3256 12556 3296
rect 12596 3256 12605 3296
rect 12835 3256 12844 3296
rect 12884 3256 12893 3296
rect 13315 3256 13324 3296
rect 13364 3256 13516 3296
rect 13556 3256 13565 3296
rect 15004 3212 15044 3508
rect 15148 3424 15340 3464
rect 15380 3424 15389 3464
rect 15497 3424 15628 3464
rect 15668 3424 15677 3464
rect 15148 3380 15188 3424
rect 16684 3413 16724 3508
rect 18892 3464 18932 3592
rect 18979 3508 18988 3548
rect 19028 3508 19412 3548
rect 24643 3508 24652 3548
rect 24692 3508 25076 3548
rect 29539 3508 29548 3548
rect 29588 3508 30068 3548
rect 31817 3508 31948 3548
rect 31988 3508 31997 3548
rect 33475 3508 33484 3548
rect 33524 3508 33908 3548
rect 35011 3508 35020 3548
rect 35060 3508 43372 3548
rect 43412 3508 43421 3548
rect 19372 3464 19412 3508
rect 25036 3464 25076 3508
rect 30028 3464 30068 3508
rect 33868 3464 33908 3508
rect 44236 3464 44276 3676
rect 44908 3464 44948 3844
rect 46278 3632 46368 3652
rect 45139 3592 45148 3632
rect 45188 3592 46368 3632
rect 46278 3572 46368 3592
rect 18019 3424 18028 3464
rect 18068 3424 18932 3464
rect 19363 3424 19372 3464
rect 19412 3424 19421 3464
rect 20515 3424 20524 3464
rect 20564 3424 20948 3464
rect 20995 3424 21004 3464
rect 21044 3424 21175 3464
rect 23020 3424 24692 3464
rect 24739 3424 24748 3464
rect 24788 3424 24796 3464
rect 24836 3424 24919 3464
rect 25027 3424 25036 3464
rect 25076 3424 25085 3464
rect 25219 3424 25228 3464
rect 25268 3424 25708 3464
rect 25748 3424 25757 3464
rect 29539 3424 29548 3464
rect 29588 3424 29788 3464
rect 29828 3424 29837 3464
rect 30019 3424 30028 3464
rect 30068 3424 30077 3464
rect 30211 3424 30220 3464
rect 30260 3424 31796 3464
rect 32131 3424 32140 3464
rect 32180 3424 33812 3464
rect 33859 3424 33868 3464
rect 33908 3424 33917 3464
rect 34819 3424 34828 3464
rect 34868 3424 37324 3464
rect 37364 3424 37373 3464
rect 37507 3424 37516 3464
rect 37556 3424 38324 3464
rect 38441 3424 38572 3464
rect 38612 3424 38621 3464
rect 39235 3424 39244 3464
rect 39284 3424 43892 3464
rect 44227 3424 44236 3464
rect 44276 3424 44285 3464
rect 44611 3424 44620 3464
rect 44660 3424 44669 3464
rect 44899 3424 44908 3464
rect 44948 3424 44957 3464
rect 16204 3380 16244 3389
rect 15130 3340 15139 3380
rect 15179 3340 15188 3380
rect 15235 3340 15244 3380
rect 15284 3340 15293 3380
rect 15593 3340 15724 3380
rect 15764 3340 15773 3380
rect 16073 3340 16204 3380
rect 16244 3340 16253 3380
rect 20908 3380 20948 3424
rect 23020 3380 23060 3424
rect 16684 3364 16724 3373
rect 16780 3340 18316 3380
rect 18356 3340 18365 3380
rect 18460 3340 18595 3380
rect 18635 3340 18644 3380
rect 18883 3340 18892 3380
rect 18932 3340 20812 3380
rect 20852 3340 20861 3380
rect 20908 3340 23060 3380
rect 23945 3340 23980 3380
rect 24020 3340 24076 3380
rect 24116 3340 24125 3380
rect 24250 3340 24259 3380
rect 24308 3340 24460 3380
rect 24500 3340 24509 3380
rect 15244 3296 15284 3340
rect 16204 3331 16244 3340
rect 15244 3256 16012 3296
rect 16052 3256 16061 3296
rect 16780 3212 16820 3340
rect 18460 3212 18500 3340
rect 24652 3296 24692 3424
rect 27628 3380 27668 3389
rect 31756 3380 31796 3424
rect 33772 3380 33812 3424
rect 37424 3380 37464 3389
rect 38284 3380 38324 3424
rect 39148 3380 39188 3389
rect 43852 3380 43892 3424
rect 44620 3380 44660 3424
rect 26249 3340 26380 3380
rect 26420 3340 26429 3380
rect 28745 3340 28876 3380
rect 28916 3340 28925 3380
rect 29033 3340 29155 3380
rect 29204 3340 29932 3380
rect 29972 3340 29981 3380
rect 30403 3340 30412 3380
rect 30452 3340 30508 3380
rect 30548 3340 30583 3380
rect 31843 3340 31852 3380
rect 31892 3340 32812 3380
rect 32852 3340 32861 3380
rect 33082 3340 33091 3380
rect 33131 3340 33292 3380
rect 33332 3340 33341 3380
rect 33772 3340 35788 3380
rect 35828 3340 35837 3380
rect 36041 3340 36172 3380
rect 36212 3340 36221 3380
rect 36940 3340 37424 3380
rect 27628 3296 27668 3340
rect 31756 3296 31796 3340
rect 18569 3256 18700 3296
rect 18740 3256 18749 3296
rect 19123 3256 19132 3296
rect 19172 3256 19372 3296
rect 19412 3256 19421 3296
rect 20140 3256 21484 3296
rect 21524 3256 21533 3296
rect 23011 3256 23020 3296
rect 23060 3256 24364 3296
rect 24404 3256 24413 3296
rect 24652 3256 29204 3296
rect 29251 3256 29260 3296
rect 29300 3256 29356 3296
rect 29396 3256 29431 3296
rect 29644 3256 31180 3296
rect 31220 3256 31229 3296
rect 31756 3256 32812 3296
rect 32852 3256 32861 3296
rect 33020 3256 33100 3296
rect 33140 3256 33180 3296
rect 33220 3256 33271 3296
rect 33619 3256 33628 3296
rect 33668 3256 33676 3296
rect 33716 3256 33799 3296
rect 20140 3212 20180 3256
rect 29164 3212 29204 3256
rect 29644 3212 29684 3256
rect 36940 3212 36980 3340
rect 37424 3331 37464 3340
rect 37612 3340 38083 3380
rect 38123 3340 38132 3380
rect 38179 3340 38188 3380
rect 38228 3340 38237 3380
rect 38284 3340 38668 3380
rect 38708 3340 38717 3380
rect 39658 3340 39667 3380
rect 39707 3340 40204 3380
rect 40244 3340 40253 3380
rect 40675 3340 40684 3380
rect 40724 3340 41356 3380
rect 41396 3340 42988 3380
rect 43028 3340 43756 3380
rect 43796 3340 43805 3380
rect 43852 3340 44660 3380
rect 37612 3296 37652 3340
rect 38188 3296 38228 3340
rect 39148 3296 39188 3340
rect 46278 3296 46368 3316
rect 37603 3256 37612 3296
rect 37652 3256 37661 3296
rect 37891 3256 37900 3296
rect 37940 3256 38228 3296
rect 38371 3256 38380 3296
rect 38420 3256 38668 3296
rect 38708 3256 39188 3296
rect 39244 3256 42604 3296
rect 42644 3256 42653 3296
rect 44131 3256 44140 3296
rect 44180 3256 44380 3296
rect 44420 3256 44429 3296
rect 45187 3256 45196 3296
rect 45236 3256 46368 3296
rect 1708 3172 8852 3212
rect 8947 3172 8956 3212
rect 8996 3172 15044 3212
rect 15427 3172 15436 3212
rect 15476 3172 16820 3212
rect 16867 3172 16876 3212
rect 16916 3172 17047 3212
rect 17657 3172 17740 3212
rect 17780 3172 17788 3212
rect 17828 3172 17837 3212
rect 18460 3172 19948 3212
rect 19988 3172 20180 3212
rect 21235 3172 21244 3212
rect 21284 3172 24692 3212
rect 25337 3172 25420 3212
rect 25460 3172 25468 3212
rect 25508 3172 25517 3212
rect 27689 3172 27820 3212
rect 27860 3172 27869 3212
rect 29164 3172 29684 3212
rect 29932 3172 35404 3212
rect 35444 3172 35453 3212
rect 35500 3172 39148 3212
rect 39188 3172 39197 3212
rect 24652 3128 24692 3172
rect 29932 3128 29972 3172
rect 35500 3128 35540 3172
rect 39244 3128 39284 3256
rect 46278 3236 46368 3256
rect 39689 3172 39820 3212
rect 39860 3172 39869 3212
rect 40195 3172 40204 3212
rect 40244 3172 41635 3212
rect 41675 3172 41684 3212
rect 41801 3172 41923 3212
rect 41972 3172 42211 3212
rect 42251 3172 42499 3212
rect 42539 3172 42787 3212
rect 42827 3172 43075 3212
rect 43124 3172 43363 3212
rect 43403 3172 43412 3212
rect 76 3088 1652 3128
rect 6019 3088 6028 3128
rect 6068 3088 8812 3128
rect 8852 3088 9292 3128
rect 9332 3088 9341 3128
rect 11587 3088 11596 3128
rect 11636 3088 12556 3128
rect 12596 3088 15244 3128
rect 15284 3088 15293 3128
rect 15715 3088 15724 3128
rect 15764 3088 24596 3128
rect 24652 3088 29972 3128
rect 31171 3088 31180 3128
rect 31220 3088 35540 3128
rect 35587 3088 35596 3128
rect 35636 3088 39284 3128
rect 39619 3088 39628 3128
rect 39668 3088 43756 3128
rect 43796 3088 43805 3128
rect 76 2980 116 3088
rect 24556 3044 24596 3088
rect 4919 3004 4928 3044
rect 4968 3004 5010 3044
rect 5050 3004 5092 3044
rect 5132 3004 5174 3044
rect 5214 3004 5256 3044
rect 5296 3004 5305 3044
rect 8899 3004 8908 3044
rect 8948 3004 15340 3044
rect 15380 3004 15389 3044
rect 15436 3004 18892 3044
rect 18932 3004 18941 3044
rect 20039 3004 20048 3044
rect 20088 3004 20130 3044
rect 20170 3004 20212 3044
rect 20252 3004 20294 3044
rect 20334 3004 20376 3044
rect 20416 3004 20425 3044
rect 24556 3004 25132 3044
rect 25172 3004 25181 3044
rect 29059 3004 29068 3044
rect 29108 3004 35020 3044
rect 35060 3004 35069 3044
rect 35159 3004 35168 3044
rect 35208 3004 35250 3044
rect 35290 3004 35332 3044
rect 35372 3004 35414 3044
rect 35454 3004 35496 3044
rect 35536 3004 35545 3044
rect 35779 3004 35788 3044
rect 35828 3004 44908 3044
rect 44948 3004 44957 3044
rect 0 2920 116 2980
rect 15436 2960 15476 3004
rect 46278 2960 46368 2980
rect 5740 2920 15476 2960
rect 16867 2920 16876 2960
rect 16916 2920 25804 2960
rect 25844 2920 25853 2960
rect 27360 2920 27436 2960
rect 27476 2920 27485 2960
rect 29251 2920 29260 2960
rect 29300 2920 39572 2960
rect 39907 2920 39916 2960
rect 39956 2920 40204 2960
rect 40244 2920 40253 2960
rect 41164 2920 41932 2960
rect 41972 2920 41981 2960
rect 42316 2920 43220 2960
rect 0 2900 90 2920
rect 5740 2876 5780 2920
rect 27436 2876 27476 2920
rect 39532 2876 39572 2920
rect 41164 2876 41204 2920
rect 42316 2876 42356 2920
rect 43180 2876 43220 2920
rect 45580 2920 46368 2960
rect 5587 2836 5596 2876
rect 5636 2836 5780 2876
rect 7171 2836 7180 2876
rect 7220 2836 7468 2876
rect 7508 2836 7517 2876
rect 8611 2836 8620 2876
rect 8660 2836 9004 2876
rect 9044 2836 9053 2876
rect 9571 2836 9580 2876
rect 9620 2836 9628 2876
rect 9668 2836 9751 2876
rect 11081 2836 11212 2876
rect 11252 2836 11261 2876
rect 11404 2836 14036 2876
rect 15305 2836 15436 2876
rect 15476 2836 15485 2876
rect 15619 2836 15628 2876
rect 15668 2836 15820 2876
rect 15860 2836 15869 2876
rect 16003 2836 16012 2876
rect 16052 2836 17068 2876
rect 17108 2836 17117 2876
rect 19564 2836 20908 2876
rect 20948 2836 20957 2876
rect 21676 2836 24844 2876
rect 24884 2836 24893 2876
rect 25123 2836 25132 2876
rect 25172 2836 27476 2876
rect 27523 2836 27532 2876
rect 27572 2836 28876 2876
rect 28916 2836 28925 2876
rect 29443 2836 29452 2876
rect 29492 2836 30028 2876
rect 30068 2836 30077 2876
rect 34051 2836 34060 2876
rect 34100 2836 34348 2876
rect 34388 2836 34397 2876
rect 35212 2836 39092 2876
rect 39532 2836 40771 2876
rect 40811 2836 41059 2876
rect 41099 2836 41204 2876
rect 41251 2836 41260 2876
rect 41300 2836 41308 2876
rect 41348 2836 41431 2876
rect 41635 2836 41644 2876
rect 41684 2836 41692 2876
rect 41732 2836 41815 2876
rect 42019 2836 42028 2876
rect 42068 2836 42356 2876
rect 42403 2836 42412 2876
rect 42452 2836 42460 2876
rect 42500 2836 42583 2876
rect 42953 2836 43075 2876
rect 43124 2836 43133 2876
rect 43180 2836 44660 2876
rect 45065 2836 45148 2876
rect 45188 2836 45196 2876
rect 45236 2836 45245 2876
rect 11404 2792 11444 2836
rect 1459 2752 1468 2792
rect 1508 2752 10636 2792
rect 10676 2752 10685 2792
rect 10732 2752 11444 2792
rect 11491 2752 11500 2792
rect 11540 2752 13748 2792
rect 5356 2668 5740 2708
rect 5780 2668 5836 2708
rect 5876 2668 6892 2708
rect 6932 2668 6941 2708
rect 6988 2699 7028 2708
rect 0 2624 90 2644
rect 5356 2624 5396 2668
rect 7433 2668 7564 2708
rect 7604 2668 7613 2708
rect 8681 2668 8812 2708
rect 8852 2668 8861 2708
rect 9641 2668 9772 2708
rect 9812 2668 9821 2708
rect 6988 2624 7028 2659
rect 8812 2650 8852 2659
rect 10732 2624 10772 2752
rect 11404 2708 11444 2752
rect 13708 2708 13748 2752
rect 13996 2708 14036 2836
rect 16492 2752 18604 2792
rect 18644 2752 18700 2792
rect 18740 2752 18804 2792
rect 19180 2752 19276 2792
rect 19316 2752 19325 2792
rect 10889 2668 11020 2708
rect 11060 2668 11069 2708
rect 11395 2668 11404 2708
rect 11444 2668 11453 2708
rect 12652 2699 12940 2708
rect 0 2584 1228 2624
rect 1268 2584 1277 2624
rect 1603 2584 1612 2624
rect 1652 2584 1661 2624
rect 1708 2584 1996 2624
rect 2036 2584 2045 2624
rect 5347 2584 5356 2624
rect 5396 2584 5405 2624
rect 6857 2584 6988 2624
rect 7028 2584 7037 2624
rect 9257 2584 9388 2624
rect 9428 2584 10772 2624
rect 11020 2624 11060 2659
rect 12692 2668 12940 2699
rect 12980 2668 12989 2708
rect 13315 2668 13324 2708
rect 13364 2668 13373 2708
rect 13444 2668 13453 2708
rect 13493 2668 13652 2708
rect 13699 2668 13708 2708
rect 13748 2668 13757 2708
rect 13987 2668 13996 2708
rect 14036 2668 14045 2708
rect 15244 2699 15284 2708
rect 12652 2624 12692 2659
rect 13324 2624 13364 2668
rect 11020 2584 12692 2624
rect 12940 2584 13228 2624
rect 13268 2584 13277 2624
rect 13324 2584 13420 2624
rect 13460 2584 13469 2624
rect 0 2564 90 2584
rect 0 2288 90 2308
rect 1612 2288 1652 2584
rect 0 2248 1652 2288
rect 0 2228 90 2248
rect 1708 2120 1748 2584
rect 6988 2540 7028 2584
rect 12940 2540 12980 2584
rect 2227 2500 2236 2540
rect 2276 2500 2860 2540
rect 2900 2500 2909 2540
rect 6988 2500 10540 2540
rect 10580 2500 11596 2540
rect 11636 2500 11645 2540
rect 11692 2500 12980 2540
rect 13612 2540 13652 2668
rect 15331 2668 15340 2708
rect 15380 2668 15715 2708
rect 15755 2668 15764 2708
rect 15811 2668 15820 2708
rect 15860 2668 16012 2708
rect 16052 2668 16061 2708
rect 16195 2668 16204 2708
rect 16244 2668 16396 2708
rect 16436 2668 16445 2708
rect 15244 2624 15284 2659
rect 16492 2624 16532 2752
rect 19180 2708 19220 2752
rect 16649 2668 16780 2708
rect 16820 2668 16829 2708
rect 16963 2668 16972 2708
rect 17012 2699 17300 2708
rect 17012 2668 17260 2699
rect 16780 2650 16820 2659
rect 18089 2668 18220 2708
rect 18260 2668 18269 2708
rect 18490 2668 18499 2708
rect 18539 2668 18988 2708
rect 19028 2668 19037 2708
rect 19162 2668 19171 2708
rect 19211 2668 19220 2708
rect 19267 2668 19276 2708
rect 19316 2668 19468 2708
rect 19508 2668 19517 2708
rect 17260 2650 17300 2659
rect 19564 2624 19604 2836
rect 21676 2792 21716 2836
rect 35212 2792 35252 2836
rect 19939 2752 19948 2792
rect 19988 2752 20180 2792
rect 20227 2752 20236 2792
rect 20276 2752 21716 2792
rect 22627 2752 22636 2792
rect 22676 2752 23156 2792
rect 24355 2752 24364 2792
rect 24404 2752 24788 2792
rect 24979 2752 24988 2792
rect 25028 2752 25036 2792
rect 25076 2752 25159 2792
rect 25315 2752 25324 2792
rect 25364 2752 26132 2792
rect 26563 2752 26572 2792
rect 26612 2752 28532 2792
rect 30115 2752 30124 2792
rect 30164 2752 30556 2792
rect 30596 2752 30605 2792
rect 30700 2752 30988 2792
rect 31028 2752 31037 2792
rect 32323 2752 32332 2792
rect 32372 2752 35252 2792
rect 35491 2752 35500 2792
rect 35540 2752 35740 2792
rect 35780 2752 35789 2792
rect 36067 2752 36076 2792
rect 36116 2752 37900 2792
rect 37940 2752 37949 2792
rect 38083 2752 38092 2792
rect 38132 2752 38141 2792
rect 38633 2752 38764 2792
rect 38804 2752 38813 2792
rect 38947 2752 38956 2792
rect 38996 2752 39005 2792
rect 20140 2708 20180 2752
rect 23116 2708 23156 2752
rect 24748 2708 24788 2752
rect 26092 2708 26132 2752
rect 19651 2668 19660 2708
rect 19700 2668 19988 2708
rect 20140 2699 20276 2708
rect 20140 2668 20236 2699
rect 19948 2624 19988 2668
rect 20585 2668 20716 2708
rect 20756 2668 20765 2708
rect 20995 2668 21004 2708
rect 21044 2668 21196 2708
rect 21236 2668 21245 2708
rect 21571 2668 21580 2708
rect 21620 2699 22924 2708
rect 21620 2668 22444 2699
rect 20236 2650 20276 2659
rect 20716 2650 20756 2659
rect 22484 2668 22924 2699
rect 22964 2668 22973 2708
rect 23098 2668 23107 2708
rect 23147 2668 23156 2708
rect 23203 2668 23212 2708
rect 23252 2668 23383 2708
rect 23587 2668 23596 2708
rect 23636 2668 23884 2708
rect 23924 2668 23933 2708
rect 24172 2699 24556 2708
rect 22444 2650 22484 2659
rect 24212 2668 24556 2699
rect 24596 2668 24605 2708
rect 24652 2699 24692 2708
rect 24172 2650 24212 2659
rect 24748 2668 25324 2708
rect 25364 2668 25373 2708
rect 25444 2668 25453 2708
rect 25493 2668 25516 2708
rect 25556 2668 25633 2708
rect 25699 2668 25708 2708
rect 25748 2668 25879 2708
rect 26083 2668 26092 2708
rect 26132 2668 26141 2708
rect 26275 2668 26284 2708
rect 26324 2699 27532 2708
rect 26324 2668 27340 2699
rect 24652 2624 24692 2659
rect 27380 2668 27532 2699
rect 27572 2668 27581 2708
rect 27811 2668 27820 2708
rect 27860 2668 28291 2708
rect 28331 2668 28340 2708
rect 28387 2668 28396 2708
rect 28436 2668 28445 2708
rect 27340 2650 27380 2659
rect 15244 2584 15628 2624
rect 15668 2584 15677 2624
rect 16195 2584 16204 2624
rect 16244 2584 16300 2624
rect 16340 2584 16532 2624
rect 17731 2584 17740 2624
rect 17780 2584 19604 2624
rect 19747 2584 19756 2624
rect 19796 2584 19805 2624
rect 19948 2584 20044 2624
rect 20084 2584 20093 2624
rect 23683 2584 23692 2624
rect 23732 2584 24076 2624
rect 24116 2584 24125 2624
rect 24652 2584 27244 2624
rect 27284 2584 27293 2624
rect 27907 2584 27916 2624
rect 27956 2584 28300 2624
rect 28340 2584 28349 2624
rect 19756 2540 19796 2584
rect 13612 2500 15724 2540
rect 15764 2500 15773 2540
rect 18979 2500 18988 2540
rect 19028 2500 19796 2540
rect 19939 2500 19948 2540
rect 19988 2500 25996 2540
rect 26036 2500 26045 2540
rect 26179 2500 26188 2540
rect 26228 2500 27676 2540
rect 27716 2500 27725 2540
rect 11692 2456 11732 2500
rect 19756 2456 19796 2500
rect 28396 2456 28436 2668
rect 28492 2624 28532 2752
rect 30700 2708 30740 2752
rect 38092 2708 38132 2752
rect 28649 2668 28780 2708
rect 28820 2668 29108 2708
rect 29155 2668 29164 2708
rect 29204 2699 29396 2708
rect 29204 2668 29356 2699
rect 29068 2624 29108 2668
rect 29356 2650 29396 2659
rect 29836 2699 30740 2708
rect 29876 2668 30740 2699
rect 31049 2668 31180 2708
rect 31220 2668 31229 2708
rect 32035 2668 32044 2708
rect 32084 2668 32428 2708
rect 32468 2668 32477 2708
rect 32611 2668 32620 2708
rect 32660 2668 32669 2708
rect 32803 2668 32812 2708
rect 32852 2699 33908 2708
rect 32852 2668 33868 2699
rect 29836 2650 29876 2659
rect 31180 2650 31220 2659
rect 32620 2624 32660 2668
rect 34793 2668 34924 2708
rect 34964 2668 34973 2708
rect 35057 2668 35116 2708
rect 35156 2668 35179 2708
rect 35219 2668 35237 2708
rect 35290 2668 35299 2708
rect 35339 2668 35348 2708
rect 36643 2668 36652 2708
rect 36692 2668 37132 2708
rect 37172 2668 37181 2708
rect 37315 2668 37324 2708
rect 37364 2699 37940 2708
rect 37364 2668 37900 2699
rect 33868 2650 33908 2659
rect 35308 2624 35348 2668
rect 36652 2624 36692 2668
rect 38092 2668 38380 2708
rect 38420 2668 38429 2708
rect 38537 2668 38659 2708
rect 38708 2668 38717 2708
rect 37900 2650 37940 2659
rect 38956 2624 38996 2752
rect 39052 2708 39092 2836
rect 39139 2752 39148 2792
rect 39188 2752 42356 2792
rect 42595 2752 42604 2792
rect 42644 2752 44564 2792
rect 39052 2668 41588 2708
rect 41548 2624 41588 2668
rect 42316 2624 42356 2752
rect 44524 2624 44564 2752
rect 44620 2624 44660 2836
rect 45580 2792 45620 2920
rect 46278 2900 46368 2920
rect 44755 2752 44764 2792
rect 44804 2752 45620 2792
rect 46278 2624 46368 2644
rect 28492 2584 28684 2624
rect 28724 2584 28876 2624
rect 28916 2584 28925 2624
rect 29068 2584 29260 2624
rect 29300 2584 29309 2624
rect 30281 2584 30412 2624
rect 30452 2584 30461 2624
rect 30691 2584 30700 2624
rect 30740 2584 30796 2624
rect 30836 2584 30871 2624
rect 31843 2584 31852 2624
rect 31892 2584 32660 2624
rect 33379 2584 33388 2624
rect 33428 2584 33812 2624
rect 34435 2584 34444 2624
rect 34484 2584 35348 2624
rect 35596 2584 35980 2624
rect 36020 2584 36029 2624
rect 36259 2584 36268 2624
rect 36308 2584 36692 2624
rect 37996 2584 38996 2624
rect 39091 2584 39100 2624
rect 39140 2584 39436 2624
rect 39476 2584 39485 2624
rect 41539 2584 41548 2624
rect 41588 2584 41597 2624
rect 41801 2584 41932 2624
rect 41972 2584 41981 2624
rect 42067 2584 42076 2624
rect 42116 2584 42124 2624
rect 42164 2584 42247 2624
rect 42307 2584 42316 2624
rect 42356 2584 42365 2624
rect 42691 2584 42700 2624
rect 42740 2584 42749 2624
rect 43075 2584 43084 2624
rect 43124 2584 43372 2624
rect 43412 2584 43421 2624
rect 43625 2584 43756 2624
rect 43796 2584 43805 2624
rect 43852 2584 44332 2624
rect 44372 2584 44381 2624
rect 44515 2584 44524 2624
rect 44564 2584 44573 2624
rect 44620 2584 44908 2624
rect 44948 2584 44957 2624
rect 45187 2584 45196 2624
rect 45236 2584 46368 2624
rect 33772 2540 33812 2584
rect 35596 2540 35636 2584
rect 37996 2540 38036 2584
rect 42700 2540 42740 2584
rect 43852 2540 43892 2584
rect 46278 2564 46368 2584
rect 31363 2500 31372 2540
rect 31412 2500 32044 2540
rect 32084 2500 32093 2540
rect 32227 2500 32236 2540
rect 32276 2500 33580 2540
rect 33620 2500 33629 2540
rect 33772 2500 34676 2540
rect 35587 2500 35596 2540
rect 35636 2500 35645 2540
rect 35692 2500 38036 2540
rect 38851 2500 38860 2540
rect 38900 2500 42740 2540
rect 43180 2500 43892 2540
rect 43987 2500 43996 2540
rect 44036 2500 45100 2540
rect 45140 2500 45149 2540
rect 34636 2456 34676 2500
rect 35692 2456 35732 2500
rect 43180 2456 43220 2500
rect 1843 2416 1852 2456
rect 1892 2416 2092 2456
rect 2132 2416 2141 2456
rect 5155 2416 5164 2456
rect 5204 2416 8428 2456
rect 8468 2416 8477 2456
rect 8707 2416 8716 2456
rect 8756 2416 11020 2456
rect 11060 2416 11069 2456
rect 11203 2416 11212 2456
rect 11252 2416 11732 2456
rect 12713 2416 12844 2456
rect 12884 2416 12893 2456
rect 12940 2416 13036 2456
rect 13076 2416 13085 2456
rect 16579 2416 16588 2456
rect 16628 2416 17491 2456
rect 17531 2416 17540 2456
rect 17971 2416 17980 2456
rect 18020 2416 18508 2456
rect 18548 2416 18557 2456
rect 18883 2416 18892 2456
rect 18932 2416 18941 2456
rect 19756 2416 23060 2456
rect 23203 2416 23212 2456
rect 23252 2416 24980 2456
rect 4108 2332 12748 2372
rect 12788 2332 12797 2372
rect 3679 2248 3688 2288
rect 3728 2248 3770 2288
rect 3810 2248 3852 2288
rect 3892 2248 3934 2288
rect 3974 2248 4016 2288
rect 4056 2248 4065 2288
rect 172 2080 1748 2120
rect 1843 2080 1852 2120
rect 1892 2080 1900 2120
rect 1940 2080 2023 2120
rect 2611 2080 2620 2120
rect 2660 2080 3532 2120
rect 3572 2080 3581 2120
rect 0 1952 90 1972
rect 172 1952 212 2080
rect 4108 2036 4148 2332
rect 12940 2288 12980 2416
rect 18892 2372 18932 2416
rect 23020 2372 23060 2416
rect 24940 2372 24980 2416
rect 25132 2416 28436 2456
rect 29827 2416 29836 2456
rect 29876 2416 30172 2456
rect 30212 2416 30221 2456
rect 34636 2416 35732 2456
rect 36499 2416 36508 2456
rect 36548 2416 38668 2456
rect 38708 2416 38717 2456
rect 38947 2416 38956 2456
rect 38996 2416 39196 2456
rect 39236 2416 39245 2456
rect 39331 2416 39340 2456
rect 39380 2416 43220 2456
rect 43529 2416 43612 2456
rect 43652 2416 43660 2456
rect 43700 2416 43709 2456
rect 43948 2416 44092 2456
rect 44132 2416 44141 2456
rect 25132 2372 25172 2416
rect 13219 2332 13228 2372
rect 13268 2332 16396 2372
rect 16436 2332 18548 2372
rect 18892 2332 19276 2372
rect 19316 2332 19325 2372
rect 19372 2332 22924 2372
rect 22964 2332 22973 2372
rect 23020 2332 24844 2372
rect 24884 2332 24893 2372
rect 24940 2332 25172 2372
rect 25507 2332 25516 2372
rect 25556 2332 29684 2372
rect 29731 2332 29740 2372
rect 29780 2332 29876 2372
rect 31555 2332 31564 2372
rect 31604 2332 33388 2372
rect 33428 2332 33437 2372
rect 33820 2332 37324 2372
rect 37364 2332 37373 2372
rect 39043 2332 39052 2372
rect 39092 2332 41932 2372
rect 41972 2332 41981 2372
rect 5827 2248 5836 2288
rect 5876 2248 12652 2288
rect 12692 2248 12701 2288
rect 12844 2248 12980 2288
rect 5452 2164 5684 2204
rect 5452 2120 5492 2164
rect 4243 2080 4252 2120
rect 4292 2080 5492 2120
rect 5644 2120 5684 2164
rect 5836 2164 7852 2204
rect 7892 2164 7901 2204
rect 8620 2164 8908 2204
rect 8948 2164 8957 2204
rect 9004 2164 11980 2204
rect 12020 2164 12029 2204
rect 5836 2120 5876 2164
rect 8620 2120 8660 2164
rect 9004 2120 9044 2164
rect 12844 2120 12884 2248
rect 18508 2204 18548 2332
rect 18799 2248 18808 2288
rect 18848 2248 18890 2288
rect 18930 2248 18972 2288
rect 19012 2248 19054 2288
rect 19094 2248 19136 2288
rect 19176 2248 19185 2288
rect 19372 2204 19412 2332
rect 19459 2248 19468 2288
rect 19508 2248 22732 2288
rect 22772 2248 22781 2288
rect 22924 2248 24940 2288
rect 24980 2248 24989 2288
rect 25123 2248 25132 2288
rect 25172 2248 28780 2288
rect 28820 2248 28829 2288
rect 22924 2204 22964 2248
rect 29644 2204 29684 2332
rect 29836 2288 29876 2332
rect 33820 2288 33860 2332
rect 43948 2288 43988 2416
rect 46278 2288 46368 2308
rect 29836 2248 33860 2288
rect 33919 2248 33928 2288
rect 33968 2248 34010 2288
rect 34050 2248 34092 2288
rect 34132 2248 34174 2288
rect 34214 2248 34256 2288
rect 34296 2248 34305 2288
rect 40291 2248 40300 2288
rect 40340 2248 41260 2288
rect 41300 2248 41309 2288
rect 41443 2248 41452 2288
rect 41492 2248 43988 2288
rect 44716 2248 46368 2288
rect 13228 2164 15340 2204
rect 15380 2164 15389 2204
rect 15523 2164 15532 2204
rect 15572 2164 16780 2204
rect 16820 2164 16829 2204
rect 16925 2164 16972 2204
rect 17012 2164 17021 2204
rect 18508 2164 19412 2204
rect 19468 2164 22964 2204
rect 23212 2164 29548 2204
rect 29588 2164 29597 2204
rect 29644 2164 33772 2204
rect 33812 2164 33821 2204
rect 34819 2164 34828 2204
rect 34868 2164 36076 2204
rect 36116 2164 36125 2204
rect 36172 2164 37612 2204
rect 37652 2164 37661 2204
rect 37891 2164 37900 2204
rect 37940 2164 42124 2204
rect 42164 2164 42173 2204
rect 42499 2164 42508 2204
rect 42548 2164 44044 2204
rect 44084 2164 44093 2204
rect 5644 2080 5876 2120
rect 5923 2080 5932 2120
rect 5972 2080 5980 2120
rect 6020 2080 6103 2120
rect 6211 2080 6220 2120
rect 6260 2080 8660 2120
rect 8755 2080 8764 2120
rect 8804 2080 9044 2120
rect 9139 2080 9148 2120
rect 9188 2080 10348 2120
rect 10388 2080 10397 2120
rect 10723 2080 10732 2120
rect 10772 2080 11500 2120
rect 11540 2080 11549 2120
rect 12844 2080 12932 2120
rect 1219 1996 1228 2036
rect 1268 1996 2420 2036
rect 3475 1996 3484 2036
rect 3524 1996 4148 2036
rect 4819 1996 4828 2036
rect 4868 1996 5836 2036
rect 5876 1996 5885 2036
rect 6124 1996 7756 2036
rect 7796 1996 7805 2036
rect 8044 1996 8660 2036
rect 9955 1996 9964 2036
rect 10004 1996 12220 2036
rect 12260 1996 12269 2036
rect 2380 1952 2420 1996
rect 6124 1952 6164 1996
rect 8044 1952 8084 1996
rect 0 1912 212 1952
rect 1219 1912 1228 1952
rect 1268 1912 1277 1952
rect 1411 1912 1420 1952
rect 1460 1912 1612 1952
rect 1652 1912 1661 1952
rect 1987 1912 1996 1952
rect 2036 1912 2045 1952
rect 2371 1912 2380 1952
rect 2420 1912 2429 1952
rect 3113 1912 3148 1952
rect 3188 1912 3244 1952
rect 3284 1912 3293 1952
rect 3881 1912 3916 1952
rect 3956 1912 4012 1952
rect 4052 1912 4061 1952
rect 4579 1912 4588 1952
rect 4628 1912 4684 1952
rect 4724 1912 4759 1952
rect 4963 1912 4972 1952
rect 5012 1912 5021 1952
rect 5155 1912 5164 1952
rect 5204 1912 5212 1952
rect 5252 1912 5335 1952
rect 5386 1912 5395 1952
rect 5435 1912 5684 1952
rect 5731 1912 5740 1952
rect 5780 1912 5911 1952
rect 6115 1912 6124 1952
rect 6164 1912 6173 1952
rect 6499 1912 6508 1952
rect 6548 1912 7564 1952
rect 7604 1912 8084 1952
rect 8515 1912 8524 1952
rect 8564 1912 8573 1952
rect 0 1892 90 1912
rect 1228 1784 1268 1912
rect 1996 1868 2036 1912
rect 1315 1828 1324 1868
rect 1364 1828 2036 1868
rect 4972 1868 5012 1912
rect 5644 1868 5684 1912
rect 4972 1828 5452 1868
rect 5492 1828 5501 1868
rect 5644 1828 6220 1868
rect 6260 1828 6269 1868
rect 6508 1784 6548 1912
rect 8140 1868 8180 1877
rect 6761 1828 6892 1868
rect 6932 1828 6941 1868
rect 8180 1828 8468 1868
rect 8140 1819 8180 1828
rect 67 1744 76 1784
rect 116 1744 1268 1784
rect 1459 1744 1468 1784
rect 1508 1744 6548 1784
rect 8428 1700 8468 1828
rect 8524 1784 8564 1912
rect 8620 1868 8660 1996
rect 12892 1952 12932 2080
rect 8899 1912 8908 1952
rect 8948 1912 10060 1952
rect 10100 1912 10109 1952
rect 10793 1912 10828 1952
rect 10868 1912 10924 1952
rect 10964 1912 10973 1952
rect 11491 1912 11500 1952
rect 11540 1912 11596 1952
rect 11636 1912 11671 1952
rect 11875 1912 11884 1952
rect 11924 1912 12404 1952
rect 12451 1912 12460 1952
rect 12500 1912 12509 1952
rect 12595 1912 12604 1952
rect 12644 1912 12652 1952
rect 12692 1912 12775 1952
rect 12835 1912 12844 1952
rect 12884 1912 12932 1952
rect 10540 1868 10580 1877
rect 12364 1868 12404 1912
rect 8620 1828 9292 1868
rect 9332 1828 9341 1868
rect 10409 1828 10540 1868
rect 10580 1828 10589 1868
rect 12355 1828 12364 1868
rect 12404 1828 12413 1868
rect 10540 1819 10580 1828
rect 12460 1784 12500 1912
rect 12835 1828 12844 1868
rect 12884 1828 13132 1868
rect 13172 1828 13181 1868
rect 8524 1744 9292 1784
rect 9332 1744 9341 1784
rect 11731 1744 11740 1784
rect 11780 1744 11980 1784
rect 12020 1744 12029 1784
rect 12115 1744 12124 1784
rect 12164 1744 12404 1784
rect 12460 1744 13132 1784
rect 13172 1744 13181 1784
rect 12364 1700 12404 1744
rect 2227 1660 2236 1700
rect 2276 1660 2804 1700
rect 5587 1660 5596 1700
rect 5636 1660 6124 1700
rect 6164 1660 6173 1700
rect 6355 1660 6364 1700
rect 6404 1660 6644 1700
rect 6739 1660 6748 1700
rect 6788 1660 7180 1700
rect 7220 1660 7229 1700
rect 8323 1660 8332 1700
rect 8372 1660 8381 1700
rect 8428 1660 8716 1700
rect 8756 1660 8765 1700
rect 11155 1660 11164 1700
rect 11204 1660 11500 1700
rect 11540 1660 11549 1700
rect 12364 1660 13036 1700
rect 13076 1660 13085 1700
rect 0 1616 90 1636
rect 0 1576 76 1616
rect 116 1576 125 1616
rect 0 1556 90 1576
rect 2764 1364 2804 1660
rect 6604 1616 6644 1660
rect 8332 1616 8372 1660
rect 13228 1616 13268 2164
rect 16972 2120 17012 2164
rect 19468 2120 19508 2164
rect 13891 2080 13900 2120
rect 13940 2080 13948 2120
rect 13988 2080 14071 2120
rect 16483 2080 16492 2120
rect 16532 2080 16540 2120
rect 16580 2080 16663 2120
rect 16963 2080 16972 2120
rect 17012 2080 17021 2120
rect 17155 2080 17164 2120
rect 17204 2080 19508 2120
rect 20585 2080 20620 2120
rect 20660 2080 20716 2120
rect 20756 2080 20765 2120
rect 20995 2080 21004 2120
rect 21044 2080 22828 2120
rect 22868 2080 22877 2120
rect 13795 1996 13804 2036
rect 13844 1996 13853 2036
rect 14611 1996 14620 2036
rect 14660 1996 16684 2036
rect 16724 1996 16733 2036
rect 17923 1996 17932 2036
rect 17972 1996 22636 2036
rect 22676 1996 22685 2036
rect 13804 1952 13844 1996
rect 23212 1952 23252 2164
rect 36172 2120 36212 2164
rect 44716 2120 44756 2248
rect 46278 2228 46368 2248
rect 25027 2080 25036 2120
rect 25076 2080 25460 2120
rect 25987 2080 25996 2120
rect 26036 2080 34060 2120
rect 34100 2080 34109 2120
rect 34243 2080 34252 2120
rect 34292 2080 34924 2120
rect 34964 2080 34973 2120
rect 35155 2080 35164 2120
rect 35204 2080 36212 2120
rect 36979 2080 36988 2120
rect 37028 2080 37804 2120
rect 37844 2080 37853 2120
rect 38083 2080 38092 2120
rect 38132 2080 39004 2120
rect 39044 2080 39053 2120
rect 40361 2080 40444 2120
rect 40484 2080 40492 2120
rect 40532 2080 40541 2120
rect 40963 2080 40972 2120
rect 41012 2080 41884 2120
rect 41924 2080 41933 2120
rect 42835 2080 42844 2120
rect 42884 2080 44756 2120
rect 24643 1996 24652 2036
rect 24692 1996 25076 2036
rect 25171 1996 25180 2036
rect 25220 1996 25228 2036
rect 25268 1996 25351 2036
rect 25036 1952 25076 1996
rect 25420 1952 25460 2080
rect 25891 1996 25900 2036
rect 25940 1996 27380 2036
rect 28675 1996 28684 2036
rect 28724 1996 30412 2036
rect 30452 1996 30461 2036
rect 31603 1996 31612 2036
rect 31652 1996 43028 2036
rect 27340 1952 27380 1996
rect 42988 1952 43028 1996
rect 43084 1996 43796 2036
rect 13411 1912 13420 1952
rect 13460 1912 13556 1952
rect 13804 1912 14188 1952
rect 14228 1912 14237 1952
rect 14371 1912 14380 1952
rect 14420 1912 14429 1952
rect 14633 1912 14668 1952
rect 14708 1912 14764 1952
rect 14804 1912 14813 1952
rect 14995 1912 15004 1952
rect 15044 1912 15436 1952
rect 15476 1912 15485 1952
rect 15619 1912 15628 1952
rect 15668 1912 15677 1952
rect 15811 1912 15820 1952
rect 15860 1912 15991 1952
rect 16195 1912 16204 1952
rect 16244 1912 16300 1952
rect 16340 1912 16375 1952
rect 16579 1912 16588 1952
rect 16628 1912 16780 1952
rect 16820 1912 16829 1952
rect 18115 1912 18124 1952
rect 18164 1912 18604 1952
rect 18644 1912 18653 1952
rect 18979 1912 18988 1952
rect 19028 1912 19037 1952
rect 19267 1912 19276 1952
rect 19316 1912 19564 1952
rect 19604 1912 19613 1952
rect 19721 1912 19756 1952
rect 19796 1912 19852 1952
rect 19892 1912 19901 1952
rect 20105 1912 20236 1952
rect 20276 1912 20285 1952
rect 21667 1912 21676 1952
rect 21716 1912 22636 1952
rect 22676 1912 22685 1952
rect 23212 1912 23251 1952
rect 23291 1912 23300 1952
rect 23369 1912 23500 1952
rect 23540 1912 23549 1952
rect 23596 1912 24116 1952
rect 24739 1912 24748 1952
rect 24788 1912 24796 1952
rect 24836 1912 24919 1952
rect 25027 1912 25036 1952
rect 25076 1912 25085 1952
rect 25411 1912 25420 1952
rect 25460 1912 25469 1952
rect 25673 1912 25804 1952
rect 25844 1912 25853 1952
rect 27340 1912 30028 1952
rect 30068 1912 30077 1952
rect 31241 1912 31372 1952
rect 31412 1912 31421 1952
rect 31721 1912 31852 1952
rect 31892 1912 31901 1952
rect 32009 1912 32092 1952
rect 32132 1912 32140 1952
rect 32180 1912 32189 1952
rect 34243 1912 34252 1952
rect 34292 1912 34924 1952
rect 34964 1912 34973 1952
rect 36163 1912 36172 1952
rect 36212 1912 36748 1952
rect 36788 1912 36797 1952
rect 37699 1912 37708 1952
rect 37748 1912 39244 1952
rect 39284 1912 39293 1952
rect 39907 1912 39916 1952
rect 39956 1912 40300 1952
rect 40340 1912 40349 1952
rect 40675 1912 40684 1952
rect 40724 1912 40733 1952
rect 40780 1912 42124 1952
rect 42164 1912 42173 1952
rect 42595 1912 42604 1952
rect 42644 1912 42653 1952
rect 42979 1912 42988 1952
rect 43028 1912 43037 1952
rect 13402 1828 13411 1868
rect 13451 1828 13460 1868
rect 13420 1784 13460 1828
rect 13516 1784 13556 1912
rect 14380 1868 14420 1912
rect 13891 1828 13900 1868
rect 13940 1828 14420 1868
rect 15628 1868 15668 1912
rect 18988 1868 19028 1912
rect 20812 1868 20852 1877
rect 23596 1868 23636 1912
rect 24076 1868 24116 1912
rect 27244 1868 27284 1877
rect 31852 1868 31892 1912
rect 34060 1868 34100 1877
rect 40684 1868 40724 1912
rect 15628 1828 16204 1868
rect 16244 1828 16253 1868
rect 17155 1828 17164 1868
rect 17204 1828 17356 1868
rect 17396 1828 17405 1868
rect 18019 1828 18028 1868
rect 18068 1828 18412 1868
rect 18452 1828 18461 1868
rect 18988 1828 19372 1868
rect 19412 1828 19421 1868
rect 20611 1828 20620 1868
rect 20660 1828 20812 1868
rect 20899 1828 20908 1868
rect 20948 1828 22060 1868
rect 22100 1828 22109 1868
rect 22243 1828 22252 1868
rect 22292 1828 23636 1868
rect 23683 1828 23692 1868
rect 23732 1828 23741 1868
rect 23849 1828 23980 1868
rect 24020 1828 24029 1868
rect 24076 1828 24235 1868
rect 24275 1828 24284 1868
rect 24346 1828 24355 1868
rect 24404 1828 24535 1868
rect 25987 1828 25996 1868
rect 26036 1828 26045 1868
rect 27084 1828 27148 1868
rect 27188 1828 27244 1868
rect 27284 1828 27820 1868
rect 27860 1828 27869 1868
rect 28003 1828 28012 1868
rect 28052 1828 28061 1868
rect 28282 1828 28291 1868
rect 28331 1828 28684 1868
rect 28724 1828 28733 1868
rect 28841 1828 28972 1868
rect 29012 1828 29021 1868
rect 29129 1828 29251 1868
rect 29300 1828 29309 1868
rect 29683 1828 29692 1868
rect 29732 1828 30700 1868
rect 30740 1828 30749 1868
rect 31852 1828 32812 1868
rect 32852 1828 32861 1868
rect 35587 1828 35596 1868
rect 35636 1828 40724 1868
rect 20812 1819 20852 1828
rect 23692 1784 23732 1828
rect 6604 1576 8276 1616
rect 8332 1576 13268 1616
rect 13324 1744 13460 1784
rect 13507 1744 13516 1784
rect 13556 1744 15532 1784
rect 15572 1744 15581 1784
rect 16435 1744 16444 1784
rect 16484 1744 16972 1784
rect 17012 1744 17021 1784
rect 19219 1744 19228 1784
rect 19268 1744 19852 1784
rect 19892 1744 19901 1784
rect 21676 1744 23596 1784
rect 23636 1744 23645 1784
rect 23692 1744 24076 1784
rect 24116 1744 24125 1784
rect 24643 1744 24652 1784
rect 24692 1744 25564 1784
rect 25604 1744 25613 1784
rect 13324 1616 13364 1744
rect 15379 1660 15388 1700
rect 15428 1660 15436 1700
rect 15476 1660 15559 1700
rect 16051 1660 16060 1700
rect 16100 1660 16204 1700
rect 16244 1660 16253 1700
rect 18835 1660 18844 1700
rect 18884 1660 19220 1700
rect 19315 1660 19324 1700
rect 19364 1660 19564 1700
rect 19604 1660 19613 1700
rect 19939 1660 19948 1700
rect 19988 1660 20092 1700
rect 20132 1660 20141 1700
rect 20467 1660 20476 1700
rect 20516 1660 21580 1700
rect 21620 1660 21629 1700
rect 19180 1616 19220 1660
rect 21676 1616 21716 1744
rect 25996 1700 26036 1828
rect 27244 1819 27284 1828
rect 28012 1784 28052 1828
rect 34060 1784 34100 1828
rect 40780 1784 40820 1912
rect 42604 1868 42644 1912
rect 43084 1868 43124 1996
rect 43756 1952 43796 1996
rect 43852 1996 44756 2036
rect 45065 1996 45148 2036
rect 45188 1996 45196 2036
rect 45236 1996 45245 2036
rect 43241 1912 43372 1952
rect 43412 1912 43421 1952
rect 43747 1912 43756 1952
rect 43796 1912 43805 1952
rect 41059 1828 41068 1868
rect 41108 1828 42644 1868
rect 42691 1828 42700 1868
rect 42740 1828 43124 1868
rect 43171 1828 43180 1868
rect 43220 1828 43756 1868
rect 43796 1828 43805 1868
rect 43852 1784 43892 1996
rect 44716 1952 44756 1996
rect 46278 1952 46368 1972
rect 44035 1912 44044 1952
rect 44084 1912 44092 1952
rect 44132 1912 44215 1952
rect 44323 1912 44332 1952
rect 44372 1912 44381 1952
rect 44707 1912 44716 1952
rect 44756 1912 44908 1952
rect 44948 1912 44957 1952
rect 45091 1912 45100 1952
rect 45140 1912 46368 1952
rect 44332 1868 44372 1912
rect 46278 1892 46368 1912
rect 43939 1828 43948 1868
rect 43988 1828 44372 1868
rect 27427 1744 27436 1784
rect 27476 1744 28052 1784
rect 28387 1744 28396 1784
rect 28436 1744 28780 1784
rect 28820 1744 29356 1784
rect 29396 1744 29405 1784
rect 29539 1744 29548 1784
rect 29588 1744 29924 1784
rect 30115 1744 30124 1784
rect 30164 1744 34100 1784
rect 34156 1744 34444 1784
rect 34484 1744 34493 1784
rect 34627 1744 34636 1784
rect 34676 1744 40820 1784
rect 42403 1744 42412 1784
rect 42452 1744 43892 1784
rect 43987 1744 43996 1784
rect 44036 1744 46196 1784
rect 29884 1700 29924 1744
rect 34156 1700 34196 1744
rect 22265 1660 22348 1700
rect 22388 1660 22396 1700
rect 22436 1660 22445 1700
rect 23059 1660 23068 1700
rect 23108 1660 23116 1700
rect 23156 1660 23239 1700
rect 23731 1660 23740 1700
rect 23780 1660 23884 1700
rect 23924 1660 23933 1700
rect 23980 1660 24748 1700
rect 24788 1660 24797 1700
rect 24844 1660 26036 1700
rect 26947 1660 26956 1700
rect 26996 1660 29788 1700
rect 29828 1660 29837 1700
rect 29884 1660 34196 1700
rect 34339 1660 34348 1700
rect 34388 1660 38764 1700
rect 38804 1660 38813 1700
rect 40282 1660 40291 1700
rect 40331 1660 41068 1700
rect 41108 1660 41356 1700
rect 41396 1660 41644 1700
rect 41684 1660 42316 1700
rect 42356 1660 42365 1700
rect 43219 1660 43228 1700
rect 43268 1660 43508 1700
rect 43603 1660 43612 1700
rect 43652 1660 43988 1700
rect 23980 1616 24020 1660
rect 24844 1616 24884 1660
rect 13324 1576 13460 1616
rect 19180 1576 19276 1616
rect 19316 1576 19325 1616
rect 19948 1576 21716 1616
rect 21763 1576 21772 1616
rect 21812 1576 24020 1616
rect 24067 1576 24076 1616
rect 24116 1576 24884 1616
rect 24931 1576 24940 1616
rect 24980 1576 32716 1616
rect 32756 1576 32765 1616
rect 33571 1576 33580 1616
rect 33620 1576 38668 1616
rect 38708 1576 38717 1616
rect 38947 1576 38956 1616
rect 38996 1576 42604 1616
rect 42644 1576 42653 1616
rect 8236 1532 8276 1576
rect 13420 1532 13460 1576
rect 19948 1532 19988 1576
rect 43468 1532 43508 1660
rect 43948 1532 43988 1660
rect 46156 1616 46196 1744
rect 46278 1616 46368 1636
rect 46156 1576 46368 1616
rect 46278 1556 46368 1576
rect 4919 1492 4928 1532
rect 4968 1492 5010 1532
rect 5050 1492 5092 1532
rect 5132 1492 5174 1532
rect 5214 1492 5256 1532
rect 5296 1492 5305 1532
rect 5731 1492 5740 1532
rect 5780 1492 6988 1532
rect 7028 1492 7037 1532
rect 8236 1492 13324 1532
rect 13364 1492 13373 1532
rect 13420 1492 19988 1532
rect 20039 1492 20048 1532
rect 20088 1492 20130 1532
rect 20170 1492 20212 1532
rect 20252 1492 20294 1532
rect 20334 1492 20376 1532
rect 20416 1492 20425 1532
rect 20515 1492 20524 1532
rect 20564 1492 23308 1532
rect 23348 1492 23357 1532
rect 23491 1492 23500 1532
rect 23540 1492 27628 1532
rect 27668 1492 27677 1532
rect 27811 1492 27820 1532
rect 27860 1492 30124 1532
rect 30164 1492 30173 1532
rect 32419 1492 32428 1532
rect 32468 1492 33236 1532
rect 35159 1492 35168 1532
rect 35208 1492 35250 1532
rect 35290 1492 35332 1532
rect 35372 1492 35414 1532
rect 35454 1492 35496 1532
rect 35536 1492 35545 1532
rect 38860 1492 42700 1532
rect 42740 1492 42749 1532
rect 43468 1492 43892 1532
rect 43948 1492 45004 1532
rect 45044 1492 45053 1532
rect 33196 1448 33236 1492
rect 7171 1408 7180 1448
rect 7220 1408 33140 1448
rect 33196 1408 34828 1448
rect 34868 1408 34877 1448
rect 33100 1364 33140 1408
rect 38860 1364 38900 1492
rect 43852 1448 43892 1492
rect 43852 1408 44812 1448
rect 44852 1408 44861 1448
rect 2764 1324 31372 1364
rect 31412 1324 31421 1364
rect 33100 1324 38900 1364
rect 0 1280 90 1300
rect 46278 1280 46368 1300
rect 0 1240 1228 1280
rect 1268 1240 1277 1280
rect 44611 1240 44620 1280
rect 44660 1240 46368 1280
rect 0 1220 90 1240
rect 46278 1220 46368 1240
rect 0 944 90 964
rect 46278 944 46368 964
rect 0 904 1324 944
rect 1364 904 1373 944
rect 44803 904 44812 944
rect 44852 904 46368 944
rect 0 884 90 904
rect 46278 884 46368 904
rect 0 608 90 628
rect 46278 608 46368 628
rect 0 568 1420 608
rect 1460 568 1469 608
rect 44995 568 45004 608
rect 45044 568 46368 608
rect 0 548 90 568
rect 46278 548 46368 568
rect 14851 148 14860 188
rect 14900 148 29260 188
rect 29300 148 29309 188
rect 27715 64 27724 104
rect 27764 64 38860 104
rect 38900 64 38909 104
<< via2 >>
rect 19948 11068 19988 11108
rect 21196 11068 21236 11108
rect 1324 10984 1364 11024
rect 44716 10984 44756 11024
rect 18412 10900 18452 10940
rect 21004 10900 21044 10940
rect 28684 10732 28724 10772
rect 32332 10732 32372 10772
rect 1132 10648 1172 10688
rect 44236 10648 44276 10688
rect 1420 10312 1460 10352
rect 34444 10312 34484 10352
rect 39148 10312 39188 10352
rect 43276 10312 43316 10352
rect 30604 10228 30644 10268
rect 34924 10228 34964 10268
rect 17644 10144 17684 10184
rect 18220 10144 18260 10184
rect 23404 10144 23444 10184
rect 3436 10060 3476 10100
rect 15820 10060 15860 10100
rect 16300 10060 16340 10100
rect 18604 10060 18644 10100
rect 21004 10060 21044 10100
rect 21484 10060 21524 10100
rect 21676 10060 21716 10100
rect 22732 10060 22772 10100
rect 24652 10060 24692 10100
rect 25804 10060 25844 10100
rect 29548 10060 29588 10100
rect 31756 10060 31796 10100
rect 36460 10060 36500 10100
rect 36652 10060 36692 10100
rect 41452 10060 41492 10100
rect 2284 9976 2324 10016
rect 12652 9976 12692 10016
rect 12844 9976 12884 10016
rect 13420 9976 13460 10016
rect 23212 9976 23252 10016
rect 33868 9976 33908 10016
rect 37900 9976 37940 10016
rect 38668 9976 38708 10016
rect 42220 9976 42260 10016
rect 44428 9976 44468 10016
rect 1324 9892 1364 9932
rect 8236 9892 8276 9932
rect 11788 9892 11828 9932
rect 12076 9892 12116 9932
rect 15052 9892 15092 9932
rect 21292 9892 21332 9932
rect 29644 9892 29684 9932
rect 31468 9892 31508 9932
rect 33772 9892 33812 9932
rect 38188 9892 38228 9932
rect 41068 9892 41108 9932
rect 41548 9892 41588 9932
rect 1420 9556 1460 9596
rect 1228 9472 1268 9512
rect 3688 9808 3728 9848
rect 3770 9808 3810 9848
rect 3852 9808 3892 9848
rect 3934 9808 3974 9848
rect 4016 9808 4056 9848
rect 10924 9808 10964 9848
rect 13324 9808 13364 9848
rect 3436 9640 3476 9680
rect 15820 9808 15860 9848
rect 18220 9808 18260 9848
rect 18808 9808 18848 9848
rect 18890 9808 18930 9848
rect 18972 9808 19012 9848
rect 19054 9808 19094 9848
rect 19136 9808 19176 9848
rect 19276 9808 19316 9848
rect 20044 9808 20084 9848
rect 23116 9808 23156 9848
rect 28588 9808 28628 9848
rect 33388 9808 33428 9848
rect 33928 9808 33968 9848
rect 34010 9808 34050 9848
rect 34092 9808 34132 9848
rect 34174 9808 34214 9848
rect 34256 9808 34296 9848
rect 39052 9808 39092 9848
rect 44140 9808 44180 9848
rect 6220 9724 6260 9764
rect 9964 9724 10004 9764
rect 17548 9724 17588 9764
rect 19372 9724 19412 9764
rect 8236 9640 8276 9680
rect 10252 9640 10292 9680
rect 12076 9640 12116 9680
rect 12844 9640 12884 9680
rect 15436 9640 15476 9680
rect 20620 9640 20660 9680
rect 21580 9640 21620 9680
rect 22060 9640 22100 9680
rect 8140 9556 8180 9596
rect 10060 9556 10100 9596
rect 18124 9556 18164 9596
rect 19948 9556 19988 9596
rect 20716 9556 20756 9596
rect 5740 9472 5780 9512
rect 7948 9472 7988 9512
rect 8812 9472 8852 9512
rect 9292 9472 9332 9512
rect 11308 9472 11348 9512
rect 11884 9472 11924 9512
rect 12268 9472 12308 9512
rect 13420 9472 13460 9512
rect 14764 9472 14804 9512
rect 15436 9472 15476 9512
rect 15820 9472 15860 9512
rect 16204 9472 16244 9512
rect 5836 9388 5876 9428
rect 2860 9220 2900 9260
rect 4204 9220 4244 9260
rect 9004 9388 9044 9428
rect 10252 9388 10292 9428
rect 12652 9388 12692 9428
rect 14284 9388 14324 9428
rect 15148 9388 15188 9428
rect 16108 9388 16148 9428
rect 8620 9304 8660 9344
rect 9484 9304 9524 9344
rect 9964 9304 10004 9344
rect 10348 9304 10388 9344
rect 10636 9304 10676 9344
rect 21676 9556 21716 9596
rect 21868 9556 21908 9596
rect 23308 9724 23348 9764
rect 27052 9724 27092 9764
rect 32140 9724 32180 9764
rect 23500 9640 23540 9680
rect 24748 9640 24788 9680
rect 25132 9640 25172 9680
rect 29068 9640 29108 9680
rect 33484 9640 33524 9680
rect 34444 9640 34484 9680
rect 37228 9640 37268 9680
rect 38764 9640 38804 9680
rect 39148 9640 39188 9680
rect 43276 9640 43316 9680
rect 44428 9640 44468 9680
rect 23692 9556 23732 9596
rect 24076 9556 24116 9596
rect 24844 9556 24884 9596
rect 30700 9556 30740 9596
rect 31468 9556 31508 9596
rect 31660 9556 31700 9596
rect 33772 9556 33812 9596
rect 35596 9556 35636 9596
rect 35980 9556 36020 9596
rect 36172 9556 36212 9596
rect 36460 9556 36500 9596
rect 39340 9556 39380 9596
rect 17548 9472 17588 9512
rect 20140 9472 20180 9512
rect 24268 9472 24308 9512
rect 25228 9472 25268 9512
rect 25804 9472 25844 9512
rect 28300 9472 28340 9512
rect 28684 9472 28724 9512
rect 28876 9472 28916 9512
rect 29452 9472 29492 9512
rect 29836 9472 29876 9512
rect 32332 9472 32372 9512
rect 32716 9472 32756 9512
rect 33868 9472 33908 9512
rect 34540 9472 34580 9512
rect 37228 9472 37268 9512
rect 37708 9472 37748 9512
rect 38668 9472 38708 9512
rect 45196 9640 45236 9680
rect 39052 9472 39092 9512
rect 42316 9472 42356 9512
rect 42604 9472 42644 9512
rect 17836 9388 17876 9428
rect 18796 9388 18836 9428
rect 19852 9388 19892 9428
rect 20908 9388 20948 9428
rect 21292 9388 21332 9428
rect 22924 9388 22964 9428
rect 23884 9388 23924 9428
rect 24556 9388 24596 9428
rect 24748 9388 24788 9428
rect 27052 9388 27092 9428
rect 27436 9388 27476 9428
rect 27628 9388 27668 9428
rect 30124 9388 30164 9428
rect 32428 9388 32468 9428
rect 32812 9388 32852 9428
rect 35980 9388 36020 9428
rect 37420 9388 37460 9428
rect 38188 9388 38228 9428
rect 39628 9388 39668 9428
rect 14188 9304 14228 9344
rect 19372 9304 19412 9344
rect 22444 9304 22484 9344
rect 24940 9304 24980 9344
rect 29068 9304 29108 9344
rect 29548 9304 29588 9344
rect 30220 9304 30260 9344
rect 8044 9220 8084 9260
rect 10444 9220 10484 9260
rect 13132 9220 13172 9260
rect 18124 9220 18164 9260
rect 18412 9220 18452 9260
rect 18604 9220 18644 9260
rect 19180 9220 19220 9260
rect 19756 9220 19796 9260
rect 20044 9220 20084 9260
rect 21292 9220 21332 9260
rect 22348 9220 22388 9260
rect 22636 9220 22676 9260
rect 23692 9220 23732 9260
rect 23884 9220 23924 9260
rect 9580 9136 9620 9176
rect 10636 9136 10676 9176
rect 13804 9136 13844 9176
rect 15148 9136 15188 9176
rect 18508 9136 18548 9176
rect 20620 9136 20660 9176
rect 35308 9304 35348 9344
rect 38764 9304 38804 9344
rect 41356 9388 41396 9428
rect 38956 9304 38996 9344
rect 42028 9304 42068 9344
rect 42412 9304 42452 9344
rect 45004 9304 45044 9344
rect 24460 9220 24500 9260
rect 25900 9220 25940 9260
rect 26092 9220 26132 9260
rect 26284 9220 26324 9260
rect 27340 9220 27380 9260
rect 27820 9220 27860 9260
rect 28780 9220 28820 9260
rect 30316 9220 30356 9260
rect 30604 9220 30644 9260
rect 31276 9220 31316 9260
rect 32044 9220 32084 9260
rect 34156 9220 34196 9260
rect 34828 9220 34868 9260
rect 35884 9220 35924 9260
rect 37516 9220 37556 9260
rect 37804 9220 37844 9260
rect 38188 9220 38228 9260
rect 40204 9220 40235 9260
rect 40235 9220 40244 9260
rect 41740 9220 41771 9260
rect 41771 9220 41780 9260
rect 43084 9220 43124 9260
rect 44332 9220 44372 9260
rect 21580 9136 21620 9176
rect 21868 9136 21908 9176
rect 34444 9136 34484 9176
rect 36940 9136 36980 9176
rect 40492 9136 40532 9176
rect 42892 9136 42932 9176
rect 4108 9052 4148 9092
rect 4928 9052 4968 9092
rect 5010 9052 5050 9092
rect 5092 9052 5132 9092
rect 5174 9052 5214 9092
rect 5256 9052 5296 9092
rect 18892 9052 18932 9092
rect 19564 9052 19604 9092
rect 20048 9052 20088 9092
rect 20130 9052 20170 9092
rect 20212 9052 20252 9092
rect 20294 9052 20334 9092
rect 20376 9052 20416 9092
rect 28396 9052 28436 9092
rect 33196 9052 33236 9092
rect 34828 9052 34868 9092
rect 35168 9052 35208 9092
rect 35250 9052 35290 9092
rect 35332 9052 35372 9092
rect 35414 9052 35454 9092
rect 35496 9052 35536 9092
rect 37996 9052 38036 9092
rect 1228 8968 1268 9008
rect 12844 8968 12884 9008
rect 15436 8968 15476 9008
rect 22444 8968 22484 9008
rect 24172 8968 24212 9008
rect 26188 8968 26228 9008
rect 28108 8968 28148 9008
rect 28588 8968 28628 9008
rect 33004 8968 33044 9008
rect 8044 8884 8084 8924
rect 9004 8884 9044 8924
rect 10732 8884 10772 8924
rect 13804 8884 13844 8924
rect 16300 8884 16340 8924
rect 18796 8884 18836 8924
rect 20332 8884 20372 8924
rect 1132 8800 1172 8840
rect 4108 8800 4148 8840
rect 8524 8800 8564 8840
rect 10252 8800 10292 8840
rect 15148 8800 15188 8840
rect 2284 8716 2324 8756
rect 3532 8716 3572 8756
rect 5644 8747 5684 8756
rect 5644 8716 5684 8747
rect 6796 8716 6836 8756
rect 9196 8716 9236 8756
rect 9484 8716 9524 8756
rect 10156 8716 10196 8756
rect 16588 8800 16628 8840
rect 18028 8800 18068 8840
rect 19180 8800 19220 8840
rect 11500 8716 11540 8756
rect 11980 8716 12020 8756
rect 12940 8716 12980 8756
rect 14188 8716 14228 8756
rect 15340 8747 15380 8756
rect 15340 8716 15380 8747
rect 15820 8716 15860 8756
rect 16108 8716 16148 8756
rect 18604 8716 18644 8756
rect 18796 8716 18836 8756
rect 18988 8716 19028 8756
rect 39244 9052 39284 9092
rect 40300 9052 40340 9092
rect 40780 8968 40820 9008
rect 23212 8884 23252 8924
rect 24844 8884 24884 8924
rect 26476 8884 26516 8924
rect 34636 8884 34676 8924
rect 35692 8884 35732 8924
rect 35980 8884 36020 8924
rect 36172 8884 36212 8924
rect 41740 8884 41771 8924
rect 41771 8884 41780 8924
rect 44236 8884 44276 8924
rect 45196 8884 45236 8924
rect 22060 8800 22100 8840
rect 27244 8800 27284 8840
rect 28396 8800 28436 8840
rect 30892 8800 30932 8840
rect 33484 8800 33524 8840
rect 33868 8800 33908 8840
rect 19756 8716 19796 8756
rect 20332 8716 20372 8756
rect 21100 8716 21140 8756
rect 1132 8632 1172 8672
rect 8524 8632 8564 8672
rect 9580 8632 9620 8672
rect 11884 8632 11924 8672
rect 12268 8632 12308 8672
rect 13132 8632 13172 8672
rect 13804 8632 13844 8672
rect 14764 8632 14804 8672
rect 15148 8632 15188 8672
rect 15916 8632 15956 8672
rect 18316 8632 18356 8672
rect 20236 8632 20276 8672
rect 8620 8548 8660 8588
rect 13228 8548 13268 8588
rect 13900 8464 13940 8504
rect 14380 8464 14420 8504
rect 15820 8464 15860 8504
rect 17260 8464 17300 8504
rect 19276 8464 19316 8504
rect 22348 8716 22388 8756
rect 22828 8716 22868 8756
rect 23788 8716 23828 8756
rect 20524 8632 20564 8672
rect 20908 8632 20948 8672
rect 21196 8632 21236 8672
rect 21676 8632 21716 8672
rect 22060 8632 22100 8672
rect 24652 8716 24692 8756
rect 25612 8747 25652 8756
rect 25612 8716 25652 8747
rect 26092 8747 26132 8756
rect 26092 8716 26132 8747
rect 24076 8548 24116 8588
rect 24364 8632 24404 8672
rect 25132 8632 25172 8672
rect 29356 8716 29396 8756
rect 30412 8716 30452 8756
rect 31468 8716 31508 8756
rect 32140 8716 32180 8756
rect 33292 8716 33332 8756
rect 33580 8716 33611 8756
rect 33611 8716 33620 8756
rect 34060 8800 34100 8840
rect 34540 8800 34580 8840
rect 34156 8716 34196 8756
rect 35980 8716 36020 8756
rect 37516 8716 37556 8756
rect 37900 8716 37940 8756
rect 38860 8716 38900 8756
rect 41260 8800 41300 8840
rect 39628 8716 39668 8756
rect 40012 8716 40052 8756
rect 27436 8632 27476 8672
rect 27820 8632 27860 8672
rect 28108 8632 28148 8672
rect 28684 8632 28724 8672
rect 29068 8632 29099 8672
rect 29099 8632 29108 8672
rect 30988 8632 31028 8672
rect 33196 8632 33236 8672
rect 33388 8632 33428 8672
rect 34924 8632 34964 8672
rect 35788 8632 35828 8672
rect 37804 8632 37844 8672
rect 38764 8632 38804 8672
rect 39148 8632 39188 8672
rect 40396 8632 40436 8672
rect 40780 8632 40820 8672
rect 43084 8632 43124 8672
rect 43468 8632 43508 8672
rect 24460 8548 24500 8588
rect 28972 8548 29012 8588
rect 29740 8548 29780 8588
rect 29932 8548 29972 8588
rect 33004 8548 33044 8588
rect 38860 8548 38900 8588
rect 41740 8548 41780 8588
rect 23788 8464 23828 8504
rect 24268 8464 24308 8504
rect 27532 8464 27572 8504
rect 28588 8464 28628 8504
rect 30220 8464 30260 8504
rect 35980 8464 36020 8504
rect 38380 8464 38420 8504
rect 41164 8464 41204 8504
rect 45772 8464 45812 8504
rect 11020 8380 11060 8420
rect 19948 8380 19988 8420
rect 20332 8380 20372 8420
rect 20620 8380 20660 8420
rect 22732 8380 22772 8420
rect 32908 8380 32948 8420
rect 34924 8380 34964 8420
rect 36268 8380 36308 8420
rect 3688 8296 3728 8336
rect 3770 8296 3810 8336
rect 3852 8296 3892 8336
rect 3934 8296 3974 8336
rect 4016 8296 4056 8336
rect 14572 8296 14612 8336
rect 18604 8296 18644 8336
rect 18808 8296 18848 8336
rect 18890 8296 18930 8336
rect 18972 8296 19012 8336
rect 19054 8296 19094 8336
rect 19136 8296 19176 8336
rect 28780 8296 28820 8336
rect 29932 8212 29972 8252
rect 32524 8296 32564 8336
rect 33928 8296 33968 8336
rect 34010 8296 34050 8336
rect 34092 8296 34132 8336
rect 34174 8296 34214 8336
rect 34256 8296 34296 8336
rect 35212 8296 35252 8336
rect 40204 8296 40244 8336
rect 30796 8212 30836 8252
rect 32716 8212 32756 8252
rect 34732 8212 34772 8252
rect 34924 8212 34964 8252
rect 10252 8128 10292 8168
rect 13612 8128 13652 8168
rect 17932 8128 17972 8168
rect 22444 8128 22484 8168
rect 25708 8128 25748 8168
rect 26092 8128 26132 8168
rect 28204 8128 28244 8168
rect 33292 8128 33332 8168
rect 1132 8044 1172 8084
rect 7180 8044 7220 8084
rect 9964 8044 10004 8084
rect 10636 8044 10676 8084
rect 11788 8044 11828 8084
rect 14092 8044 14132 8084
rect 17260 8044 17300 8084
rect 20524 8044 20564 8084
rect 21388 8044 21428 8084
rect 22156 8044 22196 8084
rect 26188 8044 26228 8084
rect 1228 7960 1268 8000
rect 4108 7960 4148 8000
rect 9484 7960 9524 8000
rect 10828 7960 10868 8000
rect 11116 7960 11156 8000
rect 11500 7960 11540 8000
rect 11980 7960 12020 8000
rect 13612 7960 13652 8000
rect 16300 7960 16340 8000
rect 17452 7960 17492 8000
rect 18796 7960 18836 8000
rect 19756 7960 19796 8000
rect 22252 7960 22292 8000
rect 23212 7960 23252 8000
rect 23404 7960 23444 8000
rect 5740 7876 5780 7916
rect 6796 7876 6836 7916
rect 26380 8044 26420 8084
rect 28108 8044 28148 8084
rect 35116 8212 35156 8252
rect 40396 8212 40436 8252
rect 35980 8128 36020 8168
rect 37420 8128 37460 8168
rect 30220 8044 30260 8084
rect 34732 8044 34772 8084
rect 37324 8044 37364 8084
rect 39148 8044 39188 8084
rect 32716 7960 32756 8000
rect 36364 7960 36404 8000
rect 36748 7960 36788 8000
rect 45004 8296 45044 8336
rect 44716 8128 44756 8168
rect 40684 7960 40724 8000
rect 41452 7960 41492 8000
rect 41740 7960 41780 8000
rect 44332 7960 44372 8000
rect 45772 7960 45812 8000
rect 10636 7907 10676 7916
rect 10636 7876 10676 7907
rect 12652 7876 12692 7916
rect 13036 7876 13076 7916
rect 14380 7876 14420 7916
rect 15340 7876 15380 7916
rect 15820 7876 15860 7916
rect 17068 7876 17108 7916
rect 18028 7876 18068 7916
rect 19948 7876 19988 7916
rect 20140 7876 20180 7916
rect 20428 7876 20468 7916
rect 21772 7876 21812 7916
rect 23788 7876 23828 7916
rect 25804 7876 25844 7916
rect 28588 7876 28628 7916
rect 29356 7876 29396 7916
rect 29740 7876 29780 7916
rect 31372 7876 31412 7916
rect 32140 7876 32180 7916
rect 32812 7876 32852 7916
rect 34156 7876 34196 7916
rect 34924 7876 34964 7916
rect 38668 7876 38708 7916
rect 39820 7876 39860 7916
rect 41260 7876 41300 7916
rect 10348 7792 10388 7832
rect 12172 7792 12212 7832
rect 14572 7792 14612 7832
rect 18220 7792 18260 7832
rect 19468 7792 19508 7832
rect 21676 7792 21716 7832
rect 22252 7792 22292 7832
rect 22828 7792 22868 7832
rect 24172 7792 24212 7832
rect 25996 7792 26036 7832
rect 27340 7792 27380 7832
rect 1708 7708 1748 7748
rect 2860 7708 2900 7748
rect 5932 7708 5972 7748
rect 4928 7540 4968 7580
rect 5010 7540 5050 7580
rect 5092 7540 5132 7580
rect 5174 7540 5214 7580
rect 5256 7540 5296 7580
rect 1228 7288 1268 7328
rect 31660 7792 31700 7832
rect 33292 7792 33332 7832
rect 35788 7792 35828 7832
rect 35980 7792 36020 7832
rect 37708 7792 37748 7832
rect 15052 7708 15092 7748
rect 15340 7708 15380 7748
rect 19852 7708 19892 7748
rect 21100 7708 21140 7748
rect 22444 7708 22484 7748
rect 24652 7708 24692 7748
rect 28396 7708 28436 7748
rect 29932 7708 29972 7748
rect 33580 7708 33620 7748
rect 11500 7624 11540 7664
rect 12172 7624 12212 7664
rect 19756 7624 19796 7664
rect 34252 7624 34292 7664
rect 9100 7540 9140 7580
rect 14764 7540 14804 7580
rect 15532 7540 15572 7580
rect 20048 7540 20088 7580
rect 20130 7540 20170 7580
rect 20212 7540 20252 7580
rect 20294 7540 20334 7580
rect 20376 7540 20416 7580
rect 27628 7540 27668 7580
rect 28396 7540 28436 7580
rect 29068 7540 29108 7580
rect 34156 7540 34196 7580
rect 15052 7456 15092 7496
rect 9676 7372 9716 7412
rect 9772 7288 9812 7328
rect 10732 7288 10772 7328
rect 18796 7372 18836 7412
rect 22444 7372 22484 7412
rect 29356 7372 29396 7412
rect 33100 7372 33140 7412
rect 33580 7372 33620 7412
rect 33964 7372 34004 7412
rect 10444 7204 10484 7244
rect 11020 7204 11060 7244
rect 76 7120 116 7160
rect 3532 7120 3572 7160
rect 6316 7120 6356 7160
rect 7180 7120 7220 7160
rect 8140 7120 8180 7160
rect 8908 7120 8948 7160
rect 10732 7120 10772 7160
rect 11692 7120 11732 7160
rect 13900 7288 13940 7328
rect 18892 7288 18932 7328
rect 19468 7288 19508 7328
rect 21964 7288 22004 7328
rect 23020 7288 23060 7328
rect 23596 7288 23636 7328
rect 25612 7288 25652 7328
rect 27724 7288 27764 7328
rect 31084 7288 31124 7328
rect 31852 7288 31892 7328
rect 34348 7288 34388 7328
rect 12940 7204 12980 7244
rect 14476 7204 14516 7244
rect 11980 7120 12020 7160
rect 12844 7120 12884 7160
rect 13036 7120 13076 7160
rect 13900 7120 13940 7160
rect 14380 7120 14420 7160
rect 14572 7120 14612 7160
rect 13516 7036 13556 7076
rect 14092 7036 14132 7076
rect 14860 7036 14900 7076
rect 76 6952 116 6992
rect 4300 6952 4340 6992
rect 10540 6952 10580 6992
rect 10732 6952 10772 6992
rect 11116 6952 11156 6992
rect 11788 6952 11828 6992
rect 12940 6952 12980 6992
rect 13708 6952 13748 6992
rect 14380 6952 14420 6992
rect 14764 6952 14804 6992
rect 9964 6868 10004 6908
rect 12748 6868 12788 6908
rect 3688 6784 3728 6824
rect 3770 6784 3810 6824
rect 3852 6784 3892 6824
rect 3934 6784 3974 6824
rect 4016 6784 4056 6824
rect 11212 6784 11252 6824
rect 13324 6784 13364 6824
rect 12748 6700 12788 6740
rect 76 6448 116 6488
rect 16492 7204 16532 7244
rect 17068 7204 17108 7244
rect 17452 7204 17492 7244
rect 15532 7120 15572 7160
rect 16108 7120 16148 7160
rect 18412 7204 18452 7244
rect 20524 7204 20564 7244
rect 21292 7204 21332 7244
rect 21580 7204 21611 7244
rect 21611 7204 21620 7244
rect 22156 7204 22196 7244
rect 16300 7120 16340 7160
rect 16684 7120 16724 7160
rect 18892 7120 18932 7160
rect 36076 7708 36116 7748
rect 38956 7708 38996 7748
rect 39244 7708 39284 7748
rect 40780 7708 40820 7748
rect 45772 7708 45812 7748
rect 35168 7540 35208 7580
rect 35250 7540 35290 7580
rect 35332 7540 35372 7580
rect 35414 7540 35454 7580
rect 35496 7540 35536 7580
rect 36748 7540 36788 7580
rect 40972 7540 41012 7580
rect 36364 7372 36404 7412
rect 41452 7372 41492 7412
rect 41836 7372 41867 7412
rect 41867 7372 41876 7412
rect 34828 7288 34868 7328
rect 36076 7288 36116 7328
rect 37900 7288 37940 7328
rect 39916 7288 39956 7328
rect 45772 7288 45812 7328
rect 27148 7204 27188 7244
rect 29068 7204 29108 7244
rect 29548 7204 29588 7244
rect 31660 7204 31700 7244
rect 32140 7204 32180 7244
rect 33676 7204 33716 7244
rect 19660 7120 19700 7160
rect 19948 7120 19988 7160
rect 20812 7120 20852 7160
rect 21964 7120 22004 7160
rect 22828 7120 22868 7160
rect 23788 7120 23828 7160
rect 25036 7120 25076 7160
rect 25324 7120 25364 7160
rect 26956 7120 26996 7160
rect 27532 7120 27572 7160
rect 29644 7120 29684 7160
rect 30412 7120 30452 7160
rect 32716 7120 32756 7160
rect 34060 7120 34100 7160
rect 34540 7120 34580 7160
rect 35980 7235 36020 7244
rect 35980 7204 36020 7235
rect 39436 7204 39476 7244
rect 40684 7235 40724 7244
rect 40684 7204 40724 7235
rect 34732 7120 34772 7160
rect 36940 7120 36980 7160
rect 37708 7120 37748 7160
rect 43276 7120 43316 7160
rect 43852 7120 43892 7160
rect 44908 7120 44948 7160
rect 17164 7036 17204 7076
rect 19852 7036 19892 7076
rect 20716 7036 20756 7076
rect 23212 7036 23252 7076
rect 25132 7036 25172 7076
rect 25420 7036 25460 7076
rect 27340 7036 27380 7076
rect 29740 7036 29780 7076
rect 30028 7036 30068 7076
rect 32620 7036 32660 7076
rect 32812 7036 32852 7076
rect 33868 7036 33908 7076
rect 35596 7036 35636 7076
rect 38092 7036 38132 7076
rect 46156 7036 46196 7076
rect 16012 6952 16052 6992
rect 16780 6952 16820 6992
rect 17068 6952 17108 6992
rect 19180 6952 19220 6992
rect 20140 6952 20180 6992
rect 20908 6952 20948 6992
rect 21580 6952 21620 6992
rect 23404 6952 23444 6992
rect 23692 6952 23732 6992
rect 24364 6952 24404 6992
rect 25900 6952 25940 6992
rect 27052 6952 27092 6992
rect 29644 6952 29684 6992
rect 31852 6952 31892 6992
rect 32236 6952 32276 6992
rect 33004 6952 33044 6992
rect 21004 6868 21044 6908
rect 26572 6868 26612 6908
rect 26764 6868 26804 6908
rect 30028 6868 30068 6908
rect 32716 6868 32756 6908
rect 33580 6868 33620 6908
rect 34636 6868 34676 6908
rect 36844 6952 36884 6992
rect 37324 6952 37364 6992
rect 41260 6952 41300 6992
rect 16396 6784 16436 6824
rect 18808 6784 18848 6824
rect 18890 6784 18930 6824
rect 18972 6784 19012 6824
rect 19054 6784 19094 6824
rect 19136 6784 19176 6824
rect 26668 6784 26708 6824
rect 29740 6784 29780 6824
rect 33928 6784 33968 6824
rect 34010 6784 34050 6824
rect 34092 6784 34132 6824
rect 34174 6784 34214 6824
rect 34256 6784 34296 6824
rect 34444 6784 34484 6824
rect 13516 6700 13556 6740
rect 14380 6700 14420 6740
rect 14668 6700 14708 6740
rect 15916 6700 15956 6740
rect 16492 6700 16532 6740
rect 22636 6700 22676 6740
rect 29836 6700 29876 6740
rect 32716 6700 32756 6740
rect 41932 6952 41972 6992
rect 11116 6616 11156 6656
rect 12556 6616 12596 6656
rect 15244 6616 15284 6656
rect 17356 6616 17396 6656
rect 17740 6616 17780 6656
rect 18700 6616 18740 6656
rect 20620 6616 20660 6656
rect 22924 6616 22964 6656
rect 23212 6616 23252 6656
rect 26668 6616 26708 6656
rect 27052 6616 27092 6656
rect 32812 6616 32852 6656
rect 33964 6616 34004 6656
rect 34828 6616 34868 6656
rect 35980 6616 36020 6656
rect 37036 6616 37076 6656
rect 42028 6616 42068 6656
rect 46252 6616 46292 6656
rect 5740 6532 5780 6572
rect 10156 6532 10196 6572
rect 12172 6532 12212 6572
rect 5932 6448 5972 6488
rect 6220 6448 6260 6488
rect 3532 6364 3572 6404
rect 6412 6364 6452 6404
rect 6796 6364 6836 6404
rect 9676 6448 9716 6488
rect 10252 6448 10292 6488
rect 11020 6448 11060 6488
rect 12268 6448 12308 6488
rect 12556 6448 12596 6488
rect 8812 6364 8852 6404
rect 9388 6364 9428 6404
rect 10156 6364 10196 6404
rect 76 6280 116 6320
rect 5644 6196 5684 6236
rect 10636 6364 10676 6404
rect 11500 6364 11540 6404
rect 12652 6364 12692 6404
rect 9196 6280 9236 6320
rect 10252 6280 10292 6320
rect 10444 6280 10484 6320
rect 23020 6532 23060 6572
rect 24268 6532 24308 6572
rect 28108 6532 28148 6572
rect 28876 6532 28916 6572
rect 32620 6532 32660 6572
rect 34348 6532 34388 6572
rect 35596 6532 35636 6572
rect 35788 6532 35828 6572
rect 37420 6532 37460 6572
rect 42412 6532 42452 6572
rect 14380 6448 14420 6488
rect 17644 6448 17684 6488
rect 18028 6448 18068 6488
rect 19948 6448 19988 6488
rect 21772 6448 21812 6488
rect 22156 6448 22196 6488
rect 24556 6448 24596 6488
rect 25324 6448 25364 6488
rect 27148 6448 27188 6488
rect 27916 6448 27956 6488
rect 28780 6448 28820 6488
rect 31468 6448 31508 6488
rect 14668 6364 14708 6404
rect 15052 6364 15092 6404
rect 16012 6364 16052 6404
rect 17260 6364 17300 6404
rect 18124 6364 18164 6404
rect 19180 6364 19220 6404
rect 20716 6364 20756 6404
rect 22060 6364 22100 6404
rect 22252 6364 22292 6404
rect 22540 6364 22580 6404
rect 23596 6364 23636 6404
rect 25900 6364 25940 6404
rect 28972 6364 29012 6404
rect 29548 6364 29588 6404
rect 31372 6364 31412 6404
rect 32044 6364 32084 6404
rect 32236 6364 32276 6404
rect 34828 6364 34868 6404
rect 35980 6364 36020 6404
rect 36748 6364 36788 6404
rect 38188 6364 38228 6404
rect 38956 6364 38996 6404
rect 13900 6280 13940 6320
rect 16108 6280 16148 6320
rect 19468 6280 19508 6320
rect 7468 6196 7508 6236
rect 11116 6196 11156 6236
rect 12268 6196 12308 6236
rect 27340 6280 27380 6320
rect 28684 6280 28724 6320
rect 33004 6280 33044 6320
rect 13996 6196 14036 6236
rect 20524 6196 20564 6236
rect 22252 6196 22292 6236
rect 25900 6196 25940 6236
rect 28300 6196 28340 6236
rect 33676 6280 33716 6320
rect 34060 6280 34100 6320
rect 34636 6280 34676 6320
rect 35788 6280 35828 6320
rect 37900 6280 37940 6320
rect 39628 6364 39668 6404
rect 40108 6364 40148 6404
rect 40588 6364 40596 6404
rect 40596 6364 40628 6404
rect 41260 6364 41300 6404
rect 42124 6364 42164 6404
rect 42412 6364 42443 6404
rect 42443 6364 42452 6404
rect 40876 6280 40916 6320
rect 40396 6196 40436 6236
rect 41740 6196 41780 6236
rect 43852 6196 43883 6236
rect 43883 6196 43892 6236
rect 9196 6112 9236 6152
rect 13324 6112 13364 6152
rect 15820 6112 15860 6152
rect 16012 6112 16052 6152
rect 19180 6112 19220 6152
rect 19660 6112 19700 6152
rect 23212 6112 23252 6152
rect 23596 6112 23636 6152
rect 31756 6112 31796 6152
rect 39628 6112 39668 6152
rect 42412 6112 42452 6152
rect 44428 6448 44468 6488
rect 4928 6028 4968 6068
rect 5010 6028 5050 6068
rect 5092 6028 5132 6068
rect 5174 6028 5214 6068
rect 5256 6028 5296 6068
rect 18412 6028 18452 6068
rect 20048 6028 20088 6068
rect 20130 6028 20170 6068
rect 20212 6028 20252 6068
rect 20294 6028 20334 6068
rect 20376 6028 20416 6068
rect 26764 6028 26804 6068
rect 35168 6028 35208 6068
rect 35250 6028 35290 6068
rect 35332 6028 35372 6068
rect 35414 6028 35454 6068
rect 35496 6028 35536 6068
rect 36364 6028 36404 6068
rect 12748 5944 12788 5984
rect 13900 5944 13940 5984
rect 20812 5944 20852 5984
rect 28876 5944 28916 5984
rect 46252 6112 46292 6152
rect 31564 5944 31604 5984
rect 41932 5944 41972 5984
rect 46252 5944 46292 5984
rect 12940 5860 12980 5900
rect 13996 5860 14036 5900
rect 22924 5860 22964 5900
rect 23116 5860 23156 5900
rect 29644 5860 29684 5900
rect 42124 5860 42164 5900
rect 5932 5776 5972 5816
rect 9676 5776 9716 5816
rect 10348 5776 10388 5816
rect 13036 5776 13076 5816
rect 16492 5776 16532 5816
rect 19276 5776 19316 5816
rect 21580 5776 21620 5816
rect 22732 5776 22772 5816
rect 39628 5776 39668 5816
rect 40780 5776 40820 5816
rect 3532 5692 3572 5732
rect 4780 5723 4820 5732
rect 4780 5692 4784 5723
rect 4784 5692 4820 5723
rect 5644 5692 5684 5732
rect 6220 5692 6260 5732
rect 9004 5692 9044 5732
rect 11020 5692 11051 5732
rect 11051 5692 11060 5732
rect 1996 5608 2036 5648
rect 9772 5608 9812 5648
rect 10060 5608 10100 5648
rect 4684 5524 4724 5564
rect 5836 5524 5876 5564
rect 6316 5524 6356 5564
rect 5452 5440 5492 5480
rect 8332 5440 8372 5480
rect 9004 5440 9044 5480
rect 10540 5440 10580 5480
rect 6028 5356 6068 5396
rect 3688 5272 3728 5312
rect 3770 5272 3810 5312
rect 3852 5272 3892 5312
rect 3934 5272 3974 5312
rect 4016 5272 4056 5312
rect 14668 5692 14708 5732
rect 15916 5723 15956 5732
rect 15916 5692 15956 5723
rect 11788 5608 11828 5648
rect 12364 5608 12404 5648
rect 13132 5608 13172 5648
rect 20044 5692 20084 5732
rect 20716 5692 20756 5732
rect 21004 5692 21044 5732
rect 21388 5692 21428 5732
rect 22540 5692 22580 5732
rect 23404 5692 23444 5732
rect 24268 5692 24308 5732
rect 25996 5692 26036 5732
rect 27532 5692 27572 5732
rect 14188 5608 14228 5648
rect 19948 5608 19988 5648
rect 22060 5608 22100 5648
rect 22444 5608 22484 5648
rect 23020 5608 23060 5648
rect 23692 5608 23732 5648
rect 25132 5608 25172 5648
rect 25708 5608 25739 5648
rect 25739 5608 25748 5648
rect 12748 5524 12788 5564
rect 12940 5524 12980 5564
rect 14668 5524 14708 5564
rect 15628 5524 15668 5564
rect 20524 5524 20564 5564
rect 21292 5524 21332 5564
rect 25612 5524 25652 5564
rect 12652 5440 12692 5480
rect 15148 5440 15188 5480
rect 15436 5440 15476 5480
rect 15916 5440 15956 5480
rect 17836 5440 17876 5480
rect 24556 5440 24596 5480
rect 22252 5356 22292 5396
rect 29260 5692 29300 5732
rect 26188 5608 26228 5648
rect 28876 5608 28916 5648
rect 29452 5608 29492 5648
rect 33676 5692 33716 5732
rect 33964 5692 34004 5732
rect 34636 5692 34676 5732
rect 34828 5692 34868 5732
rect 32908 5608 32948 5648
rect 33196 5608 33236 5648
rect 33868 5608 33872 5648
rect 33872 5608 33908 5648
rect 34060 5608 34100 5648
rect 31756 5524 31796 5564
rect 33004 5524 33044 5564
rect 33484 5524 33524 5564
rect 28972 5440 29012 5480
rect 30220 5440 30260 5480
rect 32812 5440 32852 5480
rect 33868 5440 33908 5480
rect 34444 5440 34484 5480
rect 38956 5692 38996 5732
rect 39436 5692 39476 5732
rect 39820 5723 39860 5732
rect 39820 5692 39860 5723
rect 40300 5692 40340 5732
rect 40684 5692 40724 5732
rect 35020 5608 35060 5648
rect 35596 5608 35636 5648
rect 36460 5608 36500 5648
rect 37420 5608 37460 5648
rect 37996 5608 38036 5648
rect 38860 5608 38900 5648
rect 42988 5608 43028 5648
rect 43852 5608 43892 5648
rect 36172 5524 36212 5564
rect 42412 5524 42452 5564
rect 35116 5440 35156 5480
rect 30124 5356 30164 5396
rect 31180 5356 31220 5396
rect 32716 5356 32756 5396
rect 35980 5440 36020 5480
rect 38572 5440 38612 5480
rect 40588 5440 40628 5480
rect 42508 5356 42548 5396
rect 12652 5272 12692 5312
rect 15532 5272 15572 5312
rect 17356 5272 17396 5312
rect 18124 5272 18164 5312
rect 18808 5272 18848 5312
rect 18890 5272 18930 5312
rect 18972 5272 19012 5312
rect 19054 5272 19094 5312
rect 19136 5272 19176 5312
rect 19276 5272 19316 5312
rect 22540 5272 22580 5312
rect 27532 5272 27572 5312
rect 31948 5272 31988 5312
rect 32812 5272 32852 5312
rect 33928 5272 33968 5312
rect 34010 5272 34050 5312
rect 34092 5272 34132 5312
rect 34174 5272 34214 5312
rect 34256 5272 34296 5312
rect 41644 5272 41684 5312
rect 14188 5188 14228 5228
rect 14764 5188 14804 5228
rect 29260 5188 29300 5228
rect 31660 5188 31700 5228
rect 8524 5104 8564 5144
rect 8716 5104 8756 5144
rect 11404 5104 11444 5144
rect 46252 5440 46292 5480
rect 46252 5272 46292 5312
rect 35116 5188 35156 5228
rect 12748 5104 12788 5144
rect 23596 5104 23636 5144
rect 28972 5104 29012 5144
rect 31372 5104 31412 5144
rect 33196 5104 33236 5144
rect 36076 5104 36116 5144
rect 36556 5104 36596 5144
rect 1996 5020 2036 5060
rect 6412 5020 6452 5060
rect 14188 5020 14228 5060
rect 1612 4936 1652 4976
rect 9196 4936 9236 4976
rect 9676 4936 9716 4976
rect 11692 4936 11732 4976
rect 11884 4936 11924 4976
rect 14668 5020 14708 5060
rect 17356 5020 17396 5060
rect 18412 5020 18452 5060
rect 23980 5020 24020 5060
rect 12652 4936 12692 4976
rect 14764 4936 14804 4976
rect 5452 4852 5492 4892
rect 5740 4852 5771 4892
rect 5771 4852 5780 4892
rect 6316 4852 6356 4892
rect 6700 4852 6731 4892
rect 6731 4852 6740 4892
rect 7564 4852 7604 4892
rect 8620 4852 8660 4892
rect 9772 4852 9812 4892
rect 11212 4852 11252 4892
rect 11596 4852 11636 4892
rect 12460 4852 12500 4892
rect 13900 4852 13940 4892
rect 19948 4936 19988 4976
rect 23692 4936 23732 4976
rect 15532 4852 15572 4892
rect 16492 4852 16532 4892
rect 17260 4852 17300 4892
rect 20524 4852 20564 4892
rect 22444 4852 22484 4892
rect 22636 4852 22676 4892
rect 23788 4852 23828 4892
rect 24172 5020 24212 5060
rect 33100 5020 33140 5060
rect 34732 5020 34772 5060
rect 42028 5020 42068 5060
rect 43756 5020 43796 5060
rect 24268 4936 24308 4976
rect 25996 4936 26036 4976
rect 27052 4936 27092 4976
rect 28972 4936 29012 4976
rect 29740 4936 29780 4976
rect 32524 4936 32564 4976
rect 34348 4936 34388 4976
rect 24556 4852 24596 4892
rect 27148 4852 27188 4892
rect 28588 4852 28628 4892
rect 29164 4852 29204 4892
rect 32620 4852 32660 4892
rect 33292 4852 33332 4892
rect 33868 4852 33908 4892
rect 38956 4936 38996 4976
rect 40300 4936 40340 4976
rect 40588 4936 40628 4976
rect 34924 4852 34964 4892
rect 38572 4852 38612 4892
rect 39436 4852 39476 4892
rect 41260 4936 41300 4976
rect 44236 4852 44276 4892
rect 76 4768 116 4808
rect 4396 4768 4436 4808
rect 8524 4768 8564 4808
rect 9964 4768 10004 4808
rect 15820 4768 15860 4808
rect 18412 4768 18452 4808
rect 18700 4768 18740 4808
rect 21580 4768 21620 4808
rect 24268 4768 24308 4808
rect 27052 4768 27092 4808
rect 33196 4768 33236 4808
rect 33484 4768 33524 4808
rect 33676 4768 33716 4808
rect 37996 4768 38036 4808
rect 40876 4768 40916 4808
rect 6028 4684 6068 4724
rect 11020 4684 11060 4724
rect 12172 4684 12212 4724
rect 13324 4684 13364 4724
rect 13612 4684 13652 4724
rect 18220 4684 18260 4724
rect 24076 4684 24116 4724
rect 29068 4684 29108 4724
rect 29260 4684 29300 4724
rect 29452 4684 29492 4724
rect 30124 4684 30164 4724
rect 38764 4684 38804 4724
rect 41068 4684 41108 4724
rect 76 4600 116 4640
rect 42988 4684 43019 4724
rect 43019 4684 43028 4724
rect 43852 4684 43883 4724
rect 43883 4684 43892 4724
rect 8044 4600 8084 4640
rect 9100 4600 9140 4640
rect 9484 4600 9524 4640
rect 15244 4600 15284 4640
rect 15820 4600 15860 4640
rect 22924 4600 22964 4640
rect 31660 4600 31700 4640
rect 35692 4600 35732 4640
rect 4928 4516 4968 4556
rect 5010 4516 5050 4556
rect 5092 4516 5132 4556
rect 5174 4516 5214 4556
rect 5256 4516 5296 4556
rect 17260 4516 17300 4556
rect 20048 4516 20088 4556
rect 20130 4516 20170 4556
rect 20212 4516 20252 4556
rect 20294 4516 20334 4556
rect 20376 4516 20416 4556
rect 23980 4516 24020 4556
rect 28492 4516 28532 4556
rect 35168 4516 35208 4556
rect 35250 4516 35290 4556
rect 35332 4516 35372 4556
rect 35414 4516 35454 4556
rect 35496 4516 35536 4556
rect 38188 4516 38228 4556
rect 43756 4516 43796 4556
rect 8620 4432 8660 4472
rect 9964 4432 10004 4472
rect 10540 4432 10580 4472
rect 14476 4432 14516 4472
rect 15148 4432 15188 4472
rect 32908 4432 32948 4472
rect 39916 4432 39956 4472
rect 8332 4348 8372 4388
rect 13324 4348 13364 4388
rect 15820 4348 15860 4388
rect 21388 4348 21428 4388
rect 23788 4348 23828 4388
rect 24172 4348 24212 4388
rect 24364 4348 24404 4388
rect 32236 4348 32276 4388
rect 33292 4348 33332 4388
rect 40588 4348 40628 4388
rect 1612 4264 1652 4304
rect 7948 4264 7988 4304
rect 8908 4264 8948 4304
rect 9292 4264 9332 4304
rect 9676 4264 9716 4304
rect 11692 4264 11732 4304
rect 14668 4264 14708 4304
rect 15148 4264 15188 4304
rect 18412 4264 18452 4304
rect 20908 4264 20948 4304
rect 6028 4211 6068 4220
rect 6028 4180 6068 4211
rect 6892 4180 6932 4220
rect 8044 4180 8084 4220
rect 22348 4264 22388 4304
rect 23500 4264 23540 4304
rect 32620 4264 32660 4304
rect 33100 4264 33140 4304
rect 34924 4264 34964 4304
rect 38764 4264 38804 4304
rect 38956 4264 38996 4304
rect 39148 4264 39188 4304
rect 40300 4264 40340 4304
rect 43852 4264 43892 4304
rect 8620 4211 8660 4220
rect 8620 4180 8660 4211
rect 9484 4180 9524 4220
rect 10060 4180 10100 4220
rect 11980 4180 12020 4220
rect 13132 4180 13172 4220
rect 13708 4180 13748 4220
rect 15436 4180 15476 4220
rect 15628 4180 15668 4220
rect 17932 4180 17972 4220
rect 76 4096 116 4136
rect 4108 4096 4148 4136
rect 6412 4096 6452 4136
rect 7660 4096 7700 4136
rect 9004 4096 9044 4136
rect 11020 4096 11060 4136
rect 14188 4096 14228 4136
rect 15820 4096 15860 4136
rect 76 3928 116 3968
rect 18796 4180 18836 4220
rect 24940 4180 24980 4220
rect 25132 4180 25172 4220
rect 25324 4180 25364 4220
rect 27244 4180 27284 4220
rect 28876 4211 28916 4220
rect 28876 4180 28916 4211
rect 19948 4096 19988 4136
rect 20428 4096 20468 4136
rect 22060 4096 22100 4136
rect 22252 4096 22292 4136
rect 23500 4096 23540 4136
rect 23692 4096 23732 4136
rect 24556 4096 24596 4136
rect 28588 4096 28628 4136
rect 29164 4096 29204 4136
rect 31948 4180 31988 4220
rect 32812 4180 32852 4220
rect 33292 4180 33332 4220
rect 33868 4180 33908 4220
rect 34348 4180 34388 4220
rect 37132 4180 37172 4220
rect 37996 4180 38036 4220
rect 39340 4180 39380 4220
rect 42988 4180 43028 4220
rect 33004 4096 33044 4136
rect 33388 4096 33428 4136
rect 34732 4096 34772 4136
rect 36172 4096 36212 4136
rect 37516 4096 37556 4136
rect 39532 4096 39572 4136
rect 42028 4096 42068 4136
rect 43084 4096 43124 4136
rect 44524 4096 44564 4136
rect 44908 4096 44948 4136
rect 13612 4012 13652 4052
rect 16684 4012 16724 4052
rect 19276 4012 19316 4052
rect 20140 4012 20180 4052
rect 20524 4012 20564 4052
rect 23116 4012 23156 4052
rect 23980 4012 24020 4052
rect 34636 4012 34676 4052
rect 38476 4012 38516 4052
rect 39436 4012 39476 4052
rect 13228 3928 13268 3968
rect 14860 3928 14900 3968
rect 15628 3928 15668 3968
rect 17452 3928 17492 3968
rect 20428 3928 20468 3968
rect 20908 3928 20948 3968
rect 25708 3928 25748 3968
rect 28972 3928 29012 3968
rect 29740 3928 29780 3968
rect 30220 3928 30260 3968
rect 32140 3928 32180 3968
rect 32524 3928 32564 3968
rect 35596 3928 35636 3968
rect 39628 3928 39668 3968
rect 40204 3928 40244 3968
rect 41740 3928 41780 3968
rect 3688 3760 3728 3800
rect 3770 3760 3810 3800
rect 3852 3760 3892 3800
rect 3934 3760 3974 3800
rect 4016 3760 4056 3800
rect 7852 3844 7892 3884
rect 9676 3844 9716 3884
rect 14380 3844 14420 3884
rect 18412 3844 18452 3884
rect 18604 3844 18644 3884
rect 22636 3844 22676 3884
rect 31852 3844 31892 3884
rect 32332 3844 32372 3884
rect 6892 3760 6932 3800
rect 11116 3760 11156 3800
rect 18808 3760 18848 3800
rect 18890 3760 18930 3800
rect 18972 3760 19012 3800
rect 19054 3760 19094 3800
rect 19136 3760 19176 3800
rect 19468 3760 19508 3800
rect 32524 3760 32564 3800
rect 33928 3760 33968 3800
rect 34010 3760 34050 3800
rect 34092 3760 34132 3800
rect 34174 3760 34214 3800
rect 34256 3760 34296 3800
rect 35404 3760 35444 3800
rect 44428 3760 44468 3800
rect 13708 3676 13748 3716
rect 14188 3676 14228 3716
rect 29260 3676 29300 3716
rect 30604 3676 30644 3716
rect 36940 3676 36980 3716
rect 14572 3592 14612 3632
rect 15436 3592 15476 3632
rect 15628 3592 15668 3632
rect 18796 3592 18836 3632
rect 24844 3592 24884 3632
rect 25132 3592 25172 3632
rect 29644 3592 29684 3632
rect 40684 3592 40724 3632
rect 42220 3592 42260 3632
rect 6316 3508 6356 3548
rect 12460 3508 12500 3548
rect 13612 3508 13652 3548
rect 14284 3508 14324 3548
rect 15724 3508 15764 3548
rect 18604 3508 18644 3548
rect 76 3424 116 3464
rect 76 3256 116 3296
rect 8524 3424 8564 3464
rect 12940 3424 12980 3464
rect 13516 3424 13556 3464
rect 14860 3424 14900 3464
rect 3532 3340 3572 3380
rect 4108 3340 4148 3380
rect 4780 3340 4820 3380
rect 6988 3340 7028 3380
rect 7468 3340 7508 3380
rect 7660 3340 7700 3380
rect 7852 3256 7892 3296
rect 11980 3340 12020 3380
rect 13420 3340 13451 3380
rect 13451 3340 13460 3380
rect 9292 3256 9332 3296
rect 12364 3256 12404 3296
rect 12556 3256 12596 3296
rect 13324 3256 13364 3296
rect 15340 3424 15380 3464
rect 15628 3424 15668 3464
rect 31948 3508 31988 3548
rect 35020 3508 35060 3548
rect 43372 3508 43412 3548
rect 20524 3424 20564 3464
rect 21004 3424 21044 3464
rect 24748 3424 24788 3464
rect 25228 3424 25268 3464
rect 29548 3424 29588 3464
rect 30220 3424 30260 3464
rect 32140 3424 32180 3464
rect 34828 3424 34868 3464
rect 37324 3424 37364 3464
rect 37516 3424 37556 3464
rect 38572 3424 38612 3464
rect 39244 3424 39284 3464
rect 15724 3340 15764 3380
rect 16204 3340 16244 3380
rect 18892 3340 18932 3380
rect 20812 3340 20852 3380
rect 24076 3340 24116 3380
rect 24268 3340 24299 3380
rect 24299 3340 24308 3380
rect 24460 3340 24500 3380
rect 16012 3256 16052 3296
rect 26380 3340 26420 3380
rect 28876 3340 28916 3380
rect 29164 3340 29195 3380
rect 29195 3340 29204 3380
rect 29932 3340 29972 3380
rect 30412 3340 30452 3380
rect 31852 3340 31892 3380
rect 33292 3340 33332 3380
rect 35788 3340 35828 3380
rect 36172 3340 36212 3380
rect 18700 3256 18740 3296
rect 19372 3256 19412 3296
rect 21484 3256 21524 3296
rect 23020 3256 23060 3296
rect 24364 3256 24404 3296
rect 29356 3256 29396 3296
rect 31180 3256 31220 3296
rect 32812 3256 32852 3296
rect 33100 3256 33140 3296
rect 33676 3256 33716 3296
rect 40204 3340 40244 3380
rect 40684 3340 40724 3380
rect 42988 3340 43028 3380
rect 37900 3256 37940 3296
rect 38380 3256 38420 3296
rect 38668 3256 38708 3296
rect 42604 3256 42644 3296
rect 44140 3256 44180 3296
rect 45196 3256 45236 3296
rect 15436 3172 15476 3212
rect 16876 3172 16916 3212
rect 17740 3172 17780 3212
rect 19948 3172 19988 3212
rect 25420 3172 25460 3212
rect 27820 3172 27860 3212
rect 35404 3172 35444 3212
rect 39148 3172 39188 3212
rect 39820 3172 39860 3212
rect 40204 3172 40244 3212
rect 41932 3172 41963 3212
rect 41963 3172 41972 3212
rect 43084 3172 43115 3212
rect 43115 3172 43124 3212
rect 6028 3088 6068 3128
rect 8812 3088 8852 3128
rect 9292 3088 9332 3128
rect 11596 3088 11636 3128
rect 12556 3088 12596 3128
rect 15244 3088 15284 3128
rect 15724 3088 15764 3128
rect 31180 3088 31220 3128
rect 35596 3088 35636 3128
rect 39628 3088 39668 3128
rect 43756 3088 43796 3128
rect 4928 3004 4968 3044
rect 5010 3004 5050 3044
rect 5092 3004 5132 3044
rect 5174 3004 5214 3044
rect 5256 3004 5296 3044
rect 8908 3004 8948 3044
rect 15340 3004 15380 3044
rect 18892 3004 18932 3044
rect 20048 3004 20088 3044
rect 20130 3004 20170 3044
rect 20212 3004 20252 3044
rect 20294 3004 20334 3044
rect 20376 3004 20416 3044
rect 25132 3004 25172 3044
rect 29068 3004 29108 3044
rect 35020 3004 35060 3044
rect 35168 3004 35208 3044
rect 35250 3004 35290 3044
rect 35332 3004 35372 3044
rect 35414 3004 35454 3044
rect 35496 3004 35536 3044
rect 35788 3004 35828 3044
rect 44908 3004 44948 3044
rect 16876 2920 16916 2960
rect 25804 2920 25844 2960
rect 27436 2920 27476 2960
rect 29260 2920 29300 2960
rect 39916 2920 39956 2960
rect 40204 2920 40244 2960
rect 41932 2920 41972 2960
rect 7468 2836 7508 2876
rect 8620 2836 8660 2876
rect 9580 2836 9620 2876
rect 11212 2836 11252 2876
rect 15436 2836 15476 2876
rect 15628 2836 15668 2876
rect 15820 2836 15860 2876
rect 16012 2836 16052 2876
rect 17068 2836 17108 2876
rect 25132 2836 25172 2876
rect 28876 2836 28916 2876
rect 29452 2836 29492 2876
rect 34348 2836 34388 2876
rect 41260 2836 41300 2876
rect 41644 2836 41684 2876
rect 42028 2836 42068 2876
rect 42412 2836 42452 2876
rect 43084 2836 43115 2876
rect 43115 2836 43124 2876
rect 45196 2836 45236 2876
rect 10636 2752 10676 2792
rect 11500 2752 11540 2792
rect 5836 2668 5876 2708
rect 6892 2668 6932 2708
rect 7564 2668 7604 2708
rect 8812 2699 8852 2708
rect 8812 2668 8852 2699
rect 9772 2668 9812 2708
rect 18700 2752 18740 2792
rect 19276 2752 19316 2792
rect 11020 2699 11060 2708
rect 11020 2668 11060 2699
rect 6988 2584 7028 2624
rect 9388 2584 9428 2624
rect 12940 2668 12980 2708
rect 13228 2584 13268 2624
rect 13420 2584 13460 2624
rect 2860 2500 2900 2540
rect 10540 2500 10580 2540
rect 11596 2500 11636 2540
rect 15340 2668 15380 2708
rect 16012 2668 16052 2708
rect 16396 2668 16436 2708
rect 16780 2699 16820 2708
rect 16780 2668 16820 2699
rect 16972 2668 17012 2708
rect 18220 2668 18260 2708
rect 18988 2668 19028 2708
rect 19468 2668 19508 2708
rect 19948 2752 19988 2792
rect 20236 2752 20276 2792
rect 24364 2752 24404 2792
rect 25036 2752 25076 2792
rect 25324 2752 25364 2792
rect 26572 2752 26612 2792
rect 30124 2752 30164 2792
rect 32332 2752 32372 2792
rect 35500 2752 35540 2792
rect 36076 2752 36116 2792
rect 37900 2752 37940 2792
rect 38764 2752 38804 2792
rect 38956 2752 38996 2792
rect 20716 2699 20756 2708
rect 20716 2668 20756 2699
rect 21004 2668 21044 2708
rect 21580 2668 21620 2708
rect 22924 2668 22964 2708
rect 23212 2668 23252 2708
rect 23596 2668 23636 2708
rect 23884 2668 23924 2708
rect 24556 2668 24596 2708
rect 25516 2668 25556 2708
rect 25708 2668 25748 2708
rect 26284 2668 26324 2708
rect 27532 2668 27572 2708
rect 27820 2668 27860 2708
rect 15628 2584 15668 2624
rect 16204 2584 16244 2624
rect 20044 2584 20084 2624
rect 24076 2584 24116 2624
rect 27244 2584 27284 2624
rect 28300 2584 28340 2624
rect 15724 2500 15764 2540
rect 18988 2500 19028 2540
rect 19948 2500 19988 2540
rect 25996 2500 26036 2540
rect 26188 2500 26228 2540
rect 28780 2668 28820 2708
rect 29164 2668 29204 2708
rect 31180 2699 31220 2708
rect 31180 2668 31220 2699
rect 32044 2668 32084 2708
rect 32812 2668 32852 2708
rect 34924 2668 34964 2708
rect 35116 2668 35156 2708
rect 37132 2668 37172 2708
rect 37324 2668 37364 2708
rect 38668 2668 38699 2708
rect 38699 2668 38708 2708
rect 39148 2752 39188 2792
rect 42604 2752 42644 2792
rect 28684 2584 28724 2624
rect 29260 2584 29300 2624
rect 30412 2584 30452 2624
rect 30700 2584 30740 2624
rect 31852 2584 31892 2624
rect 33388 2584 33428 2624
rect 34444 2584 34484 2624
rect 41932 2584 41972 2624
rect 42124 2584 42164 2624
rect 43756 2584 43796 2624
rect 45196 2584 45236 2624
rect 31372 2500 31412 2540
rect 32044 2500 32084 2540
rect 32236 2500 32276 2540
rect 33580 2500 33620 2540
rect 38860 2500 38900 2540
rect 45100 2500 45140 2540
rect 2092 2416 2132 2456
rect 5164 2416 5204 2456
rect 8428 2416 8468 2456
rect 8716 2416 8756 2456
rect 11020 2416 11060 2456
rect 11212 2416 11252 2456
rect 12844 2416 12884 2456
rect 16588 2416 16628 2456
rect 18508 2416 18548 2456
rect 23212 2416 23252 2456
rect 12748 2332 12788 2372
rect 3688 2248 3728 2288
rect 3770 2248 3810 2288
rect 3852 2248 3892 2288
rect 3934 2248 3974 2288
rect 4016 2248 4056 2288
rect 1900 2080 1940 2120
rect 3532 2080 3572 2120
rect 29836 2416 29876 2456
rect 38668 2416 38708 2456
rect 38956 2416 38996 2456
rect 39340 2416 39380 2456
rect 43660 2416 43700 2456
rect 13228 2332 13268 2372
rect 16396 2332 16436 2372
rect 19276 2332 19316 2372
rect 22924 2332 22964 2372
rect 24844 2332 24884 2372
rect 25516 2332 25556 2372
rect 29740 2332 29780 2372
rect 31564 2332 31604 2372
rect 33388 2332 33428 2372
rect 37324 2332 37364 2372
rect 39052 2332 39092 2372
rect 41932 2332 41972 2372
rect 5836 2248 5876 2288
rect 12652 2248 12692 2288
rect 7852 2164 7892 2204
rect 8908 2164 8948 2204
rect 11980 2164 12020 2204
rect 18808 2248 18848 2288
rect 18890 2248 18930 2288
rect 18972 2248 19012 2288
rect 19054 2248 19094 2288
rect 19136 2248 19176 2288
rect 19468 2248 19508 2288
rect 22732 2248 22772 2288
rect 24940 2248 24980 2288
rect 25132 2248 25172 2288
rect 28780 2248 28820 2288
rect 33928 2248 33968 2288
rect 34010 2248 34050 2288
rect 34092 2248 34132 2288
rect 34174 2248 34214 2288
rect 34256 2248 34296 2288
rect 40300 2248 40340 2288
rect 41260 2248 41300 2288
rect 41452 2248 41492 2288
rect 15340 2164 15380 2204
rect 15532 2164 15572 2204
rect 16780 2164 16820 2204
rect 16972 2164 17012 2204
rect 29548 2164 29588 2204
rect 33772 2164 33812 2204
rect 34828 2164 34868 2204
rect 36076 2164 36116 2204
rect 37612 2164 37652 2204
rect 37900 2164 37940 2204
rect 42124 2164 42164 2204
rect 42508 2164 42548 2204
rect 44044 2164 44084 2204
rect 5932 2080 5972 2120
rect 6220 2080 6260 2120
rect 10348 2080 10388 2120
rect 11500 2080 11540 2120
rect 1228 1996 1268 2036
rect 5836 1996 5876 2036
rect 7756 1996 7796 2036
rect 9964 1996 10004 2036
rect 1420 1912 1460 1952
rect 3148 1912 3188 1952
rect 3916 1912 3956 1952
rect 4684 1912 4724 1952
rect 5164 1912 5204 1952
rect 5740 1912 5780 1952
rect 7564 1912 7604 1952
rect 1324 1828 1364 1868
rect 5452 1828 5492 1868
rect 6220 1828 6260 1868
rect 6892 1828 6932 1868
rect 76 1744 116 1784
rect 10060 1912 10100 1952
rect 10828 1912 10868 1952
rect 11596 1912 11636 1952
rect 12652 1912 12692 1952
rect 10540 1828 10580 1868
rect 12364 1828 12404 1868
rect 12844 1828 12884 1868
rect 9292 1744 9332 1784
rect 11980 1744 12020 1784
rect 13132 1744 13172 1784
rect 6124 1660 6164 1700
rect 7180 1660 7220 1700
rect 8716 1660 8756 1700
rect 11500 1660 11540 1700
rect 13036 1660 13076 1700
rect 76 1576 116 1616
rect 13900 2080 13940 2120
rect 16492 2080 16532 2120
rect 17164 2080 17204 2120
rect 20716 2080 20756 2120
rect 21004 2080 21044 2120
rect 22828 2080 22868 2120
rect 16684 1996 16724 2036
rect 17932 1996 17972 2036
rect 22636 1996 22676 2036
rect 25036 2080 25076 2120
rect 25996 2080 26036 2120
rect 34060 2080 34100 2120
rect 34924 2080 34964 2120
rect 37804 2080 37844 2120
rect 38092 2080 38132 2120
rect 40492 2080 40532 2120
rect 40972 2080 41012 2120
rect 25228 1996 25268 2036
rect 25900 1996 25940 2036
rect 30412 1996 30452 2036
rect 13420 1912 13460 1952
rect 14668 1912 14708 1952
rect 15436 1912 15476 1952
rect 15820 1912 15860 1952
rect 16300 1912 16340 1952
rect 16588 1912 16628 1952
rect 18124 1912 18164 1952
rect 19276 1912 19316 1952
rect 19756 1912 19796 1952
rect 20236 1912 20276 1952
rect 21676 1912 21716 1952
rect 23500 1912 23540 1952
rect 24748 1912 24788 1952
rect 25804 1912 25844 1952
rect 31372 1912 31412 1952
rect 31852 1912 31892 1952
rect 32140 1912 32180 1952
rect 34252 1912 34292 1952
rect 36172 1912 36212 1952
rect 37708 1912 37748 1952
rect 39916 1912 39956 1952
rect 13900 1828 13940 1868
rect 16204 1828 16244 1868
rect 17356 1828 17396 1868
rect 18028 1828 18068 1868
rect 18412 1828 18452 1868
rect 19372 1828 19412 1868
rect 20620 1828 20660 1868
rect 20908 1828 20948 1868
rect 22252 1828 22292 1868
rect 23692 1828 23732 1868
rect 23980 1828 24020 1868
rect 24364 1828 24395 1868
rect 24395 1828 24404 1868
rect 27148 1828 27188 1868
rect 27820 1828 27860 1868
rect 28684 1828 28724 1868
rect 28972 1828 29012 1868
rect 29260 1828 29291 1868
rect 29291 1828 29300 1868
rect 30700 1828 30740 1868
rect 35596 1828 35636 1868
rect 15532 1744 15572 1784
rect 16972 1744 17012 1784
rect 19852 1744 19892 1784
rect 23596 1744 23636 1784
rect 24076 1744 24116 1784
rect 24652 1744 24692 1784
rect 15436 1660 15476 1700
rect 16204 1660 16244 1700
rect 19564 1660 19604 1700
rect 19948 1660 19988 1700
rect 21580 1660 21620 1700
rect 45196 1996 45236 2036
rect 43372 1912 43412 1952
rect 41068 1828 41108 1868
rect 42700 1828 42740 1868
rect 43180 1828 43220 1868
rect 43756 1828 43796 1868
rect 44044 1912 44084 1952
rect 45100 1912 45140 1952
rect 43948 1828 43988 1868
rect 28780 1744 28820 1784
rect 29356 1744 29396 1784
rect 29548 1744 29588 1784
rect 30124 1744 30164 1784
rect 34444 1744 34484 1784
rect 34636 1744 34676 1784
rect 22348 1660 22388 1700
rect 23116 1660 23156 1700
rect 23884 1660 23924 1700
rect 24748 1660 24788 1700
rect 26956 1660 26996 1700
rect 34348 1660 34388 1700
rect 38764 1660 38804 1700
rect 19276 1576 19316 1616
rect 21772 1576 21812 1616
rect 24076 1576 24116 1616
rect 24940 1576 24980 1616
rect 32716 1576 32756 1616
rect 33580 1576 33620 1616
rect 38668 1576 38708 1616
rect 38956 1576 38996 1616
rect 42604 1576 42644 1616
rect 4928 1492 4968 1532
rect 5010 1492 5050 1532
rect 5092 1492 5132 1532
rect 5174 1492 5214 1532
rect 5256 1492 5296 1532
rect 5740 1492 5780 1532
rect 6988 1492 7028 1532
rect 13324 1492 13364 1532
rect 20048 1492 20088 1532
rect 20130 1492 20170 1532
rect 20212 1492 20252 1532
rect 20294 1492 20334 1532
rect 20376 1492 20416 1532
rect 20524 1492 20564 1532
rect 23308 1492 23348 1532
rect 23500 1492 23540 1532
rect 27628 1492 27668 1532
rect 27820 1492 27860 1532
rect 30124 1492 30164 1532
rect 32428 1492 32468 1532
rect 35168 1492 35208 1532
rect 35250 1492 35290 1532
rect 35332 1492 35372 1532
rect 35414 1492 35454 1532
rect 35496 1492 35536 1532
rect 42700 1492 42740 1532
rect 45004 1492 45044 1532
rect 7180 1408 7220 1448
rect 34828 1408 34868 1448
rect 44812 1408 44852 1448
rect 31372 1324 31412 1364
rect 1228 1240 1268 1280
rect 44620 1240 44660 1280
rect 1324 904 1364 944
rect 44812 904 44852 944
rect 1420 568 1460 608
rect 45004 568 45044 608
rect 14860 148 14900 188
rect 29260 148 29300 188
rect 27724 64 27764 104
rect 38860 64 38900 104
<< metal3 >>
rect 10540 11780 10580 11789
rect 11000 11780 11080 11844
rect 11000 11764 11020 11780
rect 1324 11024 1364 11033
rect 1132 10688 1172 10697
rect 1132 8840 1172 10648
rect 1324 9932 1364 10984
rect 1324 9883 1364 9892
rect 1420 10352 1460 10361
rect 1420 9596 1460 10312
rect 3436 10100 3476 10109
rect 1420 9547 1460 9556
rect 2284 10016 2324 10025
rect 1228 9512 1268 9521
rect 1228 9008 1268 9472
rect 1228 8959 1268 8968
rect 1132 8791 1172 8800
rect 2284 8756 2324 9976
rect 3436 9680 3476 10060
rect 8236 9932 8276 9941
rect 3688 9848 4056 9857
rect 3728 9808 3770 9848
rect 3810 9808 3852 9848
rect 3892 9808 3934 9848
rect 3974 9808 4016 9848
rect 3688 9799 4056 9808
rect 3436 9631 3476 9640
rect 6220 9764 6260 9773
rect 5740 9512 5780 9521
rect 2860 9260 2900 9269
rect 2860 9125 2900 9220
rect 4204 9260 4244 9269
rect 4108 9092 4148 9101
rect 4108 8840 4148 9052
rect 2284 8707 2324 8716
rect 3532 8756 3572 8765
rect 1132 8672 1172 8681
rect 1132 8084 1172 8632
rect 1132 8035 1172 8044
rect 1228 8000 1268 8009
rect 1228 7328 1268 7960
rect 1708 7748 1748 7757
rect 1708 7664 1748 7708
rect 1708 7613 1748 7624
rect 2860 7748 2900 7757
rect 2860 7613 2900 7708
rect 1228 7279 1268 7288
rect 76 7160 116 7169
rect 76 6992 116 7120
rect 76 6943 116 6952
rect 3532 7160 3572 8716
rect 3688 8336 4056 8345
rect 3728 8296 3770 8336
rect 3810 8296 3852 8336
rect 3892 8296 3934 8336
rect 3974 8296 4016 8336
rect 3688 8287 4056 8296
rect 4108 8000 4148 8800
rect 4108 7951 4148 7960
rect 76 6488 116 6497
rect 76 6320 116 6448
rect 76 6271 116 6280
rect 3532 6404 3572 7120
rect 3688 6824 4056 6833
rect 3728 6784 3770 6824
rect 3810 6784 3852 6824
rect 3892 6784 3934 6824
rect 3974 6784 4016 6824
rect 3688 6775 4056 6784
rect 3532 5732 3572 6364
rect 4204 6404 4244 9220
rect 4928 9092 5296 9101
rect 4968 9052 5010 9092
rect 5050 9052 5092 9092
rect 5132 9052 5174 9092
rect 5214 9052 5256 9092
rect 4928 9043 5296 9052
rect 5644 8756 5684 8765
rect 5740 8756 5780 9472
rect 5684 8716 5780 8756
rect 5644 8707 5684 8716
rect 5740 7916 5780 8716
rect 4928 7580 5296 7589
rect 4968 7540 5010 7580
rect 5050 7540 5092 7580
rect 5132 7540 5174 7580
rect 5214 7540 5256 7580
rect 4928 7531 5296 7540
rect 4300 6992 4340 7001
rect 4300 6857 4340 6952
rect 5740 6572 5780 7876
rect 5740 6523 5780 6532
rect 5836 9428 5876 9437
rect 4204 6355 4244 6364
rect 5740 6320 5780 6329
rect 5644 6236 5684 6245
rect 4928 6068 5296 6077
rect 4968 6028 5010 6068
rect 5050 6028 5092 6068
rect 5132 6028 5174 6068
rect 5214 6028 5256 6068
rect 4928 6019 5296 6028
rect 3532 5683 3572 5692
rect 4780 5732 4820 5741
rect 1996 5648 2036 5657
rect 1996 5060 2036 5608
rect 4684 5564 4724 5573
rect 3688 5312 4056 5321
rect 3728 5272 3770 5312
rect 3810 5272 3852 5312
rect 3892 5272 3934 5312
rect 3974 5272 4016 5312
rect 3688 5263 4056 5272
rect 1996 5011 2036 5020
rect 1612 4976 1652 4985
rect 76 4808 116 4817
rect 76 4640 116 4768
rect 76 4591 116 4600
rect 1612 4304 1652 4936
rect 4396 4892 4436 4903
rect 4396 4808 4436 4852
rect 4396 4759 4436 4768
rect 1612 4255 1652 4264
rect 76 4136 116 4145
rect 76 3968 116 4096
rect 76 3919 116 3928
rect 4108 4136 4148 4145
rect 3688 3800 4056 3809
rect 3728 3760 3770 3800
rect 3810 3760 3852 3800
rect 3892 3760 3934 3800
rect 3974 3760 4016 3800
rect 3688 3751 4056 3760
rect 76 3464 116 3473
rect 76 3296 116 3424
rect 76 3247 116 3256
rect 1900 3380 1940 3389
rect 1900 2120 1940 3340
rect 3532 3380 3572 3389
rect 2860 2540 2900 2549
rect 2092 2456 2132 2465
rect 2092 2321 2132 2416
rect 2860 2405 2900 2500
rect 1900 2071 1940 2080
rect 3532 2120 3572 3340
rect 4108 3380 4148 4096
rect 4108 3331 4148 3340
rect 4684 2708 4724 5524
rect 4780 3380 4820 5692
rect 5644 5732 5684 6196
rect 5644 5683 5684 5692
rect 5452 5480 5492 5489
rect 5452 4892 5492 5440
rect 5452 4843 5492 4852
rect 5740 4892 5780 6280
rect 5740 4843 5780 4852
rect 5836 5564 5876 9388
rect 5932 7748 5972 7757
rect 5932 6488 5972 7708
rect 5932 6439 5972 6448
rect 6220 6488 6260 9724
rect 8236 9680 8276 9892
rect 9964 9764 10004 9773
rect 10004 9724 10292 9764
rect 9964 9715 10004 9724
rect 8236 9631 8276 9640
rect 10252 9680 10292 9724
rect 10252 9631 10292 9640
rect 8140 9596 8180 9605
rect 7948 9512 7988 9521
rect 7660 9176 7700 9185
rect 6796 8756 6836 8765
rect 6796 7916 6836 8716
rect 6796 7867 6836 7876
rect 7180 8084 7220 8093
rect 4928 4556 5296 4565
rect 4968 4516 5010 4556
rect 5050 4516 5092 4556
rect 5132 4516 5174 4556
rect 5214 4516 5256 4556
rect 4928 4507 5296 4516
rect 4780 3331 4820 3340
rect 4928 3044 5296 3053
rect 4968 3004 5010 3044
rect 5050 3004 5092 3044
rect 5132 3004 5174 3044
rect 5214 3004 5256 3044
rect 4928 2995 5296 3004
rect 4684 2659 4724 2668
rect 5836 2708 5876 5524
rect 5836 2659 5876 2668
rect 5932 5816 5972 5825
rect 5164 2456 5204 2465
rect 3688 2288 4056 2297
rect 3728 2248 3770 2288
rect 3810 2248 3852 2288
rect 3892 2248 3934 2288
rect 3974 2248 4016 2288
rect 3688 2239 4056 2248
rect 3532 2071 3572 2080
rect 1228 2036 1268 2045
rect 76 1784 116 1793
rect 76 1616 116 1744
rect 76 1567 116 1576
rect 1228 1280 1268 1996
rect 1420 1952 1460 1961
rect 1228 1231 1268 1240
rect 1324 1868 1364 1877
rect 1324 944 1364 1828
rect 1324 895 1364 904
rect 1420 608 1460 1912
rect 1420 559 1460 568
rect 3148 1952 3188 1961
rect 3148 80 3188 1912
rect 3916 1952 3956 1961
rect 3916 80 3956 1912
rect 4684 1952 4724 1961
rect 4684 80 4724 1912
rect 5164 1952 5204 2416
rect 5836 2288 5876 2297
rect 5836 2036 5876 2248
rect 5932 2120 5972 5776
rect 6220 5732 6260 6448
rect 6220 5683 6260 5692
rect 6316 7160 6356 7169
rect 6316 5564 6356 7120
rect 7180 7160 7220 8044
rect 7180 7111 7220 7120
rect 6412 6488 6452 6497
rect 6412 6404 6452 6448
rect 6412 6353 6452 6364
rect 6700 6488 6740 6497
rect 6316 5515 6356 5524
rect 6028 5396 6068 5405
rect 6028 4724 6068 5356
rect 6412 5060 6452 5069
rect 6028 4675 6068 4684
rect 6316 4892 6356 4901
rect 6028 4220 6068 4229
rect 6028 3128 6068 4180
rect 6316 3548 6356 4852
rect 6412 4136 6452 5020
rect 6700 4892 6740 6448
rect 6796 6404 6836 6415
rect 6796 6320 6836 6364
rect 6796 6271 6836 6280
rect 6700 4843 6740 4852
rect 7468 6236 7508 6245
rect 6412 4087 6452 4096
rect 6892 4220 6932 4229
rect 6892 3800 6932 4180
rect 6892 3751 6932 3760
rect 6316 3499 6356 3508
rect 7468 3548 7508 6196
rect 7564 4892 7604 4901
rect 7564 4757 7604 4852
rect 7468 3499 7508 3508
rect 7660 4136 7700 9136
rect 7948 6908 7988 9472
rect 8044 9260 8084 9269
rect 8044 8924 8084 9220
rect 8044 8875 8084 8884
rect 8140 7160 8180 9556
rect 10060 9596 10100 9605
rect 8812 9512 8852 9521
rect 8620 9344 8660 9353
rect 8660 9304 8756 9344
rect 8620 9295 8660 9304
rect 8524 8840 8564 8849
rect 8524 8672 8564 8800
rect 8524 8623 8564 8632
rect 8140 7111 8180 7120
rect 8620 8588 8660 8597
rect 7948 6859 7988 6868
rect 8332 5480 8372 5489
rect 8044 4640 8084 4649
rect 7948 4304 7988 4313
rect 7948 4169 7988 4264
rect 8044 4220 8084 4600
rect 8332 4388 8372 5440
rect 8524 5144 8564 5153
rect 8524 4808 8564 5104
rect 8620 4892 8660 8548
rect 8716 5144 8756 9304
rect 8812 6404 8852 9472
rect 9292 9512 9332 9521
rect 9004 9428 9044 9437
rect 9004 8924 9044 9388
rect 9004 8875 9044 8884
rect 9196 8756 9236 8765
rect 9100 7580 9140 7589
rect 8812 6355 8852 6364
rect 8908 7160 8948 7169
rect 8908 5480 8948 7120
rect 9004 5732 9044 5741
rect 9100 5732 9140 7540
rect 9044 5692 9140 5732
rect 9004 5683 9044 5692
rect 8908 5431 8948 5440
rect 9004 5480 9044 5489
rect 8716 5095 8756 5104
rect 8660 4852 8756 4892
rect 8620 4843 8660 4852
rect 8524 4724 8564 4768
rect 8524 4684 8660 4724
rect 8620 4472 8660 4684
rect 8620 4423 8660 4432
rect 8332 4339 8372 4348
rect 8044 4171 8084 4180
rect 8620 4220 8660 4229
rect 6028 3079 6068 3088
rect 6988 3380 7028 3389
rect 6892 2708 6932 2717
rect 5932 2071 5972 2080
rect 6220 2120 6260 2129
rect 6220 2036 6260 2080
rect 5836 1987 5876 1996
rect 6124 1996 6260 2036
rect 5164 1903 5204 1912
rect 5740 1952 5780 1961
rect 5452 1868 5492 1877
rect 4928 1532 5296 1541
rect 4968 1492 5010 1532
rect 5050 1492 5092 1532
rect 5132 1492 5174 1532
rect 5214 1492 5256 1532
rect 4928 1483 5296 1492
rect 5452 80 5492 1828
rect 5740 1532 5780 1912
rect 6124 1700 6164 1996
rect 6124 1651 6164 1660
rect 6220 1868 6260 1877
rect 5740 1483 5780 1492
rect 6220 80 6260 1828
rect 6892 1868 6932 2668
rect 6988 2624 7028 3340
rect 7468 3380 7508 3389
rect 7468 2876 7508 3340
rect 7660 3380 7700 4096
rect 7660 3331 7700 3340
rect 7852 3884 7892 3893
rect 7468 2827 7508 2836
rect 7852 3296 7892 3844
rect 6988 2575 7028 2584
rect 7564 2708 7604 2717
rect 7564 1952 7604 2668
rect 7852 2204 7892 3256
rect 8524 3464 8564 3473
rect 8428 2456 8468 2467
rect 8428 2372 8468 2416
rect 8428 2323 8468 2332
rect 7852 2155 7892 2164
rect 7564 1903 7604 1912
rect 7756 2036 7796 2045
rect 6892 1819 6932 1828
rect 7180 1700 7220 1709
rect 6988 1532 7028 1541
rect 6988 80 7028 1492
rect 7180 1448 7220 1660
rect 7180 1399 7220 1408
rect 7756 80 7796 1996
rect 8524 80 8564 3424
rect 8620 2876 8660 4180
rect 8620 2827 8660 2836
rect 8716 2456 8756 4852
rect 8908 4304 8948 4313
rect 8812 3128 8852 3137
rect 8812 2708 8852 3088
rect 8908 3044 8948 4264
rect 9004 4136 9044 5440
rect 9100 4640 9140 5692
rect 9100 4591 9140 4600
rect 9196 6320 9236 8716
rect 9196 6152 9236 6280
rect 9196 4976 9236 6112
rect 9196 4304 9236 4936
rect 9196 4255 9236 4264
rect 9292 4304 9332 9472
rect 9484 9344 9524 9353
rect 9484 8756 9524 9304
rect 9964 9344 10004 9353
rect 9484 8621 9524 8716
rect 9580 9176 9620 9185
rect 9580 8672 9620 9136
rect 9964 8840 10004 9304
rect 9964 8791 10004 8800
rect 9580 8623 9620 8632
rect 9964 8084 10004 8093
rect 9484 8000 9524 8009
rect 9292 4255 9332 4264
rect 9388 6404 9428 6413
rect 9004 4087 9044 4096
rect 9292 3296 9332 3305
rect 9292 3128 9332 3256
rect 9292 3079 9332 3088
rect 8908 2995 8948 3004
rect 8812 2659 8852 2668
rect 8716 1700 8756 2416
rect 8908 2624 8948 2633
rect 8908 2204 8948 2584
rect 9388 2624 9428 6364
rect 9484 4808 9524 7960
rect 9868 7580 9908 7589
rect 9676 7412 9716 7421
rect 9676 6488 9716 7372
rect 9676 6439 9716 6448
rect 9772 7328 9812 7337
rect 9484 4759 9524 4768
rect 9676 5816 9716 5825
rect 9676 4976 9716 5776
rect 9484 4640 9524 4649
rect 9484 4220 9524 4600
rect 9484 4171 9524 4180
rect 9676 4304 9716 4936
rect 9772 5648 9812 7288
rect 9772 4892 9812 5608
rect 9772 4843 9812 4852
rect 9676 3884 9716 4264
rect 9676 3835 9716 3844
rect 9580 3464 9620 3473
rect 9580 2876 9620 3424
rect 9868 3464 9908 7540
rect 9964 6908 10004 8044
rect 9964 6859 10004 6868
rect 10060 5648 10100 9556
rect 10252 9428 10292 9437
rect 10252 9293 10292 9388
rect 10348 9344 10388 9353
rect 10252 8840 10292 8849
rect 10156 8756 10196 8765
rect 10156 7916 10196 8716
rect 10252 8168 10292 8800
rect 10252 8119 10292 8128
rect 10156 7867 10196 7876
rect 10348 7832 10388 9304
rect 10156 6572 10196 6581
rect 10156 6404 10196 6532
rect 10252 6572 10292 6583
rect 10252 6488 10292 6532
rect 10252 6439 10292 6448
rect 10156 6355 10196 6364
rect 10252 6320 10292 6329
rect 10252 6152 10292 6280
rect 10252 6103 10292 6112
rect 10060 5599 10100 5608
rect 10348 5816 10388 7792
rect 10444 9260 10484 9269
rect 10444 7412 10484 9220
rect 10444 7363 10484 7372
rect 10444 7244 10484 7253
rect 10444 6320 10484 7204
rect 10540 6992 10580 11740
rect 11060 11764 11080 11780
rect 11192 11764 11272 11844
rect 11384 11764 11464 11844
rect 11576 11764 11656 11844
rect 11768 11764 11848 11844
rect 11960 11764 12040 11844
rect 12152 11764 12232 11844
rect 12344 11764 12424 11844
rect 12536 11764 12616 11844
rect 12728 11764 12808 11844
rect 12920 11764 13000 11844
rect 13112 11764 13192 11844
rect 13304 11764 13384 11844
rect 13496 11764 13576 11844
rect 13688 11764 13768 11844
rect 13880 11764 13960 11844
rect 14072 11764 14152 11844
rect 14264 11764 14344 11844
rect 14456 11764 14536 11844
rect 14648 11764 14728 11844
rect 14840 11764 14920 11844
rect 15032 11764 15112 11844
rect 15224 11764 15304 11844
rect 15416 11764 15496 11844
rect 15608 11764 15688 11844
rect 15800 11764 15880 11844
rect 15992 11764 16072 11844
rect 16184 11764 16264 11844
rect 16376 11764 16456 11844
rect 16568 11764 16648 11844
rect 16760 11764 16840 11844
rect 16952 11764 17032 11844
rect 17144 11764 17224 11844
rect 17336 11764 17416 11844
rect 17528 11764 17608 11844
rect 17720 11764 17800 11844
rect 17912 11764 17992 11844
rect 18104 11764 18184 11844
rect 18296 11764 18376 11844
rect 18488 11764 18568 11844
rect 18680 11764 18760 11844
rect 18872 11764 18952 11844
rect 19064 11764 19144 11844
rect 19256 11764 19336 11844
rect 19448 11764 19528 11844
rect 19640 11764 19720 11844
rect 19832 11764 19912 11844
rect 20024 11764 20104 11844
rect 20216 11764 20296 11844
rect 20408 11764 20488 11844
rect 20600 11764 20680 11844
rect 20792 11764 20872 11844
rect 20984 11764 21064 11844
rect 21176 11764 21256 11844
rect 21368 11764 21448 11844
rect 21560 11764 21640 11844
rect 21752 11764 21832 11844
rect 21944 11764 22024 11844
rect 22136 11764 22216 11844
rect 22328 11764 22408 11844
rect 22520 11764 22600 11844
rect 22712 11764 22792 11844
rect 22904 11764 22984 11844
rect 23096 11764 23176 11844
rect 23288 11764 23368 11844
rect 23480 11764 23560 11844
rect 23672 11764 23752 11844
rect 23864 11764 23944 11844
rect 24056 11764 24136 11844
rect 24248 11764 24328 11844
rect 24440 11764 24520 11844
rect 24632 11764 24712 11844
rect 24824 11764 24904 11844
rect 25016 11764 25096 11844
rect 25208 11764 25288 11844
rect 25400 11764 25480 11844
rect 25592 11764 25672 11844
rect 25784 11764 25864 11844
rect 25976 11764 26056 11844
rect 26168 11764 26248 11844
rect 26360 11764 26440 11844
rect 26552 11764 26632 11844
rect 26744 11764 26824 11844
rect 26936 11764 27016 11844
rect 27128 11764 27208 11844
rect 27320 11764 27400 11844
rect 27512 11764 27592 11844
rect 27704 11764 27784 11844
rect 27896 11764 27976 11844
rect 28088 11764 28168 11844
rect 28280 11764 28360 11844
rect 28472 11764 28552 11844
rect 28664 11764 28744 11844
rect 28856 11764 28936 11844
rect 29048 11764 29128 11844
rect 29240 11764 29320 11844
rect 29432 11764 29512 11844
rect 29624 11764 29704 11844
rect 29816 11764 29896 11844
rect 30008 11764 30088 11844
rect 30200 11764 30280 11844
rect 30392 11764 30472 11844
rect 30584 11764 30664 11844
rect 30776 11764 30856 11844
rect 30968 11764 31048 11844
rect 31160 11764 31240 11844
rect 31352 11764 31432 11844
rect 31544 11764 31624 11844
rect 31736 11764 31816 11844
rect 31928 11764 32008 11844
rect 32120 11764 32200 11844
rect 32312 11764 32392 11844
rect 32504 11764 32584 11844
rect 32696 11764 32776 11844
rect 32888 11764 32968 11844
rect 33080 11764 33160 11844
rect 33272 11764 33352 11844
rect 33464 11764 33544 11844
rect 33656 11764 33736 11844
rect 33848 11764 33928 11844
rect 34040 11764 34120 11844
rect 34232 11764 34312 11844
rect 34424 11764 34504 11844
rect 34616 11764 34696 11844
rect 34808 11764 34888 11844
rect 35000 11764 35080 11844
rect 11020 11731 11060 11740
rect 10636 10016 10676 10025
rect 10636 9344 10676 9976
rect 10636 9176 10676 9304
rect 10636 9127 10676 9136
rect 10924 9848 10964 9857
rect 10732 8924 10772 8933
rect 10732 8789 10772 8884
rect 10636 8084 10676 8179
rect 10636 8035 10676 8044
rect 10828 8000 10868 8009
rect 10636 7916 10676 7925
rect 10636 7781 10676 7876
rect 10732 7328 10772 7423
rect 10732 7279 10772 7288
rect 10540 6943 10580 6952
rect 10636 7244 10676 7253
rect 10636 6404 10676 7204
rect 10732 7160 10772 7169
rect 10732 6992 10772 7120
rect 10732 6943 10772 6952
rect 10636 6355 10676 6364
rect 10732 6572 10772 6581
rect 10444 6271 10484 6280
rect 9868 3415 9908 3424
rect 9964 4808 10004 4817
rect 9964 4472 10004 4768
rect 9580 2827 9620 2836
rect 9388 2575 9428 2584
rect 9772 2708 9812 2717
rect 9772 2573 9812 2668
rect 8908 2155 8948 2164
rect 9964 2036 10004 4432
rect 10060 4220 10100 4229
rect 10060 4085 10100 4180
rect 10348 2120 10388 5776
rect 10540 5480 10580 5489
rect 10540 4472 10580 5440
rect 10540 4423 10580 4432
rect 10732 4472 10772 6532
rect 10732 4423 10772 4432
rect 10828 2900 10868 7960
rect 10924 4556 10964 9808
rect 11116 8504 11156 8513
rect 11020 8420 11060 8429
rect 11020 7244 11060 8380
rect 11116 8000 11156 8464
rect 11116 7951 11156 7960
rect 11020 7195 11060 7204
rect 11020 7076 11060 7085
rect 11020 6488 11060 7036
rect 11116 6992 11156 7001
rect 11212 6992 11252 11764
rect 11156 6952 11252 6992
rect 11308 9512 11348 9521
rect 11116 6943 11156 6952
rect 11212 6824 11252 6833
rect 11116 6740 11156 6749
rect 11116 6656 11156 6700
rect 11116 6605 11156 6616
rect 11020 5732 11060 6448
rect 11020 5683 11060 5692
rect 11116 6236 11156 6245
rect 10924 4507 10964 4516
rect 11020 4724 11060 4733
rect 11020 4136 11060 4684
rect 11020 4087 11060 4096
rect 11116 3800 11156 6196
rect 11212 6068 11252 6784
rect 11212 6019 11252 6028
rect 11308 5732 11348 9472
rect 11308 5683 11348 5692
rect 11404 5144 11444 11764
rect 11500 8840 11540 8849
rect 11500 8756 11540 8800
rect 11500 8705 11540 8716
rect 11500 8084 11540 8095
rect 11500 8000 11540 8044
rect 11500 7951 11540 7960
rect 11500 7664 11540 7673
rect 11500 6572 11540 7624
rect 11596 6740 11636 11764
rect 11788 9932 11828 11764
rect 11788 9883 11828 9892
rect 11980 9680 12020 11764
rect 11788 9640 12020 9680
rect 12076 9932 12116 9941
rect 12076 9680 12116 9892
rect 11788 8084 11828 9640
rect 12076 9631 12116 9640
rect 11884 9512 11924 9521
rect 11924 9472 12116 9512
rect 11884 9463 11924 9472
rect 11980 8756 12020 8765
rect 11788 8035 11828 8044
rect 11884 8672 11924 8681
rect 11596 6691 11636 6700
rect 11692 7160 11732 7169
rect 11500 6532 11636 6572
rect 11500 6404 11540 6413
rect 11500 5816 11540 6364
rect 11500 5767 11540 5776
rect 11404 5095 11444 5104
rect 11116 3751 11156 3760
rect 11212 4892 11252 4901
rect 10636 2860 10868 2900
rect 11212 2876 11252 4852
rect 11596 4892 11636 6532
rect 11692 5144 11732 7120
rect 11788 6992 11828 7001
rect 11788 5648 11828 6952
rect 11884 6236 11924 8632
rect 11980 8420 12020 8716
rect 11980 8371 12020 8380
rect 11980 8000 12020 8009
rect 11980 7865 12020 7960
rect 11884 6187 11924 6196
rect 11980 7160 12020 7169
rect 11788 5599 11828 5608
rect 11884 6068 11924 6077
rect 11692 5095 11732 5104
rect 11596 4843 11636 4852
rect 11692 4976 11732 4985
rect 11692 4304 11732 4936
rect 11884 4976 11924 6028
rect 11980 5648 12020 7120
rect 11980 5599 12020 5608
rect 11924 4936 12020 4976
rect 11884 4927 11924 4936
rect 11692 4255 11732 4264
rect 11980 4220 12020 4936
rect 11980 3380 12020 4180
rect 11980 3331 12020 3340
rect 10636 2792 10676 2860
rect 11212 2827 11252 2836
rect 11596 3128 11636 3137
rect 10636 2743 10676 2752
rect 11500 2792 11540 2801
rect 11020 2708 11060 2717
rect 10348 2071 10388 2080
rect 10540 2540 10580 2549
rect 9964 1987 10004 1996
rect 10060 1952 10100 1961
rect 8716 1651 8756 1660
rect 9292 1784 9332 1793
rect 9292 80 9332 1744
rect 10060 80 10100 1912
rect 10540 1868 10580 2500
rect 11020 2456 11060 2668
rect 11020 2407 11060 2416
rect 11212 2456 11252 2465
rect 11212 2372 11252 2416
rect 11212 2321 11252 2332
rect 11500 2120 11540 2752
rect 11596 2540 11636 3088
rect 11596 2491 11636 2500
rect 11980 3128 12020 3137
rect 11980 2204 12020 3088
rect 12076 2900 12116 9472
rect 12172 7832 12212 11764
rect 12268 9512 12308 9521
rect 12268 8672 12308 9472
rect 12268 8623 12308 8632
rect 12172 7783 12212 7792
rect 12172 7664 12212 7673
rect 12172 6572 12212 7624
rect 12172 6523 12212 6532
rect 12268 6572 12308 6583
rect 12268 6488 12308 6532
rect 12268 6439 12308 6448
rect 12268 6236 12308 6245
rect 12172 4724 12212 4733
rect 12172 4589 12212 4684
rect 12268 4304 12308 6196
rect 12364 5648 12404 11764
rect 12460 8420 12500 8429
rect 12460 6068 12500 8380
rect 12556 6656 12596 11764
rect 12652 10016 12692 10027
rect 12652 9932 12692 9976
rect 12652 9883 12692 9892
rect 12652 9428 12692 9437
rect 12652 7916 12692 9388
rect 12652 7496 12692 7876
rect 12652 7447 12692 7456
rect 12748 6908 12788 11764
rect 12940 11444 12980 11764
rect 13132 11528 13172 11764
rect 13132 11488 13268 11528
rect 12940 11404 13172 11444
rect 12844 10016 12884 10025
rect 12844 9680 12884 9976
rect 12844 9631 12884 9640
rect 13132 9260 13172 11404
rect 13132 9211 13172 9220
rect 12844 9092 12884 9101
rect 12844 9008 12884 9052
rect 12844 8957 12884 8968
rect 13036 9092 13076 9101
rect 12940 8756 12980 8765
rect 12940 8504 12980 8716
rect 12940 8455 12980 8464
rect 13036 7916 13076 9052
rect 13228 8756 13268 11488
rect 13324 9848 13364 11764
rect 13420 10016 13460 10025
rect 13420 9881 13460 9976
rect 13324 9799 13364 9808
rect 13420 9512 13460 9521
rect 13228 8716 13364 8756
rect 13132 8672 13172 8681
rect 13132 8084 13172 8632
rect 13132 8035 13172 8044
rect 13228 8588 13268 8597
rect 13036 7832 13076 7876
rect 13036 7752 13076 7792
rect 12940 7244 12980 7339
rect 12940 7195 12980 7204
rect 13132 7328 13172 7337
rect 12748 6859 12788 6868
rect 12844 7160 12884 7169
rect 12556 6607 12596 6616
rect 12748 6740 12788 6749
rect 12748 6605 12788 6700
rect 12460 6019 12500 6028
rect 12556 6488 12596 6497
rect 12364 5599 12404 5608
rect 12556 4976 12596 6448
rect 12652 6404 12692 6413
rect 12652 6068 12692 6364
rect 12652 6019 12692 6028
rect 12748 5984 12788 5993
rect 12748 5849 12788 5944
rect 12748 5564 12788 5573
rect 12652 5480 12692 5489
rect 12652 5312 12692 5440
rect 12652 5263 12692 5272
rect 12748 5312 12788 5524
rect 12748 5263 12788 5272
rect 12748 5144 12788 5153
rect 12652 4976 12692 4985
rect 12556 4936 12652 4976
rect 12652 4927 12692 4936
rect 12460 4892 12500 4901
rect 12460 4808 12500 4852
rect 12748 4808 12788 5104
rect 12460 4768 12788 4808
rect 12268 4255 12308 4264
rect 12844 3968 12884 7120
rect 13036 7160 13076 7169
rect 12940 6992 12980 7001
rect 12940 6824 12980 6952
rect 12940 6775 12980 6784
rect 12940 5900 12980 5909
rect 12940 5765 12980 5860
rect 13036 5816 13076 7120
rect 13036 5767 13076 5776
rect 13132 5648 13172 7288
rect 13228 6320 13268 8548
rect 13324 6824 13364 8716
rect 13324 6775 13364 6784
rect 13420 6572 13460 9472
rect 13516 7076 13556 11764
rect 13708 10016 13748 11764
rect 13612 9976 13748 10016
rect 13612 8168 13652 9976
rect 13612 8119 13652 8128
rect 13708 9596 13748 9605
rect 13900 9596 13940 11764
rect 13900 9556 14036 9596
rect 13516 7027 13556 7036
rect 13612 8000 13652 8009
rect 13516 6740 13556 6749
rect 13516 6656 13556 6700
rect 13516 6605 13556 6616
rect 13324 6532 13460 6572
rect 13324 6488 13364 6532
rect 13324 6448 13460 6488
rect 13420 6404 13460 6448
rect 13420 6364 13556 6404
rect 13228 6280 13460 6320
rect 13324 6152 13364 6161
rect 13324 6017 13364 6112
rect 13132 5599 13172 5608
rect 12940 5564 12980 5573
rect 12940 5429 12980 5524
rect 13324 4724 13364 4733
rect 13324 4388 13364 4684
rect 13324 4339 13364 4348
rect 12844 3919 12884 3928
rect 13132 4220 13172 4229
rect 12364 3632 12404 3641
rect 12364 3296 12404 3592
rect 12460 3548 12500 3557
rect 12460 3464 12500 3508
rect 12460 3413 12500 3424
rect 12940 3464 12980 3473
rect 12940 3329 12980 3424
rect 12364 3247 12404 3256
rect 12556 3296 12596 3305
rect 12556 3128 12596 3256
rect 12556 3079 12596 3088
rect 12940 2960 12980 2969
rect 12076 2860 12596 2900
rect 11980 2155 12020 2164
rect 11500 2071 11540 2080
rect 10540 1819 10580 1828
rect 10828 1952 10868 1961
rect 10828 80 10868 1912
rect 11596 1952 11636 1961
rect 12556 1952 12596 2860
rect 12940 2708 12980 2920
rect 13132 2960 13172 4180
rect 13228 3968 13268 3979
rect 13228 3884 13268 3928
rect 13228 3835 13268 3844
rect 13420 3716 13460 6280
rect 13420 3667 13460 3676
rect 13420 3464 13460 3473
rect 13420 3380 13460 3424
rect 13516 3464 13556 6364
rect 13612 4724 13652 7960
rect 13708 6992 13748 9556
rect 13804 9176 13844 9185
rect 13804 8924 13844 9136
rect 13804 8875 13844 8884
rect 13708 6943 13748 6952
rect 13804 8672 13844 8681
rect 13612 4675 13652 4684
rect 13708 4220 13748 4229
rect 13612 4052 13652 4061
rect 13612 3548 13652 4012
rect 13708 4052 13748 4180
rect 13708 4003 13748 4012
rect 13708 3800 13748 3809
rect 13708 3716 13748 3760
rect 13708 3665 13748 3676
rect 13612 3499 13652 3508
rect 13516 3415 13556 3424
rect 13420 3329 13460 3340
rect 13132 2911 13172 2920
rect 13324 3296 13364 3305
rect 12940 2659 12980 2668
rect 13228 2876 13268 2885
rect 13228 2624 13268 2836
rect 13324 2624 13364 3256
rect 13804 3296 13844 8632
rect 13900 8504 13940 8513
rect 13900 7328 13940 8464
rect 13900 7279 13940 7288
rect 13900 7160 13940 7169
rect 13900 6320 13940 7120
rect 13996 6824 14036 9556
rect 14092 8084 14132 11764
rect 14284 9596 14324 11764
rect 14284 9547 14324 9556
rect 14380 9932 14420 9941
rect 14284 9428 14324 9437
rect 14188 9344 14228 9353
rect 14188 8756 14228 9304
rect 14188 8707 14228 8716
rect 14092 8035 14132 8044
rect 14188 7412 14228 7421
rect 13996 6775 14036 6784
rect 14092 7076 14132 7085
rect 13900 6271 13940 6280
rect 13996 6236 14036 6245
rect 13996 6068 14036 6196
rect 13996 6019 14036 6028
rect 13900 5984 13940 5993
rect 13900 5816 13940 5944
rect 13900 5767 13940 5776
rect 13996 5900 14036 5909
rect 13996 5765 14036 5860
rect 13900 5564 13940 5573
rect 13900 4892 13940 5524
rect 13900 4843 13940 4852
rect 13804 3247 13844 3256
rect 13420 2624 13460 2633
rect 13324 2584 13420 2624
rect 13228 2575 13268 2584
rect 12844 2456 12884 2465
rect 12748 2372 12788 2381
rect 12652 2288 12692 2299
rect 12652 2204 12692 2248
rect 12652 2155 12692 2164
rect 12748 2036 12788 2332
rect 12748 1987 12788 1996
rect 12652 1952 12692 1961
rect 12556 1912 12652 1952
rect 11500 1700 11540 1709
rect 11500 1565 11540 1660
rect 11596 80 11636 1912
rect 12652 1903 12692 1912
rect 12364 1868 12404 1877
rect 11980 1784 12020 1793
rect 11980 1649 12020 1744
rect 12364 80 12404 1828
rect 12844 1868 12884 2416
rect 13228 2372 13268 2381
rect 12940 2036 12980 2045
rect 13228 2036 13268 2332
rect 12980 1996 13268 2036
rect 12940 1987 12980 1996
rect 13420 1952 13460 2584
rect 13900 2120 13940 2215
rect 13900 2071 13940 2080
rect 12844 1819 12884 1828
rect 13036 1912 13420 1952
rect 13036 1700 13076 1912
rect 13420 1903 13460 1912
rect 13900 1868 13940 1877
rect 13036 1651 13076 1660
rect 13132 1784 13172 1793
rect 13132 80 13172 1744
rect 13324 1532 13364 1541
rect 13324 1397 13364 1492
rect 13900 80 13940 1828
rect 14092 1868 14132 7036
rect 14188 5648 14228 7372
rect 14188 5599 14228 5608
rect 14188 5228 14228 5323
rect 14188 5179 14228 5188
rect 14188 5060 14228 5069
rect 14188 4136 14228 5020
rect 14188 4087 14228 4096
rect 14188 3800 14228 3811
rect 14188 3716 14228 3760
rect 14188 3667 14228 3676
rect 14284 3548 14324 9388
rect 14380 8504 14420 9892
rect 14380 7916 14420 8464
rect 14380 7160 14420 7876
rect 14476 7244 14516 11764
rect 14572 8336 14612 8345
rect 14572 7832 14612 8296
rect 14572 7783 14612 7792
rect 14476 7195 14516 7204
rect 14380 7111 14420 7120
rect 14572 7160 14612 7169
rect 14380 6992 14420 7001
rect 14380 6740 14420 6952
rect 14380 6691 14420 6700
rect 14380 6488 14420 6497
rect 14380 3884 14420 6448
rect 14572 5900 14612 7120
rect 14668 6740 14708 11764
rect 14764 9512 14804 9521
rect 14764 8672 14804 9472
rect 14764 8623 14804 8632
rect 14764 8252 14804 8261
rect 14764 7580 14804 8212
rect 14764 7531 14804 7540
rect 14860 7076 14900 11764
rect 15052 9932 15092 11764
rect 15052 9883 15092 9892
rect 15148 9428 15188 9437
rect 15148 9176 15188 9388
rect 15148 9127 15188 9136
rect 14860 7027 14900 7036
rect 14956 8840 14996 8849
rect 14668 6691 14708 6700
rect 14764 6992 14804 7001
rect 14764 6656 14804 6952
rect 14764 6607 14804 6616
rect 14476 5860 14612 5900
rect 14668 6404 14708 6413
rect 14956 6404 14996 8800
rect 15148 8840 15188 8935
rect 15148 8791 15188 8800
rect 15148 8672 15188 8681
rect 15052 7748 15092 7757
rect 15052 7496 15092 7708
rect 15052 7447 15092 7456
rect 15052 6404 15092 6413
rect 14956 6364 15052 6404
rect 14476 4472 14516 5860
rect 14668 5732 14708 6364
rect 15052 6355 15092 6364
rect 15148 6068 15188 8632
rect 15244 6656 15284 11764
rect 15436 9680 15476 11764
rect 15436 9631 15476 9640
rect 15436 9512 15476 9521
rect 15436 9008 15476 9472
rect 15436 8959 15476 8968
rect 15628 8840 15668 11764
rect 15820 10100 15860 11764
rect 15820 10051 15860 10060
rect 15820 9848 15860 9857
rect 15820 9512 15860 9808
rect 15820 9463 15860 9472
rect 15628 8791 15668 8800
rect 15724 9092 15764 9101
rect 15340 8756 15380 8765
rect 15340 7916 15380 8716
rect 15340 7867 15380 7876
rect 15244 6607 15284 6616
rect 15340 7748 15380 7757
rect 15148 6019 15188 6028
rect 14708 5692 14804 5732
rect 14668 5683 14708 5692
rect 14668 5564 14708 5573
rect 14476 4423 14516 4432
rect 14572 5312 14612 5321
rect 14380 3835 14420 3844
rect 14572 3632 14612 5272
rect 14668 5060 14708 5524
rect 14764 5228 14804 5692
rect 14764 5179 14804 5188
rect 15148 5480 15188 5489
rect 14668 5011 14708 5020
rect 14764 4976 14804 4985
rect 14668 4388 14708 4399
rect 14668 4304 14708 4348
rect 14668 4255 14708 4264
rect 14572 3583 14612 3592
rect 14284 3499 14324 3508
rect 14764 2900 14804 4936
rect 15148 4472 15188 5440
rect 15148 4423 15188 4432
rect 15244 4640 15284 4649
rect 15148 4304 15188 4313
rect 14860 3968 14900 3977
rect 14860 3464 14900 3928
rect 14860 3415 14900 3424
rect 14764 2860 14900 2900
rect 14092 1819 14132 1828
rect 14476 2372 14516 2381
rect 14476 1532 14516 2332
rect 14476 1483 14516 1492
rect 14668 1952 14708 1961
rect 14668 80 14708 1912
rect 14860 188 14900 2860
rect 15148 2624 15188 4264
rect 15244 3128 15284 4600
rect 15340 3464 15380 7708
rect 15532 7580 15572 7589
rect 15436 7496 15476 7505
rect 15436 5480 15476 7456
rect 15532 7445 15572 7540
rect 15436 5431 15476 5440
rect 15532 7160 15572 7169
rect 15532 5312 15572 7120
rect 15628 5564 15668 5573
rect 15628 5429 15668 5524
rect 15532 5263 15572 5272
rect 15532 4892 15572 4901
rect 15436 4220 15476 4229
rect 15436 3632 15476 4180
rect 15436 3583 15476 3592
rect 15340 3415 15380 3424
rect 15244 3079 15284 3088
rect 15436 3212 15476 3221
rect 15340 3044 15380 3053
rect 15340 2909 15380 3004
rect 15436 2876 15476 3172
rect 15436 2827 15476 2836
rect 15148 2575 15188 2584
rect 15340 2708 15380 2717
rect 15340 2204 15380 2668
rect 15532 2624 15572 4852
rect 15628 4388 15668 4397
rect 15628 4220 15668 4348
rect 15628 4171 15668 4180
rect 15628 4052 15668 4063
rect 15628 3968 15668 4012
rect 15628 3919 15668 3928
rect 15628 3632 15668 3641
rect 15628 3464 15668 3592
rect 15724 3548 15764 9052
rect 15820 8756 15860 8765
rect 15820 8504 15860 8716
rect 15820 8455 15860 8464
rect 15916 8672 15956 8681
rect 15820 7916 15860 7925
rect 15820 6152 15860 7876
rect 15916 7832 15956 8632
rect 15916 7783 15956 7792
rect 15916 7160 15956 7169
rect 15916 6740 15956 7120
rect 16012 6992 16052 11764
rect 16204 9512 16244 11764
rect 16204 9463 16244 9472
rect 16300 10100 16340 10109
rect 16108 9428 16148 9437
rect 16108 8756 16148 9388
rect 16108 8707 16148 8716
rect 16204 9008 16244 9017
rect 16012 6943 16052 6952
rect 16108 7160 16148 7169
rect 16204 7160 16244 8968
rect 16300 8924 16340 10060
rect 16300 8875 16340 8884
rect 16300 8000 16340 8009
rect 16300 7328 16340 7960
rect 16300 7279 16340 7288
rect 16300 7160 16340 7169
rect 16204 7120 16300 7160
rect 15916 6691 15956 6700
rect 15820 5900 15860 6112
rect 16012 6404 16052 6413
rect 16012 6152 16052 6364
rect 16108 6320 16148 7120
rect 16300 7111 16340 7120
rect 16396 6824 16436 11764
rect 16588 8840 16628 11764
rect 16588 8791 16628 8800
rect 16780 7328 16820 11764
rect 16492 7288 16820 7328
rect 16492 7244 16532 7288
rect 16492 7195 16532 7204
rect 16684 7160 16724 7169
rect 16396 6775 16436 6784
rect 16492 7076 16532 7085
rect 16492 6740 16532 7036
rect 16492 6691 16532 6700
rect 16108 6271 16148 6280
rect 16012 6103 16052 6112
rect 15820 5851 15860 5860
rect 16492 5816 16532 5825
rect 15916 5732 15956 5741
rect 15916 5480 15956 5692
rect 15916 5431 15956 5440
rect 16492 4892 16532 5776
rect 16492 4843 16532 4852
rect 15820 4808 15860 4817
rect 15820 4640 15860 4768
rect 15820 4591 15860 4600
rect 16492 4472 16532 4481
rect 15820 4388 15860 4397
rect 15820 4136 15860 4348
rect 15820 4087 15860 4096
rect 15724 3499 15764 3508
rect 15628 3415 15668 3424
rect 16204 3464 16244 3473
rect 15724 3380 15764 3389
rect 15724 3128 15764 3340
rect 16204 3380 16244 3424
rect 16204 3329 16244 3340
rect 15628 3044 15668 3053
rect 15628 2876 15668 3004
rect 15628 2827 15668 2836
rect 15628 2624 15668 2633
rect 15532 2584 15628 2624
rect 15340 2155 15380 2164
rect 15532 2204 15572 2213
rect 15436 1952 15476 2047
rect 15436 1903 15476 1912
rect 15532 1784 15572 2164
rect 15532 1735 15572 1744
rect 14860 139 14900 148
rect 15436 1700 15476 1709
rect 15436 80 15476 1660
rect 15628 1616 15668 2584
rect 15724 2540 15764 3088
rect 16012 3296 16052 3305
rect 15724 2491 15764 2500
rect 15820 2876 15860 2885
rect 15820 1952 15860 2836
rect 16012 2876 16052 3256
rect 16012 2708 16052 2836
rect 16012 2659 16052 2668
rect 16300 3212 16340 3221
rect 16204 2624 16244 2633
rect 16204 2489 16244 2584
rect 15820 1903 15860 1912
rect 16204 2036 16244 2045
rect 16204 1868 16244 1996
rect 16300 1952 16340 3172
rect 16396 2708 16436 2717
rect 16396 2372 16436 2668
rect 16396 2323 16436 2332
rect 16492 2120 16532 4432
rect 16684 4052 16724 7120
rect 16780 6992 16820 7001
rect 16972 6992 17012 11764
rect 17068 7916 17108 7925
rect 17068 7244 17108 7876
rect 17068 7195 17108 7204
rect 17164 7076 17204 11764
rect 17260 8504 17300 8513
rect 17260 8084 17300 8464
rect 17260 8035 17300 8044
rect 17164 7027 17204 7036
rect 16820 6952 17012 6992
rect 17068 6992 17108 7001
rect 16780 6943 16820 6952
rect 17068 5060 17108 6952
rect 17356 6656 17396 11764
rect 17548 9764 17588 11764
rect 17548 9715 17588 9724
rect 17644 10184 17684 10193
rect 17548 9512 17588 9521
rect 17452 9344 17492 9353
rect 17452 8000 17492 9304
rect 17452 7951 17492 7960
rect 17356 6607 17396 6616
rect 17452 7244 17492 7253
rect 17068 5011 17108 5020
rect 17260 6404 17300 6413
rect 17260 4892 17300 6364
rect 17356 5312 17396 5321
rect 17356 5060 17396 5272
rect 17356 5011 17396 5020
rect 17260 4556 17300 4852
rect 17260 4507 17300 4516
rect 16684 4003 16724 4012
rect 17452 3968 17492 7204
rect 16876 3212 16916 3221
rect 16876 2960 16916 3172
rect 16876 2911 16916 2920
rect 17260 2960 17300 2969
rect 17260 2900 17300 2920
rect 17452 2900 17492 3928
rect 17548 3884 17588 9472
rect 17644 7244 17684 10144
rect 17644 7195 17684 7204
rect 17740 6656 17780 11764
rect 17740 6607 17780 6616
rect 17836 9428 17876 9437
rect 17548 3835 17588 3844
rect 17644 6488 17684 6497
rect 17068 2876 17300 2900
rect 17108 2860 17300 2876
rect 17356 2860 17492 2900
rect 17068 2796 17108 2836
rect 16780 2708 16820 2717
rect 16492 2071 16532 2080
rect 16588 2456 16628 2465
rect 16300 1903 16340 1912
rect 16588 1952 16628 2416
rect 16780 2204 16820 2668
rect 16780 2155 16820 2164
rect 16972 2708 17012 2717
rect 16972 2204 17012 2668
rect 16972 2155 17012 2164
rect 17164 2120 17204 2129
rect 17068 2080 17164 2120
rect 16684 2036 16724 2045
rect 17068 2036 17108 2080
rect 17164 2071 17204 2080
rect 16724 1996 17108 2036
rect 16684 1987 16724 1996
rect 16588 1903 16628 1912
rect 16204 1819 16244 1828
rect 17356 1868 17396 2860
rect 17644 2792 17684 6448
rect 17836 5480 17876 9388
rect 17932 8168 17972 11764
rect 17932 8119 17972 8128
rect 18028 9596 18068 9605
rect 18028 8840 18068 9556
rect 18124 9596 18164 11764
rect 18220 10184 18260 10193
rect 18220 9848 18260 10144
rect 18220 9799 18260 9808
rect 18124 9547 18164 9556
rect 18028 7916 18068 8800
rect 18124 9260 18164 9269
rect 18124 8504 18164 9220
rect 18316 8924 18356 11764
rect 18412 10940 18452 10949
rect 18412 9260 18452 10900
rect 18412 9211 18452 9220
rect 18508 9176 18548 11764
rect 18604 10100 18644 10109
rect 18700 10100 18740 11764
rect 18644 10060 18740 10100
rect 18604 10051 18644 10060
rect 18892 10016 18932 11764
rect 18700 9976 18932 10016
rect 19084 10016 19124 11764
rect 19276 10184 19316 11764
rect 19276 10135 19316 10144
rect 19084 9976 19412 10016
rect 18508 9127 18548 9136
rect 18604 9260 18644 9269
rect 18124 8455 18164 8464
rect 18220 8884 18356 8924
rect 18412 8924 18452 8933
rect 18604 8924 18644 9220
rect 18028 7496 18068 7876
rect 18220 7832 18260 8884
rect 18220 7783 18260 7792
rect 18316 8672 18356 8681
rect 18028 7447 18068 7456
rect 18028 6488 18068 6497
rect 18028 6152 18068 6448
rect 18028 6103 18068 6112
rect 18124 6404 18164 6413
rect 17836 5431 17876 5440
rect 18124 5312 18164 6364
rect 18124 4556 18164 5272
rect 18028 4516 18164 4556
rect 18220 4724 18260 4733
rect 17932 4220 17972 4229
rect 17932 4052 17972 4180
rect 17932 3632 17972 4012
rect 17932 3583 17972 3592
rect 17644 2743 17684 2752
rect 17740 3212 17780 3221
rect 17356 1819 17396 1828
rect 16972 1784 17012 1793
rect 15628 1567 15668 1576
rect 16204 1700 16244 1709
rect 16204 80 16244 1660
rect 16972 80 17012 1744
rect 17740 80 17780 3172
rect 17932 2036 17972 2045
rect 17932 1901 17972 1996
rect 18028 1868 18068 4516
rect 18124 4304 18164 4313
rect 18124 1952 18164 4264
rect 18220 2708 18260 4684
rect 18220 2659 18260 2668
rect 18316 2624 18356 8632
rect 18412 7496 18452 8884
rect 18412 7447 18452 7456
rect 18508 8884 18644 8924
rect 18412 7244 18452 7253
rect 18412 6068 18452 7204
rect 18412 6019 18452 6028
rect 18412 5060 18452 5069
rect 18412 4808 18452 5020
rect 18412 4759 18452 4768
rect 18412 4304 18452 4313
rect 18412 3884 18452 4264
rect 18412 3835 18452 3844
rect 18508 2960 18548 8884
rect 18604 8756 18644 8765
rect 18604 8672 18644 8716
rect 18604 8621 18644 8632
rect 18604 8336 18644 8345
rect 18604 8168 18644 8296
rect 18604 8119 18644 8128
rect 18604 7328 18644 7337
rect 18604 5396 18644 7288
rect 18700 6656 18740 9976
rect 18808 9848 19176 9857
rect 18848 9808 18890 9848
rect 18930 9808 18972 9848
rect 19012 9808 19054 9848
rect 19094 9808 19136 9848
rect 18808 9799 19176 9808
rect 19276 9848 19316 9857
rect 19180 9512 19220 9521
rect 18796 9428 18836 9437
rect 18796 8924 18836 9388
rect 19180 9260 19220 9472
rect 19180 9211 19220 9220
rect 18796 8875 18836 8884
rect 18892 9092 18932 9101
rect 18796 8756 18836 8765
rect 18892 8756 18932 9052
rect 18836 8716 18932 8756
rect 18988 8840 19028 8851
rect 18988 8756 19028 8800
rect 19180 8840 19220 8849
rect 19276 8840 19316 9808
rect 19372 9764 19412 9976
rect 19372 9715 19412 9724
rect 19372 9344 19412 9353
rect 19468 9344 19508 11764
rect 19412 9304 19508 9344
rect 19564 10184 19604 10193
rect 19564 9344 19604 10144
rect 19372 9295 19412 9304
rect 19564 9295 19604 9304
rect 19220 8800 19316 8840
rect 19468 9092 19508 9101
rect 19180 8791 19220 8800
rect 18796 8707 18836 8716
rect 18988 8707 19028 8716
rect 19372 8672 19412 8681
rect 19276 8504 19316 8513
rect 18808 8336 19176 8345
rect 18848 8296 18890 8336
rect 18930 8296 18972 8336
rect 19012 8296 19054 8336
rect 19094 8296 19136 8336
rect 18808 8287 19176 8296
rect 19276 8336 19316 8464
rect 19276 8287 19316 8296
rect 18796 8000 18836 8009
rect 18796 7412 18836 7960
rect 19180 7580 19220 7589
rect 18796 7363 18836 7372
rect 18892 7328 18932 7423
rect 18892 7279 18932 7288
rect 18892 7160 18932 7169
rect 18892 7076 18932 7120
rect 18892 7025 18932 7036
rect 19180 6992 19220 7540
rect 19180 6943 19220 6952
rect 18808 6824 19176 6833
rect 18848 6784 18890 6824
rect 18930 6784 18972 6824
rect 19012 6784 19054 6824
rect 19094 6784 19136 6824
rect 18808 6775 19176 6784
rect 18700 6607 18740 6616
rect 19276 6740 19316 6749
rect 19180 6404 19220 6413
rect 19180 6152 19220 6364
rect 19180 6103 19220 6112
rect 18604 5347 18644 5356
rect 18700 5900 18740 5909
rect 18700 4808 18740 5860
rect 19276 5816 19316 6700
rect 19276 5767 19316 5776
rect 19276 5396 19316 5405
rect 18808 5312 19176 5321
rect 18848 5272 18890 5312
rect 18930 5272 18972 5312
rect 19012 5272 19054 5312
rect 19094 5272 19136 5312
rect 18808 5263 19176 5272
rect 19276 5312 19316 5356
rect 19276 5261 19316 5272
rect 18700 4759 18740 4768
rect 18796 4556 18836 4565
rect 18796 4220 18836 4516
rect 18796 4171 18836 4180
rect 19276 4052 19316 4061
rect 18604 3884 18644 3893
rect 18604 3548 18644 3844
rect 18808 3800 19176 3809
rect 18848 3760 18890 3800
rect 18930 3760 18972 3800
rect 19012 3760 19054 3800
rect 19094 3760 19136 3800
rect 18808 3751 19176 3760
rect 18604 3499 18644 3508
rect 18796 3632 18836 3641
rect 18796 3497 18836 3592
rect 18892 3380 18932 3389
rect 18508 2911 18548 2920
rect 18700 3296 18740 3305
rect 18700 2792 18740 3256
rect 18892 3044 18932 3340
rect 18892 2995 18932 3004
rect 18700 2743 18740 2752
rect 19276 2792 19316 4012
rect 19372 3296 19412 8632
rect 19468 7832 19508 9052
rect 19468 7328 19508 7792
rect 19468 7279 19508 7288
rect 19564 9092 19604 9101
rect 19468 6320 19508 6329
rect 19468 5060 19508 6280
rect 19564 5984 19604 9052
rect 19660 7580 19700 11764
rect 19852 10100 19892 11764
rect 19852 10051 19892 10060
rect 19948 11108 19988 11117
rect 19948 9596 19988 11068
rect 20044 9848 20084 11764
rect 20044 9799 20084 9808
rect 20140 10604 20180 10613
rect 19948 9547 19988 9556
rect 20044 9512 20084 9521
rect 19852 9428 19892 9437
rect 19756 9260 19796 9269
rect 19756 8756 19796 9220
rect 19852 9092 19892 9388
rect 19852 9043 19892 9052
rect 19948 9428 19988 9437
rect 19756 8707 19796 8716
rect 19948 8420 19988 9388
rect 20044 9260 20084 9472
rect 20140 9512 20180 10564
rect 20140 9463 20180 9472
rect 20236 9344 20276 11764
rect 20428 10100 20468 11764
rect 20428 10060 20564 10100
rect 20236 9295 20276 9304
rect 20044 9211 20084 9220
rect 20048 9092 20416 9101
rect 20088 9052 20130 9092
rect 20170 9052 20212 9092
rect 20252 9052 20294 9092
rect 20334 9052 20376 9092
rect 20048 9043 20416 9052
rect 20236 8924 20276 8933
rect 20236 8672 20276 8884
rect 20332 8924 20372 8933
rect 20524 8924 20564 10060
rect 20620 9680 20660 11764
rect 20620 9631 20660 9640
rect 20716 9596 20756 9605
rect 20372 8884 20564 8924
rect 20620 9176 20660 9185
rect 20332 8875 20372 8884
rect 20620 8840 20660 9136
rect 20524 8800 20660 8840
rect 20236 8537 20276 8632
rect 20332 8756 20372 8765
rect 20332 8588 20372 8716
rect 20332 8539 20372 8548
rect 20428 8672 20468 8681
rect 19948 8371 19988 8380
rect 20236 8420 20276 8429
rect 19948 8252 19988 8261
rect 19756 8084 19796 8095
rect 19756 8000 19796 8044
rect 19756 7951 19796 7960
rect 19948 7916 19988 8212
rect 20044 8084 20084 8093
rect 20044 7916 20084 8044
rect 20140 7916 20180 7925
rect 20044 7876 20140 7916
rect 19948 7867 19988 7876
rect 20140 7867 20180 7876
rect 19852 7748 19892 7757
rect 20236 7748 20276 8380
rect 20332 8420 20372 8429
rect 20332 8084 20372 8380
rect 20332 8035 20372 8044
rect 20428 7916 20468 8632
rect 20524 8672 20564 8800
rect 20524 8623 20564 8632
rect 20620 8420 20660 8429
rect 20428 7867 20468 7876
rect 20524 8084 20564 8093
rect 19756 7708 19852 7748
rect 19756 7664 19796 7708
rect 19852 7699 19892 7708
rect 19960 7708 20276 7748
rect 19960 7664 20000 7708
rect 19756 7615 19796 7624
rect 19948 7624 20000 7664
rect 19948 7580 19988 7624
rect 19660 7531 19700 7540
rect 19900 7540 19988 7580
rect 20048 7580 20416 7589
rect 20088 7540 20130 7580
rect 20170 7540 20212 7580
rect 20252 7540 20294 7580
rect 20334 7540 20376 7580
rect 19756 7412 19796 7421
rect 19900 7412 19940 7540
rect 20048 7531 20416 7540
rect 19900 7372 20000 7412
rect 19756 7244 19796 7372
rect 19960 7328 20000 7372
rect 19948 7288 20000 7328
rect 19756 7204 19892 7244
rect 19660 7160 19700 7169
rect 19660 6152 19700 7120
rect 19660 6103 19700 6112
rect 19756 7076 19796 7085
rect 19564 5944 19700 5984
rect 19468 5020 19604 5060
rect 19372 3247 19412 3256
rect 19468 3800 19508 3809
rect 19468 3128 19508 3760
rect 19276 2743 19316 2752
rect 19372 3088 19508 3128
rect 18316 2575 18356 2584
rect 18988 2708 19028 2717
rect 18988 2540 19028 2668
rect 18988 2491 19028 2500
rect 18508 2456 18548 2465
rect 18124 1903 18164 1912
rect 18412 2036 18452 2045
rect 18028 1819 18068 1828
rect 18412 1868 18452 1996
rect 18412 1819 18452 1828
rect 18508 80 18548 2416
rect 19276 2372 19316 2381
rect 18808 2288 19176 2297
rect 18848 2248 18890 2288
rect 18930 2248 18972 2288
rect 19012 2248 19054 2288
rect 19094 2248 19136 2288
rect 18808 2239 19176 2248
rect 19276 1952 19316 2332
rect 19276 1903 19316 1912
rect 19372 1868 19412 3088
rect 19468 2960 19508 2969
rect 19468 2708 19508 2920
rect 19468 2288 19508 2668
rect 19468 2239 19508 2248
rect 19372 1819 19412 1828
rect 19564 1700 19604 5020
rect 19660 1952 19700 5944
rect 19756 4472 19796 7036
rect 19852 7076 19892 7204
rect 19948 7160 19988 7288
rect 20524 7244 20564 8044
rect 20524 7195 20564 7204
rect 19948 7111 19988 7120
rect 19852 7027 19892 7036
rect 20140 7076 20180 7087
rect 20140 6992 20180 7036
rect 20140 6943 20180 6952
rect 20620 6656 20660 8380
rect 20716 7076 20756 9556
rect 20812 7160 20852 11764
rect 21004 10940 21044 11764
rect 21196 11108 21236 11764
rect 21196 11059 21236 11068
rect 21004 10891 21044 10900
rect 21004 10100 21044 10109
rect 20908 9428 20948 9437
rect 20908 9293 20948 9388
rect 20812 7111 20852 7120
rect 20908 8672 20948 8681
rect 20716 7027 20756 7036
rect 20908 6992 20948 8632
rect 20908 6943 20948 6952
rect 21004 6908 21044 10060
rect 21292 9932 21332 9941
rect 21292 9428 21332 9892
rect 21292 9379 21332 9388
rect 21292 9260 21332 9269
rect 21100 8840 21140 8880
rect 21100 8756 21140 8800
rect 21100 8336 21140 8716
rect 21100 7748 21140 8296
rect 21100 7699 21140 7708
rect 21196 8672 21236 8681
rect 21196 7580 21236 8632
rect 21004 6859 21044 6868
rect 21100 7540 21236 7580
rect 20620 6607 20660 6616
rect 19756 4423 19796 4432
rect 19948 6488 19988 6497
rect 19948 5648 19988 6448
rect 20716 6404 20756 6413
rect 20524 6236 20564 6245
rect 20048 6068 20416 6077
rect 20088 6028 20130 6068
rect 20170 6028 20212 6068
rect 20252 6028 20294 6068
rect 20334 6028 20376 6068
rect 20048 6019 20416 6028
rect 20044 5816 20084 5825
rect 20044 5732 20084 5776
rect 20044 5681 20084 5692
rect 19948 4976 19988 5608
rect 20524 5564 20564 6196
rect 20716 5732 20756 6364
rect 20812 5984 20852 5993
rect 20812 5849 20852 5944
rect 20716 5683 20756 5692
rect 21004 5732 21044 5741
rect 20524 5515 20564 5524
rect 19948 4136 19988 4936
rect 20524 4892 20564 4901
rect 20048 4556 20416 4565
rect 20088 4516 20130 4556
rect 20170 4516 20212 4556
rect 20252 4516 20294 4556
rect 20334 4516 20376 4556
rect 20048 4507 20416 4516
rect 20524 4304 20564 4852
rect 19948 4087 19988 4096
rect 20428 4264 20564 4304
rect 20908 4304 20948 4313
rect 20428 4136 20468 4264
rect 20140 4052 20180 4061
rect 20140 3917 20180 4012
rect 20428 3968 20468 4096
rect 20428 3919 20468 3928
rect 20524 4052 20564 4061
rect 20524 3464 20564 4012
rect 20908 3968 20948 4264
rect 19948 3212 19988 3221
rect 19948 2792 19988 3172
rect 20048 3044 20416 3053
rect 20088 3004 20130 3044
rect 20170 3004 20212 3044
rect 20252 3004 20294 3044
rect 20334 3004 20376 3044
rect 20048 2995 20416 3004
rect 20524 2900 20564 3424
rect 20812 3800 20852 3809
rect 20812 3380 20852 3760
rect 20812 3331 20852 3340
rect 20524 2860 20660 2900
rect 19948 2743 19988 2752
rect 20236 2792 20276 2801
rect 20044 2624 20084 2633
rect 19948 2540 19988 2549
rect 19948 2204 19988 2500
rect 20044 2288 20084 2584
rect 20044 2239 20084 2248
rect 19948 2155 19988 2164
rect 19756 1952 19796 1961
rect 19660 1912 19756 1952
rect 19756 1903 19796 1912
rect 20236 1952 20276 2752
rect 20236 1903 20276 1912
rect 20620 1868 20660 2860
rect 20716 2708 20756 2717
rect 20716 2120 20756 2668
rect 20716 2071 20756 2080
rect 20620 1819 20660 1828
rect 20908 1868 20948 3928
rect 21004 3464 21044 5692
rect 21004 2708 21044 3424
rect 21100 2876 21140 7540
rect 21292 7412 21332 9220
rect 21388 8084 21428 11764
rect 21580 10604 21620 11764
rect 21580 10555 21620 10564
rect 21484 10100 21524 10109
rect 21484 8924 21524 10060
rect 21676 10100 21716 10109
rect 21580 9680 21620 9689
rect 21580 9545 21620 9640
rect 21676 9596 21716 10060
rect 21676 9547 21716 9556
rect 21676 9428 21716 9437
rect 21484 8875 21524 8884
rect 21580 9176 21620 9185
rect 21388 8035 21428 8044
rect 21484 8420 21524 8429
rect 21196 7372 21332 7412
rect 21196 3632 21236 7372
rect 21292 7244 21332 7253
rect 21292 5564 21332 7204
rect 21292 5515 21332 5524
rect 21388 5732 21428 5741
rect 21388 4388 21428 5692
rect 21388 4339 21428 4348
rect 21196 3583 21236 3592
rect 21484 3296 21524 8380
rect 21580 7244 21620 9136
rect 21676 8672 21716 9388
rect 21676 8623 21716 8632
rect 21676 8504 21716 8513
rect 21676 7832 21716 8464
rect 21772 7916 21812 11764
rect 21868 9596 21908 9605
rect 21868 9176 21908 9556
rect 21868 9127 21908 9136
rect 21772 7867 21812 7876
rect 21868 8924 21908 8933
rect 21676 7783 21716 7792
rect 21580 7195 21620 7204
rect 21676 7496 21716 7505
rect 21580 6992 21620 7001
rect 21580 6908 21620 6952
rect 21580 6857 21620 6868
rect 21580 5816 21620 5825
rect 21580 5228 21620 5776
rect 21580 5179 21620 5188
rect 21484 3247 21524 3256
rect 21580 4808 21620 4817
rect 21100 2827 21140 2836
rect 21292 2876 21332 2885
rect 21004 2659 21044 2668
rect 21292 2372 21332 2836
rect 21580 2708 21620 4768
rect 21580 2659 21620 2668
rect 21292 2323 21332 2332
rect 21004 2120 21044 2129
rect 21004 1952 21044 2080
rect 21004 1903 21044 1912
rect 21676 1952 21716 7456
rect 21772 6908 21812 6917
rect 21772 6488 21812 6868
rect 21772 6439 21812 6448
rect 21868 2288 21908 8884
rect 21964 7328 22004 11764
rect 22060 9848 22100 9857
rect 22060 9680 22100 9808
rect 22060 9631 22100 9640
rect 22060 9092 22100 9101
rect 22060 8840 22100 9052
rect 22060 8791 22100 8800
rect 22060 8672 22100 8681
rect 22060 7832 22100 8632
rect 22156 8084 22196 11764
rect 22348 9932 22388 11764
rect 22156 8035 22196 8044
rect 22252 9892 22388 9932
rect 22252 8000 22292 9892
rect 22540 9680 22580 11764
rect 22732 10100 22772 11764
rect 22732 10051 22772 10060
rect 22540 9631 22580 9640
rect 22924 9428 22964 11764
rect 23116 9848 23156 11764
rect 23116 9799 23156 9808
rect 23212 10016 23252 10025
rect 23212 9596 23252 9976
rect 23308 9764 23348 11764
rect 23308 9715 23348 9724
rect 23404 10184 23444 10193
rect 23404 9680 23444 10144
rect 23404 9631 23444 9640
rect 23500 9680 23540 11764
rect 23500 9631 23540 9640
rect 23212 9547 23252 9556
rect 23692 9596 23732 11764
rect 23692 9547 23732 9556
rect 22924 9379 22964 9388
rect 23884 9428 23924 11764
rect 24076 9596 24116 11764
rect 24076 9547 24116 9556
rect 24268 9512 24308 11764
rect 24460 10688 24500 11764
rect 24460 10639 24500 10648
rect 24652 10100 24692 11764
rect 24652 10051 24692 10060
rect 24268 9463 24308 9472
rect 24748 9680 24788 9689
rect 23884 9379 23924 9388
rect 24556 9428 24596 9437
rect 22444 9344 22484 9353
rect 22348 9260 22388 9269
rect 22348 8924 22388 9220
rect 22444 9008 22484 9304
rect 22444 8959 22484 8968
rect 22636 9260 22676 9269
rect 22348 8875 22388 8884
rect 22252 7951 22292 7960
rect 22348 8756 22388 8765
rect 22252 7832 22292 7841
rect 22060 7792 22252 7832
rect 22252 7783 22292 7792
rect 21964 7279 22004 7288
rect 22156 7244 22196 7253
rect 21964 7160 22004 7169
rect 21964 3632 22004 7120
rect 22156 6488 22196 7204
rect 22156 6439 22196 6448
rect 22060 6404 22100 6413
rect 22060 5648 22100 6364
rect 22252 6404 22292 6413
rect 22252 6236 22292 6364
rect 22252 6187 22292 6196
rect 22060 5599 22100 5608
rect 22252 5396 22292 5405
rect 22252 4388 22292 5356
rect 22252 4339 22292 4348
rect 22348 4304 22388 8716
rect 22540 8336 22580 8345
rect 22444 8168 22484 8177
rect 22444 8033 22484 8128
rect 22444 7748 22484 7757
rect 22444 7412 22484 7708
rect 22444 7363 22484 7372
rect 22540 7244 22580 8296
rect 22540 6404 22580 7204
rect 22636 6740 22676 9220
rect 23692 9260 23732 9269
rect 23692 9092 23732 9220
rect 23692 9043 23732 9052
rect 23884 9260 23924 9269
rect 23212 8924 23252 8933
rect 22828 8756 22868 8765
rect 22732 8420 22772 8429
rect 22732 8285 22772 8380
rect 22828 8000 22868 8716
rect 22636 6691 22676 6700
rect 22732 7960 22868 8000
rect 23212 8000 23252 8884
rect 23788 8756 23828 8765
rect 23788 8504 23828 8716
rect 23788 8455 23828 8464
rect 22732 7160 22772 7960
rect 23212 7951 23252 7960
rect 23404 8084 23444 8093
rect 23404 8000 23444 8044
rect 23404 7949 23444 7960
rect 23788 7916 23828 7925
rect 22540 6355 22580 6364
rect 22732 5816 22772 7120
rect 22732 5767 22772 5776
rect 22828 7832 22868 7841
rect 22828 7160 22868 7792
rect 23020 7328 23060 7337
rect 22828 5816 22868 7120
rect 22924 7288 23020 7328
rect 22924 6656 22964 7288
rect 23020 7260 23060 7288
rect 23596 7328 23636 7337
rect 23212 7076 23252 7171
rect 23212 7027 23252 7036
rect 23404 6992 23444 7001
rect 22924 6607 22964 6616
rect 23212 6656 23252 6665
rect 23020 6572 23060 6581
rect 23060 6532 23156 6572
rect 23020 6523 23060 6532
rect 22924 5984 22964 5995
rect 22924 5900 22964 5944
rect 22924 5851 22964 5860
rect 23116 5900 23156 6532
rect 23212 6152 23252 6616
rect 23212 6103 23252 6112
rect 23404 6068 23444 6952
rect 23596 6404 23636 7288
rect 23788 7160 23828 7876
rect 23596 6152 23636 6364
rect 23596 6103 23636 6112
rect 23692 6992 23732 7001
rect 23404 6019 23444 6028
rect 23116 5851 23156 5860
rect 23404 5900 23444 5909
rect 22540 5732 22580 5741
rect 22444 5648 22484 5657
rect 22444 4892 22484 5608
rect 22540 5312 22580 5692
rect 22540 5263 22580 5272
rect 22444 4843 22484 4852
rect 22636 4892 22676 4901
rect 22348 4255 22388 4264
rect 22060 4136 22100 4145
rect 22252 4136 22292 4145
rect 22100 4096 22252 4136
rect 22060 4087 22100 4096
rect 22252 4087 22292 4096
rect 22636 3884 22676 4852
rect 22636 3835 22676 3844
rect 21964 3583 22004 3592
rect 21868 2239 21908 2248
rect 22252 2288 22292 2297
rect 21676 1903 21716 1912
rect 20908 1819 20948 1828
rect 21772 1868 21812 1877
rect 19564 1651 19604 1660
rect 19852 1784 19892 1793
rect 19276 1616 19316 1625
rect 19276 80 19316 1576
rect 19852 188 19892 1744
rect 19948 1700 19988 1709
rect 19948 860 19988 1660
rect 21580 1700 21620 1709
rect 20524 1616 20564 1627
rect 20048 1532 20416 1541
rect 20088 1492 20130 1532
rect 20170 1492 20212 1532
rect 20252 1492 20294 1532
rect 20334 1492 20376 1532
rect 20048 1483 20416 1492
rect 20524 1532 20564 1576
rect 20524 1483 20564 1492
rect 19948 811 19988 820
rect 20812 860 20852 869
rect 19852 148 20084 188
rect 20044 80 20084 148
rect 20812 80 20852 820
rect 21580 80 21620 1660
rect 21772 1616 21812 1828
rect 22252 1868 22292 2248
rect 22732 2288 22772 2297
rect 22732 2153 22772 2248
rect 22636 2120 22676 2129
rect 22636 2036 22676 2080
rect 22828 2120 22868 5776
rect 23020 5816 23060 5825
rect 23020 5648 23060 5776
rect 23404 5732 23444 5860
rect 23404 5683 23444 5692
rect 23020 5599 23060 5608
rect 23692 5648 23732 6952
rect 23692 5599 23732 5608
rect 23212 5396 23252 5405
rect 22924 4892 22964 4901
rect 22924 4640 22964 4852
rect 22924 4591 22964 4600
rect 23116 4472 23156 4481
rect 23116 4052 23156 4432
rect 23116 4003 23156 4012
rect 23020 3296 23060 3305
rect 22924 3256 23020 3296
rect 22924 3128 22964 3256
rect 23020 3228 23060 3256
rect 22924 3079 22964 3088
rect 23212 3044 23252 5356
rect 23596 5144 23636 5153
rect 23596 4556 23636 5104
rect 23692 4976 23732 4985
rect 23692 4841 23732 4936
rect 23788 4892 23828 7120
rect 23788 4843 23828 4852
rect 23596 4507 23636 4516
rect 23788 4388 23828 4397
rect 23500 4304 23540 4313
rect 23500 4136 23540 4264
rect 23788 4253 23828 4348
rect 23500 4087 23540 4096
rect 23692 4136 23732 4145
rect 23020 3004 23252 3044
rect 23020 2792 23060 3004
rect 22924 2752 23060 2792
rect 22924 2708 22964 2752
rect 22924 2659 22964 2668
rect 23212 2708 23252 2717
rect 23212 2456 23252 2668
rect 22924 2372 22964 2381
rect 22924 2204 22964 2332
rect 23212 2288 23252 2416
rect 23212 2239 23252 2248
rect 23596 2708 23636 2717
rect 23020 2204 23060 2213
rect 22924 2164 23020 2204
rect 23020 2136 23060 2164
rect 22828 2071 22868 2080
rect 22636 1985 22676 1996
rect 22252 1819 22292 1828
rect 23500 1952 23540 1961
rect 21772 1567 21812 1576
rect 22348 1700 22388 1709
rect 22348 80 22388 1660
rect 23116 1700 23156 1709
rect 23116 80 23156 1660
rect 23308 1532 23348 1541
rect 23308 1397 23348 1492
rect 23500 1532 23540 1912
rect 23596 1784 23636 2668
rect 23692 2036 23732 4096
rect 23884 2708 23924 9220
rect 24460 9260 24500 9269
rect 24172 9008 24212 9017
rect 24172 8672 24212 8968
rect 24460 8756 24500 9220
rect 24460 8707 24500 8716
rect 24364 8672 24404 8681
rect 24172 8632 24364 8672
rect 24364 8623 24404 8632
rect 24076 8588 24116 8597
rect 23980 5060 24020 5069
rect 23980 4556 24020 5020
rect 24076 4892 24116 8548
rect 24460 8588 24500 8597
rect 24268 8504 24308 8513
rect 24268 8369 24308 8464
rect 24172 7832 24212 7841
rect 24172 5396 24212 7792
rect 24364 6992 24404 7001
rect 24268 6572 24308 6581
rect 24268 5732 24308 6532
rect 24268 5683 24308 5692
rect 24172 5347 24212 5356
rect 24076 4843 24116 4852
rect 24172 5060 24212 5069
rect 23980 4507 24020 4516
rect 24076 4724 24116 4733
rect 23884 2659 23924 2668
rect 23980 4052 24020 4061
rect 23692 1868 23732 1996
rect 23692 1819 23732 1828
rect 23980 1868 24020 4012
rect 24076 3380 24116 4684
rect 24172 4388 24212 5020
rect 24268 4976 24308 5071
rect 24268 4927 24308 4936
rect 24172 4339 24212 4348
rect 24268 4808 24308 4817
rect 24268 4388 24308 4768
rect 24268 4339 24308 4348
rect 24364 4388 24404 6952
rect 24364 4339 24404 4348
rect 24268 3380 24308 3389
rect 24076 3331 24116 3340
rect 24172 3340 24268 3380
rect 24076 2624 24116 2633
rect 24172 2624 24212 3340
rect 24268 3331 24308 3340
rect 24460 3380 24500 8548
rect 24556 8504 24596 9388
rect 24748 9428 24788 9640
rect 24844 9596 24884 11764
rect 24844 9547 24884 9556
rect 24748 9379 24788 9388
rect 24940 9344 24980 9353
rect 24844 8924 24884 8933
rect 24556 8455 24596 8464
rect 24652 8756 24692 8765
rect 24652 7748 24692 8716
rect 24652 7244 24692 7708
rect 24652 7195 24692 7204
rect 24556 6488 24596 6497
rect 24556 5480 24596 6448
rect 24556 5431 24596 5440
rect 24556 4892 24596 4901
rect 24556 4136 24596 4852
rect 24556 4087 24596 4096
rect 24748 3716 24788 3725
rect 24748 3464 24788 3676
rect 24844 3632 24884 8884
rect 24940 8840 24980 9304
rect 24940 8672 24980 8800
rect 24940 8623 24980 8632
rect 25036 7160 25076 11764
rect 25228 10856 25268 11764
rect 25228 10807 25268 10816
rect 25228 10688 25268 10697
rect 25132 9680 25172 9689
rect 25132 8672 25172 9640
rect 25228 9512 25268 10648
rect 25228 9463 25268 9472
rect 25132 8623 25172 8632
rect 25036 7111 25076 7120
rect 25324 7160 25364 7169
rect 25132 7076 25172 7085
rect 25132 6488 25172 7036
rect 25324 6908 25364 7120
rect 25420 7076 25460 11764
rect 25612 10604 25652 11764
rect 25612 10555 25652 10564
rect 25804 10352 25844 11764
rect 25996 10940 26036 11764
rect 25996 10891 26036 10900
rect 25804 10303 25844 10312
rect 25804 10100 25844 10109
rect 25804 9512 25844 10060
rect 25804 9463 25844 9472
rect 25900 9260 25940 9269
rect 25612 8756 25652 8765
rect 25612 8621 25652 8716
rect 25708 8168 25748 8177
rect 25748 8128 25844 8168
rect 25708 8119 25748 8128
rect 25804 7916 25844 8128
rect 25804 7867 25844 7876
rect 25420 7027 25460 7036
rect 25612 7328 25652 7337
rect 25324 6859 25364 6868
rect 25324 6488 25364 6497
rect 25132 6448 25324 6488
rect 25132 5648 25172 6448
rect 25324 6439 25364 6448
rect 24940 4304 24980 4315
rect 24940 4220 24980 4264
rect 24940 4171 24980 4180
rect 25132 4220 25172 5608
rect 25612 5564 25652 7288
rect 25900 7244 25940 9220
rect 26092 9260 26132 9269
rect 26092 9125 26132 9220
rect 26188 9008 26228 11764
rect 26380 11192 26420 11764
rect 26380 11143 26420 11152
rect 26188 8959 26228 8968
rect 26284 9260 26324 9269
rect 26092 8756 26132 8765
rect 26092 8168 26132 8716
rect 26092 8119 26132 8128
rect 26188 8084 26228 8093
rect 26284 8084 26324 9220
rect 26476 8924 26516 8933
rect 26476 8588 26516 8884
rect 26572 8672 26612 11764
rect 26764 11360 26804 11764
rect 26764 11311 26804 11320
rect 26572 8623 26612 8632
rect 26476 8539 26516 8548
rect 26380 8084 26420 8112
rect 26228 8044 26380 8084
rect 26188 8035 26228 8044
rect 26380 8035 26420 8044
rect 25900 7195 25940 7204
rect 25996 7832 26036 7841
rect 25900 6992 25940 7001
rect 25996 6992 26036 7792
rect 26956 7160 26996 11764
rect 27148 10100 27188 11764
rect 27148 10051 27188 10060
rect 27052 9764 27092 9773
rect 27052 9428 27092 9724
rect 27052 8756 27092 9388
rect 27340 9428 27380 11764
rect 27532 9596 27572 11764
rect 27724 10688 27764 11764
rect 27724 10648 27860 10688
rect 27724 10352 27764 10361
rect 27532 9547 27572 9556
rect 27628 10100 27668 10109
rect 27340 9379 27380 9388
rect 27436 9428 27476 9437
rect 27340 9260 27380 9269
rect 27340 9008 27380 9220
rect 27340 8959 27380 8968
rect 27052 8707 27092 8716
rect 27244 8840 27284 8849
rect 27244 8705 27284 8800
rect 27436 8840 27476 9388
rect 27628 9428 27668 10060
rect 27628 9379 27668 9388
rect 27436 8791 27476 8800
rect 27436 8672 27476 8681
rect 27724 8672 27764 10312
rect 27820 9932 27860 10648
rect 27820 9883 27860 9892
rect 27820 9260 27860 9269
rect 27820 9176 27860 9220
rect 27820 9125 27860 9136
rect 27820 8672 27860 8681
rect 27724 8632 27820 8672
rect 27340 7832 27380 7841
rect 26956 7111 26996 7120
rect 27148 7328 27188 7337
rect 27148 7244 27188 7288
rect 27340 7328 27380 7792
rect 27340 7279 27380 7288
rect 25940 6952 26036 6992
rect 27052 6992 27092 7001
rect 25900 6404 25940 6952
rect 25900 6355 25940 6364
rect 26572 6908 26612 6917
rect 25900 6236 25940 6245
rect 25708 5900 25748 5909
rect 25708 5648 25748 5860
rect 25708 5599 25748 5608
rect 25612 5515 25652 5524
rect 25132 4171 25172 4180
rect 25324 4220 25364 4229
rect 24844 3583 24884 3592
rect 25132 3632 25172 3641
rect 24748 3415 24788 3424
rect 24460 3331 24500 3340
rect 24364 3296 24404 3305
rect 24364 2792 24404 3256
rect 25132 3044 25172 3592
rect 25228 3548 25268 3559
rect 25228 3464 25268 3508
rect 25228 3415 25268 3424
rect 25132 2995 25172 3004
rect 25228 2960 25268 2969
rect 24116 2584 24212 2624
rect 24268 2708 24308 2717
rect 24076 2575 24116 2584
rect 24268 2372 24308 2668
rect 24268 2323 24308 2332
rect 23980 1819 24020 1828
rect 24364 1868 24404 2752
rect 24940 2876 25172 2900
rect 24940 2860 25132 2876
rect 24556 2708 24596 2717
rect 24556 2573 24596 2668
rect 24940 2456 24980 2860
rect 25132 2827 25172 2836
rect 24844 2416 24980 2456
rect 25036 2792 25076 2801
rect 24844 2372 24884 2416
rect 24844 2323 24884 2332
rect 24940 2288 24980 2297
rect 24364 1819 24404 1828
rect 24748 1952 24788 1961
rect 23596 1735 23636 1744
rect 24076 1784 24116 1793
rect 23500 1483 23540 1492
rect 23884 1700 23924 1709
rect 23884 80 23924 1660
rect 24076 1616 24116 1744
rect 24076 1567 24116 1576
rect 24652 1784 24692 1793
rect 24652 80 24692 1744
rect 24748 1700 24788 1912
rect 24748 1651 24788 1660
rect 24940 1616 24980 2248
rect 25036 2120 25076 2752
rect 25132 2288 25172 2299
rect 25132 2204 25172 2248
rect 25132 2155 25172 2164
rect 25036 2071 25076 2080
rect 25228 2036 25268 2920
rect 25324 2792 25364 4180
rect 25708 3968 25748 3977
rect 25324 2743 25364 2752
rect 25420 3212 25460 3221
rect 25228 1987 25268 1996
rect 24940 1567 24980 1576
rect 25420 80 25460 3172
rect 25516 2708 25556 2717
rect 25516 2372 25556 2668
rect 25708 2708 25748 3928
rect 25708 2659 25748 2668
rect 25804 2960 25844 2969
rect 25516 2323 25556 2332
rect 25804 1952 25844 2920
rect 25900 2036 25940 6196
rect 25996 5732 26036 5741
rect 25996 4976 26036 5692
rect 25996 3380 26036 4936
rect 26188 5648 26228 5657
rect 26188 4472 26228 5608
rect 26188 4423 26228 4432
rect 25996 3331 26036 3340
rect 26380 3380 26420 3389
rect 26380 3245 26420 3340
rect 26572 2792 26612 6868
rect 26764 6908 26804 6917
rect 26668 6824 26708 6833
rect 26668 6656 26708 6784
rect 26668 6607 26708 6616
rect 26764 6068 26804 6868
rect 27052 6656 27092 6952
rect 27052 6607 27092 6616
rect 27148 6488 27188 7204
rect 27340 7076 27380 7085
rect 27340 6572 27380 7036
rect 27340 6523 27380 6532
rect 27188 6448 27284 6488
rect 27148 6439 27188 6448
rect 26764 6019 26804 6028
rect 27052 4976 27092 4985
rect 27052 4808 27092 4936
rect 27052 4759 27092 4768
rect 27148 4892 27188 4901
rect 26572 2743 26612 2752
rect 26284 2708 26324 2717
rect 25996 2540 26036 2549
rect 25996 2120 26036 2500
rect 25996 2071 26036 2080
rect 26188 2540 26228 2549
rect 25900 1987 25940 1996
rect 25804 1903 25844 1912
rect 26188 80 26228 2500
rect 26284 1532 26324 2668
rect 27148 1868 27188 4852
rect 27244 4220 27284 6448
rect 27244 4171 27284 4180
rect 27340 6320 27380 6329
rect 27340 2900 27380 6280
rect 27436 2960 27476 8632
rect 27820 8623 27860 8632
rect 27532 8504 27572 8513
rect 27532 7160 27572 8464
rect 27532 7111 27572 7120
rect 27628 7580 27668 7589
rect 27532 5732 27572 5741
rect 27532 5312 27572 5692
rect 27532 5263 27572 5272
rect 27436 2911 27476 2920
rect 27244 2860 27380 2900
rect 27244 2624 27284 2860
rect 27244 2575 27284 2584
rect 27532 2708 27572 2717
rect 27532 2573 27572 2668
rect 27148 1819 27188 1828
rect 26284 1483 26324 1492
rect 26956 1700 26996 1709
rect 26956 80 26996 1660
rect 27628 1532 27668 7540
rect 27724 7580 27764 7589
rect 27724 7328 27764 7540
rect 27724 7279 27764 7288
rect 27916 6488 27956 11764
rect 28108 10100 28148 11764
rect 28300 11024 28340 11764
rect 28300 10975 28340 10984
rect 28300 10856 28340 10865
rect 28108 10060 28244 10100
rect 28108 9008 28148 9017
rect 28108 8672 28148 8968
rect 28108 8623 28148 8632
rect 28204 8168 28244 10060
rect 28300 9512 28340 10816
rect 28300 9463 28340 9472
rect 28204 8119 28244 8128
rect 28300 9176 28340 9185
rect 28108 8084 28148 8093
rect 28108 6572 28148 8044
rect 28108 6523 28148 6532
rect 27916 6439 27956 6448
rect 28300 6236 28340 9136
rect 28396 9092 28436 9101
rect 28396 8840 28436 9052
rect 28396 8791 28436 8800
rect 28492 8084 28532 11764
rect 28684 10772 28724 11764
rect 28876 11108 28916 11764
rect 28876 11068 29012 11108
rect 28684 10723 28724 10732
rect 28876 10940 28916 10949
rect 28684 10604 28724 10613
rect 28588 9848 28628 9857
rect 28588 9713 28628 9808
rect 28684 9512 28724 10564
rect 28684 9463 28724 9472
rect 28876 9512 28916 10900
rect 28876 9463 28916 9472
rect 28780 9260 28820 9269
rect 28588 9092 28628 9103
rect 28588 9008 28628 9052
rect 28588 8959 28628 8968
rect 28684 8672 28724 8681
rect 28684 8537 28724 8632
rect 28492 8035 28532 8044
rect 28588 8504 28628 8513
rect 28588 7916 28628 8464
rect 28780 8336 28820 9220
rect 28972 8588 29012 11068
rect 29068 10100 29108 11764
rect 29068 10060 29204 10100
rect 29068 9680 29108 9689
rect 29068 9545 29108 9640
rect 29068 9344 29108 9353
rect 29068 8672 29108 9304
rect 29068 8623 29108 8632
rect 28972 8539 29012 8548
rect 29164 8588 29204 10060
rect 29260 8672 29300 11764
rect 29452 11360 29492 11764
rect 29356 11320 29492 11360
rect 29356 10100 29396 11320
rect 29356 10051 29396 10060
rect 29452 11192 29492 11201
rect 29452 9512 29492 11152
rect 29644 10772 29684 11764
rect 29836 11528 29876 11764
rect 30028 11612 30068 11764
rect 29836 11479 29876 11488
rect 29932 11572 30068 11612
rect 29644 10723 29684 10732
rect 29836 11360 29876 11369
rect 29452 9463 29492 9472
rect 29548 10100 29588 10109
rect 29548 9344 29588 10060
rect 29644 9932 29684 9941
rect 29644 9797 29684 9892
rect 29836 9512 29876 11320
rect 29836 9463 29876 9472
rect 29932 9344 29972 11572
rect 29548 9295 29588 9304
rect 29836 9304 29972 9344
rect 30028 11444 30068 11453
rect 29260 8623 29300 8632
rect 29356 8756 29396 8765
rect 29164 8539 29204 8548
rect 29356 8504 29396 8716
rect 28780 8287 28820 8296
rect 29260 8464 29396 8504
rect 29644 8588 29684 8597
rect 28588 7867 28628 7876
rect 28396 7748 28436 7757
rect 28396 7580 28436 7708
rect 28396 7531 28436 7540
rect 29068 7580 29108 7589
rect 29068 7328 29108 7540
rect 29068 7244 29108 7288
rect 29068 7193 29108 7204
rect 28876 6572 28916 6581
rect 28780 6488 28820 6497
rect 28300 6187 28340 6196
rect 28396 6448 28780 6488
rect 27820 3212 27860 3221
rect 27820 2708 27860 3172
rect 28396 2900 28436 6448
rect 28780 6439 28820 6448
rect 28684 6320 28724 6329
rect 28588 4892 28628 4901
rect 27820 2659 27860 2668
rect 28300 2860 28436 2900
rect 28492 4556 28532 4565
rect 28300 2624 28340 2860
rect 28300 2575 28340 2584
rect 27628 1483 27668 1492
rect 27820 1868 27860 1877
rect 27820 1532 27860 1828
rect 27820 1483 27860 1492
rect 27724 104 27764 113
rect 3128 0 3208 80
rect 3896 0 3976 80
rect 4664 0 4744 80
rect 5432 0 5512 80
rect 6200 0 6280 80
rect 6968 0 7048 80
rect 7736 0 7816 80
rect 8504 0 8584 80
rect 9272 0 9352 80
rect 10040 0 10120 80
rect 10808 0 10888 80
rect 11576 0 11656 80
rect 12344 0 12424 80
rect 13112 0 13192 80
rect 13880 0 13960 80
rect 14648 0 14728 80
rect 15416 0 15496 80
rect 16184 0 16264 80
rect 16952 0 17032 80
rect 17720 0 17800 80
rect 18488 0 18568 80
rect 19256 0 19336 80
rect 20024 0 20104 80
rect 20792 0 20872 80
rect 21560 0 21640 80
rect 22328 0 22408 80
rect 23096 0 23176 80
rect 23864 0 23944 80
rect 24632 0 24712 80
rect 25400 0 25480 80
rect 26168 0 26248 80
rect 26936 0 27016 80
rect 27704 64 27724 80
rect 28492 80 28532 4516
rect 28588 4136 28628 4852
rect 28588 4087 28628 4096
rect 28684 3548 28724 6280
rect 28684 3499 28724 3508
rect 28780 6068 28820 6077
rect 28780 2708 28820 6028
rect 28876 5984 28916 6532
rect 28876 5935 28916 5944
rect 28972 6404 29012 6413
rect 28972 5984 29012 6364
rect 28972 5935 29012 5944
rect 29260 5900 29300 8464
rect 29356 7916 29396 7925
rect 29356 7412 29396 7876
rect 29356 7363 29396 7372
rect 29548 7244 29588 7253
rect 29548 6404 29588 7204
rect 29644 7160 29684 8548
rect 29740 8588 29780 8597
rect 29740 7916 29780 8548
rect 29740 7867 29780 7876
rect 29644 7111 29684 7120
rect 29740 7076 29780 7171
rect 29740 7027 29780 7036
rect 29548 6355 29588 6364
rect 29644 6992 29684 7001
rect 29164 5860 29300 5900
rect 29644 5900 29684 6952
rect 29836 6908 29876 9304
rect 29932 8588 29972 8597
rect 29932 8252 29972 8548
rect 29932 8203 29972 8212
rect 29836 6859 29876 6868
rect 29932 7748 29972 7757
rect 29740 6824 29780 6833
rect 29740 6689 29780 6784
rect 29836 6740 29876 6749
rect 29836 6572 29876 6700
rect 29836 6523 29876 6532
rect 28876 5648 28916 5657
rect 28876 4976 28916 5608
rect 28876 4927 28916 4936
rect 28972 5480 29012 5489
rect 28972 5144 29012 5440
rect 28972 4976 29012 5104
rect 28972 4927 29012 4936
rect 29164 4892 29204 5860
rect 29644 5851 29684 5860
rect 29836 6152 29876 6161
rect 29260 5732 29300 5741
rect 29260 5228 29300 5692
rect 29260 5179 29300 5188
rect 29452 5648 29492 5657
rect 29068 4724 29108 4733
rect 28876 4304 28916 4313
rect 28876 4220 28916 4264
rect 28876 4169 28916 4180
rect 28972 3968 29012 3977
rect 28876 3380 28916 3389
rect 28876 2876 28916 3340
rect 28876 2827 28916 2836
rect 28780 2659 28820 2668
rect 28684 2624 28724 2633
rect 28684 1868 28724 2584
rect 28684 1819 28724 1828
rect 28780 2288 28820 2297
rect 28780 1784 28820 2248
rect 28972 1868 29012 3928
rect 29068 3044 29108 4684
rect 29164 4136 29204 4852
rect 29260 4724 29300 4733
rect 29260 4304 29300 4684
rect 29452 4724 29492 5608
rect 29740 4976 29780 4985
rect 29740 4841 29780 4936
rect 29452 4675 29492 4684
rect 29260 4255 29300 4264
rect 29164 4087 29204 4096
rect 29740 3968 29780 3977
rect 29644 3800 29684 3809
rect 29260 3716 29300 3725
rect 29068 2995 29108 3004
rect 29164 3380 29204 3389
rect 29164 2708 29204 3340
rect 29260 2960 29300 3676
rect 29548 3632 29588 3641
rect 29548 3464 29588 3592
rect 29644 3632 29684 3760
rect 29644 3583 29684 3592
rect 29548 3415 29588 3424
rect 29260 2911 29300 2920
rect 29356 3296 29396 3305
rect 29164 2659 29204 2668
rect 28972 1819 29012 1828
rect 29260 2624 29300 2633
rect 29260 1868 29300 2584
rect 29260 1819 29300 1828
rect 28780 1735 28820 1744
rect 29356 1784 29396 3256
rect 29452 2876 29492 2885
rect 29452 2120 29492 2836
rect 29740 2708 29780 3928
rect 29740 2372 29780 2668
rect 29836 2456 29876 6112
rect 29932 3380 29972 7708
rect 30028 7076 30068 11404
rect 30220 10016 30260 11764
rect 30412 10688 30452 11764
rect 30412 10639 30452 10648
rect 30604 10268 30644 11764
rect 30604 10219 30644 10228
rect 30220 9967 30260 9976
rect 30700 9596 30740 9605
rect 30700 9461 30740 9556
rect 30124 9428 30164 9437
rect 30124 9293 30164 9388
rect 30220 9344 30260 9353
rect 30028 7027 30068 7036
rect 30124 9008 30164 9017
rect 30028 6908 30068 6917
rect 30028 6773 30068 6868
rect 30124 5984 30164 8968
rect 30220 8504 30260 9304
rect 30412 9344 30452 9353
rect 30220 8455 30260 8464
rect 30316 9260 30356 9269
rect 30220 8084 30260 8093
rect 30220 7949 30260 8044
rect 30316 6824 30356 9220
rect 30412 8756 30452 9304
rect 30412 8707 30452 8716
rect 30604 9260 30644 9269
rect 30316 6775 30356 6784
rect 30412 7160 30452 7169
rect 29932 3331 29972 3340
rect 30028 5944 30164 5984
rect 29836 2407 29876 2416
rect 29740 2323 29780 2332
rect 29452 2071 29492 2080
rect 29548 2204 29588 2213
rect 29356 1735 29396 1744
rect 29548 1784 29588 2164
rect 29548 1735 29588 1744
rect 29260 188 29300 197
rect 29260 80 29300 148
rect 30028 80 30068 5944
rect 30220 5480 30260 5489
rect 30124 5396 30164 5405
rect 30124 4724 30164 5356
rect 30124 4675 30164 4684
rect 30124 4556 30164 4565
rect 30124 2792 30164 4516
rect 30220 3968 30260 5440
rect 30220 3919 30260 3928
rect 30220 3548 30260 3557
rect 30220 3464 30260 3508
rect 30220 3413 30260 3424
rect 30412 3380 30452 7120
rect 30604 3716 30644 9220
rect 30796 8252 30836 11764
rect 30892 10100 30932 10109
rect 30988 10100 31028 11764
rect 30988 10060 31124 10100
rect 30892 8840 30932 10060
rect 30892 8791 30932 8800
rect 30988 8672 31028 8681
rect 30988 8537 31028 8632
rect 30796 8203 30836 8212
rect 31084 8168 31124 10060
rect 31084 8119 31124 8128
rect 31084 7328 31124 7337
rect 31084 4304 31124 7288
rect 31180 5396 31220 11764
rect 31372 10184 31412 11764
rect 31372 10135 31412 10144
rect 31468 9932 31508 9941
rect 31468 9596 31508 9892
rect 31468 9547 31508 9556
rect 31276 9260 31316 9269
rect 31276 6488 31316 9220
rect 31468 8756 31508 8765
rect 31372 7916 31412 7925
rect 31372 7664 31412 7876
rect 31372 7615 31412 7624
rect 31468 7328 31508 8716
rect 31276 6439 31316 6448
rect 31372 7288 31508 7328
rect 31180 5347 31220 5356
rect 31372 6404 31412 7288
rect 31468 6908 31508 6917
rect 31468 6488 31508 6868
rect 31468 6439 31508 6448
rect 31372 5144 31412 6364
rect 31564 5984 31604 11764
rect 31660 11024 31700 11033
rect 31660 9596 31700 10984
rect 31756 10100 31796 11764
rect 31756 10051 31796 10060
rect 31660 9547 31700 9556
rect 31852 10016 31892 10025
rect 31756 9260 31796 9269
rect 31564 5935 31604 5944
rect 31660 7832 31700 7841
rect 31660 7244 31700 7792
rect 31660 5228 31700 7204
rect 31756 6152 31796 9220
rect 31852 7328 31892 9976
rect 31852 7279 31892 7288
rect 31756 6103 31796 6112
rect 31852 6992 31892 7001
rect 31852 5900 31892 6952
rect 31852 5851 31892 5860
rect 31756 5816 31796 5825
rect 31756 5564 31796 5776
rect 31756 5515 31796 5524
rect 31948 5312 31988 11764
rect 32140 9764 32180 11764
rect 32332 11276 32372 11764
rect 32332 11227 32372 11236
rect 32140 9715 32180 9724
rect 32332 10772 32372 10781
rect 32332 9512 32372 10732
rect 32332 9463 32372 9472
rect 32428 9428 32468 9439
rect 32428 9344 32468 9388
rect 32428 9295 32468 9304
rect 32044 9260 32084 9269
rect 32044 6656 32084 9220
rect 32140 8756 32180 8765
rect 32140 7916 32180 8716
rect 32524 8336 32564 11764
rect 32716 11192 32756 11764
rect 32716 11143 32756 11152
rect 32716 9512 32756 9521
rect 32524 8287 32564 8296
rect 32620 9472 32716 9512
rect 32620 8168 32660 9472
rect 32716 9463 32756 9472
rect 32812 9428 32852 9437
rect 32524 8128 32660 8168
rect 32716 8252 32756 8261
rect 32140 7867 32180 7876
rect 32236 7916 32276 7925
rect 32140 7244 32180 7253
rect 32140 6740 32180 7204
rect 32236 6992 32276 7876
rect 32236 6943 32276 6952
rect 32140 6700 32276 6740
rect 32044 6616 32180 6656
rect 31948 5263 31988 5272
rect 32044 6404 32084 6413
rect 31660 5179 31700 5188
rect 31372 5095 31412 5104
rect 31084 4255 31124 4264
rect 31660 4640 31700 4649
rect 30604 3667 30644 3676
rect 31660 3380 31700 4600
rect 31948 4220 31988 4229
rect 31852 3884 31892 3893
rect 31852 3749 31892 3844
rect 31948 3548 31988 4180
rect 31948 3499 31988 3508
rect 31852 3380 31892 3389
rect 31660 3340 31852 3380
rect 30412 3331 30452 3340
rect 31852 3331 31892 3340
rect 30124 2743 30164 2752
rect 31180 3296 31220 3305
rect 31180 3128 31220 3256
rect 31180 2708 31220 3088
rect 31180 2659 31220 2668
rect 32044 2708 32084 6364
rect 32140 4220 32180 6616
rect 32236 6404 32276 6700
rect 32236 6355 32276 6364
rect 32428 5060 32468 5069
rect 32140 4171 32180 4180
rect 32236 4388 32276 4397
rect 32140 3968 32180 3977
rect 32140 3464 32180 3928
rect 32140 3415 32180 3424
rect 30412 2624 30452 2633
rect 30412 2036 30452 2584
rect 30412 1987 30452 1996
rect 30700 2624 30740 2633
rect 30700 1868 30740 2584
rect 31852 2624 31892 2633
rect 30700 1819 30740 1828
rect 31372 2540 31412 2549
rect 31372 1952 31412 2500
rect 30124 1784 30164 1793
rect 30124 1532 30164 1744
rect 30124 1483 30164 1492
rect 31372 1364 31412 1912
rect 31372 1315 31412 1324
rect 31564 2372 31604 2381
rect 30796 1028 30836 1037
rect 30796 80 30836 988
rect 31564 80 31604 2332
rect 31852 2372 31892 2584
rect 32044 2540 32084 2668
rect 32044 2491 32084 2500
rect 32236 2540 32276 4348
rect 32332 3884 32372 3893
rect 32332 3749 32372 3844
rect 32236 2491 32276 2500
rect 32332 2792 32372 2801
rect 31852 1952 31892 2332
rect 31852 1903 31892 1912
rect 32140 1952 32180 1961
rect 32140 1817 32180 1912
rect 32332 80 32372 2752
rect 32428 1532 32468 5020
rect 32524 4976 32564 8128
rect 32716 8000 32756 8212
rect 32716 7951 32756 7960
rect 32812 7916 32852 9388
rect 32908 8420 32948 11764
rect 33100 11444 33140 11764
rect 33100 11404 33236 11444
rect 33196 9260 33236 11404
rect 33196 9211 33236 9220
rect 33196 9092 33236 9101
rect 33004 9008 33044 9017
rect 33004 8873 33044 8968
rect 33196 8840 33236 9052
rect 33292 8924 33332 11764
rect 33388 9848 33428 9857
rect 33388 9092 33428 9808
rect 33484 9680 33524 11764
rect 33484 9631 33524 9640
rect 33388 9043 33428 9052
rect 33292 8884 33428 8924
rect 33196 8791 33236 8800
rect 33292 8756 33332 8765
rect 33196 8672 33236 8681
rect 32908 8371 32948 8380
rect 33004 8588 33044 8597
rect 33004 8420 33044 8548
rect 33004 8371 33044 8380
rect 32620 7580 32660 7589
rect 32620 7076 32660 7540
rect 32620 7027 32660 7036
rect 32716 7160 32756 7169
rect 32716 6908 32756 7120
rect 32812 7076 32852 7876
rect 33100 7412 33140 7421
rect 33100 7277 33140 7372
rect 32812 7027 32852 7036
rect 32908 7076 32948 7085
rect 32716 6859 32756 6868
rect 32620 6824 32660 6833
rect 32620 6572 32660 6784
rect 32620 6523 32660 6532
rect 32716 6740 32756 6749
rect 32716 6572 32756 6700
rect 32716 6523 32756 6532
rect 32812 6656 32852 6665
rect 32812 6488 32852 6616
rect 32812 6439 32852 6448
rect 32908 5648 32948 7036
rect 33004 6992 33044 7001
rect 33196 6992 33236 8632
rect 33292 8168 33332 8716
rect 33388 8672 33428 8884
rect 33388 8623 33428 8632
rect 33484 8840 33524 8849
rect 33292 8119 33332 8128
rect 33388 8504 33428 8513
rect 33292 7832 33332 7841
rect 33292 7160 33332 7792
rect 33292 7111 33332 7120
rect 33388 7076 33428 8464
rect 33388 7027 33428 7036
rect 33196 6952 33332 6992
rect 33004 6320 33044 6952
rect 33004 6271 33044 6280
rect 32908 5599 32948 5608
rect 33196 5648 33236 5657
rect 33004 5564 33044 5573
rect 32812 5480 32852 5489
rect 32524 4927 32564 4936
rect 32716 5396 32756 5405
rect 32620 4892 32660 4901
rect 32620 4304 32660 4852
rect 32620 4255 32660 4264
rect 32524 3968 32564 3977
rect 32524 3800 32564 3928
rect 32524 3751 32564 3760
rect 32716 1616 32756 5356
rect 32812 5312 32852 5440
rect 33004 5396 33044 5524
rect 33004 5347 33044 5356
rect 32812 5263 32852 5272
rect 33196 5144 33236 5608
rect 33196 5095 33236 5104
rect 33100 5060 33140 5069
rect 32812 4976 32852 4985
rect 32812 4220 32852 4936
rect 33100 4925 33140 5020
rect 33292 4892 33332 6952
rect 33484 6656 33524 8800
rect 33580 8756 33620 8765
rect 33580 7748 33620 8716
rect 33580 7412 33620 7708
rect 33580 7363 33620 7372
rect 33676 7244 33716 11764
rect 33868 10016 33908 11764
rect 33868 9967 33908 9976
rect 34060 10016 34100 11764
rect 34252 10016 34292 11764
rect 34444 10352 34484 11764
rect 34444 10303 34484 10312
rect 34540 10772 34580 10781
rect 34252 9976 34388 10016
rect 34060 9967 34100 9976
rect 33772 9932 33812 9941
rect 33772 9797 33812 9892
rect 33928 9848 34296 9857
rect 33968 9808 34010 9848
rect 34050 9808 34092 9848
rect 34132 9808 34174 9848
rect 34214 9808 34256 9848
rect 33928 9799 34296 9808
rect 33676 7195 33716 7204
rect 33772 9596 33812 9605
rect 33676 7076 33716 7085
rect 33580 6908 33620 6917
rect 33580 6773 33620 6868
rect 33484 6616 33620 6656
rect 33292 4843 33332 4852
rect 33388 6152 33428 6161
rect 33196 4808 33236 4817
rect 32908 4472 32948 4481
rect 32908 4337 32948 4432
rect 33100 4304 33140 4313
rect 32812 4171 32852 4180
rect 33004 4264 33100 4304
rect 33004 4136 33044 4264
rect 33100 4255 33140 4264
rect 33004 4087 33044 4096
rect 32812 3296 32852 3305
rect 32812 2708 32852 3256
rect 33100 3296 33140 3305
rect 33196 3296 33236 4768
rect 33292 4640 33332 4649
rect 33292 4388 33332 4600
rect 33292 4220 33332 4348
rect 33292 4171 33332 4180
rect 33388 4136 33428 6112
rect 33484 5564 33524 5573
rect 33484 4808 33524 5524
rect 33484 4759 33524 4768
rect 33388 3464 33428 4096
rect 33292 3424 33428 3464
rect 33292 3380 33332 3424
rect 33292 3331 33332 3340
rect 33140 3256 33236 3296
rect 33100 3228 33140 3256
rect 33196 2900 33236 3256
rect 33100 2876 33236 2900
rect 33140 2860 33236 2876
rect 33580 2900 33620 6616
rect 33676 6320 33716 7036
rect 33676 6271 33716 6280
rect 33676 5732 33716 5741
rect 33676 4976 33716 5692
rect 33676 4927 33716 4936
rect 33676 4808 33716 4817
rect 33676 4673 33716 4768
rect 33676 3296 33716 3305
rect 33676 3161 33716 3256
rect 33580 2860 33716 2900
rect 33100 2827 33140 2836
rect 32812 2659 32852 2668
rect 33388 2624 33428 2633
rect 33388 2372 33428 2584
rect 33388 2323 33428 2332
rect 33580 2540 33620 2549
rect 32716 1567 32756 1576
rect 33580 1616 33620 2500
rect 33676 1784 33716 2860
rect 33772 2204 33812 9556
rect 33868 9512 33908 9521
rect 33868 9008 33908 9472
rect 33868 8959 33908 8968
rect 34156 9260 34196 9269
rect 33868 8840 33908 8849
rect 34060 8840 34100 8849
rect 33908 8800 34060 8840
rect 33868 8791 33908 8800
rect 34060 8791 34100 8800
rect 34156 8756 34196 9220
rect 34156 8707 34196 8716
rect 33928 8336 34296 8345
rect 33968 8296 34010 8336
rect 34050 8296 34092 8336
rect 34132 8296 34174 8336
rect 34214 8296 34256 8336
rect 33928 8287 34296 8296
rect 34060 8168 34100 8177
rect 33964 7412 34004 7421
rect 33964 7244 34004 7372
rect 33964 7195 34004 7204
rect 33868 7076 33908 7171
rect 34060 7160 34100 8128
rect 34252 8168 34292 8177
rect 34060 7111 34100 7120
rect 34156 7916 34196 7925
rect 34156 7580 34196 7876
rect 34252 7664 34292 8128
rect 34348 8084 34388 9976
rect 34444 9680 34484 9689
rect 34444 9176 34484 9640
rect 34540 9512 34580 10732
rect 34540 9463 34580 9472
rect 34444 9127 34484 9136
rect 34540 9344 34580 9353
rect 34444 9008 34484 9017
rect 34444 8168 34484 8968
rect 34540 8840 34580 9304
rect 34636 8924 34676 11764
rect 34828 9260 34868 11764
rect 34828 9211 34868 9220
rect 34924 10268 34964 10277
rect 34636 8875 34676 8884
rect 34828 9092 34868 9101
rect 34540 8791 34580 8800
rect 34732 8252 34772 8261
rect 34444 8128 34580 8168
rect 34348 8044 34484 8084
rect 34252 7615 34292 7624
rect 34156 7160 34196 7540
rect 34348 7328 34388 7337
rect 34348 7193 34388 7288
rect 34156 7111 34196 7120
rect 33868 7027 33908 7036
rect 33928 6824 34296 6833
rect 33968 6784 34010 6824
rect 34050 6784 34092 6824
rect 34132 6784 34174 6824
rect 34214 6784 34256 6824
rect 33928 6775 34296 6784
rect 34444 6824 34484 8044
rect 34540 7328 34580 8128
rect 34732 8084 34772 8212
rect 34732 8035 34772 8044
rect 34828 7328 34868 9052
rect 34924 8672 34964 10228
rect 34924 8623 34964 8632
rect 34924 8420 34964 8429
rect 34924 8252 34964 8380
rect 34924 8203 34964 8212
rect 34924 7916 34964 7925
rect 34924 7580 34964 7876
rect 34924 7531 34964 7540
rect 34540 7288 34772 7328
rect 34540 7160 34580 7169
rect 34540 6908 34580 7120
rect 34732 7160 34772 7288
rect 34636 6908 34676 6917
rect 34540 6868 34636 6908
rect 34636 6859 34676 6868
rect 34444 6775 34484 6784
rect 33964 6656 34004 6665
rect 33964 5732 34004 6616
rect 34348 6572 34388 6581
rect 33964 5683 34004 5692
rect 34060 6320 34100 6329
rect 33868 5648 33908 5657
rect 33868 5480 33908 5608
rect 34060 5648 34100 6280
rect 34060 5599 34100 5608
rect 33868 5431 33908 5440
rect 33928 5312 34296 5321
rect 33968 5272 34010 5312
rect 34050 5272 34092 5312
rect 34132 5272 34174 5312
rect 34214 5272 34256 5312
rect 33928 5263 34296 5272
rect 34348 4976 34388 6532
rect 34732 6404 34772 7120
rect 34828 6656 34868 7288
rect 34828 6607 34868 6616
rect 34924 6488 34964 6497
rect 34828 6404 34868 6413
rect 34732 6364 34828 6404
rect 34828 6355 34868 6364
rect 34636 6320 34676 6329
rect 34636 5732 34676 6280
rect 34636 5683 34676 5692
rect 34828 5816 34868 5825
rect 34828 5732 34868 5776
rect 34828 5681 34868 5692
rect 34348 4927 34388 4936
rect 34444 5480 34484 5489
rect 33868 4892 33908 4901
rect 33868 4220 33908 4852
rect 33868 4171 33908 4180
rect 34348 4220 34388 4229
rect 33928 3800 34296 3809
rect 33968 3760 34010 3800
rect 34050 3760 34092 3800
rect 34132 3760 34174 3800
rect 34214 3760 34256 3800
rect 33928 3751 34296 3760
rect 34348 2876 34388 4180
rect 34348 2827 34388 2836
rect 34444 2624 34484 5440
rect 34540 5144 34580 5153
rect 34540 4052 34580 5104
rect 34732 5060 34772 5069
rect 34924 5060 34964 6448
rect 35020 5900 35060 11764
rect 37228 11276 37268 11285
rect 35980 10688 36020 10697
rect 35788 9932 35828 9941
rect 35596 9596 35636 9605
rect 35308 9344 35348 9439
rect 35308 9295 35348 9304
rect 35168 9092 35536 9101
rect 35208 9052 35250 9092
rect 35290 9052 35332 9092
rect 35372 9052 35414 9092
rect 35454 9052 35496 9092
rect 35168 9043 35536 9052
rect 35212 8420 35252 8429
rect 35212 8336 35252 8380
rect 35212 8285 35252 8296
rect 35116 8252 35156 8263
rect 35116 8168 35156 8212
rect 35116 8119 35156 8128
rect 35168 7580 35536 7589
rect 35208 7540 35250 7580
rect 35290 7540 35332 7580
rect 35372 7540 35414 7580
rect 35454 7540 35496 7580
rect 35168 7531 35536 7540
rect 35596 7076 35636 9556
rect 35596 7027 35636 7036
rect 35692 8924 35732 8933
rect 35596 6572 35636 6581
rect 35168 6068 35536 6077
rect 35208 6028 35250 6068
rect 35290 6028 35332 6068
rect 35372 6028 35414 6068
rect 35454 6028 35496 6068
rect 35168 6019 35536 6028
rect 35020 5860 35156 5900
rect 35020 5732 35060 5743
rect 35020 5648 35060 5692
rect 35020 5599 35060 5608
rect 35116 5480 35156 5860
rect 35596 5648 35636 6532
rect 35692 6320 35732 8884
rect 35788 8672 35828 9892
rect 35980 9596 36020 10648
rect 35980 9547 36020 9556
rect 36172 10184 36212 10193
rect 36172 9596 36212 10144
rect 36172 9547 36212 9556
rect 36460 10100 36500 10109
rect 36460 9596 36500 10060
rect 36652 10100 36692 10109
rect 36652 9932 36692 10060
rect 36652 9883 36692 9892
rect 37228 9680 37268 11236
rect 37228 9631 37268 9640
rect 37516 11192 37556 11201
rect 36460 9547 36500 9556
rect 37228 9512 37268 9521
rect 35980 9428 36020 9437
rect 35788 8623 35828 8632
rect 35884 9260 35924 9269
rect 35692 6271 35732 6280
rect 35788 7832 35828 7841
rect 35788 6572 35828 7792
rect 35788 6320 35828 6532
rect 35788 6271 35828 6280
rect 35596 5599 35636 5608
rect 35116 5431 35156 5440
rect 34732 4136 34772 5020
rect 34732 4087 34772 4096
rect 34828 5020 34964 5060
rect 35116 5228 35156 5237
rect 35116 5060 35156 5188
rect 34636 4052 34676 4061
rect 34540 4012 34636 4052
rect 34636 4003 34676 4012
rect 34828 3464 34868 5020
rect 35116 5011 35156 5020
rect 34924 4892 34964 4901
rect 34924 4304 34964 4852
rect 35692 4640 35732 4649
rect 35168 4556 35536 4565
rect 35208 4516 35250 4556
rect 35290 4516 35332 4556
rect 35372 4516 35414 4556
rect 35454 4516 35496 4556
rect 35168 4507 35536 4516
rect 34924 4255 34964 4264
rect 35596 3968 35636 3977
rect 35404 3800 35444 3809
rect 34828 2900 34868 3424
rect 35020 3548 35060 3557
rect 35020 3044 35060 3508
rect 35404 3212 35444 3760
rect 35404 3163 35444 3172
rect 35596 3128 35636 3928
rect 35596 3079 35636 3088
rect 35020 2995 35060 3004
rect 35168 3044 35536 3053
rect 35208 3004 35250 3044
rect 35290 3004 35332 3044
rect 35372 3004 35414 3044
rect 35454 3004 35496 3044
rect 35168 2995 35536 3004
rect 34828 2860 35156 2900
rect 33928 2288 34296 2297
rect 33968 2248 34010 2288
rect 34050 2248 34092 2288
rect 34132 2248 34174 2288
rect 34214 2248 34256 2288
rect 33928 2239 34296 2248
rect 33772 2155 33812 2164
rect 34060 2120 34100 2129
rect 34444 2120 34484 2584
rect 34924 2708 34964 2717
rect 34100 2080 34484 2120
rect 34828 2204 34868 2213
rect 34060 2071 34100 2080
rect 33676 1735 33716 1744
rect 34252 1952 34292 1961
rect 33580 1567 33620 1576
rect 32428 1483 32468 1492
rect 33100 104 33140 113
rect 27764 64 27784 80
rect 27704 0 27784 64
rect 28472 0 28552 80
rect 29240 0 29320 80
rect 30008 0 30088 80
rect 30776 0 30856 80
rect 31544 0 31624 80
rect 32312 0 32392 80
rect 33080 64 33100 80
rect 33868 104 33908 113
rect 33140 64 33160 80
rect 33080 0 33160 64
rect 33848 64 33868 80
rect 34060 104 34100 113
rect 33908 64 33928 80
rect 33848 0 33928 64
rect 34060 60 34100 64
rect 34252 60 34292 1912
rect 34348 1700 34388 2080
rect 34348 1651 34388 1660
rect 34444 1784 34484 1793
rect 34444 1649 34484 1744
rect 34636 1784 34676 1793
rect 34636 80 34676 1744
rect 34828 1448 34868 2164
rect 34924 2120 34964 2668
rect 35116 2708 35156 2860
rect 35116 2659 35156 2668
rect 35500 2792 35540 2801
rect 35500 2657 35540 2752
rect 34924 2071 34964 2080
rect 35692 1952 35732 4600
rect 35884 3464 35924 9220
rect 35980 8924 36020 9388
rect 36940 9176 36980 9185
rect 36172 8924 36212 8933
rect 35980 8875 36020 8884
rect 36076 8884 36172 8924
rect 35980 8756 36020 8765
rect 36076 8756 36116 8884
rect 36172 8875 36212 8884
rect 36020 8716 36116 8756
rect 35980 8707 36020 8716
rect 35980 8504 36020 8513
rect 35980 8168 36020 8464
rect 35980 8119 36020 8128
rect 36268 8420 36308 8429
rect 35980 7832 36020 7841
rect 35980 7697 36020 7792
rect 36076 7748 36116 7757
rect 36076 7328 36116 7708
rect 36268 7496 36308 8380
rect 36268 7447 36308 7456
rect 36364 8000 36404 8009
rect 36364 7412 36404 7960
rect 36748 8000 36788 8009
rect 36748 7580 36788 7960
rect 36748 7531 36788 7540
rect 36364 7363 36404 7372
rect 36076 7279 36116 7288
rect 35980 7244 36020 7253
rect 35980 6656 36020 7204
rect 35980 6607 36020 6616
rect 36748 7160 36788 7169
rect 36364 6572 36404 6581
rect 35980 6404 36020 6413
rect 36020 6364 36116 6404
rect 35980 6355 36020 6364
rect 35980 5480 36020 5489
rect 35980 5345 36020 5440
rect 36076 5144 36116 6364
rect 36364 6068 36404 6532
rect 36748 6404 36788 7120
rect 36940 7160 36980 9136
rect 36940 7111 36980 7120
rect 37036 7244 37076 7253
rect 36844 6992 36884 7001
rect 36844 6740 36884 6952
rect 36844 6691 36884 6700
rect 37036 6656 37076 7204
rect 37036 6607 37076 6616
rect 36748 6355 36788 6364
rect 37132 6404 37172 6413
rect 36364 6019 36404 6028
rect 36556 5900 36596 5909
rect 36460 5648 36500 5657
rect 36172 5564 36212 5573
rect 36172 5396 36212 5524
rect 36460 5513 36500 5608
rect 36172 5347 36212 5356
rect 36076 5095 36116 5104
rect 36556 5144 36596 5860
rect 36556 5095 36596 5104
rect 37132 4220 37172 6364
rect 35884 3415 35924 3424
rect 36172 4136 36212 4145
rect 35788 3380 35828 3389
rect 35788 3044 35828 3340
rect 35788 2995 35828 3004
rect 36172 3380 36212 4096
rect 36076 2792 36116 2801
rect 36076 2204 36116 2752
rect 36172 2540 36212 3340
rect 36172 2491 36212 2500
rect 36940 3716 36980 3725
rect 36076 2155 36116 2164
rect 35692 1903 35732 1912
rect 36172 1952 36212 1961
rect 35596 1868 35636 1877
rect 35168 1532 35536 1541
rect 35208 1492 35250 1532
rect 35290 1492 35332 1532
rect 35372 1492 35414 1532
rect 35454 1492 35496 1532
rect 35168 1483 35536 1492
rect 34828 1399 34868 1408
rect 35596 188 35636 1828
rect 35404 148 35636 188
rect 35404 80 35444 148
rect 36172 80 36212 1912
rect 36940 80 36980 3676
rect 37132 2708 37172 4180
rect 37132 2659 37172 2668
rect 37228 2204 37268 9472
rect 37420 9428 37460 9437
rect 37324 8756 37364 8765
rect 37324 8084 37364 8716
rect 37420 8168 37460 9388
rect 37516 9260 37556 11152
rect 44716 11024 44756 11033
rect 44236 10688 44276 10697
rect 39148 10352 39188 10361
rect 37900 10016 37940 10025
rect 37708 9512 37748 9521
rect 37516 9211 37556 9220
rect 37612 9472 37708 9512
rect 37420 8119 37460 8128
rect 37516 8756 37556 8765
rect 37324 8035 37364 8044
rect 37324 6992 37364 7001
rect 37324 6908 37364 6952
rect 37324 6857 37364 6868
rect 37420 6572 37460 6581
rect 37420 5648 37460 6532
rect 37420 5599 37460 5608
rect 37516 4136 37556 8716
rect 37516 4087 37556 4096
rect 37324 3464 37364 3473
rect 37516 3464 37556 3473
rect 37364 3424 37516 3464
rect 37324 3415 37364 3424
rect 37516 3415 37556 3424
rect 37324 2708 37364 2717
rect 37324 2372 37364 2668
rect 37324 2323 37364 2332
rect 37228 2155 37268 2164
rect 37612 2204 37652 9472
rect 37708 9463 37748 9472
rect 37804 9260 37844 9269
rect 37804 9125 37844 9220
rect 37900 8756 37940 9976
rect 38668 10016 38708 10025
rect 38188 9932 38228 9941
rect 38188 9428 38228 9892
rect 38668 9512 38708 9976
rect 38764 10016 38804 10025
rect 38764 9680 38804 9976
rect 38764 9631 38804 9640
rect 39052 9848 39092 9857
rect 38668 9463 38708 9472
rect 39052 9512 39092 9808
rect 39148 9680 39188 10312
rect 43276 10352 43316 10361
rect 41452 10100 41492 10109
rect 39148 9631 39188 9640
rect 41068 9932 41108 9941
rect 39052 9463 39092 9472
rect 39340 9596 39380 9605
rect 38188 9379 38228 9388
rect 38764 9344 38804 9353
rect 38956 9344 38996 9353
rect 38804 9304 38956 9344
rect 38764 9295 38804 9304
rect 38956 9295 38996 9304
rect 38188 9260 38228 9269
rect 37996 9220 38188 9260
rect 37996 9092 38036 9220
rect 38188 9211 38228 9220
rect 39340 9176 39380 9556
rect 39340 9127 39380 9136
rect 39628 9428 39668 9437
rect 39244 9092 39284 9101
rect 37996 9043 38036 9052
rect 38860 9052 39244 9092
rect 37900 8707 37940 8716
rect 38860 8756 38900 9052
rect 39244 9043 39284 9052
rect 38860 8707 38900 8716
rect 39628 8756 39668 9388
rect 40204 9260 40244 9269
rect 39628 8707 39668 8716
rect 40012 8756 40052 8765
rect 37804 8672 37844 8681
rect 37708 7832 37748 7841
rect 37708 7160 37748 7792
rect 37708 7111 37748 7120
rect 37612 2155 37652 2164
rect 37804 2120 37844 8632
rect 38764 8672 38804 8681
rect 38380 8504 38420 8513
rect 37900 7412 37940 7421
rect 37900 7328 37940 7372
rect 37900 7277 37940 7288
rect 38092 7076 38132 7085
rect 37900 6320 37940 6329
rect 37900 4976 37940 6280
rect 37900 3296 37940 4936
rect 37996 5648 38036 5657
rect 37996 4808 38036 5608
rect 37996 4220 38036 4768
rect 37996 4171 38036 4180
rect 37900 3247 37940 3256
rect 37900 2876 37940 2885
rect 37900 2792 37940 2836
rect 37900 2741 37940 2752
rect 37804 2071 37844 2080
rect 37900 2204 37940 2213
rect 37900 2069 37940 2164
rect 38092 2120 38132 7036
rect 38188 6404 38228 6413
rect 38188 6269 38228 6364
rect 38092 2071 38132 2080
rect 38188 4556 38228 4565
rect 37708 1952 37748 1961
rect 37708 80 37748 1912
rect 38188 188 38228 4516
rect 38380 3296 38420 8464
rect 38764 8000 38804 8632
rect 39148 8672 39188 8681
rect 38764 7951 38804 7960
rect 38860 8588 38900 8597
rect 38668 7916 38708 7925
rect 38668 7160 38708 7876
rect 38668 7111 38708 7120
rect 38860 5648 38900 8548
rect 39148 8084 39188 8632
rect 39148 8035 39188 8044
rect 39820 7916 39860 7925
rect 38956 7748 38996 7757
rect 38956 6404 38996 7708
rect 38956 6355 38996 6364
rect 39244 7748 39284 7757
rect 38860 5599 38900 5608
rect 38956 5732 38996 5741
rect 38572 5480 38612 5489
rect 38572 4892 38612 5440
rect 38956 4976 38996 5692
rect 38956 4927 38996 4936
rect 38572 4843 38612 4852
rect 38764 4724 38804 4733
rect 38572 4304 38612 4313
rect 38476 4052 38516 4061
rect 38476 3917 38516 4012
rect 38572 3464 38612 4264
rect 38764 4304 38804 4684
rect 39244 4472 39284 7708
rect 39436 7664 39476 7673
rect 39436 7244 39476 7624
rect 39436 5732 39476 7204
rect 39628 6404 39668 6413
rect 39628 6152 39668 6364
rect 39628 5816 39668 6112
rect 39628 5767 39668 5776
rect 39436 5683 39476 5692
rect 39820 5732 39860 7876
rect 39820 5683 39860 5692
rect 39916 7328 39956 7337
rect 39244 4423 39284 4432
rect 39436 4892 39476 4901
rect 38764 4255 38804 4264
rect 38956 4304 38996 4399
rect 38956 4255 38996 4264
rect 39148 4304 39188 4313
rect 39148 4220 39188 4264
rect 39052 4180 39188 4220
rect 39340 4220 39380 4229
rect 39052 4136 39092 4180
rect 39340 4136 39380 4180
rect 38572 3415 38612 3424
rect 38764 4096 39092 4136
rect 39148 4096 39380 4136
rect 38380 3247 38420 3256
rect 38668 3296 38708 3305
rect 38668 2708 38708 3256
rect 38668 2659 38708 2668
rect 38764 2792 38804 4096
rect 39148 3212 39188 4096
rect 39436 4052 39476 4852
rect 39916 4472 39956 7288
rect 39436 4003 39476 4012
rect 39532 4136 39572 4147
rect 39532 4052 39572 4096
rect 39532 4003 39572 4012
rect 39628 3968 39668 3977
rect 39148 3163 39188 3172
rect 39244 3464 39284 3473
rect 38668 2456 38708 2465
rect 38668 2288 38708 2416
rect 38668 2239 38708 2248
rect 38764 1700 38804 2752
rect 38956 2792 38996 2801
rect 39148 2792 39188 2801
rect 38996 2752 39148 2792
rect 38956 2743 38996 2752
rect 39148 2743 39188 2752
rect 38956 2624 38996 2633
rect 38764 1651 38804 1660
rect 38860 2540 38900 2549
rect 38668 1616 38708 1627
rect 38668 1532 38708 1576
rect 38668 1483 38708 1492
rect 38188 148 38516 188
rect 38476 80 38516 148
rect 38860 104 38900 2500
rect 38956 2456 38996 2584
rect 38956 2407 38996 2416
rect 39052 2372 39092 2381
rect 38956 1616 38996 1625
rect 38956 1532 38996 1576
rect 38956 1481 38996 1492
rect 39052 1028 39092 2332
rect 39052 979 39092 988
rect 34060 20 34292 60
rect 34616 0 34696 80
rect 35384 0 35464 80
rect 36152 0 36232 80
rect 36920 0 37000 80
rect 37688 0 37768 80
rect 38456 0 38536 80
rect 39244 80 39284 3424
rect 39628 3128 39668 3928
rect 39628 3079 39668 3088
rect 39820 3212 39860 3221
rect 39820 3077 39860 3172
rect 39916 2960 39956 4432
rect 39340 2456 39380 2465
rect 39340 188 39380 2416
rect 39916 1952 39956 2920
rect 39916 1903 39956 1912
rect 39340 139 39380 148
rect 40012 80 40052 8716
rect 40204 8336 40244 9220
rect 40492 9176 40532 9185
rect 40300 9092 40340 9101
rect 40300 8957 40340 9052
rect 40204 8287 40244 8296
rect 40396 8672 40436 8681
rect 40396 8252 40436 8632
rect 40396 8203 40436 8212
rect 40108 7328 40148 7337
rect 40108 6404 40148 7288
rect 40108 6355 40148 6364
rect 40396 6236 40436 6245
rect 40300 5732 40340 5741
rect 40300 4976 40340 5692
rect 40300 4304 40340 4936
rect 40204 3968 40244 3977
rect 40204 3380 40244 3928
rect 40204 3331 40244 3340
rect 40204 3212 40244 3221
rect 40204 2960 40244 3172
rect 40204 2911 40244 2920
rect 40300 2456 40340 4264
rect 40300 2407 40340 2416
rect 40300 2288 40340 2297
rect 40300 2153 40340 2248
rect 40396 1784 40436 6196
rect 40492 2120 40532 9136
rect 40780 9008 40820 9017
rect 40780 8672 40820 8968
rect 40684 8000 40724 8009
rect 40684 7244 40724 7960
rect 40780 7748 40820 8632
rect 40780 7699 40820 7708
rect 40588 6404 40628 6413
rect 40588 5480 40628 6364
rect 40684 5732 40724 7204
rect 40972 7580 41012 7589
rect 40876 6320 40916 6329
rect 40684 5683 40724 5692
rect 40780 5816 40820 5825
rect 40588 5431 40628 5440
rect 40588 4976 40628 4985
rect 40588 4388 40628 4936
rect 40588 4339 40628 4348
rect 40684 3632 40724 3641
rect 40684 3380 40724 3592
rect 40684 3331 40724 3340
rect 40492 2071 40532 2080
rect 40396 1735 40436 1744
rect 40780 80 40820 5776
rect 40876 4808 40916 6280
rect 40876 1700 40916 4768
rect 40972 2120 41012 7540
rect 41068 4892 41108 9892
rect 41356 9428 41396 9437
rect 41260 8840 41300 8849
rect 41164 8504 41204 8513
rect 41164 4976 41204 8464
rect 41260 7916 41300 8800
rect 41260 7867 41300 7876
rect 41260 6992 41300 7001
rect 41260 6404 41300 6952
rect 41260 6355 41300 6364
rect 41260 4976 41300 4985
rect 41164 4936 41260 4976
rect 41260 4927 41300 4936
rect 41068 4852 41204 4892
rect 41164 4808 41204 4852
rect 41164 4768 41300 4808
rect 40972 2071 41012 2080
rect 41068 4724 41108 4733
rect 41068 1868 41108 4684
rect 41068 1819 41108 1828
rect 41164 4640 41204 4649
rect 40876 1651 40916 1660
rect 38860 55 38900 64
rect 39224 0 39304 80
rect 39992 0 40072 80
rect 40760 0 40840 80
rect 41164 60 41204 4600
rect 41260 2876 41300 4768
rect 41260 2827 41300 2836
rect 41260 2288 41300 2297
rect 41356 2288 41396 9388
rect 41452 8000 41492 10060
rect 42220 10016 42260 10025
rect 41452 7951 41492 7960
rect 41548 9932 41588 9941
rect 41300 2248 41396 2288
rect 41452 7412 41492 7421
rect 41452 2288 41492 7372
rect 41548 4640 41588 9892
rect 42028 9344 42068 9353
rect 41740 9260 41780 9269
rect 41740 8924 41780 9220
rect 41780 8884 41876 8924
rect 41740 8875 41780 8884
rect 41740 8588 41780 8597
rect 41740 8000 41780 8548
rect 41740 7951 41780 7960
rect 41836 7412 41876 8884
rect 41836 7363 41876 7372
rect 41932 6992 41972 7001
rect 41740 6236 41780 6245
rect 41740 6101 41780 6196
rect 41932 5984 41972 6952
rect 42028 6656 42068 9304
rect 42028 6607 42068 6616
rect 41932 5935 41972 5944
rect 42124 6404 42164 6413
rect 42124 5900 42164 6364
rect 42124 5851 42164 5860
rect 41548 4591 41588 4600
rect 41644 5312 41684 5321
rect 41644 2876 41684 5272
rect 42028 5060 42068 5069
rect 42028 4136 42068 5020
rect 42028 4087 42068 4096
rect 41740 3968 41780 3977
rect 41740 3833 41780 3928
rect 42220 3632 42260 9976
rect 43276 9680 43316 10312
rect 43276 9631 43316 9640
rect 44140 9848 44180 9857
rect 42220 3583 42260 3592
rect 42316 9512 42356 9521
rect 41932 3212 41972 3221
rect 41932 2960 41972 3172
rect 41932 2911 41972 2920
rect 41644 2827 41684 2836
rect 42028 2876 42068 2885
rect 42028 2741 42068 2836
rect 41932 2624 41972 2633
rect 41932 2372 41972 2584
rect 41932 2323 41972 2332
rect 42124 2624 42164 2633
rect 41260 2239 41300 2248
rect 41452 2239 41492 2248
rect 42124 2204 42164 2584
rect 42124 2155 42164 2164
rect 41260 104 41300 113
rect 41548 104 41588 113
rect 41260 60 41300 64
rect 41164 20 41300 60
rect 41528 64 41548 80
rect 42316 80 42356 9472
rect 42604 9512 42644 9521
rect 42412 9344 42452 9353
rect 42412 6572 42452 9304
rect 42412 6523 42452 6532
rect 42412 6404 42452 6413
rect 42412 6152 42452 6364
rect 42412 6103 42452 6112
rect 42412 5564 42452 5573
rect 42412 2876 42452 5524
rect 42412 2827 42452 2836
rect 42508 5396 42548 5405
rect 42508 2204 42548 5356
rect 42604 3296 42644 9472
rect 43084 9260 43124 9269
rect 42892 9220 43084 9260
rect 42892 9176 42932 9220
rect 43084 9211 43124 9220
rect 42892 9127 42932 9136
rect 43084 8672 43124 8681
rect 43084 6656 43124 8632
rect 43468 8672 43508 8681
rect 43276 7160 43316 7169
rect 43276 6992 43316 7120
rect 43276 6943 43316 6952
rect 43084 6607 43124 6616
rect 42988 5648 43028 5657
rect 42988 4724 43028 5608
rect 43468 5564 43508 8632
rect 43468 5515 43508 5524
rect 43852 7160 43892 7169
rect 43852 6236 43892 7120
rect 43852 5648 43892 6196
rect 42988 4220 43028 4684
rect 43756 5060 43796 5069
rect 43756 4556 43796 5020
rect 43756 4507 43796 4516
rect 43852 4724 43892 5608
rect 43852 4304 43892 4684
rect 43852 4255 43892 4264
rect 42988 3380 43028 4180
rect 42988 3331 43028 3340
rect 43084 4136 43124 4145
rect 42604 3247 42644 3256
rect 43084 3212 43124 4096
rect 43084 2876 43124 3172
rect 43084 2827 43124 2836
rect 43372 3548 43412 3557
rect 42508 2155 42548 2164
rect 42604 2792 42644 2801
rect 42604 1616 42644 2752
rect 43372 1952 43412 3508
rect 44140 3296 44180 9808
rect 44236 8924 44276 10648
rect 44428 10016 44468 10025
rect 44428 9680 44468 9976
rect 44428 9631 44468 9640
rect 44332 9260 44372 9269
rect 44332 9092 44372 9220
rect 44332 9043 44372 9052
rect 44236 8875 44276 8884
rect 44716 8168 44756 10984
rect 45196 9680 45236 9689
rect 45004 9344 45044 9353
rect 45004 8336 45044 9304
rect 45196 8924 45236 9640
rect 45196 8875 45236 8884
rect 45004 8287 45044 8296
rect 45772 8504 45812 8513
rect 44716 8119 44756 8128
rect 44332 8000 44372 8009
rect 44236 4892 44276 4901
rect 44332 4892 44372 7960
rect 45772 8000 45812 8464
rect 45772 7951 45812 7960
rect 45772 7748 45812 7757
rect 45772 7328 45812 7708
rect 45772 7279 45812 7288
rect 44908 7160 44948 7169
rect 44276 4852 44372 4892
rect 44428 6488 44468 6497
rect 44236 4843 44276 4852
rect 44428 3800 44468 6448
rect 44908 4724 44948 7120
rect 46156 7076 46196 7085
rect 46156 6656 46196 7036
rect 46252 6656 46292 6665
rect 46156 6616 46252 6656
rect 46252 6607 46292 6616
rect 46252 6152 46292 6161
rect 46252 5984 46292 6112
rect 46252 5935 46292 5944
rect 46252 5480 46292 5489
rect 46252 5312 46292 5440
rect 46252 5263 46292 5272
rect 44908 4675 44948 4684
rect 44524 4136 44564 4145
rect 44524 4001 44564 4096
rect 44908 4136 44948 4145
rect 44428 3751 44468 3760
rect 44140 3247 44180 3256
rect 43756 3128 43796 3137
rect 43756 2624 43796 3088
rect 44908 3044 44948 4096
rect 44908 2995 44948 3004
rect 45196 3296 45236 3305
rect 45196 2876 45236 3256
rect 45196 2827 45236 2836
rect 43756 2575 43796 2584
rect 45196 2624 45236 2633
rect 45100 2540 45140 2549
rect 43660 2456 43700 2465
rect 43660 2321 43700 2416
rect 44620 2456 44660 2465
rect 43372 1903 43412 1912
rect 44044 2204 44084 2213
rect 44044 1952 44084 2164
rect 44044 1903 44084 1912
rect 42604 1567 42644 1576
rect 42700 1868 42740 1877
rect 42700 1532 42740 1828
rect 43180 1868 43220 1877
rect 43180 1784 43220 1828
rect 43756 1868 43796 1877
rect 43948 1868 43988 1877
rect 43796 1828 43948 1868
rect 43756 1819 43796 1828
rect 43948 1819 43988 1828
rect 42700 1483 42740 1492
rect 43084 1744 43220 1784
rect 43084 80 43124 1744
rect 44620 1280 44660 2416
rect 45100 1952 45140 2500
rect 45196 2036 45236 2584
rect 45196 1987 45236 1996
rect 45100 1903 45140 1912
rect 45004 1532 45044 1541
rect 44620 1231 44660 1240
rect 44812 1448 44852 1457
rect 44812 944 44852 1408
rect 44812 895 44852 904
rect 45004 608 45044 1492
rect 45004 559 45044 568
rect 41588 64 41608 80
rect 41528 0 41608 64
rect 42296 0 42376 80
rect 43064 0 43144 80
<< via3 >>
rect 10540 11740 10580 11780
rect 3688 9808 3728 9848
rect 3770 9808 3810 9848
rect 3852 9808 3892 9848
rect 3934 9808 3974 9848
rect 4016 9808 4056 9848
rect 2860 9220 2900 9260
rect 1708 7624 1748 7664
rect 2860 7708 2900 7748
rect 3688 8296 3728 8336
rect 3770 8296 3810 8336
rect 3852 8296 3892 8336
rect 3934 8296 3974 8336
rect 4016 8296 4056 8336
rect 3688 6784 3728 6824
rect 3770 6784 3810 6824
rect 3852 6784 3892 6824
rect 3934 6784 3974 6824
rect 4016 6784 4056 6824
rect 4928 9052 4968 9092
rect 5010 9052 5050 9092
rect 5092 9052 5132 9092
rect 5174 9052 5214 9092
rect 5256 9052 5296 9092
rect 4928 7540 4968 7580
rect 5010 7540 5050 7580
rect 5092 7540 5132 7580
rect 5174 7540 5214 7580
rect 5256 7540 5296 7580
rect 4300 6952 4340 6992
rect 4204 6364 4244 6404
rect 5740 6280 5780 6320
rect 4928 6028 4968 6068
rect 5010 6028 5050 6068
rect 5092 6028 5132 6068
rect 5174 6028 5214 6068
rect 5256 6028 5296 6068
rect 3688 5272 3728 5312
rect 3770 5272 3810 5312
rect 3852 5272 3892 5312
rect 3934 5272 3974 5312
rect 4016 5272 4056 5312
rect 4396 4852 4436 4892
rect 3688 3760 3728 3800
rect 3770 3760 3810 3800
rect 3852 3760 3892 3800
rect 3934 3760 3974 3800
rect 4016 3760 4056 3800
rect 1900 3340 1940 3380
rect 2860 2500 2900 2540
rect 2092 2416 2132 2456
rect 7660 9136 7700 9176
rect 4928 4516 4968 4556
rect 5010 4516 5050 4556
rect 5092 4516 5132 4556
rect 5174 4516 5214 4556
rect 5256 4516 5296 4556
rect 4928 3004 4968 3044
rect 5010 3004 5050 3044
rect 5092 3004 5132 3044
rect 5174 3004 5214 3044
rect 5256 3004 5296 3044
rect 4684 2668 4724 2708
rect 3688 2248 3728 2288
rect 3770 2248 3810 2288
rect 3852 2248 3892 2288
rect 3934 2248 3974 2288
rect 4016 2248 4056 2288
rect 6412 6448 6452 6488
rect 6700 6448 6740 6488
rect 6796 6280 6836 6320
rect 7564 4852 7604 4892
rect 7468 3508 7508 3548
rect 7948 6868 7988 6908
rect 7948 4264 7988 4304
rect 8908 5440 8948 5480
rect 4928 1492 4968 1532
rect 5010 1492 5050 1532
rect 5092 1492 5132 1532
rect 5174 1492 5214 1532
rect 5256 1492 5296 1532
rect 8428 2332 8468 2372
rect 9196 4264 9236 4304
rect 9484 8716 9524 8756
rect 9964 8800 10004 8840
rect 8908 2584 8948 2624
rect 9868 7540 9908 7580
rect 9484 4768 9524 4808
rect 9580 3424 9620 3464
rect 10252 9388 10292 9428
rect 10156 7876 10196 7916
rect 10252 6532 10292 6572
rect 10252 6112 10292 6152
rect 10444 7372 10484 7412
rect 11020 11740 11060 11780
rect 10636 9976 10676 10016
rect 10732 8884 10772 8924
rect 10636 8044 10676 8084
rect 10636 7876 10676 7916
rect 10732 7288 10772 7328
rect 10636 7204 10676 7244
rect 10732 6532 10772 6572
rect 9868 3424 9908 3464
rect 9772 2668 9812 2708
rect 10060 4180 10100 4220
rect 10732 4432 10772 4472
rect 11116 8464 11156 8504
rect 11020 7204 11060 7244
rect 11020 7036 11060 7076
rect 11116 6700 11156 6740
rect 10924 4516 10964 4556
rect 11212 6028 11252 6068
rect 11308 5692 11348 5732
rect 11500 8800 11540 8840
rect 11500 8044 11540 8084
rect 11596 6700 11636 6740
rect 11500 5776 11540 5816
rect 11980 8380 12020 8420
rect 11980 7960 12020 8000
rect 11884 6196 11924 6236
rect 11884 6028 11924 6068
rect 11692 5104 11732 5144
rect 11980 5608 12020 5648
rect 11212 2332 11252 2372
rect 11980 3088 12020 3128
rect 12268 6532 12308 6572
rect 12172 4684 12212 4724
rect 12460 8380 12500 8420
rect 12652 9892 12692 9932
rect 12652 7456 12692 7496
rect 12844 9052 12884 9092
rect 13036 9052 13076 9092
rect 12940 8464 12980 8504
rect 13420 9976 13460 10016
rect 13132 8044 13172 8084
rect 13036 7792 13076 7832
rect 12940 7204 12980 7244
rect 13132 7288 13172 7328
rect 12748 6700 12788 6740
rect 12460 6028 12500 6068
rect 12652 6028 12692 6068
rect 12748 5944 12788 5984
rect 12748 5272 12788 5312
rect 12268 4264 12308 4304
rect 12940 6784 12980 6824
rect 12940 5860 12980 5900
rect 13708 9556 13748 9596
rect 13516 6616 13556 6656
rect 13324 6112 13364 6152
rect 12940 5524 12980 5564
rect 12844 3928 12884 3968
rect 12364 3592 12404 3632
rect 12460 3424 12500 3464
rect 12940 3424 12980 3464
rect 12940 2920 12980 2960
rect 13228 3844 13268 3884
rect 13420 3676 13460 3716
rect 13420 3424 13460 3464
rect 13708 4012 13748 4052
rect 13708 3760 13748 3800
rect 13132 2920 13172 2960
rect 13228 2836 13268 2876
rect 14284 9556 14324 9596
rect 14380 9892 14420 9932
rect 14188 7372 14228 7412
rect 13996 6784 14036 6824
rect 13996 6028 14036 6068
rect 13900 5776 13940 5816
rect 13996 5860 14036 5900
rect 13900 5524 13940 5564
rect 13804 3256 13844 3296
rect 12652 2164 12692 2204
rect 12748 1996 12788 2036
rect 11500 1660 11540 1700
rect 11980 1744 12020 1784
rect 12940 1996 12980 2036
rect 13900 2080 13940 2120
rect 13324 1492 13364 1532
rect 14188 5188 14228 5228
rect 14188 3760 14228 3800
rect 14764 8212 14804 8252
rect 14956 8800 14996 8840
rect 14764 6616 14804 6656
rect 15148 8800 15188 8840
rect 15628 8800 15668 8840
rect 15724 9052 15764 9092
rect 15148 6028 15188 6068
rect 14572 5272 14612 5312
rect 14668 4348 14708 4388
rect 14092 1828 14132 1868
rect 14476 2332 14516 2372
rect 14476 1492 14516 1532
rect 15532 7540 15572 7580
rect 15436 7456 15476 7496
rect 15628 5524 15668 5564
rect 15340 3004 15380 3044
rect 15148 2584 15188 2624
rect 15628 4348 15668 4388
rect 15628 4012 15668 4052
rect 15916 7792 15956 7832
rect 15916 7120 15956 7160
rect 16204 8968 16244 9008
rect 16300 7288 16340 7328
rect 16492 7036 16532 7076
rect 15820 5860 15860 5900
rect 16492 4432 16532 4472
rect 16204 3424 16244 3464
rect 15628 3004 15668 3044
rect 15436 1912 15476 1952
rect 16300 3172 16340 3212
rect 16204 2584 16244 2624
rect 16204 1996 16244 2036
rect 17452 9304 17492 9344
rect 17068 5020 17108 5060
rect 17260 2920 17300 2960
rect 17644 7204 17684 7244
rect 17548 3844 17588 3884
rect 18028 9556 18068 9596
rect 19276 10144 19316 10184
rect 18124 8464 18164 8504
rect 18412 8884 18452 8924
rect 18028 7456 18068 7496
rect 18028 6112 18068 6152
rect 17932 4012 17972 4052
rect 17932 3592 17972 3632
rect 17644 2752 17684 2792
rect 15628 1576 15668 1616
rect 17932 1996 17972 2036
rect 18124 4264 18164 4304
rect 18412 7456 18452 7496
rect 18604 8632 18644 8672
rect 18604 8128 18644 8168
rect 18604 7288 18644 7328
rect 18808 9808 18848 9848
rect 18890 9808 18930 9848
rect 18972 9808 19012 9848
rect 19054 9808 19094 9848
rect 19136 9808 19176 9848
rect 19180 9472 19220 9512
rect 18988 8800 19028 8840
rect 19564 10144 19604 10184
rect 19564 9304 19604 9344
rect 19468 9052 19508 9092
rect 19372 8632 19412 8672
rect 18808 8296 18848 8336
rect 18890 8296 18930 8336
rect 18972 8296 19012 8336
rect 19054 8296 19094 8336
rect 19136 8296 19176 8336
rect 19276 8296 19316 8336
rect 19180 7540 19220 7580
rect 18892 7288 18932 7328
rect 18892 7036 18932 7076
rect 18808 6784 18848 6824
rect 18890 6784 18930 6824
rect 18972 6784 19012 6824
rect 19054 6784 19094 6824
rect 19136 6784 19176 6824
rect 19276 6700 19316 6740
rect 18604 5356 18644 5396
rect 18700 5860 18740 5900
rect 19276 5356 19316 5396
rect 18808 5272 18848 5312
rect 18890 5272 18930 5312
rect 18972 5272 19012 5312
rect 19054 5272 19094 5312
rect 19136 5272 19176 5312
rect 18796 4516 18836 4556
rect 18808 3760 18848 3800
rect 18890 3760 18930 3800
rect 18972 3760 19012 3800
rect 19054 3760 19094 3800
rect 19136 3760 19176 3800
rect 18796 3592 18836 3632
rect 18508 2920 18548 2960
rect 19852 10060 19892 10100
rect 20140 10564 20180 10604
rect 20044 9472 20084 9512
rect 19852 9052 19892 9092
rect 19948 9388 19988 9428
rect 20236 9304 20276 9344
rect 20048 9052 20088 9092
rect 20130 9052 20170 9092
rect 20212 9052 20252 9092
rect 20294 9052 20334 9092
rect 20376 9052 20416 9092
rect 20236 8884 20276 8924
rect 20236 8632 20276 8672
rect 20332 8548 20372 8588
rect 20428 8632 20468 8672
rect 20236 8380 20276 8420
rect 19948 8212 19988 8252
rect 19756 8044 19796 8084
rect 20044 8044 20084 8084
rect 20332 8044 20372 8084
rect 19660 7540 19700 7580
rect 20048 7540 20088 7580
rect 20130 7540 20170 7580
rect 20212 7540 20252 7580
rect 20294 7540 20334 7580
rect 20376 7540 20416 7580
rect 19756 7372 19796 7412
rect 19756 7036 19796 7076
rect 18316 2584 18356 2624
rect 18412 1996 18452 2036
rect 18808 2248 18848 2288
rect 18890 2248 18930 2288
rect 18972 2248 19012 2288
rect 19054 2248 19094 2288
rect 19136 2248 19176 2288
rect 19468 2920 19508 2960
rect 20140 7036 20180 7076
rect 20908 9388 20948 9428
rect 21100 8800 21140 8840
rect 21100 8296 21140 8336
rect 21196 8632 21236 8672
rect 19756 4432 19796 4472
rect 20048 6028 20088 6068
rect 20130 6028 20170 6068
rect 20212 6028 20252 6068
rect 20294 6028 20334 6068
rect 20376 6028 20416 6068
rect 20044 5776 20084 5816
rect 20812 5944 20852 5984
rect 20048 4516 20088 4556
rect 20130 4516 20170 4556
rect 20212 4516 20252 4556
rect 20294 4516 20334 4556
rect 20376 4516 20416 4556
rect 20140 4012 20180 4052
rect 20048 3004 20088 3044
rect 20130 3004 20170 3044
rect 20212 3004 20252 3044
rect 20294 3004 20334 3044
rect 20376 3004 20416 3044
rect 20812 3760 20852 3800
rect 20044 2248 20084 2288
rect 19948 2164 19988 2204
rect 21580 10564 21620 10604
rect 21580 9640 21620 9680
rect 21676 9388 21716 9428
rect 21484 8884 21524 8924
rect 21484 8380 21524 8420
rect 21196 3592 21236 3632
rect 21676 8464 21716 8504
rect 21868 8884 21908 8924
rect 21676 7456 21716 7496
rect 21580 6868 21620 6908
rect 21580 5188 21620 5228
rect 21100 2836 21140 2876
rect 21292 2836 21332 2876
rect 21292 2332 21332 2372
rect 21004 1912 21044 1952
rect 21772 6868 21812 6908
rect 22060 9808 22100 9848
rect 22060 9052 22100 9092
rect 22540 9640 22580 9680
rect 23404 9640 23444 9680
rect 23212 9556 23252 9596
rect 24460 10648 24500 10688
rect 22348 8884 22388 8924
rect 22252 4348 22292 4388
rect 22540 8296 22580 8336
rect 22444 8128 22484 8168
rect 22540 7204 22580 7244
rect 23692 9052 23732 9092
rect 22732 8380 22772 8420
rect 23404 8044 23444 8084
rect 22732 7120 22772 7160
rect 23212 7036 23252 7076
rect 22924 5944 22964 5984
rect 23404 6028 23444 6068
rect 23404 5860 23444 5900
rect 22828 5776 22868 5816
rect 21964 3592 22004 3632
rect 21868 2248 21908 2288
rect 22252 2248 22292 2288
rect 21772 1828 21812 1868
rect 20524 1576 20564 1616
rect 20048 1492 20088 1532
rect 20130 1492 20170 1532
rect 20212 1492 20252 1532
rect 20294 1492 20334 1532
rect 20376 1492 20416 1532
rect 19948 820 19988 860
rect 20812 820 20852 860
rect 22732 2248 22772 2288
rect 22636 2080 22676 2120
rect 23020 5776 23060 5816
rect 23212 5356 23252 5396
rect 22924 4852 22964 4892
rect 23116 4432 23156 4472
rect 22924 3088 22964 3128
rect 23692 4936 23732 4976
rect 23596 4516 23636 4556
rect 23788 4348 23828 4388
rect 23212 2248 23252 2288
rect 23020 2164 23060 2204
rect 23308 1492 23348 1532
rect 24460 8716 24500 8756
rect 24268 8464 24308 8504
rect 24172 5356 24212 5396
rect 24076 4852 24116 4892
rect 23692 1996 23732 2036
rect 24268 4936 24308 4976
rect 24268 4348 24308 4388
rect 24556 8464 24596 8504
rect 24652 7204 24692 7244
rect 24556 4852 24596 4892
rect 24748 3676 24788 3716
rect 24940 8800 24980 8840
rect 24940 8632 24980 8672
rect 25228 10816 25268 10856
rect 25228 10648 25268 10688
rect 25612 10564 25652 10604
rect 25996 10900 26036 10940
rect 25804 10312 25844 10352
rect 25612 8716 25652 8756
rect 25324 6868 25364 6908
rect 24940 4264 24980 4304
rect 26092 9220 26132 9260
rect 26380 11152 26420 11192
rect 26764 11320 26804 11360
rect 26572 8632 26612 8672
rect 26476 8548 26516 8588
rect 25900 7204 25940 7244
rect 27148 10060 27188 10100
rect 27724 10312 27764 10352
rect 27532 9556 27572 9596
rect 27628 10060 27668 10100
rect 27340 9388 27380 9428
rect 27340 8968 27380 9008
rect 27052 8716 27092 8756
rect 27244 8800 27284 8840
rect 27436 8800 27476 8840
rect 27820 9892 27860 9932
rect 27820 9136 27860 9176
rect 27148 7288 27188 7328
rect 27340 7288 27380 7328
rect 25708 5860 25748 5900
rect 25228 3508 25268 3548
rect 25228 2920 25268 2960
rect 24268 2668 24308 2708
rect 24268 2332 24308 2372
rect 24556 2668 24596 2708
rect 25132 2164 25172 2204
rect 25516 2668 25556 2708
rect 26188 4432 26228 4472
rect 25996 3340 26036 3380
rect 26380 3340 26420 3380
rect 27340 6532 27380 6572
rect 27532 2668 27572 2708
rect 26284 1492 26324 1532
rect 27724 7540 27764 7580
rect 28300 10984 28340 11024
rect 28300 10816 28340 10856
rect 28300 9136 28340 9176
rect 28876 10900 28916 10940
rect 28684 10564 28724 10604
rect 28588 9808 28628 9848
rect 28588 9052 28628 9092
rect 28684 8632 28724 8672
rect 28492 8044 28532 8084
rect 29068 9640 29108 9680
rect 29356 10060 29396 10100
rect 29452 11152 29492 11192
rect 29836 11488 29876 11528
rect 29644 10732 29684 10772
rect 29836 11320 29876 11360
rect 29644 9892 29684 9932
rect 30028 11404 30068 11444
rect 29260 8632 29300 8672
rect 29164 8548 29204 8588
rect 29644 8548 29684 8588
rect 29068 7288 29108 7328
rect 28684 3508 28724 3548
rect 28780 6028 28820 6068
rect 28972 5944 29012 5984
rect 29740 7036 29780 7076
rect 29836 6868 29876 6908
rect 29740 6784 29780 6824
rect 29836 6532 29876 6572
rect 28876 4936 28916 4976
rect 29836 6112 29876 6152
rect 28876 4264 28916 4304
rect 29740 4936 29780 4976
rect 29260 4264 29300 4304
rect 29644 3760 29684 3800
rect 29548 3592 29588 3632
rect 29740 2668 29780 2708
rect 30412 10648 30452 10688
rect 30220 9976 30260 10016
rect 30700 9556 30740 9596
rect 30124 9388 30164 9428
rect 30124 8968 30164 9008
rect 30028 6868 30068 6908
rect 30412 9304 30452 9344
rect 30220 8044 30260 8084
rect 30316 6784 30356 6824
rect 30412 7120 30452 7160
rect 29452 2080 29492 2120
rect 30124 4516 30164 4556
rect 30220 3508 30260 3548
rect 30892 10060 30932 10100
rect 30988 8632 31028 8672
rect 31084 8128 31124 8168
rect 31372 10144 31412 10184
rect 31372 7624 31412 7664
rect 31276 6448 31316 6488
rect 31468 6868 31508 6908
rect 31660 10984 31700 11024
rect 31852 9976 31892 10016
rect 31756 9220 31796 9260
rect 31852 5860 31892 5900
rect 31756 5776 31796 5816
rect 32332 11236 32372 11276
rect 32428 9304 32468 9344
rect 32140 8716 32180 8756
rect 32716 11152 32756 11192
rect 32236 7876 32276 7916
rect 31084 4264 31124 4304
rect 31852 3844 31892 3884
rect 32428 5020 32468 5060
rect 32140 4180 32180 4220
rect 30796 988 30836 1028
rect 32332 3844 32372 3884
rect 31852 2332 31892 2372
rect 32140 1912 32180 1952
rect 33196 9220 33236 9260
rect 33004 8968 33044 9008
rect 33388 9052 33428 9092
rect 33196 8800 33236 8840
rect 33004 8380 33044 8420
rect 32620 7540 32660 7580
rect 33100 7372 33140 7412
rect 32908 7036 32948 7076
rect 32620 6784 32660 6824
rect 32716 6532 32756 6572
rect 32812 6448 32852 6488
rect 33388 8464 33428 8504
rect 33292 7120 33332 7160
rect 33388 7036 33428 7076
rect 33004 5356 33044 5396
rect 33100 5020 33140 5060
rect 32812 4936 32852 4976
rect 34060 9976 34100 10016
rect 34540 10732 34580 10772
rect 33772 9892 33812 9932
rect 33928 9808 33968 9848
rect 34010 9808 34050 9848
rect 34092 9808 34132 9848
rect 34174 9808 34214 9848
rect 34256 9808 34296 9848
rect 33676 7036 33716 7076
rect 33580 6868 33620 6908
rect 33388 6112 33428 6152
rect 32908 4432 32948 4472
rect 33292 4600 33332 4640
rect 33100 2836 33140 2876
rect 33676 4936 33716 4976
rect 33676 4768 33716 4808
rect 33676 3256 33716 3296
rect 33868 8968 33908 9008
rect 33928 8296 33968 8336
rect 34010 8296 34050 8336
rect 34092 8296 34132 8336
rect 34174 8296 34214 8336
rect 34256 8296 34296 8336
rect 34060 8128 34100 8168
rect 33964 7204 34004 7244
rect 34252 8128 34292 8168
rect 34540 9304 34580 9344
rect 34444 8968 34484 9008
rect 34348 7288 34388 7328
rect 34156 7120 34196 7160
rect 33868 7036 33908 7076
rect 33928 6784 33968 6824
rect 34010 6784 34050 6824
rect 34092 6784 34132 6824
rect 34174 6784 34214 6824
rect 34256 6784 34296 6824
rect 34924 7540 34964 7580
rect 33928 5272 33968 5312
rect 34010 5272 34050 5312
rect 34092 5272 34132 5312
rect 34174 5272 34214 5312
rect 34256 5272 34296 5312
rect 34924 6448 34964 6488
rect 34828 5776 34868 5816
rect 33928 3760 33968 3800
rect 34010 3760 34050 3800
rect 34092 3760 34132 3800
rect 34174 3760 34214 3800
rect 34256 3760 34296 3800
rect 34540 5104 34580 5144
rect 37228 11236 37268 11276
rect 35980 10648 36020 10688
rect 35788 9892 35828 9932
rect 35308 9304 35348 9344
rect 35168 9052 35208 9092
rect 35250 9052 35290 9092
rect 35332 9052 35372 9092
rect 35414 9052 35454 9092
rect 35496 9052 35536 9092
rect 35212 8380 35252 8420
rect 35116 8128 35156 8168
rect 35168 7540 35208 7580
rect 35250 7540 35290 7580
rect 35332 7540 35372 7580
rect 35414 7540 35454 7580
rect 35496 7540 35536 7580
rect 35168 6028 35208 6068
rect 35250 6028 35290 6068
rect 35332 6028 35372 6068
rect 35414 6028 35454 6068
rect 35496 6028 35536 6068
rect 35020 5692 35060 5732
rect 36172 10144 36212 10184
rect 36652 9892 36692 9932
rect 37516 11152 37556 11192
rect 35692 6280 35732 6320
rect 35116 5020 35156 5060
rect 35168 4516 35208 4556
rect 35250 4516 35290 4556
rect 35332 4516 35372 4556
rect 35414 4516 35454 4556
rect 35496 4516 35536 4556
rect 35168 3004 35208 3044
rect 35250 3004 35290 3044
rect 35332 3004 35372 3044
rect 35414 3004 35454 3044
rect 35496 3004 35536 3044
rect 33928 2248 33968 2288
rect 34010 2248 34050 2288
rect 34092 2248 34132 2288
rect 34174 2248 34214 2288
rect 34256 2248 34296 2288
rect 33676 1744 33716 1784
rect 33100 64 33140 104
rect 33868 64 33908 104
rect 34060 64 34100 104
rect 34444 1744 34484 1784
rect 35500 2752 35540 2792
rect 35980 7792 36020 7832
rect 36268 7456 36308 7496
rect 36748 7120 36788 7160
rect 36364 6532 36404 6572
rect 35980 5440 36020 5480
rect 37036 7204 37076 7244
rect 36844 6700 36884 6740
rect 37132 6364 37172 6404
rect 36556 5860 36596 5900
rect 36460 5608 36500 5648
rect 36172 5356 36212 5396
rect 35884 3424 35924 3464
rect 36172 2500 36212 2540
rect 35692 1912 35732 1952
rect 35168 1492 35208 1532
rect 35250 1492 35290 1532
rect 35332 1492 35372 1532
rect 35414 1492 35454 1532
rect 35496 1492 35536 1532
rect 37324 8716 37364 8756
rect 37324 6868 37364 6908
rect 37228 2164 37268 2204
rect 37804 9220 37844 9260
rect 38764 9976 38804 10016
rect 39340 9136 39380 9176
rect 37900 7372 37940 7412
rect 37900 4936 37940 4976
rect 37900 2836 37940 2876
rect 37900 2164 37940 2204
rect 38188 6364 38228 6404
rect 38764 7960 38804 8000
rect 38668 7120 38708 7160
rect 38572 4264 38612 4304
rect 38476 4012 38516 4052
rect 39436 7624 39476 7664
rect 39244 4432 39284 4472
rect 38956 4264 38996 4304
rect 39532 4012 39572 4052
rect 38668 2248 38708 2288
rect 38956 2584 38996 2624
rect 38668 1492 38708 1532
rect 38956 1492 38996 1532
rect 39052 988 39092 1028
rect 39820 3172 39860 3212
rect 39340 148 39380 188
rect 40300 9052 40340 9092
rect 40108 7288 40148 7328
rect 40300 2416 40340 2456
rect 40300 2248 40340 2288
rect 40396 1744 40436 1784
rect 41164 4600 41204 4640
rect 40876 1660 40916 1700
rect 41740 6196 41780 6236
rect 41548 4600 41588 4640
rect 41740 3928 41780 3968
rect 42028 2836 42068 2876
rect 41260 64 41300 104
rect 41548 64 41588 104
rect 43276 6952 43316 6992
rect 43084 6616 43124 6656
rect 43468 5524 43508 5564
rect 44332 9052 44372 9092
rect 44908 4684 44948 4724
rect 44524 4096 44564 4136
rect 43660 2416 43700 2456
rect 44620 2416 44660 2456
<< metal4 >>
rect 10531 11740 10540 11780
rect 10580 11740 11020 11780
rect 11060 11740 11069 11780
rect 29827 11488 29836 11528
rect 29876 11488 29885 11528
rect 29836 11444 29876 11488
rect 29836 11404 30028 11444
rect 30068 11404 30077 11444
rect 26755 11320 26764 11360
rect 26804 11320 29836 11360
rect 29876 11320 29885 11360
rect 32323 11236 32332 11276
rect 32372 11236 37228 11276
rect 37268 11236 37277 11276
rect 26371 11152 26380 11192
rect 26420 11152 29452 11192
rect 29492 11152 29501 11192
rect 32707 11152 32716 11192
rect 32756 11152 37516 11192
rect 37556 11152 37565 11192
rect 28291 10984 28300 11024
rect 28340 10984 31660 11024
rect 31700 10984 31709 11024
rect 25987 10900 25996 10940
rect 26036 10900 28876 10940
rect 28916 10900 28925 10940
rect 25219 10816 25228 10856
rect 25268 10816 28300 10856
rect 28340 10816 28349 10856
rect 29635 10732 29644 10772
rect 29684 10732 34540 10772
rect 34580 10732 34589 10772
rect 24451 10648 24460 10688
rect 24500 10648 25228 10688
rect 25268 10648 25277 10688
rect 30403 10648 30412 10688
rect 30452 10648 35980 10688
rect 36020 10648 36029 10688
rect 20131 10564 20140 10604
rect 20180 10564 21580 10604
rect 21620 10564 21629 10604
rect 25603 10564 25612 10604
rect 25652 10564 28684 10604
rect 28724 10564 28733 10604
rect 25795 10312 25804 10352
rect 25844 10312 27724 10352
rect 27764 10312 27773 10352
rect 19267 10144 19276 10184
rect 19316 10144 19564 10184
rect 19604 10144 19613 10184
rect 31363 10144 31372 10184
rect 31412 10144 36172 10184
rect 36212 10144 36221 10184
rect 19757 10060 19852 10100
rect 19892 10060 19901 10100
rect 27139 10060 27148 10100
rect 27188 10060 27628 10100
rect 27668 10060 27677 10100
rect 29347 10060 29356 10100
rect 29396 10060 30892 10100
rect 30932 10060 30941 10100
rect 10627 9976 10636 10016
rect 10676 9976 13420 10016
rect 13460 9976 13469 10016
rect 30211 9976 30220 10016
rect 30260 9976 31852 10016
rect 31892 9976 31901 10016
rect 34051 9976 34060 10016
rect 34100 9976 38764 10016
rect 38804 9976 38813 10016
rect 12643 9892 12652 9932
rect 12692 9892 14380 9932
rect 14420 9892 14429 9932
rect 27811 9892 27820 9932
rect 27860 9892 29644 9932
rect 29684 9892 29693 9932
rect 33763 9892 33772 9932
rect 33812 9892 35788 9932
rect 35828 9892 36652 9932
rect 36692 9892 36701 9932
rect 3679 9808 3688 9848
rect 3728 9808 3770 9848
rect 3810 9808 3852 9848
rect 3892 9808 3934 9848
rect 3974 9808 4016 9848
rect 4056 9808 4065 9848
rect 18799 9808 18808 9848
rect 18848 9808 18890 9848
rect 18930 9808 18972 9848
rect 19012 9808 19054 9848
rect 19094 9808 19136 9848
rect 19176 9808 19185 9848
rect 22051 9808 22060 9848
rect 22100 9808 28588 9848
rect 28628 9808 28637 9848
rect 33919 9808 33928 9848
rect 33968 9808 34010 9848
rect 34050 9808 34092 9848
rect 34132 9808 34174 9848
rect 34214 9808 34256 9848
rect 34296 9808 34305 9848
rect 21571 9640 21580 9680
rect 21620 9640 22540 9680
rect 22580 9640 22589 9680
rect 23395 9640 23404 9680
rect 23444 9640 29068 9680
rect 29108 9640 29117 9680
rect 13699 9556 13708 9596
rect 13748 9556 14284 9596
rect 14324 9556 14333 9596
rect 18019 9556 18028 9596
rect 18068 9556 23212 9596
rect 23252 9556 23261 9596
rect 27523 9556 27532 9596
rect 27572 9556 30700 9596
rect 30740 9556 30749 9596
rect 19171 9472 19180 9512
rect 19220 9472 20044 9512
rect 20084 9472 20093 9512
rect 10243 9388 10252 9428
rect 10292 9388 19948 9428
rect 19988 9388 19997 9428
rect 20899 9388 20908 9428
rect 20948 9388 21676 9428
rect 21716 9388 21725 9428
rect 27331 9388 27340 9428
rect 27380 9388 30124 9428
rect 30164 9388 30173 9428
rect 17443 9304 17452 9344
rect 17492 9304 19564 9344
rect 19604 9304 19613 9344
rect 20227 9304 20236 9344
rect 20276 9304 20524 9344
rect 20564 9304 20573 9344
rect 23020 9304 30412 9344
rect 30452 9304 32428 9344
rect 32468 9304 32477 9344
rect 34531 9304 34540 9344
rect 34580 9304 35308 9344
rect 35348 9304 35357 9344
rect 23020 9260 23060 9304
rect 2851 9220 2860 9260
rect 2900 9220 23060 9260
rect 26083 9220 26092 9260
rect 26132 9220 31756 9260
rect 31796 9220 31805 9260
rect 33187 9220 33196 9260
rect 33236 9220 37804 9260
rect 37844 9220 37853 9260
rect 7651 9136 7660 9176
rect 7700 9136 27820 9176
rect 27860 9136 27869 9176
rect 28291 9136 28300 9176
rect 28340 9136 39340 9176
rect 39380 9136 39389 9176
rect 4919 9052 4928 9092
rect 4968 9052 5010 9092
rect 5050 9052 5092 9092
rect 5132 9052 5174 9092
rect 5214 9052 5256 9092
rect 5296 9052 5305 9092
rect 12835 9052 12844 9092
rect 12884 9052 13036 9092
rect 13076 9052 13085 9092
rect 15715 9052 15724 9092
rect 15764 9052 19468 9092
rect 19508 9052 19852 9092
rect 19892 9052 19901 9092
rect 20039 9052 20048 9092
rect 20088 9052 20130 9092
rect 20170 9052 20212 9092
rect 20252 9052 20294 9092
rect 20334 9052 20376 9092
rect 20416 9052 20425 9092
rect 22051 9052 22060 9092
rect 22100 9052 23692 9092
rect 23732 9052 28588 9092
rect 28628 9052 28637 9092
rect 33293 9052 33388 9092
rect 33428 9052 33437 9092
rect 35159 9052 35168 9092
rect 35208 9052 35250 9092
rect 35290 9052 35332 9092
rect 35372 9052 35414 9092
rect 35454 9052 35496 9092
rect 35536 9052 35545 9092
rect 40291 9052 40300 9092
rect 40340 9052 44332 9092
rect 44372 9052 44381 9092
rect 16195 8968 16204 9008
rect 16244 8968 27340 9008
rect 27380 8968 27389 9008
rect 30115 8968 30124 9008
rect 30164 8968 33004 9008
rect 33044 8968 33053 9008
rect 33859 8968 33868 9008
rect 33908 8968 34444 9008
rect 34484 8968 34493 9008
rect 10723 8884 10732 8924
rect 10772 8884 18412 8924
rect 18452 8884 18461 8924
rect 20227 8884 20236 8924
rect 20276 8884 21484 8924
rect 21524 8884 21533 8924
rect 21859 8884 21868 8924
rect 21908 8884 22348 8924
rect 22388 8884 22397 8924
rect 9955 8800 9964 8840
rect 10004 8800 11500 8840
rect 11540 8800 14956 8840
rect 14996 8800 15005 8840
rect 15139 8800 15148 8840
rect 15188 8800 15628 8840
rect 15668 8800 15677 8840
rect 18979 8800 18988 8840
rect 19028 8800 21100 8840
rect 21140 8800 21149 8840
rect 24931 8800 24940 8840
rect 24980 8800 27244 8840
rect 27284 8800 27436 8840
rect 27476 8800 27485 8840
rect 33187 8800 33196 8840
rect 33236 8800 33331 8840
rect 9475 8716 9484 8756
rect 9524 8716 24460 8756
rect 24500 8716 24509 8756
rect 25603 8716 25612 8756
rect 25652 8716 27052 8756
rect 27092 8716 27101 8756
rect 32131 8716 32140 8756
rect 32180 8716 37324 8756
rect 37364 8716 37373 8756
rect 18595 8632 18604 8672
rect 18644 8632 19372 8672
rect 19412 8632 19421 8672
rect 20227 8632 20236 8672
rect 20276 8632 20428 8672
rect 20468 8632 20477 8672
rect 21187 8632 21196 8672
rect 21236 8632 24940 8672
rect 24980 8632 24989 8672
rect 26563 8632 26572 8672
rect 26612 8632 28684 8672
rect 28724 8632 28733 8672
rect 29251 8632 29260 8672
rect 29300 8632 30988 8672
rect 31028 8632 31037 8672
rect 20323 8548 20332 8588
rect 20372 8548 26476 8588
rect 26516 8548 26525 8588
rect 29155 8548 29164 8588
rect 29204 8548 29644 8588
rect 29684 8548 29693 8588
rect 11107 8464 11116 8504
rect 11156 8464 12940 8504
rect 12980 8464 12989 8504
rect 18115 8464 18124 8504
rect 18164 8464 21676 8504
rect 21716 8464 21725 8504
rect 24259 8464 24268 8504
rect 24308 8464 24556 8504
rect 24596 8464 24605 8504
rect 33293 8464 33388 8504
rect 33428 8464 33437 8504
rect 11971 8380 11980 8420
rect 12020 8380 12460 8420
rect 12500 8380 12509 8420
rect 20227 8380 20236 8420
rect 20276 8380 20524 8420
rect 20564 8380 20573 8420
rect 21475 8380 21484 8420
rect 21524 8380 22732 8420
rect 22772 8380 22781 8420
rect 32995 8380 33004 8420
rect 33044 8380 35212 8420
rect 35252 8380 35261 8420
rect 3679 8296 3688 8336
rect 3728 8296 3770 8336
rect 3810 8296 3852 8336
rect 3892 8296 3934 8336
rect 3974 8296 4016 8336
rect 4056 8296 4065 8336
rect 18799 8296 18808 8336
rect 18848 8296 18890 8336
rect 18930 8296 18972 8336
rect 19012 8296 19054 8336
rect 19094 8296 19136 8336
rect 19176 8296 19185 8336
rect 19267 8296 19276 8336
rect 19316 8296 20908 8336
rect 20948 8296 20957 8336
rect 21091 8296 21100 8336
rect 21140 8296 22540 8336
rect 22580 8296 22589 8336
rect 33919 8296 33928 8336
rect 33968 8296 34010 8336
rect 34050 8296 34092 8336
rect 34132 8296 34174 8336
rect 34214 8296 34256 8336
rect 34296 8296 34305 8336
rect 14755 8212 14764 8252
rect 14804 8212 19948 8252
rect 19988 8212 19997 8252
rect 18595 8128 18604 8168
rect 18644 8128 22444 8168
rect 22484 8128 22493 8168
rect 31075 8128 31084 8168
rect 31124 8128 34060 8168
rect 34100 8128 34109 8168
rect 34243 8128 34252 8168
rect 34292 8128 35116 8168
rect 35156 8128 35165 8168
rect 10627 8044 10636 8084
rect 10676 8044 11500 8084
rect 11540 8044 11549 8084
rect 13123 8044 13132 8084
rect 13172 8044 19468 8084
rect 19508 8044 19517 8084
rect 19747 8044 19756 8084
rect 19796 8044 20044 8084
rect 20084 8044 20093 8084
rect 20323 8044 20332 8084
rect 20372 8044 23404 8084
rect 23444 8044 23453 8084
rect 28483 8044 28492 8084
rect 28532 8044 30220 8084
rect 30260 8044 30269 8084
rect 11971 7960 11980 8000
rect 12020 7960 38764 8000
rect 38804 7960 38813 8000
rect 10147 7876 10156 7916
rect 10196 7876 10636 7916
rect 10676 7876 32236 7916
rect 32276 7876 32285 7916
rect 13027 7792 13036 7832
rect 13076 7792 13171 7832
rect 15907 7792 15916 7832
rect 15956 7792 35980 7832
rect 36020 7792 36029 7832
rect 2851 7708 2860 7748
rect 2900 7708 33140 7748
rect 33100 7664 33140 7708
rect 1699 7624 1708 7664
rect 1748 7624 31372 7664
rect 31412 7624 31421 7664
rect 33100 7624 39436 7664
rect 39476 7624 39485 7664
rect 4919 7540 4928 7580
rect 4968 7540 5010 7580
rect 5050 7540 5092 7580
rect 5132 7540 5174 7580
rect 5214 7540 5256 7580
rect 5296 7540 5305 7580
rect 9859 7540 9868 7580
rect 9908 7540 15532 7580
rect 15572 7540 15581 7580
rect 19171 7540 19180 7580
rect 19220 7540 19660 7580
rect 19700 7540 19709 7580
rect 20039 7540 20048 7580
rect 20088 7540 20130 7580
rect 20170 7540 20212 7580
rect 20252 7540 20294 7580
rect 20334 7540 20376 7580
rect 20416 7540 20425 7580
rect 27715 7540 27724 7580
rect 27764 7540 30260 7580
rect 32611 7540 32620 7580
rect 32660 7540 34924 7580
rect 34964 7540 34973 7580
rect 35159 7540 35168 7580
rect 35208 7540 35250 7580
rect 35290 7540 35332 7580
rect 35372 7540 35414 7580
rect 35454 7540 35496 7580
rect 35536 7540 35545 7580
rect 30220 7496 30260 7540
rect 12643 7456 12652 7496
rect 12692 7456 15436 7496
rect 15476 7456 18028 7496
rect 18068 7456 18077 7496
rect 18403 7456 18412 7496
rect 18452 7456 21676 7496
rect 21716 7456 21725 7496
rect 30220 7456 36268 7496
rect 36308 7456 36317 7496
rect 10435 7372 10444 7412
rect 10484 7372 14188 7412
rect 14228 7372 14237 7412
rect 19747 7372 19756 7412
rect 19796 7372 19852 7412
rect 19892 7372 19901 7412
rect 33091 7372 33100 7412
rect 33140 7372 37900 7412
rect 37940 7372 37949 7412
rect 10723 7288 10732 7328
rect 10772 7288 13132 7328
rect 13172 7288 13181 7328
rect 16291 7288 16300 7328
rect 16340 7288 18604 7328
rect 18644 7288 18653 7328
rect 18883 7288 18892 7328
rect 18932 7288 27148 7328
rect 27188 7288 27197 7328
rect 27331 7288 27340 7328
rect 27380 7288 29068 7328
rect 29108 7288 29117 7328
rect 34339 7288 34348 7328
rect 34388 7288 40108 7328
rect 40148 7288 40157 7328
rect 10627 7204 10636 7244
rect 10676 7204 11020 7244
rect 11060 7204 11069 7244
rect 12845 7204 12940 7244
rect 12980 7204 12989 7244
rect 17635 7204 17644 7244
rect 17684 7204 22004 7244
rect 22531 7204 22540 7244
rect 22580 7204 24652 7244
rect 24692 7204 24701 7244
rect 25891 7204 25900 7244
rect 25940 7204 33292 7244
rect 33332 7204 33341 7244
rect 33955 7204 33964 7244
rect 34004 7204 37036 7244
rect 37076 7204 37085 7244
rect 15907 7120 15916 7160
rect 15956 7120 20180 7160
rect 20140 7076 20180 7120
rect 21964 7076 22004 7204
rect 22723 7120 22732 7160
rect 22772 7120 30412 7160
rect 30452 7120 30461 7160
rect 33283 7120 33292 7160
rect 33332 7120 33341 7160
rect 34147 7120 34156 7160
rect 34196 7120 36748 7160
rect 36788 7120 38668 7160
rect 38708 7120 38717 7160
rect 33292 7076 33332 7120
rect 11011 7036 11020 7076
rect 11060 7036 16492 7076
rect 16532 7036 16541 7076
rect 18883 7036 18892 7076
rect 18932 7036 19756 7076
rect 19796 7036 19805 7076
rect 20131 7036 20140 7076
rect 20180 7036 20189 7076
rect 21964 7036 23212 7076
rect 23252 7036 23261 7076
rect 29645 7036 29740 7076
rect 29780 7036 29789 7076
rect 32899 7036 32908 7076
rect 32948 7036 33332 7076
rect 33379 7036 33388 7076
rect 33428 7036 33676 7076
rect 33716 7036 33868 7076
rect 33908 7036 33917 7076
rect 4291 6952 4300 6992
rect 4340 6952 43276 6992
rect 43316 6952 43325 6992
rect 7939 6868 7948 6908
rect 7988 6868 21580 6908
rect 21620 6868 21629 6908
rect 21763 6868 21772 6908
rect 21812 6868 25324 6908
rect 25364 6868 25373 6908
rect 29827 6868 29836 6908
rect 29876 6868 30028 6908
rect 30068 6868 30077 6908
rect 31459 6868 31468 6908
rect 31508 6868 33580 6908
rect 33620 6868 33629 6908
rect 33676 6868 37324 6908
rect 37364 6868 37373 6908
rect 33676 6824 33716 6868
rect 3679 6784 3688 6824
rect 3728 6784 3770 6824
rect 3810 6784 3852 6824
rect 3892 6784 3934 6824
rect 3974 6784 4016 6824
rect 4056 6784 4065 6824
rect 12931 6784 12940 6824
rect 12980 6784 13996 6824
rect 14036 6784 14045 6824
rect 18799 6784 18808 6824
rect 18848 6784 18890 6824
rect 18930 6784 18972 6824
rect 19012 6784 19054 6824
rect 19094 6784 19136 6824
rect 19176 6784 19185 6824
rect 19459 6784 19468 6824
rect 19508 6784 23060 6824
rect 29731 6784 29740 6824
rect 29780 6784 30316 6824
rect 30356 6784 30365 6824
rect 32611 6784 32620 6824
rect 32660 6784 33716 6824
rect 33919 6784 33928 6824
rect 33968 6784 34010 6824
rect 34050 6784 34092 6824
rect 34132 6784 34174 6824
rect 34214 6784 34256 6824
rect 34296 6784 34305 6824
rect 23020 6740 23060 6784
rect 11107 6700 11116 6740
rect 11156 6700 11596 6740
rect 11636 6700 11645 6740
rect 12739 6700 12748 6740
rect 12788 6700 19276 6740
rect 19316 6700 19325 6740
rect 23020 6700 36844 6740
rect 36884 6700 36893 6740
rect 13421 6616 13516 6656
rect 13556 6616 13565 6656
rect 14755 6616 14764 6656
rect 14804 6616 43084 6656
rect 43124 6616 43133 6656
rect 10243 6532 10252 6572
rect 10292 6532 10732 6572
rect 10772 6532 10781 6572
rect 12259 6532 12268 6572
rect 12308 6532 27340 6572
rect 27380 6532 27389 6572
rect 29731 6532 29740 6572
rect 29780 6532 29836 6572
rect 29876 6532 29885 6572
rect 32707 6532 32716 6572
rect 32756 6532 36364 6572
rect 36404 6532 36413 6572
rect 6403 6448 6412 6488
rect 6452 6448 6700 6488
rect 6740 6448 31276 6488
rect 31316 6448 31325 6488
rect 32803 6448 32812 6488
rect 32852 6448 34924 6488
rect 34964 6448 34973 6488
rect 4195 6364 4204 6404
rect 4244 6364 37132 6404
rect 37172 6364 38188 6404
rect 38228 6364 38237 6404
rect 5731 6280 5740 6320
rect 5780 6280 6796 6320
rect 6836 6280 35692 6320
rect 35732 6280 35741 6320
rect 11875 6196 11884 6236
rect 11924 6196 41740 6236
rect 41780 6196 41789 6236
rect 10243 6112 10252 6152
rect 10292 6112 13324 6152
rect 13364 6112 13373 6152
rect 18019 6112 18028 6152
rect 18068 6112 29836 6152
rect 29876 6112 29885 6152
rect 33187 6112 33196 6152
rect 33236 6112 33388 6152
rect 33428 6112 33437 6152
rect 4919 6028 4928 6068
rect 4968 6028 5010 6068
rect 5050 6028 5092 6068
rect 5132 6028 5174 6068
rect 5214 6028 5256 6068
rect 5296 6028 5305 6068
rect 11203 6028 11212 6068
rect 11252 6028 11884 6068
rect 11924 6028 12460 6068
rect 12500 6028 12509 6068
rect 12643 6028 12652 6068
rect 12692 6028 13996 6068
rect 14036 6028 14045 6068
rect 15139 6028 15148 6068
rect 15188 6028 19604 6068
rect 20039 6028 20048 6068
rect 20088 6028 20130 6068
rect 20170 6028 20212 6068
rect 20252 6028 20294 6068
rect 20334 6028 20376 6068
rect 20416 6028 20425 6068
rect 23395 6028 23404 6068
rect 23444 6028 28780 6068
rect 28820 6028 28829 6068
rect 35159 6028 35168 6068
rect 35208 6028 35250 6068
rect 35290 6028 35332 6068
rect 35372 6028 35414 6068
rect 35454 6028 35496 6068
rect 35536 6028 35545 6068
rect 19564 5984 19604 6028
rect 12739 5944 12748 5984
rect 12788 5944 19508 5984
rect 19564 5944 20812 5984
rect 20852 5944 20861 5984
rect 22915 5944 22924 5984
rect 22964 5944 28972 5984
rect 29012 5944 29021 5984
rect 12931 5860 12940 5900
rect 12980 5860 13996 5900
rect 14036 5860 14045 5900
rect 15811 5860 15820 5900
rect 15860 5860 18700 5900
rect 18740 5860 18749 5900
rect 19468 5816 19508 5944
rect 23395 5860 23404 5900
rect 23444 5860 25708 5900
rect 25748 5860 25757 5900
rect 31843 5860 31852 5900
rect 31892 5860 36556 5900
rect 36596 5860 36605 5900
rect 11491 5776 11500 5816
rect 11540 5776 13900 5816
rect 13940 5776 13949 5816
rect 19468 5776 20044 5816
rect 20084 5776 20093 5816
rect 22819 5776 22828 5816
rect 22868 5776 23020 5816
rect 23060 5776 23069 5816
rect 31747 5776 31756 5816
rect 31796 5776 34828 5816
rect 34868 5776 34877 5816
rect 11299 5692 11308 5732
rect 11348 5692 35020 5732
rect 35060 5692 35069 5732
rect 11971 5608 11980 5648
rect 12020 5608 36460 5648
rect 36500 5608 36509 5648
rect 12912 5524 12940 5564
rect 12980 5524 13036 5564
rect 13076 5524 13900 5564
rect 13940 5524 13949 5564
rect 15619 5524 15628 5564
rect 15668 5524 43468 5564
rect 43508 5524 43517 5564
rect 8899 5440 8908 5480
rect 8948 5440 35980 5480
rect 36020 5440 36029 5480
rect 18595 5356 18604 5396
rect 18644 5356 19276 5396
rect 19316 5356 19325 5396
rect 23203 5356 23212 5396
rect 23252 5356 24172 5396
rect 24212 5356 24221 5396
rect 32995 5356 33004 5396
rect 33044 5356 36172 5396
rect 36212 5356 36221 5396
rect 3679 5272 3688 5312
rect 3728 5272 3770 5312
rect 3810 5272 3852 5312
rect 3892 5272 3934 5312
rect 3974 5272 4016 5312
rect 4056 5272 4065 5312
rect 12739 5272 12748 5312
rect 12788 5272 14572 5312
rect 14612 5272 14621 5312
rect 18799 5272 18808 5312
rect 18848 5272 18890 5312
rect 18930 5272 18972 5312
rect 19012 5272 19054 5312
rect 19094 5272 19136 5312
rect 19176 5272 19185 5312
rect 33919 5272 33928 5312
rect 33968 5272 34010 5312
rect 34050 5272 34092 5312
rect 34132 5272 34174 5312
rect 34214 5272 34256 5312
rect 34296 5272 34305 5312
rect 14179 5188 14188 5228
rect 14228 5188 21580 5228
rect 21620 5188 21629 5228
rect 11683 5104 11692 5144
rect 11732 5104 34540 5144
rect 34580 5104 34589 5144
rect 17059 5020 17068 5060
rect 17108 5020 32428 5060
rect 32468 5020 32477 5060
rect 33091 5020 33100 5060
rect 33140 5020 35116 5060
rect 35156 5020 35165 5060
rect 23683 4936 23692 4976
rect 23732 4936 24268 4976
rect 24308 4936 24317 4976
rect 28867 4936 28876 4976
rect 28916 4936 29740 4976
rect 29780 4936 29789 4976
rect 32803 4936 32812 4976
rect 32852 4936 33676 4976
rect 33716 4936 37900 4976
rect 37940 4936 37949 4976
rect 4387 4852 4396 4892
rect 4436 4852 7564 4892
rect 7604 4852 7613 4892
rect 22915 4852 22924 4892
rect 22964 4852 24076 4892
rect 24116 4852 24556 4892
rect 24596 4852 24605 4892
rect 9475 4768 9484 4808
rect 9524 4768 33676 4808
rect 33716 4768 33725 4808
rect 12163 4684 12172 4724
rect 12212 4684 44908 4724
rect 44948 4684 44957 4724
rect 33197 4600 33292 4640
rect 33332 4600 33341 4640
rect 41155 4600 41164 4640
rect 41204 4600 41548 4640
rect 41588 4600 41597 4640
rect 4919 4516 4928 4556
rect 4968 4516 5010 4556
rect 5050 4516 5092 4556
rect 5132 4516 5174 4556
rect 5214 4516 5256 4556
rect 5296 4516 5305 4556
rect 10915 4516 10924 4556
rect 10964 4516 18796 4556
rect 18836 4516 18845 4556
rect 20039 4516 20048 4556
rect 20088 4516 20130 4556
rect 20170 4516 20212 4556
rect 20252 4516 20294 4556
rect 20334 4516 20376 4556
rect 20416 4516 20425 4556
rect 23587 4516 23596 4556
rect 23636 4516 30124 4556
rect 30164 4516 30173 4556
rect 35159 4516 35168 4556
rect 35208 4516 35250 4556
rect 35290 4516 35332 4556
rect 35372 4516 35414 4556
rect 35454 4516 35496 4556
rect 35536 4516 35545 4556
rect 10723 4432 10732 4472
rect 10772 4432 16492 4472
rect 16532 4432 16541 4472
rect 19747 4432 19756 4472
rect 19796 4432 23116 4472
rect 23156 4432 23165 4472
rect 23692 4432 26188 4472
rect 26228 4432 26237 4472
rect 32899 4432 32908 4472
rect 32948 4432 39244 4472
rect 39284 4432 39293 4472
rect 23692 4388 23732 4432
rect 14659 4348 14668 4388
rect 14708 4348 15628 4388
rect 15668 4348 15677 4388
rect 22243 4348 22252 4388
rect 22292 4348 23732 4388
rect 23779 4348 23788 4388
rect 23828 4348 24268 4388
rect 24308 4348 24317 4388
rect 7939 4264 7948 4304
rect 7988 4264 9196 4304
rect 9236 4264 9245 4304
rect 12259 4264 12268 4304
rect 12308 4264 18124 4304
rect 18164 4264 18173 4304
rect 24931 4264 24940 4304
rect 24980 4264 28876 4304
rect 28916 4264 29260 4304
rect 29300 4264 29309 4304
rect 31075 4264 31084 4304
rect 31124 4264 38572 4304
rect 38612 4264 38956 4304
rect 38996 4264 39005 4304
rect 10051 4180 10060 4220
rect 10100 4180 32140 4220
rect 32180 4180 32189 4220
rect 13507 4096 13516 4136
rect 13556 4096 44524 4136
rect 44564 4096 44573 4136
rect 13699 4012 13708 4052
rect 13748 4012 15628 4052
rect 15668 4012 15677 4052
rect 17923 4012 17932 4052
rect 17972 4012 20140 4052
rect 20180 4012 20189 4052
rect 38467 4012 38476 4052
rect 38516 4012 39532 4052
rect 39572 4012 39581 4052
rect 12835 3928 12844 3968
rect 12884 3928 41740 3968
rect 41780 3928 41789 3968
rect 13219 3844 13228 3884
rect 13268 3844 17548 3884
rect 17588 3844 17597 3884
rect 31843 3844 31852 3884
rect 31892 3844 32332 3884
rect 32372 3844 32381 3884
rect 3679 3760 3688 3800
rect 3728 3760 3770 3800
rect 3810 3760 3852 3800
rect 3892 3760 3934 3800
rect 3974 3760 4016 3800
rect 4056 3760 4065 3800
rect 13699 3760 13708 3800
rect 13748 3760 14188 3800
rect 14228 3760 14237 3800
rect 18799 3760 18808 3800
rect 18848 3760 18890 3800
rect 18930 3760 18972 3800
rect 19012 3760 19054 3800
rect 19094 3760 19136 3800
rect 19176 3760 19185 3800
rect 20803 3760 20812 3800
rect 20852 3760 29644 3800
rect 29684 3760 29693 3800
rect 33919 3760 33928 3800
rect 33968 3760 34010 3800
rect 34050 3760 34092 3800
rect 34132 3760 34174 3800
rect 34214 3760 34256 3800
rect 34296 3760 34305 3800
rect 13411 3676 13420 3716
rect 13460 3676 24748 3716
rect 24788 3676 24797 3716
rect 12355 3592 12364 3632
rect 12404 3592 17932 3632
rect 17972 3592 17981 3632
rect 18787 3592 18796 3632
rect 18836 3592 21196 3632
rect 21236 3592 21245 3632
rect 21955 3592 21964 3632
rect 22004 3592 29548 3632
rect 29588 3592 29597 3632
rect 7459 3508 7468 3548
rect 7508 3508 25228 3548
rect 25268 3508 25277 3548
rect 28675 3508 28684 3548
rect 28724 3508 30220 3548
rect 30260 3508 30269 3548
rect 9571 3424 9580 3464
rect 9620 3424 9868 3464
rect 9908 3424 9917 3464
rect 12451 3424 12460 3464
rect 12500 3424 12940 3464
rect 12980 3424 12989 3464
rect 13411 3424 13420 3464
rect 13460 3424 16204 3464
rect 16244 3424 35884 3464
rect 35924 3424 35933 3464
rect 1891 3340 1900 3380
rect 1940 3340 25996 3380
rect 26036 3340 26380 3380
rect 26420 3340 26429 3380
rect 13795 3256 13804 3296
rect 13844 3256 33676 3296
rect 33716 3256 33725 3296
rect 16291 3172 16300 3212
rect 16340 3172 39820 3212
rect 39860 3172 39869 3212
rect 11971 3088 11980 3128
rect 12020 3088 22924 3128
rect 22964 3088 22973 3128
rect 4919 3004 4928 3044
rect 4968 3004 5010 3044
rect 5050 3004 5092 3044
rect 5132 3004 5174 3044
rect 5214 3004 5256 3044
rect 5296 3004 5305 3044
rect 15331 3004 15340 3044
rect 15380 3004 15628 3044
rect 15668 3004 15677 3044
rect 20039 3004 20048 3044
rect 20088 3004 20130 3044
rect 20170 3004 20212 3044
rect 20252 3004 20294 3044
rect 20334 3004 20376 3044
rect 20416 3004 20425 3044
rect 35159 3004 35168 3044
rect 35208 3004 35250 3044
rect 35290 3004 35332 3044
rect 35372 3004 35414 3044
rect 35454 3004 35496 3044
rect 35536 3004 35545 3044
rect 12931 2920 12940 2960
rect 12980 2920 13132 2960
rect 13172 2920 13181 2960
rect 17251 2920 17260 2960
rect 17300 2920 18508 2960
rect 18548 2920 19468 2960
rect 19508 2920 19517 2960
rect 20899 2920 20908 2960
rect 20948 2920 25228 2960
rect 25268 2920 25277 2960
rect 13219 2836 13228 2876
rect 13268 2836 21100 2876
rect 21140 2836 21149 2876
rect 21283 2836 21292 2876
rect 21332 2836 33100 2876
rect 33140 2836 33149 2876
rect 37891 2836 37900 2876
rect 37940 2836 42028 2876
rect 42068 2836 42077 2876
rect 17635 2752 17644 2792
rect 17684 2752 35500 2792
rect 35540 2752 35549 2792
rect 4675 2668 4684 2708
rect 4724 2668 9772 2708
rect 9812 2668 24268 2708
rect 24308 2668 24317 2708
rect 24547 2668 24556 2708
rect 24596 2668 25516 2708
rect 25556 2668 25565 2708
rect 27523 2668 27532 2708
rect 27572 2668 29740 2708
rect 29780 2668 29789 2708
rect 8899 2584 8908 2624
rect 8948 2584 15148 2624
rect 15188 2584 16204 2624
rect 16244 2584 16253 2624
rect 18307 2584 18316 2624
rect 18356 2584 38956 2624
rect 38996 2584 39005 2624
rect 2851 2500 2860 2540
rect 2900 2500 36172 2540
rect 36212 2500 36221 2540
rect 2083 2416 2092 2456
rect 2132 2416 40300 2456
rect 40340 2416 40349 2456
rect 43651 2416 43660 2456
rect 43700 2416 44620 2456
rect 44660 2416 44669 2456
rect 8419 2332 8428 2372
rect 8468 2332 11212 2372
rect 11252 2332 11261 2372
rect 14467 2332 14476 2372
rect 14516 2332 21292 2372
rect 21332 2332 21341 2372
rect 24259 2332 24268 2372
rect 24308 2332 31852 2372
rect 31892 2332 31901 2372
rect 3679 2248 3688 2288
rect 3728 2248 3770 2288
rect 3810 2248 3852 2288
rect 3892 2248 3934 2288
rect 3974 2248 4016 2288
rect 4056 2248 4065 2288
rect 18799 2248 18808 2288
rect 18848 2248 18890 2288
rect 18930 2248 18972 2288
rect 19012 2248 19054 2288
rect 19094 2248 19136 2288
rect 19176 2248 19185 2288
rect 20035 2248 20044 2288
rect 20084 2248 21868 2288
rect 21908 2248 22252 2288
rect 22292 2248 22301 2288
rect 22723 2248 22732 2288
rect 22772 2248 23212 2288
rect 23252 2248 23261 2288
rect 33919 2248 33928 2288
rect 33968 2248 34010 2288
rect 34050 2248 34092 2288
rect 34132 2248 34174 2288
rect 34214 2248 34256 2288
rect 34296 2248 34305 2288
rect 38659 2248 38668 2288
rect 38708 2248 40300 2288
rect 40340 2248 40349 2288
rect 12643 2164 12652 2204
rect 12692 2164 19948 2204
rect 19988 2164 19997 2204
rect 23011 2164 23020 2204
rect 23060 2164 25132 2204
rect 25172 2164 25181 2204
rect 37219 2164 37228 2204
rect 37268 2164 37900 2204
rect 37940 2164 37949 2204
rect 12931 2080 12940 2120
rect 12980 2080 13900 2120
rect 13940 2080 13949 2120
rect 22627 2080 22636 2120
rect 22676 2080 29452 2120
rect 29492 2080 29501 2120
rect 12739 1996 12748 2036
rect 12788 1996 12940 2036
rect 12980 1996 12989 2036
rect 16195 1996 16204 2036
rect 16244 1996 17932 2036
rect 17972 1996 17981 2036
rect 18403 1996 18412 2036
rect 18452 1996 23692 2036
rect 23732 1996 23741 2036
rect 15427 1912 15436 1952
rect 15476 1912 21004 1952
rect 21044 1912 21053 1952
rect 32131 1912 32140 1952
rect 32180 1912 35692 1952
rect 35732 1912 35741 1952
rect 14083 1828 14092 1868
rect 14132 1828 21772 1868
rect 21812 1828 21821 1868
rect 11971 1744 11980 1784
rect 12020 1744 33676 1784
rect 33716 1744 33725 1784
rect 34435 1744 34444 1784
rect 34484 1744 40396 1784
rect 40436 1744 40445 1784
rect 11491 1660 11500 1700
rect 11540 1660 40876 1700
rect 40916 1660 40925 1700
rect 15619 1576 15628 1616
rect 15668 1576 20524 1616
rect 20564 1576 20573 1616
rect 4919 1492 4928 1532
rect 4968 1492 5010 1532
rect 5050 1492 5092 1532
rect 5132 1492 5174 1532
rect 5214 1492 5256 1532
rect 5296 1492 5305 1532
rect 13315 1492 13324 1532
rect 13364 1492 14476 1532
rect 14516 1492 14525 1532
rect 20039 1492 20048 1532
rect 20088 1492 20130 1532
rect 20170 1492 20212 1532
rect 20252 1492 20294 1532
rect 20334 1492 20376 1532
rect 20416 1492 20425 1532
rect 23299 1492 23308 1532
rect 23348 1492 26284 1532
rect 26324 1492 26333 1532
rect 35159 1492 35168 1532
rect 35208 1492 35250 1532
rect 35290 1492 35332 1532
rect 35372 1492 35414 1532
rect 35454 1492 35496 1532
rect 35536 1492 35545 1532
rect 38659 1492 38668 1532
rect 38708 1492 38956 1532
rect 38996 1492 39005 1532
rect 30787 988 30796 1028
rect 30836 988 39052 1028
rect 39092 988 39101 1028
rect 19939 820 19948 860
rect 19988 820 20812 860
rect 20852 820 20861 860
rect 33100 148 39340 188
rect 39380 148 39389 188
rect 33100 104 33140 148
rect 33091 64 33100 104
rect 33140 64 33149 104
rect 33859 64 33868 104
rect 33908 64 34060 104
rect 34100 64 34109 104
rect 41251 64 41260 104
rect 41300 64 41548 104
rect 41588 64 41597 104
<< via4 >>
rect 19852 10060 19892 10100
rect 3688 9808 3728 9848
rect 3770 9808 3810 9848
rect 3852 9808 3892 9848
rect 3934 9808 3974 9848
rect 4016 9808 4056 9848
rect 18808 9808 18848 9848
rect 18890 9808 18930 9848
rect 18972 9808 19012 9848
rect 19054 9808 19094 9848
rect 19136 9808 19176 9848
rect 33928 9808 33968 9848
rect 34010 9808 34050 9848
rect 34092 9808 34132 9848
rect 34174 9808 34214 9848
rect 34256 9808 34296 9848
rect 20524 9304 20564 9344
rect 4928 9052 4968 9092
rect 5010 9052 5050 9092
rect 5092 9052 5132 9092
rect 5174 9052 5214 9092
rect 5256 9052 5296 9092
rect 20048 9052 20088 9092
rect 20130 9052 20170 9092
rect 20212 9052 20252 9092
rect 20294 9052 20334 9092
rect 20376 9052 20416 9092
rect 33388 9052 33428 9092
rect 35168 9052 35208 9092
rect 35250 9052 35290 9092
rect 35332 9052 35372 9092
rect 35414 9052 35454 9092
rect 35496 9052 35536 9092
rect 33196 8800 33236 8840
rect 33388 8464 33428 8504
rect 20524 8380 20564 8420
rect 3688 8296 3728 8336
rect 3770 8296 3810 8336
rect 3852 8296 3892 8336
rect 3934 8296 3974 8336
rect 4016 8296 4056 8336
rect 18808 8296 18848 8336
rect 18890 8296 18930 8336
rect 18972 8296 19012 8336
rect 19054 8296 19094 8336
rect 19136 8296 19176 8336
rect 20908 8296 20948 8336
rect 33928 8296 33968 8336
rect 34010 8296 34050 8336
rect 34092 8296 34132 8336
rect 34174 8296 34214 8336
rect 34256 8296 34296 8336
rect 19468 8044 19508 8084
rect 13036 7792 13076 7832
rect 4928 7540 4968 7580
rect 5010 7540 5050 7580
rect 5092 7540 5132 7580
rect 5174 7540 5214 7580
rect 5256 7540 5296 7580
rect 20048 7540 20088 7580
rect 20130 7540 20170 7580
rect 20212 7540 20252 7580
rect 20294 7540 20334 7580
rect 20376 7540 20416 7580
rect 35168 7540 35208 7580
rect 35250 7540 35290 7580
rect 35332 7540 35372 7580
rect 35414 7540 35454 7580
rect 35496 7540 35536 7580
rect 19852 7372 19892 7412
rect 12940 7204 12980 7244
rect 33292 7204 33332 7244
rect 29740 7036 29780 7076
rect 3688 6784 3728 6824
rect 3770 6784 3810 6824
rect 3852 6784 3892 6824
rect 3934 6784 3974 6824
rect 4016 6784 4056 6824
rect 18808 6784 18848 6824
rect 18890 6784 18930 6824
rect 18972 6784 19012 6824
rect 19054 6784 19094 6824
rect 19136 6784 19176 6824
rect 19468 6784 19508 6824
rect 33928 6784 33968 6824
rect 34010 6784 34050 6824
rect 34092 6784 34132 6824
rect 34174 6784 34214 6824
rect 34256 6784 34296 6824
rect 13516 6616 13556 6656
rect 29740 6532 29780 6572
rect 33196 6112 33236 6152
rect 4928 6028 4968 6068
rect 5010 6028 5050 6068
rect 5092 6028 5132 6068
rect 5174 6028 5214 6068
rect 5256 6028 5296 6068
rect 20048 6028 20088 6068
rect 20130 6028 20170 6068
rect 20212 6028 20252 6068
rect 20294 6028 20334 6068
rect 20376 6028 20416 6068
rect 35168 6028 35208 6068
rect 35250 6028 35290 6068
rect 35332 6028 35372 6068
rect 35414 6028 35454 6068
rect 35496 6028 35536 6068
rect 13036 5524 13076 5564
rect 3688 5272 3728 5312
rect 3770 5272 3810 5312
rect 3852 5272 3892 5312
rect 3934 5272 3974 5312
rect 4016 5272 4056 5312
rect 18808 5272 18848 5312
rect 18890 5272 18930 5312
rect 18972 5272 19012 5312
rect 19054 5272 19094 5312
rect 19136 5272 19176 5312
rect 33928 5272 33968 5312
rect 34010 5272 34050 5312
rect 34092 5272 34132 5312
rect 34174 5272 34214 5312
rect 34256 5272 34296 5312
rect 33292 4600 33332 4640
rect 4928 4516 4968 4556
rect 5010 4516 5050 4556
rect 5092 4516 5132 4556
rect 5174 4516 5214 4556
rect 5256 4516 5296 4556
rect 20048 4516 20088 4556
rect 20130 4516 20170 4556
rect 20212 4516 20252 4556
rect 20294 4516 20334 4556
rect 20376 4516 20416 4556
rect 35168 4516 35208 4556
rect 35250 4516 35290 4556
rect 35332 4516 35372 4556
rect 35414 4516 35454 4556
rect 35496 4516 35536 4556
rect 13516 4096 13556 4136
rect 3688 3760 3728 3800
rect 3770 3760 3810 3800
rect 3852 3760 3892 3800
rect 3934 3760 3974 3800
rect 4016 3760 4056 3800
rect 18808 3760 18848 3800
rect 18890 3760 18930 3800
rect 18972 3760 19012 3800
rect 19054 3760 19094 3800
rect 19136 3760 19176 3800
rect 33928 3760 33968 3800
rect 34010 3760 34050 3800
rect 34092 3760 34132 3800
rect 34174 3760 34214 3800
rect 34256 3760 34296 3800
rect 4928 3004 4968 3044
rect 5010 3004 5050 3044
rect 5092 3004 5132 3044
rect 5174 3004 5214 3044
rect 5256 3004 5296 3044
rect 20048 3004 20088 3044
rect 20130 3004 20170 3044
rect 20212 3004 20252 3044
rect 20294 3004 20334 3044
rect 20376 3004 20416 3044
rect 35168 3004 35208 3044
rect 35250 3004 35290 3044
rect 35332 3004 35372 3044
rect 35414 3004 35454 3044
rect 35496 3004 35536 3044
rect 20908 2920 20948 2960
rect 3688 2248 3728 2288
rect 3770 2248 3810 2288
rect 3852 2248 3892 2288
rect 3934 2248 3974 2288
rect 4016 2248 4056 2288
rect 18808 2248 18848 2288
rect 18890 2248 18930 2288
rect 18972 2248 19012 2288
rect 19054 2248 19094 2288
rect 19136 2248 19176 2288
rect 33928 2248 33968 2288
rect 34010 2248 34050 2288
rect 34092 2248 34132 2288
rect 34174 2248 34214 2288
rect 34256 2248 34296 2288
rect 12940 2080 12980 2120
rect 4928 1492 4968 1532
rect 5010 1492 5050 1532
rect 5092 1492 5132 1532
rect 5174 1492 5214 1532
rect 5256 1492 5296 1532
rect 20048 1492 20088 1532
rect 20130 1492 20170 1532
rect 20212 1492 20252 1532
rect 20294 1492 20334 1532
rect 20376 1492 20416 1532
rect 35168 1492 35208 1532
rect 35250 1492 35290 1532
rect 35332 1492 35372 1532
rect 35414 1492 35454 1532
rect 35496 1492 35536 1532
<< metal5 >>
rect 3652 9848 4092 11844
rect 3652 9808 3688 9848
rect 3728 9808 3770 9848
rect 3810 9808 3852 9848
rect 3892 9808 3934 9848
rect 3974 9808 4016 9848
rect 4056 9808 4092 9848
rect 3652 8336 4092 9808
rect 3652 8296 3688 8336
rect 3728 8296 3770 8336
rect 3810 8296 3852 8336
rect 3892 8296 3934 8336
rect 3974 8296 4016 8336
rect 4056 8296 4092 8336
rect 3652 6824 4092 8296
rect 3652 6784 3688 6824
rect 3728 6784 3770 6824
rect 3810 6784 3852 6824
rect 3892 6784 3934 6824
rect 3974 6784 4016 6824
rect 4056 6784 4092 6824
rect 3652 5312 4092 6784
rect 3652 5272 3688 5312
rect 3728 5272 3770 5312
rect 3810 5272 3852 5312
rect 3892 5272 3934 5312
rect 3974 5272 4016 5312
rect 4056 5272 4092 5312
rect 3652 3800 4092 5272
rect 3652 3760 3688 3800
rect 3728 3760 3770 3800
rect 3810 3760 3852 3800
rect 3892 3760 3934 3800
rect 3974 3760 4016 3800
rect 4056 3760 4092 3800
rect 3652 2288 4092 3760
rect 3652 2248 3688 2288
rect 3728 2248 3770 2288
rect 3810 2248 3852 2288
rect 3892 2248 3934 2288
rect 3974 2248 4016 2288
rect 4056 2248 4092 2288
rect 3652 0 4092 2248
rect 4892 9092 5332 11844
rect 4892 9052 4928 9092
rect 4968 9052 5010 9092
rect 5050 9052 5092 9092
rect 5132 9052 5174 9092
rect 5214 9052 5256 9092
rect 5296 9052 5332 9092
rect 4892 7580 5332 9052
rect 18772 9848 19212 11844
rect 18772 9808 18808 9848
rect 18848 9808 18890 9848
rect 18930 9808 18972 9848
rect 19012 9808 19054 9848
rect 19094 9808 19136 9848
rect 19176 9808 19212 9848
rect 18772 8336 19212 9808
rect 18772 8296 18808 8336
rect 18848 8296 18890 8336
rect 18930 8296 18972 8336
rect 19012 8296 19054 8336
rect 19094 8296 19136 8336
rect 19176 8296 19212 8336
rect 4892 7540 4928 7580
rect 4968 7540 5010 7580
rect 5050 7540 5092 7580
rect 5132 7540 5174 7580
rect 5214 7540 5256 7580
rect 5296 7540 5332 7580
rect 4892 6068 5332 7540
rect 13036 7832 13076 7841
rect 4892 6028 4928 6068
rect 4968 6028 5010 6068
rect 5050 6028 5092 6068
rect 5132 6028 5174 6068
rect 5214 6028 5256 6068
rect 5296 6028 5332 6068
rect 4892 4556 5332 6028
rect 4892 4516 4928 4556
rect 4968 4516 5010 4556
rect 5050 4516 5092 4556
rect 5132 4516 5174 4556
rect 5214 4516 5256 4556
rect 5296 4516 5332 4556
rect 4892 3044 5332 4516
rect 4892 3004 4928 3044
rect 4968 3004 5010 3044
rect 5050 3004 5092 3044
rect 5132 3004 5174 3044
rect 5214 3004 5256 3044
rect 5296 3004 5332 3044
rect 4892 1532 5332 3004
rect 12940 7244 12980 7253
rect 12940 2120 12980 7204
rect 13036 5564 13076 7792
rect 18772 6824 19212 8296
rect 19852 10100 19892 10109
rect 18772 6784 18808 6824
rect 18848 6784 18890 6824
rect 18930 6784 18972 6824
rect 19012 6784 19054 6824
rect 19094 6784 19136 6824
rect 19176 6784 19212 6824
rect 13036 5515 13076 5524
rect 13516 6656 13556 6665
rect 13516 4136 13556 6616
rect 13516 4087 13556 4096
rect 18772 5312 19212 6784
rect 19468 8084 19508 8093
rect 19468 6824 19508 8044
rect 19852 7412 19892 10060
rect 19852 7363 19892 7372
rect 20012 9092 20452 11844
rect 33892 9848 34332 11844
rect 33892 9808 33928 9848
rect 33968 9808 34010 9848
rect 34050 9808 34092 9848
rect 34132 9808 34174 9848
rect 34214 9808 34256 9848
rect 34296 9808 34332 9848
rect 20012 9052 20048 9092
rect 20088 9052 20130 9092
rect 20170 9052 20212 9092
rect 20252 9052 20294 9092
rect 20334 9052 20376 9092
rect 20416 9052 20452 9092
rect 20012 7580 20452 9052
rect 20524 9344 20564 9353
rect 20524 8420 20564 9304
rect 33388 9092 33428 9101
rect 20524 8371 20564 8380
rect 33196 8840 33236 8849
rect 20012 7540 20048 7580
rect 20088 7540 20130 7580
rect 20170 7540 20212 7580
rect 20252 7540 20294 7580
rect 20334 7540 20376 7580
rect 20416 7540 20452 7580
rect 19468 6775 19508 6784
rect 18772 5272 18808 5312
rect 18848 5272 18890 5312
rect 18930 5272 18972 5312
rect 19012 5272 19054 5312
rect 19094 5272 19136 5312
rect 19176 5272 19212 5312
rect 12940 2071 12980 2080
rect 18772 3800 19212 5272
rect 18772 3760 18808 3800
rect 18848 3760 18890 3800
rect 18930 3760 18972 3800
rect 19012 3760 19054 3800
rect 19094 3760 19136 3800
rect 19176 3760 19212 3800
rect 18772 2288 19212 3760
rect 18772 2248 18808 2288
rect 18848 2248 18890 2288
rect 18930 2248 18972 2288
rect 19012 2248 19054 2288
rect 19094 2248 19136 2288
rect 19176 2248 19212 2288
rect 4892 1492 4928 1532
rect 4968 1492 5010 1532
rect 5050 1492 5092 1532
rect 5132 1492 5174 1532
rect 5214 1492 5256 1532
rect 5296 1492 5332 1532
rect 4892 0 5332 1492
rect 18772 0 19212 2248
rect 20012 6068 20452 7540
rect 20012 6028 20048 6068
rect 20088 6028 20130 6068
rect 20170 6028 20212 6068
rect 20252 6028 20294 6068
rect 20334 6028 20376 6068
rect 20416 6028 20452 6068
rect 20012 4556 20452 6028
rect 20012 4516 20048 4556
rect 20088 4516 20130 4556
rect 20170 4516 20212 4556
rect 20252 4516 20294 4556
rect 20334 4516 20376 4556
rect 20416 4516 20452 4556
rect 20012 3044 20452 4516
rect 20012 3004 20048 3044
rect 20088 3004 20130 3044
rect 20170 3004 20212 3044
rect 20252 3004 20294 3044
rect 20334 3004 20376 3044
rect 20416 3004 20452 3044
rect 20012 1532 20452 3004
rect 20908 8336 20948 8345
rect 20908 2960 20948 8296
rect 29740 7076 29780 7085
rect 29740 6572 29780 7036
rect 29740 6523 29780 6532
rect 33196 6152 33236 8800
rect 33388 8504 33428 9052
rect 33388 8455 33428 8464
rect 33892 8336 34332 9808
rect 33892 8296 33928 8336
rect 33968 8296 34010 8336
rect 34050 8296 34092 8336
rect 34132 8296 34174 8336
rect 34214 8296 34256 8336
rect 34296 8296 34332 8336
rect 33196 6103 33236 6112
rect 33292 7244 33332 7253
rect 33292 4640 33332 7204
rect 33292 4591 33332 4600
rect 33892 6824 34332 8296
rect 33892 6784 33928 6824
rect 33968 6784 34010 6824
rect 34050 6784 34092 6824
rect 34132 6784 34174 6824
rect 34214 6784 34256 6824
rect 34296 6784 34332 6824
rect 33892 5312 34332 6784
rect 33892 5272 33928 5312
rect 33968 5272 34010 5312
rect 34050 5272 34092 5312
rect 34132 5272 34174 5312
rect 34214 5272 34256 5312
rect 34296 5272 34332 5312
rect 20908 2911 20948 2920
rect 33892 3800 34332 5272
rect 33892 3760 33928 3800
rect 33968 3760 34010 3800
rect 34050 3760 34092 3800
rect 34132 3760 34174 3800
rect 34214 3760 34256 3800
rect 34296 3760 34332 3800
rect 20012 1492 20048 1532
rect 20088 1492 20130 1532
rect 20170 1492 20212 1532
rect 20252 1492 20294 1532
rect 20334 1492 20376 1532
rect 20416 1492 20452 1532
rect 20012 0 20452 1492
rect 33892 2288 34332 3760
rect 33892 2248 33928 2288
rect 33968 2248 34010 2288
rect 34050 2248 34092 2288
rect 34132 2248 34174 2288
rect 34214 2248 34256 2288
rect 34296 2248 34332 2288
rect 33892 0 34332 2248
rect 35132 9092 35572 11844
rect 35132 9052 35168 9092
rect 35208 9052 35250 9092
rect 35290 9052 35332 9092
rect 35372 9052 35414 9092
rect 35454 9052 35496 9092
rect 35536 9052 35572 9092
rect 35132 7580 35572 9052
rect 35132 7540 35168 7580
rect 35208 7540 35250 7580
rect 35290 7540 35332 7580
rect 35372 7540 35414 7580
rect 35454 7540 35496 7580
rect 35536 7540 35572 7580
rect 35132 6068 35572 7540
rect 35132 6028 35168 6068
rect 35208 6028 35250 6068
rect 35290 6028 35332 6068
rect 35372 6028 35414 6068
rect 35454 6028 35496 6068
rect 35536 6028 35572 6068
rect 35132 4556 35572 6028
rect 35132 4516 35168 4556
rect 35208 4516 35250 4556
rect 35290 4516 35332 4556
rect 35372 4516 35414 4556
rect 35454 4516 35496 4556
rect 35536 4516 35572 4556
rect 35132 3044 35572 4516
rect 35132 3004 35168 3044
rect 35208 3004 35250 3044
rect 35290 3004 35332 3044
rect 35372 3004 35414 3044
rect 35454 3004 35496 3044
rect 35536 3004 35572 3044
rect 35132 1532 35572 3004
rect 35132 1492 35168 1532
rect 35208 1492 35250 1532
rect 35290 1492 35332 1532
rect 35372 1492 35414 1532
rect 35454 1492 35496 1532
rect 35536 1492 35572 1532
rect 35132 0 35572 1492
use sg13g2_mux4_1  _000_
timestamp 1677257233
transform 1 0 22272 0 1 6048
box -48 -56 2064 834
use sg13g2_mux4_1  _001_
timestamp 1677257233
transform 1 0 34272 0 -1 7560
box -48 -56 2064 834
use sg13g2_mux4_1  _002_
timestamp 1677257233
transform 1 0 5568 0 1 6048
box -48 -56 2064 834
use sg13g2_mux4_1  _003_
timestamp 1677257233
transform 1 0 14976 0 1 3024
box -48 -56 2064 834
use sg13g2_mux4_1  _004_
timestamp 1677257233
transform 1 0 27840 0 1 7560
box -48 -56 2064 834
use sg13g2_mux4_1  _005_
timestamp 1677257233
transform 1 0 38880 0 1 6048
box -48 -56 2064 834
use sg13g2_mux4_1  _006_
timestamp 1677257233
transform 1 0 8832 0 -1 9072
box -48 -56 2064 834
use sg13g2_mux4_1  _007_
timestamp 1677257233
transform 1 0 22944 0 -1 3024
box -48 -56 2064 834
use sg13g2_mux4_1  _008_
timestamp 1677257233
transform 1 0 18720 0 -1 9072
box -48 -56 2064 834
use sg13g2_mux4_1  _009_
timestamp 1677257233
transform 1 0 32448 0 -1 4536
box -48 -56 2064 834
use sg13g2_mux4_1  _010_
timestamp 1677257233
transform 1 0 10176 0 1 6048
box -48 -56 2064 834
use sg13g2_mux4_1  _011_
timestamp 1677257233
transform 1 0 19008 0 -1 3024
box -48 -56 2064 834
use sg13g2_mux4_1  _012_
timestamp 1677257233
transform 1 0 24384 0 -1 9072
box -48 -56 2064 834
use sg13g2_mux4_1  _013_
timestamp 1677257233
transform 1 0 37920 0 1 3024
box -48 -56 2064 834
use sg13g2_mux4_1  _014_
timestamp 1677257233
transform 1 0 6912 0 -1 4536
box -48 -56 2064 834
use sg13g2_mux4_1  _015_
timestamp 1677257233
transform 1 0 28128 0 -1 3024
box -48 -56 2064 834
use sg13g2_mux2_1  _016_
timestamp 1677247768
transform 1 0 28704 0 1 3024
box -48 -56 1008 834
use sg13g2_mux2_1  _017_
timestamp 1677247768
transform 1 0 9312 0 -1 4536
box -48 -56 1008 834
use sg13g2_mux2_1  _018_
timestamp 1677247768
transform 1 0 38208 0 -1 3024
box -48 -56 1008 834
use sg13g2_mux2_1  _019_
timestamp 1677247768
transform 1 0 26688 0 1 9072
box -48 -56 1008 834
use sg13g2_mux2_1  _020_
timestamp 1677247768
transform 1 0 18144 0 1 3024
box -48 -56 1008 834
use sg13g2_mux2_1  _021_
timestamp 1677247768
transform 1 0 9216 0 -1 7560
box -48 -56 1008 834
use sg13g2_mux2_1  _022_
timestamp 1677247768
transform 1 0 32928 0 1 4536
box -48 -56 1008 834
use sg13g2_mux2_1  _023_
timestamp 1677247768
transform 1 0 19296 0 1 9072
box -48 -56 1008 834
use sg13g2_mux2_1  _024_
timestamp 1677247768
transform -1 0 25920 0 -1 3024
box -48 -56 1008 834
use sg13g2_mux2_1  _025_
timestamp 1677247768
transform -1 0 11136 0 1 7560
box -48 -56 1008 834
use sg13g2_mux2_1  _026_
timestamp 1677247768
transform 1 0 40992 0 1 6048
box -48 -56 1008 834
use sg13g2_mux2_1  _027_
timestamp 1677247768
transform 1 0 33120 0 -1 9072
box -48 -56 1008 834
use sg13g2_mux2_1  _028_
timestamp 1677247768
transform 1 0 12960 0 1 3024
box -48 -56 1008 834
use sg13g2_mux2_1  _029_
timestamp 1677247768
transform 1 0 5280 0 1 4536
box -48 -56 1008 834
use sg13g2_mux2_1  _030_
timestamp 1677247768
transform 1 0 35136 0 1 7560
box -48 -56 1008 834
use sg13g2_mux2_1  _031_
timestamp 1677247768
transform 1 0 22848 0 -1 7560
box -48 -56 1008 834
use sg13g2_mux2_1  _032_
timestamp 1677247768
transform 1 0 27840 0 1 1512
box -48 -56 1008 834
use sg13g2_mux2_1  _033_
timestamp 1677247768
transform 1 0 7296 0 1 3024
box -48 -56 1008 834
use sg13g2_mux2_1  _034_
timestamp 1677247768
transform 1 0 34752 0 -1 3024
box -48 -56 1008 834
use sg13g2_mux2_1  _035_
timestamp 1677247768
transform 1 0 24384 0 1 9072
box -48 -56 1008 834
use sg13g2_mux2_1  _036_
timestamp 1677247768
transform 1 0 18048 0 -1 3024
box -48 -56 1008 834
use sg13g2_mux2_1  _037_
timestamp 1677247768
transform 1 0 10464 0 -1 7560
box -48 -56 1008 834
use sg13g2_mux2_1  _038_
timestamp 1677247768
transform 1 0 32640 0 1 3024
box -48 -56 1008 834
use sg13g2_mux2_1  _039_
timestamp 1677247768
transform 1 0 19200 0 1 7560
box -48 -56 1008 834
use sg13g2_mux2_1  _040_
timestamp 1677247768
transform 1 0 23808 0 1 3024
box -48 -56 1008 834
use sg13g2_mux2_1  _041_
timestamp 1677247768
transform -1 0 10944 0 1 9072
box -48 -56 1008 834
use sg13g2_mux2_1  _042_
timestamp 1677247768
transform 1 0 41952 0 1 6048
box -48 -56 1008 834
use sg13g2_mux2_1  _043_
timestamp 1677247768
transform 1 0 34752 0 1 9072
box -48 -56 1008 834
use sg13g2_mux2_1  _044_
timestamp 1677247768
transform -1 0 13920 0 -1 3024
box -48 -56 1008 834
use sg13g2_mux2_1  _045_
timestamp 1677247768
transform 1 0 6240 0 1 4536
box -48 -56 1008 834
use sg13g2_mux2_1  _046_
timestamp 1677247768
transform 1 0 34464 0 1 6048
box -48 -56 1008 834
use sg13g2_mux2_1  _047_
timestamp 1677247768
transform 1 0 23136 0 -1 6048
box -48 -56 1008 834
use sg13g2_mux2_1  _048_
timestamp 1677247768
transform 1 0 23808 0 1 1512
box -48 -56 1008 834
use sg13g2_mux2_1  _049_
timestamp 1677247768
transform 1 0 10560 0 -1 6048
box -48 -56 1008 834
use sg13g2_mux2_1  _050_
timestamp 1677247768
transform 1 0 40608 0 1 4536
box -48 -56 1008 834
use sg13g2_mux2_1  _051_
timestamp 1677247768
transform 1 0 34272 0 -1 9072
box -48 -56 1008 834
use sg13g2_mux2_1  _052_
timestamp 1677247768
transform 1 0 12960 0 1 1512
box -48 -56 1008 834
use sg13g2_mux2_1  _053_
timestamp 1677247768
transform -1 0 9216 0 1 9072
box -48 -56 1008 834
use sg13g2_mux2_1  _054_
timestamp 1677247768
transform 1 0 35712 0 1 6048
box -48 -56 1008 834
use sg13g2_mux2_1  _055_
timestamp 1677247768
transform 1 0 21984 0 1 7560
box -48 -56 1008 834
use sg13g2_mux2_1  _056_
timestamp 1677247768
transform 1 0 28800 0 1 1512
box -48 -56 1008 834
use sg13g2_mux2_1  _057_
timestamp 1677247768
transform -1 0 9408 0 -1 6048
box -48 -56 1008 834
use sg13g2_mux2_1  _058_
timestamp 1677247768
transform 1 0 38784 0 -1 4536
box -48 -56 1008 834
use sg13g2_mux2_1  _059_
timestamp 1677247768
transform 1 0 26688 0 -1 9072
box -48 -56 1008 834
use sg13g2_mux2_1  _060_
timestamp 1677247768
transform -1 0 15840 0 -1 4536
box -48 -56 1008 834
use sg13g2_mux2_1  _061_
timestamp 1677247768
transform 1 0 5472 0 -1 6048
box -48 -56 1008 834
use sg13g2_mux2_1  _062_
timestamp 1677247768
transform 1 0 33504 0 1 6048
box -48 -56 1008 834
use sg13g2_mux2_1  _063_
timestamp 1677247768
transform 1 0 21120 0 -1 7560
box -48 -56 1008 834
use sg13g2_mux4_1  _064_
timestamp 1677257233
transform 1 0 15552 0 -1 3024
box -48 -56 2064 834
use sg13g2_mux4_1  _065_
timestamp 1677257233
transform 1 0 9120 0 1 4536
box -48 -56 2064 834
use sg13g2_mux4_1  _066_
timestamp 1677257233
transform 1 0 33216 0 -1 6048
box -48 -56 2064 834
use sg13g2_mux4_1  _067_
timestamp 1677257233
transform 1 0 20736 0 -1 9072
box -48 -56 2064 834
use sg13g2_dlhq_1  _068_
timestamp 1678805552
transform 1 0 16992 0 -1 7560
box -50 -56 1692 834
use sg13g2_dlhq_1  _069_
timestamp 1678805552
transform 1 0 20832 0 -1 4536
box -50 -56 1692 834
use sg13g2_dlhq_1  _070_
timestamp 1678805552
transform 1 0 27552 0 -1 6048
box -50 -56 1692 834
use sg13g2_dlhq_1  _071_
timestamp 1678805552
transform 1 0 30432 0 -1 6048
box -50 -56 1692 834
use sg13g2_dlhq_1  _072_
timestamp 1678805552
transform 1 0 7488 0 1 4536
box -50 -56 1692 834
use sg13g2_dlhq_1  _073_
timestamp 1678805552
transform 1 0 9696 0 -1 3024
box -50 -56 1692 834
use sg13g2_dlhq_1  _074_
timestamp 1678805552
transform 1 0 6816 0 1 1512
box -50 -56 1692 834
use sg13g2_dlhq_1  _075_
timestamp 1678805552
transform -1 0 18528 0 1 1512
box -50 -56 1692 834
use sg13g2_dlhq_1  _076_
timestamp 1678805552
transform 1 0 19968 0 -1 6048
box -50 -56 1692 834
use sg13g2_dlhq_1  _077_
timestamp 1678805552
transform 1 0 30240 0 1 6048
box -50 -56 1692 834
use sg13g2_dlhq_1  _078_
timestamp 1678805552
transform 1 0 3648 0 1 6048
box -50 -56 1692 834
use sg13g2_dlhq_1  _079_
timestamp 1678805552
transform 1 0 12192 0 -1 4536
box -50 -56 1692 834
use sg13g2_dlhq_1  _080_
timestamp 1678805552
transform -1 0 32256 0 -1 9072
box -50 -56 1692 834
use sg13g2_dlhq_1  _081_
timestamp 1678805552
transform 1 0 37248 0 1 4536
box -50 -56 1692 834
use sg13g2_dlhq_1  _082_
timestamp 1678805552
transform -1 0 13920 0 1 4536
box -50 -56 1692 834
use sg13g2_dlhq_1  _083_
timestamp 1678805552
transform 1 0 27552 0 -1 4536
box -50 -56 1692 834
use sg13g2_dlhq_1  _084_
timestamp 1678805552
transform 1 0 16128 0 1 9072
box -50 -56 1692 834
use sg13g2_dlhq_1  _085_
timestamp 1678805552
transform 1 0 34848 0 1 4536
box -50 -56 1692 834
use sg13g2_dlhq_1  _086_
timestamp 1678805552
transform 1 0 6720 0 -1 9072
box -50 -56 1692 834
use sg13g2_dlhq_1  _087_
timestamp 1678805552
transform 1 0 11328 0 -1 3024
box -50 -56 1692 834
use sg13g2_dlhq_1  _088_
timestamp 1678805552
transform 1 0 32640 0 1 9072
box -50 -56 1692 834
use sg13g2_dlhq_1  _089_
timestamp 1678805552
transform 1 0 37152 0 -1 4536
box -50 -56 1692 834
use sg13g2_dlhq_1  _090_
timestamp 1678805552
transform -1 0 17280 0 -1 6048
box -50 -56 1692 834
use sg13g2_dlhq_1  _091_
timestamp 1678805552
transform -1 0 25728 0 -1 4536
box -50 -56 1692 834
use sg13g2_dlhq_1  _092_
timestamp 1678805552
transform -1 0 27264 0 -1 6048
box -50 -56 1692 834
use sg13g2_dlhq_1  _093_
timestamp 1678805552
transform 1 0 31872 0 1 6048
box -50 -56 1692 834
use sg13g2_dlhq_1  _094_
timestamp 1678805552
transform 1 0 3840 0 1 3024
box -50 -56 1692 834
use sg13g2_dlhq_1  _095_
timestamp 1678805552
transform 1 0 9216 0 1 1512
box -50 -56 1692 834
use sg13g2_dlhq_1  _096_
timestamp 1678805552
transform -1 0 37536 0 -1 9072
box -50 -56 1692 834
use sg13g2_dlhq_1  _097_
timestamp 1678805552
transform 1 0 40416 0 -1 6048
box -50 -56 1692 834
use sg13g2_dlhq_1  _098_
timestamp 1678805552
transform -1 0 14016 0 1 9072
box -50 -56 1692 834
use sg13g2_dlhq_1  _099_
timestamp 1678805552
transform 1 0 22848 0 1 4536
box -50 -56 1692 834
use sg13g2_dlhq_1  _100_
timestamp 1678805552
transform 1 0 17280 0 1 7560
box -50 -56 1692 834
use sg13g2_dlhq_1  _101_
timestamp 1678805552
transform 1 0 21024 0 1 4536
box -50 -56 1692 834
use sg13g2_dlhq_1  _102_
timestamp 1678805552
transform -1 0 14880 0 -1 6048
box -50 -56 1692 834
use sg13g2_dlhq_1  _103_
timestamp 1678805552
transform 1 0 16992 0 1 4536
box -50 -56 1692 834
use sg13g2_dlhq_1  _104_
timestamp 1678805552
transform 1 0 22752 0 -1 9072
box -50 -56 1692 834
use sg13g2_dlhq_1  _105_
timestamp 1678805552
transform 1 0 32736 0 1 1512
box -50 -56 1692 834
use sg13g2_dlhq_1  _106_
timestamp 1678805552
transform 1 0 5664 0 -1 3024
box -50 -56 1692 834
use sg13g2_dlhq_1  _107_
timestamp 1678805552
transform 1 0 25920 0 1 1512
box -50 -56 1692 834
use sg13g2_dlhq_1  _108_
timestamp 1678805552
transform 1 0 20640 0 1 6048
box -50 -56 1692 834
use sg13g2_dlhq_1  _109_
timestamp 1678805552
transform 1 0 30624 0 -1 7560
box -50 -56 1692 834
use sg13g2_dlhq_1  _110_
timestamp 1678805552
transform 1 0 3456 0 -1 6048
box -50 -56 1692 834
use sg13g2_dlhq_1  _111_
timestamp 1678805552
transform 1 0 11328 0 1 3024
box -50 -56 1692 834
use sg13g2_dlhq_1  _112_
timestamp 1678805552
transform 1 0 31296 0 1 7560
box -50 -56 1692 834
use sg13g2_dlhq_1  _113_
timestamp 1678805552
transform 1 0 39360 0 -1 7560
box -50 -56 1692 834
use sg13g2_dlhq_1  _114_
timestamp 1678805552
transform -1 0 13920 0 1 7560
box -50 -56 1692 834
use sg13g2_dlhq_1  _115_
timestamp 1678805552
transform -1 0 27360 0 -1 4536
box -50 -56 1692 834
use sg13g2_dlhq_1  _116_
timestamp 1678805552
transform 1 0 16224 0 -1 9072
box -50 -56 1692 834
use sg13g2_dlhq_1  _117_
timestamp 1678805552
transform 1 0 29664 0 -1 4536
box -50 -56 1692 834
use sg13g2_dlhq_1  _118_
timestamp 1678805552
transform 1 0 7488 0 1 7560
box -50 -56 1692 834
use sg13g2_dlhq_1  _119_
timestamp 1678805552
transform 1 0 13920 0 -1 3024
box -50 -56 1692 834
use sg13g2_dlhq_1  _120_
timestamp 1678805552
transform -1 0 30624 0 -1 9072
box -50 -56 1692 834
use sg13g2_dlhq_1  _121_
timestamp 1678805552
transform 1 0 36576 0 -1 3024
box -50 -56 1692 834
use sg13g2_dlhq_1  _122_
timestamp 1678805552
transform -1 0 16608 0 1 4536
box -50 -56 1692 834
use sg13g2_dlhq_1  _123_
timestamp 1678805552
transform 1 0 26016 0 -1 3024
box -50 -56 1692 834
use sg13g2_dlhq_1  _124_
timestamp 1678805552
transform 1 0 26304 0 1 3024
box -50 -56 1692 834
use sg13g2_dlhq_1  _125_
timestamp 1678805552
transform -1 0 32544 0 -1 3024
box -50 -56 1692 834
use sg13g2_dlhq_1  _126_
timestamp 1678805552
transform 1 0 4704 0 -1 4536
box -50 -56 1692 834
use sg13g2_dlhq_1  _127_
timestamp 1678805552
transform 1 0 7488 0 -1 3024
box -50 -56 1692 834
use sg13g2_dlhq_1  _128_
timestamp 1678805552
transform 1 0 36096 0 1 3024
box -50 -56 1692 834
use sg13g2_dlhq_1  _129_
timestamp 1678805552
transform -1 0 41760 0 -1 4536
box -50 -56 1692 834
use sg13g2_dlhq_1  _130_
timestamp 1678805552
transform 1 0 14016 0 -1 9072
box -50 -56 1692 834
use sg13g2_dlhq_1  _131_
timestamp 1678805552
transform 1 0 24384 0 1 7560
box -50 -56 1692 834
use sg13g2_dlhq_1  _132_
timestamp 1678805552
transform 1 0 16800 0 -1 4536
box -50 -56 1692 834
use sg13g2_dlhq_1  _133_
timestamp 1678805552
transform -1 0 22176 0 1 1512
box -50 -56 1692 834
use sg13g2_dlhq_1  _134_
timestamp 1678805552
transform -1 0 14976 0 1 6048
box -50 -56 1692 834
use sg13g2_dlhq_1  _135_
timestamp 1678805552
transform -1 0 17376 0 1 6048
box -50 -56 1692 834
use sg13g2_dlhq_1  _136_
timestamp 1678805552
transform 1 0 30432 0 1 3024
box -50 -56 1692 834
use sg13g2_dlhq_1  _137_
timestamp 1678805552
transform 1 0 32544 0 -1 3024
box -50 -56 1692 834
use sg13g2_dlhq_1  _138_
timestamp 1678805552
transform 1 0 6240 0 1 9072
box -50 -56 1692 834
use sg13g2_dlhq_1  _139_
timestamp 1678805552
transform 1 0 18528 0 1 6048
box -50 -56 1692 834
use sg13g2_dlhq_1  _140_
timestamp 1678805552
transform 1 0 21120 0 -1 3024
box -50 -56 1692 834
use sg13g2_dlhq_1  _141_
timestamp 1678805552
transform -1 0 30048 0 1 6048
box -50 -56 1692 834
use sg13g2_dlhq_1  _142_
timestamp 1678805552
transform 1 0 4320 0 -1 9072
box -50 -56 1692 834
use sg13g2_dlhq_1  _143_
timestamp 1678805552
transform -1 0 12768 0 -1 9072
box -50 -56 1692 834
use sg13g2_dlhq_1  _144_
timestamp 1678805552
transform 1 0 37440 0 1 7560
box -50 -56 1692 834
use sg13g2_dlhq_1  _145_
timestamp 1678805552
transform 1 0 38496 0 -1 6048
box -50 -56 1692 834
use sg13g2_dlhq_1  _146_
timestamp 1678805552
transform 1 0 26208 0 1 7560
box -50 -56 1692 834
use sg13g2_dlhq_1  _147_
timestamp 1678805552
transform 1 0 27840 0 -1 7560
box -50 -56 1692 834
use sg13g2_dlhq_1  _148_
timestamp 1678805552
transform 1 0 14208 0 1 7560
box -50 -56 1692 834
use sg13g2_dlhq_1  _149_
timestamp 1678805552
transform -1 0 20064 0 -1 4536
box -50 -56 1692 834
use sg13g2_dlhq_1  _150_
timestamp 1678805552
transform 1 0 4416 0 1 7560
box -50 -56 1692 834
use sg13g2_dlhq_1  _151_
timestamp 1678805552
transform -1 0 9216 0 1 6048
box -50 -56 1692 834
use sg13g2_dlhq_1  _152_
timestamp 1678805552
transform 1 0 32928 0 1 7560
box -50 -56 1692 834
use sg13g2_dlhq_1  _153_
timestamp 1678805552
transform -1 0 38304 0 1 6048
box -50 -56 1692 834
use sg13g2_dlhq_1  _154_
timestamp 1678805552
transform 1 0 17952 0 -1 6048
box -50 -56 1692 834
use sg13g2_dlhq_1  _155_
timestamp 1678805552
transform -1 0 26592 0 1 6048
box -50 -56 1692 834
use sg13g2_buf_1  _157_
timestamp 1676381911
transform 1 0 25920 0 1 4536
box -48 -56 432 834
use sg13g2_buf_1  _158_
timestamp 1676381911
transform 1 0 31296 0 1 1512
box -48 -56 432 834
use sg13g2_buf_1  _159_
timestamp 1676381911
transform 1 0 4032 0 -1 4536
box -48 -56 432 834
use sg13g2_buf_1  _160_
timestamp 1676381911
transform 1 0 6432 0 1 1512
box -48 -56 432 834
use sg13g2_buf_1  _161_
timestamp 1676381911
transform 1 0 35904 0 -1 4536
box -48 -56 432 834
use sg13g2_buf_1  _162_
timestamp 1676381911
transform 1 0 40224 0 1 4536
box -48 -56 432 834
use sg13g2_buf_1  _163_
timestamp 1676381911
transform 1 0 11136 0 1 7560
box -48 -56 432 834
use sg13g2_buf_1  _164_
timestamp 1676381911
transform 1 0 23904 0 -1 7560
box -48 -56 432 834
use sg13g2_buf_1  _165_
timestamp 1676381911
transform 1 0 16608 0 -1 7560
box -48 -56 432 834
use sg13g2_buf_1  _166_
timestamp 1676381911
transform 1 0 20448 0 -1 4536
box -48 -56 432 834
use sg13g2_buf_1  _167_
timestamp 1676381911
transform 1 0 12960 0 1 6048
box -48 -56 432 834
use sg13g2_buf_1  _168_
timestamp 1676381911
transform 1 0 29760 0 -1 6048
box -48 -56 432 834
use sg13g2_buf_1  _169_
timestamp 1676381911
transform 1 0 30240 0 -1 7560
box -48 -56 432 834
use sg13g2_buf_1  _170_
timestamp 1676381911
transform 1 0 31776 0 1 1512
box -48 -56 432 834
use sg13g2_buf_1  _171_
timestamp 1676381911
transform 1 0 5280 0 -1 3024
box -48 -56 432 834
use sg13g2_buf_1  _172_
timestamp 1676381911
transform 1 0 23712 0 -1 4536
box -48 -56 432 834
use sg13g2_buf_1  _173_
timestamp 1676381911
transform 1 0 20928 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  _174_
timestamp 1676381911
transform 1 0 29472 0 -1 7560
box -48 -56 432 834
use sg13g2_buf_1  _175_
timestamp 1676381911
transform 1 0 3456 0 -1 7560
box -48 -56 432 834
use sg13g2_buf_1  _176_
timestamp 1676381911
transform 1 0 11808 0 1 4536
box -48 -56 432 834
use sg13g2_buf_1  _177_
timestamp 1676381911
transform 1 0 39072 0 -1 9072
box -48 -56 432 834
use sg13g2_buf_1  _178_
timestamp 1676381911
transform 1 0 38880 0 1 4536
box -48 -56 432 834
use sg13g2_buf_1  _179_
timestamp 1676381911
transform 1 0 12768 0 -1 6048
box -48 -56 432 834
use sg13g2_buf_1  _180_
timestamp 1676381911
transform 1 0 27072 0 1 6048
box -48 -56 432 834
use sg13g2_buf_1  _181_
timestamp 1676381911
transform 1 0 14304 0 -1 7560
box -48 -56 432 834
use sg13g2_buf_1  _182_
timestamp 1676381911
transform 1 0 34848 0 -1 4536
box -48 -56 432 834
use sg13g2_buf_1  _183_
timestamp 1676381911
transform 1 0 4032 0 1 7560
box -48 -56 432 834
use sg13g2_buf_1  _184_
timestamp 1676381911
transform 1 0 9312 0 -1 3024
box -48 -56 432 834
use sg13g2_buf_1  _185_
timestamp 1676381911
transform 1 0 33408 0 -1 7560
box -48 -56 432 834
use sg13g2_buf_1  _186_
timestamp 1676381911
transform 1 0 36192 0 -1 3024
box -48 -56 432 834
use sg13g2_buf_1  _187_
timestamp 1676381911
transform 1 0 14880 0 -1 6048
box -48 -56 432 834
use sg13g2_buf_1  _188_
timestamp 1676381911
transform 1 0 25248 0 -1 6048
box -48 -56 432 834
use sg13g2_buf_1  _189_
timestamp 1676381911
transform -1 0 39744 0 1 7560
box -48 -56 432 834
use sg13g2_buf_1  _190_
timestamp 1676381911
transform -1 0 41568 0 1 7560
box -48 -56 432 834
use sg13g2_buf_1  _191_
timestamp 1676381911
transform -1 0 40224 0 -1 9072
box -48 -56 432 834
use sg13g2_buf_1  _192_
timestamp 1676381911
transform -1 0 42048 0 -1 3024
box -48 -56 432 834
use sg13g2_buf_1  _193_
timestamp 1676381911
transform -1 0 42432 0 -1 3024
box -48 -56 432 834
use sg13g2_buf_1  _194_
timestamp 1676381911
transform -1 0 41664 0 -1 3024
box -48 -56 432 834
use sg13g2_buf_1  _195_
timestamp 1676381911
transform -1 0 44448 0 -1 3024
box -48 -56 432 834
use sg13g2_buf_1  _196_
timestamp 1676381911
transform 1 0 34848 0 1 1512
box -48 -56 432 834
use sg13g2_buf_1  _197_
timestamp 1676381911
transform -1 0 42240 0 1 1512
box -48 -56 432 834
use sg13g2_buf_1  _198_
timestamp 1676381911
transform -1 0 40800 0 1 1512
box -48 -56 432 834
use sg13g2_buf_1  _199_
timestamp 1676381911
transform 1 0 36672 0 1 1512
box -48 -56 432 834
use sg13g2_buf_1  _200_
timestamp 1676381911
transform -1 0 44352 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  _201_
timestamp 1676381911
transform -1 0 39360 0 1 1512
box -48 -56 432 834
use sg13g2_buf_1  _202_
timestamp 1676381911
transform -1 0 44448 0 1 4536
box -48 -56 432 834
use sg13g2_buf_1  _203_
timestamp 1676381911
transform -1 0 44736 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  _204_
timestamp 1676381911
transform -1 0 41280 0 -1 9072
box -48 -56 432 834
use sg13g2_buf_1  _205_
timestamp 1676381911
transform -1 0 44352 0 1 6048
box -48 -56 432 834
use sg13g2_buf_1  _206_
timestamp 1676381911
transform -1 0 45216 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  _207_
timestamp 1676381911
transform -1 0 41376 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  _208_
timestamp 1676381911
transform -1 0 44448 0 1 1512
box -48 -56 432 834
use sg13g2_buf_1  _209_
timestamp 1676381911
transform -1 0 23328 0 1 7560
box -48 -56 432 834
use sg13g2_buf_1  _210_
timestamp 1676381911
transform -1 0 36384 0 -1 6048
box -48 -56 432 834
use sg13g2_buf_1  _211_
timestamp 1676381911
transform 1 0 10944 0 -1 4536
box -48 -56 432 834
use sg13g2_buf_1  _212_
timestamp 1676381911
transform -1 0 16896 0 1 1512
box -48 -56 432 834
use sg13g2_buf_1  _213_
timestamp 1676381911
transform -1 0 22464 0 -1 7560
box -48 -56 432 834
use sg13g2_buf_1  _214_
timestamp 1676381911
transform -1 0 34272 0 1 4536
box -48 -56 432 834
use sg13g2_buf_1  _215_
timestamp 1676381911
transform 1 0 6240 0 -1 7560
box -48 -56 432 834
use sg13g2_buf_1  _216_
timestamp 1676381911
transform -1 0 14976 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  _217_
timestamp 1676381911
transform -1 0 27840 0 -1 7560
box -48 -56 432 834
use sg13g2_buf_1  _218_
timestamp 1676381911
transform -1 0 40128 0 -1 4536
box -48 -56 432 834
use sg13g2_buf_1  _219_
timestamp 1676381911
transform 1 0 8928 0 -1 4536
box -48 -56 432 834
use sg13g2_buf_1  _220_
timestamp 1676381911
transform -1 0 30912 0 -1 3024
box -48 -56 432 834
use sg13g2_buf_1  _221_
timestamp 1676381911
transform -1 0 23712 0 1 7560
box -48 -56 432 834
use sg13g2_buf_1  _222_
timestamp 1676381911
transform -1 0 37536 0 -1 6048
box -48 -56 432 834
use sg13g2_buf_1  _223_
timestamp 1676381911
transform 1 0 8064 0 -1 7560
box -48 -56 432 834
use sg13g2_buf_1  _224_
timestamp 1676381911
transform -1 0 14304 0 1 1512
box -48 -56 432 834
use sg13g2_buf_1  _225_
timestamp 1676381911
transform -1 0 39072 0 -1 9072
box -48 -56 432 834
use sg13g2_buf_1  _226_
timestamp 1676381911
transform -1 0 42144 0 -1 4536
box -48 -56 432 834
use sg13g2_buf_1  _227_
timestamp 1676381911
transform 1 0 11520 0 -1 6048
box -48 -56 432 834
use sg13g2_buf_1  _228_
timestamp 1676381911
transform -1 0 25152 0 1 1512
box -48 -56 432 834
use sg13g2_buf_1  _229_
timestamp 1676381911
transform -1 0 24672 0 1 6048
box -48 -56 432 834
use sg13g2_buf_1  _230_
timestamp 1676381911
transform -1 0 35616 0 -1 6048
box -48 -56 432 834
use sg13g2_buf_1  _231_
timestamp 1676381911
transform 1 0 6336 0 -1 4536
box -48 -56 432 834
use sg13g2_buf_1  _232_
timestamp 1676381911
transform -1 0 12960 0 1 1512
box -48 -56 432 834
use sg13g2_buf_1  _233_
timestamp 1676381911
transform -1 0 37440 0 -1 7560
box -48 -56 432 834
use sg13g2_buf_1  _234_
timestamp 1676381911
transform -1 0 43296 0 1 6048
box -48 -56 432 834
use sg13g2_buf_1  _235_
timestamp 1676381911
transform 1 0 10176 0 -1 6048
box -48 -56 432 834
use sg13g2_buf_1  _236_
timestamp 1676381911
transform -1 0 25152 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  _237_
timestamp 1676381911
transform -1 0 20352 0 -1 7560
box -48 -56 432 834
use sg13g2_buf_1  _238_
timestamp 1676381911
transform -1 0 33984 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  _239_
timestamp 1676381911
transform 1 0 11904 0 -1 6048
box -48 -56 432 834
use sg13g2_buf_1  _240_
timestamp 1676381911
transform -1 0 19680 0 1 1512
box -48 -56 432 834
use sg13g2_buf_1  _241_
timestamp 1676381911
transform -1 0 28032 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  _242_
timestamp 1676381911
transform -1 0 36096 0 -1 3024
box -48 -56 432 834
use sg13g2_buf_1  _243_
timestamp 1676381911
transform 1 0 8256 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  _244_
timestamp 1676381911
transform -1 0 30528 0 -1 3024
box -48 -56 432 834
use sg13g2_buf_1  _245_
timestamp 1676381911
transform -1 0 24480 0 -1 6048
box -48 -56 432 834
use sg13g2_buf_1  _246_
timestamp 1676381911
transform -1 0 37824 0 -1 7560
box -48 -56 432 834
use sg13g2_buf_1  _247_
timestamp 1676381911
transform 1 0 6432 0 -1 6048
box -48 -56 432 834
use sg13g2_buf_1  _248_
timestamp 1676381911
transform 1 0 13920 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  _249_
timestamp 1676381911
transform -1 0 37248 0 1 7560
box -48 -56 432 834
use sg13g2_buf_1  _250_
timestamp 1676381911
transform -1 0 42336 0 -1 7560
box -48 -56 432 834
use sg13g2_buf_1  _251_
timestamp 1676381911
transform 1 0 8448 0 -1 9072
box -48 -56 432 834
use sg13g2_buf_1  _252_
timestamp 1676381911
transform -1 0 25536 0 1 1512
box -48 -56 432 834
use sg13g2_buf_1  _253_
timestamp 1676381911
transform -1 0 20736 0 -1 7560
box -48 -56 432 834
use sg13g2_buf_1  _254_
timestamp 1676381911
transform -1 0 34848 0 -1 4536
box -48 -56 432 834
use sg13g2_buf_1  _255_
timestamp 1676381911
transform 1 0 9408 0 1 6048
box -48 -56 432 834
use sg13g2_buf_1  _256_
timestamp 1676381911
transform -1 0 19488 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  _257_
timestamp 1676381911
transform -1 0 30720 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  _258_
timestamp 1676381911
transform -1 0 39552 0 -1 3024
box -48 -56 432 834
use sg13g2_buf_1  _259_
timestamp 1676381911
transform 1 0 10272 0 -1 4536
box -48 -56 432 834
use sg13g2_buf_1  _260_
timestamp 1676381911
transform -1 0 30144 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  _261_
timestamp 1676381911
transform -1 0 42816 0 -1 3024
box -48 -56 432 834
use sg13g2_antennanp  ANTENNA_1
timestamp 1679999689
transform 1 0 43680 0 1 3024
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_2
timestamp 1679999689
transform -1 0 44160 0 -1 7560
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_3
timestamp 1679999689
transform -1 0 43008 0 -1 9072
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_4
timestamp 1679999689
transform 1 0 42240 0 1 9072
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_5
timestamp 1679999689
transform 1 0 43776 0 1 7560
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_6
timestamp 1679999689
transform 1 0 43008 0 1 3024
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_7
timestamp 1679999689
transform -1 0 42528 0 1 1512
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_8
timestamp 1679999689
transform -1 0 43296 0 -1 6048
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_9
timestamp 1679999689
transform -1 0 43872 0 -1 7560
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_10
timestamp 1679999689
transform 1 0 43200 0 1 7560
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_11
timestamp 1679999689
transform 1 0 41952 0 1 9072
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_12
timestamp 1679999689
transform 1 0 43488 0 1 7560
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_13
timestamp 1679999689
transform 1 0 43296 0 1 3024
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_14
timestamp 1679999689
transform 1 0 42720 0 -1 4536
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_15
timestamp 1679999689
transform -1 0 43584 0 -1 6048
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_16
timestamp 1679999689
transform -1 0 43584 0 -1 7560
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_17
timestamp 1679999689
transform 1 0 42912 0 1 7560
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_18
timestamp 1679999689
transform 1 0 41664 0 1 9072
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_19
timestamp 1679999689
transform -1 0 42720 0 -1 9072
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_20
timestamp 1679999689
transform 1 0 42720 0 1 3024
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_21
timestamp 1679999689
transform 1 0 41568 0 1 3024
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_22
timestamp 1679999689
transform 1 0 42912 0 1 4536
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_23
timestamp 1679999689
transform -1 0 43296 0 -1 7560
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_24
timestamp 1679999689
transform 1 0 42624 0 1 7560
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_25
timestamp 1679999689
transform 1 0 41376 0 1 9072
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_26
timestamp 1679999689
transform -1 0 42432 0 -1 9072
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_27
timestamp 1679999689
transform 1 0 42432 0 1 3024
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_28
timestamp 1679999689
transform 1 0 42144 0 -1 4536
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_29
timestamp 1679999689
transform 1 0 43200 0 1 4536
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_30
timestamp 1679999689
transform 1 0 43392 0 1 6048
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_31
timestamp 1679999689
transform 1 0 42336 0 1 7560
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_32
timestamp 1679999689
transform 1 0 41568 0 -1 9072
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_33
timestamp 1679999689
transform -1 0 42144 0 -1 9072
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_34
timestamp 1679999689
transform -1 0 43296 0 -1 4536
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_35
timestamp 1679999689
transform -1 0 41856 0 1 1512
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_36
timestamp 1679999689
transform 1 0 41280 0 1 3024
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_37
timestamp 1679999689
transform -1 0 43968 0 -1 4536
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_38
timestamp 1679999689
transform -1 0 41568 0 -1 9072
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_39
timestamp 1679999689
transform 1 0 40704 0 1 9072
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_40
timestamp 1679999689
transform 1 0 42048 0 1 7560
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_41
timestamp 1679999689
transform 1 0 42144 0 1 3024
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_42
timestamp 1679999689
transform 1 0 42432 0 -1 4536
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_43
timestamp 1679999689
transform 1 0 43392 0 -1 4536
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_44
timestamp 1679999689
transform 1 0 43680 0 1 4536
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_45
timestamp 1679999689
transform 1 0 41760 0 1 7560
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_46
timestamp 1679999689
transform 1 0 40416 0 1 9072
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_47
timestamp 1679999689
transform 1 0 42720 0 -1 7560
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_48
timestamp 1679999689
transform 1 0 41856 0 1 3024
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_49
timestamp 1679999689
transform -1 0 41568 0 1 1512
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_50
timestamp 1679999689
transform -1 0 43008 0 -1 6048
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_51
timestamp 1679999689
transform 1 0 43680 0 -1 6048
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_52
timestamp 1679999689
transform -1 0 40896 0 -1 9072
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_53
timestamp 1679999689
transform 1 0 40128 0 1 9072
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_54
timestamp 1679999689
transform 1 0 42432 0 -1 7560
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_55
timestamp 1679999689
transform 1 0 40992 0 -1 3024
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_56
timestamp 1679999689
transform -1 0 41280 0 1 1512
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_57
timestamp 1679999689
transform 1 0 44160 0 -1 4536
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_58
timestamp 1679999689
transform 1 0 43680 0 1 6048
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_59
timestamp 1679999689
transform 1 0 40896 0 1 7560
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_60
timestamp 1679999689
transform -1 0 41952 0 -1 7560
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_61
timestamp 1679999689
transform -1 0 40608 0 -1 9072
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_62
timestamp 1679999689
transform 1 0 40704 0 -1 3024
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_63
timestamp 1679999689
transform -1 0 40416 0 1 1512
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_64
timestamp 1679999689
transform -1 0 44448 0 -1 6048
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_65
timestamp 1679999689
transform -1 0 44448 0 -1 7560
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_66
timestamp 1679999689
transform -1 0 44832 0 -1 9072
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_67
timestamp 1679999689
transform 1 0 43392 0 1 9072
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_68
timestamp 1679999689
transform -1 0 44064 0 -1 9072
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_69
timestamp 1679999689
transform 1 0 43008 0 -1 3024
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_70
timestamp 1679999689
transform -1 0 44832 0 1 1512
box -48 -56 336 834
use sg13g2_buf_1  fanout44
timestamp 1676381911
transform -1 0 14304 0 -1 4536
box -48 -56 432 834
use sg13g2_buf_1  fanout45
timestamp 1676381911
transform -1 0 29568 0 -1 6048
box -48 -56 432 834
use sg13g2_buf_1  fanout46
timestamp 1676381911
transform 1 0 37920 0 -1 6048
box -48 -56 432 834
use sg13g2_buf_1  fanout47
timestamp 1676381911
transform 1 0 39456 0 -1 9072
box -48 -56 432 834
use sg13g2_buf_1  fanout48
timestamp 1676381911
transform 1 0 29088 0 1 4536
box -48 -56 432 834
use sg13g2_buf_1  fanout49
timestamp 1676381911
transform -1 0 29568 0 -1 4536
box -48 -56 432 834
use sg13g2_buf_1  fanout50
timestamp 1676381911
transform -1 0 14592 0 1 4536
box -48 -56 432 834
use sg13g2_buf_1  fanout51
timestamp 1676381911
transform -1 0 15648 0 -1 6048
box -48 -56 432 834
use sg13g2_buf_1  fanout52
timestamp 1676381911
transform -1 0 22464 0 -1 6048
box -48 -56 432 834
use sg13g2_buf_1  fanout53
timestamp 1676381911
transform -1 0 14976 0 1 4536
box -48 -56 432 834
use sg13g2_buf_1  fanout54
timestamp 1676381911
transform 1 0 19680 0 1 4536
box -48 -56 432 834
use sg13g2_buf_1  fanout55
timestamp 1676381911
transform 1 0 20064 0 -1 4536
box -48 -56 432 834
use sg13g2_buf_1  fanout56
timestamp 1676381911
transform 1 0 25632 0 -1 7560
box -48 -56 432 834
use sg13g2_buf_1  fanout57
timestamp 1676381911
transform 1 0 20160 0 1 6048
box -48 -56 432 834
use sg13g2_buf_1  fanout58
timestamp 1676381911
transform -1 0 20448 0 1 4536
box -48 -56 432 834
use sg13g2_decap_4  FILLER_0_16
timestamp 1679577901
transform 1 0 2688 0 1 1512
box -48 -56 432 834
use sg13g2_fill_1  FILLER_0_20
timestamp 1677579658
transform 1 0 3072 0 1 1512
box -48 -56 144 834
use sg13g2_decap_4  FILLER_0_25
timestamp 1679577901
transform 1 0 3552 0 1 1512
box -48 -56 432 834
use sg13g2_fill_2  FILLER_0_33
timestamp 1677580104
transform 1 0 4320 0 1 1512
box -48 -56 240 834
use sg13g2_fill_2  FILLER_0_105
timestamp 1677580104
transform 1 0 11232 0 1 1512
box -48 -56 240 834
use sg13g2_fill_2  FILLER_0_145
timestamp 1677580104
transform 1 0 15072 0 1 1512
box -48 -56 240 834
use sg13g2_fill_1  FILLER_0_147
timestamp 1677579658
transform 1 0 15264 0 1 1512
box -48 -56 144 834
use sg13g2_fill_1  FILLER_0_193
timestamp 1677579658
transform 1 0 19680 0 1 1512
box -48 -56 144 834
use sg13g2_fill_2  FILLER_0_219
timestamp 1677580104
transform 1 0 22176 0 1 1512
box -48 -56 240 834
use sg13g2_fill_2  FILLER_0_225
timestamp 1677580104
transform 1 0 22752 0 1 1512
box -48 -56 240 834
use sg13g2_fill_1  FILLER_0_227
timestamp 1677579658
transform 1 0 22944 0 1 1512
box -48 -56 144 834
use sg13g2_fill_2  FILLER_0_275
timestamp 1677580104
transform 1 0 27552 0 1 1512
box -48 -56 240 834
use sg13g2_fill_1  FILLER_0_277
timestamp 1677579658
transform 1 0 27744 0 1 1512
box -48 -56 144 834
use sg13g2_decap_8  FILLER_0_302
timestamp 1679581782
transform 1 0 30144 0 1 1512
box -48 -56 720 834
use sg13g2_decap_4  FILLER_0_309
timestamp 1679577901
transform 1 0 30816 0 1 1512
box -48 -56 432 834
use sg13g2_fill_1  FILLER_0_313
timestamp 1677579658
transform 1 0 31200 0 1 1512
box -48 -56 144 834
use sg13g2_fill_1  FILLER_0_318
timestamp 1677579658
transform 1 0 31680 0 1 1512
box -48 -56 144 834
use sg13g2_decap_4  FILLER_0_323
timestamp 1679577901
transform 1 0 32160 0 1 1512
box -48 -56 432 834
use sg13g2_fill_2  FILLER_0_327
timestamp 1677580104
transform 1 0 32544 0 1 1512
box -48 -56 240 834
use sg13g2_decap_4  FILLER_0_346
timestamp 1679577901
transform 1 0 34368 0 1 1512
box -48 -56 432 834
use sg13g2_fill_1  FILLER_0_350
timestamp 1677579658
transform 1 0 34752 0 1 1512
box -48 -56 144 834
use sg13g2_decap_8  FILLER_0_355
timestamp 1679581782
transform 1 0 35232 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_362
timestamp 1679581782
transform 1 0 35904 0 1 1512
box -48 -56 720 834
use sg13g2_fill_1  FILLER_0_369
timestamp 1677579658
transform 1 0 36576 0 1 1512
box -48 -56 144 834
use sg13g2_decap_8  FILLER_0_374
timestamp 1679581782
transform 1 0 37056 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_381
timestamp 1679581782
transform 1 0 37728 0 1 1512
box -48 -56 720 834
use sg13g2_decap_4  FILLER_0_388
timestamp 1679577901
transform 1 0 38400 0 1 1512
box -48 -56 432 834
use sg13g2_fill_2  FILLER_0_392
timestamp 1677580104
transform 1 0 38784 0 1 1512
box -48 -56 240 834
use sg13g2_decap_8  FILLER_0_398
timestamp 1679581782
transform 1 0 39360 0 1 1512
box -48 -56 720 834
use sg13g2_fill_1  FILLER_0_405
timestamp 1677579658
transform 1 0 40032 0 1 1512
box -48 -56 144 834
use sg13g2_fill_2  FILLER_0_413
timestamp 1677580104
transform 1 0 40800 0 1 1512
box -48 -56 240 834
use sg13g2_fill_1  FILLER_0_451
timestamp 1677579658
transform 1 0 44448 0 1 1512
box -48 -56 144 834
use sg13g2_decap_8  FILLER_1_12
timestamp 1679581782
transform 1 0 2304 0 -1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_19
timestamp 1679581782
transform 1 0 2976 0 -1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_26
timestamp 1679581782
transform 1 0 3648 0 -1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_33
timestamp 1679581782
transform 1 0 4320 0 -1 3024
box -48 -56 720 834
use sg13g2_fill_2  FILLER_1_40
timestamp 1677580104
transform 1 0 4992 0 -1 3024
box -48 -56 240 834
use sg13g2_fill_1  FILLER_1_42
timestamp 1677579658
transform 1 0 5184 0 -1 3024
box -48 -56 144 834
use sg13g2_fill_2  FILLER_1_64
timestamp 1677580104
transform 1 0 7296 0 -1 3024
box -48 -56 240 834
use sg13g2_fill_2  FILLER_1_83
timestamp 1677580104
transform 1 0 9120 0 -1 3024
box -48 -56 240 834
use sg13g2_fill_1  FILLER_1_171
timestamp 1677579658
transform 1 0 17568 0 -1 3024
box -48 -56 144 834
use sg13g2_fill_1  FILLER_1_207
timestamp 1677579658
transform 1 0 21024 0 -1 3024
box -48 -56 144 834
use sg13g2_fill_2  FILLER_1_225
timestamp 1677580104
transform 1 0 22752 0 -1 3024
box -48 -56 240 834
use sg13g2_fill_1  FILLER_1_258
timestamp 1677579658
transform 1 0 25920 0 -1 3024
box -48 -56 144 834
use sg13g2_fill_1  FILLER_1_280
timestamp 1677579658
transform 1 0 28032 0 -1 3024
box -48 -56 144 834
use sg13g2_decap_4  FILLER_1_344
timestamp 1679577901
transform 1 0 34176 0 -1 3024
box -48 -56 432 834
use sg13g2_fill_2  FILLER_1_348
timestamp 1677580104
transform 1 0 34560 0 -1 3024
box -48 -56 240 834
use sg13g2_fill_1  FILLER_1_364
timestamp 1677579658
transform 1 0 36096 0 -1 3024
box -48 -56 144 834
use sg13g2_decap_8  FILLER_1_400
timestamp 1679581782
transform 1 0 39552 0 -1 3024
box -48 -56 720 834
use sg13g2_decap_4  FILLER_1_407
timestamp 1679577901
transform 1 0 40224 0 -1 3024
box -48 -56 432 834
use sg13g2_fill_1  FILLER_1_411
timestamp 1677579658
transform 1 0 40608 0 -1 3024
box -48 -56 144 834
use sg13g2_fill_2  FILLER_1_434
timestamp 1677580104
transform 1 0 42816 0 -1 3024
box -48 -56 240 834
use sg13g2_decap_8  FILLER_2_8
timestamp 1679581782
transform 1 0 1920 0 1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_15
timestamp 1679581782
transform 1 0 2592 0 1 3024
box -48 -56 720 834
use sg13g2_decap_4  FILLER_2_22
timestamp 1679577901
transform 1 0 3264 0 1 3024
box -48 -56 432 834
use sg13g2_fill_2  FILLER_2_26
timestamp 1677580104
transform 1 0 3648 0 1 3024
box -48 -56 240 834
use sg13g2_decap_8  FILLER_2_45
timestamp 1679581782
transform 1 0 5472 0 1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_52
timestamp 1679581782
transform 1 0 6144 0 1 3024
box -48 -56 720 834
use sg13g2_decap_4  FILLER_2_59
timestamp 1679577901
transform 1 0 6816 0 1 3024
box -48 -56 432 834
use sg13g2_fill_1  FILLER_2_63
timestamp 1677579658
transform 1 0 7200 0 1 3024
box -48 -56 144 834
use sg13g2_decap_8  FILLER_2_82
timestamp 1679581782
transform 1 0 9024 0 1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_89
timestamp 1679581782
transform 1 0 9696 0 1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_96
timestamp 1679581782
transform 1 0 10368 0 1 3024
box -48 -56 720 834
use sg13g2_fill_2  FILLER_2_103
timestamp 1677580104
transform 1 0 11040 0 1 3024
box -48 -56 240 834
use sg13g2_fill_1  FILLER_2_105
timestamp 1677579658
transform 1 0 11232 0 1 3024
box -48 -56 144 834
use sg13g2_fill_2  FILLER_2_137
timestamp 1677580104
transform 1 0 14304 0 1 3024
box -48 -56 240 834
use sg13g2_fill_1  FILLER_2_139
timestamp 1677579658
transform 1 0 14496 0 1 3024
box -48 -56 144 834
use sg13g2_decap_8  FILLER_2_165
timestamp 1679581782
transform 1 0 16992 0 1 3024
box -48 -56 720 834
use sg13g2_fill_1  FILLER_2_172
timestamp 1677579658
transform 1 0 17664 0 1 3024
box -48 -56 144 834
use sg13g2_decap_8  FILLER_2_191
timestamp 1679581782
transform 1 0 19488 0 1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_198
timestamp 1679581782
transform 1 0 20160 0 1 3024
box -48 -56 720 834
use sg13g2_fill_1  FILLER_2_205
timestamp 1677579658
transform 1 0 20832 0 1 3024
box -48 -56 144 834
use sg13g2_decap_8  FILLER_2_210
timestamp 1679581782
transform 1 0 21312 0 1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_217
timestamp 1679581782
transform 1 0 21984 0 1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_224
timestamp 1679581782
transform 1 0 22656 0 1 3024
box -48 -56 720 834
use sg13g2_decap_4  FILLER_2_231
timestamp 1679577901
transform 1 0 23328 0 1 3024
box -48 -56 432 834
use sg13g2_fill_1  FILLER_2_235
timestamp 1677579658
transform 1 0 23712 0 1 3024
box -48 -56 144 834
use sg13g2_fill_2  FILLER_2_250
timestamp 1677580104
transform 1 0 25152 0 1 3024
box -48 -56 240 834
use sg13g2_fill_1  FILLER_2_252
timestamp 1677579658
transform 1 0 25344 0 1 3024
box -48 -56 144 834
use sg13g2_decap_4  FILLER_2_257
timestamp 1679577901
transform 1 0 25824 0 1 3024
box -48 -56 432 834
use sg13g2_fill_1  FILLER_2_261
timestamp 1677579658
transform 1 0 26208 0 1 3024
box -48 -56 144 834
use sg13g2_decap_8  FILLER_2_279
timestamp 1679581782
transform 1 0 27936 0 1 3024
box -48 -56 720 834
use sg13g2_fill_1  FILLER_2_286
timestamp 1677579658
transform 1 0 28608 0 1 3024
box -48 -56 144 834
use sg13g2_fill_1  FILLER_2_297
timestamp 1677579658
transform 1 0 29664 0 1 3024
box -48 -56 144 834
use sg13g2_fill_2  FILLER_2_302
timestamp 1677580104
transform 1 0 30144 0 1 3024
box -48 -56 240 834
use sg13g2_fill_1  FILLER_2_304
timestamp 1677579658
transform 1 0 30336 0 1 3024
box -48 -56 144 834
use sg13g2_decap_4  FILLER_2_322
timestamp 1679577901
transform 1 0 32064 0 1 3024
box -48 -56 432 834
use sg13g2_fill_2  FILLER_2_326
timestamp 1677580104
transform 1 0 32448 0 1 3024
box -48 -56 240 834
use sg13g2_decap_8  FILLER_2_342
timestamp 1679581782
transform 1 0 33984 0 1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_349
timestamp 1679581782
transform 1 0 34656 0 1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_356
timestamp 1679581782
transform 1 0 35328 0 1 3024
box -48 -56 720 834
use sg13g2_fill_1  FILLER_2_363
timestamp 1677579658
transform 1 0 36000 0 1 3024
box -48 -56 144 834
use sg13g2_fill_2  FILLER_2_381
timestamp 1677580104
transform 1 0 37728 0 1 3024
box -48 -56 240 834
use sg13g2_decap_8  FILLER_2_404
timestamp 1679581782
transform 1 0 39936 0 1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_411
timestamp 1679581782
transform 1 0 40608 0 1 3024
box -48 -56 720 834
use sg13g2_fill_1  FILLER_2_442
timestamp 1677579658
transform 1 0 43584 0 1 3024
box -48 -56 144 834
use sg13g2_fill_1  FILLER_2_454
timestamp 1677579658
transform 1 0 44736 0 1 3024
box -48 -56 144 834
use sg13g2_decap_8  FILLER_3_8
timestamp 1679581782
transform 1 0 1920 0 -1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_15
timestamp 1679581782
transform 1 0 2592 0 -1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_22
timestamp 1679581782
transform 1 0 3264 0 -1 4536
box -48 -56 720 834
use sg13g2_fill_1  FILLER_3_29
timestamp 1677579658
transform 1 0 3936 0 -1 4536
box -48 -56 144 834
use sg13g2_fill_2  FILLER_3_34
timestamp 1677580104
transform 1 0 4416 0 -1 4536
box -48 -56 240 834
use sg13g2_fill_1  FILLER_3_36
timestamp 1677579658
transform 1 0 4608 0 -1 4536
box -48 -56 144 834
use sg13g2_fill_2  FILLER_3_58
timestamp 1677580104
transform 1 0 6720 0 -1 4536
box -48 -56 240 834
use sg13g2_fill_2  FILLER_3_99
timestamp 1677580104
transform 1 0 10656 0 -1 4536
box -48 -56 240 834
use sg13g2_fill_1  FILLER_3_101
timestamp 1677579658
transform 1 0 10848 0 -1 4536
box -48 -56 144 834
use sg13g2_decap_8  FILLER_3_106
timestamp 1679581782
transform 1 0 11328 0 -1 4536
box -48 -56 720 834
use sg13g2_fill_2  FILLER_3_113
timestamp 1677580104
transform 1 0 12000 0 -1 4536
box -48 -56 240 834
use sg13g2_fill_1  FILLER_3_132
timestamp 1677579658
transform 1 0 13824 0 -1 4536
box -48 -56 144 834
use sg13g2_decap_4  FILLER_3_137
timestamp 1679577901
transform 1 0 14304 0 -1 4536
box -48 -56 432 834
use sg13g2_fill_2  FILLER_3_141
timestamp 1677580104
transform 1 0 14688 0 -1 4536
box -48 -56 240 834
use sg13g2_decap_8  FILLER_3_153
timestamp 1679581782
transform 1 0 15840 0 -1 4536
box -48 -56 720 834
use sg13g2_fill_2  FILLER_3_160
timestamp 1677580104
transform 1 0 16512 0 -1 4536
box -48 -56 240 834
use sg13g2_fill_1  FILLER_3_162
timestamp 1677579658
transform 1 0 16704 0 -1 4536
box -48 -56 144 834
use sg13g2_decap_8  FILLER_3_222
timestamp 1679581782
transform 1 0 22464 0 -1 4536
box -48 -56 720 834
use sg13g2_decap_4  FILLER_3_229
timestamp 1679577901
transform 1 0 23136 0 -1 4536
box -48 -56 432 834
use sg13g2_fill_2  FILLER_3_233
timestamp 1677580104
transform 1 0 23520 0 -1 4536
box -48 -56 240 834
use sg13g2_fill_2  FILLER_3_273
timestamp 1677580104
transform 1 0 27360 0 -1 4536
box -48 -56 240 834
use sg13g2_fill_1  FILLER_3_296
timestamp 1677579658
transform 1 0 29568 0 -1 4536
box -48 -56 144 834
use sg13g2_decap_8  FILLER_3_314
timestamp 1679581782
transform 1 0 31296 0 -1 4536
box -48 -56 720 834
use sg13g2_decap_4  FILLER_3_321
timestamp 1679577901
transform 1 0 31968 0 -1 4536
box -48 -56 432 834
use sg13g2_fill_1  FILLER_3_325
timestamp 1677579658
transform 1 0 32352 0 -1 4536
box -48 -56 144 834
use sg13g2_decap_8  FILLER_3_355
timestamp 1679581782
transform 1 0 35232 0 -1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_366
timestamp 1679581782
transform 1 0 36288 0 -1 4536
box -48 -56 720 834
use sg13g2_fill_2  FILLER_3_373
timestamp 1677580104
transform 1 0 36960 0 -1 4536
box -48 -56 240 834
use sg13g2_fill_1  FILLER_3_439
timestamp 1677579658
transform 1 0 43296 0 -1 4536
box -48 -56 144 834
use sg13g2_fill_2  FILLER_3_446
timestamp 1677580104
transform 1 0 43968 0 -1 4536
box -48 -56 240 834
use sg13g2_decap_8  FILLER_4_8
timestamp 1679581782
transform 1 0 1920 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_15
timestamp 1679581782
transform 1 0 2592 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_22
timestamp 1679581782
transform 1 0 3264 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_29
timestamp 1679581782
transform 1 0 3936 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_36
timestamp 1679581782
transform 1 0 4608 0 1 4536
box -48 -56 720 834
use sg13g2_fill_2  FILLER_4_63
timestamp 1677580104
transform 1 0 7200 0 1 4536
box -48 -56 240 834
use sg13g2_fill_1  FILLER_4_65
timestamp 1677579658
transform 1 0 7392 0 1 4536
box -48 -56 144 834
use sg13g2_fill_2  FILLER_4_104
timestamp 1677580104
transform 1 0 11136 0 1 4536
box -48 -56 240 834
use sg13g2_fill_1  FILLER_4_106
timestamp 1677579658
transform 1 0 11328 0 1 4536
box -48 -56 144 834
use sg13g2_fill_1  FILLER_4_115
timestamp 1677579658
transform 1 0 12192 0 1 4536
box -48 -56 144 834
use sg13g2_fill_2  FILLER_4_133
timestamp 1677580104
transform 1 0 13920 0 1 4536
box -48 -56 240 834
use sg13g2_fill_1  FILLER_4_135
timestamp 1677579658
transform 1 0 14112 0 1 4536
box -48 -56 144 834
use sg13g2_decap_4  FILLER_4_161
timestamp 1679577901
transform 1 0 16608 0 1 4536
box -48 -56 432 834
use sg13g2_decap_8  FILLER_4_182
timestamp 1679581782
transform 1 0 18624 0 1 4536
box -48 -56 720 834
use sg13g2_decap_4  FILLER_4_189
timestamp 1679577901
transform 1 0 19296 0 1 4536
box -48 -56 432 834
use sg13g2_decap_4  FILLER_4_201
timestamp 1679577901
transform 1 0 20448 0 1 4536
box -48 -56 432 834
use sg13g2_fill_2  FILLER_4_205
timestamp 1677580104
transform 1 0 20832 0 1 4536
box -48 -56 240 834
use sg13g2_fill_2  FILLER_4_224
timestamp 1677580104
transform 1 0 22656 0 1 4536
box -48 -56 240 834
use sg13g2_decap_8  FILLER_4_243
timestamp 1679581782
transform 1 0 24480 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_250
timestamp 1679581782
transform 1 0 25152 0 1 4536
box -48 -56 720 834
use sg13g2_fill_1  FILLER_4_257
timestamp 1677579658
transform 1 0 25824 0 1 4536
box -48 -56 144 834
use sg13g2_decap_8  FILLER_4_262
timestamp 1679581782
transform 1 0 26304 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_269
timestamp 1679581782
transform 1 0 26976 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_276
timestamp 1679581782
transform 1 0 27648 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_283
timestamp 1679581782
transform 1 0 28320 0 1 4536
box -48 -56 720 834
use sg13g2_fill_1  FILLER_4_290
timestamp 1677579658
transform 1 0 28992 0 1 4536
box -48 -56 144 834
use sg13g2_decap_8  FILLER_4_295
timestamp 1679581782
transform 1 0 29472 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_302
timestamp 1679581782
transform 1 0 30144 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_309
timestamp 1679581782
transform 1 0 30816 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_316
timestamp 1679581782
transform 1 0 31488 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_323
timestamp 1679581782
transform 1 0 32160 0 1 4536
box -48 -56 720 834
use sg13g2_fill_1  FILLER_4_330
timestamp 1677579658
transform 1 0 32832 0 1 4536
box -48 -56 144 834
use sg13g2_decap_4  FILLER_4_345
timestamp 1679577901
transform 1 0 34272 0 1 4536
box -48 -56 432 834
use sg13g2_fill_2  FILLER_4_349
timestamp 1677580104
transform 1 0 34656 0 1 4536
box -48 -56 240 834
use sg13g2_decap_8  FILLER_4_368
timestamp 1679581782
transform 1 0 36480 0 1 4536
box -48 -56 720 834
use sg13g2_fill_1  FILLER_4_375
timestamp 1677579658
transform 1 0 37152 0 1 4536
box -48 -56 144 834
use sg13g2_decap_8  FILLER_4_397
timestamp 1679581782
transform 1 0 39264 0 1 4536
box -48 -56 720 834
use sg13g2_fill_2  FILLER_4_404
timestamp 1677580104
transform 1 0 39936 0 1 4536
box -48 -56 240 834
use sg13g2_fill_1  FILLER_4_406
timestamp 1677579658
transform 1 0 40128 0 1 4536
box -48 -56 144 834
use sg13g2_decap_8  FILLER_4_421
timestamp 1679581782
transform 1 0 41568 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_428
timestamp 1679581782
transform 1 0 42240 0 1 4536
box -48 -56 720 834
use sg13g2_fill_2  FILLER_4_441
timestamp 1677580104
transform 1 0 43488 0 1 4536
box -48 -56 240 834
use sg13g2_fill_1  FILLER_4_446
timestamp 1677579658
transform 1 0 43968 0 1 4536
box -48 -56 144 834
use sg13g2_decap_8  FILLER_5_12
timestamp 1679581782
transform 1 0 2304 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_4  FILLER_5_19
timestamp 1679577901
transform 1 0 2976 0 -1 6048
box -48 -56 432 834
use sg13g2_fill_1  FILLER_5_23
timestamp 1677579658
transform 1 0 3360 0 -1 6048
box -48 -56 144 834
use sg13g2_decap_4  FILLER_5_41
timestamp 1679577901
transform 1 0 5088 0 -1 6048
box -48 -56 432 834
use sg13g2_decap_8  FILLER_5_59
timestamp 1679581782
transform 1 0 6816 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_66
timestamp 1679581782
transform 1 0 7488 0 -1 6048
box -48 -56 720 834
use sg13g2_fill_2  FILLER_5_73
timestamp 1677580104
transform 1 0 8160 0 -1 6048
box -48 -56 240 834
use sg13g2_fill_1  FILLER_5_75
timestamp 1677579658
transform 1 0 8352 0 -1 6048
box -48 -56 144 834
use sg13g2_decap_8  FILLER_5_86
timestamp 1679581782
transform 1 0 9408 0 -1 6048
box -48 -56 720 834
use sg13g2_fill_1  FILLER_5_93
timestamp 1677579658
transform 1 0 10080 0 -1 6048
box -48 -56 144 834
use sg13g2_fill_1  FILLER_5_116
timestamp 1677579658
transform 1 0 12288 0 -1 6048
box -48 -56 144 834
use sg13g2_fill_1  FILLER_5_125
timestamp 1677579658
transform 1 0 13152 0 -1 6048
box -48 -56 144 834
use sg13g2_decap_8  FILLER_5_168
timestamp 1679581782
transform 1 0 17280 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_4  FILLER_5_192
timestamp 1679577901
transform 1 0 19584 0 -1 6048
box -48 -56 432 834
use sg13g2_decap_4  FILLER_5_213
timestamp 1679577901
transform 1 0 21600 0 -1 6048
box -48 -56 432 834
use sg13g2_fill_1  FILLER_5_217
timestamp 1677579658
transform 1 0 21984 0 -1 6048
box -48 -56 144 834
use sg13g2_decap_8  FILLER_5_222
timestamp 1679581782
transform 1 0 22464 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_243
timestamp 1679581782
transform 1 0 24480 0 -1 6048
box -48 -56 720 834
use sg13g2_fill_1  FILLER_5_250
timestamp 1677579658
transform 1 0 25152 0 -1 6048
box -48 -56 144 834
use sg13g2_fill_2  FILLER_5_272
timestamp 1677580104
transform 1 0 27264 0 -1 6048
box -48 -56 240 834
use sg13g2_fill_1  FILLER_5_274
timestamp 1677579658
transform 1 0 27456 0 -1 6048
box -48 -56 144 834
use sg13g2_fill_2  FILLER_5_296
timestamp 1677580104
transform 1 0 29568 0 -1 6048
box -48 -56 240 834
use sg13g2_fill_2  FILLER_5_302
timestamp 1677580104
transform 1 0 30144 0 -1 6048
box -48 -56 240 834
use sg13g2_fill_1  FILLER_5_304
timestamp 1677579658
transform 1 0 30336 0 -1 6048
box -48 -56 144 834
use sg13g2_decap_8  FILLER_5_367
timestamp 1679581782
transform 1 0 36384 0 -1 6048
box -48 -56 720 834
use sg13g2_fill_1  FILLER_5_374
timestamp 1677579658
transform 1 0 37056 0 -1 6048
box -48 -56 144 834
use sg13g2_decap_4  FILLER_5_379
timestamp 1679577901
transform 1 0 37536 0 -1 6048
box -48 -56 432 834
use sg13g2_fill_2  FILLER_5_387
timestamp 1677580104
transform 1 0 38304 0 -1 6048
box -48 -56 240 834
use sg13g2_fill_2  FILLER_5_406
timestamp 1677580104
transform 1 0 40128 0 -1 6048
box -48 -56 240 834
use sg13g2_fill_1  FILLER_5_408
timestamp 1677579658
transform 1 0 40320 0 -1 6048
box -48 -56 144 834
use sg13g2_decap_8  FILLER_5_426
timestamp 1679581782
transform 1 0 42048 0 -1 6048
box -48 -56 720 834
use sg13g2_fill_1  FILLER_5_442
timestamp 1677579658
transform 1 0 43584 0 -1 6048
box -48 -56 144 834
use sg13g2_fill_2  FILLER_5_446
timestamp 1677580104
transform 1 0 43968 0 -1 6048
box -48 -56 240 834
use sg13g2_decap_8  FILLER_6_8
timestamp 1679581782
transform 1 0 1920 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_15
timestamp 1679581782
transform 1 0 2592 0 1 6048
box -48 -56 720 834
use sg13g2_decap_4  FILLER_6_22
timestamp 1679577901
transform 1 0 3264 0 1 6048
box -48 -56 432 834
use sg13g2_fill_2  FILLER_6_43
timestamp 1677580104
transform 1 0 5280 0 1 6048
box -48 -56 240 834
use sg13g2_fill_1  FILLER_6_45
timestamp 1677579658
transform 1 0 5472 0 1 6048
box -48 -56 144 834
use sg13g2_fill_2  FILLER_6_84
timestamp 1677580104
transform 1 0 9216 0 1 6048
box -48 -56 240 834
use sg13g2_fill_2  FILLER_6_144
timestamp 1677580104
transform 1 0 14976 0 1 6048
box -48 -56 240 834
use sg13g2_fill_1  FILLER_6_146
timestamp 1677579658
transform 1 0 15168 0 1 6048
box -48 -56 144 834
use sg13g2_fill_1  FILLER_6_151
timestamp 1677579658
transform 1 0 15648 0 1 6048
box -48 -56 144 834
use sg13g2_fill_1  FILLER_6_202
timestamp 1677579658
transform 1 0 20544 0 1 6048
box -48 -56 144 834
use sg13g2_fill_2  FILLER_6_245
timestamp 1677580104
transform 1 0 24672 0 1 6048
box -48 -56 240 834
use sg13g2_fill_1  FILLER_6_247
timestamp 1677579658
transform 1 0 24864 0 1 6048
box -48 -56 144 834
use sg13g2_decap_4  FILLER_6_265
timestamp 1679577901
transform 1 0 26592 0 1 6048
box -48 -56 432 834
use sg13g2_fill_1  FILLER_6_269
timestamp 1677579658
transform 1 0 26976 0 1 6048
box -48 -56 144 834
use sg13g2_decap_4  FILLER_6_274
timestamp 1679577901
transform 1 0 27456 0 1 6048
box -48 -56 432 834
use sg13g2_fill_1  FILLER_6_278
timestamp 1677579658
transform 1 0 27840 0 1 6048
box -48 -56 144 834
use sg13g2_fill_1  FILLER_6_283
timestamp 1677579658
transform 1 0 28320 0 1 6048
box -48 -56 144 834
use sg13g2_fill_2  FILLER_6_301
timestamp 1677580104
transform 1 0 30048 0 1 6048
box -48 -56 240 834
use sg13g2_fill_2  FILLER_6_357
timestamp 1677580104
transform 1 0 35424 0 1 6048
box -48 -56 240 834
use sg13g2_fill_1  FILLER_6_359
timestamp 1677579658
transform 1 0 35616 0 1 6048
box -48 -56 144 834
use sg13g2_decap_4  FILLER_6_387
timestamp 1679577901
transform 1 0 38304 0 1 6048
box -48 -56 432 834
use sg13g2_fill_2  FILLER_6_391
timestamp 1677580104
transform 1 0 38688 0 1 6048
box -48 -56 240 834
use sg13g2_fill_1  FILLER_6_414
timestamp 1677579658
transform 1 0 40896 0 1 6048
box -48 -56 144 834
use sg13g2_fill_1  FILLER_6_439
timestamp 1677579658
transform 1 0 43296 0 1 6048
box -48 -56 144 834
use sg13g2_fill_1  FILLER_6_450
timestamp 1677579658
transform 1 0 44352 0 1 6048
box -48 -56 144 834
use sg13g2_decap_8  FILLER_7_8
timestamp 1679581782
transform 1 0 1920 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_15
timestamp 1679581782
transform 1 0 2592 0 -1 7560
box -48 -56 720 834
use sg13g2_fill_2  FILLER_7_22
timestamp 1677580104
transform 1 0 3264 0 -1 7560
box -48 -56 240 834
use sg13g2_decap_8  FILLER_7_28
timestamp 1679581782
transform 1 0 3840 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_35
timestamp 1679581782
transform 1 0 4512 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_42
timestamp 1679581782
transform 1 0 5184 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_4  FILLER_7_49
timestamp 1679577901
transform 1 0 5856 0 -1 7560
box -48 -56 432 834
use sg13g2_decap_8  FILLER_7_57
timestamp 1679581782
transform 1 0 6624 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_64
timestamp 1679581782
transform 1 0 7296 0 -1 7560
box -48 -56 720 834
use sg13g2_fill_1  FILLER_7_71
timestamp 1677579658
transform 1 0 7968 0 -1 7560
box -48 -56 144 834
use sg13g2_fill_2  FILLER_7_94
timestamp 1677580104
transform 1 0 10176 0 -1 7560
box -48 -56 240 834
use sg13g2_fill_1  FILLER_7_96
timestamp 1677579658
transform 1 0 10368 0 -1 7560
box -48 -56 144 834
use sg13g2_fill_2  FILLER_7_107
timestamp 1677580104
transform 1 0 11424 0 -1 7560
box -48 -56 240 834
use sg13g2_fill_2  FILLER_7_182
timestamp 1677580104
transform 1 0 18624 0 -1 7560
box -48 -56 240 834
use sg13g2_fill_1  FILLER_7_236
timestamp 1677579658
transform 1 0 23808 0 -1 7560
box -48 -56 144 834
use sg13g2_decap_8  FILLER_7_241
timestamp 1679581782
transform 1 0 24288 0 -1 7560
box -48 -56 720 834
use sg13g2_fill_1  FILLER_7_248
timestamp 1677579658
transform 1 0 24960 0 -1 7560
box -48 -56 144 834
use sg13g2_fill_2  FILLER_7_253
timestamp 1677580104
transform 1 0 25440 0 -1 7560
box -48 -56 240 834
use sg13g2_decap_4  FILLER_7_263
timestamp 1679577901
transform 1 0 26400 0 -1 7560
box -48 -56 432 834
use sg13g2_fill_2  FILLER_7_267
timestamp 1677580104
transform 1 0 26784 0 -1 7560
box -48 -56 240 834
use sg13g2_fill_1  FILLER_7_273
timestamp 1677579658
transform 1 0 27360 0 -1 7560
box -48 -56 144 834
use sg13g2_fill_1  FILLER_7_344
timestamp 1677579658
transform 1 0 34176 0 -1 7560
box -48 -56 144 834
use sg13g2_decap_8  FILLER_7_382
timestamp 1679581782
transform 1 0 37824 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_389
timestamp 1679581782
transform 1 0 38496 0 -1 7560
box -48 -56 720 834
use sg13g2_fill_2  FILLER_7_396
timestamp 1677580104
transform 1 0 39168 0 -1 7560
box -48 -56 240 834
use sg13g2_decap_8  FILLER_7_415
timestamp 1679581782
transform 1 0 40992 0 -1 7560
box -48 -56 720 834
use sg13g2_fill_1  FILLER_7_429
timestamp 1677579658
transform 1 0 42336 0 -1 7560
box -48 -56 144 834
use sg13g2_decap_8  FILLER_8_8
timestamp 1679581782
transform 1 0 1920 0 1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_15
timestamp 1679581782
transform 1 0 2592 0 1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_22
timestamp 1679581782
transform 1 0 3264 0 1 7560
box -48 -56 720 834
use sg13g2_fill_1  FILLER_8_29
timestamp 1677579658
transform 1 0 3936 0 1 7560
box -48 -56 144 834
use sg13g2_decap_8  FILLER_8_51
timestamp 1679581782
transform 1 0 6048 0 1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_58
timestamp 1679581782
transform 1 0 6720 0 1 7560
box -48 -56 720 834
use sg13g2_fill_1  FILLER_8_65
timestamp 1677579658
transform 1 0 7392 0 1 7560
box -48 -56 144 834
use sg13g2_fill_2  FILLER_8_83
timestamp 1677580104
transform 1 0 9120 0 1 7560
box -48 -56 240 834
use sg13g2_fill_1  FILLER_8_85
timestamp 1677579658
transform 1 0 9312 0 1 7560
box -48 -56 144 834
use sg13g2_fill_2  FILLER_8_133
timestamp 1677580104
transform 1 0 13920 0 1 7560
box -48 -56 240 834
use sg13g2_fill_1  FILLER_8_135
timestamp 1677579658
transform 1 0 14112 0 1 7560
box -48 -56 144 834
use sg13g2_fill_2  FILLER_8_153
timestamp 1677580104
transform 1 0 15840 0 1 7560
box -48 -56 240 834
use sg13g2_fill_1  FILLER_8_155
timestamp 1677579658
transform 1 0 16032 0 1 7560
box -48 -56 144 834
use sg13g2_fill_2  FILLER_8_185
timestamp 1677580104
transform 1 0 18912 0 1 7560
box -48 -56 240 834
use sg13g2_fill_1  FILLER_8_187
timestamp 1677579658
transform 1 0 19104 0 1 7560
box -48 -56 144 834
use sg13g2_fill_2  FILLER_8_198
timestamp 1677580104
transform 1 0 20160 0 1 7560
box -48 -56 240 834
use sg13g2_fill_1  FILLER_8_200
timestamp 1677579658
transform 1 0 20352 0 1 7560
box -48 -56 144 834
use sg13g2_decap_8  FILLER_8_235
timestamp 1679581782
transform 1 0 23712 0 1 7560
box -48 -56 720 834
use sg13g2_fill_2  FILLER_8_259
timestamp 1677580104
transform 1 0 26016 0 1 7560
box -48 -56 240 834
use sg13g2_fill_2  FILLER_8_311
timestamp 1677580104
transform 1 0 31008 0 1 7560
box -48 -56 240 834
use sg13g2_fill_1  FILLER_8_313
timestamp 1677579658
transform 1 0 31200 0 1 7560
box -48 -56 144 834
use sg13g2_fill_2  FILLER_8_352
timestamp 1677580104
transform 1 0 34944 0 1 7560
box -48 -56 240 834
use sg13g2_fill_2  FILLER_8_376
timestamp 1677580104
transform 1 0 37248 0 1 7560
box -48 -56 240 834
use sg13g2_fill_2  FILLER_8_395
timestamp 1677580104
transform 1 0 39072 0 1 7560
box -48 -56 240 834
use sg13g2_fill_1  FILLER_8_397
timestamp 1677579658
transform 1 0 39264 0 1 7560
box -48 -56 144 834
use sg13g2_decap_8  FILLER_8_402
timestamp 1679581782
transform 1 0 39744 0 1 7560
box -48 -56 720 834
use sg13g2_decap_4  FILLER_8_409
timestamp 1679577901
transform 1 0 40416 0 1 7560
box -48 -56 432 834
use sg13g2_fill_1  FILLER_8_413
timestamp 1677579658
transform 1 0 40800 0 1 7560
box -48 -56 144 834
use sg13g2_fill_2  FILLER_8_421
timestamp 1677580104
transform 1 0 41568 0 1 7560
box -48 -56 240 834
use sg13g2_decap_8  FILLER_9_16
timestamp 1679581782
transform 1 0 2688 0 -1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_23
timestamp 1679581782
transform 1 0 3360 0 -1 9072
box -48 -56 720 834
use sg13g2_fill_2  FILLER_9_30
timestamp 1677580104
transform 1 0 4032 0 -1 9072
box -48 -56 240 834
use sg13g2_fill_1  FILLER_9_32
timestamp 1677579658
transform 1 0 4224 0 -1 9072
box -48 -56 144 834
use sg13g2_decap_8  FILLER_9_50
timestamp 1679581782
transform 1 0 5952 0 -1 9072
box -48 -56 720 834
use sg13g2_fill_1  FILLER_9_57
timestamp 1677579658
transform 1 0 6624 0 -1 9072
box -48 -56 144 834
use sg13g2_fill_1  FILLER_9_75
timestamp 1677579658
transform 1 0 8352 0 -1 9072
box -48 -56 144 834
use sg13g2_fill_2  FILLER_9_101
timestamp 1677580104
transform 1 0 10848 0 -1 9072
box -48 -56 240 834
use sg13g2_fill_1  FILLER_9_103
timestamp 1677579658
transform 1 0 11040 0 -1 9072
box -48 -56 144 834
use sg13g2_fill_1  FILLER_9_121
timestamp 1677579658
transform 1 0 12768 0 -1 9072
box -48 -56 144 834
use sg13g2_fill_2  FILLER_9_151
timestamp 1677580104
transform 1 0 15648 0 -1 9072
box -48 -56 240 834
use sg13g2_fill_1  FILLER_9_174
timestamp 1677579658
transform 1 0 17856 0 -1 9072
box -48 -56 144 834
use sg13g2_fill_2  FILLER_9_263
timestamp 1677580104
transform 1 0 26400 0 -1 9072
box -48 -56 240 834
use sg13g2_fill_1  FILLER_9_265
timestamp 1677579658
transform 1 0 26592 0 -1 9072
box -48 -56 144 834
use sg13g2_fill_2  FILLER_9_288
timestamp 1677580104
transform 1 0 28800 0 -1 9072
box -48 -56 240 834
use sg13g2_fill_1  FILLER_9_332
timestamp 1677579658
transform 1 0 33024 0 -1 9072
box -48 -56 144 834
use sg13g2_fill_2  FILLER_9_343
timestamp 1677580104
transform 1 0 34080 0 -1 9072
box -48 -56 240 834
use sg13g2_fill_2  FILLER_9_359
timestamp 1677580104
transform 1 0 35616 0 -1 9072
box -48 -56 240 834
use sg13g2_fill_1  FILLER_9_361
timestamp 1677579658
transform 1 0 35808 0 -1 9072
box -48 -56 144 834
use sg13g2_fill_1  FILLER_9_407
timestamp 1677579658
transform 1 0 40224 0 -1 9072
box -48 -56 144 834
use sg13g2_fill_1  FILLER_9_451
timestamp 1677579658
transform 1 0 44448 0 -1 9072
box -48 -56 144 834
use sg13g2_decap_8  FILLER_10_24
timestamp 1679581782
transform 1 0 3456 0 1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_31
timestamp 1679581782
transform 1 0 4128 0 1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_38
timestamp 1679581782
transform 1 0 4800 0 1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_45
timestamp 1679581782
transform 1 0 5472 0 1 9072
box -48 -56 720 834
use sg13g2_fill_1  FILLER_10_52
timestamp 1677579658
transform 1 0 6144 0 1 9072
box -48 -56 144 834
use sg13g2_fill_2  FILLER_10_102
timestamp 1677580104
transform 1 0 10944 0 1 9072
box -48 -56 240 834
use sg13g2_fill_1  FILLER_10_104
timestamp 1677579658
transform 1 0 11136 0 1 9072
box -48 -56 144 834
use sg13g2_fill_2  FILLER_10_134
timestamp 1677580104
transform 1 0 14016 0 1 9072
box -48 -56 240 834
use sg13g2_fill_2  FILLER_10_199
timestamp 1677580104
transform 1 0 20256 0 1 9072
box -48 -56 240 834
use sg13g2_fill_1  FILLER_10_201
timestamp 1677579658
transform 1 0 20448 0 1 9072
box -48 -56 144 834
use sg13g2_fill_2  FILLER_10_264
timestamp 1677580104
transform 1 0 26496 0 1 9072
box -48 -56 240 834
use sg13g2_fill_1  FILLER_10_349
timestamp 1677579658
transform 1 0 34656 0 1 9072
box -48 -56 144 834
use sg13g2_fill_2  FILLER_10_404
timestamp 1677580104
transform 1 0 39936 0 1 9072
box -48 -56 240 834
use sg13g2_fill_1  FILLER_10_439
timestamp 1677579658
transform 1 0 43296 0 1 9072
box -48 -56 144 834
use sg13g2_buf_1  input1
timestamp 1676381911
transform 1 0 1536 0 1 1512
box -48 -56 432 834
use sg13g2_buf_1  input2
timestamp 1676381911
transform 1 0 1152 0 -1 4536
box -48 -56 432 834
use sg13g2_buf_1  input3
timestamp 1676381911
transform 1 0 1536 0 1 4536
box -48 -56 432 834
use sg13g2_buf_1  input4
timestamp 1676381911
transform 1 0 1152 0 1 4536
box -48 -56 432 834
use sg13g2_buf_1  input5
timestamp 1676381911
transform 1 0 1920 0 -1 6048
box -48 -56 432 834
use sg13g2_buf_1  input6
timestamp 1676381911
transform 1 0 1536 0 -1 6048
box -48 -56 432 834
use sg13g2_buf_1  input7
timestamp 1676381911
transform 1 0 1152 0 -1 6048
box -48 -56 432 834
use sg13g2_buf_1  input8
timestamp 1676381911
transform 1 0 1536 0 1 6048
box -48 -56 432 834
use sg13g2_buf_1  input9
timestamp 1676381911
transform 1 0 1152 0 1 6048
box -48 -56 432 834
use sg13g2_buf_1  input10
timestamp 1676381911
transform 1 0 1536 0 -1 7560
box -48 -56 432 834
use sg13g2_buf_1  input11
timestamp 1676381911
transform 1 0 1152 0 -1 7560
box -48 -56 432 834
use sg13g2_buf_1  input12
timestamp 1676381911
transform 1 0 1920 0 1 1512
box -48 -56 432 834
use sg13g2_buf_1  input13
timestamp 1676381911
transform 1 0 1152 0 1 7560
box -48 -56 432 834
use sg13g2_buf_1  input14
timestamp 1676381911
transform 1 0 1536 0 1 7560
box -48 -56 432 834
use sg13g2_buf_1  input15
timestamp 1676381911
transform 1 0 1152 0 -1 9072
box -48 -56 432 834
use sg13g2_buf_1  input16
timestamp 1676381911
transform 1 0 1536 0 -1 9072
box -48 -56 432 834
use sg13g2_buf_1  input17
timestamp 1676381911
transform 1 0 1920 0 -1 9072
box -48 -56 432 834
use sg13g2_buf_1  input18
timestamp 1676381911
transform 1 0 1152 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  input19
timestamp 1676381911
transform 1 0 1536 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  input20
timestamp 1676381911
transform 1 0 1920 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  input21
timestamp 1676381911
transform 1 0 2304 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  input22
timestamp 1676381911
transform 1 0 2688 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  input23
timestamp 1676381911
transform 1 0 2304 0 1 1512
box -48 -56 432 834
use sg13g2_buf_1  input24
timestamp 1676381911
transform 1 0 2304 0 -1 9072
box -48 -56 432 834
use sg13g2_buf_1  input25
timestamp 1676381911
transform 1 0 3072 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  input26
timestamp 1676381911
transform 1 0 1152 0 1 1512
box -48 -56 432 834
use sg13g2_buf_1  input27
timestamp 1676381911
transform 1 0 1920 0 -1 3024
box -48 -56 432 834
use sg13g2_buf_1  input28
timestamp 1676381911
transform 1 0 1536 0 -1 3024
box -48 -56 432 834
use sg13g2_buf_1  input29
timestamp 1676381911
transform 1 0 1152 0 -1 3024
box -48 -56 432 834
use sg13g2_buf_1  input30
timestamp 1676381911
transform 1 0 1536 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  input31
timestamp 1676381911
transform 1 0 1152 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  input32
timestamp 1676381911
transform 1 0 1536 0 -1 4536
box -48 -56 432 834
use sg13g2_buf_1  input33
timestamp 1676381911
transform 1 0 3168 0 1 1512
box -48 -56 432 834
use sg13g2_buf_1  input34
timestamp 1676381911
transform 1 0 3936 0 1 1512
box -48 -56 432 834
use sg13g2_buf_1  input35
timestamp 1676381911
transform 1 0 10848 0 1 1512
box -48 -56 432 834
use sg13g2_buf_1  input36
timestamp 1676381911
transform 1 0 11424 0 1 1512
box -48 -56 432 834
use sg13g2_buf_1  input37
timestamp 1676381911
transform 1 0 11808 0 1 1512
box -48 -56 432 834
use sg13g2_buf_1  input38
timestamp 1676381911
transform -1 0 12576 0 1 1512
box -48 -56 432 834
use sg13g2_buf_1  input39
timestamp 1676381911
transform 1 0 14304 0 1 1512
box -48 -56 432 834
use sg13g2_buf_1  input40
timestamp 1676381911
transform 1 0 14688 0 1 1512
box -48 -56 432 834
use sg13g2_buf_1  input41
timestamp 1676381911
transform 1 0 4512 0 1 1512
box -48 -56 432 834
use sg13g2_buf_1  input42
timestamp 1676381911
transform 1 0 4896 0 1 1512
box -48 -56 432 834
use sg13g2_buf_1  input43
timestamp 1676381911
transform 1 0 5280 0 1 1512
box -48 -56 432 834
use sg13g2_buf_1  input44
timestamp 1676381911
transform 1 0 5664 0 1 1512
box -48 -56 432 834
use sg13g2_buf_1  input45
timestamp 1676381911
transform 1 0 6048 0 1 1512
box -48 -56 432 834
use sg13g2_buf_1  input46
timestamp 1676381911
transform 1 0 8640 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  input47
timestamp 1676381911
transform 1 0 8448 0 1 1512
box -48 -56 432 834
use sg13g2_buf_1  input48
timestamp 1676381911
transform 1 0 8832 0 1 1512
box -48 -56 432 834
use sg13g2_buf_1  input49
timestamp 1676381911
transform -1 0 18912 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  input50
timestamp 1676381911
transform -1 0 20832 0 1 7560
box -48 -56 432 834
use sg13g2_buf_1  input51
timestamp 1676381911
transform 1 0 18912 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  input52
timestamp 1676381911
transform -1 0 21216 0 1 7560
box -48 -56 432 834
use sg13g2_buf_1  input53
timestamp 1676381911
transform -1 0 22848 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  input54
timestamp 1676381911
transform -1 0 23232 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  input55
timestamp 1676381911
transform 1 0 23232 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  input56
timestamp 1676381911
transform -1 0 24000 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  input57
timestamp 1676381911
transform -1 0 24384 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  input58
timestamp 1676381911
transform -1 0 25728 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  input59
timestamp 1676381911
transform 1 0 25728 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  input60
timestamp 1676381911
transform 1 0 26112 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  input61
timestamp 1676381911
transform 1 0 22464 0 -1 7560
box -48 -56 432 834
use sg13g2_buf_1  input62
timestamp 1676381911
transform -1 0 21600 0 1 7560
box -48 -56 432 834
use sg13g2_buf_1  input63
timestamp 1676381911
transform 1 0 21600 0 1 7560
box -48 -56 432 834
use sg13g2_buf_1  input64
timestamp 1676381911
transform 1 0 20544 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  input65
timestamp 1676381911
transform -1 0 21312 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  input66
timestamp 1676381911
transform -1 0 21696 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  input67
timestamp 1676381911
transform 1 0 21696 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  input68
timestamp 1676381911
transform -1 0 22464 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  input69
timestamp 1676381911
transform 1 0 25056 0 -1 7560
box -48 -56 432 834
use sg13g2_buf_1  input70
timestamp 1676381911
transform 1 0 26976 0 -1 7560
box -48 -56 432 834
use sg13g2_buf_1  input71
timestamp 1676381911
transform 1 0 29952 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  input72
timestamp 1676381911
transform -1 0 31104 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  input73
timestamp 1676381911
transform -1 0 31488 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  input74
timestamp 1676381911
transform 1 0 31488 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  input75
timestamp 1676381911
transform -1 0 28320 0 1 6048
box -48 -56 432 834
use sg13g2_buf_1  input76
timestamp 1676381911
transform -1 0 28416 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  input77
timestamp 1676381911
transform 1 0 26016 0 -1 7560
box -48 -56 432 834
use sg13g2_buf_1  input78
timestamp 1676381911
transform -1 0 28800 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  input79
timestamp 1676381911
transform -1 0 28032 0 -1 9072
box -48 -56 432 834
use sg13g2_buf_1  input80
timestamp 1676381911
transform -1 0 29184 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  input81
timestamp 1676381911
transform 1 0 28032 0 -1 9072
box -48 -56 432 834
use sg13g2_buf_1  input82
timestamp 1676381911
transform -1 0 29568 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  input83
timestamp 1676381911
transform -1 0 28800 0 -1 9072
box -48 -56 432 834
use sg13g2_buf_1  input84
timestamp 1676381911
transform -1 0 29952 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  input85
timestamp 1676381911
transform -1 0 30240 0 1 7560
box -48 -56 432 834
use sg13g2_buf_1  input86
timestamp 1676381911
transform 1 0 32640 0 -1 7560
box -48 -56 432 834
use sg13g2_buf_1  input87
timestamp 1676381911
transform 1 0 33024 0 -1 7560
box -48 -56 432 834
use sg13g2_buf_1  input88
timestamp 1676381911
transform -1 0 36096 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  input89
timestamp 1676381911
transform -1 0 35616 0 -1 9072
box -48 -56 432 834
use sg13g2_buf_1  input90
timestamp 1676381911
transform 1 0 34560 0 1 7560
box -48 -56 432 834
use sg13g2_buf_1  input91
timestamp 1676381911
transform -1 0 34176 0 -1 7560
box -48 -56 432 834
use sg13g2_buf_1  input92
timestamp 1676381911
transform -1 0 32256 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  input93
timestamp 1676381911
transform 1 0 30240 0 1 7560
box -48 -56 432 834
use sg13g2_buf_1  input94
timestamp 1676381911
transform -1 0 32640 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  input95
timestamp 1676381911
transform -1 0 31008 0 1 7560
box -48 -56 432 834
use sg13g2_buf_1  input96
timestamp 1676381911
transform -1 0 30240 0 -1 7560
box -48 -56 432 834
use sg13g2_buf_1  input97
timestamp 1676381911
transform 1 0 32256 0 -1 9072
box -48 -56 432 834
use sg13g2_buf_1  input98
timestamp 1676381911
transform -1 0 33024 0 -1 9072
box -48 -56 432 834
use sg13g2_buf_1  input99
timestamp 1676381911
transform -1 0 34656 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  input100
timestamp 1676381911
transform -1 0 32640 0 -1 7560
box -48 -56 432 834
use sg13g2_buf_1  output101
timestamp 1676381911
transform 1 0 43296 0 1 1512
box -48 -56 432 834
use sg13g2_buf_1  output102
timestamp 1676381911
transform 1 0 44448 0 -1 4536
box -48 -56 432 834
use sg13g2_buf_1  output103
timestamp 1676381911
transform 1 0 44832 0 -1 4536
box -48 -56 432 834
use sg13g2_buf_1  output104
timestamp 1676381911
transform 1 0 44448 0 1 4536
box -48 -56 432 834
use sg13g2_buf_1  output105
timestamp 1676381911
transform 1 0 44832 0 1 4536
box -48 -56 432 834
use sg13g2_buf_1  output106
timestamp 1676381911
transform 1 0 44448 0 -1 6048
box -48 -56 432 834
use sg13g2_buf_1  output107
timestamp 1676381911
transform 1 0 44832 0 -1 6048
box -48 -56 432 834
use sg13g2_buf_1  output108
timestamp 1676381911
transform 1 0 44448 0 1 6048
box -48 -56 432 834
use sg13g2_buf_1  output109
timestamp 1676381911
transform 1 0 44832 0 1 6048
box -48 -56 432 834
use sg13g2_buf_1  output110
timestamp 1676381911
transform 1 0 44448 0 -1 7560
box -48 -56 432 834
use sg13g2_buf_1  output111
timestamp 1676381911
transform 1 0 44832 0 -1 7560
box -48 -56 432 834
use sg13g2_buf_1  output112
timestamp 1676381911
transform 1 0 42912 0 1 1512
box -48 -56 432 834
use sg13g2_buf_1  output113
timestamp 1676381911
transform 1 0 44832 0 1 7560
box -48 -56 432 834
use sg13g2_buf_1  output114
timestamp 1676381911
transform 1 0 44448 0 1 7560
box -48 -56 432 834
use sg13g2_buf_1  output115
timestamp 1676381911
transform 1 0 44832 0 -1 9072
box -48 -56 432 834
use sg13g2_buf_1  output116
timestamp 1676381911
transform 1 0 44448 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  output117
timestamp 1676381911
transform 1 0 43008 0 -1 9072
box -48 -56 432 834
use sg13g2_buf_1  output118
timestamp 1676381911
transform 1 0 42528 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  output119
timestamp 1676381911
transform 1 0 43680 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  output120
timestamp 1676381911
transform 1 0 44064 0 -1 9072
box -48 -56 432 834
use sg13g2_buf_1  output121
timestamp 1676381911
transform 1 0 44064 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  output122
timestamp 1676381911
transform 1 0 42912 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  output123
timestamp 1676381911
transform 1 0 43296 0 -1 3024
box -48 -56 432 834
use sg13g2_buf_1  output124
timestamp 1676381911
transform 1 0 43392 0 -1 9072
box -48 -56 432 834
use sg13g2_buf_1  output125
timestamp 1676381911
transform 1 0 44064 0 1 7560
box -48 -56 432 834
use sg13g2_buf_1  output126
timestamp 1676381911
transform 1 0 43680 0 1 1512
box -48 -56 432 834
use sg13g2_buf_1  output127
timestamp 1676381911
transform 1 0 43680 0 -1 3024
box -48 -56 432 834
use sg13g2_buf_1  output128
timestamp 1676381911
transform 1 0 42528 0 1 1512
box -48 -56 432 834
use sg13g2_buf_1  output129
timestamp 1676381911
transform 1 0 44832 0 1 1512
box -48 -56 432 834
use sg13g2_buf_1  output130
timestamp 1676381911
transform 1 0 44448 0 -1 3024
box -48 -56 432 834
use sg13g2_buf_1  output131
timestamp 1676381911
transform 1 0 44832 0 -1 3024
box -48 -56 432 834
use sg13g2_buf_1  output132
timestamp 1676381911
transform 1 0 44832 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  output133
timestamp 1676381911
transform -1 0 36480 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  output134
timestamp 1676381911
transform -1 0 37920 0 -1 9072
box -48 -56 432 834
use sg13g2_buf_1  output135
timestamp 1676381911
transform -1 0 38784 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  output136
timestamp 1676381911
transform -1 0 36672 0 -1 7560
box -48 -56 432 834
use sg13g2_buf_1  output137
timestamp 1676381911
transform -1 0 38304 0 -1 9072
box -48 -56 432 834
use sg13g2_buf_1  output138
timestamp 1676381911
transform -1 0 39168 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  output139
timestamp 1676381911
transform -1 0 37056 0 -1 7560
box -48 -56 432 834
use sg13g2_buf_1  output140
timestamp 1676381911
transform -1 0 39552 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  output141
timestamp 1676381911
transform -1 0 38688 0 -1 9072
box -48 -56 432 834
use sg13g2_buf_1  output142
timestamp 1676381911
transform -1 0 39936 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  output143
timestamp 1676381911
transform -1 0 36000 0 -1 6048
box -48 -56 432 834
use sg13g2_buf_1  output144
timestamp 1676381911
transform -1 0 32832 0 -1 6048
box -48 -56 432 834
use sg13g2_buf_1  output145
timestamp 1676381911
transform -1 0 36864 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  output146
timestamp 1676381911
transform -1 0 33216 0 -1 6048
box -48 -56 432 834
use sg13g2_buf_1  output147
timestamp 1676381911
transform -1 0 37248 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  output148
timestamp 1676381911
transform -1 0 37632 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  output149
timestamp 1676381911
transform -1 0 36480 0 1 7560
box -48 -56 432 834
use sg13g2_buf_1  output150
timestamp 1676381911
transform -1 0 38016 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  output151
timestamp 1676381911
transform -1 0 36864 0 1 7560
box -48 -56 432 834
use sg13g2_buf_1  output152
timestamp 1676381911
transform -1 0 38400 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  output153
timestamp 1676381911
transform -1 0 15744 0 1 1512
box -48 -56 432 834
use sg13g2_buf_1  output154
timestamp 1676381911
transform 1 0 15744 0 1 1512
box -48 -56 432 834
use sg13g2_buf_1  output155
timestamp 1676381911
transform -1 0 23424 0 1 1512
box -48 -56 432 834
use sg13g2_buf_1  output156
timestamp 1676381911
transform 1 0 23424 0 1 1512
box -48 -56 432 834
use sg13g2_buf_1  output157
timestamp 1676381911
transform -1 0 25920 0 1 1512
box -48 -56 432 834
use sg13g2_buf_1  output158
timestamp 1676381911
transform -1 0 25824 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  output159
timestamp 1676381911
transform -1 0 28032 0 -1 3024
box -48 -56 432 834
use sg13g2_buf_1  output160
timestamp 1676381911
transform -1 0 30144 0 1 1512
box -48 -56 432 834
use sg13g2_buf_1  output161
timestamp 1676381911
transform 1 0 16128 0 1 1512
box -48 -56 432 834
use sg13g2_buf_1  output162
timestamp 1676381911
transform -1 0 18144 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  output163
timestamp 1676381911
transform 1 0 17664 0 -1 3024
box -48 -56 432 834
use sg13g2_buf_1  output164
timestamp 1676381911
transform 1 0 18528 0 1 1512
box -48 -56 432 834
use sg13g2_buf_1  output165
timestamp 1676381911
transform 1 0 18912 0 1 1512
box -48 -56 432 834
use sg13g2_buf_1  output166
timestamp 1676381911
transform 1 0 19776 0 1 1512
box -48 -56 432 834
use sg13g2_buf_1  output167
timestamp 1676381911
transform 1 0 20160 0 1 1512
box -48 -56 432 834
use sg13g2_buf_1  output168
timestamp 1676381911
transform -1 0 22752 0 1 1512
box -48 -56 432 834
use sg13g2_buf_1  output169
timestamp 1676381911
transform 1 0 8448 0 -1 7560
box -48 -56 432 834
use sg13g2_buf_1  output170
timestamp 1676381911
transform 1 0 8832 0 -1 7560
box -48 -56 432 834
use sg13g2_buf_1  output171
timestamp 1676381911
transform -1 0 11808 0 1 4536
box -48 -56 432 834
use sg13g2_buf_1  output172
timestamp 1676381911
transform 1 0 9792 0 1 6048
box -48 -56 432 834
use sg13g2_buf_1  output173
timestamp 1676381911
transform 1 0 7872 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  output174
timestamp 1676381911
transform 1 0 9408 0 1 7560
box -48 -56 432 834
use sg13g2_buf_1  output175
timestamp 1676381911
transform 1 0 9792 0 1 7560
box -48 -56 432 834
use sg13g2_buf_1  output176
timestamp 1676381911
transform -1 0 12768 0 -1 6048
box -48 -56 432 834
use sg13g2_buf_1  output177
timestamp 1676381911
transform 1 0 12192 0 1 6048
box -48 -56 432 834
use sg13g2_buf_1  output178
timestamp 1676381911
transform 1 0 11616 0 -1 7560
box -48 -56 432 834
use sg13g2_buf_1  output179
timestamp 1676381911
transform 1 0 9216 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  output180
timestamp 1676381911
transform 1 0 12576 0 1 6048
box -48 -56 432 834
use sg13g2_buf_1  output181
timestamp 1676381911
transform 1 0 9600 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  output182
timestamp 1676381911
transform 1 0 12000 0 -1 7560
box -48 -56 432 834
use sg13g2_buf_1  output183
timestamp 1676381911
transform 1 0 11520 0 1 7560
box -48 -56 432 834
use sg13g2_buf_1  output184
timestamp 1676381911
transform 1 0 12384 0 -1 7560
box -48 -56 432 834
use sg13g2_buf_1  output185
timestamp 1676381911
transform 1 0 11904 0 1 7560
box -48 -56 432 834
use sg13g2_buf_1  output186
timestamp 1676381911
transform 1 0 12768 0 -1 7560
box -48 -56 432 834
use sg13g2_buf_1  output187
timestamp 1676381911
transform 1 0 13152 0 -1 7560
box -48 -56 432 834
use sg13g2_buf_1  output188
timestamp 1676381911
transform 1 0 13536 0 -1 7560
box -48 -56 432 834
use sg13g2_buf_1  output189
timestamp 1676381911
transform 1 0 13920 0 -1 7560
box -48 -56 432 834
use sg13g2_buf_1  output190
timestamp 1676381911
transform 1 0 15456 0 -1 7560
box -48 -56 432 834
use sg13g2_buf_1  output191
timestamp 1676381911
transform 1 0 15840 0 -1 7560
box -48 -56 432 834
use sg13g2_buf_1  output192
timestamp 1676381911
transform 1 0 16224 0 -1 7560
box -48 -56 432 834
use sg13g2_buf_1  output193
timestamp 1676381911
transform -1 0 17760 0 1 6048
box -48 -56 432 834
use sg13g2_buf_1  output194
timestamp 1676381911
transform 1 0 14208 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  output195
timestamp 1676381911
transform -1 0 18144 0 1 6048
box -48 -56 432 834
use sg13g2_buf_1  output196
timestamp 1676381911
transform 1 0 11232 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  output197
timestamp 1676381911
transform -1 0 15648 0 1 6048
box -48 -56 432 834
use sg13g2_buf_1  output198
timestamp 1676381911
transform 1 0 11616 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  output199
timestamp 1676381911
transform 1 0 12864 0 -1 9072
box -48 -56 432 834
use sg13g2_buf_1  output200
timestamp 1676381911
transform 1 0 12000 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  output201
timestamp 1676381911
transform 1 0 14688 0 -1 7560
box -48 -56 432 834
use sg13g2_buf_1  output202
timestamp 1676381911
transform 1 0 13248 0 -1 9072
box -48 -56 432 834
use sg13g2_buf_1  output203
timestamp 1676381911
transform 1 0 15072 0 -1 7560
box -48 -56 432 834
use sg13g2_buf_1  output204
timestamp 1676381911
transform 1 0 13632 0 -1 9072
box -48 -56 432 834
use sg13g2_buf_1  output205
timestamp 1676381911
transform 1 0 16128 0 1 7560
box -48 -56 432 834
use sg13g2_buf_1  output206
timestamp 1676381911
transform 1 0 19200 0 -1 7560
box -48 -56 432 834
use sg13g2_buf_1  output207
timestamp 1676381911
transform 1 0 17952 0 -1 9072
box -48 -56 432 834
use sg13g2_buf_1  output208
timestamp 1676381911
transform 1 0 19584 0 -1 7560
box -48 -56 432 834
use sg13g2_buf_1  output209
timestamp 1676381911
transform 1 0 18336 0 -1 9072
box -48 -56 432 834
use sg13g2_buf_1  output210
timestamp 1676381911
transform 1 0 17760 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  output211
timestamp 1676381911
transform -1 0 21120 0 -1 7560
box -48 -56 432 834
use sg13g2_buf_1  output212
timestamp 1676381911
transform 1 0 14592 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  output213
timestamp 1676381911
transform 1 0 16512 0 1 7560
box -48 -56 432 834
use sg13g2_buf_1  output214
timestamp 1676381911
transform 1 0 14976 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  output215
timestamp 1676381911
transform 1 0 15840 0 -1 9072
box -48 -56 432 834
use sg13g2_buf_1  output216
timestamp 1676381911
transform 1 0 18144 0 1 6048
box -48 -56 432 834
use sg13g2_buf_1  output217
timestamp 1676381911
transform 1 0 15360 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  output218
timestamp 1676381911
transform 1 0 16896 0 1 7560
box -48 -56 432 834
use sg13g2_buf_1  output219
timestamp 1676381911
transform 1 0 15744 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  output220
timestamp 1676381911
transform 1 0 18816 0 -1 7560
box -48 -56 432 834
use sg13g2_buf_1  output221
timestamp 1676381911
transform -1 0 32448 0 -1 6048
box -48 -56 432 834
use sg13g2_tielo  S_CPU_IF_222
timestamp 1680000637
transform 1 0 18144 0 1 9072
box -48 -56 432 834
<< labels >>
flabel metal3 s 20984 11764 21064 11844 0 FreeSans 320 0 0 0 Co
port 0 nsew signal output
flabel metal2 s 0 548 90 628 0 FreeSans 320 0 0 0 FrameData[0]
port 1 nsew signal input
flabel metal2 s 0 3908 90 3988 0 FreeSans 320 0 0 0 FrameData[10]
port 2 nsew signal input
flabel metal2 s 0 4244 90 4324 0 FreeSans 320 0 0 0 FrameData[11]
port 3 nsew signal input
flabel metal2 s 0 4580 90 4660 0 FreeSans 320 0 0 0 FrameData[12]
port 4 nsew signal input
flabel metal2 s 0 4916 90 4996 0 FreeSans 320 0 0 0 FrameData[13]
port 5 nsew signal input
flabel metal2 s 0 5252 90 5332 0 FreeSans 320 0 0 0 FrameData[14]
port 6 nsew signal input
flabel metal2 s 0 5588 90 5668 0 FreeSans 320 0 0 0 FrameData[15]
port 7 nsew signal input
flabel metal2 s 0 5924 90 6004 0 FreeSans 320 0 0 0 FrameData[16]
port 8 nsew signal input
flabel metal2 s 0 6260 90 6340 0 FreeSans 320 0 0 0 FrameData[17]
port 9 nsew signal input
flabel metal2 s 0 6596 90 6676 0 FreeSans 320 0 0 0 FrameData[18]
port 10 nsew signal input
flabel metal2 s 0 6932 90 7012 0 FreeSans 320 0 0 0 FrameData[19]
port 11 nsew signal input
flabel metal2 s 0 884 90 964 0 FreeSans 320 0 0 0 FrameData[1]
port 12 nsew signal input
flabel metal2 s 0 7268 90 7348 0 FreeSans 320 0 0 0 FrameData[20]
port 13 nsew signal input
flabel metal2 s 0 7604 90 7684 0 FreeSans 320 0 0 0 FrameData[21]
port 14 nsew signal input
flabel metal2 s 0 7940 90 8020 0 FreeSans 320 0 0 0 FrameData[22]
port 15 nsew signal input
flabel metal2 s 0 8276 90 8356 0 FreeSans 320 0 0 0 FrameData[23]
port 16 nsew signal input
flabel metal2 s 0 8612 90 8692 0 FreeSans 320 0 0 0 FrameData[24]
port 17 nsew signal input
flabel metal2 s 0 8948 90 9028 0 FreeSans 320 0 0 0 FrameData[25]
port 18 nsew signal input
flabel metal2 s 0 9284 90 9364 0 FreeSans 320 0 0 0 FrameData[26]
port 19 nsew signal input
flabel metal2 s 0 9620 90 9700 0 FreeSans 320 0 0 0 FrameData[27]
port 20 nsew signal input
flabel metal2 s 0 9956 90 10036 0 FreeSans 320 0 0 0 FrameData[28]
port 21 nsew signal input
flabel metal2 s 0 10292 90 10372 0 FreeSans 320 0 0 0 FrameData[29]
port 22 nsew signal input
flabel metal2 s 0 1220 90 1300 0 FreeSans 320 0 0 0 FrameData[2]
port 23 nsew signal input
flabel metal2 s 0 10628 90 10708 0 FreeSans 320 0 0 0 FrameData[30]
port 24 nsew signal input
flabel metal2 s 0 10964 90 11044 0 FreeSans 320 0 0 0 FrameData[31]
port 25 nsew signal input
flabel metal2 s 0 1556 90 1636 0 FreeSans 320 0 0 0 FrameData[3]
port 26 nsew signal input
flabel metal2 s 0 1892 90 1972 0 FreeSans 320 0 0 0 FrameData[4]
port 27 nsew signal input
flabel metal2 s 0 2228 90 2308 0 FreeSans 320 0 0 0 FrameData[5]
port 28 nsew signal input
flabel metal2 s 0 2564 90 2644 0 FreeSans 320 0 0 0 FrameData[6]
port 29 nsew signal input
flabel metal2 s 0 2900 90 2980 0 FreeSans 320 0 0 0 FrameData[7]
port 30 nsew signal input
flabel metal2 s 0 3236 90 3316 0 FreeSans 320 0 0 0 FrameData[8]
port 31 nsew signal input
flabel metal2 s 0 3572 90 3652 0 FreeSans 320 0 0 0 FrameData[9]
port 32 nsew signal input
flabel metal2 s 46278 548 46368 628 0 FreeSans 320 0 0 0 FrameData_O[0]
port 33 nsew signal output
flabel metal2 s 46278 3908 46368 3988 0 FreeSans 320 0 0 0 FrameData_O[10]
port 34 nsew signal output
flabel metal2 s 46278 4244 46368 4324 0 FreeSans 320 0 0 0 FrameData_O[11]
port 35 nsew signal output
flabel metal2 s 46278 4580 46368 4660 0 FreeSans 320 0 0 0 FrameData_O[12]
port 36 nsew signal output
flabel metal2 s 46278 4916 46368 4996 0 FreeSans 320 0 0 0 FrameData_O[13]
port 37 nsew signal output
flabel metal2 s 46278 5252 46368 5332 0 FreeSans 320 0 0 0 FrameData_O[14]
port 38 nsew signal output
flabel metal2 s 46278 5588 46368 5668 0 FreeSans 320 0 0 0 FrameData_O[15]
port 39 nsew signal output
flabel metal2 s 46278 5924 46368 6004 0 FreeSans 320 0 0 0 FrameData_O[16]
port 40 nsew signal output
flabel metal2 s 46278 6260 46368 6340 0 FreeSans 320 0 0 0 FrameData_O[17]
port 41 nsew signal output
flabel metal2 s 46278 6596 46368 6676 0 FreeSans 320 0 0 0 FrameData_O[18]
port 42 nsew signal output
flabel metal2 s 46278 6932 46368 7012 0 FreeSans 320 0 0 0 FrameData_O[19]
port 43 nsew signal output
flabel metal2 s 46278 884 46368 964 0 FreeSans 320 0 0 0 FrameData_O[1]
port 44 nsew signal output
flabel metal2 s 46278 7268 46368 7348 0 FreeSans 320 0 0 0 FrameData_O[20]
port 45 nsew signal output
flabel metal2 s 46278 7604 46368 7684 0 FreeSans 320 0 0 0 FrameData_O[21]
port 46 nsew signal output
flabel metal2 s 46278 7940 46368 8020 0 FreeSans 320 0 0 0 FrameData_O[22]
port 47 nsew signal output
flabel metal2 s 46278 8276 46368 8356 0 FreeSans 320 0 0 0 FrameData_O[23]
port 48 nsew signal output
flabel metal2 s 46278 8612 46368 8692 0 FreeSans 320 0 0 0 FrameData_O[24]
port 49 nsew signal output
flabel metal2 s 46278 8948 46368 9028 0 FreeSans 320 0 0 0 FrameData_O[25]
port 50 nsew signal output
flabel metal2 s 46278 9284 46368 9364 0 FreeSans 320 0 0 0 FrameData_O[26]
port 51 nsew signal output
flabel metal2 s 46278 9620 46368 9700 0 FreeSans 320 0 0 0 FrameData_O[27]
port 52 nsew signal output
flabel metal2 s 46278 9956 46368 10036 0 FreeSans 320 0 0 0 FrameData_O[28]
port 53 nsew signal output
flabel metal2 s 46278 10292 46368 10372 0 FreeSans 320 0 0 0 FrameData_O[29]
port 54 nsew signal output
flabel metal2 s 46278 1220 46368 1300 0 FreeSans 320 0 0 0 FrameData_O[2]
port 55 nsew signal output
flabel metal2 s 46278 10628 46368 10708 0 FreeSans 320 0 0 0 FrameData_O[30]
port 56 nsew signal output
flabel metal2 s 46278 10964 46368 11044 0 FreeSans 320 0 0 0 FrameData_O[31]
port 57 nsew signal output
flabel metal2 s 46278 1556 46368 1636 0 FreeSans 320 0 0 0 FrameData_O[3]
port 58 nsew signal output
flabel metal2 s 46278 1892 46368 1972 0 FreeSans 320 0 0 0 FrameData_O[4]
port 59 nsew signal output
flabel metal2 s 46278 2228 46368 2308 0 FreeSans 320 0 0 0 FrameData_O[5]
port 60 nsew signal output
flabel metal2 s 46278 2564 46368 2644 0 FreeSans 320 0 0 0 FrameData_O[6]
port 61 nsew signal output
flabel metal2 s 46278 2900 46368 2980 0 FreeSans 320 0 0 0 FrameData_O[7]
port 62 nsew signal output
flabel metal2 s 46278 3236 46368 3316 0 FreeSans 320 0 0 0 FrameData_O[8]
port 63 nsew signal output
flabel metal2 s 46278 3572 46368 3652 0 FreeSans 320 0 0 0 FrameData_O[9]
port 64 nsew signal output
flabel metal3 s 28472 0 28552 80 0 FreeSans 320 0 0 0 FrameStrobe[0]
port 65 nsew signal input
flabel metal3 s 36152 0 36232 80 0 FreeSans 320 0 0 0 FrameStrobe[10]
port 66 nsew signal input
flabel metal3 s 36920 0 37000 80 0 FreeSans 320 0 0 0 FrameStrobe[11]
port 67 nsew signal input
flabel metal3 s 37688 0 37768 80 0 FreeSans 320 0 0 0 FrameStrobe[12]
port 68 nsew signal input
flabel metal3 s 38456 0 38536 80 0 FreeSans 320 0 0 0 FrameStrobe[13]
port 69 nsew signal input
flabel metal3 s 39224 0 39304 80 0 FreeSans 320 0 0 0 FrameStrobe[14]
port 70 nsew signal input
flabel metal3 s 39992 0 40072 80 0 FreeSans 320 0 0 0 FrameStrobe[15]
port 71 nsew signal input
flabel metal3 s 40760 0 40840 80 0 FreeSans 320 0 0 0 FrameStrobe[16]
port 72 nsew signal input
flabel metal3 s 41528 0 41608 80 0 FreeSans 320 0 0 0 FrameStrobe[17]
port 73 nsew signal input
flabel metal3 s 42296 0 42376 80 0 FreeSans 320 0 0 0 FrameStrobe[18]
port 74 nsew signal input
flabel metal3 s 43064 0 43144 80 0 FreeSans 320 0 0 0 FrameStrobe[19]
port 75 nsew signal input
flabel metal3 s 29240 0 29320 80 0 FreeSans 320 0 0 0 FrameStrobe[1]
port 76 nsew signal input
flabel metal3 s 30008 0 30088 80 0 FreeSans 320 0 0 0 FrameStrobe[2]
port 77 nsew signal input
flabel metal3 s 30776 0 30856 80 0 FreeSans 320 0 0 0 FrameStrobe[3]
port 78 nsew signal input
flabel metal3 s 31544 0 31624 80 0 FreeSans 320 0 0 0 FrameStrobe[4]
port 79 nsew signal input
flabel metal3 s 32312 0 32392 80 0 FreeSans 320 0 0 0 FrameStrobe[5]
port 80 nsew signal input
flabel metal3 s 33080 0 33160 80 0 FreeSans 320 0 0 0 FrameStrobe[6]
port 81 nsew signal input
flabel metal3 s 33848 0 33928 80 0 FreeSans 320 0 0 0 FrameStrobe[7]
port 82 nsew signal input
flabel metal3 s 34616 0 34696 80 0 FreeSans 320 0 0 0 FrameStrobe[8]
port 83 nsew signal input
flabel metal3 s 35384 0 35464 80 0 FreeSans 320 0 0 0 FrameStrobe[9]
port 84 nsew signal input
flabel metal3 s 31352 11764 31432 11844 0 FreeSans 320 0 0 0 FrameStrobe_O[0]
port 85 nsew signal output
flabel metal3 s 33272 11764 33352 11844 0 FreeSans 320 0 0 0 FrameStrobe_O[10]
port 86 nsew signal output
flabel metal3 s 33464 11764 33544 11844 0 FreeSans 320 0 0 0 FrameStrobe_O[11]
port 87 nsew signal output
flabel metal3 s 33656 11764 33736 11844 0 FreeSans 320 0 0 0 FrameStrobe_O[12]
port 88 nsew signal output
flabel metal3 s 33848 11764 33928 11844 0 FreeSans 320 0 0 0 FrameStrobe_O[13]
port 89 nsew signal output
flabel metal3 s 34040 11764 34120 11844 0 FreeSans 320 0 0 0 FrameStrobe_O[14]
port 90 nsew signal output
flabel metal3 s 34232 11764 34312 11844 0 FreeSans 320 0 0 0 FrameStrobe_O[15]
port 91 nsew signal output
flabel metal3 s 34424 11764 34504 11844 0 FreeSans 320 0 0 0 FrameStrobe_O[16]
port 92 nsew signal output
flabel metal3 s 34616 11764 34696 11844 0 FreeSans 320 0 0 0 FrameStrobe_O[17]
port 93 nsew signal output
flabel metal3 s 34808 11764 34888 11844 0 FreeSans 320 0 0 0 FrameStrobe_O[18]
port 94 nsew signal output
flabel metal3 s 35000 11764 35080 11844 0 FreeSans 320 0 0 0 FrameStrobe_O[19]
port 95 nsew signal output
flabel metal3 s 31544 11764 31624 11844 0 FreeSans 320 0 0 0 FrameStrobe_O[1]
port 96 nsew signal output
flabel metal3 s 31736 11764 31816 11844 0 FreeSans 320 0 0 0 FrameStrobe_O[2]
port 97 nsew signal output
flabel metal3 s 31928 11764 32008 11844 0 FreeSans 320 0 0 0 FrameStrobe_O[3]
port 98 nsew signal output
flabel metal3 s 32120 11764 32200 11844 0 FreeSans 320 0 0 0 FrameStrobe_O[4]
port 99 nsew signal output
flabel metal3 s 32312 11764 32392 11844 0 FreeSans 320 0 0 0 FrameStrobe_O[5]
port 100 nsew signal output
flabel metal3 s 32504 11764 32584 11844 0 FreeSans 320 0 0 0 FrameStrobe_O[6]
port 101 nsew signal output
flabel metal3 s 32696 11764 32776 11844 0 FreeSans 320 0 0 0 FrameStrobe_O[7]
port 102 nsew signal output
flabel metal3 s 32888 11764 32968 11844 0 FreeSans 320 0 0 0 FrameStrobe_O[8]
port 103 nsew signal output
flabel metal3 s 33080 11764 33160 11844 0 FreeSans 320 0 0 0 FrameStrobe_O[9]
port 104 nsew signal output
flabel metal3 s 15416 0 15496 80 0 FreeSans 320 0 0 0 I_top0
port 105 nsew signal output
flabel metal3 s 16184 0 16264 80 0 FreeSans 320 0 0 0 I_top1
port 106 nsew signal output
flabel metal3 s 23096 0 23176 80 0 FreeSans 320 0 0 0 I_top10
port 107 nsew signal output
flabel metal3 s 23864 0 23944 80 0 FreeSans 320 0 0 0 I_top11
port 108 nsew signal output
flabel metal3 s 24632 0 24712 80 0 FreeSans 320 0 0 0 I_top12
port 109 nsew signal output
flabel metal3 s 25400 0 25480 80 0 FreeSans 320 0 0 0 I_top13
port 110 nsew signal output
flabel metal3 s 26168 0 26248 80 0 FreeSans 320 0 0 0 I_top14
port 111 nsew signal output
flabel metal3 s 26936 0 27016 80 0 FreeSans 320 0 0 0 I_top15
port 112 nsew signal output
flabel metal3 s 16952 0 17032 80 0 FreeSans 320 0 0 0 I_top2
port 113 nsew signal output
flabel metal3 s 17720 0 17800 80 0 FreeSans 320 0 0 0 I_top3
port 114 nsew signal output
flabel metal3 s 18488 0 18568 80 0 FreeSans 320 0 0 0 I_top4
port 115 nsew signal output
flabel metal3 s 19256 0 19336 80 0 FreeSans 320 0 0 0 I_top5
port 116 nsew signal output
flabel metal3 s 20024 0 20104 80 0 FreeSans 320 0 0 0 I_top6
port 117 nsew signal output
flabel metal3 s 20792 0 20872 80 0 FreeSans 320 0 0 0 I_top7
port 118 nsew signal output
flabel metal3 s 21560 0 21640 80 0 FreeSans 320 0 0 0 I_top8
port 119 nsew signal output
flabel metal3 s 22328 0 22408 80 0 FreeSans 320 0 0 0 I_top9
port 120 nsew signal output
flabel metal3 s 11000 11764 11080 11844 0 FreeSans 320 0 0 0 N1BEG[0]
port 121 nsew signal output
flabel metal3 s 11192 11764 11272 11844 0 FreeSans 320 0 0 0 N1BEG[1]
port 122 nsew signal output
flabel metal3 s 11384 11764 11464 11844 0 FreeSans 320 0 0 0 N1BEG[2]
port 123 nsew signal output
flabel metal3 s 11576 11764 11656 11844 0 FreeSans 320 0 0 0 N1BEG[3]
port 124 nsew signal output
flabel metal3 s 11768 11764 11848 11844 0 FreeSans 320 0 0 0 N2BEG[0]
port 125 nsew signal output
flabel metal3 s 11960 11764 12040 11844 0 FreeSans 320 0 0 0 N2BEG[1]
port 126 nsew signal output
flabel metal3 s 12152 11764 12232 11844 0 FreeSans 320 0 0 0 N2BEG[2]
port 127 nsew signal output
flabel metal3 s 12344 11764 12424 11844 0 FreeSans 320 0 0 0 N2BEG[3]
port 128 nsew signal output
flabel metal3 s 12536 11764 12616 11844 0 FreeSans 320 0 0 0 N2BEG[4]
port 129 nsew signal output
flabel metal3 s 12728 11764 12808 11844 0 FreeSans 320 0 0 0 N2BEG[5]
port 130 nsew signal output
flabel metal3 s 12920 11764 13000 11844 0 FreeSans 320 0 0 0 N2BEG[6]
port 131 nsew signal output
flabel metal3 s 13112 11764 13192 11844 0 FreeSans 320 0 0 0 N2BEG[7]
port 132 nsew signal output
flabel metal3 s 13304 11764 13384 11844 0 FreeSans 320 0 0 0 N2BEGb[0]
port 133 nsew signal output
flabel metal3 s 13496 11764 13576 11844 0 FreeSans 320 0 0 0 N2BEGb[1]
port 134 nsew signal output
flabel metal3 s 13688 11764 13768 11844 0 FreeSans 320 0 0 0 N2BEGb[2]
port 135 nsew signal output
flabel metal3 s 13880 11764 13960 11844 0 FreeSans 320 0 0 0 N2BEGb[3]
port 136 nsew signal output
flabel metal3 s 14072 11764 14152 11844 0 FreeSans 320 0 0 0 N2BEGb[4]
port 137 nsew signal output
flabel metal3 s 14264 11764 14344 11844 0 FreeSans 320 0 0 0 N2BEGb[5]
port 138 nsew signal output
flabel metal3 s 14456 11764 14536 11844 0 FreeSans 320 0 0 0 N2BEGb[6]
port 139 nsew signal output
flabel metal3 s 14648 11764 14728 11844 0 FreeSans 320 0 0 0 N2BEGb[7]
port 140 nsew signal output
flabel metal3 s 14840 11764 14920 11844 0 FreeSans 320 0 0 0 N4BEG[0]
port 141 nsew signal output
flabel metal3 s 16760 11764 16840 11844 0 FreeSans 320 0 0 0 N4BEG[10]
port 142 nsew signal output
flabel metal3 s 16952 11764 17032 11844 0 FreeSans 320 0 0 0 N4BEG[11]
port 143 nsew signal output
flabel metal3 s 17144 11764 17224 11844 0 FreeSans 320 0 0 0 N4BEG[12]
port 144 nsew signal output
flabel metal3 s 17336 11764 17416 11844 0 FreeSans 320 0 0 0 N4BEG[13]
port 145 nsew signal output
flabel metal3 s 17528 11764 17608 11844 0 FreeSans 320 0 0 0 N4BEG[14]
port 146 nsew signal output
flabel metal3 s 17720 11764 17800 11844 0 FreeSans 320 0 0 0 N4BEG[15]
port 147 nsew signal output
flabel metal3 s 15032 11764 15112 11844 0 FreeSans 320 0 0 0 N4BEG[1]
port 148 nsew signal output
flabel metal3 s 15224 11764 15304 11844 0 FreeSans 320 0 0 0 N4BEG[2]
port 149 nsew signal output
flabel metal3 s 15416 11764 15496 11844 0 FreeSans 320 0 0 0 N4BEG[3]
port 150 nsew signal output
flabel metal3 s 15608 11764 15688 11844 0 FreeSans 320 0 0 0 N4BEG[4]
port 151 nsew signal output
flabel metal3 s 15800 11764 15880 11844 0 FreeSans 320 0 0 0 N4BEG[5]
port 152 nsew signal output
flabel metal3 s 15992 11764 16072 11844 0 FreeSans 320 0 0 0 N4BEG[6]
port 153 nsew signal output
flabel metal3 s 16184 11764 16264 11844 0 FreeSans 320 0 0 0 N4BEG[7]
port 154 nsew signal output
flabel metal3 s 16376 11764 16456 11844 0 FreeSans 320 0 0 0 N4BEG[8]
port 155 nsew signal output
flabel metal3 s 16568 11764 16648 11844 0 FreeSans 320 0 0 0 N4BEG[9]
port 156 nsew signal output
flabel metal3 s 17912 11764 17992 11844 0 FreeSans 320 0 0 0 NN4BEG[0]
port 157 nsew signal output
flabel metal3 s 19832 11764 19912 11844 0 FreeSans 320 0 0 0 NN4BEG[10]
port 158 nsew signal output
flabel metal3 s 20024 11764 20104 11844 0 FreeSans 320 0 0 0 NN4BEG[11]
port 159 nsew signal output
flabel metal3 s 20216 11764 20296 11844 0 FreeSans 320 0 0 0 NN4BEG[12]
port 160 nsew signal output
flabel metal3 s 20408 11764 20488 11844 0 FreeSans 320 0 0 0 NN4BEG[13]
port 161 nsew signal output
flabel metal3 s 20600 11764 20680 11844 0 FreeSans 320 0 0 0 NN4BEG[14]
port 162 nsew signal output
flabel metal3 s 20792 11764 20872 11844 0 FreeSans 320 0 0 0 NN4BEG[15]
port 163 nsew signal output
flabel metal3 s 18104 11764 18184 11844 0 FreeSans 320 0 0 0 NN4BEG[1]
port 164 nsew signal output
flabel metal3 s 18296 11764 18376 11844 0 FreeSans 320 0 0 0 NN4BEG[2]
port 165 nsew signal output
flabel metal3 s 18488 11764 18568 11844 0 FreeSans 320 0 0 0 NN4BEG[3]
port 166 nsew signal output
flabel metal3 s 18680 11764 18760 11844 0 FreeSans 320 0 0 0 NN4BEG[4]
port 167 nsew signal output
flabel metal3 s 18872 11764 18952 11844 0 FreeSans 320 0 0 0 NN4BEG[5]
port 168 nsew signal output
flabel metal3 s 19064 11764 19144 11844 0 FreeSans 320 0 0 0 NN4BEG[6]
port 169 nsew signal output
flabel metal3 s 19256 11764 19336 11844 0 FreeSans 320 0 0 0 NN4BEG[7]
port 170 nsew signal output
flabel metal3 s 19448 11764 19528 11844 0 FreeSans 320 0 0 0 NN4BEG[8]
port 171 nsew signal output
flabel metal3 s 19640 11764 19720 11844 0 FreeSans 320 0 0 0 NN4BEG[9]
port 172 nsew signal output
flabel metal3 s 3128 0 3208 80 0 FreeSans 320 0 0 0 O_top0
port 173 nsew signal input
flabel metal3 s 3896 0 3976 80 0 FreeSans 320 0 0 0 O_top1
port 174 nsew signal input
flabel metal3 s 10808 0 10888 80 0 FreeSans 320 0 0 0 O_top10
port 175 nsew signal input
flabel metal3 s 11576 0 11656 80 0 FreeSans 320 0 0 0 O_top11
port 176 nsew signal input
flabel metal3 s 12344 0 12424 80 0 FreeSans 320 0 0 0 O_top12
port 177 nsew signal input
flabel metal3 s 13112 0 13192 80 0 FreeSans 320 0 0 0 O_top13
port 178 nsew signal input
flabel metal3 s 13880 0 13960 80 0 FreeSans 320 0 0 0 O_top14
port 179 nsew signal input
flabel metal3 s 14648 0 14728 80 0 FreeSans 320 0 0 0 O_top15
port 180 nsew signal input
flabel metal3 s 4664 0 4744 80 0 FreeSans 320 0 0 0 O_top2
port 181 nsew signal input
flabel metal3 s 5432 0 5512 80 0 FreeSans 320 0 0 0 O_top3
port 182 nsew signal input
flabel metal3 s 6200 0 6280 80 0 FreeSans 320 0 0 0 O_top4
port 183 nsew signal input
flabel metal3 s 6968 0 7048 80 0 FreeSans 320 0 0 0 O_top5
port 184 nsew signal input
flabel metal3 s 7736 0 7816 80 0 FreeSans 320 0 0 0 O_top6
port 185 nsew signal input
flabel metal3 s 8504 0 8584 80 0 FreeSans 320 0 0 0 O_top7
port 186 nsew signal input
flabel metal3 s 9272 0 9352 80 0 FreeSans 320 0 0 0 O_top8
port 187 nsew signal input
flabel metal3 s 10040 0 10120 80 0 FreeSans 320 0 0 0 O_top9
port 188 nsew signal input
flabel metal3 s 21176 11764 21256 11844 0 FreeSans 320 0 0 0 S1END[0]
port 189 nsew signal input
flabel metal3 s 21368 11764 21448 11844 0 FreeSans 320 0 0 0 S1END[1]
port 190 nsew signal input
flabel metal3 s 21560 11764 21640 11844 0 FreeSans 320 0 0 0 S1END[2]
port 191 nsew signal input
flabel metal3 s 21752 11764 21832 11844 0 FreeSans 320 0 0 0 S1END[3]
port 192 nsew signal input
flabel metal3 s 23480 11764 23560 11844 0 FreeSans 320 0 0 0 S2END[0]
port 193 nsew signal input
flabel metal3 s 23672 11764 23752 11844 0 FreeSans 320 0 0 0 S2END[1]
port 194 nsew signal input
flabel metal3 s 23864 11764 23944 11844 0 FreeSans 320 0 0 0 S2END[2]
port 195 nsew signal input
flabel metal3 s 24056 11764 24136 11844 0 FreeSans 320 0 0 0 S2END[3]
port 196 nsew signal input
flabel metal3 s 24248 11764 24328 11844 0 FreeSans 320 0 0 0 S2END[4]
port 197 nsew signal input
flabel metal3 s 24440 11764 24520 11844 0 FreeSans 320 0 0 0 S2END[5]
port 198 nsew signal input
flabel metal3 s 24632 11764 24712 11844 0 FreeSans 320 0 0 0 S2END[6]
port 199 nsew signal input
flabel metal3 s 24824 11764 24904 11844 0 FreeSans 320 0 0 0 S2END[7]
port 200 nsew signal input
flabel metal3 s 21944 11764 22024 11844 0 FreeSans 320 0 0 0 S2MID[0]
port 201 nsew signal input
flabel metal3 s 22136 11764 22216 11844 0 FreeSans 320 0 0 0 S2MID[1]
port 202 nsew signal input
flabel metal3 s 22328 11764 22408 11844 0 FreeSans 320 0 0 0 S2MID[2]
port 203 nsew signal input
flabel metal3 s 22520 11764 22600 11844 0 FreeSans 320 0 0 0 S2MID[3]
port 204 nsew signal input
flabel metal3 s 22712 11764 22792 11844 0 FreeSans 320 0 0 0 S2MID[4]
port 205 nsew signal input
flabel metal3 s 22904 11764 22984 11844 0 FreeSans 320 0 0 0 S2MID[5]
port 206 nsew signal input
flabel metal3 s 23096 11764 23176 11844 0 FreeSans 320 0 0 0 S2MID[6]
port 207 nsew signal input
flabel metal3 s 23288 11764 23368 11844 0 FreeSans 320 0 0 0 S2MID[7]
port 208 nsew signal input
flabel metal3 s 25016 11764 25096 11844 0 FreeSans 320 0 0 0 S4END[0]
port 209 nsew signal input
flabel metal3 s 26936 11764 27016 11844 0 FreeSans 320 0 0 0 S4END[10]
port 210 nsew signal input
flabel metal3 s 27128 11764 27208 11844 0 FreeSans 320 0 0 0 S4END[11]
port 211 nsew signal input
flabel metal3 s 27320 11764 27400 11844 0 FreeSans 320 0 0 0 S4END[12]
port 212 nsew signal input
flabel metal3 s 27512 11764 27592 11844 0 FreeSans 320 0 0 0 S4END[13]
port 213 nsew signal input
flabel metal3 s 27704 11764 27784 11844 0 FreeSans 320 0 0 0 S4END[14]
port 214 nsew signal input
flabel metal3 s 27896 11764 27976 11844 0 FreeSans 320 0 0 0 S4END[15]
port 215 nsew signal input
flabel metal3 s 25208 11764 25288 11844 0 FreeSans 320 0 0 0 S4END[1]
port 216 nsew signal input
flabel metal3 s 25400 11764 25480 11844 0 FreeSans 320 0 0 0 S4END[2]
port 217 nsew signal input
flabel metal3 s 25592 11764 25672 11844 0 FreeSans 320 0 0 0 S4END[3]
port 218 nsew signal input
flabel metal3 s 25784 11764 25864 11844 0 FreeSans 320 0 0 0 S4END[4]
port 219 nsew signal input
flabel metal3 s 25976 11764 26056 11844 0 FreeSans 320 0 0 0 S4END[5]
port 220 nsew signal input
flabel metal3 s 26168 11764 26248 11844 0 FreeSans 320 0 0 0 S4END[6]
port 221 nsew signal input
flabel metal3 s 26360 11764 26440 11844 0 FreeSans 320 0 0 0 S4END[7]
port 222 nsew signal input
flabel metal3 s 26552 11764 26632 11844 0 FreeSans 320 0 0 0 S4END[8]
port 223 nsew signal input
flabel metal3 s 26744 11764 26824 11844 0 FreeSans 320 0 0 0 S4END[9]
port 224 nsew signal input
flabel metal3 s 28088 11764 28168 11844 0 FreeSans 320 0 0 0 SS4END[0]
port 225 nsew signal input
flabel metal3 s 30008 11764 30088 11844 0 FreeSans 320 0 0 0 SS4END[10]
port 226 nsew signal input
flabel metal3 s 30200 11764 30280 11844 0 FreeSans 320 0 0 0 SS4END[11]
port 227 nsew signal input
flabel metal3 s 30392 11764 30472 11844 0 FreeSans 320 0 0 0 SS4END[12]
port 228 nsew signal input
flabel metal3 s 30584 11764 30664 11844 0 FreeSans 320 0 0 0 SS4END[13]
port 229 nsew signal input
flabel metal3 s 30776 11764 30856 11844 0 FreeSans 320 0 0 0 SS4END[14]
port 230 nsew signal input
flabel metal3 s 30968 11764 31048 11844 0 FreeSans 320 0 0 0 SS4END[15]
port 231 nsew signal input
flabel metal3 s 28280 11764 28360 11844 0 FreeSans 320 0 0 0 SS4END[1]
port 232 nsew signal input
flabel metal3 s 28472 11764 28552 11844 0 FreeSans 320 0 0 0 SS4END[2]
port 233 nsew signal input
flabel metal3 s 28664 11764 28744 11844 0 FreeSans 320 0 0 0 SS4END[3]
port 234 nsew signal input
flabel metal3 s 28856 11764 28936 11844 0 FreeSans 320 0 0 0 SS4END[4]
port 235 nsew signal input
flabel metal3 s 29048 11764 29128 11844 0 FreeSans 320 0 0 0 SS4END[5]
port 236 nsew signal input
flabel metal3 s 29240 11764 29320 11844 0 FreeSans 320 0 0 0 SS4END[6]
port 237 nsew signal input
flabel metal3 s 29432 11764 29512 11844 0 FreeSans 320 0 0 0 SS4END[7]
port 238 nsew signal input
flabel metal3 s 29624 11764 29704 11844 0 FreeSans 320 0 0 0 SS4END[8]
port 239 nsew signal input
flabel metal3 s 29816 11764 29896 11844 0 FreeSans 320 0 0 0 SS4END[9]
port 240 nsew signal input
flabel metal3 s 27704 0 27784 80 0 FreeSans 320 0 0 0 UserCLK
port 241 nsew signal input
flabel metal3 s 31160 11764 31240 11844 0 FreeSans 320 0 0 0 UserCLKo
port 242 nsew signal output
flabel metal5 s 4892 0 5332 11844 0 FreeSans 2560 90 0 0 VGND
port 243 nsew ground bidirectional
flabel metal5 s 4892 0 5332 40 0 FreeSans 320 0 0 0 VGND
port 243 nsew ground bidirectional
flabel metal5 s 4892 11804 5332 11844 0 FreeSans 320 0 0 0 VGND
port 243 nsew ground bidirectional
flabel metal5 s 20012 0 20452 11844 0 FreeSans 2560 90 0 0 VGND
port 243 nsew ground bidirectional
flabel metal5 s 20012 0 20452 40 0 FreeSans 320 0 0 0 VGND
port 243 nsew ground bidirectional
flabel metal5 s 20012 11804 20452 11844 0 FreeSans 320 0 0 0 VGND
port 243 nsew ground bidirectional
flabel metal5 s 35132 0 35572 11844 0 FreeSans 2560 90 0 0 VGND
port 243 nsew ground bidirectional
flabel metal5 s 35132 0 35572 40 0 FreeSans 320 0 0 0 VGND
port 243 nsew ground bidirectional
flabel metal5 s 35132 11804 35572 11844 0 FreeSans 320 0 0 0 VGND
port 243 nsew ground bidirectional
flabel metal5 s 3652 0 4092 11844 0 FreeSans 2560 90 0 0 VPWR
port 244 nsew power bidirectional
flabel metal5 s 3652 0 4092 40 0 FreeSans 320 0 0 0 VPWR
port 244 nsew power bidirectional
flabel metal5 s 3652 11804 4092 11844 0 FreeSans 320 0 0 0 VPWR
port 244 nsew power bidirectional
flabel metal5 s 18772 0 19212 11844 0 FreeSans 2560 90 0 0 VPWR
port 244 nsew power bidirectional
flabel metal5 s 18772 0 19212 40 0 FreeSans 320 0 0 0 VPWR
port 244 nsew power bidirectional
flabel metal5 s 18772 11804 19212 11844 0 FreeSans 320 0 0 0 VPWR
port 244 nsew power bidirectional
flabel metal5 s 33892 0 34332 11844 0 FreeSans 2560 90 0 0 VPWR
port 244 nsew power bidirectional
flabel metal5 s 33892 0 34332 40 0 FreeSans 320 0 0 0 VPWR
port 244 nsew power bidirectional
flabel metal5 s 33892 11804 34332 11844 0 FreeSans 320 0 0 0 VPWR
port 244 nsew power bidirectional
rlabel metal1 23184 9072 23184 9072 0 VGND
rlabel metal1 23184 9828 23184 9828 0 VPWR
rlabel metal2 752 588 752 588 0 FrameData[0]
rlabel via2 80 3948 80 3948 0 FrameData[10]
rlabel metal2 848 4284 848 4284 0 FrameData[11]
rlabel via2 80 4620 80 4620 0 FrameData[12]
rlabel metal2 560 4956 560 4956 0 FrameData[13]
rlabel metal2 128 5292 128 5292 0 FrameData[14]
rlabel metal2 656 5628 656 5628 0 FrameData[15]
rlabel metal2 128 5964 128 5964 0 FrameData[16]
rlabel via2 80 6300 80 6300 0 FrameData[17]
rlabel metal2 128 6636 128 6636 0 FrameData[18]
rlabel via2 80 6972 80 6972 0 FrameData[19]
rlabel metal2 704 924 704 924 0 FrameData[1]
rlabel metal2 656 7308 656 7308 0 FrameData[20]
rlabel metal2 464 7644 464 7644 0 FrameData[21]
rlabel metal2 368 7980 368 7980 0 FrameData[22]
rlabel metal2 848 8316 848 8316 0 FrameData[23]
rlabel metal2 560 8652 560 8652 0 FrameData[24]
rlabel metal2 656 8988 656 8988 0 FrameData[25]
rlabel metal2 848 9324 848 9324 0 FrameData[26]
rlabel metal2 1040 9660 1040 9660 0 FrameData[27]
rlabel metal2 656 9996 656 9996 0 FrameData[28]
rlabel metal2 752 10332 752 10332 0 FrameData[29]
rlabel metal2 656 1260 656 1260 0 FrameData[2]
rlabel metal2 608 10668 608 10668 0 FrameData[30]
rlabel metal2 704 11004 704 11004 0 FrameData[31]
rlabel via2 80 1596 80 1596 0 FrameData[3]
rlabel metal2 128 1932 128 1932 0 FrameData[4]
rlabel metal2 848 2268 848 2268 0 FrameData[5]
rlabel metal2 656 2604 656 2604 0 FrameData[6]
rlabel metal2 80 2940 80 2940 0 FrameData[7]
rlabel via2 80 3276 80 3276 0 FrameData[8]
rlabel metal2 848 3612 848 3612 0 FrameData[9]
rlabel metal2 45663 588 45663 588 0 FrameData_O[0]
rlabel metal2 45951 3948 45951 3948 0 FrameData_O[10]
rlabel metal2 45735 4284 45735 4284 0 FrameData_O[11]
rlabel metal2 45543 4620 45543 4620 0 FrameData_O[12]
rlabel metal2 45735 4956 45735 4956 0 FrameData_O[13]
rlabel via2 46287 5292 46287 5292 0 FrameData_O[14]
rlabel metal2 45735 5628 45735 5628 0 FrameData_O[15]
rlabel via2 46287 5964 46287 5964 0 FrameData_O[16]
rlabel metal2 45735 6300 45735 6300 0 FrameData_O[17]
rlabel via2 46287 6636 46287 6636 0 FrameData_O[18]
rlabel metal2 45735 6972 45735 6972 0 FrameData_O[19]
rlabel metal2 45567 924 45567 924 0 FrameData_O[1]
rlabel metal2 46047 7308 46047 7308 0 FrameData_O[20]
rlabel metal2 45543 7644 45543 7644 0 FrameData_O[21]
rlabel metal2 46047 7980 46047 7980 0 FrameData_O[22]
rlabel metal2 45663 8316 45663 8316 0 FrameData_O[23]
rlabel metal2 45663 8652 45663 8652 0 FrameData_O[24]
rlabel metal2 44655 8988 44655 8988 0 FrameData_O[25]
rlabel metal2 45735 9324 45735 9324 0 FrameData_O[26]
rlabel metal2 44808 8904 44808 8904 0 FrameData_O[27]
rlabel metal2 44424 9660 44424 9660 0 FrameData_O[28]
rlabel metal2 43272 9660 43272 9660 0 FrameData_O[29]
rlabel metal2 45471 1260 45471 1260 0 FrameData_O[2]
rlabel metal2 43992 8904 43992 8904 0 FrameData_O[30]
rlabel metal2 44568 8148 44568 8148 0 FrameData_O[31]
rlabel metal2 46239 1596 46239 1596 0 FrameData_O[3]
rlabel metal2 45711 1932 45711 1932 0 FrameData_O[4]
rlabel metal2 44736 2184 44736 2184 0 FrameData_O[5]
rlabel metal2 45192 2016 45192 2016 0 FrameData_O[6]
rlabel metal2 45192 2772 45192 2772 0 FrameData_O[7]
rlabel metal2 45192 2856 45192 2856 0 FrameData_O[8]
rlabel metal2 45735 3612 45735 3612 0 FrameData_O[9]
rlabel metal2 20352 4998 20352 4998 0 FrameStrobe[0]
rlabel metal3 36192 996 36192 996 0 FrameStrobe[10]
rlabel metal3 36960 1878 36960 1878 0 FrameStrobe[11]
rlabel metal3 37728 996 37728 996 0 FrameStrobe[12]
rlabel metal3 38496 114 38496 114 0 FrameStrobe[13]
rlabel metal3 39264 1752 39264 1752 0 FrameStrobe[14]
rlabel metal2 40608 8736 40608 8736 0 FrameStrobe[15]
rlabel metal3 40800 2928 40800 2928 0 FrameStrobe[16]
rlabel via3 41568 72 41568 72 0 FrameStrobe[17]
rlabel metal2 41808 9492 41808 9492 0 FrameStrobe[18]
rlabel metal3 43104 912 43104 912 0 FrameStrobe[19]
rlabel metal3 14880 1524 14880 1524 0 FrameStrobe[1]
rlabel metal2 38496 8946 38496 8946 0 FrameStrobe[2]
rlabel metal3 41952 2478 41952 2478 0 FrameStrobe[3]
rlabel metal3 33408 2478 33408 2478 0 FrameStrobe[4]
rlabel metal2 35232 2814 35232 2814 0 FrameStrobe[5]
rlabel metal2 43200 2478 43200 2478 0 FrameStrobe[6]
rlabel via3 33888 72 33888 72 0 FrameStrobe[7]
rlabel metal3 34656 912 34656 912 0 FrameStrobe[8]
rlabel metal3 35424 114 35424 114 0 FrameStrobe[9]
rlabel metal2 36168 9576 36168 9576 0 FrameStrobe_O[0]
rlabel metal2 36936 8652 36936 8652 0 FrameStrobe_O[10]
rlabel metal2 38328 9240 38328 9240 0 FrameStrobe_O[11]
rlabel metal2 36360 6972 36360 6972 0 FrameStrobe_O[12]
rlabel metal2 37944 8652 37944 8652 0 FrameStrobe_O[13]
rlabel metal2 38808 9660 38808 9660 0 FrameStrobe_O[14]
rlabel metal2 36600 6972 36600 6972 0 FrameStrobe_O[15]
rlabel metal2 39192 9660 39192 9660 0 FrameStrobe_O[16]
rlabel metal2 37272 8904 37272 8904 0 FrameStrobe_O[17]
rlabel metal2 39288 9324 39288 9324 0 FrameStrobe_O[18]
rlabel metal2 35400 5460 35400 5460 0 FrameStrobe_O[19]
rlabel metal2 32496 5922 32496 5922 0 FrameStrobe_O[1]
rlabel metal2 36504 9576 36504 9576 0 FrameStrobe_O[2]
rlabel metal2 32856 5460 32856 5460 0 FrameStrobe_O[3]
rlabel metal2 36336 9660 36336 9660 0 FrameStrobe_O[4]
rlabel metal2 37272 9660 37272 9660 0 FrameStrobe_O[5]
rlabel metal2 35448 7980 35448 7980 0 FrameStrobe_O[6]
rlabel metal2 37608 9240 37608 9240 0 FrameStrobe_O[7]
rlabel metal2 35784 8064 35784 8064 0 FrameStrobe_O[8]
rlabel metal2 37944 9240 37944 9240 0 FrameStrobe_O[9]
rlabel metal3 15456 870 15456 870 0 I_top0
rlabel metal3 16224 870 16224 870 0 I_top1
rlabel metal3 23136 870 23136 870 0 I_top10
rlabel metal3 23904 870 23904 870 0 I_top11
rlabel metal3 24672 912 24672 912 0 I_top12
rlabel metal2 25464 3192 25464 3192 0 I_top13
rlabel metal3 26208 1290 26208 1290 0 I_top14
rlabel metal3 26976 870 26976 870 0 I_top15
rlabel metal3 16992 912 16992 912 0 I_top2
rlabel metal2 17784 3192 17784 3192 0 I_top3
rlabel metal3 18528 1248 18528 1248 0 I_top4
rlabel metal3 19296 828 19296 828 0 I_top5
rlabel metal3 20064 114 20064 114 0 I_top6
rlabel metal3 20832 450 20832 450 0 I_top7
rlabel metal3 21600 870 21600 870 0 I_top8
rlabel metal3 22368 870 22368 870 0 I_top9
rlabel metal2 28080 2688 28080 2688 0 Inst_S_CPU_IF_ConfigMem.Inst_frame0_bit0.Q
rlabel metal2 30288 2688 30288 2688 0 Inst_S_CPU_IF_ConfigMem.Inst_frame0_bit1.Q
rlabel metal2 10305 6383 10305 6383 0 Inst_S_CPU_IF_ConfigMem.Inst_frame0_bit10.Q
rlabel metal2 12312 6384 12312 6384 0 Inst_S_CPU_IF_ConfigMem.Inst_frame0_bit11.Q
rlabel metal3 31968 3864 31968 3864 0 Inst_S_CPU_IF_ConfigMem.Inst_frame0_bit12.Q
rlabel metal2 34224 2856 34224 2856 0 Inst_S_CPU_IF_ConfigMem.Inst_frame0_bit13.Q
rlabel metal2 7776 9156 7776 9156 0 Inst_S_CPU_IF_ConfigMem.Inst_frame0_bit14.Q
rlabel metal3 20640 7518 20640 7518 0 Inst_S_CPU_IF_ConfigMem.Inst_frame0_bit15.Q
rlabel metal2 23136 2730 23136 2730 0 Inst_S_CPU_IF_ConfigMem.Inst_frame0_bit16.Q
rlabel metal2 24672 2646 24672 2646 0 Inst_S_CPU_IF_ConfigMem.Inst_frame0_bit17.Q
rlabel metal2 8736 8736 8736 8736 0 Inst_S_CPU_IF_ConfigMem.Inst_frame0_bit18.Q
rlabel metal2 10896 8736 10896 8736 0 Inst_S_CPU_IF_ConfigMem.Inst_frame0_bit19.Q
rlabel metal2 7104 4242 7104 4242 0 Inst_S_CPU_IF_ConfigMem.Inst_frame0_bit2.Q
rlabel metal2 39009 6384 39009 6384 0 Inst_S_CPU_IF_ConfigMem.Inst_frame0_bit20.Q
rlabel via2 40616 6384 40616 6384 0 Inst_S_CPU_IF_ConfigMem.Inst_frame0_bit21.Q
rlabel metal2 27888 7896 27888 7896 0 Inst_S_CPU_IF_ConfigMem.Inst_frame0_bit22.Q
rlabel metal2 29480 7896 29480 7896 0 Inst_S_CPU_IF_ConfigMem.Inst_frame0_bit23.Q
rlabel metal2 15168 3402 15168 3402 0 Inst_S_CPU_IF_ConfigMem.Inst_frame0_bit24.Q
rlabel metal2 16704 3465 16704 3465 0 Inst_S_CPU_IF_ConfigMem.Inst_frame0_bit25.Q
rlabel metal2 5760 6426 5760 6426 0 Inst_S_CPU_IF_ConfigMem.Inst_frame0_bit26.Q
rlabel metal2 7512 6384 7512 6384 0 Inst_S_CPU_IF_ConfigMem.Inst_frame0_bit27.Q
rlabel metal2 34464 7476 34464 7476 0 Inst_S_CPU_IF_ConfigMem.Inst_frame0_bit28.Q
rlabel metal3 36000 6930 36000 6930 0 Inst_S_CPU_IF_ConfigMem.Inst_frame0_bit29.Q
rlabel metal2 8832 2856 8832 2856 0 Inst_S_CPU_IF_ConfigMem.Inst_frame0_bit3.Q
rlabel metal2 20016 5544 20016 5544 0 Inst_S_CPU_IF_ConfigMem.Inst_frame0_bit30.Q
rlabel metal2 24552 6384 24552 6384 0 Inst_S_CPU_IF_ConfigMem.Inst_frame0_bit31.Q
rlabel metal2 37872 3360 37872 3360 0 Inst_S_CPU_IF_ConfigMem.Inst_frame0_bit4.Q
rlabel metal2 39960 3360 39960 3360 0 Inst_S_CPU_IF_ConfigMem.Inst_frame0_bit5.Q
rlabel metal2 15552 8946 15552 8946 0 Inst_S_CPU_IF_ConfigMem.Inst_frame0_bit6.Q
rlabel metal2 26016 8148 26016 8148 0 Inst_S_CPU_IF_ConfigMem.Inst_frame0_bit7.Q
rlabel metal2 19248 2772 19248 2772 0 Inst_S_CPU_IF_ConfigMem.Inst_frame0_bit8.Q
rlabel metal2 20688 2100 20688 2100 0 Inst_S_CPU_IF_ConfigMem.Inst_frame0_bit9.Q
rlabel metal2 23376 5712 23376 5712 0 Inst_S_CPU_IF_ConfigMem.Inst_frame1_bit0.Q
rlabel metal2 34416 6384 34416 6384 0 Inst_S_CPU_IF_ConfigMem.Inst_frame1_bit1.Q
rlabel metal2 13248 5628 13248 5628 0 Inst_S_CPU_IF_ConfigMem.Inst_frame1_bit10.Q
rlabel metal2 18384 4704 18384 4704 0 Inst_S_CPU_IF_ConfigMem.Inst_frame1_bit11.Q
rlabel metal3 24576 8946 24576 8946 0 Inst_S_CPU_IF_ConfigMem.Inst_frame1_bit12.Q
rlabel metal3 34944 2394 34944 2394 0 Inst_S_CPU_IF_ConfigMem.Inst_frame1_bit13.Q
rlabel metal2 7344 2856 7344 2856 0 Inst_S_CPU_IF_ConfigMem.Inst_frame1_bit14.Q
rlabel metal2 28032 1806 28032 1806 0 Inst_S_CPU_IF_ConfigMem.Inst_frame1_bit15.Q
rlabel metal3 22944 6972 22944 6972 0 Inst_S_CPU_IF_ConfigMem.Inst_frame1_bit16.Q
rlabel metal2 35136 7896 35136 7896 0 Inst_S_CPU_IF_ConfigMem.Inst_frame1_bit17.Q
rlabel metal3 5472 5166 5472 5166 0 Inst_S_CPU_IF_ConfigMem.Inst_frame1_bit18.Q
rlabel metal2 13008 3360 13008 3360 0 Inst_S_CPU_IF_ConfigMem.Inst_frame1_bit19.Q
rlabel metal2 6384 4872 6384 4872 0 Inst_S_CPU_IF_ConfigMem.Inst_frame1_bit2.Q
rlabel metal3 33312 8442 33312 8442 0 Inst_S_CPU_IF_ConfigMem.Inst_frame1_bit20.Q
rlabel metal2 41232 6384 41232 6384 0 Inst_S_CPU_IF_ConfigMem.Inst_frame1_bit21.Q
rlabel metal2 11664 7896 11664 7896 0 Inst_S_CPU_IF_ConfigMem.Inst_frame1_bit22.Q
rlabel metal2 25776 3948 25776 3948 0 Inst_S_CPU_IF_ConfigMem.Inst_frame1_bit23.Q
rlabel metal2 19152 9408 19152 9408 0 Inst_S_CPU_IF_ConfigMem.Inst_frame1_bit24.Q
rlabel metal2 32880 4872 32880 4872 0 Inst_S_CPU_IF_ConfigMem.Inst_frame1_bit25.Q
rlabel metal2 9216 7224 9216 7224 0 Inst_S_CPU_IF_ConfigMem.Inst_frame1_bit26.Q
rlabel metal2 17568 3360 17568 3360 0 Inst_S_CPU_IF_ConfigMem.Inst_frame1_bit27.Q
rlabel metal3 29088 8988 29088 8988 0 Inst_S_CPU_IF_ConfigMem.Inst_frame1_bit28.Q
rlabel metal2 38256 2688 38256 2688 0 Inst_S_CPU_IF_ConfigMem.Inst_frame1_bit29.Q
rlabel metal2 13728 2730 13728 2730 0 Inst_S_CPU_IF_ConfigMem.Inst_frame1_bit3.Q
rlabel metal2 15072 4662 15072 4662 0 Inst_S_CPU_IF_ConfigMem.Inst_frame1_bit30.Q
rlabel metal2 28224 2856 28224 2856 0 Inst_S_CPU_IF_ConfigMem.Inst_frame1_bit31.Q
rlabel metal3 36000 9156 36000 9156 0 Inst_S_CPU_IF_ConfigMem.Inst_frame1_bit4.Q
rlabel metal3 42144 6132 42144 6132 0 Inst_S_CPU_IF_ConfigMem.Inst_frame1_bit5.Q
rlabel metal2 10752 9366 10752 9366 0 Inst_S_CPU_IF_ConfigMem.Inst_frame1_bit6.Q
rlabel metal2 24048 3360 24048 3360 0 Inst_S_CPU_IF_ConfigMem.Inst_frame1_bit7.Q
rlabel metal2 19392 7854 19392 7854 0 Inst_S_CPU_IF_ConfigMem.Inst_frame1_bit8.Q
rlabel metal2 22800 4704 22800 4704 0 Inst_S_CPU_IF_ConfigMem.Inst_frame1_bit9.Q
rlabel metal2 31872 5754 31872 5754 0 Inst_S_CPU_IF_ConfigMem.Inst_frame2_bit10.Q
rlabel metal2 34896 5712 34896 5712 0 Inst_S_CPU_IF_ConfigMem.Inst_frame2_bit11.Q
rlabel metal2 9168 4872 9168 4872 0 Inst_S_CPU_IF_ConfigMem.Inst_frame2_bit12.Q
rlabel metal2 11064 4872 11064 4872 0 Inst_S_CPU_IF_ConfigMem.Inst_frame2_bit13.Q
rlabel metal2 13248 1890 13248 1890 0 Inst_S_CPU_IF_ConfigMem.Inst_frame2_bit14.Q
rlabel metal2 16992 2142 16992 2142 0 Inst_S_CPU_IF_ConfigMem.Inst_frame2_bit15.Q
rlabel metal2 21408 5544 21408 5544 0 Inst_S_CPU_IF_ConfigMem.Inst_frame2_bit16.Q
rlabel metal2 33504 6384 33504 6384 0 Inst_S_CPU_IF_ConfigMem.Inst_frame2_bit17.Q
rlabel metal3 5664 5964 5664 5964 0 Inst_S_CPU_IF_ConfigMem.Inst_frame2_bit18.Q
rlabel metal3 15648 4284 15648 4284 0 Inst_S_CPU_IF_ConfigMem.Inst_frame2_bit19.Q
rlabel metal2 26880 8694 26880 8694 0 Inst_S_CPU_IF_ConfigMem.Inst_frame2_bit20.Q
rlabel metal2 38904 4200 38904 4200 0 Inst_S_CPU_IF_ConfigMem.Inst_frame2_bit21.Q
rlabel metal2 9936 5712 9936 5712 0 Inst_S_CPU_IF_ConfigMem.Inst_frame2_bit22.Q
rlabel metal2 29040 3948 29040 3948 0 Inst_S_CPU_IF_ConfigMem.Inst_frame2_bit23.Q
rlabel metal2 22176 7854 22176 7854 0 Inst_S_CPU_IF_ConfigMem.Inst_frame2_bit24.Q
rlabel metal2 36240 5124 36240 5124 0 Inst_S_CPU_IF_ConfigMem.Inst_frame2_bit25.Q
rlabel metal2 8640 8904 8640 8904 0 Inst_S_CPU_IF_ConfigMem.Inst_frame2_bit26.Q
rlabel metal3 12864 2142 12864 2142 0 Inst_S_CPU_IF_ConfigMem.Inst_frame2_bit27.Q
rlabel metal2 34320 8736 34320 8736 0 Inst_S_CPU_IF_ConfigMem.Inst_frame2_bit28.Q
rlabel metal2 40128 4872 40128 4872 0 Inst_S_CPU_IF_ConfigMem.Inst_frame2_bit29.Q
rlabel metal2 15744 5418 15744 5418 0 Inst_S_CPU_IF_ConfigMem.Inst_frame2_bit30.Q
rlabel metal2 24096 4032 24096 4032 0 Inst_S_CPU_IF_ConfigMem.Inst_frame2_bit31.Q
rlabel metal2 18768 6972 18768 6972 0 Inst_S_CPU_IF_ConfigMem.Inst_frame2_bit8.Q
rlabel metal3 22368 6510 22368 6510 0 Inst_S_CPU_IF_ConfigMem.Inst_frame2_bit9.Q
rlabel metal3 23232 8442 23232 8442 0 Inst_S_CPU_IF_switch_matrix.N1BEG0
rlabel metal2 36288 5670 36288 5670 0 Inst_S_CPU_IF_switch_matrix.N1BEG1
rlabel metal3 11040 4410 11040 4410 0 Inst_S_CPU_IF_switch_matrix.N1BEG2
rlabel metal2 17064 2436 17064 2436 0 Inst_S_CPU_IF_switch_matrix.N1BEG3
rlabel metal2 22368 7098 22368 7098 0 Inst_S_CPU_IF_switch_matrix.N2BEG0
rlabel metal2 34272 4956 34272 4956 0 Inst_S_CPU_IF_switch_matrix.N2BEG1
rlabel metal3 6336 6342 6336 6342 0 Inst_S_CPU_IF_switch_matrix.N2BEG2
rlabel metal3 14880 3696 14880 3696 0 Inst_S_CPU_IF_switch_matrix.N2BEG3
rlabel metal2 27648 7140 27648 7140 0 Inst_S_CPU_IF_switch_matrix.N2BEG4
rlabel metal2 40032 4074 40032 4074 0 Inst_S_CPU_IF_switch_matrix.N2BEG5
rlabel metal3 9024 4788 9024 4788 0 Inst_S_CPU_IF_switch_matrix.N2BEG6
rlabel metal2 30768 2604 30768 2604 0 Inst_S_CPU_IF_switch_matrix.N2BEG7
rlabel metal2 23616 8022 23616 8022 0 Inst_S_CPU_IF_switch_matrix.N2BEGb0
rlabel metal3 37440 6090 37440 6090 0 Inst_S_CPU_IF_switch_matrix.N2BEGb1
rlabel metal3 8160 8358 8160 8358 0 Inst_S_CPU_IF_switch_matrix.N2BEGb2
rlabel metal2 14016 1932 14016 1932 0 Inst_S_CPU_IF_switch_matrix.N2BEGb3
rlabel metal2 38976 8736 38976 8736 0 Inst_S_CPU_IF_switch_matrix.N2BEGb4
rlabel metal3 42048 4578 42048 4578 0 Inst_S_CPU_IF_switch_matrix.N2BEGb5
rlabel metal2 11616 5586 11616 5586 0 Inst_S_CPU_IF_switch_matrix.N2BEGb6
rlabel metal2 25056 1974 25056 1974 0 Inst_S_CPU_IF_switch_matrix.N2BEGb7
rlabel metal2 24288 5460 24288 5460 0 Inst_S_CPU_IF_switch_matrix.N4BEG0
rlabel metal2 35568 5628 35568 5628 0 Inst_S_CPU_IF_switch_matrix.N4BEG1
rlabel metal2 11904 5628 11904 5628 0 Inst_S_CPU_IF_switch_matrix.N4BEG10
rlabel metal2 19440 1932 19440 1932 0 Inst_S_CPU_IF_switch_matrix.N4BEG11
rlabel metal2 27264 9492 27264 9492 0 Inst_S_CPU_IF_switch_matrix.N4BEG12
rlabel metal2 35808 2604 35808 2604 0 Inst_S_CPU_IF_switch_matrix.N4BEG13
rlabel metal2 8256 3444 8256 3444 0 Inst_S_CPU_IF_switch_matrix.N4BEG14
rlabel metal3 30432 2310 30432 2310 0 Inst_S_CPU_IF_switch_matrix.N4BEG15
rlabel metal3 6432 4578 6432 4578 0 Inst_S_CPU_IF_switch_matrix.N4BEG2
rlabel metal2 12888 1932 12888 1932 0 Inst_S_CPU_IF_switch_matrix.N4BEG3
rlabel metal2 37200 7140 37200 7140 0 Inst_S_CPU_IF_switch_matrix.N4BEG4
rlabel metal2 43008 6552 43008 6552 0 Inst_S_CPU_IF_switch_matrix.N4BEG5
rlabel metal2 10176 5628 10176 5628 0 Inst_S_CPU_IF_switch_matrix.N4BEG6
rlabel metal2 25056 3486 25056 3486 0 Inst_S_CPU_IF_switch_matrix.N4BEG7
rlabel metal2 20400 7140 20400 7140 0 Inst_S_CPU_IF_switch_matrix.N4BEG8
rlabel metal2 33888 3486 33888 3486 0 Inst_S_CPU_IF_switch_matrix.N4BEG9
rlabel metal2 24048 5628 24048 5628 0 Inst_S_CPU_IF_switch_matrix.NN4BEG0
rlabel metal3 37728 7476 37728 7476 0 Inst_S_CPU_IF_switch_matrix.NN4BEG1
rlabel metal2 9600 6468 9600 6468 0 Inst_S_CPU_IF_switch_matrix.NN4BEG10
rlabel metal2 19392 3486 19392 3486 0 Inst_S_CPU_IF_switch_matrix.NN4BEG11
rlabel metal2 30624 9534 30624 9534 0 Inst_S_CPU_IF_switch_matrix.NN4BEG12
rlabel metal2 39288 2604 39288 2604 0 Inst_S_CPU_IF_switch_matrix.NN4BEG13
rlabel metal2 10296 4116 10296 4116 0 Inst_S_CPU_IF_switch_matrix.NN4BEG14
rlabel metal2 30048 3486 30048 3486 0 Inst_S_CPU_IF_switch_matrix.NN4BEG15
rlabel metal2 6480 5628 6480 5628 0 Inst_S_CPU_IF_switch_matrix.NN4BEG2
rlabel metal2 14016 3486 14016 3486 0 Inst_S_CPU_IF_switch_matrix.NN4BEG3
rlabel metal2 37152 8064 37152 8064 0 Inst_S_CPU_IF_switch_matrix.NN4BEG4
rlabel metal2 42240 7098 42240 7098 0 Inst_S_CPU_IF_switch_matrix.NN4BEG5
rlabel metal3 8544 8736 8544 8736 0 Inst_S_CPU_IF_switch_matrix.NN4BEG6
rlabel metal2 25440 2016 25440 2016 0 Inst_S_CPU_IF_switch_matrix.NN4BEG7
rlabel metal2 20640 7098 20640 7098 0 Inst_S_CPU_IF_switch_matrix.NN4BEG8
rlabel metal3 34752 4578 34752 4578 0 Inst_S_CPU_IF_switch_matrix.NN4BEG9
rlabel metal2 9672 6972 9672 6972 0 N1BEG[0]
rlabel metal2 9960 7140 9960 7140 0 N1BEG[1]
rlabel metal2 11448 5124 11448 5124 0 N1BEG[2]
rlabel metal2 10632 6636 10632 6636 0 N1BEG[3]
rlabel metal2 8232 9660 8232 9660 0 N2BEG[0]
rlabel metal2 9768 7980 9768 7980 0 N2BEG[1]
rlabel metal2 10632 7728 10632 7728 0 N2BEG[2]
rlabel metal2 12408 5628 12408 5628 0 N2BEG[3]
rlabel metal2 12552 6636 12552 6636 0 N2BEG[4]
rlabel metal2 12168 6972 12168 6972 0 N2BEG[5]
rlabel metal3 13152 10332 13152 10332 0 N2BEG[6]
rlabel metal3 13152 11646 13152 11646 0 N2BEG[7]
rlabel metal3 13344 10806 13344 10806 0 N2BEGb[0]
rlabel metal3 13536 9420 13536 9420 0 N2BEGb[1]
rlabel metal3 13728 10890 13728 10890 0 N2BEGb[2]
rlabel metal3 13920 10680 13920 10680 0 N2BEGb[3]
rlabel metal3 14112 9924 14112 9924 0 N2BEGb[4]
rlabel metal2 13416 6972 13416 6972 0 N2BEGb[5]
rlabel metal2 13512 7140 13512 7140 0 N2BEGb[6]
rlabel metal2 14136 6972 14136 6972 0 N2BEGb[7]
rlabel metal2 14568 7056 14568 7056 0 N4BEG[0]
rlabel metal2 16008 7056 16008 7056 0 N4BEG[10]
rlabel metal2 16488 6972 16488 6972 0 N4BEG[11]
rlabel metal2 16872 7056 16872 7056 0 N4BEG[12]
rlabel metal2 17400 6636 17400 6636 0 N4BEG[13]
rlabel metal2 14952 9660 14952 9660 0 N4BEG[14]
rlabel metal2 17784 6636 17784 6636 0 N4BEG[15]
rlabel metal3 15072 10848 15072 10848 0 N4BEG[1]
rlabel metal2 15288 6636 15288 6636 0 N4BEG[2]
rlabel metal3 15456 10722 15456 10722 0 N4BEG[3]
rlabel metal2 14184 8820 14184 8820 0 N4BEG[4]
rlabel metal3 15840 10932 15840 10932 0 N4BEG[5]
rlabel metal2 15048 7140 15048 7140 0 N4BEG[6]
rlabel metal2 13704 8904 13704 8904 0 N4BEG[7]
rlabel metal2 15432 6972 15432 6972 0 N4BEG[8]
rlabel metal2 14712 8904 14712 8904 0 N4BEG[9]
rlabel metal2 17208 8148 17208 8148 0 NN4BEG[0]
rlabel metal3 19872 10932 19872 10932 0 NN4BEG[10]
rlabel metal2 18744 8820 18744 8820 0 NN4BEG[11]
rlabel metal3 20256 8064 20256 8064 0 NN4BEG[12]
rlabel metal2 18984 8652 18984 8652 0 NN4BEG[13]
rlabel metal2 19368 9660 19368 9660 0 NN4BEG[14]
rlabel metal2 20808 7140 20808 7140 0 NN4BEG[15]
rlabel metal2 15720 9324 15720 9324 0 NN4BEG[1]
rlabel metal2 17544 7812 17544 7812 0 NN4BEG[2]
rlabel metal2 15432 9240 15432 9240 0 NN4BEG[3]
rlabel metal2 16248 8904 16248 8904 0 NN4BEG[4]
rlabel metal2 18600 6636 18600 6636 0 NN4BEG[5]
rlabel metal2 16680 9660 16680 9660 0 NN4BEG[6]
rlabel metal4 19440 10164 19440 10164 0 NN4BEG[7]
rlabel metal2 16824 9240 16824 9240 0 NN4BEG[8]
rlabel metal2 19176 6972 19176 6972 0 NN4BEG[9]
rlabel metal3 3168 996 3168 996 0 O_top0
rlabel metal3 3936 996 3936 996 0 O_top1
rlabel metal3 10848 996 10848 996 0 O_top10
rlabel metal3 11616 996 11616 996 0 O_top11
rlabel metal3 12384 954 12384 954 0 O_top12
rlabel metal3 13152 912 13152 912 0 O_top13
rlabel metal3 13920 954 13920 954 0 O_top14
rlabel metal3 14688 996 14688 996 0 O_top15
rlabel metal3 4704 996 4704 996 0 O_top2
rlabel metal3 5472 954 5472 954 0 O_top3
rlabel metal3 6240 954 6240 954 0 O_top4
rlabel metal3 7008 786 7008 786 0 O_top5
rlabel metal3 7776 1038 7776 1038 0 O_top6
rlabel metal2 8640 3444 8640 3444 0 O_top7
rlabel metal3 9312 912 9312 912 0 O_top8
rlabel metal3 10080 996 10080 996 0 O_top9
rlabel metal3 21216 11436 21216 11436 0 S1END[0]
rlabel metal3 21408 9924 21408 9924 0 S1END[1]
rlabel metal3 21600 11184 21600 11184 0 S1END[2]
rlabel metal3 21792 9840 21792 9840 0 S1END[3]
rlabel metal2 22896 9492 22896 9492 0 S2END[0]
rlabel metal3 23712 10680 23712 10680 0 S2END[1]
rlabel metal3 23904 10596 23904 10596 0 S2END[2]
rlabel metal3 24096 10680 24096 10680 0 S2END[3]
rlabel metal3 24288 10638 24288 10638 0 S2END[4]
rlabel metal3 24480 11226 24480 11226 0 S2END[5]
rlabel metal3 24672 10932 24672 10932 0 S2END[6]
rlabel metal3 24864 10680 24864 10680 0 S2END[7]
rlabel metal3 21984 9546 21984 9546 0 S2MID[0]
rlabel metal3 22176 9924 22176 9924 0 S2MID[1]
rlabel metal3 22368 10848 22368 10848 0 S2MID[2]
rlabel metal3 22560 10722 22560 10722 0 S2MID[3]
rlabel metal3 22752 10932 22752 10932 0 S2MID[4]
rlabel metal3 22944 10596 22944 10596 0 S2MID[5]
rlabel metal2 22704 9828 22704 9828 0 S2MID[6]
rlabel metal2 22944 9660 22944 9660 0 S2MID[7]
rlabel metal3 25056 9462 25056 9462 0 S4END[0]
rlabel metal3 26976 9462 26976 9462 0 S4END[10]
rlabel metal3 27168 10932 27168 10932 0 S4END[11]
rlabel metal3 27360 10596 27360 10596 0 S4END[12]
rlabel metal3 27552 10680 27552 10680 0 S4END[13]
rlabel metal3 27744 11226 27744 11226 0 S4END[14]
rlabel metal3 27936 9126 27936 9126 0 S4END[15]
rlabel metal3 25248 11310 25248 11310 0 S4END[1]
rlabel metal3 25440 9420 25440 9420 0 S4END[2]
rlabel metal3 25632 11184 25632 11184 0 S4END[3]
rlabel metal3 25824 11058 25824 11058 0 S4END[4]
rlabel metal3 26016 11352 26016 11352 0 S4END[5]
rlabel metal3 26208 10386 26208 10386 0 S4END[6]
rlabel metal3 26400 11478 26400 11478 0 S4END[7]
rlabel metal3 26592 10218 26592 10218 0 S4END[8]
rlabel metal3 26784 11562 26784 11562 0 S4END[9]
rlabel metal3 28128 10932 28128 10932 0 SS4END[0]
rlabel metal3 30048 11688 30048 11688 0 SS4END[10]
rlabel metal4 31056 9996 31056 9996 0 SS4END[11]
rlabel metal3 36000 10122 36000 10122 0 SS4END[12]
rlabel metal3 34944 9450 34944 9450 0 SS4END[13]
rlabel metal2 33888 8022 33888 8022 0 SS4END[14]
rlabel metal3 31008 10932 31008 10932 0 SS4END[15]
rlabel metal3 28320 11394 28320 11394 0 SS4END[1]
rlabel metal2 30288 7980 30288 7980 0 SS4END[2]
rlabel metal3 28704 11268 28704 11268 0 SS4END[3]
rlabel metal3 28896 11436 28896 11436 0 SS4END[4]
rlabel metal3 29088 10932 29088 10932 0 SS4END[5]
rlabel metal3 29280 10218 29280 10218 0 SS4END[6]
rlabel metal3 29472 11562 29472 11562 0 SS4END[7]
rlabel metal3 34560 10122 34560 10122 0 SS4END[8]
rlabel metal3 29856 11646 29856 11646 0 SS4END[9]
rlabel metal3 38880 1302 38880 1302 0 UserCLK
rlabel metal2 32088 5544 32088 5544 0 UserCLKo
rlabel metal2 1896 2100 1896 2100 0 net1
rlabel metal3 3552 7938 3552 7938 0 net10
rlabel metal2 29280 2688 29280 2688 0 net100
rlabel metal2 41472 6426 41472 6426 0 net101
rlabel metal3 33600 8232 33600 8232 0 net102
rlabel metal3 16224 3402 16224 3402 0 net103
rlabel metal3 35712 7602 35712 7602 0 net104
rlabel via1 35604 7896 35604 7896 0 net105
rlabel metal2 23568 6384 23568 6384 0 net106
rlabel metal2 9936 4200 9936 4200 0 net107
rlabel metal2 39168 3318 39168 3318 0 net108
rlabel metal2 31272 9660 31272 9660 0 net109
rlabel metal2 1728 6930 1728 6930 0 net11
rlabel metal3 21504 5838 21504 5838 0 net110
rlabel metal3 13920 5880 13920 5880 0 net111
rlabel metal2 33360 4872 33360 4872 0 net112
rlabel metal3 20352 8652 20352 8652 0 net113
rlabel metal2 34056 9576 34056 9576 0 net114
rlabel metal2 10128 8736 10128 8736 0 net115
rlabel metal3 35040 3276 35040 3276 0 net116
rlabel metal5 13536 5376 13536 5376 0 net117
rlabel metal2 33792 3402 33792 3402 0 net118
rlabel metal2 44544 5040 44544 5040 0 net119
rlabel metal2 2784 1512 2784 1512 0 net12
rlabel metal2 41280 4704 41280 4704 0 net120
rlabel metal2 41040 3360 41040 3360 0 net121
rlabel metal2 24120 4368 24120 4368 0 net122
rlabel metal3 35424 3486 35424 3486 0 net123
rlabel metal2 44064 6300 44064 6300 0 net124
rlabel metal2 4056 6972 4056 6972 0 net125
rlabel metal2 12168 4704 12168 4704 0 net126
rlabel metal2 43008 1974 43008 1974 0 net127
rlabel metal3 41280 8358 41280 8358 0 net128
rlabel metal2 41184 4956 41184 4956 0 net129
rlabel metal3 1728 7686 1728 7686 0 net13
rlabel metal3 15168 4956 15168 4956 0 net130
rlabel metal2 27864 6216 27864 6216 0 net131
rlabel metal3 14784 6804 14784 6804 0 net132
rlabel metal2 35400 3948 35400 3948 0 net133
rlabel metal3 40224 8778 40224 8778 0 net134
rlabel metal2 40464 8652 40464 8652 0 net135
rlabel metal2 33864 7392 33864 7392 0 net136
rlabel metal3 41328 2268 41328 2268 0 net137
rlabel metal2 40176 2856 40176 2856 0 net138
rlabel metal2 15432 5544 15432 5544 0 net139
rlabel metal3 39456 7434 39456 7434 0 net14
rlabel metal2 25608 5544 25608 5544 0 net140
rlabel metal2 38880 1428 38880 1428 0 net141
rlabel metal3 39648 3528 39648 3528 0 net142
rlabel metal2 41856 1848 41856 1848 0 net143
rlabel metal2 40128 1932 40128 1932 0 net144
rlabel metal3 33600 2058 33600 2058 0 net145
rlabel metal2 33216 1470 33216 1470 0 net146
rlabel metal2 22464 3990 22464 3990 0 net147
rlabel metal2 38424 8148 38424 8148 0 net148
rlabel metal2 37416 2100 37416 2100 0 net149
rlabel metal2 1488 8946 1488 8946 0 net15
rlabel metal3 42240 6804 42240 6804 0 net150
rlabel metal2 38568 2100 38568 2100 0 net151
rlabel metal3 41232 4956 41232 4956 0 net152
rlabel metal3 39072 9660 39072 9660 0 net153
rlabel metal3 36960 8148 36960 8148 0 net154
rlabel metal3 42048 7980 42048 7980 0 net155
rlabel metal3 39072 9072 39072 9072 0 net156
rlabel metal2 40440 9492 40440 9492 0 net157
rlabel metal2 39168 5376 39168 5376 0 net158
rlabel metal4 33312 7098 33312 7098 0 net159
rlabel metal3 27168 6888 27168 6888 0 net16
rlabel metal2 39768 8652 39768 8652 0 net160
rlabel metal2 41688 2856 41688 2856 0 net161
rlabel metal2 42120 2604 42120 2604 0 net162
rlabel metal2 41304 2856 41304 2856 0 net163
rlabel metal2 38928 7392 38928 7392 0 net164
rlabel metal2 35688 2100 35688 2100 0 net165
rlabel metal2 41448 2100 41448 2100 0 net166
rlabel metal2 40488 2100 40488 2100 0 net167
rlabel metal3 22656 2058 22656 2058 0 net168
rlabel metal2 15744 2856 15744 2856 0 net169
rlabel metal2 2280 8652 2280 8652 0 net17
rlabel metal2 34176 1722 34176 1722 0 net170
rlabel metal2 25584 1512 25584 1512 0 net171
rlabel metal3 16896 3066 16896 3066 0 net172
rlabel metal3 7488 4872 7488 4872 0 net173
rlabel metal2 34080 6888 34080 6888 0 net174
rlabel metal2 26640 2016 26640 2016 0 net175
rlabel metal3 16320 2562 16320 2562 0 net176
rlabel metal2 18912 3528 18912 3528 0 net177
rlabel metal2 18672 2604 18672 2604 0 net178
rlabel metal2 18384 1932 18384 1932 0 net179
rlabel metal2 1608 9240 1608 9240 0 net18
rlabel metal2 19200 1848 19200 1848 0 net180
rlabel metal3 20640 8988 20640 8988 0 net181
rlabel metal2 21696 2814 21696 2814 0 net182
rlabel metal2 22176 1932 22176 1932 0 net183
rlabel metal2 22368 8064 22368 8064 0 net184
rlabel metal2 36024 5460 36024 5460 0 net185
rlabel metal2 11496 4284 11496 4284 0 net186
rlabel metal2 16536 2100 16536 2100 0 net187
rlabel metal3 21600 6930 21600 6930 0 net188
rlabel metal2 33816 4788 33816 4788 0 net189
rlabel metal2 1872 9156 1872 9156 0 net19
rlabel metal2 6888 7140 6888 7140 0 net190
rlabel metal2 14616 3612 14616 3612 0 net191
rlabel metal3 12288 6510 12288 6510 0 net192
rlabel metal2 39672 4116 39672 4116 0 net193
rlabel metal2 9288 4284 9288 4284 0 net194
rlabel metal2 14400 5040 14400 5040 0 net195
rlabel metal2 9696 9450 9696 9450 0 net196
rlabel metal2 36840 5628 36840 5628 0 net197
rlabel metal2 8520 6972 8520 6972 0 net198
rlabel metal2 13944 2100 13944 2100 0 net199
rlabel metal2 1536 4158 1536 4158 0 net2
rlabel metal2 2496 9198 2496 9198 0 net20
rlabel metal3 38784 8316 38784 8316 0 net200
rlabel metal2 41784 3948 41784 3948 0 net201
rlabel metal2 12456 5796 12456 5796 0 net202
rlabel metal4 17952 1848 17952 1848 0 net203
rlabel metal2 20448 6258 20448 6258 0 net204
rlabel metal3 15552 6216 15552 6216 0 net205
rlabel metal2 19464 1680 19464 1680 0 net206
rlabel metal3 16224 8064 16224 8064 0 net207
rlabel metal2 35640 2772 35640 2772 0 net208
rlabel metal3 13536 4914 13536 4914 0 net209
rlabel metal2 2760 9240 2760 9240 0 net21
rlabel metal3 18048 6300 18048 6300 0 net210
rlabel metal3 35040 5670 35040 5670 0 net211
rlabel metal3 14400 5166 14400 5166 0 net212
rlabel metal2 12648 1932 12648 1932 0 net213
rlabel metal3 36864 6846 36864 6846 0 net214
rlabel metal2 42360 6216 42360 6216 0 net215
rlabel metal3 14496 5166 14496 5166 0 net216
rlabel metal2 24792 3444 24792 3444 0 net217
rlabel metal2 15216 7140 15216 7140 0 net218
rlabel metal2 33672 3276 33672 3276 0 net219
rlabel metal2 36912 2688 36912 2688 0 net22
rlabel metal2 22464 5376 22464 5376 0 net220
rlabel metal2 9984 6174 9984 6174 0 net221
rlabel metal2 19272 3276 19272 3276 0 net222
rlabel metal3 19680 6636 19680 6636 0 net223
rlabel metal3 38976 2520 38976 2520 0 net224
rlabel metal3 13248 3906 13248 3906 0 net225
rlabel metal2 29688 3444 29688 3444 0 net226
rlabel metal4 20208 5964 20208 5964 0 net227
rlabel metal3 13344 4536 13344 4536 0 net228
rlabel metal2 14280 3528 14280 3528 0 net229
rlabel metal2 3096 2100 3096 2100 0 net23
rlabel metal3 15936 8232 15936 8232 0 net230
rlabel metal3 41952 6468 41952 6468 0 net231
rlabel metal3 15456 9240 15456 9240 0 net232
rlabel metal2 25224 2016 25224 2016 0 net233
rlabel metal2 20424 6972 20424 6972 0 net234
rlabel metal3 23136 4242 23136 4242 0 net235
rlabel metal2 42456 2856 42456 2856 0 net236
rlabel metal3 21024 11352 21024 11352 0 net237
rlabel metal2 5352 8904 5352 8904 0 net24
rlabel metal3 17664 8694 17664 8694 0 net25
rlabel metal2 6528 1848 6528 1848 0 net26
rlabel metal2 36768 4116 36768 4116 0 net27
rlabel metal2 1992 2436 1992 2436 0 net28
rlabel metal2 13920 9366 13920 9366 0 net29
rlabel metal2 17328 4872 17328 4872 0 net3
rlabel metal3 22656 4368 22656 4368 0 net30
rlabel metal2 1728 3360 1728 3360 0 net31
rlabel metal2 21504 1848 21504 1848 0 net32
rlabel metal2 16320 2688 16320 2688 0 net33
rlabel metal2 4872 2100 4872 2100 0 net34
rlabel metal2 41040 4788 41040 4788 0 net35
rlabel metal3 33696 2322 33696 2322 0 net36
rlabel metal2 14544 1764 14544 1764 0 net37
rlabel metal2 11112 2016 11112 2016 0 net38
rlabel metal2 15672 2016 15672 2016 0 net39
rlabel metal3 22752 6468 22752 6468 0 net4
rlabel metal2 15240 1932 15240 1932 0 net40
rlabel metal3 34272 2100 34272 2100 0 net41
rlabel metal3 13248 2730 13248 2730 0 net42
rlabel metal2 5880 1680 5880 1680 0 net43
rlabel metal2 17284 1848 17284 1848 0 net44
rlabel metal2 21312 5754 21312 5754 0 net45
rlabel metal2 38592 4788 38592 4788 0 net46
rlabel metal3 22272 4872 22272 4872 0 net47
rlabel metal2 18336 4830 18336 4830 0 net48
rlabel metal2 15264 2646 15264 2646 0 net49
rlabel metal3 31872 2142 31872 2142 0 net5
rlabel metal2 14712 4788 14712 4788 0 net50
rlabel metal2 36192 8694 36192 8694 0 net51
rlabel metal2 22200 5628 22200 5628 0 net52
rlabel metal2 22424 4872 22424 4872 0 net53
rlabel metal3 22944 2730 22944 2730 0 net54
rlabel metal2 20736 1848 20736 1848 0 net55
rlabel metal2 25944 6972 25944 6972 0 net56
rlabel metal2 7584 9450 7584 9450 0 net57
rlabel metal2 19872 4956 19872 4956 0 net58
rlabel metal2 5976 2100 5976 2100 0 net59
rlabel metal2 6336 2688 6336 2688 0 net6
rlabel metal4 13920 1512 13920 1512 0 net60
rlabel metal4 21312 9408 21312 9408 0 net61
rlabel metal3 22944 3192 22944 3192 0 net62
rlabel metal2 9768 2100 9768 2100 0 net63
rlabel metal2 15936 2688 15936 2688 0 net64
rlabel metal2 9408 4914 9408 4914 0 net65
rlabel metal2 20880 9156 20880 9156 0 net66
rlabel metal3 24672 8232 24672 8232 0 net67
rlabel metal4 20976 2268 20976 2268 0 net68
rlabel metal3 22656 7980 22656 7980 0 net69
rlabel metal3 18432 1932 18432 1932 0 net7
rlabel metal3 33312 4284 33312 4284 0 net70
rlabel metal2 19392 8778 19392 8778 0 net71
rlabel metal2 21696 1680 21696 1680 0 net72
rlabel metal2 8736 9366 8736 9366 0 net73
rlabel metal2 26088 9240 26088 9240 0 net74
rlabel metal2 26376 9240 26376 9240 0 net75
rlabel metal3 28800 4368 28800 4368 0 net76
rlabel metal2 8997 5712 8997 5712 0 net77
rlabel metal3 22464 7560 22464 7560 0 net78
rlabel metal3 22464 9156 22464 9156 0 net79
rlabel metal2 21120 2688 21120 2688 0 net8
rlabel metal3 15648 3528 15648 3528 0 net80
rlabel metal2 21336 9492 21336 9492 0 net81
rlabel metal2 33888 6384 33888 6384 0 net82
rlabel metal3 21600 8190 21600 8190 0 net83
rlabel via2 28704 2604 28704 2604 0 net84
rlabel metal3 39648 6090 39648 6090 0 net85
rlabel metal2 35232 9366 35232 9366 0 net86
rlabel metal2 14688 2520 14688 2520 0 net87
rlabel metal2 6384 6384 6384 6384 0 net88
rlabel metal2 34896 7140 34896 7140 0 net89
rlabel metal2 1536 6048 1536 6048 0 net9
rlabel metal2 23952 5712 23952 5712 0 net90
rlabel metal3 7680 6636 7680 6636 0 net91
rlabel metal2 35172 2688 35172 2688 0 net92
rlabel metal2 24816 9408 24816 9408 0 net93
rlabel metal2 23040 2394 23040 2394 0 net94
rlabel metal3 28800 8778 28800 8778 0 net95
rlabel metal2 33312 4116 33312 4116 0 net96
rlabel metal2 22224 10164 22224 10164 0 net97
rlabel metal2 24384 3360 24384 3360 0 net98
rlabel metal2 10560 9408 10560 9408 0 net99
<< properties >>
string FIXED_BBOX 0 0 46368 11844
<< end >>
