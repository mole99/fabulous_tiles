magic
tech ihp-sg13g2
magscale 1 2
timestamp 1743691081
<< metal1 >>
rect 1152 95276 20452 95300
rect 1152 95236 4928 95276
rect 4968 95236 5010 95276
rect 5050 95236 5092 95276
rect 5132 95236 5174 95276
rect 5214 95236 5256 95276
rect 5296 95236 20048 95276
rect 20088 95236 20130 95276
rect 20170 95236 20212 95276
rect 20252 95236 20294 95276
rect 20334 95236 20376 95276
rect 20416 95236 20452 95276
rect 1152 95212 20452 95236
rect 7323 95108 7365 95117
rect 7323 95068 7324 95108
rect 7364 95068 7365 95108
rect 7323 95059 7365 95068
rect 1563 95024 1605 95033
rect 1563 94984 1564 95024
rect 1604 94984 1605 95024
rect 1563 94975 1605 94984
rect 2715 95024 2757 95033
rect 2715 94984 2716 95024
rect 2756 94984 2757 95024
rect 2715 94975 2757 94984
rect 3483 95024 3525 95033
rect 3483 94984 3484 95024
rect 3524 94984 3525 95024
rect 3483 94975 3525 94984
rect 4635 95024 4677 95033
rect 4635 94984 4636 95024
rect 4676 94984 4677 95024
rect 4635 94975 4677 94984
rect 5019 95024 5061 95033
rect 5019 94984 5020 95024
rect 5060 94984 5061 95024
rect 5019 94975 5061 94984
rect 5787 95024 5829 95033
rect 5787 94984 5788 95024
rect 5828 94984 5829 95024
rect 5787 94975 5829 94984
rect 6939 95024 6981 95033
rect 6939 94984 6940 95024
rect 6980 94984 6981 95024
rect 6939 94975 6981 94984
rect 8091 95024 8133 95033
rect 8091 94984 8092 95024
rect 8132 94984 8133 95024
rect 8091 94975 8133 94984
rect 15675 95024 15717 95033
rect 15675 94984 15676 95024
rect 15716 94984 15717 95024
rect 15675 94975 15717 94984
rect 16059 95024 16101 95033
rect 16059 94984 16060 95024
rect 16100 94984 16101 95024
rect 16059 94975 16101 94984
rect 16827 95024 16869 95033
rect 16827 94984 16828 95024
rect 16868 94984 16869 95024
rect 16827 94975 16869 94984
rect 17211 95024 17253 95033
rect 17211 94984 17212 95024
rect 17252 94984 17253 95024
rect 17211 94975 17253 94984
rect 18363 95024 18405 95033
rect 18363 94984 18364 95024
rect 18404 94984 18405 95024
rect 18363 94975 18405 94984
rect 18747 95024 18789 95033
rect 18747 94984 18748 95024
rect 18788 94984 18789 95024
rect 18747 94975 18789 94984
rect 19899 95024 19941 95033
rect 19899 94984 19900 95024
rect 19940 94984 19941 95024
rect 19899 94975 19941 94984
rect 1323 94856 1365 94865
rect 1323 94816 1324 94856
rect 1364 94816 1365 94856
rect 1323 94807 1365 94816
rect 1707 94856 1749 94865
rect 1707 94816 1708 94856
rect 1748 94816 1749 94856
rect 1707 94807 1749 94816
rect 2091 94856 2133 94865
rect 2091 94816 2092 94856
rect 2132 94816 2133 94856
rect 2091 94807 2133 94816
rect 2475 94856 2517 94865
rect 2475 94816 2476 94856
rect 2516 94816 2517 94856
rect 2475 94807 2517 94816
rect 2859 94856 2901 94865
rect 2859 94816 2860 94856
rect 2900 94816 2901 94856
rect 2859 94807 2901 94816
rect 3243 94856 3285 94865
rect 3243 94816 3244 94856
rect 3284 94816 3285 94856
rect 3243 94807 3285 94816
rect 3627 94856 3669 94865
rect 3627 94816 3628 94856
rect 3668 94816 3669 94856
rect 3627 94807 3669 94816
rect 4011 94856 4053 94865
rect 4011 94816 4012 94856
rect 4052 94816 4053 94856
rect 4011 94807 4053 94816
rect 4395 94856 4437 94865
rect 4395 94816 4396 94856
rect 4436 94816 4437 94856
rect 4395 94807 4437 94816
rect 4779 94856 4821 94865
rect 4779 94816 4780 94856
rect 4820 94816 4821 94856
rect 4779 94807 4821 94816
rect 5163 94856 5205 94865
rect 5163 94816 5164 94856
rect 5204 94816 5205 94856
rect 5163 94807 5205 94816
rect 5547 94856 5589 94865
rect 5547 94816 5548 94856
rect 5588 94816 5589 94856
rect 5547 94807 5589 94816
rect 5931 94856 5973 94865
rect 5931 94816 5932 94856
rect 5972 94816 5973 94856
rect 5931 94807 5973 94816
rect 6315 94856 6357 94865
rect 6315 94816 6316 94856
rect 6356 94816 6357 94856
rect 6315 94807 6357 94816
rect 6699 94856 6741 94865
rect 6699 94816 6700 94856
rect 6740 94816 6741 94856
rect 6699 94807 6741 94816
rect 7083 94856 7125 94865
rect 7083 94816 7084 94856
rect 7124 94816 7125 94856
rect 7083 94807 7125 94816
rect 7467 94856 7509 94865
rect 7467 94816 7468 94856
rect 7508 94816 7509 94856
rect 7467 94807 7509 94816
rect 7851 94856 7893 94865
rect 7851 94816 7852 94856
rect 7892 94816 7893 94856
rect 7851 94807 7893 94816
rect 8235 94856 8277 94865
rect 8235 94816 8236 94856
rect 8276 94816 8277 94856
rect 8235 94807 8277 94816
rect 8619 94856 8661 94865
rect 8619 94816 8620 94856
rect 8660 94816 8661 94856
rect 8619 94807 8661 94816
rect 9195 94856 9237 94865
rect 9195 94816 9196 94856
rect 9236 94816 9237 94856
rect 9195 94807 9237 94816
rect 9579 94856 9621 94865
rect 9579 94816 9580 94856
rect 9620 94816 9621 94856
rect 9579 94807 9621 94816
rect 9963 94856 10005 94865
rect 9963 94816 9964 94856
rect 10004 94816 10005 94856
rect 9963 94807 10005 94816
rect 10155 94856 10197 94865
rect 10155 94816 10156 94856
rect 10196 94816 10197 94856
rect 10155 94807 10197 94816
rect 10731 94856 10773 94865
rect 10731 94816 10732 94856
rect 10772 94816 10773 94856
rect 10731 94807 10773 94816
rect 10923 94856 10965 94865
rect 10923 94816 10924 94856
rect 10964 94816 10965 94856
rect 10923 94807 10965 94816
rect 11307 94856 11349 94865
rect 11307 94816 11308 94856
rect 11348 94816 11349 94856
rect 11307 94807 11349 94816
rect 11883 94856 11925 94865
rect 11883 94816 11884 94856
rect 11924 94816 11925 94856
rect 11883 94807 11925 94816
rect 12075 94856 12117 94865
rect 12075 94816 12076 94856
rect 12116 94816 12117 94856
rect 12075 94807 12117 94816
rect 12651 94856 12693 94865
rect 12651 94816 12652 94856
rect 12692 94816 12693 94856
rect 12651 94807 12693 94816
rect 12843 94856 12885 94865
rect 12843 94816 12844 94856
rect 12884 94816 12885 94856
rect 12843 94807 12885 94816
rect 13419 94856 13461 94865
rect 13419 94816 13420 94856
rect 13460 94816 13461 94856
rect 13419 94807 13461 94816
rect 13611 94856 13653 94865
rect 13611 94816 13612 94856
rect 13652 94816 13653 94856
rect 13611 94807 13653 94816
rect 14187 94856 14229 94865
rect 14187 94816 14188 94856
rect 14228 94816 14229 94856
rect 14187 94807 14229 94816
rect 14379 94856 14421 94865
rect 14379 94816 14380 94856
rect 14420 94816 14421 94856
rect 14379 94807 14421 94816
rect 14955 94856 14997 94865
rect 14955 94816 14956 94856
rect 14996 94816 14997 94856
rect 14955 94807 14997 94816
rect 15915 94856 15957 94865
rect 15915 94816 15916 94856
rect 15956 94816 15957 94856
rect 15915 94807 15957 94816
rect 16347 94856 16389 94865
rect 16347 94816 16348 94856
rect 16388 94816 16389 94856
rect 16347 94807 16389 94816
rect 16683 94856 16725 94865
rect 16683 94816 16684 94856
rect 16724 94816 16725 94856
rect 16683 94807 16725 94816
rect 17067 94856 17109 94865
rect 17067 94816 17068 94856
rect 17108 94816 17109 94856
rect 17067 94807 17109 94816
rect 17451 94856 17493 94865
rect 17451 94816 17452 94856
rect 17492 94816 17493 94856
rect 17451 94807 17493 94816
rect 17835 94856 17877 94865
rect 17835 94816 17836 94856
rect 17876 94816 17877 94856
rect 17835 94807 17877 94816
rect 18219 94856 18261 94865
rect 18219 94816 18220 94856
rect 18260 94816 18261 94856
rect 18219 94807 18261 94816
rect 18603 94856 18645 94865
rect 18603 94816 18604 94856
rect 18644 94816 18645 94856
rect 18603 94807 18645 94816
rect 18987 94856 19029 94865
rect 18987 94816 18988 94856
rect 19028 94816 19029 94856
rect 18987 94807 19029 94816
rect 19371 94856 19413 94865
rect 19371 94816 19372 94856
rect 19412 94816 19413 94856
rect 19371 94807 19413 94816
rect 19755 94856 19797 94865
rect 19755 94816 19756 94856
rect 19796 94816 19797 94856
rect 19755 94807 19797 94816
rect 20139 94856 20181 94865
rect 20139 94816 20140 94856
rect 20180 94816 20181 94856
rect 20139 94807 20181 94816
rect 1947 94772 1989 94781
rect 1947 94732 1948 94772
rect 1988 94732 1989 94772
rect 1947 94723 1989 94732
rect 3099 94772 3141 94781
rect 3099 94732 3100 94772
rect 3140 94732 3141 94772
rect 3099 94723 3141 94732
rect 3867 94772 3909 94781
rect 3867 94732 3868 94772
rect 3908 94732 3909 94772
rect 3867 94723 3909 94732
rect 5403 94772 5445 94781
rect 5403 94732 5404 94772
rect 5444 94732 5445 94772
rect 5403 94723 5445 94732
rect 6171 94772 6213 94781
rect 6171 94732 6172 94772
rect 6212 94732 6213 94772
rect 6171 94723 6213 94732
rect 7707 94772 7749 94781
rect 7707 94732 7708 94772
rect 7748 94732 7749 94772
rect 7707 94723 7749 94732
rect 8859 94772 8901 94781
rect 8859 94732 8860 94772
rect 8900 94732 8901 94772
rect 8859 94723 8901 94732
rect 10395 94772 10437 94781
rect 10395 94732 10396 94772
rect 10436 94732 10437 94772
rect 10395 94723 10437 94732
rect 11547 94772 11589 94781
rect 11547 94732 11548 94772
rect 11588 94732 11589 94772
rect 11547 94723 11589 94732
rect 12315 94772 12357 94781
rect 12315 94732 12316 94772
rect 12356 94732 12357 94772
rect 12315 94723 12357 94732
rect 13083 94772 13125 94781
rect 13083 94732 13084 94772
rect 13124 94732 13125 94772
rect 13083 94723 13125 94732
rect 13851 94772 13893 94781
rect 13851 94732 13852 94772
rect 13892 94732 13893 94772
rect 13851 94723 13893 94732
rect 14619 94772 14661 94781
rect 14619 94732 14620 94772
rect 14660 94732 14661 94772
rect 14619 94723 14661 94732
rect 2331 94688 2373 94697
rect 2331 94648 2332 94688
rect 2372 94648 2373 94688
rect 2331 94639 2373 94648
rect 4251 94688 4293 94697
rect 4251 94648 4252 94688
rect 4292 94648 4293 94688
rect 4251 94639 4293 94648
rect 6555 94688 6597 94697
rect 6555 94648 6556 94688
rect 6596 94648 6597 94688
rect 6555 94639 6597 94648
rect 8475 94688 8517 94697
rect 8475 94648 8476 94688
rect 8516 94648 8517 94688
rect 8475 94639 8517 94648
rect 8955 94688 8997 94697
rect 8955 94648 8956 94688
rect 8996 94648 8997 94688
rect 8955 94639 8997 94648
rect 9339 94688 9381 94697
rect 9339 94648 9340 94688
rect 9380 94648 9381 94688
rect 9339 94639 9381 94648
rect 9723 94688 9765 94697
rect 9723 94648 9724 94688
rect 9764 94648 9765 94688
rect 9723 94639 9765 94648
rect 10491 94688 10533 94697
rect 10491 94648 10492 94688
rect 10532 94648 10533 94688
rect 10491 94639 10533 94648
rect 11163 94688 11205 94697
rect 11163 94648 11164 94688
rect 11204 94648 11205 94688
rect 11163 94639 11205 94648
rect 11643 94688 11685 94697
rect 11643 94648 11644 94688
rect 11684 94648 11685 94688
rect 11643 94639 11685 94648
rect 12411 94688 12453 94697
rect 12411 94648 12412 94688
rect 12452 94648 12453 94688
rect 12411 94639 12453 94648
rect 13179 94688 13221 94697
rect 13179 94648 13180 94688
rect 13220 94648 13221 94688
rect 13179 94639 13221 94648
rect 13947 94688 13989 94697
rect 13947 94648 13948 94688
rect 13988 94648 13989 94688
rect 13947 94639 13989 94648
rect 14715 94688 14757 94697
rect 14715 94648 14716 94688
rect 14756 94648 14757 94688
rect 14715 94639 14757 94648
rect 16443 94688 16485 94697
rect 16443 94648 16444 94688
rect 16484 94648 16485 94688
rect 16443 94639 16485 94648
rect 17595 94688 17637 94697
rect 17595 94648 17596 94688
rect 17636 94648 17637 94688
rect 17595 94639 17637 94648
rect 17979 94688 18021 94697
rect 17979 94648 17980 94688
rect 18020 94648 18021 94688
rect 17979 94639 18021 94648
rect 19131 94688 19173 94697
rect 19131 94648 19132 94688
rect 19172 94648 19173 94688
rect 19131 94639 19173 94648
rect 19515 94688 19557 94697
rect 19515 94648 19516 94688
rect 19556 94648 19557 94688
rect 19515 94639 19557 94648
rect 1152 94520 20448 94544
rect 1152 94480 3688 94520
rect 3728 94480 3770 94520
rect 3810 94480 3852 94520
rect 3892 94480 3934 94520
rect 3974 94480 4016 94520
rect 4056 94480 18808 94520
rect 18848 94480 18890 94520
rect 18930 94480 18972 94520
rect 19012 94480 19054 94520
rect 19094 94480 19136 94520
rect 19176 94480 20448 94520
rect 1152 94456 20448 94480
rect 2235 94352 2277 94361
rect 2235 94312 2236 94352
rect 2276 94312 2277 94352
rect 2235 94303 2277 94312
rect 2619 94352 2661 94361
rect 2619 94312 2620 94352
rect 2660 94312 2661 94352
rect 2619 94303 2661 94312
rect 3003 94352 3045 94361
rect 3003 94312 3004 94352
rect 3044 94312 3045 94352
rect 3003 94303 3045 94312
rect 3579 94352 3621 94361
rect 3579 94312 3580 94352
rect 3620 94312 3621 94352
rect 3579 94303 3621 94312
rect 3963 94352 4005 94361
rect 3963 94312 3964 94352
rect 4004 94312 4005 94352
rect 3963 94303 4005 94312
rect 4347 94352 4389 94361
rect 4347 94312 4348 94352
rect 4388 94312 4389 94352
rect 4347 94303 4389 94312
rect 4731 94352 4773 94361
rect 4731 94312 4732 94352
rect 4772 94312 4773 94352
rect 4731 94303 4773 94312
rect 5115 94352 5157 94361
rect 5115 94312 5116 94352
rect 5156 94312 5157 94352
rect 5115 94303 5157 94312
rect 5883 94352 5925 94361
rect 5883 94312 5884 94352
rect 5924 94312 5925 94352
rect 5883 94303 5925 94312
rect 6267 94352 6309 94361
rect 6267 94312 6268 94352
rect 6308 94312 6309 94352
rect 6267 94303 6309 94312
rect 6651 94352 6693 94361
rect 6651 94312 6652 94352
rect 6692 94312 6693 94352
rect 6651 94303 6693 94312
rect 7035 94352 7077 94361
rect 7035 94312 7036 94352
rect 7076 94312 7077 94352
rect 7035 94303 7077 94312
rect 7419 94352 7461 94361
rect 7419 94312 7420 94352
rect 7460 94312 7461 94352
rect 7419 94303 7461 94312
rect 7803 94352 7845 94361
rect 7803 94312 7804 94352
rect 7844 94312 7845 94352
rect 7803 94303 7845 94312
rect 8571 94352 8613 94361
rect 8571 94312 8572 94352
rect 8612 94312 8613 94352
rect 8571 94303 8613 94312
rect 16443 94352 16485 94361
rect 16443 94312 16444 94352
rect 16484 94312 16485 94352
rect 16443 94303 16485 94312
rect 1851 94268 1893 94277
rect 1851 94228 1852 94268
rect 1892 94228 1893 94268
rect 1851 94219 1893 94228
rect 3387 94268 3429 94277
rect 3387 94228 3388 94268
rect 3428 94228 3429 94268
rect 3387 94219 3429 94228
rect 5499 94268 5541 94277
rect 5499 94228 5500 94268
rect 5540 94228 5541 94268
rect 5499 94219 5541 94228
rect 8187 94268 8229 94277
rect 8187 94228 8188 94268
rect 8228 94228 8229 94268
rect 8187 94219 8229 94228
rect 17211 94268 17253 94277
rect 17211 94228 17212 94268
rect 17252 94228 17253 94268
rect 17211 94219 17253 94228
rect 1227 94184 1269 94193
rect 1227 94144 1228 94184
rect 1268 94144 1269 94184
rect 1227 94135 1269 94144
rect 1611 94184 1653 94193
rect 1611 94144 1612 94184
rect 1652 94144 1653 94184
rect 1611 94135 1653 94144
rect 1995 94184 2037 94193
rect 1995 94144 1996 94184
rect 2036 94144 2037 94184
rect 1995 94135 2037 94144
rect 2379 94184 2421 94193
rect 2379 94144 2380 94184
rect 2420 94144 2421 94184
rect 2379 94135 2421 94144
rect 2763 94184 2805 94193
rect 2763 94144 2764 94184
rect 2804 94144 2805 94184
rect 2763 94135 2805 94144
rect 3147 94184 3189 94193
rect 3147 94144 3148 94184
rect 3188 94144 3189 94184
rect 3147 94135 3189 94144
rect 3819 94184 3861 94193
rect 3819 94144 3820 94184
rect 3860 94144 3861 94184
rect 3819 94135 3861 94144
rect 4203 94184 4245 94193
rect 4203 94144 4204 94184
rect 4244 94144 4245 94184
rect 4203 94135 4245 94144
rect 4587 94184 4629 94193
rect 4587 94144 4588 94184
rect 4628 94144 4629 94184
rect 4587 94135 4629 94144
rect 4971 94184 5013 94193
rect 4971 94144 4972 94184
rect 5012 94144 5013 94184
rect 4971 94135 5013 94144
rect 5355 94184 5397 94193
rect 5355 94144 5356 94184
rect 5396 94144 5397 94184
rect 5355 94135 5397 94144
rect 5739 94184 5781 94193
rect 5739 94144 5740 94184
rect 5780 94144 5781 94184
rect 5739 94135 5781 94144
rect 6123 94184 6165 94193
rect 6123 94144 6124 94184
rect 6164 94144 6165 94184
rect 6123 94135 6165 94144
rect 6507 94184 6549 94193
rect 6507 94144 6508 94184
rect 6548 94144 6549 94184
rect 6507 94135 6549 94144
rect 6891 94184 6933 94193
rect 6891 94144 6892 94184
rect 6932 94144 6933 94184
rect 6891 94135 6933 94144
rect 7275 94184 7317 94193
rect 7275 94144 7276 94184
rect 7316 94144 7317 94184
rect 7275 94135 7317 94144
rect 7659 94184 7701 94193
rect 7659 94144 7660 94184
rect 7700 94144 7701 94184
rect 7659 94135 7701 94144
rect 8043 94184 8085 94193
rect 8043 94144 8044 94184
rect 8084 94144 8085 94184
rect 8043 94135 8085 94144
rect 8427 94184 8469 94193
rect 8427 94144 8428 94184
rect 8468 94144 8469 94184
rect 8427 94135 8469 94144
rect 8811 94184 8853 94193
rect 8811 94144 8812 94184
rect 8852 94144 8853 94184
rect 8811 94135 8853 94144
rect 9003 94184 9045 94193
rect 9003 94144 9004 94184
rect 9044 94144 9045 94184
rect 9003 94135 9045 94144
rect 9579 94184 9621 94193
rect 9579 94144 9580 94184
rect 9620 94144 9621 94184
rect 9579 94135 9621 94144
rect 9771 94184 9813 94193
rect 9771 94144 9772 94184
rect 9812 94144 9813 94184
rect 9771 94135 9813 94144
rect 10347 94184 10389 94193
rect 10347 94144 10348 94184
rect 10388 94144 10389 94184
rect 10347 94135 10389 94144
rect 10539 94184 10581 94193
rect 10539 94144 10540 94184
rect 10580 94144 10581 94184
rect 10539 94135 10581 94144
rect 11115 94184 11157 94193
rect 11115 94144 11116 94184
rect 11156 94144 11157 94184
rect 11115 94135 11157 94144
rect 12843 94184 12885 94193
rect 12843 94144 12844 94184
rect 12884 94144 12885 94184
rect 12843 94135 12885 94144
rect 13035 94184 13077 94193
rect 13035 94144 13036 94184
rect 13076 94144 13077 94184
rect 13035 94135 13077 94144
rect 13611 94184 13653 94193
rect 13611 94144 13612 94184
rect 13652 94144 13653 94184
rect 13611 94135 13653 94144
rect 13803 94184 13845 94193
rect 13803 94144 13804 94184
rect 13844 94144 13845 94184
rect 13803 94135 13845 94144
rect 14571 94184 14613 94193
rect 14571 94144 14572 94184
rect 14612 94144 14613 94184
rect 14571 94135 14613 94144
rect 14955 94184 14997 94193
rect 14955 94144 14956 94184
rect 14996 94144 14997 94184
rect 14955 94135 14997 94144
rect 15339 94184 15381 94193
rect 15339 94144 15340 94184
rect 15380 94144 15381 94184
rect 15339 94135 15381 94144
rect 16203 94184 16245 94193
rect 16203 94144 16204 94184
rect 16244 94144 16245 94184
rect 16203 94135 16245 94144
rect 16779 94184 16821 94193
rect 16779 94144 16780 94184
rect 16820 94144 16821 94184
rect 16779 94135 16821 94144
rect 16971 94184 17013 94193
rect 16971 94144 16972 94184
rect 17012 94144 17013 94184
rect 16971 94135 17013 94144
rect 17355 94184 17397 94193
rect 17355 94144 17356 94184
rect 17396 94144 17397 94184
rect 17355 94135 17397 94144
rect 17595 94184 17637 94193
rect 17595 94144 17596 94184
rect 17636 94144 17637 94184
rect 17595 94135 17637 94144
rect 17931 94184 17973 94193
rect 17931 94144 17932 94184
rect 17972 94144 17973 94184
rect 17931 94135 17973 94144
rect 18123 94184 18165 94193
rect 18123 94144 18124 94184
rect 18164 94144 18165 94184
rect 18123 94135 18165 94144
rect 18699 94184 18741 94193
rect 18699 94144 18700 94184
rect 18740 94144 18741 94184
rect 18699 94135 18741 94144
rect 18843 94184 18885 94193
rect 18843 94144 18844 94184
rect 18884 94144 18885 94184
rect 18843 94135 18885 94144
rect 19083 94184 19125 94193
rect 19083 94144 19084 94184
rect 19124 94144 19125 94184
rect 19083 94135 19125 94144
rect 19467 94184 19509 94193
rect 19467 94144 19468 94184
rect 19508 94144 19509 94184
rect 19467 94135 19509 94144
rect 19851 94184 19893 94193
rect 19851 94144 19852 94184
rect 19892 94144 19893 94184
rect 19851 94135 19893 94144
rect 20235 94184 20277 94193
rect 20235 94144 20236 94184
rect 20276 94144 20277 94184
rect 20235 94135 20277 94144
rect 9243 94016 9285 94025
rect 9243 93976 9244 94016
rect 9284 93976 9285 94016
rect 9243 93967 9285 93976
rect 10011 94016 10053 94025
rect 10011 93976 10012 94016
rect 10052 93976 10053 94016
rect 10011 93967 10053 93976
rect 10779 94016 10821 94025
rect 10779 93976 10780 94016
rect 10820 93976 10821 94016
rect 10779 93967 10821 93976
rect 13275 94016 13317 94025
rect 13275 93976 13276 94016
rect 13316 93976 13317 94016
rect 13275 93967 13317 93976
rect 18363 94016 18405 94025
rect 18363 93976 18364 94016
rect 18404 93976 18405 94016
rect 18363 93967 18405 93976
rect 1467 93932 1509 93941
rect 1467 93892 1468 93932
rect 1508 93892 1509 93932
rect 1467 93883 1509 93892
rect 9339 93932 9381 93941
rect 9339 93892 9340 93932
rect 9380 93892 9381 93932
rect 9339 93883 9381 93892
rect 10107 93932 10149 93941
rect 10107 93892 10108 93932
rect 10148 93892 10149 93932
rect 10107 93883 10149 93892
rect 10875 93932 10917 93941
rect 10875 93892 10876 93932
rect 10916 93892 10917 93932
rect 10875 93883 10917 93892
rect 12603 93932 12645 93941
rect 12603 93892 12604 93932
rect 12644 93892 12645 93932
rect 12603 93883 12645 93892
rect 13371 93932 13413 93941
rect 13371 93892 13372 93932
rect 13412 93892 13413 93932
rect 13371 93883 13413 93892
rect 14043 93932 14085 93941
rect 14043 93892 14044 93932
rect 14084 93892 14085 93932
rect 14043 93883 14085 93892
rect 14331 93932 14373 93941
rect 14331 93892 14332 93932
rect 14372 93892 14373 93932
rect 14331 93883 14373 93892
rect 14715 93932 14757 93941
rect 14715 93892 14716 93932
rect 14756 93892 14757 93932
rect 14715 93883 14757 93892
rect 15099 93932 15141 93941
rect 15099 93892 15100 93932
rect 15140 93892 15141 93932
rect 15099 93883 15141 93892
rect 16539 93932 16581 93941
rect 16539 93892 16540 93932
rect 16580 93892 16581 93932
rect 16539 93883 16581 93892
rect 17691 93932 17733 93941
rect 17691 93892 17692 93932
rect 17732 93892 17733 93932
rect 17691 93883 17733 93892
rect 18459 93932 18501 93941
rect 18459 93892 18460 93932
rect 18500 93892 18501 93932
rect 18459 93883 18501 93892
rect 19227 93932 19269 93941
rect 19227 93892 19228 93932
rect 19268 93892 19269 93932
rect 19227 93883 19269 93892
rect 19611 93932 19653 93941
rect 19611 93892 19612 93932
rect 19652 93892 19653 93932
rect 19611 93883 19653 93892
rect 19995 93932 20037 93941
rect 19995 93892 19996 93932
rect 20036 93892 20037 93932
rect 19995 93883 20037 93892
rect 1152 93764 20452 93788
rect 1152 93724 4928 93764
rect 4968 93724 5010 93764
rect 5050 93724 5092 93764
rect 5132 93724 5174 93764
rect 5214 93724 5256 93764
rect 5296 93724 20048 93764
rect 20088 93724 20130 93764
rect 20170 93724 20212 93764
rect 20252 93724 20294 93764
rect 20334 93724 20376 93764
rect 20416 93724 20452 93764
rect 1152 93700 20452 93724
rect 2715 93596 2757 93605
rect 2715 93556 2716 93596
rect 2756 93556 2757 93596
rect 2715 93547 2757 93556
rect 18555 93596 18597 93605
rect 18555 93556 18556 93596
rect 18596 93556 18597 93596
rect 18555 93547 18597 93556
rect 19707 93596 19749 93605
rect 19707 93556 19708 93596
rect 19748 93556 19749 93596
rect 19707 93547 19749 93556
rect 2619 93512 2661 93521
rect 2619 93472 2620 93512
rect 2660 93472 2661 93512
rect 2619 93463 2661 93472
rect 18459 93512 18501 93521
rect 18459 93472 18460 93512
rect 18500 93472 18501 93512
rect 18459 93463 18501 93472
rect 1227 93344 1269 93353
rect 1227 93304 1228 93344
rect 1268 93304 1269 93344
rect 1227 93295 1269 93304
rect 1611 93344 1653 93353
rect 1611 93304 1612 93344
rect 1652 93304 1653 93344
rect 1611 93295 1653 93304
rect 1995 93344 2037 93353
rect 1995 93304 1996 93344
rect 2036 93304 2037 93344
rect 1995 93295 2037 93304
rect 2379 93344 2421 93353
rect 2379 93304 2380 93344
rect 2420 93304 2421 93344
rect 2379 93295 2421 93304
rect 2955 93344 2997 93353
rect 2955 93304 2956 93344
rect 2996 93304 2997 93344
rect 2955 93295 2997 93304
rect 3147 93344 3189 93353
rect 3147 93304 3148 93344
rect 3188 93304 3189 93344
rect 3147 93295 3189 93304
rect 17835 93344 17877 93353
rect 17835 93304 17836 93344
rect 17876 93304 17877 93344
rect 17835 93295 17877 93304
rect 18219 93344 18261 93353
rect 18219 93304 18220 93344
rect 18260 93304 18261 93344
rect 18219 93295 18261 93304
rect 18795 93344 18837 93353
rect 18795 93304 18796 93344
rect 18836 93304 18837 93344
rect 18795 93295 18837 93304
rect 18987 93344 19029 93353
rect 18987 93304 18988 93344
rect 19028 93304 19029 93344
rect 18987 93295 19029 93304
rect 19563 93344 19605 93353
rect 19563 93304 19564 93344
rect 19604 93304 19605 93344
rect 19563 93295 19605 93304
rect 19947 93344 19989 93353
rect 19947 93304 19948 93344
rect 19988 93304 19989 93344
rect 19947 93295 19989 93304
rect 20139 93344 20181 93353
rect 20139 93304 20140 93344
rect 20180 93304 20181 93344
rect 20139 93295 20181 93304
rect 18075 93260 18117 93269
rect 18075 93220 18076 93260
rect 18116 93220 18117 93260
rect 18075 93211 18117 93220
rect 19227 93260 19269 93269
rect 19227 93220 19228 93260
rect 19268 93220 19269 93260
rect 19227 93211 19269 93220
rect 1467 93176 1509 93185
rect 1467 93136 1468 93176
rect 1508 93136 1509 93176
rect 1467 93127 1509 93136
rect 1851 93176 1893 93185
rect 1851 93136 1852 93176
rect 1892 93136 1893 93176
rect 1851 93127 1893 93136
rect 2235 93176 2277 93185
rect 2235 93136 2236 93176
rect 2276 93136 2277 93176
rect 2235 93127 2277 93136
rect 3387 93176 3429 93185
rect 3387 93136 3388 93176
rect 3428 93136 3429 93176
rect 3387 93127 3429 93136
rect 19323 93176 19365 93185
rect 19323 93136 19324 93176
rect 19364 93136 19365 93176
rect 19323 93127 19365 93136
rect 20379 93176 20421 93185
rect 20379 93136 20380 93176
rect 20420 93136 20421 93176
rect 20379 93127 20421 93136
rect 1152 93008 20448 93032
rect 1152 92968 3688 93008
rect 3728 92968 3770 93008
rect 3810 92968 3852 93008
rect 3892 92968 3934 93008
rect 3974 92968 4016 93008
rect 4056 92968 18808 93008
rect 18848 92968 18890 93008
rect 18930 92968 18972 93008
rect 19012 92968 19054 93008
rect 19094 92968 19136 93008
rect 19176 92968 20448 93008
rect 1152 92944 20448 92968
rect 2715 92840 2757 92849
rect 2715 92800 2716 92840
rect 2756 92800 2757 92840
rect 2715 92791 2757 92800
rect 18939 92840 18981 92849
rect 18939 92800 18940 92840
rect 18980 92800 18981 92840
rect 18939 92791 18981 92800
rect 18843 92756 18885 92765
rect 18843 92716 18844 92756
rect 18884 92716 18885 92756
rect 18843 92707 18885 92716
rect 1227 92672 1269 92681
rect 1227 92632 1228 92672
rect 1268 92632 1269 92672
rect 1227 92623 1269 92632
rect 1611 92672 1653 92681
rect 1611 92632 1612 92672
rect 1652 92632 1653 92672
rect 1611 92623 1653 92632
rect 1995 92672 2037 92681
rect 1995 92632 1996 92672
rect 2036 92632 2037 92672
rect 1995 92623 2037 92632
rect 2235 92672 2277 92681
rect 2235 92632 2236 92672
rect 2276 92632 2277 92672
rect 2235 92623 2277 92632
rect 2379 92672 2421 92681
rect 2379 92632 2380 92672
rect 2420 92632 2421 92672
rect 2379 92623 2421 92632
rect 2955 92672 2997 92681
rect 2955 92632 2956 92672
rect 2996 92632 2997 92672
rect 2955 92623 2997 92632
rect 18603 92672 18645 92681
rect 18603 92632 18604 92672
rect 18644 92632 18645 92672
rect 18603 92623 18645 92632
rect 19179 92672 19221 92681
rect 19179 92632 19180 92672
rect 19220 92632 19221 92672
rect 19179 92623 19221 92632
rect 19563 92672 19605 92681
rect 19563 92632 19564 92672
rect 19604 92632 19605 92672
rect 19563 92623 19605 92632
rect 19755 92672 19797 92681
rect 19755 92632 19756 92672
rect 19796 92632 19797 92672
rect 19755 92623 19797 92632
rect 20139 92672 20181 92681
rect 20139 92632 20140 92672
rect 20180 92632 20181 92672
rect 20139 92623 20181 92632
rect 2619 92504 2661 92513
rect 2619 92464 2620 92504
rect 2660 92464 2661 92504
rect 2619 92455 2661 92464
rect 19323 92504 19365 92513
rect 19323 92464 19324 92504
rect 19364 92464 19365 92504
rect 19323 92455 19365 92464
rect 1467 92420 1509 92429
rect 1467 92380 1468 92420
rect 1508 92380 1509 92420
rect 1467 92371 1509 92380
rect 1851 92420 1893 92429
rect 1851 92380 1852 92420
rect 1892 92380 1893 92420
rect 1851 92371 1893 92380
rect 19995 92420 20037 92429
rect 19995 92380 19996 92420
rect 20036 92380 20037 92420
rect 19995 92371 20037 92380
rect 20379 92420 20421 92429
rect 20379 92380 20380 92420
rect 20420 92380 20421 92420
rect 20379 92371 20421 92380
rect 1152 92252 20452 92276
rect 1152 92212 4928 92252
rect 4968 92212 5010 92252
rect 5050 92212 5092 92252
rect 5132 92212 5174 92252
rect 5214 92212 5256 92252
rect 5296 92212 20048 92252
rect 20088 92212 20130 92252
rect 20170 92212 20212 92252
rect 20252 92212 20294 92252
rect 20334 92212 20376 92252
rect 20416 92212 20452 92252
rect 1152 92188 20452 92212
rect 7803 92084 7845 92093
rect 7803 92044 7804 92084
rect 7844 92044 7845 92084
rect 7803 92035 7845 92044
rect 19323 92084 19365 92093
rect 19323 92044 19324 92084
rect 19364 92044 19365 92084
rect 19323 92035 19365 92044
rect 1227 91832 1269 91841
rect 1227 91792 1228 91832
rect 1268 91792 1269 91832
rect 1227 91783 1269 91792
rect 1611 91832 1653 91841
rect 1611 91792 1612 91832
rect 1652 91792 1653 91832
rect 1611 91783 1653 91792
rect 1995 91832 2037 91841
rect 1995 91792 1996 91832
rect 2036 91792 2037 91832
rect 1995 91783 2037 91792
rect 2379 91832 2421 91841
rect 2379 91792 2380 91832
rect 2420 91792 2421 91832
rect 2379 91783 2421 91792
rect 2763 91832 2805 91841
rect 2763 91792 2764 91832
rect 2804 91792 2805 91832
rect 2763 91783 2805 91792
rect 8043 91832 8085 91841
rect 8043 91792 8044 91832
rect 8084 91792 8085 91832
rect 8043 91783 8085 91792
rect 19563 91832 19605 91841
rect 19563 91792 19564 91832
rect 19604 91792 19605 91832
rect 19563 91783 19605 91792
rect 19755 91832 19797 91841
rect 19755 91792 19756 91832
rect 19796 91792 19797 91832
rect 19755 91783 19797 91792
rect 20139 91832 20181 91841
rect 20139 91792 20140 91832
rect 20180 91792 20181 91832
rect 20139 91783 20181 91792
rect 1467 91664 1509 91673
rect 1467 91624 1468 91664
rect 1508 91624 1509 91664
rect 1467 91615 1509 91624
rect 1851 91664 1893 91673
rect 1851 91624 1852 91664
rect 1892 91624 1893 91664
rect 1851 91615 1893 91624
rect 2235 91664 2277 91673
rect 2235 91624 2236 91664
rect 2276 91624 2277 91664
rect 2235 91615 2277 91624
rect 2619 91664 2661 91673
rect 2619 91624 2620 91664
rect 2660 91624 2661 91664
rect 2619 91615 2661 91624
rect 3003 91664 3045 91673
rect 3003 91624 3004 91664
rect 3044 91624 3045 91664
rect 3003 91615 3045 91624
rect 19995 91664 20037 91673
rect 19995 91624 19996 91664
rect 20036 91624 20037 91664
rect 19995 91615 20037 91624
rect 20379 91664 20421 91673
rect 20379 91624 20380 91664
rect 20420 91624 20421 91664
rect 20379 91615 20421 91624
rect 1152 91496 20448 91520
rect 1152 91456 3688 91496
rect 3728 91456 3770 91496
rect 3810 91456 3852 91496
rect 3892 91456 3934 91496
rect 3974 91456 4016 91496
rect 4056 91456 18808 91496
rect 18848 91456 18890 91496
rect 18930 91456 18972 91496
rect 19012 91456 19054 91496
rect 19094 91456 19136 91496
rect 19176 91456 20448 91496
rect 1152 91432 20448 91456
rect 7707 91328 7749 91337
rect 7707 91288 7708 91328
rect 7748 91288 7749 91328
rect 7707 91279 7749 91288
rect 8091 91244 8133 91253
rect 8091 91204 8092 91244
rect 8132 91204 8133 91244
rect 8091 91195 8133 91204
rect 1227 91160 1269 91169
rect 1227 91120 1228 91160
rect 1268 91120 1269 91160
rect 1227 91111 1269 91120
rect 1611 91160 1653 91169
rect 1611 91120 1612 91160
rect 1652 91120 1653 91160
rect 1611 91111 1653 91120
rect 1995 91160 2037 91169
rect 1995 91120 1996 91160
rect 2036 91120 2037 91160
rect 1995 91111 2037 91120
rect 2379 91160 2421 91169
rect 2379 91120 2380 91160
rect 2420 91120 2421 91160
rect 2379 91111 2421 91120
rect 2763 91160 2805 91169
rect 2763 91120 2764 91160
rect 2804 91120 2805 91160
rect 2763 91111 2805 91120
rect 7947 91160 7989 91169
rect 7947 91120 7948 91160
rect 7988 91120 7989 91160
rect 7947 91111 7989 91120
rect 8331 91160 8373 91169
rect 8331 91120 8332 91160
rect 8372 91120 8373 91160
rect 8331 91111 8373 91120
rect 19755 91160 19797 91169
rect 19755 91120 19756 91160
rect 19796 91120 19797 91160
rect 19755 91111 19797 91120
rect 20139 91160 20181 91169
rect 20139 91120 20140 91160
rect 20180 91120 20181 91160
rect 20139 91111 20181 91120
rect 2235 90992 2277 91001
rect 2235 90952 2236 90992
rect 2276 90952 2277 90992
rect 2235 90943 2277 90952
rect 19995 90992 20037 91001
rect 19995 90952 19996 90992
rect 20036 90952 20037 90992
rect 19995 90943 20037 90952
rect 1467 90908 1509 90917
rect 1467 90868 1468 90908
rect 1508 90868 1509 90908
rect 1467 90859 1509 90868
rect 1851 90908 1893 90917
rect 1851 90868 1852 90908
rect 1892 90868 1893 90908
rect 1851 90859 1893 90868
rect 2619 90908 2661 90917
rect 2619 90868 2620 90908
rect 2660 90868 2661 90908
rect 2619 90859 2661 90868
rect 3003 90908 3045 90917
rect 3003 90868 3004 90908
rect 3044 90868 3045 90908
rect 3003 90859 3045 90868
rect 20379 90908 20421 90917
rect 20379 90868 20380 90908
rect 20420 90868 20421 90908
rect 20379 90859 20421 90868
rect 1152 90740 20452 90764
rect 1152 90700 4928 90740
rect 4968 90700 5010 90740
rect 5050 90700 5092 90740
rect 5132 90700 5174 90740
rect 5214 90700 5256 90740
rect 5296 90700 20048 90740
rect 20088 90700 20130 90740
rect 20170 90700 20212 90740
rect 20252 90700 20294 90740
rect 20334 90700 20376 90740
rect 20416 90700 20452 90740
rect 1152 90676 20452 90700
rect 17019 90572 17061 90581
rect 17019 90532 17020 90572
rect 17060 90532 17061 90572
rect 17019 90523 17061 90532
rect 11403 90404 11445 90413
rect 14379 90404 14421 90413
rect 11403 90364 11404 90404
rect 11444 90364 11445 90404
rect 11403 90355 11445 90364
rect 12651 90395 12693 90404
rect 12651 90355 12652 90395
rect 12692 90355 12693 90395
rect 14379 90364 14380 90404
rect 14420 90364 14421 90404
rect 14379 90355 14421 90364
rect 15627 90395 15669 90404
rect 15627 90355 15628 90395
rect 15668 90355 15669 90395
rect 12651 90346 12693 90355
rect 15627 90346 15669 90355
rect 1227 90320 1269 90329
rect 1227 90280 1228 90320
rect 1268 90280 1269 90320
rect 1227 90271 1269 90280
rect 1467 90320 1509 90329
rect 1467 90280 1468 90320
rect 1508 90280 1509 90320
rect 1467 90271 1509 90280
rect 1611 90320 1653 90329
rect 1611 90280 1612 90320
rect 1652 90280 1653 90320
rect 1611 90271 1653 90280
rect 1995 90320 2037 90329
rect 1995 90280 1996 90320
rect 2036 90280 2037 90320
rect 1995 90271 2037 90280
rect 2379 90320 2421 90329
rect 2379 90280 2380 90320
rect 2420 90280 2421 90320
rect 2379 90271 2421 90280
rect 2763 90320 2805 90329
rect 2763 90280 2764 90320
rect 2804 90280 2805 90320
rect 2763 90271 2805 90280
rect 3339 90320 3381 90329
rect 3339 90280 3340 90320
rect 3380 90280 3381 90320
rect 3339 90271 3381 90280
rect 3531 90320 3573 90329
rect 3531 90280 3532 90320
rect 3572 90280 3573 90320
rect 3531 90271 3573 90280
rect 3915 90320 3957 90329
rect 3915 90280 3916 90320
rect 3956 90280 3957 90320
rect 3915 90271 3957 90280
rect 17259 90320 17301 90329
rect 17259 90280 17260 90320
rect 17300 90280 17301 90320
rect 17259 90271 17301 90280
rect 19371 90320 19413 90329
rect 19371 90280 19372 90320
rect 19412 90280 19413 90320
rect 19371 90271 19413 90280
rect 19755 90320 19797 90329
rect 19755 90280 19756 90320
rect 19796 90280 19797 90320
rect 19755 90271 19797 90280
rect 20139 90320 20181 90329
rect 20139 90280 20140 90320
rect 20180 90280 20181 90320
rect 20139 90271 20181 90280
rect 1851 90236 1893 90245
rect 1851 90196 1852 90236
rect 1892 90196 1893 90236
rect 1851 90187 1893 90196
rect 3003 90236 3045 90245
rect 3003 90196 3004 90236
rect 3044 90196 3045 90236
rect 3003 90187 3045 90196
rect 20379 90236 20421 90245
rect 20379 90196 20380 90236
rect 20420 90196 20421 90236
rect 20379 90187 20421 90196
rect 2235 90152 2277 90161
rect 2235 90112 2236 90152
rect 2276 90112 2277 90152
rect 2235 90103 2277 90112
rect 2619 90152 2661 90161
rect 2619 90112 2620 90152
rect 2660 90112 2661 90152
rect 2619 90103 2661 90112
rect 3099 90152 3141 90161
rect 3099 90112 3100 90152
rect 3140 90112 3141 90152
rect 3099 90103 3141 90112
rect 3771 90152 3813 90161
rect 3771 90112 3772 90152
rect 3812 90112 3813 90152
rect 3771 90103 3813 90112
rect 4155 90152 4197 90161
rect 4155 90112 4156 90152
rect 4196 90112 4197 90152
rect 4155 90103 4197 90112
rect 12843 90152 12885 90161
rect 12843 90112 12844 90152
rect 12884 90112 12885 90152
rect 12843 90103 12885 90112
rect 15819 90152 15861 90161
rect 15819 90112 15820 90152
rect 15860 90112 15861 90152
rect 15819 90103 15861 90112
rect 19611 90152 19653 90161
rect 19611 90112 19612 90152
rect 19652 90112 19653 90152
rect 19611 90103 19653 90112
rect 19995 90152 20037 90161
rect 19995 90112 19996 90152
rect 20036 90112 20037 90152
rect 19995 90103 20037 90112
rect 1152 89984 20448 90008
rect 1152 89944 3688 89984
rect 3728 89944 3770 89984
rect 3810 89944 3852 89984
rect 3892 89944 3934 89984
rect 3974 89944 4016 89984
rect 4056 89944 18808 89984
rect 18848 89944 18890 89984
rect 18930 89944 18972 89984
rect 19012 89944 19054 89984
rect 19094 89944 19136 89984
rect 19176 89944 20448 89984
rect 1152 89920 20448 89944
rect 2619 89816 2661 89825
rect 2619 89776 2620 89816
rect 2660 89776 2661 89816
rect 2619 89767 2661 89776
rect 3771 89816 3813 89825
rect 3771 89776 3772 89816
rect 3812 89776 3813 89816
rect 3771 89767 3813 89776
rect 4155 89816 4197 89825
rect 4155 89776 4156 89816
rect 4196 89776 4197 89816
rect 4155 89767 4197 89776
rect 3003 89732 3045 89741
rect 3003 89692 3004 89732
rect 3044 89692 3045 89732
rect 3003 89683 3045 89692
rect 19995 89732 20037 89741
rect 19995 89692 19996 89732
rect 20036 89692 20037 89732
rect 19995 89683 20037 89692
rect 1227 89648 1269 89657
rect 1227 89608 1228 89648
rect 1268 89608 1269 89648
rect 1227 89599 1269 89608
rect 1611 89648 1653 89657
rect 1611 89608 1612 89648
rect 1652 89608 1653 89648
rect 1611 89599 1653 89608
rect 1995 89648 2037 89657
rect 1995 89608 1996 89648
rect 2036 89608 2037 89648
rect 1995 89599 2037 89608
rect 2379 89648 2421 89657
rect 2379 89608 2380 89648
rect 2420 89608 2421 89648
rect 2379 89599 2421 89608
rect 2763 89648 2805 89657
rect 2763 89608 2764 89648
rect 2804 89608 2805 89648
rect 2763 89599 2805 89608
rect 3147 89648 3189 89657
rect 3147 89608 3148 89648
rect 3188 89608 3189 89648
rect 3147 89599 3189 89608
rect 3531 89648 3573 89657
rect 3531 89608 3532 89648
rect 3572 89608 3573 89648
rect 3531 89599 3573 89608
rect 3915 89648 3957 89657
rect 3915 89608 3916 89648
rect 3956 89608 3957 89648
rect 3915 89599 3957 89608
rect 4299 89648 4341 89657
rect 4299 89608 4300 89648
rect 4340 89608 4341 89648
rect 4299 89599 4341 89608
rect 13611 89648 13653 89657
rect 13611 89608 13612 89648
rect 13652 89608 13653 89648
rect 13611 89599 13653 89608
rect 15034 89648 15092 89649
rect 15034 89608 15043 89648
rect 15083 89608 15092 89648
rect 15034 89607 15092 89608
rect 18987 89648 19029 89657
rect 18987 89608 18988 89648
rect 19028 89608 19029 89648
rect 18987 89599 19029 89608
rect 19371 89648 19413 89657
rect 19371 89608 19372 89648
rect 19412 89608 19413 89648
rect 19371 89599 19413 89608
rect 19755 89648 19797 89657
rect 19755 89608 19756 89648
rect 19796 89608 19797 89648
rect 19755 89599 19797 89608
rect 20139 89648 20181 89657
rect 20139 89608 20140 89648
rect 20180 89608 20181 89648
rect 20139 89599 20181 89608
rect 4683 89564 4725 89573
rect 4683 89524 4684 89564
rect 4724 89524 4725 89564
rect 4683 89515 4725 89524
rect 5923 89564 5981 89565
rect 5923 89524 5932 89564
rect 5972 89524 5981 89564
rect 5923 89523 5981 89524
rect 11403 89564 11445 89573
rect 11403 89524 11404 89564
rect 11444 89524 11445 89564
rect 11403 89515 11445 89524
rect 12643 89564 12701 89565
rect 12643 89524 12652 89564
rect 12692 89524 12701 89564
rect 12643 89523 12701 89524
rect 13114 89564 13172 89565
rect 13114 89524 13123 89564
rect 13163 89524 13172 89564
rect 13114 89523 13172 89524
rect 13227 89564 13269 89573
rect 13227 89524 13228 89564
rect 13268 89524 13269 89564
rect 13227 89515 13269 89524
rect 13707 89564 13749 89573
rect 13707 89524 13708 89564
rect 13748 89524 13749 89564
rect 13707 89515 13749 89524
rect 14179 89564 14237 89565
rect 14179 89524 14188 89564
rect 14228 89524 14237 89564
rect 14179 89523 14237 89524
rect 14698 89564 14756 89565
rect 14698 89524 14707 89564
rect 14747 89524 14756 89564
rect 14698 89523 14756 89524
rect 15235 89564 15293 89565
rect 15235 89524 15244 89564
rect 15284 89524 15293 89564
rect 15235 89523 15293 89524
rect 16491 89564 16533 89573
rect 16491 89524 16492 89564
rect 16532 89524 16533 89564
rect 16491 89515 16533 89524
rect 16875 89564 16917 89573
rect 16875 89524 16876 89564
rect 16916 89524 16917 89564
rect 16875 89515 16917 89524
rect 18115 89564 18173 89565
rect 18115 89524 18124 89564
rect 18164 89524 18173 89564
rect 18115 89523 18173 89524
rect 2235 89480 2277 89489
rect 2235 89440 2236 89480
rect 2276 89440 2277 89480
rect 2235 89431 2277 89440
rect 19227 89480 19269 89489
rect 19227 89440 19228 89480
rect 19268 89440 19269 89480
rect 19227 89431 19269 89440
rect 1467 89396 1509 89405
rect 1467 89356 1468 89396
rect 1508 89356 1509 89396
rect 1467 89347 1509 89356
rect 1851 89396 1893 89405
rect 1851 89356 1852 89396
rect 1892 89356 1893 89396
rect 1851 89347 1893 89356
rect 3387 89396 3429 89405
rect 3387 89356 3388 89396
rect 3428 89356 3429 89396
rect 3387 89347 3429 89356
rect 4539 89396 4581 89405
rect 4539 89356 4540 89396
rect 4580 89356 4581 89396
rect 4539 89347 4581 89356
rect 6123 89396 6165 89405
rect 6123 89356 6124 89396
rect 6164 89356 6165 89396
rect 6123 89347 6165 89356
rect 12843 89396 12885 89405
rect 12843 89356 12844 89396
rect 12884 89356 12885 89396
rect 12843 89347 12885 89356
rect 14859 89396 14901 89405
rect 14859 89356 14860 89396
rect 14900 89356 14901 89396
rect 14859 89347 14901 89356
rect 18315 89396 18357 89405
rect 18315 89356 18316 89396
rect 18356 89356 18357 89396
rect 18315 89347 18357 89356
rect 19611 89396 19653 89405
rect 19611 89356 19612 89396
rect 19652 89356 19653 89396
rect 19611 89347 19653 89356
rect 20379 89396 20421 89405
rect 20379 89356 20380 89396
rect 20420 89356 20421 89396
rect 20379 89347 20421 89356
rect 1152 89228 20452 89252
rect 1152 89188 4928 89228
rect 4968 89188 5010 89228
rect 5050 89188 5092 89228
rect 5132 89188 5174 89228
rect 5214 89188 5256 89228
rect 5296 89188 20048 89228
rect 20088 89188 20130 89228
rect 20170 89188 20212 89228
rect 20252 89188 20294 89228
rect 20334 89188 20376 89228
rect 20416 89188 20452 89228
rect 1152 89164 20452 89188
rect 2619 89060 2661 89069
rect 2619 89020 2620 89060
rect 2660 89020 2661 89060
rect 2619 89011 2661 89020
rect 9435 89060 9477 89069
rect 9435 89020 9436 89060
rect 9476 89020 9477 89060
rect 9435 89011 9477 89020
rect 14283 89060 14325 89069
rect 14283 89020 14284 89060
rect 14324 89020 14325 89060
rect 14283 89011 14325 89020
rect 16299 89060 16341 89069
rect 16299 89020 16300 89060
rect 16340 89020 16341 89060
rect 16299 89011 16341 89020
rect 12267 88976 12309 88985
rect 12267 88936 12268 88976
rect 12308 88936 12309 88976
rect 12267 88927 12309 88936
rect 19995 88976 20037 88985
rect 19995 88936 19996 88976
rect 20036 88936 20037 88976
rect 19995 88927 20037 88936
rect 2763 88892 2805 88901
rect 4491 88892 4533 88901
rect 8523 88892 8565 88901
rect 2763 88852 2764 88892
rect 2804 88852 2805 88892
rect 2763 88843 2805 88852
rect 4011 88883 4053 88892
rect 4011 88843 4012 88883
rect 4052 88843 4053 88883
rect 4491 88852 4492 88892
rect 4532 88852 4533 88892
rect 4491 88843 4533 88852
rect 5739 88883 5781 88892
rect 5739 88843 5740 88883
rect 5780 88843 5781 88883
rect 4011 88834 4053 88843
rect 5739 88834 5781 88843
rect 7275 88883 7317 88892
rect 7275 88843 7276 88883
rect 7316 88843 7317 88883
rect 8523 88852 8524 88892
rect 8564 88852 8565 88892
rect 8523 88843 8565 88852
rect 10827 88892 10869 88901
rect 12538 88892 12596 88893
rect 10827 88852 10828 88892
rect 10868 88852 10869 88892
rect 10827 88843 10869 88852
rect 12075 88883 12117 88892
rect 12075 88843 12076 88883
rect 12116 88843 12117 88883
rect 12538 88852 12547 88892
rect 12587 88852 12596 88892
rect 12538 88851 12596 88852
rect 12651 88892 12693 88901
rect 12651 88852 12652 88892
rect 12692 88852 12693 88892
rect 12651 88843 12693 88852
rect 13035 88892 13077 88901
rect 14554 88892 14612 88893
rect 13035 88852 13036 88892
rect 13076 88852 13077 88892
rect 13035 88843 13077 88852
rect 13611 88883 13653 88892
rect 13611 88843 13612 88883
rect 13652 88843 13653 88883
rect 7275 88834 7317 88843
rect 12075 88834 12117 88843
rect 13611 88834 13653 88843
rect 14091 88883 14133 88892
rect 14091 88843 14092 88883
rect 14132 88843 14133 88883
rect 14554 88852 14563 88892
rect 14603 88852 14612 88892
rect 14554 88851 14612 88852
rect 14667 88892 14709 88901
rect 14667 88852 14668 88892
rect 14708 88852 14709 88892
rect 14667 88843 14709 88852
rect 15051 88892 15093 88901
rect 16875 88892 16917 88901
rect 15051 88852 15052 88892
rect 15092 88852 15093 88892
rect 15051 88843 15093 88852
rect 15627 88883 15669 88892
rect 15627 88843 15628 88883
rect 15668 88843 15669 88883
rect 14091 88834 14133 88843
rect 15627 88834 15669 88843
rect 16107 88883 16149 88892
rect 16107 88843 16108 88883
rect 16148 88843 16149 88883
rect 16875 88852 16876 88892
rect 16916 88852 16917 88892
rect 16875 88843 16917 88852
rect 18123 88883 18165 88892
rect 18123 88843 18124 88883
rect 18164 88843 18165 88883
rect 16107 88834 16149 88843
rect 18123 88834 18165 88843
rect 1227 88808 1269 88817
rect 1227 88768 1228 88808
rect 1268 88768 1269 88808
rect 1227 88759 1269 88768
rect 1611 88808 1653 88817
rect 1611 88768 1612 88808
rect 1652 88768 1653 88808
rect 1611 88759 1653 88768
rect 1995 88808 2037 88817
rect 1995 88768 1996 88808
rect 2036 88768 2037 88808
rect 1995 88759 2037 88768
rect 2379 88808 2421 88817
rect 2379 88768 2380 88808
rect 2420 88768 2421 88808
rect 2379 88759 2421 88768
rect 6123 88808 6165 88817
rect 6123 88768 6124 88808
rect 6164 88768 6165 88808
rect 6123 88759 6165 88768
rect 9195 88808 9237 88817
rect 9195 88768 9196 88808
rect 9236 88768 9237 88808
rect 9195 88759 9237 88768
rect 9531 88808 9573 88817
rect 9531 88768 9532 88808
rect 9572 88768 9573 88808
rect 9531 88759 9573 88768
rect 9771 88808 9813 88817
rect 9771 88768 9772 88808
rect 9812 88768 9813 88808
rect 9771 88759 9813 88768
rect 10155 88808 10197 88817
rect 10155 88768 10156 88808
rect 10196 88768 10197 88808
rect 10155 88759 10197 88768
rect 10635 88808 10677 88817
rect 10635 88768 10636 88808
rect 10676 88768 10677 88808
rect 10635 88759 10677 88768
rect 13131 88808 13173 88817
rect 13131 88768 13132 88808
rect 13172 88768 13173 88808
rect 13131 88759 13173 88768
rect 15147 88808 15189 88817
rect 15147 88768 15148 88808
rect 15188 88768 15189 88808
rect 15147 88759 15189 88768
rect 18603 88808 18645 88817
rect 18603 88768 18604 88808
rect 18644 88768 18645 88808
rect 18603 88759 18645 88768
rect 18987 88808 19029 88817
rect 18987 88768 18988 88808
rect 19028 88768 19029 88808
rect 18987 88759 19029 88768
rect 19371 88808 19413 88817
rect 19371 88768 19372 88808
rect 19412 88768 19413 88808
rect 19371 88759 19413 88768
rect 19755 88808 19797 88817
rect 19755 88768 19756 88808
rect 19796 88768 19797 88808
rect 19755 88759 19797 88768
rect 20139 88808 20181 88817
rect 20139 88768 20140 88808
rect 20180 88768 20181 88808
rect 20139 88759 20181 88768
rect 20379 88808 20421 88817
rect 20379 88768 20380 88808
rect 20420 88768 20421 88808
rect 20379 88759 20421 88768
rect 2235 88724 2277 88733
rect 2235 88684 2236 88724
rect 2276 88684 2277 88724
rect 2235 88675 2277 88684
rect 18843 88724 18885 88733
rect 18843 88684 18844 88724
rect 18884 88684 18885 88724
rect 18843 88675 18885 88684
rect 1467 88640 1509 88649
rect 1467 88600 1468 88640
rect 1508 88600 1509 88640
rect 1467 88591 1509 88600
rect 1851 88640 1893 88649
rect 1851 88600 1852 88640
rect 1892 88600 1893 88640
rect 1851 88591 1893 88600
rect 4203 88640 4245 88649
rect 4203 88600 4204 88640
rect 4244 88600 4245 88640
rect 4203 88591 4245 88600
rect 5931 88640 5973 88649
rect 5931 88600 5932 88640
rect 5972 88600 5973 88640
rect 5931 88591 5973 88600
rect 6363 88640 6405 88649
rect 6363 88600 6364 88640
rect 6404 88600 6405 88640
rect 6363 88591 6405 88600
rect 7083 88640 7125 88649
rect 7083 88600 7084 88640
rect 7124 88600 7125 88640
rect 7083 88591 7125 88600
rect 9915 88640 9957 88649
rect 9915 88600 9916 88640
rect 9956 88600 9957 88640
rect 9915 88591 9957 88600
rect 10395 88640 10437 88649
rect 10395 88600 10396 88640
rect 10436 88600 10437 88640
rect 10395 88591 10437 88600
rect 18315 88640 18357 88649
rect 18315 88600 18316 88640
rect 18356 88600 18357 88640
rect 18315 88591 18357 88600
rect 19227 88640 19269 88649
rect 19227 88600 19228 88640
rect 19268 88600 19269 88640
rect 19227 88591 19269 88600
rect 19611 88640 19653 88649
rect 19611 88600 19612 88640
rect 19652 88600 19653 88640
rect 19611 88591 19653 88600
rect 1152 88472 20448 88496
rect 1152 88432 3688 88472
rect 3728 88432 3770 88472
rect 3810 88432 3852 88472
rect 3892 88432 3934 88472
rect 3974 88432 4016 88472
rect 4056 88432 18808 88472
rect 18848 88432 18890 88472
rect 18930 88432 18972 88472
rect 19012 88432 19054 88472
rect 19094 88432 19136 88472
rect 19176 88432 20448 88472
rect 1152 88408 20448 88432
rect 8667 88304 8709 88313
rect 8667 88264 8668 88304
rect 8708 88264 8709 88304
rect 8667 88255 8709 88264
rect 12171 88304 12213 88313
rect 12171 88264 12172 88304
rect 12212 88264 12213 88304
rect 12171 88255 12213 88264
rect 12795 88304 12837 88313
rect 12795 88264 12796 88304
rect 12836 88264 12837 88304
rect 12795 88255 12837 88264
rect 9099 88220 9141 88229
rect 9099 88180 9100 88220
rect 9140 88180 9141 88220
rect 9099 88171 9141 88180
rect 1227 88136 1269 88145
rect 1227 88096 1228 88136
rect 1268 88096 1269 88136
rect 1227 88087 1269 88096
rect 1899 88136 1941 88145
rect 1899 88096 1900 88136
rect 1940 88096 1941 88136
rect 1899 88087 1941 88096
rect 2283 88136 2325 88145
rect 2283 88096 2284 88136
rect 2324 88096 2325 88136
rect 2283 88087 2325 88096
rect 4395 88136 4437 88145
rect 4395 88096 4396 88136
rect 4436 88096 4437 88136
rect 4395 88087 4437 88096
rect 5355 88136 5397 88145
rect 5355 88096 5356 88136
rect 5396 88096 5397 88136
rect 5355 88087 5397 88096
rect 8907 88136 8949 88145
rect 8907 88096 8908 88136
rect 8948 88096 8949 88136
rect 8907 88087 8949 88096
rect 12555 88136 12597 88145
rect 12555 88096 12556 88136
rect 12596 88096 12597 88136
rect 12555 88087 12597 88096
rect 13515 88136 13557 88145
rect 13515 88096 13516 88136
rect 13556 88096 13557 88136
rect 13515 88087 13557 88096
rect 18219 88136 18261 88145
rect 18219 88096 18220 88136
rect 18260 88096 18261 88136
rect 18219 88087 18261 88096
rect 2763 88052 2805 88061
rect 2763 88012 2764 88052
rect 2804 88012 2805 88052
rect 2763 88003 2805 88012
rect 4003 88052 4061 88053
rect 4003 88012 4012 88052
rect 4052 88012 4061 88052
rect 4003 88011 4061 88012
rect 4858 88052 4916 88053
rect 4858 88012 4867 88052
rect 4907 88012 4916 88052
rect 4858 88011 4916 88012
rect 4971 88052 5013 88061
rect 4971 88012 4972 88052
rect 5012 88012 5013 88052
rect 4971 88003 5013 88012
rect 5451 88052 5493 88061
rect 5451 88012 5452 88052
rect 5492 88012 5493 88052
rect 5451 88003 5493 88012
rect 5923 88052 5981 88053
rect 5923 88012 5932 88052
rect 5972 88012 5981 88052
rect 5923 88011 5981 88012
rect 6411 88052 6469 88053
rect 6411 88012 6420 88052
rect 6460 88012 6469 88052
rect 6411 88011 6469 88012
rect 6979 88052 7037 88053
rect 6979 88012 6988 88052
rect 7028 88012 7037 88052
rect 6979 88011 7037 88012
rect 8235 88052 8277 88061
rect 8235 88012 8236 88052
rect 8276 88012 8277 88052
rect 8235 88003 8277 88012
rect 9283 88052 9341 88053
rect 9283 88012 9292 88052
rect 9332 88012 9341 88052
rect 9283 88011 9341 88012
rect 10539 88052 10581 88061
rect 10539 88012 10540 88052
rect 10580 88012 10581 88052
rect 10539 88003 10581 88012
rect 10731 88052 10773 88061
rect 10731 88012 10732 88052
rect 10772 88012 10773 88052
rect 10731 88003 10773 88012
rect 11979 88052 12037 88053
rect 11979 88012 11988 88052
rect 12028 88012 12037 88052
rect 11979 88011 12037 88012
rect 13018 88052 13076 88053
rect 13018 88012 13027 88052
rect 13067 88012 13076 88052
rect 13018 88011 13076 88012
rect 13131 88052 13173 88061
rect 13131 88012 13132 88052
rect 13172 88012 13173 88052
rect 13131 88003 13173 88012
rect 13611 88052 13653 88061
rect 13611 88012 13612 88052
rect 13652 88012 13653 88052
rect 13611 88003 13653 88012
rect 14083 88052 14141 88053
rect 14083 88012 14092 88052
rect 14132 88012 14141 88052
rect 14083 88011 14141 88012
rect 14602 88052 14660 88053
rect 14602 88012 14611 88052
rect 14651 88012 14660 88052
rect 14602 88011 14660 88012
rect 15139 88052 15197 88053
rect 15139 88012 15148 88052
rect 15188 88012 15197 88052
rect 15139 88011 15197 88012
rect 16395 88052 16437 88061
rect 16395 88012 16396 88052
rect 16436 88012 16437 88052
rect 16395 88003 16437 88012
rect 16587 88052 16629 88061
rect 16587 88012 16588 88052
rect 16628 88012 16629 88052
rect 16587 88003 16629 88012
rect 17827 88052 17885 88053
rect 17827 88012 17836 88052
rect 17876 88012 17885 88052
rect 17827 88011 17885 88012
rect 18603 88052 18645 88061
rect 18603 88012 18604 88052
rect 18644 88012 18645 88052
rect 18603 88003 18645 88012
rect 19843 88052 19901 88053
rect 19843 88012 19852 88052
rect 19892 88012 19901 88052
rect 19843 88011 19901 88012
rect 2139 87968 2181 87977
rect 2139 87928 2140 87968
rect 2180 87928 2181 87968
rect 2139 87919 2181 87928
rect 4203 87968 4245 87977
rect 4203 87928 4204 87968
rect 4244 87928 4245 87968
rect 4203 87919 4245 87928
rect 14955 87968 14997 87977
rect 14955 87928 14956 87968
rect 14996 87928 14997 87968
rect 14955 87919 14997 87928
rect 18027 87968 18069 87977
rect 18027 87928 18028 87968
rect 18068 87928 18069 87968
rect 18027 87919 18069 87928
rect 1467 87884 1509 87893
rect 1467 87844 1468 87884
rect 1508 87844 1509 87884
rect 1467 87835 1509 87844
rect 2523 87884 2565 87893
rect 2523 87844 2524 87884
rect 2564 87844 2565 87884
rect 2523 87835 2565 87844
rect 4635 87884 4677 87893
rect 4635 87844 4636 87884
rect 4676 87844 4677 87884
rect 4635 87835 4677 87844
rect 6603 87884 6645 87893
rect 6603 87844 6604 87884
rect 6644 87844 6645 87884
rect 6603 87835 6645 87844
rect 6795 87884 6837 87893
rect 6795 87844 6796 87884
rect 6836 87844 6837 87884
rect 6795 87835 6837 87844
rect 14763 87884 14805 87893
rect 14763 87844 14764 87884
rect 14804 87844 14805 87884
rect 14763 87835 14805 87844
rect 18459 87884 18501 87893
rect 18459 87844 18460 87884
rect 18500 87844 18501 87884
rect 18459 87835 18501 87844
rect 20043 87884 20085 87893
rect 20043 87844 20044 87884
rect 20084 87844 20085 87884
rect 20043 87835 20085 87844
rect 1152 87716 20452 87740
rect 1152 87676 4928 87716
rect 4968 87676 5010 87716
rect 5050 87676 5092 87716
rect 5132 87676 5174 87716
rect 5214 87676 5256 87716
rect 5296 87676 20048 87716
rect 20088 87676 20130 87716
rect 20170 87676 20212 87716
rect 20252 87676 20294 87716
rect 20334 87676 20376 87716
rect 20416 87676 20452 87716
rect 1152 87652 20452 87676
rect 6603 87548 6645 87557
rect 6603 87508 6604 87548
rect 6644 87508 6645 87548
rect 6603 87499 6645 87508
rect 8715 87548 8757 87557
rect 8715 87508 8716 87548
rect 8756 87508 8757 87548
rect 8715 87499 8757 87508
rect 13515 87548 13557 87557
rect 13515 87508 13516 87548
rect 13556 87508 13557 87548
rect 13515 87499 13557 87508
rect 3867 87464 3909 87473
rect 3867 87424 3868 87464
rect 3908 87424 3909 87464
rect 3867 87415 3909 87424
rect 8907 87464 8949 87473
rect 8907 87424 8908 87464
rect 8948 87424 8949 87464
rect 8907 87415 8949 87424
rect 17434 87464 17492 87465
rect 17434 87424 17443 87464
rect 17483 87424 17492 87464
rect 17434 87423 17492 87424
rect 1611 87380 1653 87389
rect 4845 87380 4887 87389
rect 1611 87340 1612 87380
rect 1652 87340 1653 87380
rect 1611 87331 1653 87340
rect 2859 87371 2901 87380
rect 2859 87331 2860 87371
rect 2900 87331 2901 87371
rect 4845 87340 4846 87380
rect 4886 87340 4887 87380
rect 4845 87331 4887 87340
rect 4971 87380 5013 87389
rect 4971 87340 4972 87380
rect 5012 87340 5013 87380
rect 4971 87331 5013 87340
rect 5355 87380 5397 87389
rect 6970 87380 7028 87381
rect 5355 87340 5356 87380
rect 5396 87340 5397 87380
rect 5355 87331 5397 87340
rect 5931 87371 5973 87380
rect 5931 87331 5932 87371
rect 5972 87331 5973 87371
rect 2859 87322 2901 87331
rect 5931 87322 5973 87331
rect 6411 87371 6453 87380
rect 6411 87331 6412 87371
rect 6452 87331 6453 87371
rect 6970 87340 6979 87380
rect 7019 87340 7028 87380
rect 6970 87339 7028 87340
rect 7083 87380 7125 87389
rect 7083 87340 7084 87380
rect 7124 87340 7125 87380
rect 7083 87331 7125 87340
rect 7467 87380 7509 87389
rect 10347 87380 10389 87389
rect 7467 87340 7468 87380
rect 7508 87340 7509 87380
rect 7467 87331 7509 87340
rect 8043 87371 8085 87380
rect 8043 87331 8044 87371
rect 8084 87331 8085 87371
rect 6411 87322 6453 87331
rect 8043 87322 8085 87331
rect 8523 87371 8565 87380
rect 8523 87331 8524 87371
rect 8564 87331 8565 87371
rect 8523 87322 8565 87331
rect 9099 87371 9141 87380
rect 9099 87331 9100 87371
rect 9140 87331 9141 87371
rect 10347 87340 10348 87380
rect 10388 87340 10389 87380
rect 10347 87331 10389 87340
rect 11115 87380 11157 87389
rect 12747 87380 12789 87389
rect 11115 87340 11116 87380
rect 11156 87340 11157 87380
rect 11115 87331 11157 87340
rect 12363 87371 12405 87380
rect 12363 87331 12364 87371
rect 12404 87331 12405 87371
rect 12747 87340 12748 87380
rect 12788 87340 12789 87380
rect 12747 87331 12789 87340
rect 12862 87380 12904 87389
rect 12862 87340 12863 87380
rect 12903 87340 12904 87380
rect 12862 87331 12904 87340
rect 13035 87380 13077 87389
rect 13035 87340 13036 87380
rect 13076 87340 13077 87380
rect 13035 87331 13077 87340
rect 13258 87380 13316 87381
rect 13258 87340 13267 87380
rect 13307 87340 13316 87380
rect 15723 87380 15765 87389
rect 17626 87380 17684 87381
rect 18603 87380 18645 87389
rect 13258 87339 13316 87340
rect 13360 87348 13418 87349
rect 9099 87322 9141 87331
rect 12363 87322 12405 87331
rect 13360 87308 13369 87348
rect 13409 87308 13418 87348
rect 15723 87340 15724 87380
rect 15764 87340 15765 87380
rect 15723 87331 15765 87340
rect 16971 87371 17013 87380
rect 16971 87331 16972 87371
rect 17012 87331 17013 87371
rect 17626 87340 17635 87380
rect 17675 87340 17684 87380
rect 17626 87339 17684 87340
rect 18123 87371 18165 87380
rect 16971 87322 17013 87331
rect 18123 87331 18124 87371
rect 18164 87331 18165 87371
rect 18603 87340 18604 87380
rect 18644 87340 18645 87380
rect 18603 87331 18645 87340
rect 19083 87380 19125 87389
rect 19083 87340 19084 87380
rect 19124 87340 19125 87380
rect 19083 87331 19125 87340
rect 19193 87380 19251 87381
rect 19193 87340 19202 87380
rect 19242 87340 19251 87380
rect 19193 87339 19251 87340
rect 18123 87322 18165 87331
rect 13360 87307 13418 87308
rect 1227 87296 1269 87305
rect 1227 87256 1228 87296
rect 1268 87256 1269 87296
rect 1227 87247 1269 87256
rect 3435 87296 3477 87305
rect 3435 87256 3436 87296
rect 3476 87256 3477 87296
rect 3435 87247 3477 87256
rect 3627 87296 3669 87305
rect 3627 87256 3628 87296
rect 3668 87256 3669 87296
rect 3627 87247 3669 87256
rect 4011 87296 4053 87305
rect 4011 87256 4012 87296
rect 4052 87256 4053 87296
rect 4011 87247 4053 87256
rect 4587 87296 4629 87305
rect 4587 87256 4588 87296
rect 4628 87256 4629 87296
rect 4587 87247 4629 87256
rect 5451 87296 5493 87305
rect 5451 87256 5452 87296
rect 5492 87256 5493 87296
rect 5451 87247 5493 87256
rect 7563 87296 7605 87305
rect 7563 87256 7564 87296
rect 7604 87256 7605 87296
rect 7563 87247 7605 87256
rect 10731 87296 10773 87305
rect 10731 87256 10732 87296
rect 10772 87256 10773 87296
rect 10731 87247 10773 87256
rect 18699 87296 18741 87305
rect 18699 87256 18700 87296
rect 18740 87256 18741 87296
rect 18699 87247 18741 87256
rect 19755 87296 19797 87305
rect 19755 87256 19756 87296
rect 19796 87256 19797 87296
rect 19755 87247 19797 87256
rect 20139 87296 20181 87305
rect 20139 87256 20140 87296
rect 20180 87256 20181 87296
rect 20139 87247 20181 87256
rect 20379 87296 20421 87305
rect 20379 87256 20380 87296
rect 20420 87256 20421 87296
rect 20379 87247 20421 87256
rect 4251 87212 4293 87221
rect 4251 87172 4252 87212
rect 4292 87172 4293 87212
rect 4251 87163 4293 87172
rect 12555 87212 12597 87221
rect 12555 87172 12556 87212
rect 12596 87172 12597 87212
rect 12555 87163 12597 87172
rect 1467 87128 1509 87137
rect 1467 87088 1468 87128
rect 1508 87088 1509 87128
rect 1467 87079 1509 87088
rect 3051 87128 3093 87137
rect 3051 87088 3052 87128
rect 3092 87088 3093 87128
rect 3051 87079 3093 87088
rect 3195 87128 3237 87137
rect 3195 87088 3196 87128
rect 3236 87088 3237 87128
rect 3195 87079 3237 87088
rect 4347 87128 4389 87137
rect 4347 87088 4348 87128
rect 4388 87088 4389 87128
rect 4347 87079 4389 87088
rect 10971 87128 11013 87137
rect 10971 87088 10972 87128
rect 11012 87088 11013 87128
rect 10971 87079 11013 87088
rect 12747 87128 12789 87137
rect 12747 87088 12748 87128
rect 12788 87088 12789 87128
rect 12747 87079 12789 87088
rect 17163 87128 17205 87137
rect 17163 87088 17164 87128
rect 17204 87088 17205 87128
rect 17163 87079 17205 87088
rect 19995 87128 20037 87137
rect 19995 87088 19996 87128
rect 20036 87088 20037 87128
rect 19995 87079 20037 87088
rect 1152 86960 20448 86984
rect 1152 86920 3688 86960
rect 3728 86920 3770 86960
rect 3810 86920 3852 86960
rect 3892 86920 3934 86960
rect 3974 86920 4016 86960
rect 4056 86920 18808 86960
rect 18848 86920 18890 86960
rect 18930 86920 18972 86960
rect 19012 86920 19054 86960
rect 19094 86920 19136 86960
rect 19176 86920 20448 86960
rect 1152 86896 20448 86920
rect 2763 86792 2805 86801
rect 2763 86752 2764 86792
rect 2804 86752 2805 86792
rect 2763 86743 2805 86752
rect 6843 86792 6885 86801
rect 6843 86752 6844 86792
rect 6884 86752 6885 86792
rect 6843 86743 6885 86752
rect 9226 86792 9284 86793
rect 9226 86752 9235 86792
rect 9275 86752 9284 86792
rect 9226 86751 9284 86752
rect 9627 86792 9669 86801
rect 9627 86752 9628 86792
rect 9668 86752 9669 86792
rect 9627 86743 9669 86752
rect 10299 86792 10341 86801
rect 10299 86752 10300 86792
rect 10340 86752 10341 86792
rect 10299 86743 10341 86752
rect 10683 86792 10725 86801
rect 10683 86752 10684 86792
rect 10724 86752 10725 86792
rect 10683 86743 10725 86752
rect 12267 86792 12309 86801
rect 12267 86752 12268 86792
rect 12308 86752 12309 86792
rect 12267 86743 12309 86752
rect 5163 86624 5205 86633
rect 5163 86584 5164 86624
rect 5204 86584 5205 86624
rect 5163 86575 5205 86584
rect 6603 86624 6645 86633
rect 6603 86584 6604 86624
rect 6644 86584 6645 86624
rect 6603 86575 6645 86584
rect 6987 86624 7029 86633
rect 6987 86584 6988 86624
rect 7028 86584 7029 86624
rect 6987 86575 7029 86584
rect 7947 86624 7989 86633
rect 7947 86584 7948 86624
rect 7988 86584 7989 86624
rect 7947 86575 7989 86584
rect 9387 86624 9429 86633
rect 9387 86584 9388 86624
rect 9428 86584 9429 86624
rect 9387 86575 9429 86584
rect 10059 86624 10101 86633
rect 10059 86584 10060 86624
rect 10100 86584 10101 86624
rect 10059 86575 10101 86584
rect 10443 86624 10485 86633
rect 10443 86584 10444 86624
rect 10484 86584 10485 86624
rect 10443 86575 10485 86584
rect 12459 86624 12501 86633
rect 12459 86584 12460 86624
rect 12500 86584 12501 86624
rect 12459 86575 12501 86584
rect 18027 86624 18069 86633
rect 18027 86584 18028 86624
rect 18068 86584 18069 86624
rect 18027 86575 18069 86584
rect 19755 86624 19797 86633
rect 19755 86584 19756 86624
rect 19796 86584 19797 86624
rect 19755 86575 19797 86584
rect 20139 86624 20181 86633
rect 20139 86584 20140 86624
rect 20180 86584 20181 86624
rect 20139 86575 20181 86584
rect 1323 86540 1365 86549
rect 1323 86500 1324 86540
rect 1364 86500 1365 86540
rect 1323 86491 1365 86500
rect 2563 86540 2621 86541
rect 2563 86500 2572 86540
rect 2612 86500 2621 86540
rect 2563 86499 2621 86500
rect 2955 86540 2997 86549
rect 2955 86500 2956 86540
rect 2996 86500 2997 86540
rect 2955 86491 2997 86500
rect 4195 86540 4253 86541
rect 4195 86500 4204 86540
rect 4244 86500 4253 86540
rect 4195 86499 4253 86500
rect 4666 86540 4724 86541
rect 4666 86500 4675 86540
rect 4715 86500 4724 86540
rect 4666 86499 4724 86500
rect 4779 86540 4821 86549
rect 4779 86500 4780 86540
rect 4820 86500 4821 86540
rect 4779 86491 4821 86500
rect 5259 86540 5301 86549
rect 5259 86500 5260 86540
rect 5300 86500 5301 86540
rect 5259 86491 5301 86500
rect 5731 86540 5789 86541
rect 5731 86500 5740 86540
rect 5780 86500 5789 86540
rect 5731 86499 5789 86500
rect 6219 86540 6277 86541
rect 6219 86500 6228 86540
rect 6268 86500 6277 86540
rect 6219 86499 6277 86500
rect 7437 86540 7479 86549
rect 7437 86500 7438 86540
rect 7478 86500 7479 86540
rect 7437 86491 7479 86500
rect 7563 86540 7605 86549
rect 7563 86500 7564 86540
rect 7604 86500 7605 86540
rect 7563 86491 7605 86500
rect 8043 86540 8085 86549
rect 8043 86500 8044 86540
rect 8084 86500 8085 86540
rect 8043 86491 8085 86500
rect 8514 86540 8572 86541
rect 8514 86500 8523 86540
rect 8563 86500 8572 86540
rect 8514 86499 8572 86500
rect 9003 86540 9061 86541
rect 9003 86500 9012 86540
rect 9052 86500 9061 86540
rect 9003 86499 9061 86500
rect 10827 86540 10869 86549
rect 10827 86500 10828 86540
rect 10868 86500 10869 86540
rect 10827 86491 10869 86500
rect 12067 86540 12125 86541
rect 12067 86500 12076 86540
rect 12116 86500 12125 86540
rect 12067 86499 12125 86500
rect 12826 86540 12884 86541
rect 12826 86500 12835 86540
rect 12875 86500 12884 86540
rect 12826 86499 12884 86500
rect 12944 86540 13002 86541
rect 12944 86500 12953 86540
rect 12993 86500 13002 86540
rect 12944 86499 13002 86500
rect 13076 86540 13134 86541
rect 13076 86500 13085 86540
rect 13125 86500 13134 86540
rect 13076 86499 13134 86500
rect 13210 86540 13268 86541
rect 13210 86500 13219 86540
rect 13259 86500 13268 86540
rect 13210 86499 13268 86500
rect 13354 86540 13412 86541
rect 13354 86500 13363 86540
rect 13403 86500 13412 86540
rect 13354 86499 13412 86500
rect 13899 86540 13941 86549
rect 13899 86500 13900 86540
rect 13940 86500 13941 86540
rect 13899 86491 13941 86500
rect 15139 86540 15197 86541
rect 15139 86500 15148 86540
rect 15188 86500 15197 86540
rect 15139 86499 15197 86500
rect 15531 86540 15573 86549
rect 15531 86500 15532 86540
rect 15572 86500 15573 86540
rect 15531 86491 15573 86500
rect 16771 86540 16829 86541
rect 16771 86500 16780 86540
rect 16820 86500 16829 86540
rect 16771 86499 16829 86500
rect 17530 86540 17588 86541
rect 17530 86500 17539 86540
rect 17579 86500 17588 86540
rect 17530 86499 17588 86500
rect 17643 86540 17685 86549
rect 17643 86500 17644 86540
rect 17684 86500 17685 86540
rect 17643 86491 17685 86500
rect 18123 86540 18165 86549
rect 18123 86500 18124 86540
rect 18164 86500 18165 86540
rect 18123 86491 18165 86500
rect 18595 86540 18653 86541
rect 18595 86500 18604 86540
rect 18644 86500 18653 86540
rect 18595 86499 18653 86500
rect 19083 86540 19141 86541
rect 19083 86500 19092 86540
rect 19132 86500 19141 86540
rect 19083 86499 19141 86500
rect 4395 86456 4437 86465
rect 4395 86416 4396 86456
rect 4436 86416 4437 86456
rect 4395 86407 4437 86416
rect 12267 86456 12309 86465
rect 12267 86416 12268 86456
rect 12308 86416 12309 86456
rect 12267 86407 12309 86416
rect 15339 86456 15381 86465
rect 15339 86416 15340 86456
rect 15380 86416 15381 86456
rect 15339 86407 15381 86416
rect 16971 86456 17013 86465
rect 16971 86416 16972 86456
rect 17012 86416 17013 86456
rect 16971 86407 17013 86416
rect 20379 86456 20421 86465
rect 20379 86416 20380 86456
rect 20420 86416 20421 86456
rect 20379 86407 20421 86416
rect 6411 86372 6453 86381
rect 6411 86332 6412 86372
rect 6452 86332 6453 86372
rect 6411 86323 6453 86332
rect 7227 86372 7269 86381
rect 7227 86332 7228 86372
rect 7268 86332 7269 86372
rect 7227 86323 7269 86332
rect 12699 86372 12741 86381
rect 12699 86332 12700 86372
rect 12740 86332 12741 86372
rect 12699 86323 12741 86332
rect 13035 86372 13077 86381
rect 13035 86332 13036 86372
rect 13076 86332 13077 86372
rect 13035 86323 13077 86332
rect 19275 86372 19317 86381
rect 19275 86332 19276 86372
rect 19316 86332 19317 86372
rect 19275 86323 19317 86332
rect 19995 86372 20037 86381
rect 19995 86332 19996 86372
rect 20036 86332 20037 86372
rect 19995 86323 20037 86332
rect 1152 86204 20452 86228
rect 1152 86164 4928 86204
rect 4968 86164 5010 86204
rect 5050 86164 5092 86204
rect 5132 86164 5174 86204
rect 5214 86164 5256 86204
rect 5296 86164 20048 86204
rect 20088 86164 20130 86204
rect 20170 86164 20212 86204
rect 20252 86164 20294 86204
rect 20334 86164 20376 86204
rect 20416 86164 20452 86204
rect 1152 86140 20452 86164
rect 3963 86036 4005 86045
rect 3963 85996 3964 86036
rect 4004 85996 4005 86036
rect 3963 85987 4005 85996
rect 5835 86036 5877 86045
rect 5835 85996 5836 86036
rect 5876 85996 5877 86036
rect 5835 85987 5877 85996
rect 6747 86036 6789 86045
rect 6747 85996 6748 86036
rect 6788 85996 6789 86036
rect 6747 85987 6789 85996
rect 8619 86036 8661 86045
rect 8619 85996 8620 86036
rect 8660 85996 8661 86036
rect 8619 85987 8661 85996
rect 12507 86036 12549 86045
rect 12507 85996 12508 86036
rect 12548 85996 12549 86036
rect 12507 85987 12549 85996
rect 3579 85952 3621 85961
rect 3579 85912 3580 85952
rect 3620 85912 3621 85952
rect 3579 85903 3621 85912
rect 18171 85952 18213 85961
rect 18171 85912 18172 85952
rect 18212 85912 18213 85952
rect 18171 85903 18213 85912
rect 1707 85868 1749 85877
rect 4395 85868 4437 85877
rect 7179 85868 7221 85877
rect 8811 85868 8853 85877
rect 10443 85868 10485 85877
rect 12363 85868 12405 85877
rect 1707 85828 1708 85868
rect 1748 85828 1749 85868
rect 1707 85819 1749 85828
rect 2955 85859 2997 85868
rect 2955 85819 2956 85859
rect 2996 85819 2997 85859
rect 4395 85828 4396 85868
rect 4436 85828 4437 85868
rect 4395 85819 4437 85828
rect 5643 85859 5685 85868
rect 5643 85819 5644 85859
rect 5684 85819 5685 85859
rect 7179 85828 7180 85868
rect 7220 85828 7221 85868
rect 7179 85819 7221 85828
rect 8427 85859 8469 85868
rect 8427 85819 8428 85859
rect 8468 85819 8469 85859
rect 8811 85828 8812 85868
rect 8852 85828 8853 85868
rect 8811 85819 8853 85828
rect 10059 85859 10101 85868
rect 10059 85819 10060 85859
rect 10100 85819 10101 85859
rect 10443 85828 10444 85868
rect 10484 85828 10485 85868
rect 10443 85819 10485 85828
rect 11691 85859 11733 85868
rect 11691 85819 11692 85859
rect 11732 85819 11733 85859
rect 12363 85828 12364 85868
rect 12404 85828 12405 85868
rect 12363 85819 12405 85828
rect 12651 85868 12693 85877
rect 12651 85828 12652 85868
rect 12692 85828 12693 85868
rect 12651 85819 12693 85828
rect 12826 85868 12884 85869
rect 12826 85828 12835 85868
rect 12875 85828 12884 85868
rect 12826 85827 12884 85828
rect 13131 85868 13173 85877
rect 13131 85828 13132 85868
rect 13172 85828 13173 85868
rect 13131 85819 13173 85828
rect 13360 85868 13418 85869
rect 13360 85828 13369 85868
rect 13409 85828 13418 85868
rect 13360 85827 13418 85828
rect 13515 85868 13557 85877
rect 13515 85828 13516 85868
rect 13556 85828 13557 85868
rect 13515 85819 13557 85828
rect 13803 85868 13845 85877
rect 15435 85868 15477 85877
rect 18603 85868 18645 85877
rect 13803 85828 13804 85868
rect 13844 85828 13845 85868
rect 13803 85819 13845 85828
rect 15051 85859 15093 85868
rect 15051 85819 15052 85859
rect 15092 85819 15093 85859
rect 15435 85828 15436 85868
rect 15476 85828 15477 85868
rect 15435 85819 15477 85828
rect 16683 85859 16725 85868
rect 16683 85819 16684 85859
rect 16724 85819 16725 85859
rect 18603 85828 18604 85868
rect 18644 85828 18645 85868
rect 18603 85819 18645 85828
rect 19851 85859 19893 85868
rect 19851 85819 19852 85859
rect 19892 85819 19893 85859
rect 2955 85810 2997 85819
rect 5643 85810 5685 85819
rect 8427 85810 8469 85819
rect 10059 85810 10101 85819
rect 11691 85810 11733 85819
rect 15051 85810 15093 85819
rect 16683 85810 16725 85819
rect 19851 85810 19893 85819
rect 1227 85784 1269 85793
rect 1227 85744 1228 85784
rect 1268 85744 1269 85784
rect 1227 85735 1269 85744
rect 3339 85784 3381 85793
rect 3339 85744 3340 85784
rect 3380 85744 3381 85784
rect 3339 85735 3381 85744
rect 3723 85784 3765 85793
rect 3723 85744 3724 85784
rect 3764 85744 3765 85784
rect 3723 85735 3765 85744
rect 6075 85784 6117 85793
rect 6075 85744 6076 85784
rect 6116 85744 6117 85784
rect 6075 85735 6117 85744
rect 6315 85784 6357 85793
rect 6315 85744 6316 85784
rect 6356 85744 6357 85784
rect 6315 85735 6357 85744
rect 6507 85784 6549 85793
rect 6507 85744 6508 85784
rect 6548 85744 6549 85784
rect 6507 85735 6549 85744
rect 13035 85784 13077 85793
rect 17259 85784 17301 85793
rect 13035 85744 13036 85784
rect 13076 85744 13077 85784
rect 13035 85735 13077 85744
rect 13266 85775 13312 85784
rect 13266 85735 13267 85775
rect 13307 85735 13312 85775
rect 17259 85744 17260 85784
rect 17300 85744 17301 85784
rect 17259 85735 17301 85744
rect 17451 85784 17493 85793
rect 17451 85744 17452 85784
rect 17492 85744 17493 85784
rect 17451 85735 17493 85744
rect 17835 85784 17877 85793
rect 17835 85744 17836 85784
rect 17876 85744 17877 85784
rect 17835 85735 17877 85744
rect 18411 85784 18453 85793
rect 18411 85744 18412 85784
rect 18452 85744 18453 85784
rect 18411 85735 18453 85744
rect 13266 85726 13312 85735
rect 17019 85700 17061 85709
rect 17019 85660 17020 85700
rect 17060 85660 17061 85700
rect 17019 85651 17061 85660
rect 18075 85700 18117 85709
rect 18075 85660 18076 85700
rect 18116 85660 18117 85700
rect 18075 85651 18117 85660
rect 1467 85616 1509 85625
rect 1467 85576 1468 85616
rect 1508 85576 1509 85616
rect 1467 85567 1509 85576
rect 3147 85616 3189 85625
rect 3147 85576 3148 85616
rect 3188 85576 3189 85616
rect 3147 85567 3189 85576
rect 10251 85616 10293 85625
rect 10251 85576 10252 85616
rect 10292 85576 10293 85616
rect 10251 85567 10293 85576
rect 11883 85616 11925 85625
rect 11883 85576 11884 85616
rect 11924 85576 11925 85616
rect 11883 85567 11925 85576
rect 12826 85616 12884 85617
rect 12826 85576 12835 85616
rect 12875 85576 12884 85616
rect 12826 85575 12884 85576
rect 13659 85616 13701 85625
rect 13659 85576 13660 85616
rect 13700 85576 13701 85616
rect 13659 85567 13701 85576
rect 15243 85616 15285 85625
rect 15243 85576 15244 85616
rect 15284 85576 15285 85616
rect 15243 85567 15285 85576
rect 16875 85616 16917 85625
rect 16875 85576 16876 85616
rect 16916 85576 16917 85616
rect 16875 85567 16917 85576
rect 17691 85616 17733 85625
rect 17691 85576 17692 85616
rect 17732 85576 17733 85616
rect 17691 85567 17733 85576
rect 20043 85616 20085 85625
rect 20043 85576 20044 85616
rect 20084 85576 20085 85616
rect 20043 85567 20085 85576
rect 1152 85448 20448 85472
rect 1152 85408 3688 85448
rect 3728 85408 3770 85448
rect 3810 85408 3852 85448
rect 3892 85408 3934 85448
rect 3974 85408 4016 85448
rect 4056 85408 18808 85448
rect 18848 85408 18890 85448
rect 18930 85408 18972 85448
rect 19012 85408 19054 85448
rect 19094 85408 19136 85448
rect 19176 85408 20448 85448
rect 1152 85384 20448 85408
rect 8187 85280 8229 85289
rect 8187 85240 8188 85280
rect 8228 85240 8229 85280
rect 8187 85231 8229 85240
rect 8859 85280 8901 85289
rect 8859 85240 8860 85280
rect 8900 85240 8901 85280
rect 8859 85231 8901 85240
rect 4875 85196 4917 85205
rect 4875 85156 4876 85196
rect 4916 85156 4917 85196
rect 4875 85147 4917 85156
rect 14283 85196 14325 85205
rect 14283 85156 14284 85196
rect 14324 85156 14325 85196
rect 14283 85147 14325 85156
rect 3051 85112 3093 85121
rect 3051 85072 3052 85112
rect 3092 85072 3093 85112
rect 3051 85063 3093 85072
rect 7467 85112 7509 85121
rect 7467 85072 7468 85112
rect 7508 85072 7509 85112
rect 7467 85063 7509 85072
rect 7707 85112 7749 85121
rect 7707 85072 7708 85112
rect 7748 85072 7749 85112
rect 7707 85063 7749 85072
rect 8427 85112 8469 85121
rect 8427 85072 8428 85112
rect 8468 85072 8469 85112
rect 8427 85063 8469 85072
rect 8619 85112 8661 85121
rect 8619 85072 8620 85112
rect 8660 85072 8661 85112
rect 8619 85063 8661 85072
rect 12843 85112 12885 85121
rect 12843 85072 12844 85112
rect 12884 85072 12885 85112
rect 12843 85063 12885 85072
rect 15627 85112 15669 85121
rect 15627 85072 15628 85112
rect 15668 85072 15669 85112
rect 15627 85063 15669 85072
rect 1419 85028 1461 85037
rect 1419 84988 1420 85028
rect 1460 84988 1461 85028
rect 1419 84979 1461 84988
rect 2659 85028 2717 85029
rect 2659 84988 2668 85028
rect 2708 84988 2717 85028
rect 2659 84987 2717 84988
rect 3435 85028 3477 85037
rect 3435 84988 3436 85028
rect 3476 84988 3477 85028
rect 3435 84979 3477 84988
rect 4675 85028 4733 85029
rect 4675 84988 4684 85028
rect 4724 84988 4733 85028
rect 4675 84987 4733 84988
rect 5259 85028 5301 85037
rect 5259 84988 5260 85028
rect 5300 84988 5301 85028
rect 5259 84979 5301 84988
rect 6499 85028 6557 85029
rect 6499 84988 6508 85028
rect 6548 84988 6557 85028
rect 6499 84987 6557 84988
rect 6874 85028 6932 85029
rect 6874 84988 6883 85028
rect 6923 84988 6932 85028
rect 6874 84987 6932 84988
rect 7851 85028 7893 85037
rect 7851 84988 7852 85028
rect 7892 84988 7893 85028
rect 7851 84979 7893 84988
rect 8043 85028 8085 85037
rect 8043 84988 8044 85028
rect 8084 84988 8085 85028
rect 8043 84979 8085 84988
rect 9003 85028 9045 85037
rect 9003 84988 9004 85028
rect 9044 84988 9045 85028
rect 9003 84979 9045 84988
rect 10243 85028 10301 85029
rect 10243 84988 10252 85028
rect 10292 84988 10301 85028
rect 10243 84987 10301 84988
rect 10635 85028 10677 85037
rect 10635 84988 10636 85028
rect 10676 84988 10677 85028
rect 10635 84979 10677 84988
rect 11875 85028 11933 85029
rect 11875 84988 11884 85028
rect 11924 84988 11933 85028
rect 11875 84987 11933 84988
rect 12346 85028 12404 85029
rect 12346 84988 12355 85028
rect 12395 84988 12404 85028
rect 12346 84987 12404 84988
rect 12459 85028 12501 85037
rect 12459 84988 12460 85028
rect 12500 84988 12501 85028
rect 12459 84979 12501 84988
rect 12939 85028 12981 85037
rect 12939 84988 12940 85028
rect 12980 84988 12981 85028
rect 12939 84979 12981 84988
rect 13411 85028 13469 85029
rect 13411 84988 13420 85028
rect 13460 84988 13469 85028
rect 13411 84987 13469 84988
rect 13899 85028 13957 85029
rect 13899 84988 13908 85028
rect 13948 84988 13957 85028
rect 13899 84987 13957 84988
rect 14283 85028 14325 85037
rect 14283 84988 14284 85028
rect 14324 84988 14325 85028
rect 14283 84979 14325 84988
rect 14571 85028 14613 85037
rect 14571 84988 14572 85028
rect 14612 84988 14613 85028
rect 14571 84979 14613 84988
rect 15130 85028 15188 85029
rect 15130 84988 15139 85028
rect 15179 84988 15188 85028
rect 15130 84987 15188 84988
rect 15243 85028 15285 85037
rect 15243 84988 15244 85028
rect 15284 84988 15285 85028
rect 15243 84979 15285 84988
rect 15723 85028 15765 85037
rect 15723 84988 15724 85028
rect 15764 84988 15765 85028
rect 15723 84979 15765 84988
rect 16195 85028 16253 85029
rect 16195 84988 16204 85028
rect 16244 84988 16253 85028
rect 16195 84987 16253 84988
rect 16714 85028 16772 85029
rect 16714 84988 16723 85028
rect 16763 84988 16772 85028
rect 16714 84987 16772 84988
rect 17067 85028 17109 85037
rect 17067 84988 17068 85028
rect 17108 84988 17109 85028
rect 17067 84979 17109 84988
rect 18307 85028 18365 85029
rect 18307 84988 18316 85028
rect 18356 84988 18365 85028
rect 18307 84987 18365 84988
rect 18699 85028 18741 85037
rect 18699 84988 18700 85028
rect 18740 84988 18741 85028
rect 18699 84979 18741 84988
rect 19939 85028 19997 85029
rect 19939 84988 19948 85028
rect 19988 84988 19997 85028
rect 19939 84987 19997 84988
rect 3291 84944 3333 84953
rect 3291 84904 3292 84944
rect 3332 84904 3333 84944
rect 3291 84895 3333 84904
rect 7083 84944 7125 84953
rect 7083 84904 7084 84944
rect 7124 84904 7125 84944
rect 7083 84895 7125 84904
rect 7193 84944 7235 84953
rect 7193 84904 7194 84944
rect 7234 84904 7235 84944
rect 7193 84895 7235 84904
rect 7947 84944 7989 84953
rect 7947 84904 7948 84944
rect 7988 84904 7989 84944
rect 7947 84895 7989 84904
rect 2859 84860 2901 84869
rect 2859 84820 2860 84860
rect 2900 84820 2901 84860
rect 2859 84811 2901 84820
rect 6699 84860 6741 84869
rect 6699 84820 6700 84860
rect 6740 84820 6741 84860
rect 6699 84811 6741 84820
rect 6970 84860 7028 84861
rect 6970 84820 6979 84860
rect 7019 84820 7028 84860
rect 6970 84819 7028 84820
rect 10443 84860 10485 84869
rect 10443 84820 10444 84860
rect 10484 84820 10485 84860
rect 10443 84811 10485 84820
rect 12075 84860 12117 84869
rect 12075 84820 12076 84860
rect 12116 84820 12117 84860
rect 12075 84811 12117 84820
rect 14091 84860 14133 84869
rect 14091 84820 14092 84860
rect 14132 84820 14133 84860
rect 14091 84811 14133 84820
rect 16875 84860 16917 84869
rect 16875 84820 16876 84860
rect 16916 84820 16917 84860
rect 16875 84811 16917 84820
rect 18507 84860 18549 84869
rect 18507 84820 18508 84860
rect 18548 84820 18549 84860
rect 18507 84811 18549 84820
rect 20139 84860 20181 84869
rect 20139 84820 20140 84860
rect 20180 84820 20181 84860
rect 20139 84811 20181 84820
rect 1152 84692 20452 84716
rect 1152 84652 4928 84692
rect 4968 84652 5010 84692
rect 5050 84652 5092 84692
rect 5132 84652 5174 84692
rect 5214 84652 5256 84692
rect 5296 84652 20048 84692
rect 20088 84652 20130 84692
rect 20170 84652 20212 84692
rect 20252 84652 20294 84692
rect 20334 84652 20376 84692
rect 20416 84652 20452 84692
rect 1152 84628 20452 84652
rect 4491 84524 4533 84533
rect 4491 84484 4492 84524
rect 4532 84484 4533 84524
rect 4491 84475 4533 84484
rect 7659 84524 7701 84533
rect 7659 84484 7660 84524
rect 7700 84484 7701 84524
rect 7659 84475 7701 84484
rect 8427 84524 8469 84533
rect 8427 84484 8428 84524
rect 8468 84484 8469 84524
rect 8427 84475 8469 84484
rect 9147 84524 9189 84533
rect 9147 84484 9148 84524
rect 9188 84484 9189 84524
rect 9147 84475 9189 84484
rect 12363 84524 12405 84533
rect 12363 84484 12364 84524
rect 12404 84484 12405 84524
rect 12363 84475 12405 84484
rect 12747 84524 12789 84533
rect 12747 84484 12748 84524
rect 12788 84484 12789 84524
rect 12747 84475 12789 84484
rect 14379 84524 14421 84533
rect 14379 84484 14380 84524
rect 14420 84484 14421 84524
rect 14379 84475 14421 84484
rect 14763 84524 14805 84533
rect 14763 84484 14764 84524
rect 14804 84484 14805 84524
rect 14763 84475 14805 84484
rect 16875 84524 16917 84533
rect 16875 84484 16876 84524
rect 16916 84484 16917 84524
rect 16875 84475 16917 84484
rect 19563 84524 19605 84533
rect 19563 84484 19564 84524
rect 19604 84484 19605 84524
rect 19563 84475 19605 84484
rect 5691 84440 5733 84449
rect 5691 84400 5692 84440
rect 5732 84400 5733 84440
rect 5691 84391 5733 84400
rect 13707 84440 13749 84449
rect 13707 84400 13708 84440
rect 13748 84400 13749 84440
rect 13707 84391 13749 84400
rect 14173 84440 14215 84449
rect 14173 84400 14174 84440
rect 14214 84400 14215 84440
rect 14173 84391 14215 84400
rect 14266 84440 14324 84441
rect 14266 84400 14275 84440
rect 14315 84400 14324 84440
rect 14266 84399 14324 84400
rect 2746 84356 2804 84357
rect 2746 84316 2755 84356
rect 2795 84316 2804 84356
rect 2746 84315 2804 84316
rect 2859 84356 2901 84365
rect 2859 84316 2860 84356
rect 2900 84316 2901 84356
rect 2859 84307 2901 84316
rect 3243 84356 3285 84365
rect 5914 84356 5972 84357
rect 3243 84316 3244 84356
rect 3284 84316 3285 84356
rect 3243 84307 3285 84316
rect 3819 84347 3861 84356
rect 3819 84307 3820 84347
rect 3860 84307 3861 84347
rect 3819 84298 3861 84307
rect 4299 84347 4341 84356
rect 4299 84307 4300 84347
rect 4340 84307 4341 84347
rect 5914 84316 5923 84356
rect 5963 84316 5972 84356
rect 5914 84315 5972 84316
rect 6027 84356 6069 84365
rect 6027 84316 6028 84356
rect 6068 84316 6069 84356
rect 6027 84307 6069 84316
rect 6411 84356 6453 84365
rect 7947 84356 7989 84365
rect 6411 84316 6412 84356
rect 6452 84316 6453 84356
rect 6411 84307 6453 84316
rect 6987 84347 7029 84356
rect 6987 84307 6988 84347
rect 7028 84307 7029 84347
rect 4299 84298 4341 84307
rect 6987 84298 7029 84307
rect 7467 84347 7509 84356
rect 7467 84307 7468 84347
rect 7508 84307 7509 84347
rect 7947 84316 7948 84356
rect 7988 84316 7989 84356
rect 7947 84307 7989 84316
rect 8178 84356 8220 84365
rect 8178 84316 8179 84356
rect 8219 84316 8220 84356
rect 8178 84307 8220 84316
rect 8332 84356 8374 84365
rect 8332 84316 8333 84356
rect 8373 84316 8374 84356
rect 8332 84307 8374 84316
rect 8523 84356 8565 84365
rect 8523 84316 8524 84356
rect 8564 84316 8565 84356
rect 8523 84307 8565 84316
rect 9291 84356 9333 84365
rect 10923 84356 10965 84365
rect 12843 84356 12885 84365
rect 9291 84316 9292 84356
rect 9332 84316 9333 84356
rect 9291 84307 9333 84316
rect 10539 84347 10581 84356
rect 10539 84307 10540 84347
rect 10580 84307 10581 84347
rect 10923 84316 10924 84356
rect 10964 84316 10965 84356
rect 10923 84307 10965 84316
rect 12171 84347 12213 84356
rect 12171 84307 12172 84347
rect 12212 84307 12213 84347
rect 12843 84316 12844 84356
rect 12884 84316 12885 84356
rect 12843 84307 12885 84316
rect 13072 84356 13130 84357
rect 13072 84316 13081 84356
rect 13121 84316 13130 84356
rect 13072 84315 13130 84316
rect 13323 84356 13365 84365
rect 13323 84316 13324 84356
rect 13364 84316 13365 84356
rect 13323 84307 13365 84316
rect 13594 84356 13652 84357
rect 13594 84316 13603 84356
rect 13643 84316 13652 84356
rect 14667 84356 14709 84365
rect 13594 84315 13652 84316
rect 14473 84331 14531 84332
rect 7467 84298 7509 84307
rect 10539 84298 10581 84307
rect 12171 84298 12213 84307
rect 14473 84291 14482 84331
rect 14522 84291 14531 84331
rect 14667 84316 14668 84356
rect 14708 84316 14709 84356
rect 14667 84307 14709 84316
rect 14859 84356 14901 84365
rect 14859 84316 14860 84356
rect 14900 84316 14901 84356
rect 14859 84307 14901 84316
rect 15130 84356 15188 84357
rect 15130 84316 15139 84356
rect 15179 84316 15188 84356
rect 15130 84315 15188 84316
rect 15243 84356 15285 84365
rect 15243 84316 15244 84356
rect 15284 84316 15285 84356
rect 15243 84307 15285 84316
rect 15627 84356 15669 84365
rect 17818 84356 17876 84357
rect 15627 84316 15628 84356
rect 15668 84316 15669 84356
rect 15627 84307 15669 84316
rect 16203 84347 16245 84356
rect 16203 84307 16204 84347
rect 16244 84307 16245 84347
rect 16203 84298 16245 84307
rect 16683 84347 16725 84356
rect 16683 84307 16684 84347
rect 16724 84307 16725 84347
rect 17818 84316 17827 84356
rect 17867 84316 17876 84356
rect 17818 84315 17876 84316
rect 17931 84356 17973 84365
rect 17931 84316 17932 84356
rect 17972 84316 17973 84356
rect 17931 84307 17973 84316
rect 18315 84356 18357 84365
rect 18315 84316 18316 84356
rect 18356 84316 18357 84356
rect 18315 84307 18357 84316
rect 18891 84347 18933 84356
rect 18891 84307 18892 84347
rect 18932 84307 18933 84347
rect 16683 84298 16725 84307
rect 18891 84298 18933 84307
rect 19371 84347 19413 84356
rect 19371 84307 19372 84347
rect 19412 84307 19413 84347
rect 19371 84298 19413 84307
rect 14473 84290 14531 84291
rect 1227 84272 1269 84281
rect 1227 84232 1228 84272
rect 1268 84232 1269 84272
rect 1227 84223 1269 84232
rect 1611 84272 1653 84281
rect 1611 84232 1612 84272
rect 1652 84232 1653 84272
rect 1611 84223 1653 84232
rect 1995 84272 2037 84281
rect 1995 84232 1996 84272
rect 2036 84232 2037 84272
rect 1995 84223 2037 84232
rect 3339 84272 3381 84281
rect 3339 84232 3340 84272
rect 3380 84232 3381 84272
rect 3339 84223 3381 84232
rect 4683 84272 4725 84281
rect 4683 84232 4684 84272
rect 4724 84232 4725 84272
rect 4683 84223 4725 84232
rect 5067 84272 5109 84281
rect 5067 84232 5068 84272
rect 5108 84232 5109 84272
rect 5067 84223 5109 84232
rect 5451 84272 5493 84281
rect 5451 84232 5452 84272
rect 5492 84232 5493 84272
rect 5451 84223 5493 84232
rect 6507 84272 6549 84281
rect 6507 84232 6508 84272
rect 6548 84232 6549 84272
rect 6507 84223 6549 84232
rect 7851 84272 7893 84281
rect 7851 84232 7852 84272
rect 7892 84232 7893 84272
rect 7851 84223 7893 84232
rect 8066 84272 8108 84281
rect 8066 84232 8067 84272
rect 8107 84232 8108 84272
rect 8066 84223 8108 84232
rect 8907 84272 8949 84281
rect 15723 84272 15765 84281
rect 8907 84232 8908 84272
rect 8948 84232 8949 84272
rect 8907 84223 8949 84232
rect 12978 84263 13024 84272
rect 12978 84223 12979 84263
rect 13019 84223 13024 84263
rect 15723 84232 15724 84272
rect 15764 84232 15765 84272
rect 15723 84223 15765 84232
rect 17067 84272 17109 84281
rect 17067 84232 17068 84272
rect 17108 84232 17109 84272
rect 17067 84223 17109 84232
rect 18411 84272 18453 84281
rect 18411 84232 18412 84272
rect 18452 84232 18453 84272
rect 18411 84223 18453 84232
rect 19755 84272 19797 84281
rect 19755 84232 19756 84272
rect 19796 84232 19797 84272
rect 19755 84223 19797 84232
rect 20139 84272 20181 84281
rect 20139 84232 20140 84272
rect 20180 84232 20181 84272
rect 20139 84223 20181 84232
rect 12978 84214 13024 84223
rect 5307 84188 5349 84197
rect 5307 84148 5308 84188
rect 5348 84148 5349 84188
rect 5307 84139 5349 84148
rect 13995 84188 14037 84197
rect 13995 84148 13996 84188
rect 14036 84148 14037 84188
rect 13995 84139 14037 84148
rect 1467 84104 1509 84113
rect 1467 84064 1468 84104
rect 1508 84064 1509 84104
rect 1467 84055 1509 84064
rect 1851 84104 1893 84113
rect 1851 84064 1852 84104
rect 1892 84064 1893 84104
rect 1851 84055 1893 84064
rect 2235 84104 2277 84113
rect 2235 84064 2236 84104
rect 2276 84064 2277 84104
rect 2235 84055 2277 84064
rect 4923 84104 4965 84113
rect 4923 84064 4924 84104
rect 4964 84064 4965 84104
rect 4923 84055 4965 84064
rect 9147 84104 9189 84113
rect 9147 84064 9148 84104
rect 9188 84064 9189 84104
rect 9147 84055 9189 84064
rect 10731 84104 10773 84113
rect 10731 84064 10732 84104
rect 10772 84064 10773 84104
rect 10731 84055 10773 84064
rect 17307 84104 17349 84113
rect 17307 84064 17308 84104
rect 17348 84064 17349 84104
rect 17307 84055 17349 84064
rect 19995 84104 20037 84113
rect 19995 84064 19996 84104
rect 20036 84064 20037 84104
rect 19995 84055 20037 84064
rect 20379 84104 20421 84113
rect 20379 84064 20380 84104
rect 20420 84064 20421 84104
rect 20379 84055 20421 84064
rect 1152 83936 20448 83960
rect 1152 83896 3688 83936
rect 3728 83896 3770 83936
rect 3810 83896 3852 83936
rect 3892 83896 3934 83936
rect 3974 83896 4016 83936
rect 4056 83896 18808 83936
rect 18848 83896 18890 83936
rect 18930 83896 18972 83936
rect 19012 83896 19054 83936
rect 19094 83896 19136 83936
rect 19176 83896 20448 83936
rect 1152 83872 20448 83896
rect 5307 83768 5349 83777
rect 5307 83728 5308 83768
rect 5348 83728 5349 83768
rect 5307 83719 5349 83728
rect 5883 83768 5925 83777
rect 5883 83728 5884 83768
rect 5924 83728 5925 83768
rect 5883 83719 5925 83728
rect 7659 83768 7701 83777
rect 7659 83728 7660 83768
rect 7700 83728 7701 83768
rect 7659 83719 7701 83728
rect 9339 83768 9381 83777
rect 9339 83728 9340 83768
rect 9380 83728 9381 83768
rect 9339 83719 9381 83728
rect 13066 83768 13124 83769
rect 13066 83728 13075 83768
rect 13115 83728 13124 83768
rect 13066 83727 13124 83728
rect 14811 83768 14853 83777
rect 14811 83728 14812 83768
rect 14852 83728 14853 83768
rect 14811 83719 14853 83728
rect 19594 83768 19652 83769
rect 19594 83728 19603 83768
rect 19643 83728 19652 83768
rect 19594 83727 19652 83728
rect 7467 83684 7509 83693
rect 7467 83644 7468 83684
rect 7508 83644 7509 83684
rect 7467 83635 7509 83644
rect 11019 83684 11061 83693
rect 11019 83644 11020 83684
rect 11060 83644 11061 83684
rect 11019 83635 11061 83644
rect 19755 83684 19797 83693
rect 19755 83644 19756 83684
rect 19796 83644 19797 83684
rect 19755 83635 19797 83644
rect 3915 83600 3957 83609
rect 3915 83560 3916 83600
rect 3956 83560 3957 83600
rect 3915 83551 3957 83560
rect 5547 83600 5589 83609
rect 5547 83560 5548 83600
rect 5588 83560 5589 83600
rect 5547 83551 5589 83560
rect 8907 83600 8949 83609
rect 8907 83560 8908 83600
rect 8948 83560 8949 83600
rect 8907 83551 8949 83560
rect 9099 83600 9141 83609
rect 9099 83560 9100 83600
rect 9140 83560 9141 83600
rect 9099 83551 9141 83560
rect 11787 83600 11829 83609
rect 11787 83560 11788 83600
rect 11828 83560 11829 83600
rect 11787 83551 11829 83560
rect 13611 83600 13653 83609
rect 13611 83560 13612 83600
rect 13652 83560 13653 83600
rect 13611 83551 13653 83560
rect 13851 83600 13893 83609
rect 13851 83560 13852 83600
rect 13892 83560 13893 83600
rect 13851 83551 13893 83560
rect 14187 83600 14229 83609
rect 14187 83560 14188 83600
rect 14228 83560 14229 83600
rect 14187 83551 14229 83560
rect 14523 83600 14565 83609
rect 14523 83560 14524 83600
rect 14564 83560 14565 83600
rect 14523 83551 14565 83560
rect 15675 83600 15717 83609
rect 15675 83560 15676 83600
rect 15716 83560 15717 83600
rect 15675 83551 15717 83560
rect 15915 83600 15957 83609
rect 15915 83560 15916 83600
rect 15956 83560 15957 83600
rect 15915 83551 15957 83560
rect 18315 83600 18357 83609
rect 18315 83560 18316 83600
rect 18356 83560 18357 83600
rect 18315 83551 18357 83560
rect 20139 83600 20181 83609
rect 20139 83560 20140 83600
rect 20180 83560 20181 83600
rect 20139 83551 20181 83560
rect 20379 83600 20421 83609
rect 20379 83560 20380 83600
rect 20420 83560 20421 83600
rect 20379 83551 20421 83560
rect 1515 83516 1557 83525
rect 1515 83476 1516 83516
rect 1556 83476 1557 83516
rect 1515 83467 1557 83476
rect 2755 83516 2813 83517
rect 2755 83476 2764 83516
rect 2804 83476 2813 83516
rect 2755 83475 2813 83476
rect 3418 83516 3476 83517
rect 3418 83476 3427 83516
rect 3467 83476 3476 83516
rect 3418 83475 3476 83476
rect 3531 83516 3573 83525
rect 3531 83476 3532 83516
rect 3572 83476 3573 83516
rect 3531 83467 3573 83476
rect 4011 83516 4053 83525
rect 4011 83476 4012 83516
rect 4052 83476 4053 83516
rect 4011 83467 4053 83476
rect 4483 83516 4541 83517
rect 4483 83476 4492 83516
rect 4532 83476 4541 83516
rect 4483 83475 4541 83476
rect 4971 83516 5029 83517
rect 4971 83476 4980 83516
rect 5020 83476 5029 83516
rect 4971 83475 5029 83476
rect 5739 83516 5781 83525
rect 5739 83476 5740 83516
rect 5780 83476 5781 83516
rect 5739 83467 5781 83476
rect 6027 83516 6069 83525
rect 6027 83476 6028 83516
rect 6068 83476 6069 83516
rect 6027 83467 6069 83476
rect 7267 83516 7325 83517
rect 8331 83516 8373 83525
rect 7267 83476 7276 83516
rect 7316 83476 7325 83516
rect 7267 83475 7325 83476
rect 8043 83507 8085 83516
rect 8043 83467 8044 83507
rect 8084 83467 8085 83507
rect 8331 83476 8332 83516
rect 8372 83476 8373 83516
rect 8331 83467 8373 83476
rect 8566 83516 8608 83525
rect 8566 83476 8567 83516
rect 8607 83476 8608 83516
rect 8566 83467 8608 83476
rect 8698 83516 8756 83517
rect 8698 83476 8707 83516
rect 8747 83476 8756 83516
rect 8698 83475 8756 83476
rect 8811 83516 8853 83525
rect 8811 83476 8812 83516
rect 8852 83476 8853 83516
rect 8811 83467 8853 83476
rect 9579 83516 9621 83525
rect 9579 83476 9580 83516
rect 9620 83476 9621 83516
rect 9579 83467 9621 83476
rect 10819 83516 10877 83517
rect 10819 83476 10828 83516
rect 10868 83476 10877 83516
rect 10819 83475 10877 83476
rect 11277 83516 11319 83525
rect 11277 83476 11278 83516
rect 11318 83476 11319 83516
rect 11277 83467 11319 83476
rect 11403 83516 11445 83525
rect 11403 83476 11404 83516
rect 11444 83476 11445 83516
rect 11403 83467 11445 83476
rect 11883 83516 11925 83525
rect 11883 83476 11884 83516
rect 11924 83476 11925 83516
rect 11883 83467 11925 83476
rect 12355 83516 12413 83517
rect 12355 83476 12364 83516
rect 12404 83476 12413 83516
rect 12355 83475 12413 83476
rect 12843 83516 12901 83517
rect 12843 83476 12852 83516
rect 12892 83476 12901 83516
rect 12843 83475 12901 83476
rect 14938 83516 14996 83517
rect 14938 83476 14947 83516
rect 14987 83476 14996 83516
rect 14938 83475 14996 83476
rect 15257 83516 15299 83525
rect 15257 83476 15258 83516
rect 15298 83476 15299 83516
rect 15257 83467 15299 83476
rect 16107 83516 16149 83525
rect 16107 83476 16108 83516
rect 16148 83476 16149 83516
rect 16107 83467 16149 83476
rect 17347 83516 17405 83517
rect 17347 83476 17356 83516
rect 17396 83476 17405 83516
rect 17347 83475 17405 83476
rect 17818 83516 17876 83517
rect 17818 83476 17827 83516
rect 17867 83476 17876 83516
rect 17818 83475 17876 83476
rect 17931 83516 17973 83525
rect 17931 83476 17932 83516
rect 17972 83476 17973 83516
rect 17931 83467 17973 83476
rect 18411 83516 18453 83525
rect 18411 83476 18412 83516
rect 18452 83476 18453 83516
rect 18411 83467 18453 83476
rect 18883 83516 18941 83517
rect 18883 83476 18892 83516
rect 18932 83476 18941 83516
rect 18883 83475 18941 83476
rect 19402 83516 19460 83517
rect 19402 83476 19411 83516
rect 19451 83476 19460 83516
rect 19402 83475 19460 83476
rect 19755 83516 19797 83525
rect 19755 83476 19756 83516
rect 19796 83476 19797 83516
rect 19755 83467 19797 83476
rect 19947 83516 19989 83525
rect 19947 83476 19948 83516
rect 19988 83476 19989 83516
rect 19947 83467 19989 83476
rect 8043 83458 8085 83467
rect 7947 83432 7989 83441
rect 7947 83392 7948 83432
rect 7988 83392 7989 83432
rect 7947 83383 7989 83392
rect 13947 83432 13989 83441
rect 13947 83392 13948 83432
rect 13988 83392 13989 83432
rect 13947 83383 13989 83392
rect 15051 83432 15093 83441
rect 15051 83392 15052 83432
rect 15092 83392 15093 83432
rect 15051 83383 15093 83392
rect 17547 83432 17589 83441
rect 17547 83392 17548 83432
rect 17588 83392 17589 83432
rect 17547 83383 17589 83392
rect 2955 83348 2997 83357
rect 2955 83308 2956 83348
rect 2996 83308 2997 83348
rect 2955 83299 2997 83308
rect 5163 83348 5205 83357
rect 5163 83308 5164 83348
rect 5204 83308 5205 83348
rect 5163 83299 5205 83308
rect 15147 83348 15189 83357
rect 15147 83308 15148 83348
rect 15188 83308 15189 83348
rect 15147 83299 15189 83308
rect 1152 83180 20452 83204
rect 1152 83140 4928 83180
rect 4968 83140 5010 83180
rect 5050 83140 5092 83180
rect 5132 83140 5174 83180
rect 5214 83140 5256 83180
rect 5296 83140 20048 83180
rect 20088 83140 20130 83180
rect 20170 83140 20212 83180
rect 20252 83140 20294 83180
rect 20334 83140 20376 83180
rect 20416 83140 20452 83180
rect 1152 83116 20452 83140
rect 4971 83012 5013 83021
rect 4971 82972 4972 83012
rect 5012 82972 5013 83012
rect 4971 82963 5013 82972
rect 8427 83012 8469 83021
rect 8427 82972 8428 83012
rect 8468 82972 8469 83012
rect 8427 82963 8469 82972
rect 13131 83012 13173 83021
rect 13131 82972 13132 83012
rect 13172 82972 13173 83012
rect 13131 82963 13173 82972
rect 14475 83012 14517 83021
rect 14475 82972 14476 83012
rect 14516 82972 14517 83012
rect 14475 82963 14517 82972
rect 14907 83012 14949 83021
rect 14907 82972 14908 83012
rect 14948 82972 14949 83012
rect 14907 82963 14949 82972
rect 5163 82928 5205 82937
rect 5163 82888 5164 82928
rect 5204 82888 5205 82928
rect 5163 82879 5205 82888
rect 16011 82928 16053 82937
rect 16011 82888 16012 82928
rect 16052 82888 16053 82928
rect 16011 82879 16053 82888
rect 1515 82844 1557 82853
rect 3226 82844 3284 82845
rect 1515 82804 1516 82844
rect 1556 82804 1557 82844
rect 1515 82795 1557 82804
rect 2763 82835 2805 82844
rect 2763 82795 2764 82835
rect 2804 82795 2805 82835
rect 3226 82804 3235 82844
rect 3275 82804 3284 82844
rect 3226 82803 3284 82804
rect 3339 82844 3381 82853
rect 3339 82804 3340 82844
rect 3380 82804 3381 82844
rect 3339 82795 3381 82804
rect 3723 82844 3765 82853
rect 6603 82844 6645 82853
rect 3723 82804 3724 82844
rect 3764 82804 3765 82844
rect 3723 82795 3765 82804
rect 4299 82835 4341 82844
rect 4299 82795 4300 82835
rect 4340 82795 4341 82835
rect 2763 82786 2805 82795
rect 4299 82786 4341 82795
rect 4779 82835 4821 82844
rect 4779 82795 4780 82835
rect 4820 82795 4821 82835
rect 4779 82786 4821 82795
rect 5355 82835 5397 82844
rect 5355 82795 5356 82835
rect 5396 82795 5397 82835
rect 6603 82804 6604 82844
rect 6644 82804 6645 82844
rect 6603 82795 6645 82804
rect 6987 82844 7029 82853
rect 8619 82844 8661 82853
rect 11386 82844 11444 82845
rect 6987 82804 6988 82844
rect 7028 82804 7029 82844
rect 6987 82795 7029 82804
rect 8235 82835 8277 82844
rect 8235 82795 8236 82835
rect 8276 82795 8277 82835
rect 8619 82804 8620 82844
rect 8660 82804 8661 82844
rect 8619 82795 8661 82804
rect 9867 82835 9909 82844
rect 9867 82795 9868 82835
rect 9908 82795 9909 82835
rect 11386 82804 11395 82844
rect 11435 82804 11444 82844
rect 11386 82803 11444 82804
rect 11499 82844 11541 82853
rect 11499 82804 11500 82844
rect 11540 82804 11541 82844
rect 11499 82795 11541 82804
rect 11883 82844 11925 82853
rect 14571 82844 14613 82853
rect 11883 82804 11884 82844
rect 11924 82804 11925 82844
rect 11883 82795 11925 82804
rect 12459 82835 12501 82844
rect 12459 82795 12460 82835
rect 12500 82795 12501 82835
rect 5355 82786 5397 82795
rect 8235 82786 8277 82795
rect 9867 82786 9909 82795
rect 12459 82786 12501 82795
rect 12939 82835 12981 82844
rect 12939 82795 12940 82835
rect 12980 82795 12981 82835
rect 14571 82804 14572 82844
rect 14612 82804 14613 82844
rect 14571 82795 14613 82804
rect 14800 82844 14858 82845
rect 14800 82804 14809 82844
rect 14849 82804 14858 82844
rect 14800 82803 14858 82804
rect 15243 82844 15285 82853
rect 15243 82804 15244 82844
rect 15284 82804 15285 82844
rect 15243 82795 15285 82804
rect 15344 82844 15402 82845
rect 15344 82804 15353 82844
rect 15393 82804 15402 82844
rect 15344 82803 15402 82804
rect 15627 82844 15669 82853
rect 15627 82804 15628 82844
rect 15668 82804 15669 82844
rect 15627 82795 15669 82804
rect 15915 82844 15957 82853
rect 15915 82804 15916 82844
rect 15956 82804 15957 82844
rect 15915 82795 15957 82804
rect 16107 82844 16149 82853
rect 16107 82804 16108 82844
rect 16148 82804 16149 82844
rect 16107 82795 16149 82804
rect 16299 82844 16341 82853
rect 16299 82804 16300 82844
rect 16340 82804 16341 82844
rect 16299 82795 16341 82804
rect 16491 82844 16533 82853
rect 16491 82804 16492 82844
rect 16532 82804 16533 82844
rect 16491 82795 16533 82804
rect 16875 82844 16917 82853
rect 19947 82844 19989 82853
rect 16875 82804 16876 82844
rect 16916 82804 16917 82844
rect 16875 82795 16917 82804
rect 18123 82835 18165 82844
rect 18123 82795 18124 82835
rect 18164 82795 18165 82835
rect 12939 82786 12981 82795
rect 18123 82786 18165 82795
rect 18699 82835 18741 82844
rect 18699 82795 18700 82835
rect 18740 82795 18741 82835
rect 19947 82804 19948 82844
rect 19988 82804 19989 82844
rect 19947 82795 19989 82804
rect 18699 82786 18741 82795
rect 3850 82760 3908 82761
rect 3850 82720 3859 82760
rect 3899 82720 3908 82760
rect 3850 82719 3908 82720
rect 11979 82760 12021 82769
rect 11979 82720 11980 82760
rect 12020 82720 12021 82760
rect 11979 82711 12021 82720
rect 13419 82760 13461 82769
rect 13419 82720 13420 82760
rect 13460 82720 13461 82760
rect 13419 82711 13461 82720
rect 14091 82760 14133 82769
rect 14091 82720 14092 82760
rect 14132 82720 14133 82760
rect 14091 82711 14133 82720
rect 14690 82760 14732 82769
rect 14690 82720 14691 82760
rect 14731 82720 14732 82760
rect 14690 82711 14732 82720
rect 20139 82760 20181 82769
rect 20139 82720 20140 82760
rect 20180 82720 20181 82760
rect 20139 82711 20181 82720
rect 13659 82676 13701 82685
rect 13659 82636 13660 82676
rect 13700 82636 13701 82676
rect 13659 82627 13701 82636
rect 16299 82676 16341 82685
rect 16299 82636 16300 82676
rect 16340 82636 16341 82676
rect 16299 82627 16341 82636
rect 20379 82676 20421 82685
rect 20379 82636 20380 82676
rect 20420 82636 20421 82676
rect 20379 82627 20421 82636
rect 2955 82592 2997 82601
rect 2955 82552 2956 82592
rect 2996 82552 2997 82592
rect 2955 82543 2997 82552
rect 10059 82592 10101 82601
rect 10059 82552 10060 82592
rect 10100 82552 10101 82592
rect 10059 82543 10101 82552
rect 14331 82592 14373 82601
rect 14331 82552 14332 82592
rect 14372 82552 14373 82592
rect 14331 82543 14373 82552
rect 18315 82592 18357 82601
rect 18315 82552 18316 82592
rect 18356 82552 18357 82592
rect 18315 82543 18357 82552
rect 18507 82592 18549 82601
rect 18507 82552 18508 82592
rect 18548 82552 18549 82592
rect 18507 82543 18549 82552
rect 1152 82424 20448 82448
rect 1152 82384 3688 82424
rect 3728 82384 3770 82424
rect 3810 82384 3852 82424
rect 3892 82384 3934 82424
rect 3974 82384 4016 82424
rect 4056 82384 18808 82424
rect 18848 82384 18890 82424
rect 18930 82384 18972 82424
rect 19012 82384 19054 82424
rect 19094 82384 19136 82424
rect 19176 82384 20448 82424
rect 1152 82360 20448 82384
rect 7275 82256 7317 82265
rect 7275 82216 7276 82256
rect 7316 82216 7317 82256
rect 7275 82207 7317 82216
rect 13659 82256 13701 82265
rect 13659 82216 13660 82256
rect 13700 82216 13701 82256
rect 13659 82207 13701 82216
rect 6603 82172 6645 82181
rect 6603 82132 6604 82172
rect 6644 82132 6645 82172
rect 6603 82123 6645 82132
rect 3723 82088 3765 82097
rect 3723 82048 3724 82088
rect 3764 82048 3765 82088
rect 3723 82039 3765 82048
rect 8427 82088 8469 82097
rect 8427 82048 8428 82088
rect 8468 82048 8469 82088
rect 8427 82039 8469 82048
rect 8619 82088 8661 82097
rect 8619 82048 8620 82088
rect 8660 82048 8661 82088
rect 8619 82039 8661 82048
rect 11691 82088 11733 82097
rect 11691 82048 11692 82088
rect 11732 82048 11733 82088
rect 11691 82039 11733 82048
rect 13419 82088 13461 82097
rect 13419 82048 13420 82088
rect 13460 82048 13461 82088
rect 13419 82039 13461 82048
rect 14379 82088 14421 82097
rect 14379 82048 14380 82088
rect 14420 82048 14421 82088
rect 14379 82039 14421 82048
rect 16251 82088 16293 82097
rect 16251 82048 16252 82088
rect 16292 82048 16293 82088
rect 16251 82039 16293 82048
rect 18891 82088 18933 82097
rect 18891 82048 18892 82088
rect 18932 82048 18933 82088
rect 18891 82039 18933 82048
rect 1515 82004 1557 82013
rect 1515 81964 1516 82004
rect 1556 81964 1557 82004
rect 1515 81955 1557 81964
rect 2755 82004 2813 82005
rect 2755 81964 2764 82004
rect 2804 81964 2813 82004
rect 2755 81963 2813 81964
rect 3226 82004 3284 82005
rect 3226 81964 3235 82004
rect 3275 81964 3284 82004
rect 3226 81963 3284 81964
rect 3339 82004 3381 82013
rect 3339 81964 3340 82004
rect 3380 81964 3381 82004
rect 3339 81955 3381 81964
rect 3819 82004 3861 82013
rect 3819 81964 3820 82004
rect 3860 81964 3861 82004
rect 3819 81955 3861 81964
rect 4291 82004 4349 82005
rect 4291 81964 4300 82004
rect 4340 81964 4349 82004
rect 4291 81963 4349 81964
rect 4779 82004 4837 82005
rect 4779 81964 4788 82004
rect 4828 81964 4837 82004
rect 4779 81963 4837 81964
rect 5163 82004 5205 82013
rect 5163 81964 5164 82004
rect 5204 81964 5205 82004
rect 5163 81955 5205 81964
rect 6403 82004 6461 82005
rect 6403 81964 6412 82004
rect 6452 81964 6461 82004
rect 6403 81963 6461 81964
rect 6742 82004 6784 82013
rect 6742 81964 6743 82004
rect 6783 81964 6784 82004
rect 6742 81955 6784 81964
rect 6874 82004 6932 82005
rect 6874 81964 6883 82004
rect 6923 81964 6932 82004
rect 6874 81963 6932 81964
rect 6987 82004 7029 82013
rect 6987 81964 6988 82004
rect 7028 81964 7029 82004
rect 6987 81955 7029 81964
rect 7275 82004 7317 82013
rect 7275 81964 7276 82004
rect 7316 81964 7317 82004
rect 7275 81955 7317 81964
rect 7563 82004 7605 82013
rect 7563 81964 7564 82004
rect 7604 81964 7605 82004
rect 7563 81955 7605 81964
rect 7755 82004 7797 82013
rect 7755 81964 7756 82004
rect 7796 81964 7797 82004
rect 7755 81955 7797 81964
rect 7930 82004 7988 82005
rect 7930 81964 7939 82004
rect 7979 81964 7988 82004
rect 7930 81963 7988 81964
rect 9099 82004 9141 82013
rect 9099 81964 9100 82004
rect 9140 81964 9141 82004
rect 9099 81955 9141 81964
rect 9291 82004 9333 82013
rect 9291 81964 9292 82004
rect 9332 81964 9333 82004
rect 9291 81955 9333 81964
rect 10531 82004 10589 82005
rect 10531 81964 10540 82004
rect 10580 81964 10589 82004
rect 10531 81963 10589 81964
rect 11194 82004 11252 82005
rect 11194 81964 11203 82004
rect 11243 81964 11252 82004
rect 11194 81963 11252 81964
rect 11307 82004 11349 82013
rect 11307 81964 11308 82004
rect 11348 81964 11349 82004
rect 11307 81955 11349 81964
rect 11787 82004 11829 82013
rect 11787 81964 11788 82004
rect 11828 81964 11829 82004
rect 11787 81955 11829 81964
rect 12259 82004 12317 82005
rect 12259 81964 12268 82004
rect 12308 81964 12317 82004
rect 12259 81963 12317 81964
rect 12747 82004 12805 82005
rect 12747 81964 12756 82004
rect 12796 81964 12805 82004
rect 12747 81963 12805 81964
rect 13882 82004 13940 82005
rect 13882 81964 13891 82004
rect 13931 81964 13940 82004
rect 13882 81963 13940 81964
rect 13995 82004 14037 82013
rect 13995 81964 13996 82004
rect 14036 81964 14037 82004
rect 13995 81955 14037 81964
rect 14475 82004 14517 82013
rect 14475 81964 14476 82004
rect 14516 81964 14517 82004
rect 14475 81955 14517 81964
rect 14947 82004 15005 82005
rect 14947 81964 14956 82004
rect 14996 81964 15005 82004
rect 14947 81963 15005 81964
rect 15435 82004 15493 82005
rect 15435 81964 15444 82004
rect 15484 81964 15493 82004
rect 15435 81963 15493 81964
rect 15802 82004 15860 82005
rect 15802 81964 15811 82004
rect 15851 81964 15860 82004
rect 15802 81963 15860 81964
rect 16107 82004 16149 82013
rect 16107 81964 16108 82004
rect 16148 81964 16149 82004
rect 16107 81955 16149 81964
rect 16395 82004 16437 82013
rect 16395 81964 16396 82004
rect 16436 81964 16437 82004
rect 16395 81955 16437 81964
rect 16587 82004 16629 82013
rect 16587 81964 16588 82004
rect 16628 81964 16629 82004
rect 16587 81955 16629 81964
rect 17827 82004 17885 82005
rect 17827 81964 17836 82004
rect 17876 81964 17885 82004
rect 17827 81963 17885 81964
rect 18381 82004 18423 82013
rect 18381 81964 18382 82004
rect 18422 81964 18423 82004
rect 18381 81955 18423 81964
rect 18512 82004 18554 82013
rect 18512 81964 18513 82004
rect 18553 81964 18554 82004
rect 18512 81955 18554 81964
rect 18987 82004 19029 82013
rect 18987 81964 18988 82004
rect 19028 81964 19029 82004
rect 18987 81955 19029 81964
rect 19459 82004 19517 82005
rect 19459 81964 19468 82004
rect 19508 81964 19517 82004
rect 19459 81963 19517 81964
rect 19947 82004 20005 82005
rect 19947 81964 19956 82004
rect 19996 81964 20005 82004
rect 19947 81963 20005 81964
rect 7851 81920 7893 81929
rect 7851 81880 7852 81920
rect 7892 81880 7893 81920
rect 7851 81871 7893 81880
rect 8859 81920 8901 81929
rect 8859 81880 8860 81920
rect 8900 81880 8901 81920
rect 8859 81871 8901 81880
rect 10731 81920 10773 81929
rect 10731 81880 10732 81920
rect 10772 81880 10773 81920
rect 10731 81871 10773 81880
rect 16011 81920 16053 81929
rect 16011 81880 16012 81920
rect 16052 81880 16053 81920
rect 16011 81871 16053 81880
rect 2955 81836 2997 81845
rect 2955 81796 2956 81836
rect 2996 81796 2997 81836
rect 2955 81787 2997 81796
rect 4971 81836 5013 81845
rect 4971 81796 4972 81836
rect 5012 81796 5013 81836
rect 4971 81787 5013 81796
rect 7066 81836 7124 81837
rect 7066 81796 7075 81836
rect 7115 81796 7124 81836
rect 7066 81795 7124 81796
rect 8187 81836 8229 81845
rect 8187 81796 8188 81836
rect 8228 81796 8229 81836
rect 8187 81787 8229 81796
rect 8955 81836 8997 81845
rect 8955 81796 8956 81836
rect 8996 81796 8997 81836
rect 8955 81787 8997 81796
rect 12939 81836 12981 81845
rect 12939 81796 12940 81836
rect 12980 81796 12981 81836
rect 12939 81787 12981 81796
rect 13659 81836 13701 81845
rect 13659 81796 13660 81836
rect 13700 81796 13701 81836
rect 13659 81787 13701 81796
rect 15627 81836 15669 81845
rect 15627 81796 15628 81836
rect 15668 81796 15669 81836
rect 15627 81787 15669 81796
rect 18027 81836 18069 81845
rect 18027 81796 18028 81836
rect 18068 81796 18069 81836
rect 18027 81787 18069 81796
rect 20139 81836 20181 81845
rect 20139 81796 20140 81836
rect 20180 81796 20181 81836
rect 20139 81787 20181 81796
rect 1152 81668 20452 81692
rect 1152 81628 4928 81668
rect 4968 81628 5010 81668
rect 5050 81628 5092 81668
rect 5132 81628 5174 81668
rect 5214 81628 5256 81668
rect 5296 81628 20048 81668
rect 20088 81628 20130 81668
rect 20170 81628 20212 81668
rect 20252 81628 20294 81668
rect 20334 81628 20376 81668
rect 20416 81628 20452 81668
rect 1152 81604 20452 81628
rect 4635 81500 4677 81509
rect 4635 81460 4636 81500
rect 4676 81460 4677 81500
rect 4635 81451 4677 81460
rect 6603 81500 6645 81509
rect 6603 81460 6604 81500
rect 6644 81460 6645 81500
rect 6603 81451 6645 81460
rect 7834 81500 7892 81501
rect 7834 81460 7843 81500
rect 7883 81460 7892 81500
rect 7834 81459 7892 81460
rect 8859 81500 8901 81509
rect 8859 81460 8860 81500
rect 8900 81460 8901 81500
rect 8859 81451 8901 81460
rect 10971 81500 11013 81509
rect 10971 81460 10972 81500
rect 11012 81460 11013 81500
rect 10971 81451 11013 81460
rect 13035 81500 13077 81509
rect 13035 81460 13036 81500
rect 13076 81460 13077 81500
rect 13035 81451 13077 81460
rect 17050 81500 17108 81501
rect 17050 81460 17059 81500
rect 17099 81460 17108 81500
rect 17050 81459 17108 81460
rect 17499 81500 17541 81509
rect 17499 81460 17500 81500
rect 17540 81460 17541 81500
rect 17499 81451 17541 81460
rect 20139 81500 20181 81509
rect 20139 81460 20140 81500
rect 20180 81460 20181 81500
rect 20139 81451 20181 81460
rect 7275 81416 7317 81425
rect 7275 81376 7276 81416
rect 7316 81376 7317 81416
rect 7275 81367 7317 81376
rect 7947 81416 7989 81425
rect 7947 81376 7948 81416
rect 7988 81376 7989 81416
rect 7947 81367 7989 81376
rect 10539 81416 10581 81425
rect 10539 81376 10540 81416
rect 10580 81376 10581 81416
rect 10539 81367 10581 81376
rect 14955 81416 14997 81425
rect 14955 81376 14956 81416
rect 14996 81376 14997 81416
rect 14955 81367 14997 81376
rect 1611 81332 1653 81341
rect 4858 81332 4916 81333
rect 1611 81292 1612 81332
rect 1652 81292 1653 81332
rect 1611 81283 1653 81292
rect 2859 81323 2901 81332
rect 2859 81283 2860 81323
rect 2900 81283 2901 81323
rect 4858 81292 4867 81332
rect 4907 81292 4916 81332
rect 4858 81291 4916 81292
rect 4971 81332 5013 81341
rect 4971 81292 4972 81332
rect 5012 81292 5013 81332
rect 4971 81283 5013 81292
rect 5355 81332 5397 81341
rect 6891 81332 6933 81341
rect 5355 81292 5356 81332
rect 5396 81292 5397 81332
rect 5355 81283 5397 81292
rect 5931 81323 5973 81332
rect 5931 81283 5932 81323
rect 5972 81283 5973 81323
rect 2859 81274 2901 81283
rect 5931 81274 5973 81283
rect 6411 81323 6453 81332
rect 6411 81283 6412 81323
rect 6452 81283 6453 81323
rect 6891 81292 6892 81332
rect 6932 81292 6933 81332
rect 6891 81283 6933 81292
rect 7162 81332 7220 81333
rect 7162 81292 7171 81332
rect 7211 81292 7220 81332
rect 7162 81291 7220 81292
rect 7738 81332 7796 81333
rect 7738 81292 7747 81332
rect 7787 81292 7796 81332
rect 7738 81291 7796 81292
rect 8054 81332 8096 81341
rect 8054 81292 8055 81332
rect 8095 81292 8096 81332
rect 8054 81283 8096 81292
rect 8235 81332 8277 81341
rect 8235 81292 8236 81332
rect 8276 81292 8277 81332
rect 8235 81283 8277 81292
rect 8410 81332 8468 81333
rect 8410 81292 8419 81332
rect 8459 81292 8468 81332
rect 8410 81291 8468 81292
rect 9099 81332 9141 81341
rect 11290 81332 11348 81333
rect 9099 81292 9100 81332
rect 9140 81292 9141 81332
rect 9099 81283 9141 81292
rect 10347 81323 10389 81332
rect 10347 81283 10348 81323
rect 10388 81283 10389 81323
rect 11290 81292 11299 81332
rect 11339 81292 11348 81332
rect 11290 81291 11348 81292
rect 11403 81332 11445 81341
rect 11403 81292 11404 81332
rect 11444 81292 11445 81332
rect 11403 81283 11445 81292
rect 11787 81332 11829 81341
rect 13515 81332 13557 81341
rect 16587 81332 16629 81341
rect 11787 81292 11788 81332
rect 11828 81292 11829 81332
rect 11787 81283 11829 81292
rect 12363 81323 12405 81332
rect 12363 81283 12364 81323
rect 12404 81283 12405 81323
rect 6411 81274 6453 81283
rect 10347 81274 10389 81283
rect 12363 81274 12405 81283
rect 12843 81323 12885 81332
rect 12843 81283 12844 81323
rect 12884 81283 12885 81323
rect 13515 81292 13516 81332
rect 13556 81292 13557 81332
rect 13515 81283 13557 81292
rect 14763 81323 14805 81332
rect 14763 81283 14764 81323
rect 14804 81283 14805 81323
rect 12843 81274 12885 81283
rect 14763 81274 14805 81283
rect 15339 81323 15381 81332
rect 15339 81283 15340 81323
rect 15380 81283 15381 81323
rect 16587 81292 16588 81332
rect 16628 81292 16629 81332
rect 16971 81332 17013 81341
rect 16587 81283 16629 81292
rect 16731 81290 16773 81299
rect 15339 81274 15381 81283
rect 1227 81248 1269 81257
rect 1227 81208 1228 81248
rect 1268 81208 1269 81248
rect 1227 81199 1269 81208
rect 3243 81248 3285 81257
rect 3243 81208 3244 81248
rect 3284 81208 3285 81248
rect 3243 81199 3285 81208
rect 3627 81248 3669 81257
rect 3627 81208 3628 81248
rect 3668 81208 3669 81248
rect 3627 81199 3669 81208
rect 3963 81248 4005 81257
rect 3963 81208 3964 81248
rect 4004 81208 4005 81248
rect 3963 81199 4005 81208
rect 4203 81248 4245 81257
rect 4203 81208 4204 81248
rect 4244 81208 4245 81248
rect 4203 81199 4245 81208
rect 4395 81248 4437 81257
rect 4395 81208 4396 81248
rect 4436 81208 4437 81248
rect 4395 81199 4437 81208
rect 5451 81248 5493 81257
rect 5451 81208 5452 81248
rect 5492 81208 5493 81248
rect 5451 81199 5493 81208
rect 8619 81248 8661 81257
rect 8619 81208 8620 81248
rect 8660 81208 8661 81248
rect 8619 81199 8661 81208
rect 10731 81248 10773 81257
rect 10731 81208 10732 81248
rect 10772 81208 10773 81248
rect 10731 81199 10773 81208
rect 11883 81248 11925 81257
rect 11883 81208 11884 81248
rect 11924 81208 11925 81248
rect 16731 81250 16732 81290
rect 16772 81250 16773 81290
rect 16971 81292 16972 81332
rect 17012 81292 17013 81332
rect 16971 81283 17013 81292
rect 18394 81332 18452 81333
rect 18394 81292 18403 81332
rect 18443 81292 18452 81332
rect 18394 81291 18452 81292
rect 18507 81332 18549 81341
rect 18507 81292 18508 81332
rect 18548 81292 18549 81332
rect 18507 81283 18549 81292
rect 18891 81332 18933 81341
rect 18891 81292 18892 81332
rect 18932 81292 18933 81332
rect 18891 81283 18933 81292
rect 19467 81323 19509 81332
rect 19467 81283 19468 81323
rect 19508 81283 19509 81323
rect 19467 81274 19509 81283
rect 19947 81323 19989 81332
rect 19947 81283 19948 81323
rect 19988 81283 19989 81323
rect 19947 81274 19989 81283
rect 16731 81241 16773 81250
rect 16858 81248 16916 81249
rect 11883 81199 11925 81208
rect 16858 81208 16867 81248
rect 16907 81208 16916 81248
rect 16858 81207 16916 81208
rect 17739 81248 17781 81257
rect 17739 81208 17740 81248
rect 17780 81208 17781 81248
rect 17739 81199 17781 81208
rect 17931 81248 17973 81257
rect 17931 81208 17932 81248
rect 17972 81208 17973 81248
rect 17931 81199 17973 81208
rect 18987 81248 19029 81257
rect 18987 81208 18988 81248
rect 19028 81208 19029 81248
rect 18987 81199 19029 81208
rect 3867 81164 3909 81173
rect 3867 81124 3868 81164
rect 3908 81124 3909 81164
rect 3867 81115 3909 81124
rect 7563 81164 7605 81173
rect 7563 81124 7564 81164
rect 7604 81124 7605 81164
rect 7563 81115 7605 81124
rect 8410 81164 8468 81165
rect 8410 81124 8419 81164
rect 8459 81124 8468 81164
rect 8410 81123 8468 81124
rect 1467 81080 1509 81089
rect 1467 81040 1468 81080
rect 1508 81040 1509 81080
rect 1467 81031 1509 81040
rect 3051 81080 3093 81089
rect 3051 81040 3052 81080
rect 3092 81040 3093 81080
rect 3051 81031 3093 81040
rect 3483 81080 3525 81089
rect 3483 81040 3484 81080
rect 3524 81040 3525 81080
rect 3483 81031 3525 81040
rect 15147 81080 15189 81089
rect 15147 81040 15148 81080
rect 15188 81040 15189 81080
rect 15147 81031 15189 81040
rect 18171 81080 18213 81089
rect 18171 81040 18172 81080
rect 18212 81040 18213 81080
rect 18171 81031 18213 81040
rect 1152 80912 20448 80936
rect 1152 80872 3688 80912
rect 3728 80872 3770 80912
rect 3810 80872 3852 80912
rect 3892 80872 3934 80912
rect 3974 80872 4016 80912
rect 4056 80872 18808 80912
rect 18848 80872 18890 80912
rect 18930 80872 18972 80912
rect 19012 80872 19054 80912
rect 19094 80872 19136 80912
rect 19176 80872 20448 80912
rect 1152 80848 20448 80872
rect 5931 80744 5973 80753
rect 5931 80704 5932 80744
rect 5972 80704 5973 80744
rect 5931 80695 5973 80704
rect 4347 80660 4389 80669
rect 4347 80620 4348 80660
rect 4388 80620 4389 80660
rect 4347 80611 4389 80620
rect 1227 80576 1269 80585
rect 1227 80536 1228 80576
rect 1268 80536 1269 80576
rect 1227 80527 1269 80536
rect 3339 80576 3381 80585
rect 3339 80536 3340 80576
rect 3380 80536 3381 80576
rect 3339 80527 3381 80536
rect 3723 80576 3765 80585
rect 3723 80536 3724 80576
rect 3764 80536 3765 80576
rect 3723 80527 3765 80536
rect 4107 80576 4149 80585
rect 4107 80536 4108 80576
rect 4148 80536 4149 80576
rect 4107 80527 4149 80536
rect 6682 80576 6740 80577
rect 6682 80536 6691 80576
rect 6731 80536 6740 80576
rect 6682 80535 6740 80536
rect 10347 80576 10389 80585
rect 10347 80536 10348 80576
rect 10388 80536 10389 80576
rect 10347 80527 10389 80536
rect 12459 80576 12501 80585
rect 12459 80536 12460 80576
rect 12500 80536 12501 80576
rect 12459 80527 12501 80536
rect 12843 80576 12885 80585
rect 12843 80536 12844 80576
rect 12884 80536 12885 80576
rect 12843 80527 12885 80536
rect 17163 80576 17205 80585
rect 17163 80536 17164 80576
rect 17204 80536 17205 80576
rect 17163 80527 17205 80536
rect 1707 80492 1749 80501
rect 1707 80452 1708 80492
rect 1748 80452 1749 80492
rect 1707 80443 1749 80452
rect 2947 80492 3005 80493
rect 2947 80452 2956 80492
rect 2996 80452 3005 80492
rect 2947 80451 3005 80452
rect 4491 80492 4533 80501
rect 4491 80452 4492 80492
rect 4532 80452 4533 80492
rect 4491 80443 4533 80452
rect 5731 80492 5789 80493
rect 5731 80452 5740 80492
rect 5780 80452 5789 80492
rect 5731 80451 5789 80452
rect 6106 80492 6164 80493
rect 6106 80452 6115 80492
rect 6155 80452 6164 80492
rect 6106 80451 6164 80452
rect 6411 80492 6453 80501
rect 6411 80452 6412 80492
rect 6452 80452 6453 80492
rect 6411 80443 6453 80452
rect 6550 80492 6592 80501
rect 6550 80452 6551 80492
rect 6591 80452 6592 80492
rect 6550 80443 6592 80452
rect 6795 80492 6837 80501
rect 6795 80452 6796 80492
rect 6836 80452 6837 80492
rect 6795 80443 6837 80452
rect 7083 80492 7125 80501
rect 7083 80452 7084 80492
rect 7124 80452 7125 80492
rect 7083 80443 7125 80452
rect 8323 80492 8381 80493
rect 8323 80452 8332 80492
rect 8372 80452 8381 80492
rect 8323 80451 8381 80452
rect 8899 80492 8957 80493
rect 8899 80452 8908 80492
rect 8948 80452 8957 80492
rect 8899 80451 8957 80452
rect 10155 80492 10197 80501
rect 10155 80452 10156 80492
rect 10196 80452 10197 80492
rect 10155 80443 10197 80452
rect 10731 80492 10773 80501
rect 10731 80452 10732 80492
rect 10772 80452 10773 80492
rect 10731 80443 10773 80452
rect 11971 80492 12029 80493
rect 11971 80452 11980 80492
rect 12020 80452 12029 80492
rect 11971 80451 12029 80452
rect 13227 80492 13269 80501
rect 13227 80452 13228 80492
rect 13268 80452 13269 80492
rect 13227 80443 13269 80452
rect 14467 80492 14525 80493
rect 14467 80452 14476 80492
rect 14516 80452 14525 80492
rect 14467 80451 14525 80452
rect 14955 80492 14997 80501
rect 14955 80452 14956 80492
rect 14996 80452 14997 80492
rect 14955 80443 14997 80452
rect 16195 80492 16253 80493
rect 16195 80452 16204 80492
rect 16244 80452 16253 80492
rect 16195 80451 16253 80452
rect 16666 80492 16724 80493
rect 16666 80452 16675 80492
rect 16715 80452 16724 80492
rect 16666 80451 16724 80452
rect 16779 80492 16821 80501
rect 16779 80452 16780 80492
rect 16820 80452 16821 80492
rect 16779 80443 16821 80452
rect 17259 80492 17301 80501
rect 17259 80452 17260 80492
rect 17300 80452 17301 80492
rect 17259 80443 17301 80452
rect 17731 80492 17789 80493
rect 17731 80452 17740 80492
rect 17780 80452 17789 80492
rect 17731 80451 17789 80452
rect 18219 80492 18277 80493
rect 18219 80452 18228 80492
rect 18268 80452 18277 80492
rect 18219 80451 18277 80452
rect 18603 80492 18645 80501
rect 18603 80452 18604 80492
rect 18644 80452 18645 80492
rect 18603 80443 18645 80452
rect 19843 80492 19901 80493
rect 19843 80452 19852 80492
rect 19892 80452 19901 80492
rect 19843 80451 19901 80452
rect 3579 80408 3621 80417
rect 3579 80368 3580 80408
rect 3620 80368 3621 80408
rect 3579 80359 3621 80368
rect 6315 80408 6357 80417
rect 6315 80368 6316 80408
rect 6356 80368 6357 80408
rect 6315 80359 6357 80368
rect 6874 80408 6932 80409
rect 6874 80368 6883 80408
rect 6923 80368 6932 80408
rect 6874 80367 6932 80368
rect 12171 80408 12213 80417
rect 12171 80368 12172 80408
rect 12212 80368 12213 80408
rect 12171 80359 12213 80368
rect 14667 80408 14709 80417
rect 14667 80368 14668 80408
rect 14708 80368 14709 80408
rect 14667 80359 14709 80368
rect 16395 80408 16437 80417
rect 16395 80368 16396 80408
rect 16436 80368 16437 80408
rect 16395 80359 16437 80368
rect 1467 80324 1509 80333
rect 1467 80284 1468 80324
rect 1508 80284 1509 80324
rect 1467 80275 1509 80284
rect 3147 80324 3189 80333
rect 3147 80284 3148 80324
rect 3188 80284 3189 80324
rect 3147 80275 3189 80284
rect 3963 80324 4005 80333
rect 3963 80284 3964 80324
rect 4004 80284 4005 80324
rect 3963 80275 4005 80284
rect 8523 80324 8565 80333
rect 8523 80284 8524 80324
rect 8564 80284 8565 80324
rect 8523 80275 8565 80284
rect 8715 80324 8757 80333
rect 8715 80284 8716 80324
rect 8756 80284 8757 80324
rect 8715 80275 8757 80284
rect 10587 80324 10629 80333
rect 10587 80284 10588 80324
rect 10628 80284 10629 80324
rect 10587 80275 10629 80284
rect 12699 80324 12741 80333
rect 12699 80284 12700 80324
rect 12740 80284 12741 80324
rect 12699 80275 12741 80284
rect 13083 80324 13125 80333
rect 13083 80284 13084 80324
rect 13124 80284 13125 80324
rect 13083 80275 13125 80284
rect 18411 80324 18453 80333
rect 18411 80284 18412 80324
rect 18452 80284 18453 80324
rect 18411 80275 18453 80284
rect 20043 80324 20085 80333
rect 20043 80284 20044 80324
rect 20084 80284 20085 80324
rect 20043 80275 20085 80284
rect 1152 80156 20452 80180
rect 1152 80116 4928 80156
rect 4968 80116 5010 80156
rect 5050 80116 5092 80156
rect 5132 80116 5174 80156
rect 5214 80116 5256 80156
rect 5296 80116 20048 80156
rect 20088 80116 20130 80156
rect 20170 80116 20212 80156
rect 20252 80116 20294 80156
rect 20334 80116 20376 80156
rect 20416 80116 20452 80156
rect 1152 80092 20452 80116
rect 3610 79988 3668 79989
rect 3610 79948 3619 79988
rect 3659 79948 3668 79988
rect 3610 79947 3668 79948
rect 7467 79988 7509 79997
rect 7467 79948 7468 79988
rect 7508 79948 7509 79988
rect 7467 79939 7509 79948
rect 9483 79988 9525 79997
rect 9483 79948 9484 79988
rect 9524 79948 9525 79988
rect 9483 79939 9525 79948
rect 10299 79988 10341 79997
rect 10299 79948 10300 79988
rect 10340 79948 10341 79988
rect 10299 79939 10341 79948
rect 17019 79988 17061 79997
rect 17019 79948 17020 79988
rect 17060 79948 17061 79988
rect 17019 79939 17061 79948
rect 5835 79904 5877 79913
rect 3426 79895 3472 79904
rect 3426 79855 3427 79895
rect 3467 79855 3472 79895
rect 5835 79864 5836 79904
rect 5876 79864 5877 79904
rect 5835 79855 5877 79864
rect 9915 79904 9957 79913
rect 9915 79864 9916 79904
rect 9956 79864 9957 79904
rect 9915 79855 9957 79864
rect 12507 79904 12549 79913
rect 12507 79864 12508 79904
rect 12548 79864 12549 79904
rect 12507 79855 12549 79864
rect 3426 79846 3472 79855
rect 1515 79820 1557 79829
rect 3130 79820 3188 79821
rect 3514 79820 3572 79821
rect 1515 79780 1516 79820
rect 1556 79780 1557 79820
rect 1515 79771 1557 79780
rect 2763 79811 2805 79820
rect 2763 79771 2764 79811
rect 2804 79771 2805 79811
rect 3130 79780 3139 79820
rect 3179 79780 3188 79820
rect 3130 79779 3188 79780
rect 3243 79811 3285 79820
rect 2763 79762 2805 79771
rect 3243 79771 3244 79811
rect 3284 79771 3285 79811
rect 3514 79780 3523 79820
rect 3563 79780 3572 79820
rect 3514 79779 3572 79780
rect 3648 79820 3706 79821
rect 3648 79780 3657 79820
rect 3697 79780 3706 79820
rect 3648 79779 3706 79780
rect 4395 79820 4437 79829
rect 6027 79820 6069 79829
rect 7738 79820 7796 79821
rect 4395 79780 4396 79820
rect 4436 79780 4437 79820
rect 4395 79771 4437 79780
rect 5643 79811 5685 79820
rect 5643 79771 5644 79811
rect 5684 79771 5685 79811
rect 6027 79780 6028 79820
rect 6068 79780 6069 79820
rect 6027 79771 6069 79780
rect 7275 79811 7317 79820
rect 7275 79771 7276 79811
rect 7316 79771 7317 79811
rect 7738 79780 7747 79820
rect 7787 79780 7796 79820
rect 7738 79779 7796 79780
rect 7851 79820 7893 79829
rect 7851 79780 7852 79820
rect 7892 79780 7893 79820
rect 7851 79771 7893 79780
rect 8235 79820 8277 79829
rect 12171 79820 12213 79829
rect 8235 79780 8236 79820
rect 8276 79780 8277 79820
rect 8235 79771 8277 79780
rect 8811 79811 8853 79820
rect 8811 79771 8812 79811
rect 8852 79771 8853 79811
rect 3243 79762 3285 79771
rect 5643 79762 5685 79771
rect 7275 79762 7317 79771
rect 8811 79762 8853 79771
rect 9291 79811 9333 79820
rect 9291 79771 9292 79811
rect 9332 79771 9333 79811
rect 12171 79780 12172 79820
rect 12212 79780 12213 79820
rect 12637 79820 12679 79829
rect 12171 79771 12213 79780
rect 12299 79796 12341 79805
rect 9291 79762 9333 79771
rect 12299 79756 12300 79796
rect 12340 79756 12341 79796
rect 12637 79780 12638 79820
rect 12678 79780 12679 79820
rect 12637 79771 12679 79780
rect 12747 79820 12789 79829
rect 12747 79780 12748 79820
rect 12788 79780 12789 79820
rect 12747 79771 12789 79780
rect 12939 79820 12981 79829
rect 12939 79780 12940 79820
rect 12980 79780 12981 79820
rect 12939 79771 12981 79780
rect 13131 79820 13173 79829
rect 14763 79820 14805 79829
rect 17451 79820 17493 79829
rect 13131 79780 13132 79820
rect 13172 79780 13173 79820
rect 13131 79771 13173 79780
rect 14379 79811 14421 79820
rect 14379 79771 14380 79811
rect 14420 79771 14421 79811
rect 14763 79780 14764 79820
rect 14804 79780 14805 79820
rect 14763 79771 14805 79780
rect 16011 79811 16053 79820
rect 16011 79771 16012 79811
rect 16052 79771 16053 79811
rect 17451 79780 17452 79820
rect 17492 79780 17493 79820
rect 17451 79771 17493 79780
rect 18699 79811 18741 79820
rect 18699 79771 18700 79811
rect 18740 79771 18741 79811
rect 14379 79762 14421 79771
rect 16011 79762 16053 79771
rect 18699 79762 18741 79771
rect 12299 79747 12341 79756
rect 3915 79736 3957 79745
rect 3915 79696 3916 79736
rect 3956 79696 3957 79736
rect 3915 79687 3957 79696
rect 8331 79736 8373 79745
rect 8331 79696 8332 79736
rect 8372 79696 8373 79736
rect 8331 79687 8373 79696
rect 9675 79736 9717 79745
rect 9675 79696 9676 79736
rect 9716 79696 9717 79736
rect 9675 79687 9717 79696
rect 10059 79736 10101 79745
rect 10059 79696 10060 79736
rect 10100 79696 10101 79736
rect 10059 79687 10101 79696
rect 10635 79736 10677 79745
rect 10635 79696 10636 79736
rect 10676 79696 10677 79736
rect 10635 79687 10677 79696
rect 11115 79736 11157 79745
rect 11115 79696 11116 79736
rect 11156 79696 11157 79736
rect 11115 79687 11157 79696
rect 11787 79736 11829 79745
rect 11787 79696 11788 79736
rect 11828 79696 11829 79736
rect 11787 79687 11829 79696
rect 16683 79736 16725 79745
rect 16683 79696 16684 79736
rect 16724 79696 16725 79736
rect 16683 79687 16725 79696
rect 17259 79736 17301 79745
rect 17259 79696 17260 79736
rect 17300 79696 17301 79736
rect 17259 79687 17301 79696
rect 19371 79736 19413 79745
rect 19371 79696 19372 79736
rect 19412 79696 19413 79736
rect 19371 79687 19413 79696
rect 19755 79736 19797 79745
rect 19755 79696 19756 79736
rect 19796 79696 19797 79736
rect 19755 79687 19797 79696
rect 20139 79736 20181 79745
rect 20139 79696 20140 79736
rect 20180 79696 20181 79736
rect 20139 79687 20181 79696
rect 12747 79652 12789 79661
rect 12747 79612 12748 79652
rect 12788 79612 12789 79652
rect 12747 79603 12789 79612
rect 19611 79652 19653 79661
rect 19611 79612 19612 79652
rect 19652 79612 19653 79652
rect 19611 79603 19653 79612
rect 20379 79652 20421 79661
rect 20379 79612 20380 79652
rect 20420 79612 20421 79652
rect 20379 79603 20421 79612
rect 2955 79568 2997 79577
rect 2955 79528 2956 79568
rect 2996 79528 2997 79568
rect 2955 79519 2997 79528
rect 4155 79568 4197 79577
rect 4155 79528 4156 79568
rect 4196 79528 4197 79568
rect 4155 79519 4197 79528
rect 10395 79568 10437 79577
rect 10395 79528 10396 79568
rect 10436 79528 10437 79568
rect 10395 79519 10437 79528
rect 11355 79568 11397 79577
rect 11355 79528 11356 79568
rect 11396 79528 11397 79568
rect 11355 79519 11397 79528
rect 12027 79568 12069 79577
rect 12027 79528 12028 79568
rect 12068 79528 12069 79568
rect 12027 79519 12069 79528
rect 14571 79568 14613 79577
rect 14571 79528 14572 79568
rect 14612 79528 14613 79568
rect 14571 79519 14613 79528
rect 16203 79568 16245 79577
rect 16203 79528 16204 79568
rect 16244 79528 16245 79568
rect 16203 79519 16245 79528
rect 16923 79568 16965 79577
rect 16923 79528 16924 79568
rect 16964 79528 16965 79568
rect 16923 79519 16965 79528
rect 18891 79568 18933 79577
rect 18891 79528 18892 79568
rect 18932 79528 18933 79568
rect 18891 79519 18933 79528
rect 19995 79568 20037 79577
rect 19995 79528 19996 79568
rect 20036 79528 20037 79568
rect 19995 79519 20037 79528
rect 1152 79400 20448 79424
rect 1152 79360 3688 79400
rect 3728 79360 3770 79400
rect 3810 79360 3852 79400
rect 3892 79360 3934 79400
rect 3974 79360 4016 79400
rect 4056 79360 18808 79400
rect 18848 79360 18890 79400
rect 18930 79360 18972 79400
rect 19012 79360 19054 79400
rect 19094 79360 19136 79400
rect 19176 79360 20448 79400
rect 1152 79336 20448 79360
rect 3243 79232 3285 79241
rect 3243 79192 3244 79232
rect 3284 79192 3285 79232
rect 3243 79183 3285 79192
rect 5499 79148 5541 79157
rect 5499 79108 5500 79148
rect 5540 79108 5541 79148
rect 5499 79099 5541 79108
rect 17931 79148 17973 79157
rect 17931 79108 17932 79148
rect 17972 79108 17973 79148
rect 17931 79099 17973 79108
rect 1227 79064 1269 79073
rect 1227 79024 1228 79064
rect 1268 79024 1269 79064
rect 1227 79015 1269 79024
rect 8139 79064 8181 79073
rect 8139 79024 8140 79064
rect 8180 79024 8181 79064
rect 8139 79015 8181 79024
rect 9771 79064 9813 79073
rect 9771 79024 9772 79064
rect 9812 79024 9813 79064
rect 9771 79015 9813 79024
rect 9963 79064 10005 79073
rect 9963 79024 9964 79064
rect 10004 79024 10005 79064
rect 9963 79015 10005 79024
rect 10731 79064 10773 79073
rect 10731 79024 10732 79064
rect 10772 79024 10773 79064
rect 10731 79015 10773 79024
rect 14283 79064 14325 79073
rect 14283 79024 14284 79064
rect 14324 79024 14325 79064
rect 14283 79015 14325 79024
rect 15562 79064 15620 79065
rect 15562 79024 15571 79064
rect 15611 79024 15620 79064
rect 15562 79023 15620 79024
rect 15915 79064 15957 79073
rect 15915 79024 15916 79064
rect 15956 79024 15957 79064
rect 15915 79015 15957 79024
rect 16107 79064 16149 79073
rect 16107 79024 16108 79064
rect 16148 79024 16149 79064
rect 16107 79015 16149 79024
rect 12843 78991 12885 79000
rect 1611 78980 1653 78989
rect 1611 78940 1612 78980
rect 1652 78940 1653 78980
rect 1611 78931 1653 78940
rect 2851 78980 2909 78981
rect 2851 78940 2860 78980
rect 2900 78940 2909 78980
rect 2851 78939 2909 78940
rect 3243 78980 3285 78989
rect 3243 78940 3244 78980
rect 3284 78940 3285 78980
rect 3243 78931 3285 78940
rect 3358 78980 3400 78989
rect 3358 78940 3359 78980
rect 3399 78940 3400 78980
rect 3358 78931 3400 78940
rect 3531 78980 3573 78989
rect 3531 78940 3532 78980
rect 3572 78940 3573 78980
rect 3531 78931 3573 78940
rect 3915 78980 3957 78989
rect 3915 78940 3916 78980
rect 3956 78940 3957 78980
rect 3915 78931 3957 78940
rect 5155 78980 5213 78981
rect 5155 78940 5164 78980
rect 5204 78940 5213 78980
rect 5155 78939 5213 78940
rect 5643 78980 5685 78989
rect 5643 78940 5644 78980
rect 5684 78940 5685 78980
rect 5643 78931 5685 78940
rect 5835 78980 5877 78989
rect 5835 78940 5836 78980
rect 5876 78940 5877 78980
rect 5835 78931 5877 78940
rect 7075 78980 7133 78981
rect 7075 78940 7084 78980
rect 7124 78940 7133 78980
rect 7075 78939 7133 78940
rect 7642 78980 7700 78981
rect 7642 78940 7651 78980
rect 7691 78940 7700 78980
rect 7642 78939 7700 78940
rect 7755 78980 7797 78989
rect 7755 78940 7756 78980
rect 7796 78940 7797 78980
rect 7755 78931 7797 78940
rect 8235 78980 8277 78989
rect 8235 78940 8236 78980
rect 8276 78940 8277 78980
rect 8235 78931 8277 78940
rect 8710 78980 8768 78981
rect 8710 78940 8719 78980
rect 8759 78940 8768 78980
rect 8710 78939 8768 78940
rect 9195 78980 9253 78981
rect 9195 78940 9204 78980
rect 9244 78940 9253 78980
rect 9195 78939 9253 78940
rect 11115 78980 11157 78989
rect 11115 78940 11116 78980
rect 11156 78940 11157 78980
rect 11115 78931 11157 78940
rect 12355 78980 12413 78981
rect 12355 78940 12364 78980
rect 12404 78940 12413 78980
rect 12355 78939 12413 78940
rect 12730 78980 12788 78981
rect 12730 78940 12739 78980
rect 12779 78940 12788 78980
rect 12843 78951 12844 78991
rect 12884 78951 12885 78991
rect 12843 78942 12885 78951
rect 12980 78980 13038 78981
rect 12730 78939 12788 78940
rect 12980 78940 12989 78980
rect 13029 78940 13038 78980
rect 12980 78939 13038 78940
rect 13114 78980 13172 78981
rect 13114 78940 13123 78980
rect 13163 78940 13172 78980
rect 13114 78939 13172 78940
rect 13248 78980 13306 78981
rect 13248 78940 13257 78980
rect 13297 78940 13306 78980
rect 13248 78939 13306 78940
rect 13786 78980 13844 78981
rect 13786 78940 13795 78980
rect 13835 78940 13844 78980
rect 13786 78939 13844 78940
rect 13899 78980 13941 78989
rect 13899 78940 13900 78980
rect 13940 78940 13941 78980
rect 13899 78931 13941 78940
rect 14379 78980 14421 78989
rect 14379 78940 14380 78980
rect 14420 78940 14421 78980
rect 14379 78931 14421 78940
rect 14851 78980 14909 78981
rect 14851 78940 14860 78980
rect 14900 78940 14909 78980
rect 14851 78939 14909 78940
rect 15339 78980 15397 78981
rect 15339 78940 15348 78980
rect 15388 78940 15397 78980
rect 15339 78939 15397 78940
rect 16491 78980 16533 78989
rect 16491 78940 16492 78980
rect 16532 78940 16533 78980
rect 16491 78931 16533 78940
rect 17731 78980 17789 78981
rect 17731 78940 17740 78980
rect 17780 78940 17789 78980
rect 17731 78939 17789 78940
rect 18123 78980 18165 78989
rect 18123 78940 18124 78980
rect 18164 78940 18165 78980
rect 18123 78931 18165 78940
rect 19363 78980 19421 78981
rect 19363 78940 19372 78980
rect 19412 78940 19421 78980
rect 19363 78939 19421 78940
rect 19702 78980 19744 78989
rect 19702 78940 19703 78980
rect 19743 78940 19744 78980
rect 19702 78931 19744 78940
rect 19834 78980 19892 78981
rect 19834 78940 19843 78980
rect 19883 78940 19892 78980
rect 19834 78939 19892 78940
rect 19947 78980 19989 78989
rect 19947 78940 19948 78980
rect 19988 78940 19989 78980
rect 19947 78931 19989 78940
rect 7275 78896 7317 78905
rect 7275 78856 7276 78896
rect 7316 78856 7317 78896
rect 7275 78847 7317 78856
rect 9531 78896 9573 78905
rect 9531 78856 9532 78896
rect 9572 78856 9573 78896
rect 9531 78847 9573 78856
rect 12555 78896 12597 78905
rect 12555 78856 12556 78896
rect 12596 78856 12597 78896
rect 12555 78847 12597 78856
rect 1467 78812 1509 78821
rect 1467 78772 1468 78812
rect 1508 78772 1509 78812
rect 1467 78763 1509 78772
rect 3051 78812 3093 78821
rect 3051 78772 3052 78812
rect 3092 78772 3093 78812
rect 3051 78763 3093 78772
rect 5355 78812 5397 78821
rect 5355 78772 5356 78812
rect 5396 78772 5397 78812
rect 5355 78763 5397 78772
rect 9387 78812 9429 78821
rect 9387 78772 9388 78812
rect 9428 78772 9429 78812
rect 9387 78763 9429 78772
rect 10203 78812 10245 78821
rect 10203 78772 10204 78812
rect 10244 78772 10245 78812
rect 10203 78763 10245 78772
rect 10491 78812 10533 78821
rect 10491 78772 10492 78812
rect 10532 78772 10533 78812
rect 10491 78763 10533 78772
rect 13210 78812 13268 78813
rect 13210 78772 13219 78812
rect 13259 78772 13268 78812
rect 13210 78771 13268 78772
rect 15675 78812 15717 78821
rect 15675 78772 15676 78812
rect 15716 78772 15717 78812
rect 15675 78763 15717 78772
rect 16347 78812 16389 78821
rect 16347 78772 16348 78812
rect 16388 78772 16389 78812
rect 16347 78763 16389 78772
rect 19563 78812 19605 78821
rect 19563 78772 19564 78812
rect 19604 78772 19605 78812
rect 19563 78763 19605 78772
rect 20026 78812 20084 78813
rect 20026 78772 20035 78812
rect 20075 78772 20084 78812
rect 20026 78771 20084 78772
rect 1152 78644 20452 78668
rect 1152 78604 4928 78644
rect 4968 78604 5010 78644
rect 5050 78604 5092 78644
rect 5132 78604 5174 78644
rect 5214 78604 5256 78644
rect 5296 78604 20048 78644
rect 20088 78604 20130 78644
rect 20170 78604 20212 78644
rect 20252 78604 20294 78644
rect 20334 78604 20376 78644
rect 20416 78604 20452 78644
rect 1152 78580 20452 78604
rect 3034 78476 3092 78477
rect 3034 78436 3043 78476
rect 3083 78436 3092 78476
rect 3034 78435 3092 78436
rect 5355 78476 5397 78485
rect 5355 78436 5356 78476
rect 5396 78436 5397 78476
rect 5355 78427 5397 78436
rect 8715 78476 8757 78485
rect 8715 78436 8716 78476
rect 8756 78436 8757 78476
rect 8715 78427 8757 78436
rect 11979 78476 12021 78485
rect 11979 78436 11980 78476
rect 12020 78436 12021 78476
rect 11979 78427 12021 78436
rect 12315 78476 12357 78485
rect 12315 78436 12316 78476
rect 12356 78436 12357 78476
rect 12315 78427 12357 78436
rect 13899 78476 13941 78485
rect 13899 78436 13900 78476
rect 13940 78436 13941 78476
rect 13899 78427 13941 78436
rect 14859 78476 14901 78485
rect 14859 78436 14860 78476
rect 14900 78436 14901 78476
rect 14859 78427 14901 78436
rect 16971 78476 17013 78485
rect 16971 78436 16972 78476
rect 17012 78436 17013 78476
rect 16971 78427 17013 78436
rect 20314 78476 20372 78477
rect 20314 78436 20323 78476
rect 20363 78436 20372 78476
rect 20314 78435 20372 78436
rect 17530 78392 17588 78393
rect 17530 78352 17539 78392
rect 17579 78352 17588 78392
rect 17530 78351 17588 78352
rect 1227 78308 1269 78317
rect 3339 78308 3381 78317
rect 1227 78268 1228 78308
rect 1268 78268 1269 78308
rect 1227 78259 1269 78268
rect 2475 78299 2517 78308
rect 2475 78259 2476 78299
rect 2516 78259 2517 78299
rect 2475 78250 2517 78259
rect 3195 78294 3253 78295
rect 3195 78254 3204 78294
rect 3244 78254 3253 78294
rect 3339 78268 3340 78308
rect 3380 78268 3381 78308
rect 3339 78259 3381 78268
rect 3597 78308 3639 78317
rect 3597 78268 3598 78308
rect 3638 78268 3639 78308
rect 3597 78259 3639 78268
rect 3723 78308 3765 78317
rect 3723 78268 3724 78308
rect 3764 78268 3765 78308
rect 3723 78259 3765 78268
rect 4107 78308 4149 78317
rect 6987 78308 7029 78317
rect 4107 78268 4108 78308
rect 4148 78268 4149 78308
rect 4107 78259 4149 78268
rect 4683 78299 4725 78308
rect 4683 78259 4684 78299
rect 4724 78259 4725 78299
rect 3195 78253 3253 78254
rect 4683 78250 4725 78259
rect 5163 78299 5205 78308
rect 5163 78259 5164 78299
rect 5204 78259 5205 78299
rect 5163 78250 5205 78259
rect 5739 78299 5781 78308
rect 5739 78259 5740 78299
rect 5780 78259 5781 78299
rect 6987 78268 6988 78308
rect 7028 78268 7029 78308
rect 6987 78259 7029 78268
rect 7275 78308 7317 78317
rect 7275 78268 7276 78308
rect 7316 78268 7317 78308
rect 8907 78308 8949 78317
rect 10539 78308 10581 78317
rect 12171 78308 12213 78317
rect 7275 78259 7317 78268
rect 8523 78287 8565 78296
rect 5739 78250 5781 78259
rect 8523 78247 8524 78287
rect 8564 78247 8565 78287
rect 8907 78268 8908 78308
rect 8948 78268 8949 78308
rect 8907 78259 8949 78268
rect 10155 78299 10197 78308
rect 10155 78259 10156 78299
rect 10196 78259 10197 78299
rect 10539 78268 10540 78308
rect 10580 78268 10581 78308
rect 10539 78259 10581 78268
rect 11787 78299 11829 78308
rect 11787 78259 11788 78299
rect 11828 78259 11829 78299
rect 12171 78268 12172 78308
rect 12212 78268 12213 78308
rect 12171 78259 12213 78268
rect 12459 78308 12501 78317
rect 14763 78308 14805 78317
rect 12459 78268 12460 78308
rect 12500 78268 12501 78308
rect 12459 78259 12501 78268
rect 13707 78299 13749 78308
rect 13707 78259 13708 78299
rect 13748 78259 13749 78299
rect 14763 78268 14764 78308
rect 14804 78268 14805 78308
rect 14763 78259 14805 78268
rect 14938 78308 14996 78309
rect 14938 78268 14947 78308
rect 14987 78268 14996 78308
rect 14938 78267 14996 78268
rect 15226 78308 15284 78309
rect 15226 78268 15235 78308
rect 15275 78268 15284 78308
rect 15226 78267 15284 78268
rect 15339 78308 15381 78317
rect 15339 78268 15340 78308
rect 15380 78268 15381 78308
rect 15339 78259 15381 78268
rect 15723 78308 15765 78317
rect 17722 78308 17780 78309
rect 15723 78268 15724 78308
rect 15764 78268 15765 78308
rect 15723 78259 15765 78268
rect 16299 78299 16341 78308
rect 16299 78259 16300 78299
rect 16340 78259 16341 78299
rect 10155 78250 10197 78259
rect 11787 78250 11829 78259
rect 13707 78250 13749 78259
rect 16299 78250 16341 78259
rect 16779 78299 16821 78308
rect 16779 78259 16780 78299
rect 16820 78259 16821 78299
rect 17722 78268 17731 78308
rect 17771 78268 17780 78308
rect 18699 78308 18741 78317
rect 17722 78267 17780 78268
rect 18219 78288 18261 78297
rect 16779 78250 16821 78259
rect 8523 78238 8565 78247
rect 18219 78248 18220 78288
rect 18260 78248 18261 78288
rect 18699 78268 18700 78308
rect 18740 78268 18741 78308
rect 18699 78259 18741 78268
rect 19179 78308 19221 78317
rect 19179 78268 19180 78308
rect 19220 78268 19221 78308
rect 19179 78259 19221 78268
rect 19289 78308 19347 78309
rect 19289 78268 19298 78308
rect 19338 78268 19347 78308
rect 19289 78267 19347 78268
rect 19563 78308 19605 78317
rect 19563 78268 19564 78308
rect 19604 78268 19605 78308
rect 19563 78259 19605 78268
rect 19851 78308 19893 78317
rect 19851 78268 19852 78308
rect 19892 78268 19893 78308
rect 19851 78259 19893 78268
rect 19990 78308 20032 78317
rect 19990 78268 19991 78308
rect 20031 78268 20032 78308
rect 19990 78259 20032 78268
rect 20235 78308 20277 78317
rect 20235 78268 20236 78308
rect 20276 78268 20277 78308
rect 20235 78259 20277 78268
rect 18219 78239 18261 78248
rect 4203 78224 4245 78233
rect 4203 78184 4204 78224
rect 4244 78184 4245 78224
rect 4203 78175 4245 78184
rect 14091 78224 14133 78233
rect 14091 78184 14092 78224
rect 14132 78184 14133 78224
rect 14091 78175 14133 78184
rect 15819 78224 15861 78233
rect 15819 78184 15820 78224
rect 15860 78184 15861 78224
rect 15819 78175 15861 78184
rect 17163 78224 17205 78233
rect 17163 78184 17164 78224
rect 17204 78184 17205 78224
rect 17163 78175 17205 78184
rect 18795 78224 18837 78233
rect 18795 78184 18796 78224
rect 18836 78184 18837 78224
rect 18795 78175 18837 78184
rect 20122 78224 20180 78225
rect 20122 78184 20131 78224
rect 20171 78184 20180 78224
rect 20122 78183 20180 78184
rect 5547 78140 5589 78149
rect 5547 78100 5548 78140
rect 5588 78100 5589 78140
rect 5547 78091 5589 78100
rect 10347 78140 10389 78149
rect 10347 78100 10348 78140
rect 10388 78100 10389 78140
rect 10347 78091 10389 78100
rect 19563 78140 19605 78149
rect 19563 78100 19564 78140
rect 19604 78100 19605 78140
rect 19563 78091 19605 78100
rect 2667 78056 2709 78065
rect 2667 78016 2668 78056
rect 2708 78016 2709 78056
rect 2667 78007 2709 78016
rect 14331 78056 14373 78065
rect 14331 78016 14332 78056
rect 14372 78016 14373 78056
rect 14331 78007 14373 78016
rect 17403 78056 17445 78065
rect 17403 78016 17404 78056
rect 17444 78016 17445 78056
rect 17403 78007 17445 78016
rect 1152 77888 20448 77912
rect 1152 77848 3688 77888
rect 3728 77848 3770 77888
rect 3810 77848 3852 77888
rect 3892 77848 3934 77888
rect 3974 77848 4016 77888
rect 4056 77848 18808 77888
rect 18848 77848 18890 77888
rect 18930 77848 18972 77888
rect 19012 77848 19054 77888
rect 19094 77848 19136 77888
rect 19176 77848 20448 77888
rect 1152 77824 20448 77848
rect 10539 77720 10581 77729
rect 10539 77680 10540 77720
rect 10580 77680 10581 77720
rect 10539 77671 10581 77680
rect 15291 77720 15333 77729
rect 15291 77680 15292 77720
rect 15332 77680 15333 77720
rect 15291 77671 15333 77680
rect 20026 77720 20084 77721
rect 20026 77680 20035 77720
rect 20075 77680 20084 77720
rect 20026 77679 20084 77680
rect 1467 77636 1509 77645
rect 1467 77596 1468 77636
rect 1508 77596 1509 77636
rect 1467 77587 1509 77596
rect 14571 77636 14613 77645
rect 14571 77596 14572 77636
rect 14612 77596 14613 77636
rect 14571 77587 14613 77596
rect 19851 77636 19893 77645
rect 19851 77596 19852 77636
rect 19892 77596 19893 77636
rect 19851 77587 19893 77596
rect 1227 77552 1269 77561
rect 1227 77512 1228 77552
rect 1268 77512 1269 77552
rect 1227 77503 1269 77512
rect 1611 77552 1653 77561
rect 1611 77512 1612 77552
rect 1652 77512 1653 77552
rect 1611 77503 1653 77512
rect 12555 77552 12597 77561
rect 12555 77512 12556 77552
rect 12596 77512 12597 77552
rect 12555 77503 12597 77512
rect 12747 77552 12789 77561
rect 12747 77512 12748 77552
rect 12788 77512 12789 77552
rect 12747 77503 12789 77512
rect 15051 77552 15093 77561
rect 15051 77512 15052 77552
rect 15092 77512 15093 77552
rect 15051 77503 15093 77512
rect 16011 77552 16053 77561
rect 16011 77512 16012 77552
rect 16052 77512 16053 77552
rect 16011 77503 16053 77512
rect 2187 77468 2229 77477
rect 2187 77428 2188 77468
rect 2228 77428 2229 77468
rect 2187 77419 2229 77428
rect 3427 77468 3485 77469
rect 3427 77428 3436 77468
rect 3476 77428 3485 77468
rect 3427 77427 3485 77428
rect 3819 77468 3861 77477
rect 3819 77428 3820 77468
rect 3860 77428 3861 77468
rect 3819 77419 3861 77428
rect 5059 77468 5117 77469
rect 5059 77428 5068 77468
rect 5108 77428 5117 77468
rect 5059 77427 5117 77428
rect 5739 77468 5781 77477
rect 5739 77428 5740 77468
rect 5780 77428 5781 77468
rect 5739 77419 5781 77428
rect 6979 77468 7037 77469
rect 6979 77428 6988 77468
rect 7028 77428 7037 77468
rect 6979 77427 7037 77428
rect 7555 77468 7613 77469
rect 7555 77428 7564 77468
rect 7604 77428 7613 77468
rect 7555 77427 7613 77428
rect 8811 77468 8853 77477
rect 8811 77428 8812 77468
rect 8852 77428 8853 77468
rect 8811 77419 8853 77428
rect 9099 77468 9141 77477
rect 9099 77428 9100 77468
rect 9140 77428 9141 77468
rect 9099 77419 9141 77428
rect 10339 77468 10397 77469
rect 10339 77428 10348 77468
rect 10388 77428 10397 77468
rect 10339 77427 10397 77428
rect 10731 77468 10773 77477
rect 10731 77428 10732 77468
rect 10772 77428 10773 77468
rect 10731 77419 10773 77428
rect 11971 77468 12029 77469
rect 11971 77428 11980 77468
rect 12020 77428 12029 77468
rect 11971 77427 12029 77428
rect 13131 77468 13173 77477
rect 13131 77428 13132 77468
rect 13172 77428 13173 77468
rect 13131 77419 13173 77428
rect 14371 77468 14429 77469
rect 14371 77428 14380 77468
rect 14420 77428 14429 77468
rect 14371 77427 14429 77428
rect 15514 77468 15572 77469
rect 15514 77428 15523 77468
rect 15563 77428 15572 77468
rect 15514 77427 15572 77428
rect 15627 77468 15669 77477
rect 15627 77428 15628 77468
rect 15668 77428 15669 77468
rect 15627 77419 15669 77428
rect 16107 77468 16149 77477
rect 16107 77428 16108 77468
rect 16148 77428 16149 77468
rect 16107 77419 16149 77428
rect 16579 77468 16637 77469
rect 16579 77428 16588 77468
rect 16628 77428 16637 77468
rect 16579 77427 16637 77428
rect 17098 77468 17156 77469
rect 17098 77428 17107 77468
rect 17147 77428 17156 77468
rect 17098 77427 17156 77428
rect 17635 77468 17693 77469
rect 17635 77428 17644 77468
rect 17684 77428 17693 77468
rect 17635 77427 17693 77428
rect 18891 77468 18933 77477
rect 18891 77428 18892 77468
rect 18932 77428 18933 77468
rect 18891 77419 18933 77428
rect 19179 77468 19221 77477
rect 19179 77428 19180 77468
rect 19220 77428 19221 77468
rect 19179 77419 19221 77428
rect 19450 77468 19508 77469
rect 19450 77428 19459 77468
rect 19499 77428 19508 77468
rect 19450 77427 19508 77428
rect 20029 77468 20071 77477
rect 20029 77428 20030 77468
rect 20070 77428 20071 77468
rect 20029 77419 20071 77428
rect 20323 77468 20381 77469
rect 20323 77428 20332 77468
rect 20372 77428 20381 77468
rect 20323 77427 20381 77428
rect 12315 77384 12357 77393
rect 12315 77344 12316 77384
rect 12356 77344 12357 77384
rect 12315 77335 12357 77344
rect 12987 77384 13029 77393
rect 12987 77344 12988 77384
rect 13028 77344 13029 77384
rect 12987 77335 13029 77344
rect 17451 77384 17493 77393
rect 17451 77344 17452 77384
rect 17492 77344 17493 77384
rect 17451 77335 17493 77344
rect 19563 77384 19605 77393
rect 19563 77344 19564 77384
rect 19604 77344 19605 77384
rect 19563 77335 19605 77344
rect 1851 77300 1893 77309
rect 1851 77260 1852 77300
rect 1892 77260 1893 77300
rect 1851 77251 1893 77260
rect 3627 77300 3669 77309
rect 3627 77260 3628 77300
rect 3668 77260 3669 77300
rect 3627 77251 3669 77260
rect 5259 77300 5301 77309
rect 5259 77260 5260 77300
rect 5300 77260 5301 77300
rect 5259 77251 5301 77260
rect 7179 77300 7221 77309
rect 7179 77260 7180 77300
rect 7220 77260 7221 77300
rect 7179 77251 7221 77260
rect 7371 77300 7413 77309
rect 7371 77260 7372 77300
rect 7412 77260 7413 77300
rect 7371 77251 7413 77260
rect 12171 77300 12213 77309
rect 12171 77260 12172 77300
rect 12212 77260 12213 77300
rect 12171 77251 12213 77260
rect 17259 77300 17301 77309
rect 17259 77260 17260 77300
rect 17300 77260 17301 77300
rect 17259 77251 17301 77260
rect 20235 77300 20277 77309
rect 20235 77260 20236 77300
rect 20276 77260 20277 77300
rect 20235 77251 20277 77260
rect 1152 77132 20452 77156
rect 1152 77092 4928 77132
rect 4968 77092 5010 77132
rect 5050 77092 5092 77132
rect 5132 77092 5174 77132
rect 5214 77092 5256 77132
rect 5296 77092 20048 77132
rect 20088 77092 20130 77132
rect 20170 77092 20212 77132
rect 20252 77092 20294 77132
rect 20334 77092 20376 77132
rect 20416 77092 20452 77132
rect 1152 77068 20452 77092
rect 4875 76964 4917 76973
rect 4875 76924 4876 76964
rect 4916 76924 4917 76964
rect 4875 76915 4917 76924
rect 10203 76964 10245 76973
rect 10203 76924 10204 76964
rect 10244 76924 10245 76964
rect 10203 76915 10245 76924
rect 15243 76964 15285 76973
rect 15243 76924 15244 76964
rect 15284 76924 15285 76964
rect 15243 76915 15285 76924
rect 15771 76964 15813 76973
rect 15771 76924 15772 76964
rect 15812 76924 15813 76964
rect 15771 76915 15813 76924
rect 19995 76964 20037 76973
rect 19995 76924 19996 76964
rect 20036 76924 20037 76964
rect 19995 76915 20037 76924
rect 10971 76880 11013 76889
rect 10971 76840 10972 76880
rect 11012 76840 11013 76880
rect 10971 76831 11013 76840
rect 13035 76880 13077 76889
rect 13035 76840 13036 76880
rect 13076 76840 13077 76880
rect 13035 76831 13077 76840
rect 15675 76880 15717 76889
rect 15675 76840 15676 76880
rect 15716 76840 15717 76880
rect 15675 76831 15717 76840
rect 1419 76796 1461 76805
rect 3130 76796 3188 76797
rect 1419 76756 1420 76796
rect 1460 76756 1461 76796
rect 1419 76747 1461 76756
rect 2667 76787 2709 76796
rect 2667 76747 2668 76787
rect 2708 76747 2709 76787
rect 3130 76756 3139 76796
rect 3179 76756 3188 76796
rect 3130 76755 3188 76756
rect 3243 76796 3285 76805
rect 3243 76756 3244 76796
rect 3284 76756 3285 76796
rect 3243 76747 3285 76756
rect 3627 76796 3669 76805
rect 6123 76796 6165 76805
rect 3627 76756 3628 76796
rect 3668 76756 3669 76796
rect 3627 76747 3669 76756
rect 4203 76787 4245 76796
rect 4203 76747 4204 76787
rect 4244 76747 4245 76787
rect 2667 76738 2709 76747
rect 4203 76738 4245 76747
rect 4683 76787 4725 76796
rect 4683 76747 4684 76787
rect 4724 76747 4725 76787
rect 6123 76756 6124 76796
rect 6164 76756 6165 76796
rect 6123 76747 6165 76756
rect 6298 76796 6356 76797
rect 6298 76756 6307 76796
rect 6347 76756 6356 76796
rect 6298 76755 6356 76756
rect 6411 76796 6453 76805
rect 6411 76756 6412 76796
rect 6452 76756 6453 76796
rect 6411 76747 6453 76756
rect 6603 76796 6645 76805
rect 8314 76796 8372 76797
rect 6603 76756 6604 76796
rect 6644 76756 6645 76796
rect 6603 76747 6645 76756
rect 7851 76787 7893 76796
rect 7851 76747 7852 76787
rect 7892 76747 7893 76787
rect 8314 76756 8323 76796
rect 8363 76756 8372 76796
rect 8314 76755 8372 76756
rect 8427 76796 8469 76805
rect 8427 76756 8428 76796
rect 8468 76756 8469 76796
rect 8427 76747 8469 76756
rect 8811 76796 8853 76805
rect 11595 76796 11637 76805
rect 13498 76796 13556 76797
rect 8811 76756 8812 76796
rect 8852 76756 8853 76796
rect 8811 76747 8853 76756
rect 9387 76787 9429 76796
rect 9387 76747 9388 76787
rect 9428 76747 9429 76787
rect 4683 76738 4725 76747
rect 7851 76738 7893 76747
rect 9387 76738 9429 76747
rect 9867 76787 9909 76796
rect 9867 76747 9868 76787
rect 9908 76747 9909 76787
rect 11595 76756 11596 76796
rect 11636 76756 11637 76796
rect 11595 76747 11637 76756
rect 12843 76787 12885 76796
rect 12843 76747 12844 76787
rect 12884 76747 12885 76787
rect 13498 76756 13507 76796
rect 13547 76756 13556 76796
rect 13498 76755 13556 76756
rect 13611 76796 13653 76805
rect 13611 76756 13612 76796
rect 13652 76756 13653 76796
rect 13611 76747 13653 76756
rect 13995 76796 14037 76805
rect 16203 76796 16245 76805
rect 18219 76796 18261 76805
rect 19851 76796 19893 76805
rect 13995 76756 13996 76796
rect 14036 76756 14037 76796
rect 13995 76747 14037 76756
rect 14571 76787 14613 76796
rect 14571 76747 14572 76787
rect 14612 76747 14613 76787
rect 9867 76738 9909 76747
rect 12843 76738 12885 76747
rect 14571 76738 14613 76747
rect 15051 76787 15093 76796
rect 15051 76747 15052 76787
rect 15092 76747 15093 76787
rect 16203 76756 16204 76796
rect 16244 76756 16245 76796
rect 16203 76747 16245 76756
rect 17451 76787 17493 76796
rect 17451 76747 17452 76787
rect 17492 76747 17493 76787
rect 18219 76756 18220 76796
rect 18260 76756 18261 76796
rect 18219 76747 18261 76756
rect 19467 76787 19509 76796
rect 19467 76747 19468 76787
rect 19508 76747 19509 76787
rect 19851 76756 19852 76796
rect 19892 76756 19893 76796
rect 19851 76747 19893 76756
rect 15051 76738 15093 76747
rect 17451 76738 17493 76747
rect 19467 76738 19509 76747
rect 3723 76712 3765 76721
rect 3723 76672 3724 76712
rect 3764 76672 3765 76712
rect 3723 76663 3765 76672
rect 5067 76712 5109 76721
rect 5067 76672 5068 76712
rect 5108 76672 5109 76712
rect 5067 76663 5109 76672
rect 5643 76712 5685 76721
rect 5643 76672 5644 76712
rect 5684 76672 5685 76712
rect 5643 76663 5685 76672
rect 8907 76712 8949 76721
rect 8907 76672 8908 76712
rect 8948 76672 8949 76712
rect 8907 76663 8949 76672
rect 10090 76712 10148 76713
rect 10090 76672 10099 76712
rect 10139 76672 10148 76712
rect 10090 76671 10148 76672
rect 10443 76712 10485 76721
rect 10443 76672 10444 76712
rect 10484 76672 10485 76712
rect 10443 76663 10485 76672
rect 10587 76712 10629 76721
rect 10587 76672 10588 76712
rect 10628 76672 10629 76712
rect 10587 76663 10629 76672
rect 11211 76712 11253 76721
rect 11211 76672 11212 76712
rect 11252 76672 11253 76712
rect 11211 76663 11253 76672
rect 14091 76712 14133 76721
rect 14091 76672 14092 76712
rect 14132 76672 14133 76712
rect 14091 76663 14133 76672
rect 15435 76712 15477 76721
rect 15435 76672 15436 76712
rect 15476 76672 15477 76712
rect 15435 76663 15477 76672
rect 16011 76712 16053 76721
rect 16011 76672 16012 76712
rect 16052 76672 16053 76712
rect 16011 76663 16053 76672
rect 17835 76712 17877 76721
rect 17835 76672 17836 76712
rect 17876 76672 17877 76712
rect 17835 76663 17877 76672
rect 20139 76712 20181 76721
rect 20139 76672 20140 76712
rect 20180 76672 20181 76712
rect 20139 76663 20181 76672
rect 20379 76712 20421 76721
rect 20379 76672 20380 76712
rect 20420 76672 20421 76712
rect 20379 76663 20421 76672
rect 5403 76628 5445 76637
rect 5403 76588 5404 76628
rect 5444 76588 5445 76628
rect 5403 76579 5445 76588
rect 8043 76628 8085 76637
rect 8043 76588 8044 76628
rect 8084 76588 8085 76628
rect 8043 76579 8085 76588
rect 10875 76628 10917 76637
rect 10875 76588 10876 76628
rect 10916 76588 10917 76628
rect 10875 76579 10917 76588
rect 18075 76628 18117 76637
rect 18075 76588 18076 76628
rect 18116 76588 18117 76628
rect 18075 76579 18117 76588
rect 2859 76544 2901 76553
rect 2859 76504 2860 76544
rect 2900 76504 2901 76544
rect 2859 76495 2901 76504
rect 5307 76544 5349 76553
rect 5307 76504 5308 76544
rect 5348 76504 5349 76544
rect 5307 76495 5349 76504
rect 6411 76544 6453 76553
rect 6411 76504 6412 76544
rect 6452 76504 6453 76544
rect 6411 76495 6453 76504
rect 17643 76544 17685 76553
rect 17643 76504 17644 76544
rect 17684 76504 17685 76544
rect 17643 76495 17685 76504
rect 19659 76544 19701 76553
rect 19659 76504 19660 76544
rect 19700 76504 19701 76544
rect 19659 76495 19701 76504
rect 1152 76376 20448 76400
rect 1152 76336 3688 76376
rect 3728 76336 3770 76376
rect 3810 76336 3852 76376
rect 3892 76336 3934 76376
rect 3974 76336 4016 76376
rect 4056 76336 18808 76376
rect 18848 76336 18890 76376
rect 18930 76336 18972 76376
rect 19012 76336 19054 76376
rect 19094 76336 19136 76376
rect 19176 76336 20448 76376
rect 1152 76312 20448 76336
rect 5979 76208 6021 76217
rect 5979 76168 5980 76208
rect 6020 76168 6021 76208
rect 5979 76159 6021 76168
rect 8331 76208 8373 76217
rect 8331 76168 8332 76208
rect 8372 76168 8373 76208
rect 8331 76159 8373 76168
rect 9963 76208 10005 76217
rect 9963 76168 9964 76208
rect 10004 76168 10005 76208
rect 9963 76159 10005 76168
rect 11931 76208 11973 76217
rect 11931 76168 11932 76208
rect 11972 76168 11973 76208
rect 11931 76159 11973 76168
rect 18363 76208 18405 76217
rect 18363 76168 18364 76208
rect 18404 76168 18405 76208
rect 18363 76159 18405 76168
rect 11691 76124 11733 76133
rect 11691 76084 11692 76124
rect 11732 76084 11733 76124
rect 11691 76075 11733 76084
rect 2859 76040 2901 76049
rect 2859 76000 2860 76040
rect 2900 76000 2901 76040
rect 2859 75991 2901 76000
rect 3915 76040 3957 76049
rect 3915 76000 3916 76040
rect 3956 76000 3957 76040
rect 3915 75991 3957 76000
rect 5547 76040 5589 76049
rect 5547 76000 5548 76040
rect 5588 76000 5589 76040
rect 5547 75991 5589 76000
rect 5739 76040 5781 76049
rect 5739 76000 5740 76040
rect 5780 76000 5781 76040
rect 5739 75991 5781 76000
rect 6123 76040 6165 76049
rect 6123 76000 6124 76040
rect 6164 76000 6165 76040
rect 6123 75991 6165 76000
rect 6507 76040 6549 76049
rect 6507 76000 6508 76040
rect 6548 76000 6549 76040
rect 6507 75991 6549 76000
rect 13131 76040 13173 76049
rect 13131 76000 13132 76040
rect 13172 76000 13173 76040
rect 13131 75991 13173 76000
rect 18123 76040 18165 76049
rect 18123 76000 18124 76040
rect 18164 76000 18165 76040
rect 18123 75991 18165 76000
rect 20139 76040 20181 76049
rect 20139 76000 20140 76040
rect 20180 76000 20181 76040
rect 20139 75991 20181 76000
rect 1227 75956 1269 75965
rect 1227 75916 1228 75956
rect 1268 75916 1269 75956
rect 1227 75907 1269 75916
rect 2467 75956 2525 75957
rect 2467 75916 2476 75956
rect 2516 75916 2525 75956
rect 2467 75915 2525 75916
rect 3405 75956 3447 75965
rect 3405 75916 3406 75956
rect 3446 75916 3447 75956
rect 3405 75907 3447 75916
rect 3531 75956 3573 75965
rect 3531 75916 3532 75956
rect 3572 75916 3573 75956
rect 3531 75907 3573 75916
rect 4011 75956 4053 75965
rect 4011 75916 4012 75956
rect 4052 75916 4053 75956
rect 4011 75907 4053 75916
rect 4483 75956 4541 75957
rect 4483 75916 4492 75956
rect 4532 75916 4541 75956
rect 4483 75915 4541 75916
rect 5002 75956 5060 75957
rect 5002 75916 5011 75956
rect 5051 75916 5060 75956
rect 5002 75915 5060 75916
rect 6891 75956 6933 75965
rect 6891 75916 6892 75956
rect 6932 75916 6933 75956
rect 6891 75907 6933 75916
rect 8131 75956 8189 75957
rect 8131 75916 8140 75956
rect 8180 75916 8189 75956
rect 8131 75915 8189 75916
rect 8523 75956 8565 75965
rect 8523 75916 8524 75956
rect 8564 75916 8565 75956
rect 8523 75907 8565 75916
rect 9763 75956 9821 75957
rect 9763 75916 9772 75956
rect 9812 75916 9821 75956
rect 9763 75915 9821 75916
rect 10251 75956 10293 75965
rect 10251 75916 10252 75956
rect 10292 75916 10293 75956
rect 10251 75907 10293 75916
rect 11491 75956 11549 75957
rect 11491 75916 11500 75956
rect 11540 75916 11549 75956
rect 11491 75915 11549 75916
rect 12154 75956 12212 75957
rect 12154 75916 12163 75956
rect 12203 75916 12212 75956
rect 12154 75915 12212 75916
rect 12648 75956 12706 75957
rect 12648 75916 12657 75956
rect 12697 75916 12706 75956
rect 12648 75915 12706 75916
rect 13227 75956 13269 75965
rect 13227 75916 13228 75956
rect 13268 75916 13269 75956
rect 13227 75907 13269 75916
rect 13611 75956 13653 75965
rect 13611 75916 13612 75956
rect 13652 75916 13653 75956
rect 13611 75907 13653 75916
rect 13724 75956 13766 75965
rect 13724 75916 13725 75956
rect 13765 75916 13766 75956
rect 13724 75907 13766 75916
rect 14091 75956 14133 75965
rect 14091 75916 14092 75956
rect 14132 75916 14133 75956
rect 14091 75907 14133 75916
rect 15331 75956 15389 75957
rect 15331 75916 15340 75956
rect 15380 75916 15389 75956
rect 15331 75915 15389 75916
rect 15723 75956 15765 75965
rect 15723 75916 15724 75956
rect 15764 75916 15765 75956
rect 15723 75907 15765 75916
rect 16963 75956 17021 75957
rect 16963 75916 16972 75956
rect 17012 75916 17021 75956
rect 16963 75915 17021 75916
rect 17338 75956 17396 75957
rect 17338 75916 17347 75956
rect 17387 75916 17396 75956
rect 17338 75915 17396 75916
rect 17482 75956 17540 75957
rect 17482 75916 17491 75956
rect 17531 75916 17540 75956
rect 17482 75915 17540 75916
rect 17622 75956 17680 75957
rect 17622 75916 17631 75956
rect 17671 75916 17680 75956
rect 17622 75915 17680 75916
rect 17722 75956 17780 75957
rect 17722 75916 17731 75956
rect 17771 75916 17780 75956
rect 17722 75915 17780 75916
rect 17856 75956 17914 75957
rect 17856 75916 17865 75956
rect 17905 75916 17914 75956
rect 17856 75915 17914 75916
rect 18507 75956 18549 75965
rect 18507 75916 18508 75956
rect 18548 75916 18549 75956
rect 18507 75907 18549 75916
rect 19747 75956 19805 75957
rect 19747 75916 19756 75956
rect 19796 75916 19805 75956
rect 19747 75915 19805 75916
rect 2667 75788 2709 75797
rect 2667 75748 2668 75788
rect 2708 75748 2709 75788
rect 2667 75739 2709 75748
rect 3099 75788 3141 75797
rect 3099 75748 3100 75788
rect 3140 75748 3141 75788
rect 3099 75739 3141 75748
rect 5163 75788 5205 75797
rect 5163 75748 5164 75788
rect 5204 75748 5205 75788
rect 5163 75739 5205 75748
rect 5307 75788 5349 75797
rect 5307 75748 5308 75788
rect 5348 75748 5349 75788
rect 5307 75739 5349 75748
rect 6363 75788 6405 75797
rect 6363 75748 6364 75788
rect 6404 75748 6405 75788
rect 6363 75739 6405 75748
rect 6747 75788 6789 75797
rect 6747 75748 6748 75788
rect 6788 75748 6789 75788
rect 6747 75739 6789 75748
rect 15531 75788 15573 75797
rect 15531 75748 15532 75788
rect 15572 75748 15573 75788
rect 15531 75739 15573 75748
rect 17163 75788 17205 75797
rect 17163 75748 17164 75788
rect 17204 75748 17205 75788
rect 17163 75739 17205 75748
rect 17547 75788 17589 75797
rect 17547 75748 17548 75788
rect 17588 75748 17589 75788
rect 17547 75739 17589 75748
rect 19947 75788 19989 75797
rect 19947 75748 19948 75788
rect 19988 75748 19989 75788
rect 19947 75739 19989 75748
rect 20379 75788 20421 75797
rect 20379 75748 20380 75788
rect 20420 75748 20421 75788
rect 20379 75739 20421 75748
rect 1152 75620 20452 75644
rect 1152 75580 4928 75620
rect 4968 75580 5010 75620
rect 5050 75580 5092 75620
rect 5132 75580 5174 75620
rect 5214 75580 5256 75620
rect 5296 75580 20048 75620
rect 20088 75580 20130 75620
rect 20170 75580 20212 75620
rect 20252 75580 20294 75620
rect 20334 75580 20376 75620
rect 20416 75580 20452 75620
rect 1152 75556 20452 75580
rect 2235 75452 2277 75461
rect 2235 75412 2236 75452
rect 2276 75412 2277 75452
rect 2235 75403 2277 75412
rect 9003 75452 9045 75461
rect 9003 75412 9004 75452
rect 9044 75412 9045 75452
rect 9003 75403 9045 75412
rect 11163 75452 11205 75461
rect 11163 75412 11164 75452
rect 11204 75412 11205 75452
rect 11163 75403 11205 75412
rect 14043 75452 14085 75461
rect 14043 75412 14044 75452
rect 14084 75412 14085 75452
rect 14043 75403 14085 75412
rect 16683 75452 16725 75461
rect 16683 75412 16684 75452
rect 16724 75412 16725 75452
rect 16683 75403 16725 75412
rect 10731 75368 10773 75377
rect 10731 75328 10732 75368
rect 10772 75328 10773 75368
rect 10731 75319 10773 75328
rect 2667 75284 2709 75293
rect 4683 75284 4725 75293
rect 6315 75284 6357 75293
rect 7930 75284 7988 75285
rect 8353 75284 8411 75285
rect 2667 75244 2668 75284
rect 2708 75244 2709 75284
rect 2667 75235 2709 75244
rect 3915 75275 3957 75284
rect 3915 75235 3916 75275
rect 3956 75235 3957 75275
rect 4683 75244 4684 75284
rect 4724 75244 4725 75284
rect 4683 75235 4725 75244
rect 5931 75275 5973 75284
rect 5931 75235 5932 75275
rect 5972 75235 5973 75275
rect 6315 75244 6316 75284
rect 6356 75244 6357 75284
rect 6315 75235 6357 75244
rect 7563 75275 7605 75284
rect 7563 75235 7564 75275
rect 7604 75235 7605 75275
rect 7930 75244 7939 75284
rect 7979 75244 7988 75284
rect 7930 75243 7988 75244
rect 8043 75275 8085 75284
rect 3915 75226 3957 75235
rect 5931 75226 5973 75235
rect 7563 75226 7605 75235
rect 8043 75235 8044 75275
rect 8084 75235 8085 75275
rect 8043 75226 8085 75235
rect 8187 75275 8229 75284
rect 8187 75235 8188 75275
rect 8228 75235 8229 75275
rect 8353 75244 8362 75284
rect 8402 75244 8411 75284
rect 8353 75243 8411 75244
rect 8491 75284 8549 75285
rect 8491 75244 8500 75284
rect 8540 75244 8549 75284
rect 8491 75243 8549 75244
rect 8715 75284 8757 75293
rect 8715 75244 8716 75284
rect 8756 75244 8757 75284
rect 8715 75235 8757 75244
rect 8849 75284 8907 75285
rect 8849 75244 8858 75284
rect 8898 75244 8907 75284
rect 8849 75243 8907 75244
rect 9291 75284 9333 75293
rect 14938 75284 14996 75285
rect 9291 75244 9292 75284
rect 9332 75244 9333 75284
rect 9291 75235 9333 75244
rect 10539 75275 10581 75284
rect 10539 75235 10540 75275
rect 10580 75235 10581 75275
rect 14938 75244 14947 75284
rect 14987 75244 14996 75284
rect 14938 75243 14996 75244
rect 15051 75284 15093 75293
rect 15051 75244 15052 75284
rect 15092 75244 15093 75284
rect 15051 75235 15093 75244
rect 15435 75284 15477 75293
rect 16875 75284 16917 75293
rect 18891 75284 18933 75293
rect 15435 75244 15436 75284
rect 15476 75244 15477 75284
rect 15435 75235 15477 75244
rect 16011 75275 16053 75284
rect 16011 75235 16012 75275
rect 16052 75235 16053 75275
rect 8187 75226 8229 75235
rect 10539 75226 10581 75235
rect 16011 75226 16053 75235
rect 16491 75275 16533 75284
rect 16491 75235 16492 75275
rect 16532 75235 16533 75275
rect 16875 75244 16876 75284
rect 16916 75244 16917 75284
rect 16875 75235 16917 75244
rect 18123 75275 18165 75284
rect 18123 75235 18124 75275
rect 18164 75235 18165 75275
rect 18891 75244 18892 75284
rect 18932 75244 18933 75284
rect 18891 75235 18933 75244
rect 20139 75275 20181 75284
rect 20139 75235 20140 75275
rect 20180 75235 20181 75275
rect 16491 75226 16533 75235
rect 18123 75226 18165 75235
rect 20139 75226 20181 75235
rect 1227 75200 1269 75209
rect 1227 75160 1228 75200
rect 1268 75160 1269 75200
rect 1227 75151 1269 75160
rect 1611 75200 1653 75209
rect 1611 75160 1612 75200
rect 1652 75160 1653 75200
rect 1611 75151 1653 75160
rect 1995 75200 2037 75209
rect 1995 75160 1996 75200
rect 2036 75160 2037 75200
rect 1995 75151 2037 75160
rect 4491 75200 4533 75209
rect 4491 75160 4492 75200
rect 4532 75160 4533 75200
rect 4491 75151 4533 75160
rect 10923 75200 10965 75209
rect 10923 75160 10924 75200
rect 10964 75160 10965 75200
rect 10923 75151 10965 75160
rect 12747 75200 12789 75209
rect 12747 75160 12748 75200
rect 12788 75160 12789 75200
rect 12747 75151 12789 75160
rect 12939 75200 12981 75209
rect 12939 75160 12940 75200
rect 12980 75160 12981 75200
rect 12939 75151 12981 75160
rect 13179 75200 13221 75209
rect 13179 75160 13180 75200
rect 13220 75160 13221 75200
rect 13179 75151 13221 75160
rect 13323 75200 13365 75209
rect 13323 75160 13324 75200
rect 13364 75160 13365 75200
rect 13323 75151 13365 75160
rect 13707 75200 13749 75209
rect 13707 75160 13708 75200
rect 13748 75160 13749 75200
rect 13707 75151 13749 75160
rect 14283 75200 14325 75209
rect 14283 75160 14284 75200
rect 14324 75160 14325 75200
rect 14283 75151 14325 75160
rect 14475 75200 14517 75209
rect 14475 75160 14476 75200
rect 14516 75160 14517 75200
rect 14475 75151 14517 75160
rect 15531 75200 15573 75209
rect 15531 75160 15532 75200
rect 15572 75160 15573 75200
rect 15531 75151 15573 75160
rect 18507 75200 18549 75209
rect 18507 75160 18508 75200
rect 18548 75160 18549 75200
rect 18507 75151 18549 75160
rect 4251 75116 4293 75125
rect 4251 75076 4252 75116
rect 4292 75076 4293 75116
rect 4251 75067 4293 75076
rect 13563 75116 13605 75125
rect 13563 75076 13564 75116
rect 13604 75076 13605 75116
rect 13563 75067 13605 75076
rect 13947 75116 13989 75125
rect 13947 75076 13948 75116
rect 13988 75076 13989 75116
rect 13947 75067 13989 75076
rect 1467 75032 1509 75041
rect 1467 74992 1468 75032
rect 1508 74992 1509 75032
rect 1467 74983 1509 74992
rect 1851 75032 1893 75041
rect 1851 74992 1852 75032
rect 1892 74992 1893 75032
rect 1851 74983 1893 74992
rect 4107 75032 4149 75041
rect 4107 74992 4108 75032
rect 4148 74992 4149 75032
rect 4107 74983 4149 74992
rect 6123 75032 6165 75041
rect 6123 74992 6124 75032
rect 6164 74992 6165 75032
rect 6123 74983 6165 74992
rect 7755 75032 7797 75041
rect 7755 74992 7756 75032
rect 7796 74992 7797 75032
rect 7755 74983 7797 74992
rect 7930 75032 7988 75033
rect 7930 74992 7939 75032
rect 7979 74992 7988 75032
rect 7930 74991 7988 74992
rect 12507 75032 12549 75041
rect 12507 74992 12508 75032
rect 12548 74992 12549 75032
rect 12507 74983 12549 74992
rect 14715 75032 14757 75041
rect 14715 74992 14716 75032
rect 14756 74992 14757 75032
rect 14715 74983 14757 74992
rect 18315 75032 18357 75041
rect 18315 74992 18316 75032
rect 18356 74992 18357 75032
rect 18315 74983 18357 74992
rect 18747 75032 18789 75041
rect 18747 74992 18748 75032
rect 18788 74992 18789 75032
rect 18747 74983 18789 74992
rect 20331 75032 20373 75041
rect 20331 74992 20332 75032
rect 20372 74992 20373 75032
rect 20331 74983 20373 74992
rect 1152 74864 20448 74888
rect 1152 74824 3688 74864
rect 3728 74824 3770 74864
rect 3810 74824 3852 74864
rect 3892 74824 3934 74864
rect 3974 74824 4016 74864
rect 4056 74824 18808 74864
rect 18848 74824 18890 74864
rect 18930 74824 18972 74864
rect 19012 74824 19054 74864
rect 19094 74824 19136 74864
rect 19176 74824 20448 74864
rect 1152 74800 20448 74824
rect 5499 74696 5541 74705
rect 5499 74656 5500 74696
rect 5540 74656 5541 74696
rect 5499 74647 5541 74656
rect 11691 74696 11733 74705
rect 11691 74656 11692 74696
rect 11732 74656 11733 74696
rect 11691 74647 11733 74656
rect 17355 74696 17397 74705
rect 17355 74656 17356 74696
rect 17396 74656 17397 74696
rect 17355 74647 17397 74656
rect 17691 74696 17733 74705
rect 17691 74656 17692 74696
rect 17732 74656 17733 74696
rect 17691 74647 17733 74656
rect 10059 74612 10101 74621
rect 10059 74572 10060 74612
rect 10100 74572 10101 74612
rect 10059 74563 10101 74572
rect 2859 74528 2901 74537
rect 2859 74488 2860 74528
rect 2900 74488 2901 74528
rect 2859 74479 2901 74488
rect 3915 74528 3957 74537
rect 3915 74488 3916 74528
rect 3956 74488 3957 74528
rect 3915 74479 3957 74488
rect 6219 74528 6261 74537
rect 6219 74488 6220 74528
rect 6260 74488 6261 74528
rect 6219 74479 6261 74488
rect 7851 74528 7893 74537
rect 7851 74488 7852 74528
rect 7892 74488 7893 74528
rect 7851 74479 7893 74488
rect 8427 74528 8469 74537
rect 8427 74488 8428 74528
rect 8468 74488 8469 74528
rect 8427 74479 8469 74488
rect 13611 74528 13653 74537
rect 13611 74488 13612 74528
rect 13652 74488 13653 74528
rect 13611 74479 13653 74488
rect 14859 74528 14901 74537
rect 14859 74488 14860 74528
rect 14900 74488 14901 74528
rect 14859 74479 14901 74488
rect 18411 74528 18453 74537
rect 18411 74488 18412 74528
rect 18452 74488 18453 74528
rect 18411 74479 18453 74488
rect 20139 74528 20181 74537
rect 20139 74488 20140 74528
rect 20180 74488 20181 74528
rect 20139 74479 20181 74488
rect 17058 74470 17104 74479
rect 1227 74444 1269 74453
rect 1227 74404 1228 74444
rect 1268 74404 1269 74444
rect 1227 74395 1269 74404
rect 2467 74444 2525 74445
rect 2467 74404 2476 74444
rect 2516 74404 2525 74444
rect 2467 74403 2525 74404
rect 3418 74444 3476 74445
rect 3418 74404 3427 74444
rect 3467 74404 3476 74444
rect 3418 74403 3476 74404
rect 3531 74444 3573 74453
rect 3531 74404 3532 74444
rect 3572 74404 3573 74444
rect 3531 74395 3573 74404
rect 4011 74444 4053 74453
rect 4011 74404 4012 74444
rect 4052 74404 4053 74444
rect 4011 74395 4053 74404
rect 4483 74444 4541 74445
rect 4483 74404 4492 74444
rect 4532 74404 4541 74444
rect 4483 74403 4541 74404
rect 5002 74444 5060 74445
rect 5002 74404 5011 74444
rect 5051 74404 5060 74444
rect 5002 74403 5060 74404
rect 5355 74444 5397 74453
rect 5355 74404 5356 74444
rect 5396 74404 5397 74444
rect 5355 74395 5397 74404
rect 5722 74444 5780 74445
rect 5722 74404 5731 74444
rect 5771 74404 5780 74444
rect 5722 74403 5780 74404
rect 5835 74444 5877 74453
rect 5835 74404 5836 74444
rect 5876 74404 5877 74444
rect 5835 74395 5877 74404
rect 6315 74444 6357 74453
rect 6315 74404 6316 74444
rect 6356 74404 6357 74444
rect 6315 74395 6357 74404
rect 6787 74444 6845 74445
rect 6787 74404 6796 74444
rect 6836 74404 6845 74444
rect 6787 74403 6845 74404
rect 7275 74444 7333 74445
rect 7275 74404 7284 74444
rect 7324 74404 7333 74444
rect 7275 74403 7333 74404
rect 8619 74444 8661 74453
rect 8619 74404 8620 74444
rect 8660 74404 8661 74444
rect 8619 74395 8661 74404
rect 9859 74444 9917 74445
rect 9859 74404 9868 74444
rect 9908 74404 9917 74444
rect 9859 74403 9917 74404
rect 10251 74444 10293 74453
rect 10251 74404 10252 74444
rect 10292 74404 10293 74444
rect 10251 74395 10293 74404
rect 11491 74444 11549 74445
rect 11491 74404 11500 74444
rect 11540 74404 11549 74444
rect 11491 74403 11549 74404
rect 11979 74444 12021 74453
rect 11979 74404 11980 74444
rect 12020 74404 12021 74444
rect 11979 74395 12021 74404
rect 13219 74444 13277 74445
rect 13219 74404 13228 74444
rect 13268 74404 13277 74444
rect 13219 74403 13277 74404
rect 14362 74444 14420 74445
rect 14362 74404 14371 74444
rect 14411 74404 14420 74444
rect 14362 74403 14420 74404
rect 14475 74444 14517 74453
rect 14475 74404 14476 74444
rect 14516 74404 14517 74444
rect 14475 74395 14517 74404
rect 14955 74444 14997 74453
rect 14955 74404 14956 74444
rect 14996 74404 14997 74444
rect 14955 74395 14997 74404
rect 15427 74444 15485 74445
rect 15427 74404 15436 74444
rect 15476 74404 15485 74444
rect 15427 74403 15485 74404
rect 15915 74444 15973 74445
rect 15915 74404 15924 74444
rect 15964 74404 15973 74444
rect 15915 74403 15973 74404
rect 16731 74444 16773 74453
rect 16731 74404 16732 74444
rect 16772 74404 16773 74444
rect 16731 74395 16773 74404
rect 16875 74444 16917 74453
rect 16875 74404 16876 74444
rect 16916 74404 16917 74444
rect 17058 74430 17059 74470
rect 17099 74430 17104 74470
rect 17058 74421 17104 74430
rect 17242 74444 17300 74445
rect 16875 74395 16917 74404
rect 17242 74404 17251 74444
rect 17291 74404 17300 74444
rect 17242 74403 17300 74404
rect 17355 74444 17397 74453
rect 17355 74404 17356 74444
rect 17396 74404 17397 74444
rect 17355 74395 17397 74404
rect 17547 74444 17589 74453
rect 17547 74404 17548 74444
rect 17588 74404 17589 74444
rect 17547 74395 17589 74404
rect 17914 74444 17972 74445
rect 17914 74404 17923 74444
rect 17963 74404 17972 74444
rect 17914 74403 17972 74404
rect 18027 74444 18069 74453
rect 18027 74404 18028 74444
rect 18068 74404 18069 74444
rect 18027 74395 18069 74404
rect 18507 74444 18549 74453
rect 18507 74404 18508 74444
rect 18548 74404 18549 74444
rect 18507 74395 18549 74404
rect 18979 74444 19037 74445
rect 18979 74404 18988 74444
rect 19028 74404 19037 74444
rect 18979 74403 19037 74404
rect 19498 74444 19556 74445
rect 19498 74404 19507 74444
rect 19547 74404 19556 74444
rect 19498 74403 19556 74404
rect 8091 74360 8133 74369
rect 8091 74320 8092 74360
rect 8132 74320 8133 74360
rect 8091 74311 8133 74320
rect 13851 74360 13893 74369
rect 13851 74320 13852 74360
rect 13892 74320 13893 74360
rect 13851 74311 13893 74320
rect 2667 74276 2709 74285
rect 2667 74236 2668 74276
rect 2708 74236 2709 74276
rect 2667 74227 2709 74236
rect 3099 74276 3141 74285
rect 3099 74236 3100 74276
rect 3140 74236 3141 74276
rect 3099 74227 3141 74236
rect 5163 74276 5205 74285
rect 5163 74236 5164 74276
rect 5204 74236 5205 74276
rect 5163 74227 5205 74236
rect 7467 74276 7509 74285
rect 7467 74236 7468 74276
rect 7508 74236 7509 74276
rect 7467 74227 7509 74236
rect 8187 74276 8229 74285
rect 8187 74236 8188 74276
rect 8228 74236 8229 74276
rect 8187 74227 8229 74236
rect 13419 74276 13461 74285
rect 13419 74236 13420 74276
rect 13460 74236 13461 74276
rect 13419 74227 13461 74236
rect 16107 74276 16149 74285
rect 16107 74236 16108 74276
rect 16148 74236 16149 74276
rect 16107 74227 16149 74236
rect 16570 74276 16628 74277
rect 16570 74236 16579 74276
rect 16619 74236 16628 74276
rect 16570 74235 16628 74236
rect 19659 74276 19701 74285
rect 19659 74236 19660 74276
rect 19700 74236 19701 74276
rect 19659 74227 19701 74236
rect 20379 74276 20421 74285
rect 20379 74236 20380 74276
rect 20420 74236 20421 74276
rect 20379 74227 20421 74236
rect 1152 74108 20452 74132
rect 1152 74068 4928 74108
rect 4968 74068 5010 74108
rect 5050 74068 5092 74108
rect 5132 74068 5174 74108
rect 5214 74068 5256 74108
rect 5296 74068 20048 74108
rect 20088 74068 20130 74108
rect 20170 74068 20212 74108
rect 20252 74068 20294 74108
rect 20334 74068 20376 74108
rect 20416 74068 20452 74108
rect 1152 74044 20452 74068
rect 4779 73940 4821 73949
rect 4779 73900 4780 73940
rect 4820 73900 4821 73940
rect 4779 73891 4821 73900
rect 6603 73940 6645 73949
rect 6603 73900 6604 73940
rect 6644 73900 6645 73940
rect 6603 73891 6645 73900
rect 12219 73940 12261 73949
rect 12219 73900 12220 73940
rect 12260 73900 12261 73940
rect 12219 73891 12261 73900
rect 14475 73940 14517 73949
rect 14475 73900 14476 73940
rect 14516 73900 14517 73940
rect 14475 73891 14517 73900
rect 12075 73856 12117 73865
rect 12075 73816 12076 73856
rect 12116 73816 12117 73856
rect 12075 73807 12117 73816
rect 1323 73772 1365 73781
rect 3034 73772 3092 73773
rect 1323 73732 1324 73772
rect 1364 73732 1365 73772
rect 1323 73723 1365 73732
rect 2571 73763 2613 73772
rect 2571 73723 2572 73763
rect 2612 73723 2613 73763
rect 3034 73732 3043 73772
rect 3083 73732 3092 73772
rect 3034 73731 3092 73732
rect 3147 73772 3189 73781
rect 3147 73732 3148 73772
rect 3188 73732 3189 73772
rect 3147 73723 3189 73732
rect 3531 73772 3573 73781
rect 5163 73772 5205 73781
rect 6970 73772 7028 73773
rect 7947 73772 7989 73781
rect 3531 73732 3532 73772
rect 3572 73732 3573 73772
rect 3531 73723 3573 73732
rect 4107 73763 4149 73772
rect 4107 73723 4108 73763
rect 4148 73723 4149 73763
rect 2571 73714 2613 73723
rect 4107 73714 4149 73723
rect 4587 73763 4629 73772
rect 4587 73723 4588 73763
rect 4628 73723 4629 73763
rect 5163 73732 5164 73772
rect 5204 73732 5205 73772
rect 5163 73723 5205 73732
rect 6411 73763 6453 73772
rect 6411 73723 6412 73763
rect 6452 73723 6453 73763
rect 6970 73732 6979 73772
rect 7019 73732 7028 73772
rect 6970 73731 7028 73732
rect 7467 73763 7509 73772
rect 4587 73714 4629 73723
rect 6411 73714 6453 73723
rect 7467 73723 7468 73763
rect 7508 73723 7509 73763
rect 7947 73732 7948 73772
rect 7988 73732 7989 73772
rect 7947 73723 7989 73732
rect 8427 73772 8469 73781
rect 8427 73732 8428 73772
rect 8468 73732 8469 73772
rect 8427 73723 8469 73732
rect 8528 73772 8570 73781
rect 8528 73732 8529 73772
rect 8569 73732 8570 73772
rect 8528 73723 8570 73732
rect 8995 73772 9053 73773
rect 8995 73732 9004 73772
rect 9044 73732 9053 73772
rect 8995 73731 9053 73732
rect 10251 73772 10293 73781
rect 10251 73732 10252 73772
rect 10292 73732 10293 73772
rect 10251 73723 10293 73732
rect 10635 73772 10677 73781
rect 12730 73772 12788 73773
rect 10635 73732 10636 73772
rect 10676 73732 10677 73772
rect 10635 73723 10677 73732
rect 11883 73763 11925 73772
rect 11883 73723 11884 73763
rect 11924 73723 11925 73763
rect 12730 73732 12739 73772
rect 12779 73732 12788 73772
rect 12730 73731 12788 73732
rect 12843 73772 12885 73781
rect 12843 73732 12844 73772
rect 12884 73732 12885 73772
rect 12843 73723 12885 73732
rect 13227 73772 13269 73781
rect 16395 73772 16437 73781
rect 18603 73772 18645 73781
rect 20331 73772 20373 73781
rect 13227 73732 13228 73772
rect 13268 73732 13269 73772
rect 13227 73723 13269 73732
rect 13803 73763 13845 73772
rect 13803 73723 13804 73763
rect 13844 73723 13845 73763
rect 7467 73714 7509 73723
rect 11883 73714 11925 73723
rect 13803 73714 13845 73723
rect 14283 73763 14325 73772
rect 14283 73723 14284 73763
rect 14324 73723 14325 73763
rect 16395 73732 16396 73772
rect 16436 73732 16437 73772
rect 16395 73723 16437 73732
rect 17643 73763 17685 73772
rect 17643 73723 17644 73763
rect 17684 73723 17685 73763
rect 18603 73732 18604 73772
rect 18644 73732 18645 73772
rect 18603 73723 18645 73732
rect 19851 73763 19893 73772
rect 19851 73723 19852 73763
rect 19892 73723 19893 73763
rect 20331 73732 20332 73772
rect 20372 73732 20373 73772
rect 20331 73723 20373 73732
rect 14283 73714 14325 73723
rect 17643 73714 17685 73723
rect 19851 73714 19893 73723
rect 3627 73688 3669 73697
rect 3627 73648 3628 73688
rect 3668 73648 3669 73688
rect 3627 73639 3669 73648
rect 6747 73688 6789 73697
rect 6747 73648 6748 73688
rect 6788 73648 6789 73688
rect 6747 73639 6789 73648
rect 8043 73688 8085 73697
rect 8043 73648 8044 73688
rect 8084 73648 8085 73688
rect 8043 73639 8085 73648
rect 12459 73688 12501 73697
rect 12459 73648 12460 73688
rect 12500 73648 12501 73688
rect 12459 73639 12501 73648
rect 13323 73688 13365 73697
rect 13323 73648 13324 73688
rect 13364 73648 13365 73688
rect 13323 73639 13365 73648
rect 14859 73688 14901 73697
rect 14859 73648 14860 73688
rect 14900 73648 14901 73688
rect 14859 73639 14901 73648
rect 15099 73688 15141 73697
rect 15099 73648 15100 73688
rect 15140 73648 15141 73688
rect 15099 73639 15141 73648
rect 15483 73688 15525 73697
rect 15483 73648 15484 73688
rect 15524 73648 15525 73688
rect 15483 73639 15525 73648
rect 15723 73688 15765 73697
rect 15723 73648 15724 73688
rect 15764 73648 15765 73688
rect 15723 73639 15765 73648
rect 15915 73688 15957 73697
rect 15915 73648 15916 73688
rect 15956 73648 15957 73688
rect 15915 73639 15957 73648
rect 18219 73688 18261 73697
rect 18219 73648 18220 73688
rect 18260 73648 18261 73688
rect 18219 73639 18261 73648
rect 15387 73604 15429 73613
rect 15387 73564 15388 73604
rect 15428 73564 15429 73604
rect 15387 73555 15429 73564
rect 20187 73604 20229 73613
rect 20187 73564 20188 73604
rect 20228 73564 20229 73604
rect 20187 73555 20229 73564
rect 2763 73520 2805 73529
rect 2763 73480 2764 73520
rect 2804 73480 2805 73520
rect 2763 73471 2805 73480
rect 8811 73520 8853 73529
rect 8811 73480 8812 73520
rect 8852 73480 8853 73520
rect 8811 73471 8853 73480
rect 14619 73520 14661 73529
rect 14619 73480 14620 73520
rect 14660 73480 14661 73520
rect 14619 73471 14661 73480
rect 16155 73520 16197 73529
rect 16155 73480 16156 73520
rect 16196 73480 16197 73520
rect 16155 73471 16197 73480
rect 17835 73520 17877 73529
rect 17835 73480 17836 73520
rect 17876 73480 17877 73520
rect 17835 73471 17877 73480
rect 18459 73520 18501 73529
rect 18459 73480 18460 73520
rect 18500 73480 18501 73520
rect 18459 73471 18501 73480
rect 20043 73520 20085 73529
rect 20043 73480 20044 73520
rect 20084 73480 20085 73520
rect 20043 73471 20085 73480
rect 1152 73352 20448 73376
rect 1152 73312 3688 73352
rect 3728 73312 3770 73352
rect 3810 73312 3852 73352
rect 3892 73312 3934 73352
rect 3974 73312 4016 73352
rect 4056 73312 18808 73352
rect 18848 73312 18890 73352
rect 18930 73312 18972 73352
rect 19012 73312 19054 73352
rect 19094 73312 19136 73352
rect 19176 73312 20448 73352
rect 1152 73288 20448 73312
rect 4827 73184 4869 73193
rect 4827 73144 4828 73184
rect 4868 73144 4869 73184
rect 4827 73135 4869 73144
rect 6939 73184 6981 73193
rect 6939 73144 6940 73184
rect 6980 73144 6981 73184
rect 6939 73135 6981 73144
rect 17451 73184 17493 73193
rect 17451 73144 17452 73184
rect 17492 73144 17493 73184
rect 17451 73135 17493 73144
rect 19258 73184 19316 73185
rect 19258 73144 19267 73184
rect 19307 73144 19316 73184
rect 19258 73143 19316 73144
rect 15483 73100 15525 73109
rect 15483 73060 15484 73100
rect 15524 73060 15525 73100
rect 15483 73051 15525 73060
rect 19083 73100 19125 73109
rect 19083 73060 19084 73100
rect 19124 73060 19125 73100
rect 19083 73051 19125 73060
rect 4587 73016 4629 73025
rect 4587 72976 4588 73016
rect 4628 72976 4629 73016
rect 4587 72967 4629 72976
rect 6699 73016 6741 73025
rect 6699 72976 6700 73016
rect 6740 72976 6741 73016
rect 6699 72967 6741 72976
rect 8187 73016 8229 73025
rect 8187 72976 8188 73016
rect 8228 72976 8229 73016
rect 8187 72967 8229 72976
rect 8322 73016 8380 73017
rect 8322 72976 8331 73016
rect 8371 72976 8380 73016
rect 8322 72975 8380 72976
rect 13419 73016 13461 73025
rect 13419 72976 13420 73016
rect 13460 72976 13461 73016
rect 13419 72967 13461 72976
rect 14859 73016 14901 73025
rect 14859 72976 14860 73016
rect 14900 72976 14901 73016
rect 14859 72967 14901 72976
rect 15243 73016 15285 73025
rect 15243 72976 15244 73016
rect 15284 72976 15285 73016
rect 15243 72967 15285 72976
rect 15627 73016 15669 73025
rect 15627 72976 15628 73016
rect 15668 72976 15669 73016
rect 15627 72967 15669 72976
rect 20139 73016 20181 73025
rect 20139 72976 20140 73016
rect 20180 72976 20181 73016
rect 20139 72967 20181 72976
rect 19371 72943 19413 72952
rect 1323 72932 1365 72941
rect 1323 72892 1324 72932
rect 1364 72892 1365 72932
rect 1323 72883 1365 72892
rect 2563 72932 2621 72933
rect 2563 72892 2572 72932
rect 2612 72892 2621 72932
rect 2563 72891 2621 72892
rect 2955 72932 2997 72941
rect 2955 72892 2956 72932
rect 2996 72892 2997 72932
rect 2955 72883 2997 72892
rect 4195 72932 4253 72933
rect 4195 72892 4204 72932
rect 4244 72892 4253 72932
rect 4195 72891 4253 72892
rect 4971 72932 5013 72941
rect 4971 72892 4972 72932
rect 5012 72892 5013 72932
rect 4971 72883 5013 72892
rect 6211 72932 6269 72933
rect 6211 72892 6220 72932
rect 6260 72892 6269 72932
rect 6211 72891 6269 72892
rect 7258 72932 7316 72933
rect 7258 72892 7267 72932
rect 7307 72892 7316 72932
rect 7258 72891 7316 72892
rect 7747 72932 7805 72933
rect 7747 72892 7756 72932
rect 7796 72892 7805 72932
rect 7747 72891 7805 72892
rect 8715 72932 8757 72941
rect 8715 72892 8716 72932
rect 8756 72892 8757 72932
rect 8715 72883 8757 72892
rect 8825 72932 8883 72933
rect 8825 72892 8834 72932
rect 8874 72892 8883 72932
rect 8825 72891 8883 72892
rect 9571 72932 9629 72933
rect 9571 72892 9580 72932
rect 9620 72892 9629 72932
rect 9571 72891 9629 72892
rect 10827 72932 10869 72941
rect 10827 72892 10828 72932
rect 10868 72892 10869 72932
rect 10827 72883 10869 72892
rect 11019 72932 11061 72941
rect 11019 72892 11020 72932
rect 11060 72892 11061 72932
rect 11019 72883 11061 72892
rect 12259 72932 12317 72933
rect 12259 72892 12268 72932
rect 12308 72892 12317 72932
rect 12259 72891 12317 72892
rect 12922 72932 12980 72933
rect 12922 72892 12931 72932
rect 12971 72892 12980 72932
rect 12922 72891 12980 72892
rect 13035 72932 13077 72941
rect 13035 72892 13036 72932
rect 13076 72892 13077 72932
rect 13035 72883 13077 72892
rect 13515 72932 13557 72941
rect 13515 72892 13516 72932
rect 13556 72892 13557 72932
rect 13515 72883 13557 72892
rect 13987 72932 14045 72933
rect 13987 72892 13996 72932
rect 14036 72892 14045 72932
rect 13987 72891 14045 72892
rect 14506 72932 14564 72933
rect 14506 72892 14515 72932
rect 14555 72892 14564 72932
rect 14506 72891 14564 72892
rect 16011 72932 16053 72941
rect 16011 72892 16012 72932
rect 16052 72892 16053 72932
rect 16011 72883 16053 72892
rect 17251 72932 17309 72933
rect 17251 72892 17260 72932
rect 17300 72892 17309 72932
rect 17251 72891 17309 72892
rect 17643 72932 17685 72941
rect 17643 72892 17644 72932
rect 17684 72892 17685 72932
rect 17643 72883 17685 72892
rect 18883 72932 18941 72933
rect 18883 72892 18892 72932
rect 18932 72892 18941 72932
rect 18883 72891 18941 72892
rect 19258 72932 19316 72933
rect 19258 72892 19267 72932
rect 19307 72892 19316 72932
rect 19371 72903 19372 72943
rect 19412 72903 19413 72943
rect 19776 72943 19818 72952
rect 19371 72894 19413 72903
rect 19508 72932 19566 72933
rect 19258 72891 19316 72892
rect 19508 72892 19517 72932
rect 19557 72892 19566 72932
rect 19508 72891 19566 72892
rect 19638 72932 19696 72933
rect 19638 72892 19647 72932
rect 19687 72892 19696 72932
rect 19776 72903 19777 72943
rect 19817 72903 19818 72943
rect 19776 72894 19818 72903
rect 19638 72891 19696 72892
rect 7066 72848 7124 72849
rect 7066 72808 7075 72848
rect 7115 72808 7124 72848
rect 7066 72807 7124 72808
rect 12459 72848 12501 72857
rect 12459 72808 12460 72848
rect 12500 72808 12501 72848
rect 12459 72799 12501 72808
rect 15099 72848 15141 72857
rect 15099 72808 15100 72848
rect 15140 72808 15141 72848
rect 15099 72799 15141 72808
rect 2763 72764 2805 72773
rect 2763 72724 2764 72764
rect 2804 72724 2805 72764
rect 2763 72715 2805 72724
rect 4395 72764 4437 72773
rect 4395 72724 4396 72764
rect 4436 72724 4437 72764
rect 4395 72715 4437 72724
rect 6411 72764 6453 72773
rect 6411 72724 6412 72764
rect 6452 72724 6453 72764
rect 6411 72715 6453 72724
rect 9387 72764 9429 72773
rect 9387 72724 9388 72764
rect 9428 72724 9429 72764
rect 9387 72715 9429 72724
rect 14667 72764 14709 72773
rect 14667 72724 14668 72764
rect 14708 72724 14709 72764
rect 14667 72715 14709 72724
rect 15867 72764 15909 72773
rect 15867 72724 15868 72764
rect 15908 72724 15909 72764
rect 15867 72715 15909 72724
rect 17451 72764 17493 72773
rect 17451 72724 17452 72764
rect 17492 72724 17493 72764
rect 17451 72715 17493 72724
rect 19083 72764 19125 72773
rect 19083 72724 19084 72764
rect 19124 72724 19125 72764
rect 19083 72715 19125 72724
rect 20379 72764 20421 72773
rect 20379 72724 20380 72764
rect 20420 72724 20421 72764
rect 20379 72715 20421 72724
rect 1152 72596 20452 72620
rect 1152 72556 4928 72596
rect 4968 72556 5010 72596
rect 5050 72556 5092 72596
rect 5132 72556 5174 72596
rect 5214 72556 5256 72596
rect 5296 72556 20048 72596
rect 20088 72556 20130 72596
rect 20170 72556 20212 72596
rect 20252 72556 20294 72596
rect 20334 72556 20376 72596
rect 20416 72556 20452 72596
rect 1152 72532 20452 72556
rect 10491 72428 10533 72437
rect 10491 72388 10492 72428
rect 10532 72388 10533 72428
rect 10491 72379 10533 72388
rect 11259 72428 11301 72437
rect 11259 72388 11260 72428
rect 11300 72388 11301 72428
rect 11259 72379 11301 72388
rect 15051 72428 15093 72437
rect 15051 72388 15052 72428
rect 15092 72388 15093 72428
rect 15051 72379 15093 72388
rect 17146 72428 17204 72429
rect 17146 72388 17155 72428
rect 17195 72388 17204 72428
rect 17146 72387 17204 72388
rect 20139 72428 20181 72437
rect 20139 72388 20140 72428
rect 20180 72388 20181 72428
rect 20139 72379 20181 72388
rect 2331 72344 2373 72353
rect 2331 72304 2332 72344
rect 2372 72304 2373 72344
rect 2331 72295 2373 72304
rect 5115 72344 5157 72353
rect 5115 72304 5116 72344
rect 5156 72304 5157 72344
rect 5115 72295 5157 72304
rect 5499 72344 5541 72353
rect 5499 72304 5500 72344
rect 5540 72304 5541 72344
rect 5499 72295 5541 72304
rect 10107 72344 10149 72353
rect 10107 72304 10108 72344
rect 10148 72304 10149 72344
rect 10107 72295 10149 72304
rect 2842 72260 2900 72261
rect 2842 72220 2851 72260
rect 2891 72220 2900 72260
rect 2842 72219 2900 72220
rect 2955 72260 2997 72269
rect 2955 72220 2956 72260
rect 2996 72220 2997 72260
rect 2955 72211 2997 72220
rect 3339 72260 3381 72269
rect 4618 72260 4676 72261
rect 3339 72220 3340 72260
rect 3380 72220 3381 72260
rect 3339 72211 3381 72220
rect 3915 72251 3957 72260
rect 3915 72211 3916 72251
rect 3956 72211 3957 72251
rect 3915 72202 3957 72211
rect 4395 72251 4437 72260
rect 4395 72211 4396 72251
rect 4436 72211 4437 72251
rect 4618 72220 4627 72260
rect 4667 72220 4676 72260
rect 4618 72219 4676 72220
rect 6285 72260 6327 72269
rect 6285 72220 6286 72260
rect 6326 72220 6327 72260
rect 6285 72211 6327 72220
rect 6411 72260 6453 72269
rect 6411 72220 6412 72260
rect 6452 72220 6453 72260
rect 6411 72211 6453 72220
rect 6795 72260 6837 72269
rect 11979 72260 12021 72269
rect 13611 72260 13653 72269
rect 15243 72260 15285 72269
rect 17307 72260 17349 72269
rect 6795 72220 6796 72260
rect 6836 72220 6837 72260
rect 6795 72211 6837 72220
rect 7371 72251 7413 72260
rect 7371 72211 7372 72251
rect 7412 72211 7413 72251
rect 4395 72202 4437 72211
rect 7371 72202 7413 72211
rect 7851 72251 7893 72260
rect 7851 72211 7852 72251
rect 7892 72211 7893 72251
rect 11979 72220 11980 72260
rect 12020 72220 12021 72260
rect 11979 72211 12021 72220
rect 13227 72251 13269 72260
rect 13227 72211 13228 72251
rect 13268 72211 13269 72251
rect 13611 72220 13612 72260
rect 13652 72220 13653 72260
rect 13611 72211 13653 72220
rect 14859 72251 14901 72260
rect 14859 72211 14860 72251
rect 14900 72211 14901 72251
rect 15243 72220 15244 72260
rect 15284 72220 15285 72260
rect 15243 72211 15285 72220
rect 16491 72251 16533 72260
rect 16491 72211 16492 72251
rect 16532 72211 16533 72251
rect 17307 72220 17308 72260
rect 17348 72220 17349 72260
rect 17307 72211 17349 72220
rect 17451 72260 17493 72269
rect 17451 72220 17452 72260
rect 17492 72220 17493 72260
rect 17451 72211 17493 72220
rect 17643 72260 17685 72269
rect 17643 72220 17644 72260
rect 17684 72220 17685 72260
rect 17643 72211 17685 72220
rect 17818 72260 17876 72261
rect 17818 72220 17827 72260
rect 17867 72220 17876 72260
rect 17818 72219 17876 72220
rect 17931 72260 17973 72269
rect 17931 72220 17932 72260
rect 17972 72220 17973 72260
rect 17931 72211 17973 72220
rect 18381 72260 18423 72269
rect 18381 72220 18382 72260
rect 18422 72220 18423 72260
rect 18381 72211 18423 72220
rect 18512 72260 18554 72269
rect 18512 72220 18513 72260
rect 18553 72220 18554 72260
rect 18512 72211 18554 72220
rect 18891 72260 18933 72269
rect 18891 72220 18892 72260
rect 18932 72220 18933 72260
rect 18891 72211 18933 72220
rect 19467 72251 19509 72260
rect 19467 72211 19468 72251
rect 19508 72211 19509 72251
rect 7851 72202 7893 72211
rect 13227 72202 13269 72211
rect 14859 72202 14901 72211
rect 16491 72202 16533 72211
rect 19467 72202 19509 72211
rect 19947 72251 19989 72260
rect 19947 72211 19948 72251
rect 19988 72211 19989 72251
rect 19947 72202 19989 72211
rect 1419 72176 1461 72185
rect 1419 72136 1420 72176
rect 1460 72136 1461 72176
rect 1419 72127 1461 72136
rect 1803 72176 1845 72185
rect 1803 72136 1804 72176
rect 1844 72136 1845 72176
rect 1803 72127 1845 72136
rect 2187 72176 2229 72185
rect 2187 72136 2188 72176
rect 2228 72136 2229 72176
rect 2187 72127 2229 72136
rect 2571 72176 2613 72185
rect 2571 72136 2572 72176
rect 2612 72136 2613 72176
rect 2571 72127 2613 72136
rect 3435 72176 3477 72185
rect 3435 72136 3436 72176
rect 3476 72136 3477 72176
rect 3435 72127 3477 72136
rect 4731 72176 4773 72185
rect 4731 72136 4732 72176
rect 4772 72136 4773 72176
rect 4731 72127 4773 72136
rect 4971 72176 5013 72185
rect 4971 72136 4972 72176
rect 5012 72136 5013 72176
rect 4971 72127 5013 72136
rect 5355 72176 5397 72185
rect 5355 72136 5356 72176
rect 5396 72136 5397 72176
rect 5355 72127 5397 72136
rect 5739 72176 5781 72185
rect 5739 72136 5740 72176
rect 5780 72136 5781 72176
rect 5739 72127 5781 72136
rect 6891 72176 6933 72185
rect 6891 72136 6892 72176
rect 6932 72136 6933 72176
rect 6891 72127 6933 72136
rect 8074 72176 8132 72177
rect 8074 72136 8083 72176
rect 8123 72136 8132 72176
rect 8074 72135 8132 72136
rect 8427 72176 8469 72185
rect 8427 72136 8428 72176
rect 8468 72136 8469 72176
rect 8427 72127 8469 72136
rect 8619 72176 8661 72185
rect 8619 72136 8620 72176
rect 8660 72136 8661 72176
rect 8619 72127 8661 72136
rect 8955 72176 8997 72185
rect 8955 72136 8956 72176
rect 8996 72136 8997 72176
rect 8955 72127 8997 72136
rect 9195 72176 9237 72185
rect 9195 72136 9196 72176
rect 9236 72136 9237 72176
rect 9195 72127 9237 72136
rect 9387 72176 9429 72185
rect 9387 72136 9388 72176
rect 9428 72136 9429 72176
rect 9387 72127 9429 72136
rect 9963 72176 10005 72185
rect 9963 72136 9964 72176
rect 10004 72136 10005 72176
rect 9963 72127 10005 72136
rect 10347 72176 10389 72185
rect 10347 72136 10348 72176
rect 10388 72136 10389 72176
rect 10347 72127 10389 72136
rect 10731 72176 10773 72185
rect 10731 72136 10732 72176
rect 10772 72136 10773 72176
rect 10731 72127 10773 72136
rect 11499 72176 11541 72185
rect 11499 72136 11500 72176
rect 11540 72136 11541 72176
rect 11499 72127 11541 72136
rect 18987 72176 19029 72185
rect 18987 72136 18988 72176
rect 19028 72136 19029 72176
rect 18987 72127 19029 72136
rect 1179 72092 1221 72101
rect 1179 72052 1180 72092
rect 1220 72052 1221 72092
rect 1179 72043 1221 72052
rect 1563 72092 1605 72101
rect 1563 72052 1564 72092
rect 1604 72052 1605 72092
rect 1563 72043 1605 72052
rect 1947 72092 1989 72101
rect 1947 72052 1948 72092
rect 1988 72052 1989 72092
rect 1947 72043 1989 72052
rect 8187 72092 8229 72101
rect 8187 72052 8188 72092
rect 8228 72052 8229 72092
rect 8187 72043 8229 72052
rect 8859 72092 8901 72101
rect 8859 72052 8860 72092
rect 8900 72052 8901 72092
rect 8859 72043 8901 72052
rect 9627 72092 9669 72101
rect 9627 72052 9628 72092
rect 9668 72052 9669 72092
rect 9627 72043 9669 72052
rect 17931 72092 17973 72101
rect 17931 72052 17932 72092
rect 17972 72052 17973 72092
rect 17931 72043 17973 72052
rect 9723 72008 9765 72017
rect 9723 71968 9724 72008
rect 9764 71968 9765 72008
rect 9723 71959 9765 71968
rect 13419 72008 13461 72017
rect 13419 71968 13420 72008
rect 13460 71968 13461 72008
rect 13419 71959 13461 71968
rect 16683 72008 16725 72017
rect 16683 71968 16684 72008
rect 16724 71968 16725 72008
rect 16683 71959 16725 71968
rect 1152 71840 20448 71864
rect 1152 71800 3688 71840
rect 3728 71800 3770 71840
rect 3810 71800 3852 71840
rect 3892 71800 3934 71840
rect 3974 71800 4016 71840
rect 4056 71800 18808 71840
rect 18848 71800 18890 71840
rect 18930 71800 18972 71840
rect 19012 71800 19054 71840
rect 19094 71800 19136 71840
rect 19176 71800 20448 71840
rect 1152 71776 20448 71800
rect 2139 71672 2181 71681
rect 2139 71632 2140 71672
rect 2180 71632 2181 71672
rect 2139 71623 2181 71632
rect 8139 71672 8181 71681
rect 8139 71632 8140 71672
rect 8180 71632 8181 71672
rect 8139 71623 8181 71632
rect 1419 71504 1461 71513
rect 1419 71464 1420 71504
rect 1460 71464 1461 71504
rect 1419 71455 1461 71464
rect 1899 71504 1941 71513
rect 1899 71464 1900 71504
rect 1940 71464 1941 71504
rect 1899 71455 1941 71464
rect 2283 71504 2325 71513
rect 2283 71464 2284 71504
rect 2324 71464 2325 71504
rect 2283 71455 2325 71464
rect 3339 71504 3381 71513
rect 3339 71464 3340 71504
rect 3380 71464 3381 71504
rect 3339 71455 3381 71464
rect 12459 71504 12501 71513
rect 12459 71464 12460 71504
rect 12500 71464 12501 71504
rect 12459 71455 12501 71464
rect 13738 71504 13796 71505
rect 13738 71464 13747 71504
rect 13787 71464 13796 71504
rect 13738 71463 13796 71464
rect 14091 71504 14133 71513
rect 14091 71464 14092 71504
rect 14132 71464 14133 71504
rect 14091 71455 14133 71464
rect 14763 71504 14805 71513
rect 14763 71464 14764 71504
rect 14804 71464 14805 71504
rect 14763 71455 14805 71464
rect 15531 71504 15573 71513
rect 15531 71464 15532 71504
rect 15572 71464 15573 71504
rect 15531 71455 15573 71464
rect 17259 71504 17301 71513
rect 17259 71464 17260 71504
rect 17300 71464 17301 71504
rect 17259 71455 17301 71464
rect 17643 71504 17685 71513
rect 17643 71464 17644 71504
rect 17684 71464 17685 71504
rect 17643 71455 17685 71464
rect 18603 71504 18645 71513
rect 18603 71464 18604 71504
rect 18644 71464 18645 71504
rect 18603 71455 18645 71464
rect 20139 71504 20181 71513
rect 20139 71464 20140 71504
rect 20180 71464 20181 71504
rect 20139 71455 20181 71464
rect 2829 71420 2871 71429
rect 2829 71380 2830 71420
rect 2870 71380 2871 71420
rect 2829 71371 2871 71380
rect 2955 71420 2997 71429
rect 2955 71380 2956 71420
rect 2996 71380 2997 71420
rect 2955 71371 2997 71380
rect 3435 71420 3477 71429
rect 3435 71380 3436 71420
rect 3476 71380 3477 71420
rect 3435 71371 3477 71380
rect 3907 71420 3965 71421
rect 3907 71380 3916 71420
rect 3956 71380 3965 71420
rect 3907 71379 3965 71380
rect 4395 71420 4453 71421
rect 4395 71380 4404 71420
rect 4444 71380 4453 71420
rect 4395 71379 4453 71380
rect 4779 71420 4821 71429
rect 4779 71380 4780 71420
rect 4820 71380 4821 71420
rect 4779 71371 4821 71380
rect 6019 71420 6077 71421
rect 6019 71380 6028 71420
rect 6068 71380 6077 71420
rect 6019 71379 6077 71380
rect 6699 71420 6741 71429
rect 6699 71380 6700 71420
rect 6740 71380 6741 71420
rect 6699 71371 6741 71380
rect 7939 71420 7997 71421
rect 7939 71380 7948 71420
rect 7988 71380 7997 71420
rect 7939 71379 7997 71380
rect 8619 71420 8661 71429
rect 8619 71380 8620 71420
rect 8660 71380 8661 71420
rect 8619 71371 8661 71380
rect 9859 71420 9917 71421
rect 9859 71380 9868 71420
rect 9908 71380 9917 71420
rect 9859 71379 9917 71380
rect 10251 71420 10293 71429
rect 10251 71380 10252 71420
rect 10292 71380 10293 71420
rect 10251 71371 10293 71380
rect 11491 71420 11549 71421
rect 11491 71380 11500 71420
rect 11540 71380 11549 71420
rect 11491 71379 11549 71380
rect 11962 71420 12020 71421
rect 11962 71380 11971 71420
rect 12011 71380 12020 71420
rect 11962 71379 12020 71380
rect 12075 71420 12117 71429
rect 12075 71380 12076 71420
rect 12116 71380 12117 71420
rect 12075 71371 12117 71380
rect 12555 71420 12597 71429
rect 12555 71380 12556 71420
rect 12596 71380 12597 71420
rect 12555 71371 12597 71380
rect 13027 71420 13085 71421
rect 13027 71380 13036 71420
rect 13076 71380 13085 71420
rect 13027 71379 13085 71380
rect 13515 71420 13573 71421
rect 13515 71380 13524 71420
rect 13564 71380 13573 71420
rect 13515 71379 13573 71380
rect 15034 71420 15092 71421
rect 15034 71380 15043 71420
rect 15083 71380 15092 71420
rect 15034 71379 15092 71380
rect 15147 71420 15189 71429
rect 15147 71380 15148 71420
rect 15188 71380 15189 71420
rect 15147 71371 15189 71380
rect 15627 71420 15669 71429
rect 15627 71380 15628 71420
rect 15668 71380 15669 71420
rect 15627 71371 15669 71380
rect 16099 71420 16157 71421
rect 16099 71380 16108 71420
rect 16148 71380 16157 71420
rect 16099 71379 16157 71380
rect 16618 71420 16676 71421
rect 16618 71380 16627 71420
rect 16667 71380 16676 71420
rect 16618 71379 16676 71380
rect 18106 71420 18164 71421
rect 18106 71380 18115 71420
rect 18155 71380 18164 71420
rect 18106 71379 18164 71380
rect 18219 71420 18261 71429
rect 18219 71380 18220 71420
rect 18260 71380 18261 71420
rect 18219 71371 18261 71380
rect 18699 71420 18741 71429
rect 18699 71380 18700 71420
rect 18740 71380 18741 71420
rect 18699 71371 18741 71380
rect 19171 71420 19229 71421
rect 19171 71380 19180 71420
rect 19220 71380 19229 71420
rect 19171 71379 19229 71380
rect 19690 71420 19748 71421
rect 19690 71380 19699 71420
rect 19739 71380 19748 71420
rect 19690 71379 19748 71380
rect 2523 71336 2565 71345
rect 2523 71296 2524 71336
rect 2564 71296 2565 71336
rect 2523 71287 2565 71296
rect 11691 71336 11733 71345
rect 11691 71296 11692 71336
rect 11732 71296 11733 71336
rect 11691 71287 11733 71296
rect 1179 71252 1221 71261
rect 1179 71212 1180 71252
rect 1220 71212 1221 71252
rect 1179 71203 1221 71212
rect 4587 71252 4629 71261
rect 4587 71212 4588 71252
rect 4628 71212 4629 71252
rect 4587 71203 4629 71212
rect 6219 71252 6261 71261
rect 6219 71212 6220 71252
rect 6260 71212 6261 71252
rect 6219 71203 6261 71212
rect 10059 71252 10101 71261
rect 10059 71212 10060 71252
rect 10100 71212 10101 71252
rect 10059 71203 10101 71212
rect 13851 71252 13893 71261
rect 13851 71212 13852 71252
rect 13892 71212 13893 71252
rect 13851 71203 13893 71212
rect 14523 71252 14565 71261
rect 14523 71212 14524 71252
rect 14564 71212 14565 71252
rect 14523 71203 14565 71212
rect 16779 71252 16821 71261
rect 16779 71212 16780 71252
rect 16820 71212 16821 71252
rect 16779 71203 16821 71212
rect 17499 71252 17541 71261
rect 17499 71212 17500 71252
rect 17540 71212 17541 71252
rect 17499 71203 17541 71212
rect 17883 71252 17925 71261
rect 17883 71212 17884 71252
rect 17924 71212 17925 71252
rect 17883 71203 17925 71212
rect 19851 71252 19893 71261
rect 19851 71212 19852 71252
rect 19892 71212 19893 71252
rect 19851 71203 19893 71212
rect 20379 71252 20421 71261
rect 20379 71212 20380 71252
rect 20420 71212 20421 71252
rect 20379 71203 20421 71212
rect 1152 71084 20452 71108
rect 1152 71044 4928 71084
rect 4968 71044 5010 71084
rect 5050 71044 5092 71084
rect 5132 71044 5174 71084
rect 5214 71044 5256 71084
rect 5296 71044 20048 71084
rect 20088 71044 20130 71084
rect 20170 71044 20212 71084
rect 20252 71044 20294 71084
rect 20334 71044 20376 71084
rect 20416 71044 20452 71084
rect 1152 71020 20452 71044
rect 1563 70916 1605 70925
rect 1563 70876 1564 70916
rect 1604 70876 1605 70916
rect 1563 70867 1605 70876
rect 7467 70916 7509 70925
rect 7467 70876 7468 70916
rect 7508 70876 7509 70916
rect 7467 70867 7509 70876
rect 13419 70916 13461 70925
rect 13419 70876 13420 70916
rect 13460 70876 13461 70916
rect 13419 70867 13461 70876
rect 15243 70916 15285 70925
rect 15243 70876 15244 70916
rect 15284 70876 15285 70916
rect 15243 70867 15285 70876
rect 18363 70916 18405 70925
rect 18363 70876 18364 70916
rect 18404 70876 18405 70916
rect 18363 70867 18405 70876
rect 10923 70832 10965 70841
rect 10923 70792 10924 70832
rect 10964 70792 10965 70832
rect 10923 70783 10965 70792
rect 1995 70748 2037 70757
rect 4378 70748 4436 70749
rect 1995 70708 1996 70748
rect 2036 70708 2037 70748
rect 1995 70699 2037 70708
rect 3243 70739 3285 70748
rect 3243 70699 3244 70739
rect 3284 70699 3285 70739
rect 4378 70708 4387 70748
rect 4427 70708 4436 70748
rect 4378 70707 4436 70708
rect 4491 70748 4533 70757
rect 4491 70708 4492 70748
rect 4532 70708 4533 70748
rect 4491 70699 4533 70708
rect 4875 70748 4917 70757
rect 7179 70748 7221 70757
rect 4875 70708 4876 70748
rect 4916 70708 4917 70748
rect 4875 70699 4917 70708
rect 5451 70739 5493 70748
rect 5451 70699 5452 70739
rect 5492 70699 5493 70739
rect 3243 70690 3285 70699
rect 5451 70690 5493 70699
rect 5931 70739 5973 70748
rect 5931 70699 5932 70739
rect 5972 70699 5973 70739
rect 7179 70708 7180 70748
rect 7220 70708 7221 70748
rect 7179 70699 7221 70708
rect 7313 70748 7371 70749
rect 9099 70748 9141 70757
rect 7313 70708 7322 70748
rect 7362 70708 7371 70748
rect 7313 70707 7371 70708
rect 7851 70739 7893 70748
rect 7851 70699 7852 70739
rect 7892 70699 7893 70739
rect 9099 70708 9100 70748
rect 9140 70708 9141 70748
rect 9099 70699 9141 70708
rect 9483 70748 9525 70757
rect 11674 70748 11732 70749
rect 9483 70708 9484 70748
rect 9524 70708 9525 70748
rect 9483 70699 9525 70708
rect 10731 70739 10773 70748
rect 10731 70699 10732 70739
rect 10772 70699 10773 70739
rect 11674 70708 11683 70748
rect 11723 70708 11732 70748
rect 11674 70707 11732 70708
rect 11787 70748 11829 70757
rect 11787 70708 11788 70748
rect 11828 70708 11829 70748
rect 11787 70699 11829 70708
rect 12171 70748 12213 70757
rect 13803 70748 13845 70757
rect 16107 70748 16149 70757
rect 18795 70748 18837 70757
rect 12171 70708 12172 70748
rect 12212 70708 12213 70748
rect 12171 70699 12213 70708
rect 12747 70739 12789 70748
rect 12747 70699 12748 70739
rect 12788 70699 12789 70739
rect 5931 70690 5973 70699
rect 7851 70690 7893 70699
rect 10731 70690 10773 70699
rect 12747 70690 12789 70699
rect 13227 70739 13269 70748
rect 13227 70699 13228 70739
rect 13268 70699 13269 70739
rect 13803 70708 13804 70748
rect 13844 70708 13845 70748
rect 13803 70699 13845 70708
rect 15051 70739 15093 70748
rect 15051 70699 15052 70739
rect 15092 70699 15093 70739
rect 16107 70708 16108 70748
rect 16148 70708 16149 70748
rect 16107 70699 16149 70708
rect 17355 70739 17397 70748
rect 17355 70699 17356 70739
rect 17396 70699 17397 70739
rect 18795 70708 18796 70748
rect 18836 70708 18837 70748
rect 18795 70699 18837 70708
rect 20043 70739 20085 70748
rect 20043 70699 20044 70739
rect 20084 70699 20085 70739
rect 13227 70690 13269 70699
rect 15051 70690 15093 70699
rect 17355 70690 17397 70699
rect 20043 70690 20085 70699
rect 1419 70664 1461 70673
rect 1419 70624 1420 70664
rect 1460 70624 1461 70664
rect 1419 70615 1461 70624
rect 1803 70664 1845 70673
rect 1803 70624 1804 70664
rect 1844 70624 1845 70664
rect 1803 70615 1845 70624
rect 3819 70664 3861 70673
rect 3819 70624 3820 70664
rect 3860 70624 3861 70664
rect 3819 70615 3861 70624
rect 4971 70664 5013 70673
rect 4971 70624 4972 70664
rect 5012 70624 5013 70664
rect 4971 70615 5013 70624
rect 6315 70664 6357 70673
rect 6315 70624 6316 70664
rect 6356 70624 6357 70664
rect 6315 70615 6357 70624
rect 6891 70664 6933 70673
rect 6891 70624 6892 70664
rect 6932 70624 6933 70664
rect 6891 70615 6933 70624
rect 11067 70664 11109 70673
rect 11067 70624 11068 70664
rect 11108 70624 11109 70664
rect 11067 70615 11109 70624
rect 11307 70664 11349 70673
rect 11307 70624 11308 70664
rect 11348 70624 11349 70664
rect 11307 70615 11349 70624
rect 12267 70664 12309 70673
rect 12267 70624 12268 70664
rect 12308 70624 12309 70664
rect 12267 70615 12309 70624
rect 15915 70664 15957 70673
rect 15915 70624 15916 70664
rect 15956 70624 15957 70664
rect 15915 70615 15957 70624
rect 18027 70664 18069 70673
rect 18027 70624 18028 70664
rect 18068 70624 18069 70664
rect 18027 70615 18069 70624
rect 18603 70664 18645 70673
rect 18603 70624 18604 70664
rect 18644 70624 18645 70664
rect 18603 70615 18645 70624
rect 1179 70580 1221 70589
rect 1179 70540 1180 70580
rect 1220 70540 1221 70580
rect 1179 70531 1221 70540
rect 3579 70580 3621 70589
rect 3579 70540 3580 70580
rect 3620 70540 3621 70580
rect 3579 70531 3621 70540
rect 6171 70580 6213 70589
rect 6171 70540 6172 70580
rect 6212 70540 6213 70580
rect 6171 70531 6213 70540
rect 6651 70580 6693 70589
rect 6651 70540 6652 70580
rect 6692 70540 6693 70580
rect 6651 70531 6693 70540
rect 15675 70580 15717 70589
rect 15675 70540 15676 70580
rect 15716 70540 15717 70580
rect 15675 70531 15717 70540
rect 18267 70580 18309 70589
rect 18267 70540 18268 70580
rect 18308 70540 18309 70580
rect 18267 70531 18309 70540
rect 20235 70580 20277 70589
rect 20235 70540 20236 70580
rect 20276 70540 20277 70580
rect 20235 70531 20277 70540
rect 3435 70496 3477 70505
rect 3435 70456 3436 70496
rect 3476 70456 3477 70496
rect 3435 70447 3477 70456
rect 6555 70496 6597 70505
rect 6555 70456 6556 70496
rect 6596 70456 6597 70496
rect 6555 70447 6597 70456
rect 7659 70496 7701 70505
rect 7659 70456 7660 70496
rect 7700 70456 7701 70496
rect 7659 70447 7701 70456
rect 17547 70496 17589 70505
rect 17547 70456 17548 70496
rect 17588 70456 17589 70496
rect 17547 70447 17589 70456
rect 1152 70328 20448 70352
rect 1152 70288 3688 70328
rect 3728 70288 3770 70328
rect 3810 70288 3852 70328
rect 3892 70288 3934 70328
rect 3974 70288 4016 70328
rect 4056 70288 18808 70328
rect 18848 70288 18890 70328
rect 18930 70288 18972 70328
rect 19012 70288 19054 70328
rect 19094 70288 19136 70328
rect 19176 70288 20448 70328
rect 1152 70264 20448 70288
rect 12603 70160 12645 70169
rect 12603 70120 12604 70160
rect 12644 70120 12645 70160
rect 12603 70111 12645 70120
rect 16059 70160 16101 70169
rect 16059 70120 16060 70160
rect 16100 70120 16101 70160
rect 16059 70111 16101 70120
rect 17403 70160 17445 70169
rect 17403 70120 17404 70160
rect 17444 70120 17445 70160
rect 17403 70111 17445 70120
rect 16731 70076 16773 70085
rect 16731 70036 16732 70076
rect 16772 70036 16773 70076
rect 16731 70027 16773 70036
rect 3531 69992 3573 70001
rect 3531 69952 3532 69992
rect 3572 69952 3573 69992
rect 3531 69943 3573 69952
rect 8139 69992 8181 70001
rect 8139 69952 8140 69992
rect 8180 69952 8181 69992
rect 8139 69943 8181 69952
rect 9195 69992 9237 70001
rect 9195 69952 9196 69992
rect 9236 69952 9237 69992
rect 9195 69943 9237 69952
rect 9562 69992 9620 69993
rect 9562 69952 9571 69992
rect 9611 69952 9620 69992
rect 9562 69951 9620 69952
rect 11211 69992 11253 70001
rect 11211 69952 11212 69992
rect 11252 69952 11253 69992
rect 11211 69943 11253 69952
rect 12363 69992 12405 70001
rect 12363 69952 12364 69992
rect 12404 69952 12405 69992
rect 12363 69943 12405 69952
rect 16299 69992 16341 70001
rect 16299 69952 16300 69992
rect 16340 69952 16341 69992
rect 16299 69943 16341 69952
rect 16971 69992 17013 70001
rect 16971 69952 16972 69992
rect 17012 69952 17013 69992
rect 16971 69943 17013 69952
rect 17163 69992 17205 70001
rect 17163 69952 17164 69992
rect 17204 69952 17205 69992
rect 17163 69943 17205 69952
rect 18123 69992 18165 70001
rect 18123 69952 18124 69992
rect 18164 69952 18165 69992
rect 18123 69943 18165 69952
rect 19755 69992 19797 70001
rect 19755 69952 19756 69992
rect 19796 69952 19797 69992
rect 19755 69943 19797 69952
rect 20139 69992 20181 70001
rect 20139 69952 20140 69992
rect 20180 69952 20181 69992
rect 20139 69943 20181 69952
rect 1515 69908 1557 69917
rect 1515 69868 1516 69908
rect 1556 69868 1557 69908
rect 1515 69859 1557 69868
rect 2755 69908 2813 69909
rect 2755 69868 2764 69908
rect 2804 69868 2813 69908
rect 2755 69867 2813 69868
rect 3907 69908 3965 69909
rect 3907 69868 3916 69908
rect 3956 69868 3965 69908
rect 3907 69867 3965 69868
rect 5163 69908 5205 69917
rect 5163 69868 5164 69908
rect 5204 69868 5205 69908
rect 5163 69859 5205 69868
rect 5355 69908 5397 69917
rect 5355 69868 5356 69908
rect 5396 69868 5397 69908
rect 5355 69859 5397 69868
rect 6595 69908 6653 69909
rect 6595 69868 6604 69908
rect 6644 69868 6653 69908
rect 6595 69867 6653 69868
rect 7162 69908 7220 69909
rect 7162 69868 7171 69908
rect 7211 69868 7220 69908
rect 7162 69867 7220 69868
rect 7651 69908 7709 69909
rect 7651 69868 7660 69908
rect 7700 69868 7709 69908
rect 7651 69867 7709 69868
rect 8235 69908 8277 69917
rect 8235 69868 8236 69908
rect 8276 69868 8277 69908
rect 8235 69859 8277 69868
rect 8619 69908 8661 69917
rect 8619 69868 8620 69908
rect 8660 69868 8661 69908
rect 8619 69859 8661 69868
rect 8729 69908 8787 69909
rect 8729 69868 8738 69908
rect 8778 69868 8787 69908
rect 8729 69867 8787 69868
rect 9763 69908 9821 69909
rect 9763 69868 9772 69908
rect 9812 69868 9821 69908
rect 9763 69867 9821 69868
rect 11019 69908 11061 69917
rect 11019 69868 11020 69908
rect 11060 69868 11061 69908
rect 11019 69859 11061 69868
rect 12747 69908 12789 69917
rect 12747 69868 12748 69908
rect 12788 69868 12789 69908
rect 12747 69859 12789 69868
rect 13987 69908 14045 69909
rect 13987 69868 13996 69908
rect 14036 69868 14045 69908
rect 13987 69867 14045 69868
rect 14475 69908 14517 69917
rect 14475 69868 14476 69908
rect 14516 69868 14517 69908
rect 14475 69859 14517 69868
rect 15715 69908 15773 69909
rect 15715 69868 15724 69908
rect 15764 69868 15773 69908
rect 15715 69867 15773 69868
rect 17613 69908 17655 69917
rect 17613 69868 17614 69908
rect 17654 69868 17655 69908
rect 17613 69859 17655 69868
rect 17739 69908 17781 69917
rect 17739 69868 17740 69908
rect 17780 69868 17781 69908
rect 17739 69859 17781 69868
rect 18219 69908 18261 69917
rect 18219 69868 18220 69908
rect 18260 69868 18261 69908
rect 18219 69859 18261 69868
rect 18691 69908 18749 69909
rect 18691 69868 18700 69908
rect 18740 69868 18749 69908
rect 18691 69867 18749 69868
rect 19210 69908 19268 69909
rect 19210 69868 19219 69908
rect 19259 69868 19268 69908
rect 19210 69867 19268 69868
rect 19995 69824 20037 69833
rect 19995 69784 19996 69824
rect 20036 69784 20037 69824
rect 19995 69775 20037 69784
rect 2955 69740 2997 69749
rect 2955 69700 2956 69740
rect 2996 69700 2997 69740
rect 2955 69691 2997 69700
rect 3291 69740 3333 69749
rect 3291 69700 3292 69740
rect 3332 69700 3333 69740
rect 3291 69691 3333 69700
rect 3723 69740 3765 69749
rect 3723 69700 3724 69740
rect 3764 69700 3765 69740
rect 3723 69691 3765 69700
rect 6795 69740 6837 69749
rect 6795 69700 6796 69740
rect 6836 69700 6837 69740
rect 6795 69691 6837 69700
rect 6987 69740 7029 69749
rect 6987 69700 6988 69740
rect 7028 69700 7029 69740
rect 6987 69691 7029 69700
rect 8955 69740 8997 69749
rect 8955 69700 8956 69740
rect 8996 69700 8997 69740
rect 8955 69691 8997 69700
rect 11451 69740 11493 69749
rect 11451 69700 11452 69740
rect 11492 69700 11493 69740
rect 11451 69691 11493 69700
rect 14187 69740 14229 69749
rect 14187 69700 14188 69740
rect 14228 69700 14229 69740
rect 14187 69691 14229 69700
rect 15915 69740 15957 69749
rect 15915 69700 15916 69740
rect 15956 69700 15957 69740
rect 15915 69691 15957 69700
rect 19371 69740 19413 69749
rect 19371 69700 19372 69740
rect 19412 69700 19413 69740
rect 19371 69691 19413 69700
rect 20379 69740 20421 69749
rect 20379 69700 20380 69740
rect 20420 69700 20421 69740
rect 20379 69691 20421 69700
rect 1152 69572 20452 69596
rect 1152 69532 4928 69572
rect 4968 69532 5010 69572
rect 5050 69532 5092 69572
rect 5132 69532 5174 69572
rect 5214 69532 5256 69572
rect 5296 69532 20048 69572
rect 20088 69532 20130 69572
rect 20170 69532 20212 69572
rect 20252 69532 20294 69572
rect 20334 69532 20376 69572
rect 20416 69532 20452 69572
rect 1152 69508 20452 69532
rect 4875 69404 4917 69413
rect 4875 69364 4876 69404
rect 4916 69364 4917 69404
rect 4875 69355 4917 69364
rect 7546 69404 7604 69405
rect 7546 69364 7555 69404
rect 7595 69364 7604 69404
rect 7546 69363 7604 69364
rect 16011 69404 16053 69413
rect 16011 69364 16012 69404
rect 16052 69364 16053 69404
rect 16011 69355 16053 69364
rect 20043 69404 20085 69413
rect 20043 69364 20044 69404
rect 20084 69364 20085 69404
rect 20043 69355 20085 69364
rect 5019 69320 5061 69329
rect 10683 69320 10725 69329
rect 5019 69280 5020 69320
rect 5060 69280 5061 69320
rect 5019 69271 5061 69280
rect 7842 69311 7888 69320
rect 7842 69271 7843 69311
rect 7883 69271 7888 69311
rect 10683 69280 10684 69320
rect 10724 69280 10725 69320
rect 10683 69271 10725 69280
rect 18027 69320 18069 69329
rect 18027 69280 18028 69320
rect 18068 69280 18069 69320
rect 18027 69271 18069 69280
rect 7842 69262 7888 69271
rect 1419 69236 1461 69245
rect 3117 69236 3159 69245
rect 1419 69196 1420 69236
rect 1460 69196 1461 69236
rect 1419 69187 1461 69196
rect 2667 69227 2709 69236
rect 2667 69187 2668 69227
rect 2708 69187 2709 69227
rect 3117 69196 3118 69236
rect 3158 69196 3159 69236
rect 3117 69187 3159 69196
rect 3243 69236 3285 69245
rect 3243 69196 3244 69236
rect 3284 69196 3285 69236
rect 3243 69187 3285 69196
rect 3627 69236 3669 69245
rect 5451 69236 5493 69245
rect 3627 69196 3628 69236
rect 3668 69196 3669 69236
rect 3627 69187 3669 69196
rect 4203 69227 4245 69236
rect 4203 69187 4204 69227
rect 4244 69187 4245 69227
rect 2667 69178 2709 69187
rect 4203 69178 4245 69187
rect 4683 69227 4725 69236
rect 4683 69187 4684 69227
rect 4724 69187 4725 69227
rect 5451 69196 5452 69236
rect 5492 69196 5493 69236
rect 5451 69187 5493 69196
rect 5626 69236 5684 69237
rect 5626 69196 5635 69236
rect 5675 69196 5684 69236
rect 5626 69195 5684 69196
rect 5739 69236 5781 69245
rect 5739 69196 5740 69236
rect 5780 69196 5781 69236
rect 5739 69187 5781 69196
rect 5931 69236 5973 69245
rect 7546 69236 7604 69237
rect 7930 69236 7988 69237
rect 5931 69196 5932 69236
rect 5972 69196 5973 69236
rect 5931 69187 5973 69196
rect 7179 69227 7221 69236
rect 7179 69187 7180 69227
rect 7220 69187 7221 69227
rect 7546 69196 7555 69236
rect 7595 69196 7604 69236
rect 7546 69195 7604 69196
rect 7659 69227 7701 69236
rect 4683 69178 4725 69187
rect 7179 69178 7221 69187
rect 7659 69187 7660 69227
rect 7700 69187 7701 69227
rect 7930 69196 7939 69236
rect 7979 69196 7988 69236
rect 7930 69195 7988 69196
rect 8064 69236 8122 69237
rect 8064 69196 8073 69236
rect 8113 69196 8122 69236
rect 8064 69195 8122 69196
rect 8427 69236 8469 69245
rect 11499 69236 11541 69245
rect 14266 69236 14324 69237
rect 8427 69196 8428 69236
rect 8468 69196 8469 69236
rect 8427 69187 8469 69196
rect 9675 69227 9717 69236
rect 9675 69187 9676 69227
rect 9716 69187 9717 69227
rect 11499 69196 11500 69236
rect 11540 69196 11541 69236
rect 11499 69187 11541 69196
rect 12747 69227 12789 69236
rect 12747 69187 12748 69227
rect 12788 69187 12789 69227
rect 14266 69196 14275 69236
rect 14315 69196 14324 69236
rect 14266 69195 14324 69196
rect 14379 69236 14421 69245
rect 14379 69196 14380 69236
rect 14420 69196 14421 69236
rect 14379 69187 14421 69196
rect 14859 69236 14901 69245
rect 16587 69236 16629 69245
rect 18298 69236 18356 69237
rect 14859 69196 14860 69236
rect 14900 69196 14901 69236
rect 14859 69187 14901 69196
rect 15339 69227 15381 69236
rect 15339 69187 15340 69227
rect 15380 69187 15381 69227
rect 7659 69178 7701 69187
rect 9675 69178 9717 69187
rect 12747 69178 12789 69187
rect 15339 69178 15381 69187
rect 15819 69227 15861 69236
rect 15819 69187 15820 69227
rect 15860 69187 15861 69227
rect 16587 69196 16588 69236
rect 16628 69196 16629 69236
rect 16587 69187 16629 69196
rect 17835 69227 17877 69236
rect 17835 69187 17836 69227
rect 17876 69187 17877 69227
rect 18298 69196 18307 69236
rect 18347 69196 18356 69236
rect 18298 69195 18356 69196
rect 18411 69236 18453 69245
rect 18411 69196 18412 69236
rect 18452 69196 18453 69236
rect 18411 69187 18453 69196
rect 18795 69236 18837 69245
rect 18795 69196 18796 69236
rect 18836 69196 18837 69236
rect 18795 69187 18837 69196
rect 19371 69227 19413 69236
rect 19371 69187 19372 69227
rect 19412 69187 19413 69227
rect 15819 69178 15861 69187
rect 17835 69178 17877 69187
rect 19371 69178 19413 69187
rect 19851 69227 19893 69236
rect 19851 69187 19852 69227
rect 19892 69187 19893 69227
rect 19851 69178 19893 69187
rect 3723 69152 3765 69161
rect 3723 69112 3724 69152
rect 3764 69112 3765 69152
rect 3723 69103 3765 69112
rect 5259 69152 5301 69161
rect 5259 69112 5260 69152
rect 5300 69112 5301 69152
rect 5259 69103 5301 69112
rect 10251 69152 10293 69161
rect 10251 69112 10252 69152
rect 10292 69112 10293 69152
rect 10251 69103 10293 69112
rect 10443 69152 10485 69161
rect 10443 69112 10444 69152
rect 10484 69112 10485 69152
rect 10443 69103 10485 69112
rect 13323 69152 13365 69161
rect 13323 69112 13324 69152
rect 13364 69112 13365 69152
rect 13323 69103 13365 69112
rect 13803 69152 13845 69161
rect 13803 69112 13804 69152
rect 13844 69112 13845 69152
rect 13803 69103 13845 69112
rect 14043 69152 14085 69161
rect 14043 69112 14044 69152
rect 14084 69112 14085 69152
rect 14043 69103 14085 69112
rect 14763 69152 14805 69161
rect 14763 69112 14764 69152
rect 14804 69112 14805 69152
rect 14763 69103 14805 69112
rect 16155 69152 16197 69161
rect 16155 69112 16156 69152
rect 16196 69112 16197 69152
rect 16155 69103 16197 69112
rect 16395 69152 16437 69161
rect 16395 69112 16396 69152
rect 16436 69112 16437 69152
rect 16395 69103 16437 69112
rect 18891 69152 18933 69161
rect 18891 69112 18892 69152
rect 18932 69112 18933 69152
rect 18891 69103 18933 69112
rect 7371 69068 7413 69077
rect 7371 69028 7372 69068
rect 7412 69028 7413 69068
rect 7371 69019 7413 69028
rect 13563 69068 13605 69077
rect 13563 69028 13564 69068
rect 13604 69028 13605 69068
rect 13563 69019 13605 69028
rect 2859 68984 2901 68993
rect 2859 68944 2860 68984
rect 2900 68944 2901 68984
rect 2859 68935 2901 68944
rect 5739 68984 5781 68993
rect 5739 68944 5740 68984
rect 5780 68944 5781 68984
rect 5739 68935 5781 68944
rect 9867 68984 9909 68993
rect 9867 68944 9868 68984
rect 9908 68944 9909 68984
rect 9867 68935 9909 68944
rect 10011 68984 10053 68993
rect 10011 68944 10012 68984
rect 10052 68944 10053 68984
rect 10011 68935 10053 68944
rect 12939 68984 12981 68993
rect 12939 68944 12940 68984
rect 12980 68944 12981 68984
rect 12939 68935 12981 68944
rect 1152 68816 20448 68840
rect 1152 68776 3688 68816
rect 3728 68776 3770 68816
rect 3810 68776 3852 68816
rect 3892 68776 3934 68816
rect 3974 68776 4016 68816
rect 4056 68776 18808 68816
rect 18848 68776 18890 68816
rect 18930 68776 18972 68816
rect 19012 68776 19054 68816
rect 19094 68776 19136 68816
rect 19176 68776 20448 68816
rect 1152 68752 20448 68776
rect 3195 68648 3237 68657
rect 3195 68608 3196 68648
rect 3236 68608 3237 68648
rect 3195 68599 3237 68608
rect 10011 68648 10053 68657
rect 10011 68608 10012 68648
rect 10052 68608 10053 68648
rect 10011 68599 10053 68608
rect 16827 68648 16869 68657
rect 16827 68608 16828 68648
rect 16868 68608 16869 68648
rect 16827 68599 16869 68608
rect 18987 68648 19029 68657
rect 18987 68608 18988 68648
rect 19028 68608 19029 68648
rect 18987 68599 19029 68608
rect 2811 68564 2853 68573
rect 2811 68524 2812 68564
rect 2852 68524 2853 68564
rect 2811 68515 2853 68524
rect 19419 68564 19461 68573
rect 19419 68524 19420 68564
rect 19460 68524 19461 68564
rect 19419 68515 19461 68524
rect 3051 68480 3093 68489
rect 3051 68440 3052 68480
rect 3092 68440 3093 68480
rect 3051 68431 3093 68440
rect 3435 68480 3477 68489
rect 3435 68440 3436 68480
rect 3476 68440 3477 68480
rect 3435 68431 3477 68440
rect 4299 68480 4341 68489
rect 4299 68440 4300 68480
rect 4340 68440 4341 68480
rect 4299 68431 4341 68440
rect 7371 68480 7413 68489
rect 7371 68440 7372 68480
rect 7412 68440 7413 68480
rect 7371 68431 7413 68440
rect 8331 68480 8373 68489
rect 8331 68440 8332 68480
rect 8372 68440 8373 68480
rect 8331 68431 8373 68440
rect 8458 68480 8516 68481
rect 8458 68440 8467 68480
rect 8507 68440 8516 68480
rect 8458 68439 8516 68440
rect 9771 68480 9813 68489
rect 9771 68440 9772 68480
rect 9812 68440 9813 68480
rect 9771 68431 9813 68440
rect 12747 68480 12789 68489
rect 12747 68440 12748 68480
rect 12788 68440 12789 68480
rect 12747 68431 12789 68440
rect 14026 68480 14084 68481
rect 14026 68440 14035 68480
rect 14075 68440 14084 68480
rect 14026 68439 14084 68440
rect 14379 68480 14421 68489
rect 14379 68440 14380 68480
rect 14420 68440 14421 68480
rect 14379 68431 14421 68440
rect 15339 68480 15381 68489
rect 15339 68440 15340 68480
rect 15380 68440 15381 68480
rect 15339 68431 15381 68440
rect 17067 68480 17109 68489
rect 17067 68440 17068 68480
rect 17108 68440 17109 68480
rect 17067 68431 17109 68440
rect 19659 68480 19701 68489
rect 19659 68440 19660 68480
rect 19700 68440 19701 68480
rect 19659 68431 19701 68440
rect 20139 68480 20181 68489
rect 20139 68440 20140 68480
rect 20180 68440 20181 68480
rect 20139 68431 20181 68440
rect 1227 68396 1269 68405
rect 1227 68356 1228 68396
rect 1268 68356 1269 68396
rect 1227 68347 1269 68356
rect 2467 68396 2525 68397
rect 2467 68356 2476 68396
rect 2516 68356 2525 68396
rect 2467 68355 2525 68356
rect 3802 68396 3860 68397
rect 3802 68356 3811 68396
rect 3851 68356 3860 68396
rect 3802 68355 3860 68356
rect 3915 68396 3957 68405
rect 3915 68356 3916 68396
rect 3956 68356 3957 68396
rect 3915 68347 3957 68356
rect 4395 68396 4437 68405
rect 4395 68356 4396 68396
rect 4436 68356 4437 68396
rect 4395 68347 4437 68356
rect 4867 68396 4925 68397
rect 4867 68356 4876 68396
rect 4916 68356 4925 68396
rect 4867 68355 4925 68356
rect 5386 68396 5444 68397
rect 5386 68356 5395 68396
rect 5435 68356 5444 68396
rect 5386 68355 5444 68356
rect 5923 68396 5981 68397
rect 5923 68356 5932 68396
rect 5972 68356 5981 68396
rect 5923 68355 5981 68356
rect 7179 68396 7221 68405
rect 7179 68356 7180 68396
rect 7220 68356 7221 68396
rect 7179 68347 7221 68356
rect 7834 68396 7892 68397
rect 7834 68356 7843 68396
rect 7883 68356 7892 68396
rect 7834 68355 7892 68356
rect 7947 68396 7989 68405
rect 7947 68356 7948 68396
rect 7988 68356 7989 68396
rect 7947 68347 7989 68356
rect 8899 68396 8957 68397
rect 8899 68356 8908 68396
rect 8948 68356 8957 68396
rect 8899 68355 8957 68356
rect 9418 68396 9476 68397
rect 9418 68356 9427 68396
rect 9467 68356 9476 68396
rect 9418 68355 9476 68356
rect 10443 68396 10485 68405
rect 10443 68356 10444 68396
rect 10484 68356 10485 68396
rect 10443 68347 10485 68356
rect 11683 68396 11741 68397
rect 11683 68356 11692 68396
rect 11732 68356 11741 68396
rect 11683 68355 11741 68356
rect 12250 68396 12308 68397
rect 12250 68356 12259 68396
rect 12299 68356 12308 68396
rect 12250 68355 12308 68356
rect 12363 68396 12405 68405
rect 12363 68356 12364 68396
rect 12404 68356 12405 68396
rect 12363 68347 12405 68356
rect 12843 68396 12885 68405
rect 12843 68356 12844 68396
rect 12884 68356 12885 68396
rect 12843 68347 12885 68356
rect 13315 68396 13373 68397
rect 13315 68356 13324 68396
rect 13364 68356 13373 68396
rect 13315 68355 13373 68356
rect 13803 68396 13861 68397
rect 13803 68356 13812 68396
rect 13852 68356 13861 68396
rect 13803 68355 13861 68356
rect 14842 68396 14900 68397
rect 14842 68356 14851 68396
rect 14891 68356 14900 68396
rect 14842 68355 14900 68356
rect 14955 68396 14997 68405
rect 14955 68356 14956 68396
rect 14996 68356 14997 68396
rect 14955 68347 14997 68356
rect 15435 68396 15477 68405
rect 15435 68356 15436 68396
rect 15476 68356 15477 68396
rect 15435 68347 15477 68356
rect 15907 68396 15965 68397
rect 15907 68356 15916 68396
rect 15956 68356 15965 68396
rect 15907 68355 15965 68356
rect 16395 68396 16453 68397
rect 16395 68356 16404 68396
rect 16444 68356 16453 68396
rect 16395 68355 16453 68356
rect 17547 68396 17589 68405
rect 17547 68356 17548 68396
rect 17588 68356 17589 68396
rect 17547 68347 17589 68356
rect 18787 68396 18845 68397
rect 18787 68356 18796 68396
rect 18836 68356 18845 68396
rect 18787 68355 18845 68356
rect 5739 68312 5781 68321
rect 5739 68272 5740 68312
rect 5780 68272 5781 68312
rect 5739 68263 5781 68272
rect 11883 68312 11925 68321
rect 11883 68272 11884 68312
rect 11924 68272 11925 68312
rect 11883 68263 11925 68272
rect 2667 68228 2709 68237
rect 2667 68188 2668 68228
rect 2708 68188 2709 68228
rect 2667 68179 2709 68188
rect 5547 68228 5589 68237
rect 5547 68188 5548 68228
rect 5588 68188 5589 68228
rect 5547 68179 5589 68188
rect 7611 68228 7653 68237
rect 7611 68188 7612 68228
rect 7652 68188 7653 68228
rect 7611 68179 7653 68188
rect 9579 68228 9621 68237
rect 9579 68188 9580 68228
rect 9620 68188 9621 68228
rect 9579 68179 9621 68188
rect 14139 68228 14181 68237
rect 14139 68188 14140 68228
rect 14180 68188 14181 68228
rect 14139 68179 14181 68188
rect 16587 68228 16629 68237
rect 16587 68188 16588 68228
rect 16628 68188 16629 68228
rect 16587 68179 16629 68188
rect 20379 68228 20421 68237
rect 20379 68188 20380 68228
rect 20420 68188 20421 68228
rect 20379 68179 20421 68188
rect 1152 68060 20452 68084
rect 1152 68020 4928 68060
rect 4968 68020 5010 68060
rect 5050 68020 5092 68060
rect 5132 68020 5174 68060
rect 5214 68020 5256 68060
rect 5296 68020 20048 68060
rect 20088 68020 20130 68060
rect 20170 68020 20212 68060
rect 20252 68020 20294 68060
rect 20334 68020 20376 68060
rect 20416 68020 20452 68060
rect 1152 67996 20452 68020
rect 16203 67892 16245 67901
rect 16203 67852 16204 67892
rect 16244 67852 16245 67892
rect 16203 67843 16245 67852
rect 1323 67724 1365 67733
rect 3034 67724 3092 67725
rect 1323 67684 1324 67724
rect 1364 67684 1365 67724
rect 1323 67675 1365 67684
rect 2571 67715 2613 67724
rect 2571 67675 2572 67715
rect 2612 67675 2613 67715
rect 3034 67684 3043 67724
rect 3083 67684 3092 67724
rect 3034 67683 3092 67684
rect 3147 67724 3189 67733
rect 3147 67684 3148 67724
rect 3188 67684 3189 67724
rect 3147 67675 3189 67684
rect 3531 67724 3573 67733
rect 5355 67724 5397 67733
rect 3531 67684 3532 67724
rect 3572 67684 3573 67724
rect 3531 67675 3573 67684
rect 4107 67715 4149 67724
rect 4107 67675 4108 67715
rect 4148 67675 4149 67715
rect 2571 67666 2613 67675
rect 4107 67666 4149 67675
rect 4587 67715 4629 67724
rect 4587 67675 4588 67715
rect 4628 67675 4629 67715
rect 5355 67684 5356 67724
rect 5396 67684 5397 67724
rect 5355 67675 5397 67684
rect 5643 67724 5685 67733
rect 7371 67724 7413 67733
rect 9483 67724 9525 67733
rect 11115 67724 11157 67733
rect 12747 67724 12789 67733
rect 14763 67724 14805 67733
rect 16971 67724 17013 67733
rect 18603 67724 18645 67733
rect 5643 67684 5644 67724
rect 5684 67684 5685 67724
rect 5643 67675 5685 67684
rect 6891 67715 6933 67724
rect 6891 67675 6892 67715
rect 6932 67675 6933 67715
rect 7371 67684 7372 67724
rect 7412 67684 7413 67724
rect 7371 67675 7413 67684
rect 8619 67715 8661 67724
rect 8619 67675 8620 67715
rect 8660 67675 8661 67715
rect 9483 67684 9484 67724
rect 9524 67684 9525 67724
rect 9483 67675 9525 67684
rect 10731 67715 10773 67724
rect 10731 67675 10732 67715
rect 10772 67675 10773 67715
rect 11115 67684 11116 67724
rect 11156 67684 11157 67724
rect 11115 67675 11157 67684
rect 12363 67715 12405 67724
rect 12363 67675 12364 67715
rect 12404 67675 12405 67715
rect 12747 67684 12748 67724
rect 12788 67684 12789 67724
rect 12747 67675 12789 67684
rect 13995 67715 14037 67724
rect 13995 67675 13996 67715
rect 14036 67675 14037 67715
rect 14763 67684 14764 67724
rect 14804 67684 14805 67724
rect 14763 67675 14805 67684
rect 16011 67715 16053 67724
rect 16011 67675 16012 67715
rect 16052 67675 16053 67715
rect 16971 67684 16972 67724
rect 17012 67684 17013 67724
rect 16971 67675 17013 67684
rect 18219 67715 18261 67724
rect 18219 67675 18220 67715
rect 18260 67675 18261 67715
rect 18603 67684 18604 67724
rect 18644 67684 18645 67724
rect 18603 67675 18645 67684
rect 19851 67715 19893 67724
rect 19851 67675 19852 67715
rect 19892 67675 19893 67715
rect 4587 67666 4629 67675
rect 6891 67666 6933 67675
rect 8619 67666 8661 67675
rect 10731 67666 10773 67675
rect 12363 67666 12405 67675
rect 13995 67666 14037 67675
rect 16011 67666 16053 67675
rect 18219 67666 18261 67675
rect 19851 67666 19893 67675
rect 3627 67640 3669 67649
rect 3627 67600 3628 67640
rect 3668 67600 3669 67640
rect 3627 67591 3669 67600
rect 5163 67640 5205 67649
rect 5163 67600 5164 67640
rect 5204 67600 5205 67640
rect 5163 67591 5205 67600
rect 9003 67640 9045 67649
rect 9003 67600 9004 67640
rect 9044 67600 9045 67640
rect 9003 67591 9045 67600
rect 9243 67640 9285 67649
rect 9243 67600 9244 67640
rect 9284 67600 9285 67640
rect 9243 67591 9285 67600
rect 14379 67640 14421 67649
rect 14379 67600 14380 67640
rect 14420 67600 14421 67640
rect 14379 67591 14421 67600
rect 16587 67640 16629 67649
rect 16587 67600 16588 67640
rect 16628 67600 16629 67640
rect 16587 67591 16629 67600
rect 16827 67640 16869 67649
rect 16827 67600 16828 67640
rect 16868 67600 16869 67640
rect 16827 67591 16869 67600
rect 4827 67556 4869 67565
rect 4827 67516 4828 67556
rect 4868 67516 4869 67556
rect 4827 67507 4869 67516
rect 5499 67556 5541 67565
rect 5499 67516 5500 67556
rect 5540 67516 5541 67556
rect 5499 67507 5541 67516
rect 14187 67556 14229 67565
rect 14187 67516 14188 67556
rect 14228 67516 14229 67556
rect 14187 67507 14229 67516
rect 2763 67472 2805 67481
rect 2763 67432 2764 67472
rect 2804 67432 2805 67472
rect 2763 67423 2805 67432
rect 4923 67472 4965 67481
rect 4923 67432 4924 67472
rect 4964 67432 4965 67472
rect 4923 67423 4965 67432
rect 7083 67472 7125 67481
rect 7083 67432 7084 67472
rect 7124 67432 7125 67472
rect 7083 67423 7125 67432
rect 8811 67472 8853 67481
rect 8811 67432 8812 67472
rect 8852 67432 8853 67472
rect 8811 67423 8853 67432
rect 10923 67472 10965 67481
rect 10923 67432 10924 67472
rect 10964 67432 10965 67472
rect 10923 67423 10965 67432
rect 12555 67472 12597 67481
rect 12555 67432 12556 67472
rect 12596 67432 12597 67472
rect 12555 67423 12597 67432
rect 14619 67472 14661 67481
rect 14619 67432 14620 67472
rect 14660 67432 14661 67472
rect 14619 67423 14661 67432
rect 18411 67472 18453 67481
rect 18411 67432 18412 67472
rect 18452 67432 18453 67472
rect 18411 67423 18453 67432
rect 20043 67472 20085 67481
rect 20043 67432 20044 67472
rect 20084 67432 20085 67472
rect 20043 67423 20085 67432
rect 1152 67304 20448 67328
rect 1152 67264 3688 67304
rect 3728 67264 3770 67304
rect 3810 67264 3852 67304
rect 3892 67264 3934 67304
rect 3974 67264 4016 67304
rect 4056 67264 18808 67304
rect 18848 67264 18890 67304
rect 18930 67264 18972 67304
rect 19012 67264 19054 67304
rect 19094 67264 19136 67304
rect 19176 67264 20448 67304
rect 1152 67240 20448 67264
rect 8955 67136 8997 67145
rect 8955 67096 8956 67136
rect 8996 67096 8997 67136
rect 8955 67087 8997 67096
rect 13371 67136 13413 67145
rect 13371 67096 13372 67136
rect 13412 67096 13413 67136
rect 13371 67087 13413 67096
rect 15483 67136 15525 67145
rect 15483 67096 15484 67136
rect 15524 67096 15525 67136
rect 15483 67087 15525 67096
rect 5211 67052 5253 67061
rect 5211 67012 5212 67052
rect 5252 67012 5253 67052
rect 5211 67003 5253 67012
rect 15867 67052 15909 67061
rect 15867 67012 15868 67052
rect 15908 67012 15909 67052
rect 15867 67003 15909 67012
rect 1419 66968 1461 66977
rect 1419 66928 1420 66968
rect 1460 66928 1461 66968
rect 1419 66919 1461 66928
rect 4971 66968 5013 66977
rect 4971 66928 4972 66968
rect 5012 66928 5013 66968
rect 4971 66919 5013 66928
rect 7563 66968 7605 66977
rect 7563 66928 7564 66968
rect 7604 66928 7605 66968
rect 7563 66919 7605 66928
rect 9195 66968 9237 66977
rect 9195 66928 9196 66968
rect 9236 66928 9237 66968
rect 9195 66919 9237 66928
rect 11691 66968 11733 66977
rect 11691 66928 11692 66968
rect 11732 66928 11733 66968
rect 11691 66919 11733 66928
rect 13131 66968 13173 66977
rect 13131 66928 13132 66968
rect 13172 66928 13173 66968
rect 13131 66919 13173 66928
rect 15243 66968 15285 66977
rect 15243 66928 15244 66968
rect 15284 66928 15285 66968
rect 15243 66919 15285 66928
rect 15627 66968 15669 66977
rect 15627 66928 15628 66968
rect 15668 66928 15669 66968
rect 15627 66919 15669 66928
rect 16011 66968 16053 66977
rect 16011 66928 16012 66968
rect 16052 66928 16053 66968
rect 16011 66919 16053 66928
rect 18603 66968 18645 66977
rect 18603 66928 18604 66968
rect 18644 66928 18645 66968
rect 18603 66919 18645 66928
rect 20235 66968 20277 66977
rect 20235 66928 20236 66968
rect 20276 66928 20277 66968
rect 20235 66919 20277 66928
rect 1707 66884 1749 66893
rect 1707 66844 1708 66884
rect 1748 66844 1749 66884
rect 1707 66835 1749 66844
rect 2947 66884 3005 66885
rect 2947 66844 2956 66884
rect 2996 66844 3005 66884
rect 2947 66843 3005 66844
rect 3523 66884 3581 66885
rect 3523 66844 3532 66884
rect 3572 66844 3581 66884
rect 3523 66843 3581 66844
rect 4779 66884 4821 66893
rect 4779 66844 4780 66884
rect 4820 66844 4821 66884
rect 4779 66835 4821 66844
rect 5355 66884 5397 66893
rect 5355 66844 5356 66884
rect 5396 66844 5397 66884
rect 5355 66835 5397 66844
rect 6595 66884 6653 66885
rect 6595 66844 6604 66884
rect 6644 66844 6653 66884
rect 6595 66843 6653 66844
rect 7066 66884 7124 66885
rect 7066 66844 7075 66884
rect 7115 66844 7124 66884
rect 7066 66843 7124 66844
rect 7179 66884 7221 66893
rect 7179 66844 7180 66884
rect 7220 66844 7221 66884
rect 7179 66835 7221 66844
rect 7659 66884 7701 66893
rect 7659 66844 7660 66884
rect 7700 66844 7701 66884
rect 7659 66835 7701 66844
rect 8131 66884 8189 66885
rect 8131 66844 8140 66884
rect 8180 66844 8189 66884
rect 8131 66843 8189 66844
rect 8650 66884 8708 66885
rect 8650 66844 8659 66884
rect 8699 66844 8708 66884
rect 8650 66843 8708 66844
rect 9483 66884 9525 66893
rect 9483 66844 9484 66884
rect 9524 66844 9525 66884
rect 9483 66835 9525 66844
rect 10723 66884 10781 66885
rect 10723 66844 10732 66884
rect 10772 66844 10781 66884
rect 10723 66843 10781 66844
rect 11194 66884 11252 66885
rect 11194 66844 11203 66884
rect 11243 66844 11252 66884
rect 11194 66843 11252 66844
rect 11307 66884 11349 66893
rect 11307 66844 11308 66884
rect 11348 66844 11349 66884
rect 11307 66835 11349 66844
rect 11787 66884 11829 66893
rect 11787 66844 11788 66884
rect 11828 66844 11829 66884
rect 11787 66835 11829 66844
rect 12259 66884 12317 66885
rect 12259 66844 12268 66884
rect 12308 66844 12317 66884
rect 12259 66843 12317 66844
rect 12747 66884 12805 66885
rect 12747 66844 12756 66884
rect 12796 66844 12805 66884
rect 12747 66843 12805 66844
rect 13611 66884 13653 66893
rect 13611 66844 13612 66884
rect 13652 66844 13653 66884
rect 13611 66835 13653 66844
rect 14851 66884 14909 66885
rect 14851 66844 14860 66884
rect 14900 66844 14909 66884
rect 14851 66843 14909 66844
rect 16395 66884 16437 66893
rect 16395 66844 16396 66884
rect 16436 66844 16437 66884
rect 16395 66835 16437 66844
rect 17635 66884 17693 66885
rect 17635 66844 17644 66884
rect 17684 66844 17693 66884
rect 17635 66843 17693 66844
rect 18106 66884 18164 66885
rect 18106 66844 18115 66884
rect 18155 66844 18164 66884
rect 18106 66843 18164 66844
rect 18219 66884 18261 66893
rect 18219 66844 18220 66884
rect 18260 66844 18261 66884
rect 18219 66835 18261 66844
rect 18699 66884 18741 66893
rect 18699 66844 18700 66884
rect 18740 66844 18741 66884
rect 18699 66835 18741 66844
rect 19171 66884 19229 66885
rect 19171 66844 19180 66884
rect 19220 66844 19229 66884
rect 19171 66843 19229 66844
rect 19690 66884 19748 66885
rect 19690 66844 19699 66884
rect 19739 66844 19748 66884
rect 19690 66843 19748 66844
rect 6795 66800 6837 66809
rect 6795 66760 6796 66800
rect 6836 66760 6837 66800
rect 6795 66751 6837 66760
rect 1179 66716 1221 66725
rect 1179 66676 1180 66716
rect 1220 66676 1221 66716
rect 1179 66667 1221 66676
rect 3147 66716 3189 66725
rect 3147 66676 3148 66716
rect 3188 66676 3189 66716
rect 3147 66667 3189 66676
rect 3339 66716 3381 66725
rect 3339 66676 3340 66716
rect 3380 66676 3381 66716
rect 3339 66667 3381 66676
rect 8811 66716 8853 66725
rect 8811 66676 8812 66716
rect 8852 66676 8853 66716
rect 8811 66667 8853 66676
rect 10923 66716 10965 66725
rect 10923 66676 10924 66716
rect 10964 66676 10965 66716
rect 10923 66667 10965 66676
rect 12939 66716 12981 66725
rect 12939 66676 12940 66716
rect 12980 66676 12981 66716
rect 12939 66667 12981 66676
rect 15051 66716 15093 66725
rect 15051 66676 15052 66716
rect 15092 66676 15093 66716
rect 15051 66667 15093 66676
rect 16251 66716 16293 66725
rect 16251 66676 16252 66716
rect 16292 66676 16293 66716
rect 16251 66667 16293 66676
rect 17835 66716 17877 66725
rect 17835 66676 17836 66716
rect 17876 66676 17877 66716
rect 17835 66667 17877 66676
rect 19851 66716 19893 66725
rect 19851 66676 19852 66716
rect 19892 66676 19893 66716
rect 19851 66667 19893 66676
rect 19995 66716 20037 66725
rect 19995 66676 19996 66716
rect 20036 66676 20037 66716
rect 19995 66667 20037 66676
rect 1152 66548 20452 66572
rect 1152 66508 4928 66548
rect 4968 66508 5010 66548
rect 5050 66508 5092 66548
rect 5132 66508 5174 66548
rect 5214 66508 5256 66548
rect 5296 66508 20048 66548
rect 20088 66508 20130 66548
rect 20170 66508 20212 66548
rect 20252 66508 20294 66548
rect 20334 66508 20376 66548
rect 20416 66508 20452 66548
rect 1152 66484 20452 66508
rect 4395 66380 4437 66389
rect 4395 66340 4396 66380
rect 4436 66340 4437 66380
rect 4395 66331 4437 66340
rect 17115 66380 17157 66389
rect 17115 66340 17116 66380
rect 17156 66340 17157 66380
rect 17115 66331 17157 66340
rect 20331 66380 20373 66389
rect 20331 66340 20332 66380
rect 20372 66340 20373 66380
rect 20331 66331 20373 66340
rect 6843 66296 6885 66305
rect 6843 66256 6844 66296
rect 6884 66256 6885 66296
rect 6843 66247 6885 66256
rect 16731 66296 16773 66305
rect 16731 66256 16732 66296
rect 16772 66256 16773 66296
rect 16731 66247 16773 66256
rect 2637 66212 2679 66221
rect 2637 66172 2638 66212
rect 2678 66172 2679 66212
rect 2637 66163 2679 66172
rect 2763 66212 2805 66221
rect 2763 66172 2764 66212
rect 2804 66172 2805 66212
rect 2763 66163 2805 66172
rect 3147 66212 3189 66221
rect 4779 66212 4821 66221
rect 7947 66212 7989 66221
rect 9867 66212 9909 66221
rect 13035 66212 13077 66221
rect 14842 66212 14900 66213
rect 3147 66172 3148 66212
rect 3188 66172 3189 66212
rect 3147 66163 3189 66172
rect 3723 66203 3765 66212
rect 3723 66163 3724 66203
rect 3764 66163 3765 66203
rect 3723 66154 3765 66163
rect 4203 66203 4245 66212
rect 4203 66163 4204 66203
rect 4244 66163 4245 66203
rect 4779 66172 4780 66212
rect 4820 66172 4821 66212
rect 4779 66163 4821 66172
rect 6027 66203 6069 66212
rect 6027 66163 6028 66203
rect 6068 66163 6069 66203
rect 7947 66172 7948 66212
rect 7988 66172 7989 66212
rect 7947 66163 7989 66172
rect 9195 66203 9237 66212
rect 9195 66163 9196 66203
rect 9236 66163 9237 66203
rect 9867 66172 9868 66212
rect 9908 66172 9909 66212
rect 9867 66163 9909 66172
rect 11115 66203 11157 66212
rect 11115 66163 11116 66203
rect 11156 66163 11157 66203
rect 13035 66172 13036 66212
rect 13076 66172 13077 66212
rect 13035 66163 13077 66172
rect 14283 66203 14325 66212
rect 14283 66163 14284 66203
rect 14324 66163 14325 66203
rect 14842 66172 14851 66212
rect 14891 66172 14900 66212
rect 14842 66171 14900 66172
rect 14955 66212 14997 66221
rect 14955 66172 14956 66212
rect 14996 66172 14997 66212
rect 14955 66163 14997 66172
rect 15339 66212 15381 66221
rect 18202 66212 18260 66213
rect 15339 66172 15340 66212
rect 15380 66172 15381 66212
rect 15339 66163 15381 66172
rect 15915 66203 15957 66212
rect 15915 66163 15916 66203
rect 15956 66163 15957 66203
rect 4203 66154 4245 66163
rect 6027 66154 6069 66163
rect 9195 66154 9237 66163
rect 11115 66154 11157 66163
rect 14283 66154 14325 66163
rect 15915 66154 15957 66163
rect 16395 66203 16437 66212
rect 16395 66163 16396 66203
rect 16436 66163 16437 66203
rect 18202 66172 18211 66212
rect 18251 66172 18260 66212
rect 18202 66171 18260 66172
rect 18315 66212 18357 66221
rect 18315 66172 18316 66212
rect 18356 66172 18357 66212
rect 18315 66163 18357 66172
rect 18699 66212 18741 66221
rect 18699 66172 18700 66212
rect 18740 66172 18741 66212
rect 18699 66163 18741 66172
rect 19275 66203 19317 66212
rect 19275 66163 19276 66203
rect 19316 66163 19317 66203
rect 16395 66154 16437 66163
rect 19275 66154 19317 66163
rect 19755 66203 19797 66212
rect 19755 66163 19756 66203
rect 19796 66163 19797 66203
rect 19755 66154 19797 66163
rect 1419 66128 1461 66137
rect 1419 66088 1420 66128
rect 1460 66088 1461 66128
rect 1419 66079 1461 66088
rect 1803 66128 1845 66137
rect 1803 66088 1804 66128
rect 1844 66088 1845 66128
rect 1803 66079 1845 66088
rect 2187 66128 2229 66137
rect 2187 66088 2188 66128
rect 2228 66088 2229 66128
rect 2187 66079 2229 66088
rect 3243 66128 3285 66137
rect 3243 66088 3244 66128
rect 3284 66088 3285 66128
rect 3243 66079 3285 66088
rect 6634 66128 6692 66129
rect 6634 66088 6643 66128
rect 6683 66088 6692 66128
rect 6634 66087 6692 66088
rect 6987 66128 7029 66137
rect 6987 66088 6988 66128
rect 7028 66088 7029 66128
rect 6987 66079 7029 66088
rect 7563 66128 7605 66137
rect 7563 66088 7564 66128
rect 7604 66088 7605 66128
rect 7563 66079 7605 66088
rect 12843 66128 12885 66137
rect 12843 66088 12844 66128
rect 12884 66088 12885 66128
rect 12843 66079 12885 66088
rect 15435 66128 15477 66137
rect 15435 66088 15436 66128
rect 15476 66088 15477 66128
rect 15435 66079 15477 66088
rect 16618 66128 16676 66129
rect 16618 66088 16627 66128
rect 16667 66088 16676 66128
rect 16618 66087 16676 66088
rect 16971 66128 17013 66137
rect 16971 66088 16972 66128
rect 17012 66088 17013 66128
rect 16971 66079 17013 66088
rect 17355 66128 17397 66137
rect 17355 66088 17356 66128
rect 17396 66088 17397 66128
rect 17355 66079 17397 66088
rect 17739 66128 17781 66137
rect 17739 66088 17740 66128
rect 17780 66088 17781 66128
rect 17739 66079 17781 66088
rect 18795 66128 18837 66137
rect 18795 66088 18796 66128
rect 18836 66088 18837 66128
rect 18795 66079 18837 66088
rect 7227 66044 7269 66053
rect 7227 66004 7228 66044
rect 7268 66004 7269 66044
rect 7227 65995 7269 66004
rect 14475 66044 14517 66053
rect 14475 66004 14476 66044
rect 14516 66004 14517 66044
rect 14475 65995 14517 66004
rect 19995 66044 20037 66053
rect 19995 66004 19996 66044
rect 20036 66004 20037 66044
rect 19995 65995 20037 66004
rect 1179 65960 1221 65969
rect 1179 65920 1180 65960
rect 1220 65920 1221 65960
rect 1179 65911 1221 65920
rect 1563 65960 1605 65969
rect 1563 65920 1564 65960
rect 1604 65920 1605 65960
rect 1563 65911 1605 65920
rect 1947 65960 1989 65969
rect 1947 65920 1948 65960
rect 1988 65920 1989 65960
rect 1947 65911 1989 65920
rect 6219 65960 6261 65969
rect 6219 65920 6220 65960
rect 6260 65920 6261 65960
rect 6219 65911 6261 65920
rect 7323 65960 7365 65969
rect 7323 65920 7324 65960
rect 7364 65920 7365 65960
rect 7323 65911 7365 65920
rect 9387 65960 9429 65969
rect 9387 65920 9388 65960
rect 9428 65920 9429 65960
rect 9387 65911 9429 65920
rect 11307 65960 11349 65969
rect 11307 65920 11308 65960
rect 11348 65920 11349 65960
rect 11307 65911 11349 65920
rect 12603 65960 12645 65969
rect 12603 65920 12604 65960
rect 12644 65920 12645 65960
rect 12603 65911 12645 65920
rect 17979 65960 18021 65969
rect 17979 65920 17980 65960
rect 18020 65920 18021 65960
rect 17979 65911 18021 65920
rect 1152 65792 20448 65816
rect 1152 65752 3688 65792
rect 3728 65752 3770 65792
rect 3810 65752 3852 65792
rect 3892 65752 3934 65792
rect 3974 65752 4016 65792
rect 4056 65752 18808 65792
rect 18848 65752 18890 65792
rect 18930 65752 18972 65792
rect 19012 65752 19054 65792
rect 19094 65752 19136 65792
rect 19176 65752 20448 65792
rect 1152 65728 20448 65752
rect 3099 65624 3141 65633
rect 3099 65584 3100 65624
rect 3140 65584 3141 65624
rect 3099 65575 3141 65584
rect 12027 65624 12069 65633
rect 12027 65584 12028 65624
rect 12068 65584 12069 65624
rect 12027 65575 12069 65584
rect 16906 65624 16964 65625
rect 16906 65584 16915 65624
rect 16955 65584 16964 65624
rect 16906 65583 16964 65584
rect 20139 65624 20181 65633
rect 20139 65584 20140 65624
rect 20180 65584 20181 65624
rect 20139 65575 20181 65584
rect 17067 65540 17109 65549
rect 17067 65500 17068 65540
rect 17108 65500 17109 65540
rect 17067 65491 17109 65500
rect 3339 65456 3381 65465
rect 3339 65416 3340 65456
rect 3380 65416 3381 65456
rect 3339 65407 3381 65416
rect 3723 65456 3765 65465
rect 3723 65416 3724 65456
rect 3764 65416 3765 65456
rect 3723 65407 3765 65416
rect 4299 65456 4341 65465
rect 4299 65416 4300 65456
rect 4340 65416 4341 65456
rect 4299 65407 4341 65416
rect 9963 65456 10005 65465
rect 9963 65416 9964 65456
rect 10004 65416 10005 65456
rect 9963 65407 10005 65416
rect 11787 65456 11829 65465
rect 11787 65416 11788 65456
rect 11828 65416 11829 65456
rect 11787 65407 11829 65416
rect 12123 65456 12165 65465
rect 12123 65416 12124 65456
rect 12164 65416 12165 65456
rect 12123 65407 12165 65416
rect 12363 65456 12405 65465
rect 12363 65416 12364 65456
rect 12404 65416 12405 65456
rect 12363 65407 12405 65416
rect 13131 65456 13173 65465
rect 13131 65416 13132 65456
rect 13172 65416 13173 65456
rect 13131 65407 13173 65416
rect 14410 65456 14468 65457
rect 14410 65416 14419 65456
rect 14459 65416 14468 65456
rect 14410 65415 14468 65416
rect 14763 65456 14805 65465
rect 14763 65416 14764 65456
rect 14804 65416 14805 65456
rect 14763 65407 14805 65416
rect 15627 65456 15669 65465
rect 15627 65416 15628 65456
rect 15668 65416 15669 65456
rect 15627 65407 15669 65416
rect 1515 65372 1557 65381
rect 1515 65332 1516 65372
rect 1556 65332 1557 65372
rect 1515 65323 1557 65332
rect 2763 65372 2821 65373
rect 2763 65332 2772 65372
rect 2812 65332 2821 65372
rect 2763 65331 2821 65332
rect 4491 65372 4533 65381
rect 4491 65332 4492 65372
rect 4532 65332 4533 65372
rect 4491 65323 4533 65332
rect 5731 65372 5789 65373
rect 5731 65332 5740 65372
rect 5780 65332 5789 65372
rect 5731 65331 5789 65332
rect 6123 65372 6165 65381
rect 6123 65332 6124 65372
rect 6164 65332 6165 65372
rect 6123 65323 6165 65332
rect 7363 65372 7421 65373
rect 7363 65332 7372 65372
rect 7412 65332 7421 65372
rect 7363 65331 7421 65332
rect 7755 65372 7797 65381
rect 7755 65332 7756 65372
rect 7796 65332 7797 65372
rect 7755 65323 7797 65332
rect 8995 65372 9053 65373
rect 8995 65332 9004 65372
rect 9044 65332 9053 65372
rect 8995 65331 9053 65332
rect 9466 65372 9524 65373
rect 9466 65332 9475 65372
rect 9515 65332 9524 65372
rect 9466 65331 9524 65332
rect 9579 65372 9621 65381
rect 9579 65332 9580 65372
rect 9620 65332 9621 65372
rect 9579 65323 9621 65332
rect 10059 65372 10101 65381
rect 10059 65332 10060 65372
rect 10100 65332 10101 65372
rect 10059 65323 10101 65332
rect 10531 65372 10589 65373
rect 10531 65332 10540 65372
rect 10580 65332 10589 65372
rect 10531 65331 10589 65332
rect 11019 65372 11077 65373
rect 11019 65332 11028 65372
rect 11068 65332 11077 65372
rect 11019 65331 11077 65332
rect 12634 65372 12692 65373
rect 12634 65332 12643 65372
rect 12683 65332 12692 65372
rect 12634 65331 12692 65332
rect 12747 65372 12789 65381
rect 12747 65332 12748 65372
rect 12788 65332 12789 65372
rect 12747 65323 12789 65332
rect 13227 65372 13269 65381
rect 13227 65332 13228 65372
rect 13268 65332 13269 65372
rect 13227 65323 13269 65332
rect 13699 65372 13757 65373
rect 13699 65332 13708 65372
rect 13748 65332 13757 65372
rect 13699 65331 13757 65332
rect 14187 65372 14245 65373
rect 14187 65332 14196 65372
rect 14236 65332 14245 65372
rect 14187 65331 14245 65332
rect 15117 65372 15159 65381
rect 15117 65332 15118 65372
rect 15158 65332 15159 65372
rect 15117 65323 15159 65332
rect 15243 65371 15285 65380
rect 15243 65331 15244 65371
rect 15284 65331 15285 65371
rect 15243 65322 15285 65331
rect 15723 65372 15765 65381
rect 15723 65332 15724 65372
rect 15764 65332 15765 65372
rect 15723 65323 15765 65332
rect 16195 65372 16253 65373
rect 16195 65332 16204 65372
rect 16244 65332 16253 65372
rect 16195 65331 16253 65332
rect 16683 65372 16741 65373
rect 16683 65332 16692 65372
rect 16732 65332 16741 65372
rect 16683 65331 16741 65332
rect 17251 65372 17309 65373
rect 17251 65332 17260 65372
rect 17300 65332 17309 65372
rect 17251 65331 17309 65332
rect 18507 65372 18549 65381
rect 18507 65332 18508 65372
rect 18548 65332 18549 65372
rect 18507 65323 18549 65332
rect 18699 65372 18741 65381
rect 18699 65332 18700 65372
rect 18740 65332 18741 65372
rect 18699 65323 18741 65332
rect 19939 65372 19997 65373
rect 19939 65332 19948 65372
rect 19988 65332 19997 65372
rect 19939 65331 19997 65332
rect 3483 65288 3525 65297
rect 3483 65248 3484 65288
rect 3524 65248 3525 65288
rect 3483 65239 3525 65248
rect 14523 65288 14565 65297
rect 14523 65248 14524 65288
rect 14564 65248 14565 65288
rect 14523 65239 14565 65248
rect 2955 65204 2997 65213
rect 2955 65164 2956 65204
rect 2996 65164 2997 65204
rect 2955 65155 2997 65164
rect 4059 65204 4101 65213
rect 4059 65164 4060 65204
rect 4100 65164 4101 65204
rect 4059 65155 4101 65164
rect 5931 65204 5973 65213
rect 5931 65164 5932 65204
rect 5972 65164 5973 65204
rect 5931 65155 5973 65164
rect 7563 65204 7605 65213
rect 7563 65164 7564 65204
rect 7604 65164 7605 65204
rect 7563 65155 7605 65164
rect 9195 65204 9237 65213
rect 9195 65164 9196 65204
rect 9236 65164 9237 65204
rect 9195 65155 9237 65164
rect 11211 65204 11253 65213
rect 11211 65164 11212 65204
rect 11252 65164 11253 65204
rect 11211 65155 11253 65164
rect 12027 65204 12069 65213
rect 12027 65164 12028 65204
rect 12068 65164 12069 65204
rect 12027 65155 12069 65164
rect 1152 65036 20452 65060
rect 1152 64996 4928 65036
rect 4968 64996 5010 65036
rect 5050 64996 5092 65036
rect 5132 64996 5174 65036
rect 5214 64996 5256 65036
rect 5296 64996 20048 65036
rect 20088 64996 20130 65036
rect 20170 64996 20212 65036
rect 20252 64996 20294 65036
rect 20334 64996 20376 65036
rect 20416 64996 20452 65036
rect 1152 64972 20452 64996
rect 14091 64868 14133 64877
rect 14091 64828 14092 64868
rect 14132 64828 14133 64868
rect 14091 64819 14133 64828
rect 16107 64868 16149 64877
rect 16107 64828 16108 64868
rect 16148 64828 16149 64868
rect 16107 64819 16149 64828
rect 2170 64784 2228 64785
rect 2170 64744 2179 64784
rect 2219 64744 2228 64784
rect 2170 64743 2228 64744
rect 8331 64784 8373 64793
rect 8331 64744 8332 64784
rect 8372 64744 8373 64784
rect 8331 64735 8373 64744
rect 14523 64784 14565 64793
rect 14523 64744 14524 64784
rect 14564 64744 14565 64784
rect 14523 64735 14565 64744
rect 2362 64700 2420 64701
rect 3339 64700 3381 64709
rect 2362 64660 2371 64700
rect 2411 64660 2420 64700
rect 2362 64659 2420 64660
rect 2859 64691 2901 64700
rect 2859 64651 2860 64691
rect 2900 64651 2901 64691
rect 3339 64660 3340 64700
rect 3380 64660 3381 64700
rect 3339 64651 3381 64660
rect 3819 64700 3861 64709
rect 3819 64660 3820 64700
rect 3860 64660 3861 64700
rect 3819 64651 3861 64660
rect 3929 64700 3987 64701
rect 3929 64660 3938 64700
rect 3978 64660 3987 64700
rect 3929 64659 3987 64660
rect 4282 64700 4340 64701
rect 4282 64660 4291 64700
rect 4331 64660 4340 64700
rect 4282 64659 4340 64660
rect 4395 64700 4437 64709
rect 4395 64660 4396 64700
rect 4436 64660 4437 64700
rect 4395 64651 4437 64660
rect 4779 64700 4821 64709
rect 6891 64700 6933 64709
rect 8506 64700 8564 64701
rect 4779 64660 4780 64700
rect 4820 64660 4821 64700
rect 4779 64651 4821 64660
rect 5355 64691 5397 64700
rect 5355 64651 5356 64691
rect 5396 64651 5397 64691
rect 2859 64642 2901 64651
rect 5355 64642 5397 64651
rect 5835 64691 5877 64700
rect 5835 64651 5836 64691
rect 5876 64651 5877 64691
rect 6891 64660 6892 64700
rect 6932 64660 6933 64700
rect 6891 64651 6933 64660
rect 8139 64691 8181 64700
rect 8139 64651 8140 64691
rect 8180 64651 8181 64691
rect 8506 64660 8515 64700
rect 8555 64660 8564 64700
rect 8506 64659 8564 64660
rect 8811 64700 8853 64709
rect 8811 64660 8812 64700
rect 8852 64660 8853 64700
rect 8811 64651 8853 64660
rect 9099 64700 9141 64709
rect 9099 64660 9100 64700
rect 9140 64660 9141 64700
rect 9099 64651 9141 64660
rect 9562 64700 9620 64701
rect 9562 64660 9571 64700
rect 9611 64660 9620 64700
rect 9562 64659 9620 64660
rect 9680 64700 9722 64709
rect 9680 64660 9681 64700
rect 9721 64660 9722 64700
rect 9680 64651 9722 64660
rect 10059 64700 10101 64709
rect 12651 64700 12693 64709
rect 14667 64700 14709 64709
rect 16587 64700 16629 64709
rect 18315 64700 18357 64709
rect 10059 64660 10060 64700
rect 10100 64660 10101 64700
rect 10059 64651 10101 64660
rect 10635 64691 10677 64700
rect 10635 64651 10636 64691
rect 10676 64651 10677 64691
rect 5835 64642 5877 64651
rect 8139 64642 8181 64651
rect 10635 64642 10677 64651
rect 11115 64691 11157 64700
rect 11115 64651 11116 64691
rect 11156 64651 11157 64691
rect 12651 64660 12652 64700
rect 12692 64660 12693 64700
rect 12651 64651 12693 64660
rect 13899 64691 13941 64700
rect 13899 64651 13900 64691
rect 13940 64651 13941 64691
rect 14667 64660 14668 64700
rect 14708 64660 14709 64700
rect 14667 64651 14709 64660
rect 15915 64691 15957 64700
rect 15915 64651 15916 64691
rect 15956 64651 15957 64691
rect 16587 64660 16588 64700
rect 16628 64660 16629 64700
rect 16587 64651 16629 64660
rect 17835 64691 17877 64700
rect 17835 64651 17836 64691
rect 17876 64651 17877 64691
rect 18315 64660 18316 64700
rect 18356 64660 18357 64700
rect 18315 64651 18357 64660
rect 19563 64691 19605 64700
rect 19563 64651 19564 64691
rect 19604 64651 19605 64691
rect 11115 64642 11157 64651
rect 13899 64642 13941 64651
rect 15915 64642 15957 64651
rect 17835 64642 17877 64651
rect 19563 64642 19605 64651
rect 1419 64616 1461 64625
rect 1419 64576 1420 64616
rect 1460 64576 1461 64616
rect 1419 64567 1461 64576
rect 1803 64616 1845 64625
rect 1803 64576 1804 64616
rect 1844 64576 1845 64616
rect 1803 64567 1845 64576
rect 3435 64616 3477 64625
rect 3435 64576 3436 64616
rect 3476 64576 3477 64616
rect 3435 64567 3477 64576
rect 4875 64616 4917 64625
rect 4875 64576 4876 64616
rect 4916 64576 4917 64616
rect 4875 64567 4917 64576
rect 6058 64616 6116 64617
rect 6058 64576 6067 64616
rect 6107 64576 6116 64616
rect 6058 64575 6116 64576
rect 6411 64616 6453 64625
rect 6411 64576 6412 64616
rect 6452 64576 6453 64616
rect 6411 64567 6453 64576
rect 10155 64616 10197 64625
rect 10155 64576 10156 64616
rect 10196 64576 10197 64616
rect 10155 64567 10197 64576
rect 12267 64616 12309 64625
rect 12267 64576 12268 64616
rect 12308 64576 12309 64616
rect 12267 64567 12309 64576
rect 12507 64616 12549 64625
rect 12507 64576 12508 64616
rect 12548 64576 12549 64616
rect 12507 64567 12549 64576
rect 14283 64616 14325 64625
rect 14283 64576 14284 64616
rect 14324 64576 14325 64616
rect 14283 64567 14325 64576
rect 20139 64616 20181 64625
rect 20139 64576 20140 64616
rect 20180 64576 20181 64616
rect 20139 64567 20181 64576
rect 6171 64532 6213 64541
rect 6171 64492 6172 64532
rect 6212 64492 6213 64532
rect 6171 64483 6213 64492
rect 8955 64532 8997 64541
rect 8955 64492 8956 64532
rect 8996 64492 8997 64532
rect 8955 64483 8997 64492
rect 1179 64448 1221 64457
rect 1179 64408 1180 64448
rect 1220 64408 1221 64448
rect 1179 64399 1221 64408
rect 1563 64448 1605 64457
rect 1563 64408 1564 64448
rect 1604 64408 1605 64448
rect 1563 64399 1605 64408
rect 8811 64448 8853 64457
rect 8811 64408 8812 64448
rect 8852 64408 8853 64448
rect 8811 64399 8853 64408
rect 11338 64448 11396 64449
rect 11338 64408 11347 64448
rect 11387 64408 11396 64448
rect 11338 64407 11396 64408
rect 18027 64448 18069 64457
rect 18027 64408 18028 64448
rect 18068 64408 18069 64448
rect 18027 64399 18069 64408
rect 19755 64448 19797 64457
rect 19755 64408 19756 64448
rect 19796 64408 19797 64448
rect 19755 64399 19797 64408
rect 20379 64448 20421 64457
rect 20379 64408 20380 64448
rect 20420 64408 20421 64448
rect 20379 64399 20421 64408
rect 1152 64280 20448 64304
rect 1152 64240 3688 64280
rect 3728 64240 3770 64280
rect 3810 64240 3852 64280
rect 3892 64240 3934 64280
rect 3974 64240 4016 64280
rect 4056 64240 18808 64280
rect 18848 64240 18890 64280
rect 18930 64240 18972 64280
rect 19012 64240 19054 64280
rect 19094 64240 19136 64280
rect 19176 64240 20448 64280
rect 1152 64216 20448 64240
rect 5691 64112 5733 64121
rect 5691 64072 5692 64112
rect 5732 64072 5733 64112
rect 5691 64063 5733 64072
rect 9435 64112 9477 64121
rect 9435 64072 9436 64112
rect 9476 64072 9477 64112
rect 9435 64063 9477 64072
rect 15003 64112 15045 64121
rect 15003 64072 15004 64112
rect 15044 64072 15045 64112
rect 15003 64063 15045 64072
rect 19995 64112 20037 64121
rect 19995 64072 19996 64112
rect 20036 64072 20037 64112
rect 19995 64063 20037 64072
rect 2955 64028 2997 64037
rect 2955 63988 2956 64028
rect 2996 63988 2997 64028
rect 2955 63979 2997 63988
rect 6075 64028 6117 64037
rect 6075 63988 6076 64028
rect 6116 63988 6117 64028
rect 6075 63979 6117 63988
rect 15483 64028 15525 64037
rect 15483 63988 15484 64028
rect 15524 63988 15525 64028
rect 15483 63979 15525 63988
rect 3339 63944 3381 63953
rect 3339 63904 3340 63944
rect 3380 63904 3381 63944
rect 3339 63895 3381 63904
rect 3723 63944 3765 63953
rect 3723 63904 3724 63944
rect 3764 63904 3765 63944
rect 3723 63895 3765 63904
rect 5931 63944 5973 63953
rect 5931 63904 5932 63944
rect 5972 63904 5973 63944
rect 5931 63895 5973 63904
rect 6315 63944 6357 63953
rect 6315 63904 6316 63944
rect 6356 63904 6357 63944
rect 6315 63895 6357 63904
rect 6699 63944 6741 63953
rect 6699 63904 6700 63944
rect 6740 63904 6741 63944
rect 6699 63895 6741 63904
rect 9082 63944 9140 63945
rect 9082 63904 9091 63944
rect 9131 63904 9140 63944
rect 9082 63903 9140 63904
rect 9675 63944 9717 63953
rect 9675 63904 9676 63944
rect 9716 63904 9717 63944
rect 9675 63895 9717 63904
rect 11691 63944 11733 63953
rect 11691 63904 11692 63944
rect 11732 63904 11733 63944
rect 11691 63895 11733 63904
rect 12555 63944 12597 63953
rect 12555 63904 12556 63944
rect 12596 63904 12597 63944
rect 12555 63895 12597 63904
rect 14571 63944 14613 63953
rect 14571 63904 14572 63944
rect 14612 63904 14613 63944
rect 14571 63895 14613 63904
rect 14763 63944 14805 63953
rect 14763 63904 14764 63944
rect 14804 63904 14805 63944
rect 14763 63895 14805 63904
rect 15147 63944 15189 63953
rect 15147 63904 15148 63944
rect 15188 63904 15189 63944
rect 15147 63895 15189 63904
rect 15723 63944 15765 63953
rect 15723 63904 15724 63944
rect 15764 63904 15765 63944
rect 15723 63895 15765 63904
rect 16203 63944 16245 63953
rect 16203 63904 16204 63944
rect 16244 63904 16245 63944
rect 16203 63895 16245 63904
rect 18603 63944 18645 63953
rect 18603 63904 18604 63944
rect 18644 63904 18645 63944
rect 18603 63895 18645 63904
rect 20235 63944 20277 63953
rect 20235 63904 20236 63944
rect 20276 63904 20277 63944
rect 20235 63895 20277 63904
rect 1515 63860 1557 63869
rect 1515 63820 1516 63860
rect 1556 63820 1557 63860
rect 1515 63811 1557 63820
rect 2755 63860 2813 63861
rect 2755 63820 2764 63860
rect 2804 63820 2813 63860
rect 2755 63819 2813 63820
rect 3915 63860 3957 63869
rect 3915 63820 3916 63860
rect 3956 63820 3957 63860
rect 3915 63811 3957 63820
rect 5155 63860 5213 63861
rect 5155 63820 5164 63860
rect 5204 63820 5213 63860
rect 5155 63819 5213 63820
rect 6891 63860 6933 63869
rect 6891 63820 6892 63860
rect 6932 63820 6933 63860
rect 6891 63811 6933 63820
rect 8131 63860 8189 63861
rect 8131 63820 8140 63860
rect 8180 63820 8189 63860
rect 8131 63819 8189 63820
rect 8506 63860 8564 63861
rect 8506 63820 8515 63860
rect 8555 63820 8564 63860
rect 8506 63819 8564 63820
rect 8950 63860 8992 63869
rect 8950 63820 8951 63860
rect 8991 63820 8992 63860
rect 8950 63811 8992 63820
rect 9195 63860 9237 63869
rect 9195 63820 9196 63860
rect 9236 63820 9237 63860
rect 9195 63811 9237 63820
rect 10059 63860 10101 63869
rect 10059 63820 10060 63860
rect 10100 63820 10101 63860
rect 10059 63811 10101 63820
rect 11299 63860 11357 63861
rect 11299 63820 11308 63860
rect 11348 63820 11357 63860
rect 11299 63819 11357 63820
rect 12747 63860 12789 63869
rect 12747 63820 12748 63860
rect 12788 63820 12789 63860
rect 12747 63811 12789 63820
rect 13987 63860 14045 63861
rect 13987 63820 13996 63860
rect 14036 63820 14045 63860
rect 13987 63819 14045 63820
rect 16395 63860 16437 63869
rect 16395 63820 16396 63860
rect 16436 63820 16437 63860
rect 16395 63811 16437 63820
rect 17635 63860 17693 63861
rect 17635 63820 17644 63860
rect 17684 63820 17693 63860
rect 17635 63819 17693 63820
rect 18106 63860 18164 63861
rect 18106 63820 18115 63860
rect 18155 63820 18164 63860
rect 18106 63819 18164 63820
rect 18219 63860 18261 63869
rect 18219 63820 18220 63860
rect 18260 63820 18261 63860
rect 18219 63811 18261 63820
rect 18699 63860 18741 63869
rect 18699 63820 18700 63860
rect 18740 63820 18741 63860
rect 18699 63811 18741 63820
rect 19171 63860 19229 63861
rect 19171 63820 19180 63860
rect 19220 63820 19229 63860
rect 19171 63819 19229 63820
rect 19663 63860 19721 63861
rect 19663 63820 19672 63860
rect 19712 63820 19721 63860
rect 19663 63819 19721 63820
rect 3099 63776 3141 63785
rect 3099 63736 3100 63776
rect 3140 63736 3141 63776
rect 3099 63727 3141 63736
rect 6459 63776 6501 63785
rect 6459 63736 6460 63776
rect 6500 63736 6501 63776
rect 6459 63727 6501 63736
rect 8825 63776 8867 63785
rect 8825 63736 8826 63776
rect 8866 63736 8867 63776
rect 8825 63727 8867 63736
rect 11931 63776 11973 63785
rect 11931 63736 11932 63776
rect 11972 63736 11973 63776
rect 11931 63727 11973 63736
rect 14331 63776 14373 63785
rect 14331 63736 14332 63776
rect 14372 63736 14373 63776
rect 14331 63727 14373 63736
rect 15387 63776 15429 63785
rect 15387 63736 15388 63776
rect 15428 63736 15429 63776
rect 15387 63727 15429 63736
rect 17835 63776 17877 63785
rect 17835 63736 17836 63776
rect 17876 63736 17877 63776
rect 17835 63727 17877 63736
rect 3483 63692 3525 63701
rect 3483 63652 3484 63692
rect 3524 63652 3525 63692
rect 3483 63643 3525 63652
rect 5355 63692 5397 63701
rect 5355 63652 5356 63692
rect 5396 63652 5397 63692
rect 5355 63643 5397 63652
rect 8331 63692 8373 63701
rect 8331 63652 8332 63692
rect 8372 63652 8373 63692
rect 8331 63643 8373 63652
rect 8602 63692 8660 63693
rect 8602 63652 8611 63692
rect 8651 63652 8660 63692
rect 8602 63651 8660 63652
rect 8715 63692 8757 63701
rect 8715 63652 8716 63692
rect 8756 63652 8757 63692
rect 8715 63643 8757 63652
rect 9274 63692 9332 63693
rect 9274 63652 9283 63692
rect 9323 63652 9332 63692
rect 9274 63651 9332 63652
rect 11499 63692 11541 63701
rect 11499 63652 11500 63692
rect 11540 63652 11541 63692
rect 11499 63643 11541 63652
rect 12315 63692 12357 63701
rect 12315 63652 12316 63692
rect 12356 63652 12357 63692
rect 12315 63643 12357 63652
rect 14187 63692 14229 63701
rect 14187 63652 14188 63692
rect 14228 63652 14229 63692
rect 14187 63643 14229 63652
rect 15963 63692 16005 63701
rect 15963 63652 15964 63692
rect 16004 63652 16005 63692
rect 15963 63643 16005 63652
rect 19851 63692 19893 63701
rect 19851 63652 19852 63692
rect 19892 63652 19893 63692
rect 19851 63643 19893 63652
rect 1152 63524 20452 63548
rect 1152 63484 4928 63524
rect 4968 63484 5010 63524
rect 5050 63484 5092 63524
rect 5132 63484 5174 63524
rect 5214 63484 5256 63524
rect 5296 63484 20048 63524
rect 20088 63484 20130 63524
rect 20170 63484 20212 63524
rect 20252 63484 20294 63524
rect 20334 63484 20376 63524
rect 20416 63484 20452 63524
rect 1152 63460 20452 63484
rect 5547 63356 5589 63365
rect 5547 63316 5548 63356
rect 5588 63316 5589 63356
rect 5547 63307 5589 63316
rect 9178 63356 9236 63357
rect 9178 63316 9187 63356
rect 9227 63316 9236 63356
rect 9178 63315 9236 63316
rect 9483 63356 9525 63365
rect 9483 63316 9484 63356
rect 9524 63316 9525 63356
rect 9483 63307 9525 63316
rect 12411 63356 12453 63365
rect 12411 63316 12412 63356
rect 12452 63316 12453 63356
rect 12411 63307 12453 63316
rect 13563 63356 13605 63365
rect 13563 63316 13564 63356
rect 13604 63316 13605 63356
rect 13563 63307 13605 63316
rect 15531 63356 15573 63365
rect 15531 63316 15532 63356
rect 15572 63316 15573 63356
rect 15531 63307 15573 63316
rect 19851 63356 19893 63365
rect 19851 63316 19852 63356
rect 19892 63316 19893 63356
rect 19851 63307 19893 63316
rect 8427 63272 8469 63281
rect 8427 63232 8428 63272
rect 8468 63232 8469 63272
rect 8427 63223 8469 63232
rect 9867 63272 9909 63281
rect 9867 63232 9868 63272
rect 9908 63232 9909 63272
rect 9867 63223 9909 63232
rect 1707 63188 1749 63197
rect 3915 63188 3957 63197
rect 6987 63188 7029 63197
rect 1707 63148 1708 63188
rect 1748 63148 1749 63188
rect 1707 63139 1749 63148
rect 2955 63179 2997 63188
rect 2955 63139 2956 63179
rect 2996 63139 2997 63179
rect 3915 63148 3916 63188
rect 3956 63148 3957 63188
rect 3915 63139 3957 63148
rect 5163 63179 5205 63188
rect 5163 63139 5164 63179
rect 5204 63139 5205 63179
rect 2955 63130 2997 63139
rect 5163 63130 5205 63139
rect 5739 63179 5781 63188
rect 5739 63139 5740 63179
rect 5780 63139 5781 63179
rect 6987 63148 6988 63188
rect 7028 63148 7029 63188
rect 6987 63139 7029 63148
rect 8043 63188 8085 63197
rect 8043 63148 8044 63188
rect 8084 63148 8085 63188
rect 8043 63139 8085 63148
rect 8290 63188 8348 63189
rect 8290 63148 8299 63188
rect 8339 63148 8348 63188
rect 8290 63147 8348 63148
rect 8854 63188 8896 63197
rect 8854 63148 8855 63188
rect 8895 63148 8896 63188
rect 8854 63139 8896 63148
rect 9099 63188 9141 63197
rect 9099 63148 9100 63188
rect 9140 63148 9141 63188
rect 9099 63139 9141 63148
rect 9387 63188 9429 63197
rect 9387 63148 9388 63188
rect 9428 63148 9429 63188
rect 9387 63139 9429 63148
rect 9562 63188 9620 63189
rect 9562 63148 9571 63188
rect 9611 63148 9620 63188
rect 9562 63147 9620 63148
rect 9771 63188 9813 63197
rect 9771 63148 9772 63188
rect 9812 63148 9813 63188
rect 9771 63139 9813 63148
rect 9963 63188 10005 63197
rect 9963 63148 9964 63188
rect 10004 63148 10005 63188
rect 9963 63139 10005 63148
rect 10347 63188 10389 63197
rect 13786 63188 13844 63189
rect 10347 63148 10348 63188
rect 10388 63148 10389 63188
rect 10347 63139 10389 63148
rect 11595 63179 11637 63188
rect 11595 63139 11596 63179
rect 11636 63139 11637 63179
rect 13786 63148 13795 63188
rect 13835 63148 13844 63188
rect 13786 63147 13844 63148
rect 13899 63188 13941 63197
rect 13899 63148 13900 63188
rect 13940 63148 13941 63188
rect 13899 63139 13941 63148
rect 14283 63188 14325 63197
rect 17163 63188 17205 63197
rect 14283 63148 14284 63188
rect 14324 63148 14325 63188
rect 14283 63139 14325 63148
rect 14859 63179 14901 63188
rect 14859 63139 14860 63179
rect 14900 63139 14901 63179
rect 5739 63130 5781 63139
rect 11595 63130 11637 63139
rect 14859 63130 14901 63139
rect 15339 63179 15381 63188
rect 15339 63139 15340 63179
rect 15380 63139 15381 63179
rect 15339 63130 15381 63139
rect 15915 63179 15957 63188
rect 15915 63139 15916 63179
rect 15956 63139 15957 63179
rect 17163 63148 17164 63188
rect 17204 63148 17205 63188
rect 17163 63139 17205 63148
rect 18093 63188 18135 63197
rect 18093 63148 18094 63188
rect 18134 63148 18135 63188
rect 18093 63139 18135 63148
rect 18217 63188 18259 63197
rect 18217 63148 18218 63188
rect 18258 63148 18259 63188
rect 18217 63139 18259 63148
rect 18603 63188 18645 63197
rect 18603 63148 18604 63188
rect 18644 63148 18645 63188
rect 18603 63139 18645 63148
rect 19179 63179 19221 63188
rect 19179 63139 19180 63179
rect 19220 63139 19221 63179
rect 15915 63130 15957 63139
rect 19179 63130 19221 63139
rect 19659 63179 19701 63188
rect 19659 63139 19660 63179
rect 19700 63139 19701 63179
rect 19659 63130 19701 63139
rect 1419 63104 1461 63113
rect 1419 63064 1420 63104
rect 1460 63064 1461 63104
rect 1419 63055 1461 63064
rect 3531 63104 3573 63113
rect 3531 63064 3532 63104
rect 3572 63064 3573 63104
rect 3531 63055 3573 63064
rect 7371 63104 7413 63113
rect 7371 63064 7372 63104
rect 7412 63064 7413 63104
rect 7371 63055 7413 63064
rect 7755 63104 7797 63113
rect 7755 63064 7756 63104
rect 7796 63064 7797 63104
rect 7755 63055 7797 63064
rect 8986 63104 9044 63105
rect 8986 63064 8995 63104
rect 9035 63064 9044 63104
rect 8986 63063 9044 63064
rect 12171 63104 12213 63113
rect 12171 63064 12172 63104
rect 12212 63064 12213 63104
rect 12171 63055 12213 63064
rect 12939 63104 12981 63113
rect 12939 63064 12940 63104
rect 12980 63064 12981 63104
rect 12939 63055 12981 63064
rect 13323 63104 13365 63113
rect 13323 63064 13324 63104
rect 13364 63064 13365 63104
rect 13323 63055 13365 63064
rect 14379 63104 14421 63113
rect 14379 63064 14380 63104
rect 14420 63064 14421 63104
rect 14379 63055 14421 63064
rect 17643 63104 17685 63113
rect 17643 63064 17644 63104
rect 17684 63064 17685 63104
rect 17643 63055 17685 63064
rect 18699 63104 18741 63113
rect 18699 63064 18700 63104
rect 18740 63064 18741 63104
rect 18699 63055 18741 63064
rect 20139 63104 20181 63113
rect 20139 63064 20140 63104
rect 20180 63064 20181 63104
rect 20139 63055 20181 63064
rect 3291 63020 3333 63029
rect 3291 62980 3292 63020
rect 3332 62980 3333 63020
rect 3291 62971 3333 62980
rect 5355 63020 5397 63029
rect 5355 62980 5356 63020
rect 5396 62980 5397 63020
rect 5355 62971 5397 62980
rect 8715 63020 8757 63029
rect 8715 62980 8716 63020
rect 8756 62980 8757 63020
rect 8715 62971 8757 62980
rect 13179 63020 13221 63029
rect 13179 62980 13180 63020
rect 13220 62980 13221 63020
rect 13179 62971 13221 62980
rect 1179 62936 1221 62945
rect 1179 62896 1180 62936
rect 1220 62896 1221 62936
rect 1179 62887 1221 62896
rect 3147 62936 3189 62945
rect 3147 62896 3148 62936
rect 3188 62896 3189 62936
rect 3147 62887 3189 62896
rect 7131 62936 7173 62945
rect 7131 62896 7132 62936
rect 7172 62896 7173 62936
rect 7131 62887 7173 62896
rect 7515 62936 7557 62945
rect 7515 62896 7516 62936
rect 7556 62896 7557 62936
rect 7515 62887 7557 62896
rect 11787 62936 11829 62945
rect 11787 62896 11788 62936
rect 11828 62896 11829 62936
rect 11787 62887 11829 62896
rect 15723 62936 15765 62945
rect 15723 62896 15724 62936
rect 15764 62896 15765 62936
rect 15723 62887 15765 62896
rect 17883 62936 17925 62945
rect 17883 62896 17884 62936
rect 17924 62896 17925 62936
rect 17883 62887 17925 62896
rect 20379 62936 20421 62945
rect 20379 62896 20380 62936
rect 20420 62896 20421 62936
rect 20379 62887 20421 62896
rect 1152 62768 20448 62792
rect 1152 62728 3688 62768
rect 3728 62728 3770 62768
rect 3810 62728 3852 62768
rect 3892 62728 3934 62768
rect 3974 62728 4016 62768
rect 4056 62728 18808 62768
rect 18848 62728 18890 62768
rect 18930 62728 18972 62768
rect 19012 62728 19054 62768
rect 19094 62728 19136 62768
rect 19176 62728 20448 62768
rect 1152 62704 20448 62728
rect 9514 62600 9572 62601
rect 9514 62560 9523 62600
rect 9563 62560 9572 62600
rect 9514 62559 9572 62560
rect 13515 62600 13557 62609
rect 13515 62560 13516 62600
rect 13556 62560 13557 62600
rect 13515 62551 13557 62560
rect 14331 62600 14373 62609
rect 14331 62560 14332 62600
rect 14372 62560 14373 62600
rect 14331 62551 14373 62560
rect 19851 62600 19893 62609
rect 19851 62560 19852 62600
rect 19892 62560 19893 62600
rect 19851 62551 19893 62560
rect 3051 62432 3093 62441
rect 3051 62392 3052 62432
rect 3092 62392 3093 62432
rect 3051 62383 3093 62392
rect 3915 62432 3957 62441
rect 3915 62392 3916 62432
rect 3956 62392 3957 62432
rect 3915 62383 3957 62392
rect 6219 62432 6261 62441
rect 6219 62392 6220 62432
rect 6260 62392 6261 62432
rect 6219 62383 6261 62392
rect 8235 62432 8277 62441
rect 8235 62392 8236 62432
rect 8276 62392 8277 62432
rect 8235 62383 8277 62392
rect 10443 62432 10485 62441
rect 10443 62392 10444 62432
rect 10484 62392 10485 62432
rect 10443 62383 10485 62392
rect 13707 62432 13749 62441
rect 13707 62392 13708 62432
rect 13748 62392 13749 62432
rect 13707 62383 13749 62392
rect 14091 62432 14133 62441
rect 14091 62392 14092 62432
rect 14132 62392 14133 62432
rect 14091 62383 14133 62392
rect 15243 62432 15285 62441
rect 15243 62392 15244 62432
rect 15284 62392 15285 62432
rect 15243 62383 15285 62392
rect 20139 62432 20181 62441
rect 20139 62392 20140 62432
rect 20180 62392 20181 62432
rect 20139 62383 20181 62392
rect 1227 62348 1269 62357
rect 1227 62308 1228 62348
rect 1268 62308 1269 62348
rect 1227 62299 1269 62308
rect 2467 62348 2525 62349
rect 2467 62308 2476 62348
rect 2516 62308 2525 62348
rect 2467 62307 2525 62308
rect 3418 62348 3476 62349
rect 3418 62308 3427 62348
rect 3467 62308 3476 62348
rect 3418 62307 3476 62308
rect 3531 62348 3573 62357
rect 3531 62308 3532 62348
rect 3572 62308 3573 62348
rect 3531 62299 3573 62308
rect 4011 62348 4053 62357
rect 4011 62308 4012 62348
rect 4052 62308 4053 62348
rect 4011 62299 4053 62308
rect 4483 62348 4541 62349
rect 4483 62308 4492 62348
rect 4532 62308 4541 62348
rect 4483 62307 4541 62308
rect 5002 62348 5060 62349
rect 5002 62308 5011 62348
rect 5051 62308 5060 62348
rect 5002 62307 5060 62308
rect 5718 62348 5776 62349
rect 5718 62308 5727 62348
rect 5767 62308 5776 62348
rect 5718 62307 5776 62308
rect 5835 62348 5877 62357
rect 5835 62308 5836 62348
rect 5876 62308 5877 62348
rect 5835 62299 5877 62308
rect 6315 62348 6357 62357
rect 6315 62308 6316 62348
rect 6356 62308 6357 62348
rect 6315 62299 6357 62308
rect 6787 62348 6845 62349
rect 6787 62308 6796 62348
rect 6836 62308 6845 62348
rect 6787 62307 6845 62308
rect 7306 62348 7364 62349
rect 7306 62308 7315 62348
rect 7355 62308 7364 62348
rect 7306 62307 7364 62308
rect 7738 62348 7796 62349
rect 7738 62308 7747 62348
rect 7787 62308 7796 62348
rect 7738 62307 7796 62308
rect 7851 62348 7893 62357
rect 7851 62308 7852 62348
rect 7892 62308 7893 62348
rect 7851 62299 7893 62308
rect 8331 62348 8373 62357
rect 8331 62308 8332 62348
rect 8372 62308 8373 62348
rect 8331 62299 8373 62308
rect 8803 62348 8861 62349
rect 8803 62308 8812 62348
rect 8852 62308 8861 62348
rect 8803 62307 8861 62308
rect 9322 62348 9380 62349
rect 9322 62308 9331 62348
rect 9371 62308 9380 62348
rect 9322 62307 9380 62308
rect 9946 62348 10004 62349
rect 9946 62308 9955 62348
rect 9995 62308 10004 62348
rect 9946 62307 10004 62308
rect 10059 62348 10101 62357
rect 10059 62308 10060 62348
rect 10100 62308 10101 62348
rect 10059 62299 10101 62308
rect 10539 62348 10581 62357
rect 10539 62308 10540 62348
rect 10580 62308 10581 62348
rect 10539 62299 10581 62308
rect 11011 62348 11069 62349
rect 11011 62308 11020 62348
rect 11060 62308 11069 62348
rect 11011 62307 11069 62308
rect 11530 62348 11588 62349
rect 11530 62308 11539 62348
rect 11579 62308 11588 62348
rect 11530 62307 11588 62308
rect 12075 62348 12117 62357
rect 12075 62308 12076 62348
rect 12116 62308 12117 62348
rect 12075 62299 12117 62308
rect 13315 62348 13373 62349
rect 13315 62308 13324 62348
rect 13364 62308 13373 62348
rect 13315 62307 13373 62308
rect 14746 62348 14804 62349
rect 14746 62308 14755 62348
rect 14795 62308 14804 62348
rect 14746 62307 14804 62308
rect 14859 62348 14901 62357
rect 14859 62308 14860 62348
rect 14900 62308 14901 62348
rect 14859 62299 14901 62308
rect 15339 62348 15381 62357
rect 15339 62308 15340 62348
rect 15380 62308 15381 62348
rect 15339 62299 15381 62308
rect 15811 62348 15869 62349
rect 15811 62308 15820 62348
rect 15860 62308 15869 62348
rect 15811 62307 15869 62308
rect 16299 62348 16357 62349
rect 16299 62308 16308 62348
rect 16348 62308 16357 62348
rect 16299 62307 16357 62308
rect 16683 62348 16725 62357
rect 16683 62308 16684 62348
rect 16724 62308 16725 62348
rect 16683 62299 16725 62308
rect 17923 62348 17981 62349
rect 17923 62308 17932 62348
rect 17972 62308 17981 62348
rect 17923 62307 17981 62308
rect 18411 62348 18453 62357
rect 18411 62308 18412 62348
rect 18452 62308 18453 62348
rect 18411 62299 18453 62308
rect 19651 62348 19709 62349
rect 19651 62308 19660 62348
rect 19700 62308 19709 62348
rect 19651 62307 19709 62308
rect 13947 62264 13989 62273
rect 13947 62224 13948 62264
rect 13988 62224 13989 62264
rect 13947 62215 13989 62224
rect 2667 62180 2709 62189
rect 2667 62140 2668 62180
rect 2708 62140 2709 62180
rect 2667 62131 2709 62140
rect 2811 62180 2853 62189
rect 2811 62140 2812 62180
rect 2852 62140 2853 62180
rect 2811 62131 2853 62140
rect 5163 62180 5205 62189
rect 5163 62140 5164 62180
rect 5204 62140 5205 62180
rect 5163 62131 5205 62140
rect 7467 62180 7509 62189
rect 7467 62140 7468 62180
rect 7508 62140 7509 62180
rect 7467 62131 7509 62140
rect 11691 62180 11733 62189
rect 11691 62140 11692 62180
rect 11732 62140 11733 62180
rect 11691 62131 11733 62140
rect 16491 62180 16533 62189
rect 16491 62140 16492 62180
rect 16532 62140 16533 62180
rect 16491 62131 16533 62140
rect 18123 62180 18165 62189
rect 18123 62140 18124 62180
rect 18164 62140 18165 62180
rect 18123 62131 18165 62140
rect 20379 62180 20421 62189
rect 20379 62140 20380 62180
rect 20420 62140 20421 62180
rect 20379 62131 20421 62140
rect 1152 62012 20452 62036
rect 1152 61972 4928 62012
rect 4968 61972 5010 62012
rect 5050 61972 5092 62012
rect 5132 61972 5174 62012
rect 5214 61972 5256 62012
rect 5296 61972 20048 62012
rect 20088 61972 20130 62012
rect 20170 61972 20212 62012
rect 20252 61972 20294 62012
rect 20334 61972 20376 62012
rect 20416 61972 20452 62012
rect 1152 61948 20452 61972
rect 5307 61844 5349 61853
rect 5307 61804 5308 61844
rect 5348 61804 5349 61844
rect 5307 61795 5349 61804
rect 7371 61844 7413 61853
rect 7371 61804 7372 61844
rect 7412 61804 7413 61844
rect 7371 61795 7413 61804
rect 11403 61844 11445 61853
rect 11403 61804 11404 61844
rect 11444 61804 11445 61844
rect 11403 61795 11445 61804
rect 11739 61844 11781 61853
rect 11739 61804 11740 61844
rect 11780 61804 11781 61844
rect 11739 61795 11781 61804
rect 13611 61844 13653 61853
rect 13611 61804 13612 61844
rect 13652 61804 13653 61844
rect 13611 61795 13653 61804
rect 15243 61844 15285 61853
rect 15243 61804 15244 61844
rect 15284 61804 15285 61844
rect 15243 61795 15285 61804
rect 18123 61844 18165 61853
rect 18123 61804 18124 61844
rect 18164 61804 18165 61844
rect 18123 61795 18165 61804
rect 20139 61844 20181 61853
rect 20139 61804 20140 61844
rect 20180 61804 20181 61844
rect 20139 61795 20181 61804
rect 7515 61760 7557 61769
rect 7515 61720 7516 61760
rect 7556 61720 7557 61760
rect 7515 61711 7557 61720
rect 9387 61760 9429 61769
rect 9387 61720 9388 61760
rect 9428 61720 9429 61760
rect 9387 61711 9429 61720
rect 1707 61676 1749 61685
rect 3405 61676 3447 61685
rect 1707 61636 1708 61676
rect 1748 61636 1749 61676
rect 1707 61627 1749 61636
rect 2955 61667 2997 61676
rect 2955 61627 2956 61667
rect 2996 61627 2997 61667
rect 3405 61636 3406 61676
rect 3446 61636 3447 61676
rect 3405 61627 3447 61636
rect 3531 61676 3573 61685
rect 3531 61636 3532 61676
rect 3572 61636 3573 61676
rect 3531 61627 3573 61636
rect 3915 61676 3957 61685
rect 5931 61676 5973 61685
rect 7947 61676 7989 61685
rect 9658 61676 9716 61677
rect 3915 61636 3916 61676
rect 3956 61636 3957 61676
rect 3915 61627 3957 61636
rect 4491 61667 4533 61676
rect 4491 61627 4492 61667
rect 4532 61627 4533 61667
rect 2955 61618 2997 61627
rect 4491 61618 4533 61627
rect 4971 61667 5013 61676
rect 4971 61627 4972 61667
rect 5012 61627 5013 61667
rect 5931 61636 5932 61676
rect 5972 61636 5973 61676
rect 5931 61627 5973 61636
rect 7179 61667 7221 61676
rect 7179 61627 7180 61667
rect 7220 61627 7221 61667
rect 7947 61636 7948 61676
rect 7988 61636 7989 61676
rect 7947 61627 7989 61636
rect 9195 61667 9237 61676
rect 9195 61627 9196 61667
rect 9236 61627 9237 61667
rect 9658 61636 9667 61676
rect 9707 61636 9716 61676
rect 9658 61635 9716 61636
rect 9771 61676 9813 61685
rect 9771 61636 9772 61676
rect 9812 61636 9813 61676
rect 9771 61627 9813 61636
rect 10155 61676 10197 61685
rect 12171 61676 12213 61685
rect 13803 61676 13845 61685
rect 16378 61676 16436 61677
rect 10155 61636 10156 61676
rect 10196 61636 10197 61676
rect 10155 61627 10197 61636
rect 10731 61667 10773 61676
rect 10731 61627 10732 61667
rect 10772 61627 10773 61667
rect 4971 61618 5013 61627
rect 7179 61618 7221 61627
rect 9195 61618 9237 61627
rect 10731 61618 10773 61627
rect 11211 61667 11253 61676
rect 11211 61627 11212 61667
rect 11252 61627 11253 61667
rect 12171 61636 12172 61676
rect 12212 61636 12213 61676
rect 12171 61627 12213 61636
rect 13419 61667 13461 61676
rect 13419 61627 13420 61667
rect 13460 61627 13461 61667
rect 13803 61636 13804 61676
rect 13844 61636 13845 61676
rect 13803 61627 13845 61636
rect 15051 61667 15093 61676
rect 15051 61627 15052 61667
rect 15092 61627 15093 61667
rect 16378 61636 16387 61676
rect 16427 61636 16436 61676
rect 16378 61635 16436 61636
rect 16491 61676 16533 61685
rect 16491 61636 16492 61676
rect 16532 61636 16533 61676
rect 16491 61627 16533 61636
rect 16875 61676 16917 61685
rect 18394 61676 18452 61677
rect 16875 61636 16876 61676
rect 16916 61636 16917 61676
rect 16875 61627 16917 61636
rect 17451 61667 17493 61676
rect 17451 61627 17452 61667
rect 17492 61627 17493 61667
rect 11211 61618 11253 61627
rect 13419 61618 13461 61627
rect 15051 61618 15093 61627
rect 17451 61618 17493 61627
rect 17931 61667 17973 61676
rect 17931 61627 17932 61667
rect 17972 61627 17973 61667
rect 18394 61636 18403 61676
rect 18443 61636 18452 61676
rect 18394 61635 18452 61636
rect 18507 61676 18549 61685
rect 18507 61636 18508 61676
rect 18548 61636 18549 61676
rect 18507 61627 18549 61636
rect 18891 61676 18933 61685
rect 18891 61636 18892 61676
rect 18932 61636 18933 61676
rect 18891 61627 18933 61636
rect 19467 61667 19509 61676
rect 19467 61627 19468 61667
rect 19508 61627 19509 61667
rect 17931 61618 17973 61627
rect 19467 61618 19509 61627
rect 19947 61667 19989 61676
rect 19947 61627 19948 61667
rect 19988 61627 19989 61667
rect 19947 61618 19989 61627
rect 1419 61592 1461 61601
rect 1419 61552 1420 61592
rect 1460 61552 1461 61592
rect 1419 61543 1461 61552
rect 4011 61592 4053 61601
rect 4011 61552 4012 61592
rect 4052 61552 4053 61592
rect 4011 61543 4053 61552
rect 5547 61592 5589 61601
rect 5547 61552 5548 61592
rect 5588 61552 5589 61592
rect 5547 61543 5589 61552
rect 7755 61592 7797 61601
rect 7755 61552 7756 61592
rect 7796 61552 7797 61592
rect 7755 61543 7797 61552
rect 10251 61592 10293 61601
rect 10251 61552 10252 61592
rect 10292 61552 10293 61592
rect 10251 61543 10293 61552
rect 11979 61592 12021 61601
rect 11979 61552 11980 61592
rect 12020 61552 12021 61592
rect 11979 61543 12021 61552
rect 15723 61592 15765 61601
rect 15723 61552 15724 61592
rect 15764 61552 15765 61592
rect 15723 61543 15765 61552
rect 16107 61592 16149 61601
rect 16107 61552 16108 61592
rect 16148 61552 16149 61592
rect 16107 61543 16149 61552
rect 16971 61592 17013 61601
rect 16971 61552 16972 61592
rect 17012 61552 17013 61592
rect 16971 61543 17013 61552
rect 18987 61592 19029 61601
rect 18987 61552 18988 61592
rect 19028 61552 19029 61592
rect 18987 61543 19029 61552
rect 15867 61508 15909 61517
rect 15867 61468 15868 61508
rect 15908 61468 15909 61508
rect 15867 61459 15909 61468
rect 1179 61424 1221 61433
rect 1179 61384 1180 61424
rect 1220 61384 1221 61424
rect 1179 61375 1221 61384
rect 3147 61424 3189 61433
rect 3147 61384 3148 61424
rect 3188 61384 3189 61424
rect 3147 61375 3189 61384
rect 5194 61424 5252 61425
rect 5194 61384 5203 61424
rect 5243 61384 5252 61424
rect 5194 61383 5252 61384
rect 15483 61424 15525 61433
rect 15483 61384 15484 61424
rect 15524 61384 15525 61424
rect 15483 61375 15525 61384
rect 1152 61256 20448 61280
rect 1152 61216 3688 61256
rect 3728 61216 3770 61256
rect 3810 61216 3852 61256
rect 3892 61216 3934 61256
rect 3974 61216 4016 61256
rect 4056 61216 18808 61256
rect 18848 61216 18890 61256
rect 18930 61216 18972 61256
rect 19012 61216 19054 61256
rect 19094 61216 19136 61256
rect 19176 61216 20448 61256
rect 1152 61192 20448 61216
rect 11499 61088 11541 61097
rect 11499 61048 11500 61088
rect 11540 61048 11541 61088
rect 11499 61039 11541 61048
rect 14139 61088 14181 61097
rect 14139 61048 14140 61088
rect 14180 61048 14181 61088
rect 14139 61039 14181 61048
rect 16491 61088 16533 61097
rect 16491 61048 16492 61088
rect 16532 61048 16533 61088
rect 16491 61039 16533 61048
rect 18123 61088 18165 61097
rect 18123 61048 18124 61088
rect 18164 61048 18165 61088
rect 18123 61039 18165 61048
rect 20043 61088 20085 61097
rect 20043 61048 20044 61088
rect 20084 61048 20085 61088
rect 20043 61039 20085 61048
rect 5499 61004 5541 61013
rect 5499 60964 5500 61004
rect 5540 60964 5541 61004
rect 5499 60955 5541 60964
rect 12555 61004 12597 61013
rect 12555 60964 12556 61004
rect 12596 60964 12597 61004
rect 12555 60955 12597 60964
rect 3051 60920 3093 60929
rect 3051 60880 3052 60920
rect 3092 60880 3093 60920
rect 3051 60871 3093 60880
rect 4107 60920 4149 60929
rect 4107 60880 4108 60920
rect 4148 60880 4149 60920
rect 4107 60871 4149 60880
rect 5386 60920 5444 60921
rect 5386 60880 5395 60920
rect 5435 60880 5444 60920
rect 5386 60879 5444 60880
rect 5739 60920 5781 60929
rect 5739 60880 5740 60920
rect 5780 60880 5781 60920
rect 5739 60871 5781 60880
rect 6123 60920 6165 60929
rect 6123 60880 6124 60920
rect 6164 60880 6165 60920
rect 6123 60871 6165 60880
rect 8523 60920 8565 60929
rect 8523 60880 8524 60920
rect 8564 60880 8565 60920
rect 8523 60871 8565 60880
rect 12171 60920 12213 60929
rect 12171 60880 12172 60920
rect 12212 60880 12213 60920
rect 12171 60871 12213 60880
rect 14379 60920 14421 60929
rect 14379 60880 14380 60920
rect 14420 60880 14421 60920
rect 14379 60871 14421 60880
rect 14667 60920 14709 60929
rect 14667 60880 14668 60920
rect 14708 60880 14709 60920
rect 14667 60871 14709 60880
rect 1227 60836 1269 60845
rect 1227 60796 1228 60836
rect 1268 60796 1269 60836
rect 1227 60787 1269 60796
rect 2467 60836 2525 60837
rect 2467 60796 2476 60836
rect 2516 60796 2525 60836
rect 2467 60795 2525 60796
rect 3610 60836 3668 60837
rect 3610 60796 3619 60836
rect 3659 60796 3668 60836
rect 3610 60795 3668 60796
rect 3723 60836 3765 60845
rect 3723 60796 3724 60836
rect 3764 60796 3765 60836
rect 3723 60787 3765 60796
rect 4203 60836 4245 60845
rect 4203 60796 4204 60836
rect 4244 60796 4245 60836
rect 4203 60787 4245 60796
rect 4675 60836 4733 60837
rect 4675 60796 4684 60836
rect 4724 60796 4733 60836
rect 4675 60795 4733 60796
rect 5194 60836 5252 60837
rect 5194 60796 5203 60836
rect 5243 60796 5252 60836
rect 5194 60795 5252 60796
rect 6315 60836 6357 60845
rect 6315 60796 6316 60836
rect 6356 60796 6357 60836
rect 6315 60787 6357 60796
rect 7555 60836 7613 60837
rect 7555 60796 7564 60836
rect 7604 60796 7613 60836
rect 7555 60795 7613 60796
rect 8026 60836 8084 60837
rect 8026 60796 8035 60836
rect 8075 60796 8084 60836
rect 8026 60795 8084 60796
rect 8139 60836 8181 60845
rect 8139 60796 8140 60836
rect 8180 60796 8181 60836
rect 8139 60787 8181 60796
rect 8619 60836 8661 60845
rect 8619 60796 8620 60836
rect 8660 60796 8661 60836
rect 8619 60787 8661 60796
rect 9091 60836 9149 60837
rect 9091 60796 9100 60836
rect 9140 60796 9149 60836
rect 9091 60795 9149 60796
rect 9610 60836 9668 60837
rect 9610 60796 9619 60836
rect 9659 60796 9668 60836
rect 9610 60795 9668 60796
rect 10059 60836 10101 60845
rect 10059 60796 10060 60836
rect 10100 60796 10101 60836
rect 10059 60787 10101 60796
rect 11299 60836 11357 60837
rect 11299 60796 11308 60836
rect 11348 60796 11357 60836
rect 11299 60795 11357 60796
rect 12739 60836 12797 60837
rect 12739 60796 12748 60836
rect 12788 60796 12797 60836
rect 12739 60795 12797 60796
rect 13995 60836 14037 60845
rect 13995 60796 13996 60836
rect 14036 60796 14037 60836
rect 13995 60787 14037 60796
rect 15051 60836 15093 60845
rect 15051 60796 15052 60836
rect 15092 60796 15093 60836
rect 15051 60787 15093 60796
rect 16291 60836 16349 60837
rect 16291 60796 16300 60836
rect 16340 60796 16349 60836
rect 16291 60795 16349 60796
rect 16683 60836 16725 60845
rect 16683 60796 16684 60836
rect 16724 60796 16725 60836
rect 16683 60787 16725 60796
rect 17923 60836 17981 60837
rect 17923 60796 17932 60836
rect 17972 60796 17981 60836
rect 17923 60795 17981 60796
rect 18603 60836 18645 60845
rect 18603 60796 18604 60836
rect 18644 60796 18645 60836
rect 18603 60787 18645 60796
rect 19843 60836 19901 60837
rect 19843 60796 19852 60836
rect 19892 60796 19901 60836
rect 19843 60795 19901 60796
rect 7755 60752 7797 60761
rect 7755 60712 7756 60752
rect 7796 60712 7797 60752
rect 7755 60703 7797 60712
rect 2667 60668 2709 60677
rect 2667 60628 2668 60668
rect 2708 60628 2709 60668
rect 2667 60619 2709 60628
rect 2811 60668 2853 60677
rect 2811 60628 2812 60668
rect 2852 60628 2853 60668
rect 2811 60619 2853 60628
rect 5883 60668 5925 60677
rect 5883 60628 5884 60668
rect 5924 60628 5925 60668
rect 5883 60619 5925 60628
rect 9771 60668 9813 60677
rect 9771 60628 9772 60668
rect 9812 60628 9813 60668
rect 9771 60619 9813 60628
rect 12411 60668 12453 60677
rect 12411 60628 12412 60668
rect 12452 60628 12453 60668
rect 12411 60619 12453 60628
rect 14907 60668 14949 60677
rect 14907 60628 14908 60668
rect 14948 60628 14949 60668
rect 14907 60619 14949 60628
rect 1152 60500 20452 60524
rect 1152 60460 4928 60500
rect 4968 60460 5010 60500
rect 5050 60460 5092 60500
rect 5132 60460 5174 60500
rect 5214 60460 5256 60500
rect 5296 60460 20048 60500
rect 20088 60460 20130 60500
rect 20170 60460 20212 60500
rect 20252 60460 20294 60500
rect 20334 60460 20376 60500
rect 20416 60460 20452 60500
rect 1152 60436 20452 60460
rect 5547 60332 5589 60341
rect 5547 60292 5548 60332
rect 5588 60292 5589 60332
rect 5547 60283 5589 60292
rect 7899 60332 7941 60341
rect 7899 60292 7900 60332
rect 7940 60292 7941 60332
rect 7899 60283 7941 60292
rect 12603 60332 12645 60341
rect 12603 60292 12604 60332
rect 12644 60292 12645 60332
rect 12603 60283 12645 60292
rect 14139 60332 14181 60341
rect 14139 60292 14140 60332
rect 14180 60292 14181 60332
rect 14139 60283 14181 60292
rect 14907 60332 14949 60341
rect 14907 60292 14908 60332
rect 14948 60292 14949 60332
rect 14907 60283 14949 60292
rect 15435 60332 15477 60341
rect 15435 60292 15436 60332
rect 15476 60292 15477 60332
rect 15435 60283 15477 60292
rect 16011 60248 16053 60257
rect 16011 60208 16012 60248
rect 16052 60208 16053 60248
rect 16011 60199 16053 60208
rect 17163 60248 17205 60257
rect 17163 60208 17164 60248
rect 17204 60208 17205 60248
rect 17163 60199 17205 60208
rect 2170 60164 2228 60165
rect 2170 60124 2179 60164
rect 2219 60124 2228 60164
rect 2170 60123 2228 60124
rect 2283 60164 2325 60173
rect 2283 60124 2284 60164
rect 2324 60124 2325 60164
rect 2283 60115 2325 60124
rect 2667 60164 2709 60173
rect 4107 60164 4149 60173
rect 5835 60164 5877 60173
rect 9099 60164 9141 60173
rect 10731 60164 10773 60173
rect 15531 60164 15573 60173
rect 2667 60124 2668 60164
rect 2708 60124 2709 60164
rect 2667 60115 2709 60124
rect 3243 60155 3285 60164
rect 3243 60115 3244 60155
rect 3284 60115 3285 60155
rect 3243 60106 3285 60115
rect 3723 60155 3765 60164
rect 3723 60115 3724 60155
rect 3764 60115 3765 60155
rect 4107 60124 4108 60164
rect 4148 60124 4149 60164
rect 4107 60115 4149 60124
rect 5355 60155 5397 60164
rect 5355 60115 5356 60155
rect 5396 60115 5397 60155
rect 5835 60124 5836 60164
rect 5876 60124 5877 60164
rect 5835 60115 5877 60124
rect 7083 60155 7125 60164
rect 7083 60115 7084 60155
rect 7124 60115 7125 60155
rect 9099 60124 9100 60164
rect 9140 60124 9141 60164
rect 9099 60115 9141 60124
rect 10347 60155 10389 60164
rect 10347 60115 10348 60155
rect 10388 60115 10389 60155
rect 10731 60124 10732 60164
rect 10772 60124 10773 60164
rect 10731 60115 10773 60124
rect 11979 60155 12021 60164
rect 11979 60115 11980 60155
rect 12020 60115 12021 60155
rect 15531 60124 15532 60164
rect 15572 60124 15573 60164
rect 15531 60115 15573 60124
rect 15760 60164 15818 60165
rect 15760 60124 15769 60164
rect 15809 60124 15818 60164
rect 15760 60123 15818 60124
rect 15914 60164 15956 60173
rect 15914 60124 15915 60164
rect 15955 60124 15956 60164
rect 15914 60115 15956 60124
rect 16206 60164 16248 60173
rect 16206 60124 16207 60164
rect 16247 60124 16248 60164
rect 16206 60115 16248 60124
rect 16395 60164 16437 60173
rect 16395 60124 16396 60164
rect 16436 60124 16437 60164
rect 16395 60115 16437 60124
rect 16779 60164 16821 60173
rect 16779 60124 16780 60164
rect 16820 60124 16821 60164
rect 16779 60115 16821 60124
rect 17050 60164 17108 60165
rect 17050 60124 17059 60164
rect 17099 60124 17108 60164
rect 17050 60123 17108 60124
rect 17643 60164 17685 60173
rect 17643 60124 17644 60164
rect 17684 60124 17685 60164
rect 17643 60115 17685 60124
rect 17818 60164 17876 60165
rect 17818 60124 17827 60164
rect 17867 60124 17876 60164
rect 17818 60123 17876 60124
rect 18699 60164 18741 60173
rect 18699 60124 18700 60164
rect 18740 60124 18741 60164
rect 18699 60115 18741 60124
rect 19947 60155 19989 60164
rect 19947 60115 19948 60155
rect 19988 60115 19989 60155
rect 3723 60106 3765 60115
rect 5355 60106 5397 60115
rect 7083 60106 7125 60115
rect 10347 60106 10389 60115
rect 11979 60106 12021 60115
rect 19947 60106 19989 60115
rect 1179 60080 1221 60089
rect 1179 60040 1180 60080
rect 1220 60040 1221 60080
rect 1179 60031 1221 60040
rect 1419 60080 1461 60089
rect 1419 60040 1420 60080
rect 1460 60040 1461 60080
rect 1419 60031 1461 60040
rect 1803 60080 1845 60089
rect 1803 60040 1804 60080
rect 1844 60040 1845 60080
rect 1803 60031 1845 60040
rect 2763 60080 2805 60089
rect 2763 60040 2764 60080
rect 2804 60040 2805 60080
rect 2763 60031 2805 60040
rect 7659 60080 7701 60089
rect 7659 60040 7660 60080
rect 7700 60040 7701 60080
rect 7659 60031 7701 60040
rect 12363 60080 12405 60089
rect 12363 60040 12364 60080
rect 12404 60040 12405 60080
rect 12363 60031 12405 60040
rect 13035 60080 13077 60089
rect 13035 60040 13036 60080
rect 13076 60040 13077 60080
rect 13035 60031 13077 60040
rect 13419 60080 13461 60089
rect 13419 60040 13420 60080
rect 13460 60040 13461 60080
rect 13419 60031 13461 60040
rect 14379 60080 14421 60089
rect 14379 60040 14380 60080
rect 14420 60040 14421 60080
rect 14379 60031 14421 60040
rect 14667 60080 14709 60089
rect 14667 60040 14668 60080
rect 14708 60040 14709 60080
rect 14667 60031 14709 60040
rect 15051 60080 15093 60089
rect 18315 60080 18357 60089
rect 15051 60040 15052 60080
rect 15092 60040 15093 60080
rect 15051 60031 15093 60040
rect 15666 60071 15712 60080
rect 15666 60031 15667 60071
rect 15707 60031 15712 60071
rect 18315 60040 18316 60080
rect 18356 60040 18357 60080
rect 18315 60031 18357 60040
rect 15666 60022 15712 60031
rect 12795 59996 12837 60005
rect 12795 59956 12796 59996
rect 12836 59956 12837 59996
rect 12795 59947 12837 59956
rect 13995 59996 14037 60005
rect 13995 59956 13996 59996
rect 14036 59956 14037 59996
rect 13995 59947 14037 59956
rect 16539 59996 16581 60005
rect 16539 59956 16540 59996
rect 16580 59956 16581 59996
rect 16539 59947 16581 59956
rect 1563 59912 1605 59921
rect 1563 59872 1564 59912
rect 1604 59872 1605 59912
rect 1563 59863 1605 59872
rect 3946 59912 4004 59913
rect 3946 59872 3955 59912
rect 3995 59872 4004 59912
rect 3946 59871 4004 59872
rect 7275 59912 7317 59921
rect 7275 59872 7276 59912
rect 7316 59872 7317 59912
rect 7275 59863 7317 59872
rect 10539 59912 10581 59921
rect 10539 59872 10540 59912
rect 10580 59872 10581 59912
rect 10539 59863 10581 59872
rect 12171 59912 12213 59921
rect 12171 59872 12172 59912
rect 12212 59872 12213 59912
rect 12171 59863 12213 59872
rect 13179 59912 13221 59921
rect 13179 59872 13180 59912
rect 13220 59872 13221 59912
rect 13179 59863 13221 59872
rect 15291 59912 15333 59921
rect 15291 59872 15292 59912
rect 15332 59872 15333 59912
rect 15291 59863 15333 59872
rect 17451 59912 17493 59921
rect 17451 59872 17452 59912
rect 17492 59872 17493 59912
rect 17451 59863 17493 59872
rect 17818 59912 17876 59913
rect 17818 59872 17827 59912
rect 17867 59872 17876 59912
rect 17818 59871 17876 59872
rect 18555 59912 18597 59921
rect 18555 59872 18556 59912
rect 18596 59872 18597 59912
rect 18555 59863 18597 59872
rect 20139 59912 20181 59921
rect 20139 59872 20140 59912
rect 20180 59872 20181 59912
rect 20139 59863 20181 59872
rect 1152 59744 20448 59768
rect 1152 59704 3688 59744
rect 3728 59704 3770 59744
rect 3810 59704 3852 59744
rect 3892 59704 3934 59744
rect 3974 59704 4016 59744
rect 4056 59704 18808 59744
rect 18848 59704 18890 59744
rect 18930 59704 18972 59744
rect 19012 59704 19054 59744
rect 19094 59704 19136 59744
rect 19176 59704 20448 59744
rect 1152 59680 20448 59704
rect 3675 59576 3717 59585
rect 3675 59536 3676 59576
rect 3716 59536 3717 59576
rect 3675 59527 3717 59536
rect 7803 59576 7845 59585
rect 7803 59536 7804 59576
rect 7844 59536 7845 59576
rect 7803 59527 7845 59536
rect 8187 59576 8229 59585
rect 8187 59536 8188 59576
rect 8228 59536 8229 59576
rect 8187 59527 8229 59536
rect 14667 59576 14709 59585
rect 14667 59536 14668 59576
rect 14708 59536 14709 59576
rect 14667 59527 14709 59536
rect 16299 59492 16341 59501
rect 16299 59452 16300 59492
rect 16340 59452 16341 59492
rect 16299 59443 16341 59452
rect 1419 59408 1461 59417
rect 1419 59368 1420 59408
rect 1460 59368 1461 59408
rect 1419 59359 1461 59368
rect 3531 59408 3573 59417
rect 3531 59368 3532 59408
rect 3572 59368 3573 59408
rect 3531 59359 3573 59368
rect 3915 59408 3957 59417
rect 3915 59368 3916 59408
rect 3956 59368 3957 59408
rect 3915 59359 3957 59368
rect 6315 59408 6357 59417
rect 6315 59368 6316 59408
rect 6356 59368 6357 59408
rect 6315 59359 6357 59368
rect 8043 59408 8085 59417
rect 8043 59368 8044 59408
rect 8084 59368 8085 59408
rect 8043 59359 8085 59368
rect 8427 59408 8469 59417
rect 8427 59368 8428 59408
rect 8468 59368 8469 59408
rect 8427 59359 8469 59368
rect 11211 59408 11253 59417
rect 11211 59368 11212 59408
rect 11252 59368 11253 59408
rect 11211 59359 11253 59368
rect 12490 59408 12548 59409
rect 12490 59368 12499 59408
rect 12539 59368 12548 59408
rect 12490 59367 12548 59368
rect 12843 59408 12885 59417
rect 12843 59368 12844 59408
rect 12884 59368 12885 59408
rect 12843 59359 12885 59368
rect 18891 59408 18933 59417
rect 18891 59368 18892 59408
rect 18932 59368 18933 59408
rect 18891 59359 18933 59368
rect 1611 59324 1653 59333
rect 1611 59284 1612 59324
rect 1652 59284 1653 59324
rect 1611 59275 1653 59284
rect 2851 59324 2909 59325
rect 2851 59284 2860 59324
rect 2900 59284 2909 59324
rect 2851 59283 2909 59284
rect 4107 59324 4149 59333
rect 4107 59284 4108 59324
rect 4148 59284 4149 59324
rect 4107 59275 4149 59284
rect 5347 59324 5405 59325
rect 5347 59284 5356 59324
rect 5396 59284 5405 59324
rect 5347 59283 5405 59284
rect 5818 59324 5876 59325
rect 5818 59284 5827 59324
rect 5867 59284 5876 59324
rect 5818 59283 5876 59284
rect 5931 59324 5973 59333
rect 5931 59284 5932 59324
rect 5972 59284 5973 59324
rect 5931 59275 5973 59284
rect 6411 59324 6453 59333
rect 6411 59284 6412 59324
rect 6452 59284 6453 59324
rect 6411 59275 6453 59284
rect 6883 59324 6941 59325
rect 6883 59284 6892 59324
rect 6932 59284 6941 59324
rect 6883 59283 6941 59284
rect 7371 59324 7429 59325
rect 7371 59284 7380 59324
rect 7420 59284 7429 59324
rect 7371 59283 7429 59284
rect 8995 59324 9053 59325
rect 8995 59284 9004 59324
rect 9044 59284 9053 59324
rect 8995 59283 9053 59284
rect 10251 59324 10293 59333
rect 10251 59284 10252 59324
rect 10292 59284 10293 59324
rect 10251 59275 10293 59284
rect 10714 59324 10772 59325
rect 10714 59284 10723 59324
rect 10763 59284 10772 59324
rect 10714 59283 10772 59284
rect 10827 59324 10869 59333
rect 10827 59284 10828 59324
rect 10868 59284 10869 59324
rect 10827 59275 10869 59284
rect 11307 59324 11349 59333
rect 11307 59284 11308 59324
rect 11348 59284 11349 59324
rect 11307 59275 11349 59284
rect 11782 59324 11840 59325
rect 11782 59284 11791 59324
rect 11831 59284 11840 59324
rect 11782 59283 11840 59284
rect 12298 59324 12356 59325
rect 12298 59284 12307 59324
rect 12347 59284 12356 59324
rect 12298 59283 12356 59284
rect 13227 59324 13269 59333
rect 13227 59284 13228 59324
rect 13268 59284 13269 59324
rect 13227 59275 13269 59284
rect 14467 59324 14525 59325
rect 14467 59284 14476 59324
rect 14516 59284 14525 59324
rect 14467 59283 14525 59284
rect 14859 59324 14901 59333
rect 14859 59284 14860 59324
rect 14900 59284 14901 59324
rect 14859 59275 14901 59284
rect 16099 59324 16157 59325
rect 16099 59284 16108 59324
rect 16148 59284 16157 59324
rect 16099 59283 16157 59284
rect 16683 59324 16725 59333
rect 16683 59284 16684 59324
rect 16724 59284 16725 59324
rect 16683 59275 16725 59284
rect 17923 59324 17981 59325
rect 17923 59284 17932 59324
rect 17972 59284 17981 59324
rect 17923 59283 17981 59284
rect 18394 59324 18452 59325
rect 18394 59284 18403 59324
rect 18443 59284 18452 59324
rect 18394 59283 18452 59284
rect 18507 59324 18549 59333
rect 18507 59284 18508 59324
rect 18548 59284 18549 59324
rect 18507 59275 18549 59284
rect 18987 59324 19029 59333
rect 18987 59284 18988 59324
rect 19028 59284 19029 59324
rect 18987 59275 19029 59284
rect 19459 59324 19517 59325
rect 19459 59284 19468 59324
rect 19508 59284 19517 59324
rect 19459 59283 19517 59284
rect 19978 59324 20036 59325
rect 19978 59284 19987 59324
rect 20027 59284 20036 59324
rect 19978 59283 20036 59284
rect 3051 59240 3093 59249
rect 3051 59200 3052 59240
rect 3092 59200 3093 59240
rect 3051 59191 3093 59200
rect 5547 59240 5589 59249
rect 5547 59200 5548 59240
rect 5588 59200 5589 59240
rect 5547 59191 5589 59200
rect 18123 59240 18165 59249
rect 18123 59200 18124 59240
rect 18164 59200 18165 59240
rect 18123 59191 18165 59200
rect 1179 59156 1221 59165
rect 1179 59116 1180 59156
rect 1220 59116 1221 59156
rect 1179 59107 1221 59116
rect 3291 59156 3333 59165
rect 3291 59116 3292 59156
rect 3332 59116 3333 59156
rect 3291 59107 3333 59116
rect 7563 59156 7605 59165
rect 7563 59116 7564 59156
rect 7604 59116 7605 59156
rect 7563 59107 7605 59116
rect 8811 59156 8853 59165
rect 8811 59116 8812 59156
rect 8852 59116 8853 59156
rect 8811 59107 8853 59116
rect 12603 59156 12645 59165
rect 12603 59116 12604 59156
rect 12644 59116 12645 59156
rect 12603 59107 12645 59116
rect 16299 59156 16341 59165
rect 16299 59116 16300 59156
rect 16340 59116 16341 59156
rect 16299 59107 16341 59116
rect 20139 59156 20181 59165
rect 20139 59116 20140 59156
rect 20180 59116 20181 59156
rect 20139 59107 20181 59116
rect 1152 58988 20452 59012
rect 1152 58948 4928 58988
rect 4968 58948 5010 58988
rect 5050 58948 5092 58988
rect 5132 58948 5174 58988
rect 5214 58948 5256 58988
rect 5296 58948 20048 58988
rect 20088 58948 20130 58988
rect 20170 58948 20212 58988
rect 20252 58948 20294 58988
rect 20334 58948 20376 58988
rect 20416 58948 20452 58988
rect 1152 58924 20452 58948
rect 4011 58820 4053 58829
rect 4011 58780 4012 58820
rect 4052 58780 4053 58820
rect 4011 58771 4053 58780
rect 5787 58820 5829 58829
rect 5787 58780 5788 58820
rect 5828 58780 5829 58820
rect 5787 58771 5829 58780
rect 8235 58820 8277 58829
rect 8235 58780 8236 58820
rect 8276 58780 8277 58820
rect 8235 58771 8277 58780
rect 10714 58820 10772 58821
rect 10714 58780 10723 58820
rect 10763 58780 10772 58820
rect 10714 58779 10772 58780
rect 12987 58820 13029 58829
rect 12987 58780 12988 58820
rect 13028 58780 13029 58820
rect 12987 58771 13029 58780
rect 15051 58820 15093 58829
rect 15051 58780 15052 58820
rect 15092 58780 15093 58820
rect 15051 58771 15093 58780
rect 17163 58820 17205 58829
rect 17163 58780 17164 58820
rect 17204 58780 17205 58820
rect 17163 58771 17205 58780
rect 17931 58820 17973 58829
rect 17931 58780 17932 58820
rect 17972 58780 17973 58820
rect 17931 58771 17973 58780
rect 8410 58736 8468 58737
rect 8410 58696 8419 58736
rect 8459 58696 8468 58736
rect 8410 58695 8468 58696
rect 11259 58736 11301 58745
rect 11259 58696 11260 58736
rect 11300 58696 11301 58736
rect 11259 58687 11301 58696
rect 17341 58736 17383 58745
rect 17341 58696 17342 58736
rect 17382 58696 17383 58736
rect 17341 58687 17383 58696
rect 10172 58672 10214 58681
rect 2266 58652 2324 58653
rect 2266 58612 2275 58652
rect 2315 58612 2324 58652
rect 2266 58611 2324 58612
rect 2379 58652 2421 58661
rect 2379 58612 2380 58652
rect 2420 58612 2421 58652
rect 2379 58603 2421 58612
rect 2763 58652 2805 58661
rect 4203 58652 4245 58661
rect 6795 58652 6837 58661
rect 8602 58652 8660 58653
rect 9579 58652 9621 58661
rect 2763 58612 2764 58652
rect 2804 58612 2805 58652
rect 2763 58603 2805 58612
rect 3339 58643 3381 58652
rect 3339 58603 3340 58643
rect 3380 58603 3381 58643
rect 3339 58594 3381 58603
rect 3819 58643 3861 58652
rect 3819 58603 3820 58643
rect 3860 58603 3861 58643
rect 4203 58612 4204 58652
rect 4244 58612 4245 58652
rect 4203 58603 4245 58612
rect 5451 58643 5493 58652
rect 5451 58603 5452 58643
rect 5492 58603 5493 58643
rect 6795 58612 6796 58652
rect 6836 58612 6837 58652
rect 6795 58603 6837 58612
rect 8043 58643 8085 58652
rect 8043 58603 8044 58643
rect 8084 58603 8085 58643
rect 8602 58612 8611 58652
rect 8651 58612 8660 58652
rect 8602 58611 8660 58612
rect 9099 58643 9141 58652
rect 3819 58594 3861 58603
rect 5451 58594 5493 58603
rect 8043 58594 8085 58603
rect 9099 58603 9100 58643
rect 9140 58603 9141 58643
rect 9579 58612 9580 58652
rect 9620 58612 9621 58652
rect 9579 58603 9621 58612
rect 10059 58652 10101 58661
rect 10059 58612 10060 58652
rect 10100 58612 10101 58652
rect 10172 58632 10173 58672
rect 10213 58632 10214 58672
rect 10172 58623 10214 58632
rect 10555 58652 10613 58653
rect 10059 58603 10101 58612
rect 10555 58612 10564 58652
rect 10604 58612 10613 58652
rect 10555 58611 10613 58612
rect 10714 58652 10772 58653
rect 10714 58612 10723 58652
rect 10763 58612 10772 58652
rect 10714 58611 10772 58612
rect 10858 58652 10916 58653
rect 10858 58612 10867 58652
rect 10907 58612 10916 58652
rect 11104 58652 11162 58653
rect 10858 58611 10916 58612
rect 11002 58641 11060 58642
rect 9099 58594 9141 58603
rect 11002 58601 11011 58641
rect 11051 58601 11060 58641
rect 11104 58612 11113 58652
rect 11153 58612 11162 58652
rect 11104 58611 11162 58612
rect 11403 58652 11445 58661
rect 11403 58612 11404 58652
rect 11444 58612 11445 58652
rect 11403 58603 11445 58612
rect 13611 58652 13653 58661
rect 15418 58652 15476 58653
rect 13611 58612 13612 58652
rect 13652 58612 13653 58652
rect 13611 58603 13653 58612
rect 14859 58643 14901 58652
rect 14859 58603 14860 58643
rect 14900 58603 14901 58643
rect 15418 58612 15427 58652
rect 15467 58612 15476 58652
rect 15418 58611 15476 58612
rect 15531 58652 15573 58661
rect 15531 58612 15532 58652
rect 15572 58612 15573 58652
rect 15531 58603 15573 58612
rect 15915 58652 15957 58661
rect 17547 58652 17589 58661
rect 17835 58652 17877 58661
rect 15915 58612 15916 58652
rect 15956 58612 15957 58652
rect 15915 58603 15957 58612
rect 16491 58643 16533 58652
rect 16491 58603 16492 58643
rect 16532 58603 16533 58643
rect 11002 58600 11060 58601
rect 14859 58594 14901 58603
rect 16491 58594 16533 58603
rect 16971 58643 17013 58652
rect 16971 58603 16972 58643
rect 17012 58603 17013 58643
rect 17547 58612 17548 58652
rect 17588 58612 17589 58652
rect 17547 58603 17589 58612
rect 17643 58643 17685 58652
rect 17643 58603 17644 58643
rect 17684 58603 17685 58643
rect 17835 58612 17836 58652
rect 17876 58612 17877 58652
rect 17835 58603 17877 58612
rect 18027 58652 18069 58661
rect 18027 58612 18028 58652
rect 18068 58612 18069 58652
rect 18027 58603 18069 58612
rect 18699 58652 18741 58661
rect 18699 58612 18700 58652
rect 18740 58612 18741 58652
rect 18699 58603 18741 58612
rect 19947 58643 19989 58652
rect 19947 58603 19948 58643
rect 19988 58603 19989 58643
rect 16971 58594 17013 58603
rect 17643 58594 17685 58603
rect 19947 58594 19989 58603
rect 1419 58568 1461 58577
rect 1419 58528 1420 58568
rect 1460 58528 1461 58568
rect 1419 58519 1461 58528
rect 1803 58568 1845 58577
rect 1803 58528 1804 58568
rect 1844 58528 1845 58568
rect 1803 58519 1845 58528
rect 2859 58568 2901 58577
rect 2859 58528 2860 58568
rect 2900 58528 2901 58568
rect 2859 58519 2901 58528
rect 6027 58568 6069 58577
rect 6027 58528 6028 58568
rect 6068 58528 6069 58568
rect 6027 58519 6069 58528
rect 6411 58568 6453 58577
rect 6411 58528 6412 58568
rect 6452 58528 6453 58568
rect 6411 58519 6453 58528
rect 9675 58568 9717 58577
rect 9675 58528 9676 58568
rect 9716 58528 9717 58568
rect 9675 58519 9717 58528
rect 11787 58568 11829 58577
rect 11787 58528 11788 58568
rect 11828 58528 11829 58568
rect 11787 58519 11829 58528
rect 12747 58568 12789 58577
rect 12747 58528 12748 58568
rect 12788 58528 12789 58568
rect 12747 58519 12789 58528
rect 13131 58568 13173 58577
rect 13131 58528 13132 58568
rect 13172 58528 13173 58568
rect 13131 58519 13173 58528
rect 16011 58568 16053 58577
rect 16011 58528 16012 58568
rect 16052 58528 16053 58568
rect 16011 58519 16053 58528
rect 18411 58568 18453 58577
rect 18411 58528 18412 58568
rect 18452 58528 18453 58568
rect 18411 58519 18453 58528
rect 6171 58484 6213 58493
rect 6171 58444 6172 58484
rect 6212 58444 6213 58484
rect 6171 58435 6213 58444
rect 1179 58400 1221 58409
rect 1179 58360 1180 58400
rect 1220 58360 1221 58400
rect 1179 58351 1221 58360
rect 1563 58400 1605 58409
rect 1563 58360 1564 58400
rect 1604 58360 1605 58400
rect 1563 58351 1605 58360
rect 5643 58400 5685 58409
rect 5643 58360 5644 58400
rect 5684 58360 5685 58400
rect 5643 58351 5685 58360
rect 12027 58400 12069 58409
rect 12027 58360 12028 58400
rect 12068 58360 12069 58400
rect 12027 58351 12069 58360
rect 13371 58400 13413 58409
rect 13371 58360 13372 58400
rect 13412 58360 13413 58400
rect 13371 58351 13413 58360
rect 17338 58400 17396 58401
rect 17338 58360 17347 58400
rect 17387 58360 17396 58400
rect 17338 58359 17396 58360
rect 18171 58400 18213 58409
rect 18171 58360 18172 58400
rect 18212 58360 18213 58400
rect 18171 58351 18213 58360
rect 20139 58400 20181 58409
rect 20139 58360 20140 58400
rect 20180 58360 20181 58400
rect 20139 58351 20181 58360
rect 1152 58232 20448 58256
rect 1152 58192 3688 58232
rect 3728 58192 3770 58232
rect 3810 58192 3852 58232
rect 3892 58192 3934 58232
rect 3974 58192 4016 58232
rect 4056 58192 18808 58232
rect 18848 58192 18890 58232
rect 18930 58192 18972 58232
rect 19012 58192 19054 58232
rect 19094 58192 19136 58232
rect 19176 58192 20448 58232
rect 1152 58168 20448 58192
rect 5290 58064 5348 58065
rect 5290 58024 5299 58064
rect 5339 58024 5348 58064
rect 5290 58023 5348 58024
rect 11307 58064 11349 58073
rect 11307 58024 11308 58064
rect 11348 58024 11349 58064
rect 11307 58015 11349 58024
rect 11499 58064 11541 58073
rect 11499 58024 11500 58064
rect 11540 58024 11541 58064
rect 11499 58015 11541 58024
rect 14331 58064 14373 58073
rect 14331 58024 14332 58064
rect 14372 58024 14373 58064
rect 14331 58015 14373 58024
rect 15003 58064 15045 58073
rect 15003 58024 15004 58064
rect 15044 58024 15045 58064
rect 15003 58015 15045 58024
rect 15387 58064 15429 58073
rect 15387 58024 15388 58064
rect 15428 58024 15429 58064
rect 15387 58015 15429 58024
rect 14907 57980 14949 57989
rect 14907 57940 14908 57980
rect 14948 57940 14949 57980
rect 14907 57931 14949 57940
rect 4011 57896 4053 57905
rect 4011 57856 4012 57896
rect 4052 57856 4053 57896
rect 4011 57847 4053 57856
rect 7083 57896 7125 57905
rect 7083 57856 7084 57896
rect 7124 57856 7125 57896
rect 5067 57845 5109 57854
rect 7083 57847 7125 57856
rect 14091 57896 14133 57905
rect 14091 57856 14092 57896
rect 14132 57856 14133 57896
rect 1515 57812 1557 57821
rect 1515 57772 1516 57812
rect 1556 57772 1557 57812
rect 1515 57763 1557 57772
rect 2755 57812 2813 57813
rect 2755 57772 2764 57812
rect 2804 57772 2813 57812
rect 2755 57771 2813 57772
rect 3514 57812 3572 57813
rect 3514 57772 3523 57812
rect 3563 57772 3572 57812
rect 3514 57771 3572 57772
rect 3627 57812 3669 57821
rect 3627 57772 3628 57812
rect 3668 57772 3669 57812
rect 3627 57763 3669 57772
rect 4107 57812 4149 57821
rect 4107 57772 4108 57812
rect 4148 57772 4149 57812
rect 4107 57763 4149 57772
rect 4579 57812 4637 57813
rect 4579 57772 4588 57812
rect 4628 57772 4637 57812
rect 5067 57805 5068 57845
rect 5108 57805 5109 57845
rect 12118 57845 12160 57854
rect 14091 57847 14133 57856
rect 14667 57896 14709 57905
rect 14667 57856 14668 57896
rect 14708 57856 14709 57896
rect 14667 57847 14709 57856
rect 15243 57896 15285 57905
rect 15243 57856 15244 57896
rect 15284 57856 15285 57896
rect 15243 57847 15285 57856
rect 15627 57896 15669 57905
rect 15627 57856 15628 57896
rect 15668 57856 15669 57896
rect 15627 57847 15669 57856
rect 15819 57896 15861 57905
rect 18795 57896 18837 57905
rect 15819 57856 15820 57896
rect 15860 57856 15861 57896
rect 15819 57847 15861 57856
rect 16050 57887 16096 57896
rect 16050 57847 16051 57887
rect 16091 57847 16096 57887
rect 18795 57856 18796 57896
rect 18836 57856 18837 57896
rect 18795 57847 18837 57856
rect 5067 57796 5109 57805
rect 5627 57812 5685 57813
rect 4579 57771 4637 57772
rect 5627 57772 5636 57812
rect 5676 57772 5685 57812
rect 5627 57771 5685 57772
rect 6891 57812 6933 57821
rect 6891 57772 6892 57812
rect 6932 57772 6933 57812
rect 6891 57763 6933 57772
rect 7467 57812 7509 57821
rect 7467 57772 7468 57812
rect 7508 57772 7509 57812
rect 7467 57763 7509 57772
rect 8707 57812 8765 57813
rect 8707 57772 8716 57812
rect 8756 57772 8765 57812
rect 8707 57771 8765 57772
rect 9867 57812 9909 57821
rect 9867 57772 9868 57812
rect 9908 57772 9909 57812
rect 9867 57763 9909 57772
rect 11107 57812 11165 57813
rect 11107 57772 11116 57812
rect 11156 57772 11165 57812
rect 11107 57771 11165 57772
rect 11499 57812 11541 57821
rect 11499 57772 11500 57812
rect 11540 57772 11541 57812
rect 11499 57763 11541 57772
rect 11614 57812 11656 57821
rect 11614 57772 11615 57812
rect 11655 57772 11656 57812
rect 11614 57763 11656 57772
rect 11787 57812 11829 57821
rect 11787 57772 11788 57812
rect 11828 57772 11829 57812
rect 11787 57763 11829 57772
rect 11979 57812 12021 57821
rect 11979 57772 11980 57812
rect 12020 57772 12021 57812
rect 12118 57805 12119 57845
rect 12159 57805 12160 57845
rect 16050 57838 16096 57847
rect 12118 57796 12160 57805
rect 12459 57812 12501 57821
rect 11979 57763 12021 57772
rect 12459 57772 12460 57812
rect 12500 57772 12501 57812
rect 12459 57763 12501 57772
rect 13699 57812 13757 57813
rect 13699 57772 13708 57812
rect 13748 57772 13757 57812
rect 13699 57771 13757 57772
rect 15915 57812 15957 57821
rect 15915 57772 15916 57812
rect 15956 57772 15957 57812
rect 15915 57763 15957 57772
rect 16144 57812 16202 57813
rect 16144 57772 16153 57812
rect 16193 57772 16202 57812
rect 16144 57771 16202 57772
rect 16587 57812 16629 57821
rect 16587 57772 16588 57812
rect 16628 57772 16629 57812
rect 16587 57763 16629 57772
rect 17827 57812 17885 57813
rect 17827 57772 17836 57812
rect 17876 57772 17885 57812
rect 17827 57771 17885 57772
rect 18298 57812 18356 57813
rect 18298 57772 18307 57812
rect 18347 57772 18356 57812
rect 18298 57771 18356 57772
rect 18411 57812 18453 57821
rect 18411 57772 18412 57812
rect 18452 57772 18453 57812
rect 18411 57763 18453 57772
rect 18891 57812 18933 57821
rect 18891 57772 18892 57812
rect 18932 57772 18933 57812
rect 18891 57763 18933 57772
rect 19363 57812 19421 57813
rect 19363 57772 19372 57812
rect 19412 57772 19421 57812
rect 19363 57771 19421 57772
rect 19882 57812 19940 57813
rect 19882 57772 19891 57812
rect 19931 57772 19940 57812
rect 19882 57771 19940 57772
rect 2955 57728 2997 57737
rect 2955 57688 2956 57728
rect 2996 57688 2997 57728
rect 2955 57679 2997 57688
rect 18027 57728 18069 57737
rect 18027 57688 18028 57728
rect 18068 57688 18069 57728
rect 18027 57679 18069 57688
rect 5451 57644 5493 57653
rect 5451 57604 5452 57644
rect 5492 57604 5493 57644
rect 5451 57595 5493 57604
rect 7323 57644 7365 57653
rect 7323 57604 7324 57644
rect 7364 57604 7365 57644
rect 7323 57595 7365 57604
rect 8907 57644 8949 57653
rect 8907 57604 8908 57644
rect 8948 57604 8949 57644
rect 8907 57595 8949 57604
rect 11307 57644 11349 57653
rect 11307 57604 11308 57644
rect 11348 57604 11349 57644
rect 11307 57595 11349 57604
rect 12267 57644 12309 57653
rect 12267 57604 12268 57644
rect 12308 57604 12309 57644
rect 12267 57595 12309 57604
rect 13899 57644 13941 57653
rect 13899 57604 13900 57644
rect 13940 57604 13941 57644
rect 13899 57595 13941 57604
rect 20043 57644 20085 57653
rect 20043 57604 20044 57644
rect 20084 57604 20085 57644
rect 20043 57595 20085 57604
rect 1152 57476 20452 57500
rect 1152 57436 4928 57476
rect 4968 57436 5010 57476
rect 5050 57436 5092 57476
rect 5132 57436 5174 57476
rect 5214 57436 5256 57476
rect 5296 57436 20048 57476
rect 20088 57436 20130 57476
rect 20170 57436 20212 57476
rect 20252 57436 20294 57476
rect 20334 57436 20376 57476
rect 20416 57436 20452 57476
rect 1152 57412 20452 57436
rect 2235 57308 2277 57317
rect 2235 57268 2236 57308
rect 2276 57268 2277 57308
rect 2235 57259 2277 57268
rect 6747 57308 6789 57317
rect 6747 57268 6748 57308
rect 6788 57268 6789 57308
rect 6747 57259 6789 57268
rect 11307 57308 11349 57317
rect 11307 57268 11308 57308
rect 11348 57268 11349 57308
rect 11307 57259 11349 57268
rect 14955 57308 14997 57317
rect 14955 57268 14956 57308
rect 14996 57268 14997 57308
rect 14955 57259 14997 57268
rect 4203 57224 4245 57233
rect 4203 57184 4204 57224
rect 4244 57184 4245 57224
rect 4203 57175 4245 57184
rect 12939 57224 12981 57233
rect 12939 57184 12940 57224
rect 12980 57184 12981 57224
rect 12939 57175 12981 57184
rect 2763 57140 2805 57149
rect 4858 57140 4916 57141
rect 2763 57100 2764 57140
rect 2804 57100 2805 57140
rect 2763 57091 2805 57100
rect 4011 57131 4053 57140
rect 4011 57091 4012 57131
rect 4052 57091 4053 57131
rect 4858 57100 4867 57140
rect 4907 57100 4916 57140
rect 4858 57099 4916 57100
rect 4971 57140 5013 57149
rect 4971 57100 4972 57140
rect 5012 57100 5013 57140
rect 4971 57091 5013 57100
rect 5355 57140 5397 57149
rect 7738 57140 7796 57141
rect 5355 57100 5356 57140
rect 5396 57100 5397 57140
rect 5355 57091 5397 57100
rect 5931 57131 5973 57140
rect 5931 57091 5932 57131
rect 5972 57091 5973 57131
rect 4011 57082 4053 57091
rect 5931 57082 5973 57091
rect 6411 57131 6453 57140
rect 6411 57091 6412 57131
rect 6452 57091 6453 57131
rect 7738 57100 7747 57140
rect 7787 57100 7796 57140
rect 7738 57099 7796 57100
rect 7851 57140 7893 57149
rect 7851 57100 7852 57140
rect 7892 57100 7893 57140
rect 7851 57091 7893 57100
rect 8235 57140 8277 57149
rect 9867 57140 9909 57149
rect 11499 57140 11541 57149
rect 13210 57140 13268 57141
rect 8235 57100 8236 57140
rect 8276 57100 8277 57140
rect 8235 57091 8277 57100
rect 8811 57131 8853 57140
rect 8811 57091 8812 57131
rect 8852 57091 8853 57131
rect 6411 57082 6453 57091
rect 8811 57082 8853 57091
rect 9291 57131 9333 57140
rect 9291 57091 9292 57131
rect 9332 57091 9333 57131
rect 9867 57100 9868 57140
rect 9908 57100 9909 57140
rect 9867 57091 9909 57100
rect 11115 57131 11157 57140
rect 11115 57091 11116 57131
rect 11156 57091 11157 57131
rect 11499 57100 11500 57140
rect 11540 57100 11541 57140
rect 11499 57091 11541 57100
rect 12747 57131 12789 57140
rect 12747 57091 12748 57131
rect 12788 57091 12789 57131
rect 13210 57100 13219 57140
rect 13259 57100 13268 57140
rect 13210 57099 13268 57100
rect 13323 57140 13365 57149
rect 13323 57100 13324 57140
rect 13364 57100 13365 57140
rect 13323 57091 13365 57100
rect 13707 57140 13749 57149
rect 15339 57140 15381 57149
rect 16971 57140 17013 57149
rect 18603 57140 18645 57149
rect 13707 57100 13708 57140
rect 13748 57100 13749 57140
rect 13707 57091 13749 57100
rect 14283 57131 14325 57140
rect 14283 57091 14284 57131
rect 14324 57091 14325 57131
rect 9291 57082 9333 57091
rect 11115 57082 11157 57091
rect 12747 57082 12789 57091
rect 14283 57082 14325 57091
rect 14763 57131 14805 57140
rect 14763 57091 14764 57131
rect 14804 57091 14805 57131
rect 15339 57100 15340 57140
rect 15380 57100 15381 57140
rect 15339 57091 15381 57100
rect 16587 57131 16629 57140
rect 16587 57091 16588 57131
rect 16628 57091 16629 57131
rect 16971 57100 16972 57140
rect 17012 57100 17013 57140
rect 16971 57091 17013 57100
rect 18219 57131 18261 57140
rect 18219 57091 18220 57131
rect 18260 57091 18261 57131
rect 18603 57100 18604 57140
rect 18644 57100 18645 57140
rect 18603 57091 18645 57100
rect 19851 57131 19893 57140
rect 19851 57091 19852 57131
rect 19892 57091 19893 57131
rect 14763 57082 14805 57091
rect 16587 57082 16629 57091
rect 18219 57082 18261 57091
rect 19851 57082 19893 57091
rect 1419 57056 1461 57065
rect 1419 57016 1420 57056
rect 1460 57016 1461 57056
rect 1419 57007 1461 57016
rect 1803 57056 1845 57065
rect 1803 57016 1804 57056
rect 1844 57016 1845 57056
rect 1803 57007 1845 57016
rect 1995 57056 2037 57065
rect 1995 57016 1996 57056
rect 2036 57016 2037 57056
rect 1995 57007 2037 57016
rect 2571 57056 2613 57065
rect 2571 57016 2572 57056
rect 2612 57016 2613 57056
rect 2571 57007 2613 57016
rect 4587 57056 4629 57065
rect 4587 57016 4588 57056
rect 4628 57016 4629 57056
rect 4587 57007 4629 57016
rect 5451 57056 5493 57065
rect 5451 57016 5452 57056
rect 5492 57016 5493 57056
rect 5451 57007 5493 57016
rect 6634 57056 6692 57057
rect 6634 57016 6643 57056
rect 6683 57016 6692 57056
rect 6634 57015 6692 57016
rect 6987 57056 7029 57065
rect 6987 57016 6988 57056
rect 7028 57016 7029 57056
rect 6987 57007 7029 57016
rect 8331 57056 8373 57065
rect 8331 57016 8332 57056
rect 8372 57016 8373 57056
rect 8331 57007 8373 57016
rect 13803 57056 13845 57065
rect 13803 57016 13804 57056
rect 13844 57016 13845 57056
rect 13803 57007 13845 57016
rect 1179 56888 1221 56897
rect 1179 56848 1180 56888
rect 1220 56848 1221 56888
rect 1179 56839 1221 56848
rect 1563 56888 1605 56897
rect 1563 56848 1564 56888
rect 1604 56848 1605 56888
rect 1563 56839 1605 56848
rect 2331 56888 2373 56897
rect 2331 56848 2332 56888
rect 2372 56848 2373 56888
rect 2331 56839 2373 56848
rect 4347 56888 4389 56897
rect 4347 56848 4348 56888
rect 4388 56848 4389 56888
rect 4347 56839 4389 56848
rect 9514 56888 9572 56889
rect 9514 56848 9523 56888
rect 9563 56848 9572 56888
rect 9514 56847 9572 56848
rect 16779 56888 16821 56897
rect 16779 56848 16780 56888
rect 16820 56848 16821 56888
rect 16779 56839 16821 56848
rect 18411 56888 18453 56897
rect 18411 56848 18412 56888
rect 18452 56848 18453 56888
rect 18411 56839 18453 56848
rect 20043 56888 20085 56897
rect 20043 56848 20044 56888
rect 20084 56848 20085 56888
rect 20043 56839 20085 56848
rect 1152 56720 20448 56744
rect 1152 56680 3688 56720
rect 3728 56680 3770 56720
rect 3810 56680 3852 56720
rect 3892 56680 3934 56720
rect 3974 56680 4016 56720
rect 4056 56680 18808 56720
rect 18848 56680 18890 56720
rect 18930 56680 18972 56720
rect 19012 56680 19054 56720
rect 19094 56680 19136 56720
rect 19176 56680 20448 56720
rect 1152 56656 20448 56680
rect 8043 56552 8085 56561
rect 8043 56512 8044 56552
rect 8084 56512 8085 56552
rect 8043 56503 8085 56512
rect 10107 56552 10149 56561
rect 10107 56512 10108 56552
rect 10148 56512 10149 56552
rect 10107 56503 10149 56512
rect 13035 56552 13077 56561
rect 13035 56512 13036 56552
rect 13076 56512 13077 56552
rect 13035 56503 13077 56512
rect 17979 56552 18021 56561
rect 17979 56512 17980 56552
rect 18020 56512 18021 56552
rect 17979 56503 18021 56512
rect 5403 56468 5445 56477
rect 5403 56428 5404 56468
rect 5444 56428 5445 56468
rect 5403 56419 5445 56428
rect 17307 56468 17349 56477
rect 17307 56428 17308 56468
rect 17348 56428 17349 56468
rect 17307 56419 17349 56428
rect 1419 56384 1461 56393
rect 1419 56344 1420 56384
rect 1460 56344 1461 56384
rect 1419 56335 1461 56344
rect 4011 56384 4053 56393
rect 4011 56344 4012 56384
rect 4052 56344 4053 56384
rect 4011 56335 4053 56344
rect 5290 56384 5348 56385
rect 5290 56344 5299 56384
rect 5339 56344 5348 56384
rect 5290 56343 5348 56344
rect 5643 56384 5685 56393
rect 5643 56344 5644 56384
rect 5684 56344 5685 56384
rect 5643 56335 5685 56344
rect 6411 56384 6453 56393
rect 6411 56344 6412 56384
rect 6452 56344 6453 56384
rect 6411 56335 6453 56344
rect 10347 56384 10389 56393
rect 10347 56344 10348 56384
rect 10388 56344 10389 56384
rect 10347 56335 10389 56344
rect 13803 56384 13845 56393
rect 13803 56344 13804 56384
rect 13844 56344 13845 56384
rect 13803 56335 13845 56344
rect 15819 56384 15861 56393
rect 15819 56344 15820 56384
rect 15860 56344 15861 56384
rect 15819 56335 15861 56344
rect 17547 56384 17589 56393
rect 17547 56344 17548 56384
rect 17588 56344 17589 56384
rect 17547 56335 17589 56344
rect 17739 56384 17781 56393
rect 17739 56344 17740 56384
rect 17780 56344 17781 56384
rect 17739 56335 17781 56344
rect 18699 56384 18741 56393
rect 18699 56344 18700 56384
rect 18740 56344 18741 56384
rect 18699 56335 18741 56344
rect 20139 56384 20181 56393
rect 20139 56344 20140 56384
rect 20180 56344 20181 56384
rect 19755 56333 19797 56342
rect 20139 56335 20181 56344
rect 1707 56300 1749 56309
rect 1707 56260 1708 56300
rect 1748 56260 1749 56300
rect 1707 56251 1749 56260
rect 2947 56300 3005 56301
rect 2947 56260 2956 56300
rect 2996 56260 3005 56300
rect 2947 56259 3005 56260
rect 3514 56300 3572 56301
rect 3514 56260 3523 56300
rect 3563 56260 3572 56300
rect 3514 56259 3572 56260
rect 3627 56300 3669 56309
rect 3627 56260 3628 56300
rect 3668 56260 3669 56300
rect 3627 56251 3669 56260
rect 4107 56300 4149 56309
rect 4107 56260 4108 56300
rect 4148 56260 4149 56300
rect 4107 56251 4149 56260
rect 4579 56300 4637 56301
rect 4579 56260 4588 56300
rect 4628 56260 4637 56300
rect 4579 56259 4637 56260
rect 5098 56300 5156 56301
rect 5098 56260 5107 56300
rect 5147 56260 5156 56300
rect 5098 56259 5156 56260
rect 6608 56300 6650 56309
rect 6608 56260 6609 56300
rect 6649 56260 6650 56300
rect 6608 56251 6650 56260
rect 7843 56300 7901 56301
rect 7843 56260 7852 56300
rect 7892 56260 7901 56300
rect 7843 56259 7901 56260
rect 8523 56300 8565 56309
rect 8523 56260 8524 56300
rect 8564 56260 8565 56300
rect 8523 56251 8565 56260
rect 9763 56300 9821 56301
rect 9763 56260 9772 56300
rect 9812 56260 9821 56300
rect 9763 56259 9821 56260
rect 11595 56300 11637 56309
rect 11595 56260 11596 56300
rect 11636 56260 11637 56300
rect 11595 56251 11637 56260
rect 12835 56300 12893 56301
rect 12835 56260 12844 56300
rect 12884 56260 12893 56300
rect 12835 56259 12893 56260
rect 13306 56300 13364 56301
rect 13306 56260 13315 56300
rect 13355 56260 13364 56300
rect 13306 56259 13364 56260
rect 13419 56300 13461 56309
rect 13419 56260 13420 56300
rect 13460 56260 13461 56300
rect 13419 56251 13461 56260
rect 13899 56300 13941 56309
rect 13899 56260 13900 56300
rect 13940 56260 13941 56300
rect 13899 56251 13941 56260
rect 14371 56300 14429 56301
rect 14371 56260 14380 56300
rect 14420 56260 14429 56300
rect 14371 56259 14429 56260
rect 14859 56300 14917 56301
rect 14859 56260 14868 56300
rect 14908 56260 14917 56300
rect 14859 56259 14917 56260
rect 15322 56300 15380 56301
rect 15322 56260 15331 56300
rect 15371 56260 15380 56300
rect 15322 56259 15380 56260
rect 15435 56300 15477 56309
rect 15435 56260 15436 56300
rect 15476 56260 15477 56300
rect 15435 56251 15477 56260
rect 15915 56300 15957 56309
rect 15915 56260 15916 56300
rect 15956 56260 15957 56300
rect 15915 56251 15957 56260
rect 16387 56300 16445 56301
rect 16387 56260 16396 56300
rect 16436 56260 16445 56300
rect 16387 56259 16445 56260
rect 16875 56300 16933 56301
rect 16875 56260 16884 56300
rect 16924 56260 16933 56300
rect 16875 56259 16933 56260
rect 18202 56300 18260 56301
rect 18202 56260 18211 56300
rect 18251 56260 18260 56300
rect 18202 56259 18260 56260
rect 18315 56300 18357 56309
rect 18315 56260 18316 56300
rect 18356 56260 18357 56300
rect 18315 56251 18357 56260
rect 18795 56300 18837 56309
rect 18795 56260 18796 56300
rect 18836 56260 18837 56300
rect 18795 56251 18837 56260
rect 19267 56300 19325 56301
rect 19267 56260 19276 56300
rect 19316 56260 19325 56300
rect 19755 56293 19756 56333
rect 19796 56293 19797 56333
rect 19755 56284 19797 56293
rect 19267 56259 19325 56260
rect 1179 56216 1221 56225
rect 1179 56176 1180 56216
rect 1220 56176 1221 56216
rect 1179 56167 1221 56176
rect 3147 56216 3189 56225
rect 3147 56176 3148 56216
rect 3188 56176 3189 56216
rect 3147 56167 3189 56176
rect 20379 56216 20421 56225
rect 20379 56176 20380 56216
rect 20420 56176 20421 56216
rect 20379 56167 20421 56176
rect 6171 56132 6213 56141
rect 6171 56092 6172 56132
rect 6212 56092 6213 56132
rect 6171 56083 6213 56092
rect 9963 56132 10005 56141
rect 9963 56092 9964 56132
rect 10004 56092 10005 56132
rect 9963 56083 10005 56092
rect 15051 56132 15093 56141
rect 15051 56092 15052 56132
rect 15092 56092 15093 56132
rect 15051 56083 15093 56092
rect 17067 56132 17109 56141
rect 17067 56092 17068 56132
rect 17108 56092 17109 56132
rect 17067 56083 17109 56092
rect 19947 56132 19989 56141
rect 19947 56092 19948 56132
rect 19988 56092 19989 56132
rect 19947 56083 19989 56092
rect 1152 55964 20452 55988
rect 1152 55924 4928 55964
rect 4968 55924 5010 55964
rect 5050 55924 5092 55964
rect 5132 55924 5174 55964
rect 5214 55924 5256 55964
rect 5296 55924 20048 55964
rect 20088 55924 20130 55964
rect 20170 55924 20212 55964
rect 20252 55924 20294 55964
rect 20334 55924 20376 55964
rect 20416 55924 20452 55964
rect 1152 55900 20452 55924
rect 3291 55796 3333 55805
rect 3291 55756 3292 55796
rect 3332 55756 3333 55796
rect 3291 55747 3333 55756
rect 5355 55796 5397 55805
rect 5355 55756 5356 55796
rect 5396 55756 5397 55796
rect 5355 55747 5397 55756
rect 5499 55796 5541 55805
rect 5499 55756 5500 55796
rect 5540 55756 5541 55796
rect 5499 55747 5541 55756
rect 17067 55796 17109 55805
rect 17067 55756 17068 55796
rect 17108 55756 17109 55796
rect 17067 55747 17109 55756
rect 17211 55796 17253 55805
rect 17211 55756 17212 55796
rect 17252 55756 17253 55796
rect 17211 55747 17253 55756
rect 2859 55712 2901 55721
rect 2859 55672 2860 55712
rect 2900 55672 2901 55712
rect 2859 55663 2901 55672
rect 8043 55712 8085 55721
rect 8043 55672 8044 55712
rect 8084 55672 8085 55712
rect 8043 55663 8085 55672
rect 15051 55712 15093 55721
rect 15051 55672 15052 55712
rect 15092 55672 15093 55712
rect 15051 55663 15093 55672
rect 1419 55628 1461 55637
rect 3915 55628 3957 55637
rect 6603 55628 6645 55637
rect 8410 55628 8468 55629
rect 1419 55588 1420 55628
rect 1460 55588 1461 55628
rect 1419 55579 1461 55588
rect 2667 55619 2709 55628
rect 2667 55579 2668 55619
rect 2708 55579 2709 55619
rect 3915 55588 3916 55628
rect 3956 55588 3957 55628
rect 3915 55579 3957 55588
rect 5163 55619 5205 55628
rect 5163 55579 5164 55619
rect 5204 55579 5205 55619
rect 6603 55588 6604 55628
rect 6644 55588 6645 55628
rect 6603 55579 6645 55588
rect 7851 55619 7893 55628
rect 7851 55579 7852 55619
rect 7892 55579 7893 55619
rect 8410 55588 8419 55628
rect 8459 55588 8468 55628
rect 8410 55587 8468 55588
rect 8523 55628 8565 55637
rect 8523 55588 8524 55628
rect 8564 55588 8565 55628
rect 8523 55579 8565 55588
rect 8907 55628 8949 55637
rect 12075 55628 12117 55637
rect 8907 55588 8908 55628
rect 8948 55588 8949 55628
rect 8907 55579 8949 55588
rect 9483 55619 9525 55628
rect 9483 55579 9484 55619
rect 9524 55579 9525 55619
rect 2667 55570 2709 55579
rect 5163 55570 5205 55579
rect 7851 55570 7893 55579
rect 9483 55570 9525 55579
rect 9963 55619 10005 55628
rect 9963 55579 9964 55619
rect 10004 55579 10005 55619
rect 9963 55570 10005 55579
rect 10827 55619 10869 55628
rect 10827 55579 10828 55619
rect 10868 55579 10869 55619
rect 12075 55588 12076 55628
rect 12116 55588 12117 55628
rect 12075 55579 12117 55588
rect 13611 55628 13653 55637
rect 15322 55628 15380 55629
rect 13611 55588 13612 55628
rect 13652 55588 13653 55628
rect 13611 55579 13653 55588
rect 14859 55619 14901 55628
rect 14859 55579 14860 55619
rect 14900 55579 14901 55619
rect 15322 55588 15331 55628
rect 15371 55588 15380 55628
rect 15322 55587 15380 55588
rect 15435 55628 15477 55637
rect 15435 55588 15436 55628
rect 15476 55588 15477 55628
rect 15435 55579 15477 55588
rect 15819 55628 15861 55637
rect 18027 55628 18069 55637
rect 15819 55588 15820 55628
rect 15860 55588 15861 55628
rect 15819 55579 15861 55588
rect 16395 55619 16437 55628
rect 16395 55579 16396 55619
rect 16436 55579 16437 55619
rect 10827 55570 10869 55579
rect 14859 55570 14901 55579
rect 16395 55570 16437 55579
rect 16875 55619 16917 55628
rect 16875 55579 16876 55619
rect 16916 55579 16917 55619
rect 18027 55588 18028 55628
rect 18068 55588 18069 55628
rect 18027 55579 18069 55588
rect 19275 55619 19317 55628
rect 19275 55579 19276 55619
rect 19316 55579 19317 55619
rect 16875 55570 16917 55579
rect 19275 55570 19317 55579
rect 3051 55544 3093 55553
rect 3051 55504 3052 55544
rect 3092 55504 3093 55544
rect 3051 55495 3093 55504
rect 3627 55544 3669 55553
rect 3627 55504 3628 55544
rect 3668 55504 3669 55544
rect 3627 55495 3669 55504
rect 5739 55544 5781 55553
rect 5739 55504 5740 55544
rect 5780 55504 5781 55544
rect 5739 55495 5781 55504
rect 5931 55544 5973 55553
rect 5931 55504 5932 55544
rect 5972 55504 5973 55544
rect 5931 55495 5973 55504
rect 9003 55544 9045 55553
rect 9003 55504 9004 55544
rect 9044 55504 9045 55544
rect 9003 55495 9045 55504
rect 12267 55544 12309 55553
rect 12267 55504 12268 55544
rect 12308 55504 12309 55544
rect 12267 55495 12309 55504
rect 15915 55544 15957 55553
rect 15915 55504 15916 55544
rect 15956 55504 15957 55544
rect 15915 55495 15957 55504
rect 17451 55544 17493 55553
rect 17451 55504 17452 55544
rect 17492 55504 17493 55544
rect 17451 55495 17493 55504
rect 17643 55544 17685 55553
rect 17643 55504 17644 55544
rect 17684 55504 17685 55544
rect 17643 55495 17685 55504
rect 19755 55544 19797 55553
rect 19755 55504 19756 55544
rect 19796 55504 19797 55544
rect 19755 55495 19797 55504
rect 20139 55544 20181 55553
rect 20139 55504 20140 55544
rect 20180 55504 20181 55544
rect 20139 55495 20181 55504
rect 3387 55460 3429 55469
rect 3387 55420 3388 55460
rect 3428 55420 3429 55460
rect 3387 55411 3429 55420
rect 19995 55460 20037 55469
rect 19995 55420 19996 55460
rect 20036 55420 20037 55460
rect 19995 55411 20037 55420
rect 6171 55376 6213 55385
rect 6171 55336 6172 55376
rect 6212 55336 6213 55376
rect 6171 55327 6213 55336
rect 10186 55376 10244 55377
rect 10186 55336 10195 55376
rect 10235 55336 10244 55376
rect 10186 55335 10244 55336
rect 10635 55376 10677 55385
rect 10635 55336 10636 55376
rect 10676 55336 10677 55376
rect 10635 55327 10677 55336
rect 12507 55376 12549 55385
rect 12507 55336 12508 55376
rect 12548 55336 12549 55376
rect 12507 55327 12549 55336
rect 17883 55376 17925 55385
rect 17883 55336 17884 55376
rect 17924 55336 17925 55376
rect 17883 55327 17925 55336
rect 19467 55376 19509 55385
rect 19467 55336 19468 55376
rect 19508 55336 19509 55376
rect 19467 55327 19509 55336
rect 20379 55376 20421 55385
rect 20379 55336 20380 55376
rect 20420 55336 20421 55376
rect 20379 55327 20421 55336
rect 1152 55208 20448 55232
rect 1152 55168 3688 55208
rect 3728 55168 3770 55208
rect 3810 55168 3852 55208
rect 3892 55168 3934 55208
rect 3974 55168 4016 55208
rect 4056 55168 18808 55208
rect 18848 55168 18890 55208
rect 18930 55168 18972 55208
rect 19012 55168 19054 55208
rect 19094 55168 19136 55208
rect 19176 55168 20448 55208
rect 1152 55144 20448 55168
rect 13419 55040 13461 55049
rect 13419 55000 13420 55040
rect 13460 55000 13461 55040
rect 13419 54991 13461 55000
rect 15051 55040 15093 55049
rect 15051 55000 15052 55040
rect 15092 55000 15093 55040
rect 15051 54991 15093 55000
rect 16779 55040 16821 55049
rect 16779 55000 16780 55040
rect 16820 55000 16821 55040
rect 16779 54991 16821 55000
rect 20331 54956 20373 54965
rect 20331 54916 20332 54956
rect 20372 54916 20373 54956
rect 20331 54907 20373 54916
rect 10059 54872 10101 54881
rect 10059 54832 10060 54872
rect 10100 54832 10101 54872
rect 10059 54823 10101 54832
rect 11338 54872 11396 54873
rect 11338 54832 11347 54872
rect 11387 54832 11396 54872
rect 11338 54831 11396 54832
rect 1419 54788 1461 54797
rect 1419 54748 1420 54788
rect 1460 54748 1461 54788
rect 1419 54739 1461 54748
rect 2659 54788 2717 54789
rect 2659 54748 2668 54788
rect 2708 54748 2717 54788
rect 2659 54747 2717 54748
rect 3051 54788 3093 54797
rect 3051 54748 3052 54788
rect 3092 54748 3093 54788
rect 3051 54739 3093 54748
rect 3190 54788 3232 54797
rect 3190 54748 3191 54788
rect 3231 54748 3232 54788
rect 3190 54739 3232 54748
rect 3531 54788 3573 54797
rect 3531 54748 3532 54788
rect 3572 54748 3573 54788
rect 3531 54739 3573 54748
rect 3706 54788 3764 54789
rect 3706 54748 3715 54788
rect 3755 54748 3764 54788
rect 3706 54747 3764 54748
rect 3819 54788 3861 54797
rect 3819 54748 3820 54788
rect 3860 54748 3861 54788
rect 3819 54739 3861 54748
rect 4011 54788 4053 54797
rect 4011 54748 4012 54788
rect 4052 54748 4053 54788
rect 4011 54739 4053 54748
rect 4299 54788 4341 54797
rect 4299 54748 4300 54788
rect 4340 54748 4341 54788
rect 4299 54739 4341 54748
rect 5539 54788 5597 54789
rect 5539 54748 5548 54788
rect 5588 54748 5597 54788
rect 5539 54747 5597 54748
rect 6219 54788 6261 54797
rect 6219 54748 6220 54788
rect 6260 54748 6261 54788
rect 6219 54739 6261 54748
rect 7459 54788 7517 54789
rect 7459 54748 7468 54788
rect 7508 54748 7517 54788
rect 7459 54747 7517 54748
rect 7851 54788 7893 54797
rect 7851 54748 7852 54788
rect 7892 54748 7893 54788
rect 7851 54739 7893 54748
rect 9091 54788 9149 54789
rect 9091 54748 9100 54788
rect 9140 54748 9149 54788
rect 9091 54747 9149 54748
rect 9562 54788 9620 54789
rect 9562 54748 9571 54788
rect 9611 54748 9620 54788
rect 9562 54747 9620 54748
rect 9675 54788 9717 54797
rect 9675 54748 9676 54788
rect 9716 54748 9717 54788
rect 9675 54739 9717 54748
rect 10155 54788 10197 54797
rect 10155 54748 10156 54788
rect 10196 54748 10197 54788
rect 10155 54739 10197 54748
rect 10627 54788 10685 54789
rect 10627 54748 10636 54788
rect 10676 54748 10685 54788
rect 10627 54747 10685 54748
rect 11146 54788 11204 54789
rect 11146 54748 11155 54788
rect 11195 54748 11204 54788
rect 11146 54747 11204 54748
rect 11979 54788 12021 54797
rect 11979 54748 11980 54788
rect 12020 54748 12021 54788
rect 11979 54739 12021 54748
rect 13219 54788 13277 54789
rect 13219 54748 13228 54788
rect 13268 54748 13277 54788
rect 13219 54747 13277 54748
rect 13611 54788 13653 54797
rect 13611 54748 13612 54788
rect 13652 54748 13653 54788
rect 13611 54739 13653 54748
rect 14851 54788 14909 54789
rect 14851 54748 14860 54788
rect 14900 54748 14909 54788
rect 14851 54747 14909 54748
rect 15339 54788 15381 54797
rect 15339 54748 15340 54788
rect 15380 54748 15381 54788
rect 15339 54739 15381 54748
rect 16579 54788 16637 54789
rect 16579 54748 16588 54788
rect 16628 54748 16637 54788
rect 16579 54747 16637 54748
rect 17067 54788 17109 54797
rect 17067 54748 17068 54788
rect 17108 54748 17109 54788
rect 17067 54739 17109 54748
rect 18307 54788 18365 54789
rect 18307 54748 18316 54788
rect 18356 54748 18365 54788
rect 18307 54747 18365 54748
rect 18891 54788 18933 54797
rect 18891 54748 18892 54788
rect 18932 54748 18933 54788
rect 18891 54739 18933 54748
rect 20131 54788 20189 54789
rect 20131 54748 20140 54788
rect 20180 54748 20189 54788
rect 20131 54747 20189 54748
rect 3610 54704 3668 54705
rect 3610 54664 3619 54704
rect 3659 54664 3668 54704
rect 3610 54663 3668 54664
rect 2859 54620 2901 54629
rect 2859 54580 2860 54620
rect 2900 54580 2901 54620
rect 2859 54571 2901 54580
rect 3339 54620 3381 54629
rect 3339 54580 3340 54620
rect 3380 54580 3381 54620
rect 3339 54571 3381 54580
rect 4155 54620 4197 54629
rect 4155 54580 4156 54620
rect 4196 54580 4197 54620
rect 4155 54571 4197 54580
rect 5739 54620 5781 54629
rect 5739 54580 5740 54620
rect 5780 54580 5781 54620
rect 5739 54571 5781 54580
rect 7659 54620 7701 54629
rect 7659 54580 7660 54620
rect 7700 54580 7701 54620
rect 7659 54571 7701 54580
rect 9291 54620 9333 54629
rect 9291 54580 9292 54620
rect 9332 54580 9333 54620
rect 9291 54571 9333 54580
rect 18507 54620 18549 54629
rect 18507 54580 18508 54620
rect 18548 54580 18549 54620
rect 18507 54571 18549 54580
rect 1152 54452 20452 54476
rect 1152 54412 4928 54452
rect 4968 54412 5010 54452
rect 5050 54412 5092 54452
rect 5132 54412 5174 54452
rect 5214 54412 5256 54452
rect 5296 54412 20048 54452
rect 20088 54412 20130 54452
rect 20170 54412 20212 54452
rect 20252 54412 20294 54452
rect 20334 54412 20376 54452
rect 20416 54412 20452 54452
rect 1152 54388 20452 54412
rect 1947 54284 1989 54293
rect 1947 54244 1948 54284
rect 1988 54244 1989 54284
rect 1947 54235 1989 54244
rect 7947 54284 7989 54293
rect 7947 54244 7948 54284
rect 7988 54244 7989 54284
rect 7947 54235 7989 54244
rect 11307 54284 11349 54293
rect 11307 54244 11308 54284
rect 11348 54244 11349 54284
rect 11307 54235 11349 54244
rect 12891 54284 12933 54293
rect 12891 54244 12892 54284
rect 12932 54244 12933 54284
rect 12891 54235 12933 54244
rect 17019 54284 17061 54293
rect 17019 54244 17020 54284
rect 17060 54244 17061 54284
rect 17019 54235 17061 54244
rect 17691 54284 17733 54293
rect 17691 54244 17692 54284
rect 17732 54244 17733 54284
rect 17691 54235 17733 54244
rect 20043 54284 20085 54293
rect 20043 54244 20044 54284
rect 20084 54244 20085 54284
rect 20043 54235 20085 54244
rect 14859 54200 14901 54209
rect 4002 54191 4048 54200
rect 4002 54151 4003 54191
rect 4043 54151 4048 54191
rect 14859 54160 14860 54200
rect 14900 54160 14901 54200
rect 14859 54151 14901 54160
rect 17787 54200 17829 54209
rect 17787 54160 17788 54200
rect 17828 54160 17829 54200
rect 17787 54151 17829 54160
rect 4002 54142 4048 54151
rect 2091 54116 2133 54125
rect 4090 54116 4148 54117
rect 2091 54076 2092 54116
rect 2132 54076 2133 54116
rect 2091 54067 2133 54076
rect 3339 54107 3381 54116
rect 3339 54067 3340 54107
rect 3380 54067 3381 54107
rect 3339 54058 3381 54067
rect 3698 54105 3740 54114
rect 3698 54065 3699 54105
rect 3739 54065 3740 54105
rect 3698 54056 3740 54065
rect 3819 54107 3861 54116
rect 3819 54067 3820 54107
rect 3860 54067 3861 54107
rect 4090 54076 4099 54116
rect 4139 54076 4148 54116
rect 4090 54075 4148 54076
rect 4224 54116 4282 54117
rect 4224 54076 4233 54116
rect 4273 54076 4282 54116
rect 4224 54075 4282 54076
rect 4491 54116 4533 54125
rect 6202 54116 6260 54117
rect 4491 54076 4492 54116
rect 4532 54076 4533 54116
rect 4491 54067 4533 54076
rect 5739 54107 5781 54116
rect 5739 54067 5740 54107
rect 5780 54067 5781 54107
rect 6202 54076 6211 54116
rect 6251 54076 6260 54116
rect 6202 54075 6260 54076
rect 6315 54116 6357 54125
rect 6315 54076 6316 54116
rect 6356 54076 6357 54116
rect 6315 54067 6357 54076
rect 6699 54116 6741 54125
rect 9370 54116 9428 54117
rect 6699 54076 6700 54116
rect 6740 54076 6741 54116
rect 6699 54067 6741 54076
rect 7275 54107 7317 54116
rect 7275 54067 7276 54107
rect 7316 54067 7317 54107
rect 3819 54058 3861 54067
rect 5739 54058 5781 54067
rect 7275 54058 7317 54067
rect 7755 54107 7797 54116
rect 7755 54067 7756 54107
rect 7796 54067 7797 54107
rect 9370 54076 9379 54116
rect 9419 54076 9428 54116
rect 9370 54075 9428 54076
rect 9488 54116 9530 54125
rect 9488 54076 9489 54116
rect 9529 54076 9530 54116
rect 9488 54067 9530 54076
rect 9867 54116 9909 54125
rect 12747 54116 12789 54125
rect 9867 54076 9868 54116
rect 9908 54076 9909 54116
rect 9867 54067 9909 54076
rect 10443 54107 10485 54116
rect 10443 54067 10444 54107
rect 10484 54067 10485 54107
rect 7755 54058 7797 54067
rect 10443 54058 10485 54067
rect 10923 54107 10965 54116
rect 10923 54067 10924 54107
rect 10964 54067 10965 54107
rect 10923 54058 10965 54067
rect 11499 54107 11541 54116
rect 11499 54067 11500 54107
rect 11540 54067 11541 54107
rect 12747 54076 12748 54116
rect 12788 54076 12789 54116
rect 12747 54067 12789 54076
rect 13419 54116 13461 54125
rect 15130 54116 15188 54117
rect 13419 54076 13420 54116
rect 13460 54076 13461 54116
rect 13419 54067 13461 54076
rect 14667 54107 14709 54116
rect 14667 54067 14668 54107
rect 14708 54067 14709 54107
rect 15130 54076 15139 54116
rect 15179 54076 15188 54116
rect 15130 54075 15188 54076
rect 15243 54116 15285 54125
rect 15243 54076 15244 54116
rect 15284 54076 15285 54116
rect 15243 54067 15285 54076
rect 15627 54116 15669 54125
rect 18298 54116 18356 54117
rect 15627 54076 15628 54116
rect 15668 54076 15669 54116
rect 15627 54067 15669 54076
rect 16203 54107 16245 54116
rect 16203 54067 16204 54107
rect 16244 54067 16245 54107
rect 11499 54058 11541 54067
rect 14667 54058 14709 54067
rect 16203 54058 16245 54067
rect 16683 54107 16725 54116
rect 16683 54067 16684 54107
rect 16724 54067 16725 54107
rect 18298 54076 18307 54116
rect 18347 54076 18356 54116
rect 18298 54075 18356 54076
rect 18411 54116 18453 54125
rect 18411 54076 18412 54116
rect 18452 54076 18453 54116
rect 18411 54067 18453 54076
rect 18795 54116 18837 54125
rect 18795 54076 18796 54116
rect 18836 54076 18837 54116
rect 18795 54067 18837 54076
rect 19371 54107 19413 54116
rect 19371 54067 19372 54107
rect 19412 54067 19413 54107
rect 16683 54058 16725 54067
rect 19371 54058 19413 54067
rect 19851 54107 19893 54116
rect 19851 54067 19852 54107
rect 19892 54067 19893 54107
rect 19851 54058 19893 54067
rect 1419 54032 1461 54041
rect 1419 53992 1420 54032
rect 1460 53992 1461 54032
rect 1419 53983 1461 53992
rect 1707 54032 1749 54041
rect 1707 53992 1708 54032
rect 1748 53992 1749 54032
rect 1707 53983 1749 53992
rect 6795 54032 6837 54041
rect 6795 53992 6796 54032
rect 6836 53992 6837 54032
rect 6795 53983 6837 53992
rect 9963 54032 10005 54041
rect 9963 53992 9964 54032
rect 10004 53992 10005 54032
rect 9963 53983 10005 53992
rect 13131 54032 13173 54041
rect 13131 53992 13132 54032
rect 13172 53992 13173 54032
rect 13131 53983 13173 53992
rect 15723 54032 15765 54041
rect 15723 53992 15724 54032
rect 15764 53992 15765 54032
rect 15723 53983 15765 53992
rect 16906 54032 16964 54033
rect 16906 53992 16915 54032
rect 16955 53992 16964 54032
rect 16906 53991 16964 53992
rect 17259 54032 17301 54041
rect 17259 53992 17260 54032
rect 17300 53992 17301 54032
rect 17259 53983 17301 53992
rect 17451 54032 17493 54041
rect 17451 53992 17452 54032
rect 17492 53992 17493 54032
rect 17451 53983 17493 53992
rect 18027 54032 18069 54041
rect 18027 53992 18028 54032
rect 18068 53992 18069 54032
rect 18027 53983 18069 53992
rect 18891 54032 18933 54041
rect 18891 53992 18892 54032
rect 18932 53992 18933 54032
rect 18891 53983 18933 53992
rect 3531 53948 3573 53957
rect 3531 53908 3532 53948
rect 3572 53908 3573 53948
rect 3531 53899 3573 53908
rect 1179 53864 1221 53873
rect 1179 53824 1180 53864
rect 1220 53824 1221 53864
rect 1179 53815 1221 53824
rect 3706 53864 3764 53865
rect 3706 53824 3715 53864
rect 3755 53824 3764 53864
rect 3706 53823 3764 53824
rect 5931 53864 5973 53873
rect 5931 53824 5932 53864
rect 5972 53824 5973 53864
rect 5931 53815 5973 53824
rect 11146 53864 11204 53865
rect 11146 53824 11155 53864
rect 11195 53824 11204 53864
rect 11146 53823 11204 53824
rect 1152 53696 20448 53720
rect 1152 53656 3688 53696
rect 3728 53656 3770 53696
rect 3810 53656 3852 53696
rect 3892 53656 3934 53696
rect 3974 53656 4016 53696
rect 4056 53656 18808 53696
rect 18848 53656 18890 53696
rect 18930 53656 18972 53696
rect 19012 53656 19054 53696
rect 19094 53656 19136 53696
rect 19176 53656 20448 53696
rect 1152 53632 20448 53656
rect 2139 53528 2181 53537
rect 2139 53488 2140 53528
rect 2180 53488 2181 53528
rect 2139 53479 2181 53488
rect 8458 53528 8516 53529
rect 8458 53488 8467 53528
rect 8507 53488 8516 53528
rect 8458 53487 8516 53488
rect 10491 53528 10533 53537
rect 10491 53488 10492 53528
rect 10532 53488 10533 53528
rect 10491 53479 10533 53488
rect 12411 53528 12453 53537
rect 12411 53488 12412 53528
rect 12452 53488 12453 53528
rect 12411 53479 12453 53488
rect 15243 53528 15285 53537
rect 15243 53488 15244 53528
rect 15284 53488 15285 53528
rect 15243 53479 15285 53488
rect 17787 53528 17829 53537
rect 17787 53488 17788 53528
rect 17828 53488 17829 53528
rect 17787 53479 17829 53488
rect 10059 53444 10101 53453
rect 10059 53404 10060 53444
rect 10100 53404 10101 53444
rect 10059 53395 10101 53404
rect 12507 53444 12549 53453
rect 12507 53404 12508 53444
rect 12548 53404 12549 53444
rect 12507 53395 12549 53404
rect 17307 53444 17349 53453
rect 17307 53404 17308 53444
rect 17348 53404 17349 53444
rect 17307 53395 17349 53404
rect 1179 53360 1221 53369
rect 1179 53320 1180 53360
rect 1220 53320 1221 53360
rect 1179 53311 1221 53320
rect 1419 53360 1461 53369
rect 1419 53320 1420 53360
rect 1460 53320 1461 53360
rect 1419 53311 1461 53320
rect 1899 53360 1941 53369
rect 1899 53320 1900 53360
rect 1940 53320 1941 53360
rect 1899 53311 1941 53320
rect 3147 53360 3189 53369
rect 3147 53320 3148 53360
rect 3188 53320 3189 53360
rect 3147 53311 3189 53320
rect 7179 53360 7221 53369
rect 7179 53320 7180 53360
rect 7220 53320 7221 53360
rect 7179 53311 7221 53320
rect 10251 53360 10293 53369
rect 10251 53320 10252 53360
rect 10292 53320 10293 53360
rect 10251 53311 10293 53320
rect 10587 53360 10629 53369
rect 10587 53320 10588 53360
rect 10628 53320 10629 53360
rect 10587 53311 10629 53320
rect 12171 53360 12213 53369
rect 12171 53320 12172 53360
rect 12212 53320 12213 53360
rect 12171 53311 12213 53320
rect 12747 53360 12789 53369
rect 12747 53320 12748 53360
rect 12788 53320 12789 53360
rect 12747 53311 12789 53320
rect 16011 53360 16053 53369
rect 16011 53320 16012 53360
rect 16052 53320 16053 53360
rect 16011 53311 16053 53320
rect 17403 53360 17445 53369
rect 17403 53320 17404 53360
rect 17444 53320 17445 53360
rect 17403 53311 17445 53320
rect 17643 53360 17685 53369
rect 17643 53320 17644 53360
rect 17684 53320 17685 53360
rect 17643 53311 17685 53320
rect 18027 53360 18069 53369
rect 18027 53320 18028 53360
rect 18068 53320 18069 53360
rect 18027 53311 18069 53320
rect 18987 53360 19029 53369
rect 18987 53320 18988 53360
rect 19028 53320 19029 53360
rect 18987 53311 19029 53320
rect 2650 53276 2708 53277
rect 2650 53236 2659 53276
rect 2699 53236 2708 53276
rect 2650 53235 2708 53236
rect 2763 53276 2805 53285
rect 2763 53236 2764 53276
rect 2804 53236 2805 53276
rect 2763 53227 2805 53236
rect 3243 53276 3285 53285
rect 3243 53236 3244 53276
rect 3284 53236 3285 53276
rect 3243 53227 3285 53236
rect 3715 53276 3773 53277
rect 3715 53236 3724 53276
rect 3764 53236 3773 53276
rect 3715 53235 3773 53236
rect 4203 53276 4261 53277
rect 4203 53236 4212 53276
rect 4252 53236 4261 53276
rect 4203 53235 4261 53236
rect 4875 53276 4917 53285
rect 4875 53236 4876 53276
rect 4916 53236 4917 53276
rect 4875 53227 4917 53236
rect 6115 53276 6173 53277
rect 6115 53236 6124 53276
rect 6164 53236 6173 53276
rect 6115 53235 6173 53236
rect 6669 53276 6711 53285
rect 6669 53236 6670 53276
rect 6710 53236 6711 53276
rect 6669 53227 6711 53236
rect 6795 53276 6837 53285
rect 6795 53236 6796 53276
rect 6836 53236 6837 53276
rect 6795 53227 6837 53236
rect 7275 53276 7317 53285
rect 7275 53236 7276 53276
rect 7316 53236 7317 53276
rect 7275 53227 7317 53236
rect 7747 53276 7805 53277
rect 7747 53236 7756 53276
rect 7796 53236 7805 53276
rect 7747 53235 7805 53236
rect 8235 53276 8293 53277
rect 8235 53236 8244 53276
rect 8284 53236 8293 53276
rect 8235 53235 8293 53236
rect 8715 53276 8757 53285
rect 8715 53236 8716 53276
rect 8756 53236 8757 53276
rect 8715 53227 8757 53236
rect 9003 53276 9045 53285
rect 9003 53236 9004 53276
rect 9044 53236 9045 53276
rect 9003 53227 9045 53236
rect 9387 53276 9429 53285
rect 9387 53236 9388 53276
rect 9428 53236 9429 53276
rect 9387 53227 9429 53236
rect 9634 53276 9692 53277
rect 9634 53236 9643 53276
rect 9683 53236 9692 53276
rect 9634 53235 9692 53236
rect 9754 53276 9812 53277
rect 9754 53236 9763 53276
rect 9803 53236 9812 53276
rect 9754 53235 9812 53236
rect 10731 53276 10773 53285
rect 10731 53236 10732 53276
rect 10772 53236 10773 53276
rect 10731 53227 10773 53236
rect 13803 53276 13845 53285
rect 13803 53236 13804 53276
rect 13844 53236 13845 53276
rect 13803 53227 13845 53236
rect 15043 53276 15101 53277
rect 15043 53236 15052 53276
rect 15092 53236 15101 53276
rect 15043 53235 15101 53236
rect 15514 53276 15572 53277
rect 15514 53236 15523 53276
rect 15563 53236 15572 53276
rect 15514 53235 15572 53236
rect 15627 53276 15669 53285
rect 15627 53236 15628 53276
rect 15668 53236 15669 53276
rect 15627 53227 15669 53236
rect 16107 53276 16149 53285
rect 16107 53236 16108 53276
rect 16148 53236 16149 53276
rect 16107 53227 16149 53236
rect 16579 53276 16637 53277
rect 16579 53236 16588 53276
rect 16628 53236 16637 53276
rect 16579 53235 16637 53236
rect 17098 53276 17156 53277
rect 17098 53236 17107 53276
rect 17147 53236 17156 53276
rect 17098 53235 17156 53236
rect 18490 53276 18548 53277
rect 18490 53236 18499 53276
rect 18539 53236 18548 53276
rect 18490 53235 18548 53236
rect 18603 53276 18645 53285
rect 18603 53236 18604 53276
rect 18644 53236 18645 53276
rect 18603 53227 18645 53236
rect 19083 53276 19125 53285
rect 19083 53236 19084 53276
rect 19124 53236 19125 53276
rect 19083 53227 19125 53236
rect 19555 53276 19613 53277
rect 19555 53236 19564 53276
rect 19604 53236 19613 53276
rect 19555 53235 19613 53236
rect 20043 53276 20101 53277
rect 20043 53236 20052 53276
rect 20092 53236 20101 53276
rect 20043 53235 20101 53236
rect 4395 53108 4437 53117
rect 4395 53068 4396 53108
rect 4436 53068 4437 53108
rect 4395 53059 4437 53068
rect 6315 53108 6357 53117
rect 6315 53068 6316 53108
rect 6356 53068 6357 53108
rect 6315 53059 6357 53068
rect 8794 53108 8852 53109
rect 8794 53068 8803 53108
rect 8843 53068 8852 53108
rect 8794 53067 8852 53068
rect 20235 53108 20277 53117
rect 20235 53068 20236 53108
rect 20276 53068 20277 53108
rect 20235 53059 20277 53068
rect 1152 52940 20452 52964
rect 1152 52900 4928 52940
rect 4968 52900 5010 52940
rect 5050 52900 5092 52940
rect 5132 52900 5174 52940
rect 5214 52900 5256 52940
rect 5296 52900 20048 52940
rect 20088 52900 20130 52940
rect 20170 52900 20212 52940
rect 20252 52900 20294 52940
rect 20334 52900 20376 52940
rect 20416 52900 20452 52940
rect 1152 52876 20452 52900
rect 2667 52772 2709 52781
rect 2667 52732 2668 52772
rect 2708 52732 2709 52772
rect 2667 52723 2709 52732
rect 9867 52772 9909 52781
rect 9867 52732 9868 52772
rect 9908 52732 9909 52772
rect 9867 52723 9909 52732
rect 10635 52772 10677 52781
rect 10635 52732 10636 52772
rect 10676 52732 10677 52772
rect 10635 52723 10677 52732
rect 10923 52772 10965 52781
rect 10923 52732 10924 52772
rect 10964 52732 10965 52772
rect 10923 52723 10965 52732
rect 12555 52772 12597 52781
rect 12555 52732 12556 52772
rect 12596 52732 12597 52772
rect 12555 52723 12597 52732
rect 15627 52772 15669 52781
rect 15627 52732 15628 52772
rect 15668 52732 15669 52772
rect 15627 52723 15669 52732
rect 17259 52772 17301 52781
rect 17259 52732 17260 52772
rect 17300 52732 17301 52772
rect 17259 52723 17301 52732
rect 18891 52772 18933 52781
rect 18891 52732 18892 52772
rect 18932 52732 18933 52772
rect 18891 52723 18933 52732
rect 19035 52772 19077 52781
rect 19035 52732 19036 52772
rect 19076 52732 19077 52772
rect 19035 52723 19077 52732
rect 5067 52688 5109 52697
rect 5067 52648 5068 52688
rect 5108 52648 5109 52688
rect 5067 52639 5109 52648
rect 19419 52688 19461 52697
rect 19419 52648 19420 52688
rect 19460 52648 19461 52688
rect 19419 52639 19461 52648
rect 1227 52604 1269 52613
rect 3627 52604 3669 52613
rect 5338 52604 5396 52605
rect 1227 52564 1228 52604
rect 1268 52564 1269 52604
rect 1227 52555 1269 52564
rect 2475 52595 2517 52604
rect 2475 52555 2476 52595
rect 2516 52555 2517 52595
rect 3627 52564 3628 52604
rect 3668 52564 3669 52604
rect 3627 52555 3669 52564
rect 4875 52595 4917 52604
rect 4875 52555 4876 52595
rect 4916 52555 4917 52595
rect 5338 52564 5347 52604
rect 5387 52564 5396 52604
rect 5338 52563 5396 52564
rect 5451 52604 5493 52613
rect 5451 52564 5452 52604
rect 5492 52564 5493 52604
rect 5451 52555 5493 52564
rect 5835 52604 5877 52613
rect 8122 52604 8180 52605
rect 5835 52564 5836 52604
rect 5876 52564 5877 52604
rect 5835 52555 5877 52564
rect 6411 52595 6453 52604
rect 6411 52555 6412 52595
rect 6452 52555 6453 52595
rect 2475 52546 2517 52555
rect 4875 52546 4917 52555
rect 6411 52546 6453 52555
rect 6891 52595 6933 52604
rect 6891 52555 6892 52595
rect 6932 52555 6933 52595
rect 8122 52564 8131 52604
rect 8171 52564 8180 52604
rect 8122 52563 8180 52564
rect 8235 52604 8277 52613
rect 8235 52564 8236 52604
rect 8276 52564 8277 52604
rect 8235 52555 8277 52564
rect 8619 52604 8661 52613
rect 10006 52604 10048 52613
rect 8619 52564 8620 52604
rect 8660 52564 8661 52604
rect 8619 52555 8661 52564
rect 9195 52595 9237 52604
rect 9195 52555 9196 52595
rect 9236 52555 9237 52595
rect 6891 52546 6933 52555
rect 9195 52546 9237 52555
rect 9675 52595 9717 52604
rect 9675 52555 9676 52595
rect 9716 52555 9717 52595
rect 10006 52564 10007 52604
rect 10047 52564 10048 52604
rect 10006 52555 10048 52564
rect 10251 52604 10293 52613
rect 10251 52564 10252 52604
rect 10292 52564 10293 52604
rect 10251 52555 10293 52564
rect 10539 52604 10581 52613
rect 10539 52564 10540 52604
rect 10580 52564 10581 52604
rect 10539 52555 10581 52564
rect 10714 52604 10772 52605
rect 12363 52604 12405 52613
rect 13995 52604 14037 52613
rect 10714 52564 10723 52604
rect 10763 52564 10772 52604
rect 10714 52563 10772 52564
rect 11115 52595 11157 52604
rect 11115 52555 11116 52595
rect 11156 52555 11157 52595
rect 12363 52564 12364 52604
rect 12404 52564 12405 52604
rect 12363 52555 12405 52564
rect 12747 52595 12789 52604
rect 12747 52555 12748 52595
rect 12788 52555 12789 52595
rect 13995 52564 13996 52604
rect 14036 52564 14037 52604
rect 13995 52555 14037 52564
rect 14187 52604 14229 52613
rect 15819 52604 15861 52613
rect 17451 52604 17493 52613
rect 14187 52564 14188 52604
rect 14228 52564 14229 52604
rect 14187 52555 14229 52564
rect 15435 52595 15477 52604
rect 15435 52555 15436 52595
rect 15476 52555 15477 52595
rect 15819 52564 15820 52604
rect 15860 52564 15861 52604
rect 15819 52555 15861 52564
rect 17067 52595 17109 52604
rect 17067 52555 17068 52595
rect 17108 52555 17109 52595
rect 17451 52564 17452 52604
rect 17492 52564 17493 52604
rect 17451 52555 17493 52564
rect 18699 52595 18741 52604
rect 18699 52555 18700 52595
rect 18740 52555 18741 52595
rect 9675 52546 9717 52555
rect 11115 52546 11157 52555
rect 12747 52546 12789 52555
rect 15435 52546 15477 52555
rect 17067 52546 17109 52555
rect 18699 52546 18741 52555
rect 3051 52520 3093 52529
rect 3051 52480 3052 52520
rect 3092 52480 3093 52520
rect 3051 52471 3093 52480
rect 5931 52520 5973 52529
rect 5931 52480 5932 52520
rect 5972 52480 5973 52520
rect 5931 52471 5973 52480
rect 8715 52520 8757 52529
rect 8715 52480 8716 52520
rect 8756 52480 8757 52520
rect 8715 52471 8757 52480
rect 10138 52520 10196 52521
rect 10138 52480 10147 52520
rect 10187 52480 10196 52520
rect 10138 52479 10196 52480
rect 10347 52520 10389 52529
rect 10347 52480 10348 52520
rect 10388 52480 10389 52520
rect 10347 52471 10389 52480
rect 19275 52520 19317 52529
rect 19275 52480 19276 52520
rect 19316 52480 19317 52520
rect 19275 52471 19317 52480
rect 19659 52520 19701 52529
rect 19659 52480 19660 52520
rect 19700 52480 19701 52520
rect 19659 52471 19701 52480
rect 20139 52520 20181 52529
rect 20139 52480 20140 52520
rect 20180 52480 20181 52520
rect 20139 52471 20181 52480
rect 2811 52352 2853 52361
rect 2811 52312 2812 52352
rect 2852 52312 2853 52352
rect 2811 52303 2853 52312
rect 7114 52352 7172 52353
rect 7114 52312 7123 52352
rect 7163 52312 7172 52352
rect 7114 52311 7172 52312
rect 20379 52352 20421 52361
rect 20379 52312 20380 52352
rect 20420 52312 20421 52352
rect 20379 52303 20421 52312
rect 1152 52184 20448 52208
rect 1152 52144 3688 52184
rect 3728 52144 3770 52184
rect 3810 52144 3852 52184
rect 3892 52144 3934 52184
rect 3974 52144 4016 52184
rect 4056 52144 18808 52184
rect 18848 52144 18890 52184
rect 18930 52144 18972 52184
rect 19012 52144 19054 52184
rect 19094 52144 19136 52184
rect 19176 52144 20448 52184
rect 1152 52120 20448 52144
rect 7851 52016 7893 52025
rect 7851 51976 7852 52016
rect 7892 51976 7893 52016
rect 7851 51967 7893 51976
rect 10347 52016 10389 52025
rect 10347 51976 10348 52016
rect 10388 51976 10389 52016
rect 10347 51967 10389 51976
rect 10539 52016 10581 52025
rect 10539 51976 10540 52016
rect 10580 51976 10581 52016
rect 10539 51967 10581 51976
rect 10923 52016 10965 52025
rect 10923 51976 10924 52016
rect 10964 51976 10965 52016
rect 10923 51967 10965 51976
rect 1419 51848 1461 51857
rect 1419 51808 1420 51848
rect 1460 51808 1461 51848
rect 1419 51799 1461 51808
rect 1803 51848 1845 51857
rect 1803 51808 1804 51848
rect 1844 51808 1845 51848
rect 1803 51799 1845 51808
rect 2091 51848 2133 51857
rect 2091 51808 2092 51848
rect 2132 51808 2133 51848
rect 2091 51799 2133 51808
rect 2475 51848 2517 51857
rect 2475 51808 2476 51848
rect 2516 51808 2517 51848
rect 2475 51799 2517 51808
rect 2715 51848 2757 51857
rect 2715 51808 2716 51848
rect 2756 51808 2757 51848
rect 2715 51799 2757 51808
rect 4011 51848 4053 51857
rect 4011 51808 4012 51848
rect 4052 51808 4053 51848
rect 4011 51799 4053 51808
rect 5067 51848 5109 51857
rect 5067 51808 5068 51848
rect 5108 51808 5109 51848
rect 5067 51799 5109 51808
rect 6411 51848 6453 51857
rect 6411 51808 6412 51848
rect 6452 51808 6453 51848
rect 6411 51799 6453 51808
rect 9867 51848 9909 51857
rect 9867 51808 9868 51848
rect 9908 51808 9909 51848
rect 9867 51799 9909 51808
rect 12555 51848 12597 51857
rect 12555 51808 12556 51848
rect 12596 51808 12597 51848
rect 12555 51799 12597 51808
rect 20139 51848 20181 51857
rect 20139 51808 20140 51848
rect 20180 51808 20181 51848
rect 20139 51799 20181 51808
rect 3034 51764 3092 51765
rect 3034 51724 3043 51764
rect 3083 51724 3092 51764
rect 3034 51723 3092 51724
rect 3523 51764 3581 51765
rect 3523 51724 3532 51764
rect 3572 51724 3581 51764
rect 3523 51723 3581 51724
rect 4107 51764 4149 51773
rect 4107 51724 4108 51764
rect 4148 51724 4149 51764
rect 4107 51715 4149 51724
rect 4491 51764 4533 51773
rect 4491 51724 4492 51764
rect 4532 51724 4533 51764
rect 4491 51715 4533 51724
rect 4601 51764 4659 51765
rect 4601 51724 4610 51764
rect 4650 51724 4659 51764
rect 4601 51723 4659 51724
rect 5914 51764 5972 51765
rect 5914 51724 5923 51764
rect 5963 51724 5972 51764
rect 5914 51723 5972 51724
rect 6027 51764 6069 51773
rect 6027 51724 6028 51764
rect 6068 51724 6069 51764
rect 6027 51715 6069 51724
rect 6507 51764 6549 51773
rect 6507 51724 6508 51764
rect 6548 51724 6549 51764
rect 6507 51715 6549 51724
rect 6979 51764 7037 51765
rect 6979 51724 6988 51764
rect 7028 51724 7037 51764
rect 6979 51723 7037 51724
rect 7471 51764 7529 51765
rect 7471 51724 7480 51764
rect 7520 51724 7529 51764
rect 7471 51723 7529 51724
rect 8035 51764 8093 51765
rect 8035 51724 8044 51764
rect 8084 51724 8093 51764
rect 8035 51723 8093 51724
rect 9291 51764 9333 51773
rect 9291 51724 9292 51764
rect 9332 51724 9333 51764
rect 9291 51715 9333 51724
rect 9526 51764 9568 51773
rect 9526 51724 9527 51764
rect 9567 51724 9568 51764
rect 9526 51715 9568 51724
rect 9658 51764 9716 51765
rect 9658 51724 9667 51764
rect 9707 51724 9716 51764
rect 9658 51723 9716 51724
rect 9771 51764 9813 51773
rect 9771 51724 9772 51764
rect 9812 51724 9813 51764
rect 9771 51715 9813 51724
rect 10042 51764 10100 51765
rect 10042 51724 10051 51764
rect 10091 51724 10100 51764
rect 10042 51723 10100 51724
rect 10358 51764 10400 51773
rect 10358 51724 10359 51764
rect 10399 51724 10400 51764
rect 10358 51715 10400 51724
rect 10539 51764 10581 51773
rect 10539 51724 10540 51764
rect 10580 51724 10581 51764
rect 10539 51715 10581 51724
rect 10720 51764 10778 51765
rect 10720 51724 10729 51764
rect 10769 51724 10778 51764
rect 10720 51723 10778 51724
rect 11107 51764 11165 51765
rect 11107 51724 11116 51764
rect 11156 51724 11165 51764
rect 11107 51723 11165 51724
rect 12363 51764 12405 51773
rect 12363 51724 12364 51764
rect 12404 51724 12405 51764
rect 12363 51715 12405 51724
rect 13411 51764 13469 51765
rect 13411 51724 13420 51764
rect 13460 51724 13469 51764
rect 13411 51723 13469 51724
rect 14667 51764 14709 51773
rect 14667 51724 14668 51764
rect 14708 51724 14709 51764
rect 14667 51715 14709 51724
rect 14859 51764 14901 51773
rect 14859 51724 14860 51764
rect 14900 51724 14901 51764
rect 14859 51715 14901 51724
rect 16099 51764 16157 51765
rect 16099 51724 16108 51764
rect 16148 51724 16157 51764
rect 16099 51723 16157 51724
rect 16675 51764 16733 51765
rect 16675 51724 16684 51764
rect 16724 51724 16733 51764
rect 16675 51723 16733 51724
rect 17931 51764 17973 51773
rect 17931 51724 17932 51764
rect 17972 51724 17973 51764
rect 17931 51715 17973 51724
rect 18219 51764 18261 51773
rect 18219 51724 18220 51764
rect 18260 51724 18261 51764
rect 18219 51715 18261 51724
rect 19459 51764 19517 51765
rect 19459 51724 19468 51764
rect 19508 51724 19517 51764
rect 19459 51723 19517 51724
rect 2331 51680 2373 51689
rect 2331 51640 2332 51680
rect 2372 51640 2373 51680
rect 2331 51631 2373 51640
rect 4827 51680 4869 51689
rect 4827 51640 4828 51680
rect 4868 51640 4869 51680
rect 4827 51631 4869 51640
rect 10155 51680 10197 51689
rect 10155 51640 10156 51680
rect 10196 51640 10197 51680
rect 10155 51631 10197 51640
rect 10923 51680 10965 51689
rect 10923 51640 10924 51680
rect 10964 51640 10965 51680
rect 10923 51631 10965 51640
rect 12795 51680 12837 51689
rect 12795 51640 12796 51680
rect 12836 51640 12837 51680
rect 12795 51631 12837 51640
rect 1179 51596 1221 51605
rect 1179 51556 1180 51596
rect 1220 51556 1221 51596
rect 1179 51547 1221 51556
rect 1563 51596 1605 51605
rect 1563 51556 1564 51596
rect 1604 51556 1605 51596
rect 1563 51547 1605 51556
rect 2859 51596 2901 51605
rect 2859 51556 2860 51596
rect 2900 51556 2901 51596
rect 2859 51547 2901 51556
rect 7659 51596 7701 51605
rect 7659 51556 7660 51596
rect 7700 51556 7701 51596
rect 7659 51547 7701 51556
rect 13227 51596 13269 51605
rect 13227 51556 13228 51596
rect 13268 51556 13269 51596
rect 13227 51547 13269 51556
rect 16299 51596 16341 51605
rect 16299 51556 16300 51596
rect 16340 51556 16341 51596
rect 16299 51547 16341 51556
rect 16491 51596 16533 51605
rect 16491 51556 16492 51596
rect 16532 51556 16533 51596
rect 16491 51547 16533 51556
rect 19659 51596 19701 51605
rect 19659 51556 19660 51596
rect 19700 51556 19701 51596
rect 19659 51547 19701 51556
rect 20379 51596 20421 51605
rect 20379 51556 20380 51596
rect 20420 51556 20421 51596
rect 20379 51547 20421 51556
rect 1152 51428 20452 51452
rect 1152 51388 4928 51428
rect 4968 51388 5010 51428
rect 5050 51388 5092 51428
rect 5132 51388 5174 51428
rect 5214 51388 5256 51428
rect 5296 51388 20048 51428
rect 20088 51388 20130 51428
rect 20170 51388 20212 51428
rect 20252 51388 20294 51428
rect 20334 51388 20376 51428
rect 20416 51388 20452 51428
rect 1152 51364 20452 51388
rect 1179 51260 1221 51269
rect 1179 51220 1180 51260
rect 1220 51220 1221 51260
rect 1179 51211 1221 51220
rect 1563 51260 1605 51269
rect 1563 51220 1564 51260
rect 1604 51220 1605 51260
rect 1563 51211 1605 51220
rect 5931 51260 5973 51269
rect 5931 51220 5932 51260
rect 5972 51220 5973 51260
rect 5931 51211 5973 51220
rect 7563 51260 7605 51269
rect 7563 51220 7564 51260
rect 7604 51220 7605 51260
rect 7563 51211 7605 51220
rect 12123 51260 12165 51269
rect 12123 51220 12124 51260
rect 12164 51220 12165 51260
rect 12123 51211 12165 51220
rect 17451 51260 17493 51269
rect 17451 51220 17452 51260
rect 17492 51220 17493 51260
rect 17451 51211 17493 51220
rect 19611 51260 19653 51269
rect 19611 51220 19612 51260
rect 19652 51220 19653 51260
rect 19611 51211 19653 51220
rect 13323 51176 13365 51185
rect 13323 51136 13324 51176
rect 13364 51136 13365 51176
rect 13323 51127 13365 51136
rect 4491 51092 4533 51101
rect 6123 51092 6165 51101
rect 8907 51092 8949 51101
rect 10539 51092 10581 51101
rect 14763 51092 14805 51101
rect 4491 51052 4492 51092
rect 4532 51052 4533 51092
rect 4491 51043 4533 51052
rect 5739 51083 5781 51092
rect 5739 51043 5740 51083
rect 5780 51043 5781 51083
rect 6123 51052 6124 51092
rect 6164 51052 6165 51092
rect 6123 51043 6165 51052
rect 7371 51083 7413 51092
rect 7371 51043 7372 51083
rect 7412 51043 7413 51083
rect 8907 51052 8908 51092
rect 8948 51052 8949 51092
rect 8907 51043 8949 51052
rect 10155 51083 10197 51092
rect 10155 51043 10156 51083
rect 10196 51043 10197 51083
rect 10539 51052 10540 51092
rect 10580 51052 10581 51092
rect 10539 51043 10581 51052
rect 11787 51083 11829 51092
rect 11787 51043 11788 51083
rect 11828 51043 11829 51083
rect 5739 51034 5781 51043
rect 7371 51034 7413 51043
rect 10155 51034 10197 51043
rect 11787 51034 11829 51043
rect 13515 51083 13557 51092
rect 13515 51043 13516 51083
rect 13556 51043 13557 51083
rect 14763 51052 14764 51092
rect 14804 51052 14805 51092
rect 14763 51043 14805 51052
rect 15706 51092 15764 51093
rect 15706 51052 15715 51092
rect 15755 51052 15764 51092
rect 15706 51051 15764 51052
rect 15819 51092 15861 51101
rect 15819 51052 15820 51092
rect 15860 51052 15861 51092
rect 15819 51043 15861 51052
rect 16203 51092 16245 51101
rect 17643 51092 17685 51101
rect 16203 51052 16204 51092
rect 16244 51052 16245 51092
rect 16203 51043 16245 51052
rect 16779 51083 16821 51092
rect 16779 51043 16780 51083
rect 16820 51043 16821 51083
rect 13515 51034 13557 51043
rect 16779 51034 16821 51043
rect 17259 51083 17301 51092
rect 17259 51043 17260 51083
rect 17300 51043 17301 51083
rect 17643 51052 17644 51092
rect 17684 51052 17685 51092
rect 17643 51043 17685 51052
rect 18891 51083 18933 51092
rect 18891 51043 18892 51083
rect 18932 51043 18933 51083
rect 17259 51034 17301 51043
rect 18891 51034 18933 51043
rect 1419 51008 1461 51017
rect 1419 50968 1420 51008
rect 1460 50968 1461 51008
rect 1419 50959 1461 50968
rect 1803 51008 1845 51017
rect 1803 50968 1804 51008
rect 1844 50968 1845 51008
rect 1803 50959 1845 50968
rect 2763 51008 2805 51017
rect 2763 50968 2764 51008
rect 2804 50968 2805 51008
rect 2763 50959 2805 50968
rect 12363 51008 12405 51017
rect 12363 50968 12364 51008
rect 12404 50968 12405 51008
rect 12363 50959 12405 50968
rect 16299 51008 16341 51017
rect 16299 50968 16300 51008
rect 16340 50968 16341 51008
rect 16299 50959 16341 50968
rect 19371 51008 19413 51017
rect 19371 50968 19372 51008
rect 19412 50968 19413 51008
rect 19371 50959 19413 50968
rect 19755 51008 19797 51017
rect 19755 50968 19756 51008
rect 19796 50968 19797 51008
rect 19755 50959 19797 50968
rect 20139 51008 20181 51017
rect 20139 50968 20140 51008
rect 20180 50968 20181 51008
rect 20139 50959 20181 50968
rect 19995 50924 20037 50933
rect 19995 50884 19996 50924
rect 20036 50884 20037 50924
rect 19995 50875 20037 50884
rect 2523 50840 2565 50849
rect 2523 50800 2524 50840
rect 2564 50800 2565 50840
rect 2523 50791 2565 50800
rect 10347 50840 10389 50849
rect 10347 50800 10348 50840
rect 10388 50800 10389 50840
rect 10347 50791 10389 50800
rect 11979 50840 12021 50849
rect 11979 50800 11980 50840
rect 12020 50800 12021 50840
rect 11979 50791 12021 50800
rect 19083 50840 19125 50849
rect 19083 50800 19084 50840
rect 19124 50800 19125 50840
rect 19083 50791 19125 50800
rect 20379 50840 20421 50849
rect 20379 50800 20380 50840
rect 20420 50800 20421 50840
rect 20379 50791 20421 50800
rect 1152 50672 20448 50696
rect 1152 50632 3688 50672
rect 3728 50632 3770 50672
rect 3810 50632 3852 50672
rect 3892 50632 3934 50672
rect 3974 50632 4016 50672
rect 4056 50632 18808 50672
rect 18848 50632 18890 50672
rect 18930 50632 18972 50672
rect 19012 50632 19054 50672
rect 19094 50632 19136 50672
rect 19176 50632 20448 50672
rect 1152 50608 20448 50632
rect 8907 50420 8949 50429
rect 8907 50380 8908 50420
rect 8948 50380 8949 50420
rect 8907 50371 8949 50380
rect 11931 50420 11973 50429
rect 11931 50380 11932 50420
rect 11972 50380 11973 50420
rect 11931 50371 11973 50380
rect 18459 50420 18501 50429
rect 18459 50380 18460 50420
rect 18500 50380 18501 50420
rect 18459 50371 18501 50380
rect 9675 50336 9717 50345
rect 9675 50296 9676 50336
rect 9716 50296 9717 50336
rect 9675 50287 9717 50296
rect 11403 50336 11445 50345
rect 11403 50296 11404 50336
rect 11444 50296 11445 50336
rect 11403 50287 11445 50296
rect 11691 50336 11733 50345
rect 11691 50296 11692 50336
rect 11732 50296 11733 50336
rect 11691 50287 11733 50296
rect 12267 50336 12309 50345
rect 12267 50296 12268 50336
rect 12308 50296 12309 50336
rect 12267 50287 12309 50296
rect 16395 50336 16437 50345
rect 16395 50296 16396 50336
rect 16436 50296 16437 50336
rect 16395 50287 16437 50296
rect 19659 50336 19701 50345
rect 19659 50296 19660 50336
rect 19700 50296 19701 50336
rect 19659 50287 19701 50296
rect 2091 50252 2133 50261
rect 2091 50212 2092 50252
rect 2132 50212 2133 50252
rect 2091 50203 2133 50212
rect 3331 50252 3389 50253
rect 3331 50212 3340 50252
rect 3380 50212 3389 50252
rect 3331 50211 3389 50212
rect 4011 50252 4053 50261
rect 4011 50212 4012 50252
rect 4052 50212 4053 50252
rect 4011 50203 4053 50212
rect 5251 50252 5309 50253
rect 5251 50212 5260 50252
rect 5300 50212 5309 50252
rect 5251 50211 5309 50212
rect 7467 50252 7509 50261
rect 7467 50212 7468 50252
rect 7508 50212 7509 50252
rect 7467 50203 7509 50212
rect 8707 50252 8765 50253
rect 8707 50212 8716 50252
rect 8756 50212 8765 50252
rect 8707 50211 8765 50212
rect 9178 50252 9236 50253
rect 9178 50212 9187 50252
rect 9227 50212 9236 50252
rect 9178 50211 9236 50212
rect 9291 50252 9333 50261
rect 9291 50212 9292 50252
rect 9332 50212 9333 50252
rect 9291 50203 9333 50212
rect 9771 50252 9813 50261
rect 9771 50212 9772 50252
rect 9812 50212 9813 50252
rect 9771 50203 9813 50212
rect 10243 50252 10301 50253
rect 10243 50212 10252 50252
rect 10292 50212 10301 50252
rect 10243 50211 10301 50212
rect 10731 50252 10789 50253
rect 10731 50212 10740 50252
rect 10780 50212 10789 50252
rect 10731 50211 10789 50212
rect 12555 50252 12597 50261
rect 12555 50212 12556 50252
rect 12596 50212 12597 50252
rect 12555 50203 12597 50212
rect 13795 50252 13853 50253
rect 13795 50212 13804 50252
rect 13844 50212 13853 50252
rect 13795 50211 13853 50212
rect 14187 50252 14229 50261
rect 14187 50212 14188 50252
rect 14228 50212 14229 50252
rect 14187 50203 14229 50212
rect 15427 50252 15485 50253
rect 15427 50212 15436 50252
rect 15476 50212 15485 50252
rect 15427 50211 15485 50212
rect 15898 50252 15956 50253
rect 15898 50212 15907 50252
rect 15947 50212 15956 50252
rect 15898 50211 15956 50212
rect 16011 50252 16053 50261
rect 16011 50212 16012 50252
rect 16052 50212 16053 50252
rect 16011 50203 16053 50212
rect 16491 50252 16533 50261
rect 16491 50212 16492 50252
rect 16532 50212 16533 50252
rect 16491 50203 16533 50212
rect 16963 50252 17021 50253
rect 16963 50212 16972 50252
rect 17012 50212 17021 50252
rect 16963 50211 17021 50212
rect 17451 50252 17509 50253
rect 17451 50212 17460 50252
rect 17500 50212 17509 50252
rect 17451 50211 17509 50212
rect 18682 50252 18740 50253
rect 18682 50212 18691 50252
rect 18731 50212 18740 50252
rect 18682 50211 18740 50212
rect 19171 50252 19229 50253
rect 19171 50212 19180 50252
rect 19220 50212 19229 50252
rect 19171 50211 19229 50212
rect 19755 50252 19797 50261
rect 19755 50212 19756 50252
rect 19796 50212 19797 50252
rect 19755 50203 19797 50212
rect 20139 50252 20181 50261
rect 20139 50212 20140 50252
rect 20180 50212 20181 50252
rect 20139 50203 20181 50212
rect 20240 50252 20282 50261
rect 20240 50212 20241 50252
rect 20281 50212 20282 50252
rect 20240 50203 20282 50212
rect 3531 50084 3573 50093
rect 3531 50044 3532 50084
rect 3572 50044 3573 50084
rect 3531 50035 3573 50044
rect 5451 50084 5493 50093
rect 5451 50044 5452 50084
rect 5492 50044 5493 50084
rect 5451 50035 5493 50044
rect 10923 50084 10965 50093
rect 10923 50044 10924 50084
rect 10964 50044 10965 50084
rect 10923 50035 10965 50044
rect 11163 50084 11205 50093
rect 11163 50044 11164 50084
rect 11204 50044 11205 50084
rect 11163 50035 11205 50044
rect 12027 50084 12069 50093
rect 12027 50044 12028 50084
rect 12068 50044 12069 50084
rect 12027 50035 12069 50044
rect 13995 50084 14037 50093
rect 13995 50044 13996 50084
rect 14036 50044 14037 50084
rect 13995 50035 14037 50044
rect 15627 50084 15669 50093
rect 15627 50044 15628 50084
rect 15668 50044 15669 50084
rect 15627 50035 15669 50044
rect 17643 50084 17685 50093
rect 17643 50044 17644 50084
rect 17684 50044 17685 50084
rect 17643 50035 17685 50044
rect 1152 49916 20452 49940
rect 1152 49876 4928 49916
rect 4968 49876 5010 49916
rect 5050 49876 5092 49916
rect 5132 49876 5174 49916
rect 5214 49876 5256 49916
rect 5296 49876 20048 49916
rect 20088 49876 20130 49916
rect 20170 49876 20212 49916
rect 20252 49876 20294 49916
rect 20334 49876 20376 49916
rect 20416 49876 20452 49916
rect 1152 49852 20452 49876
rect 9195 49748 9237 49757
rect 9195 49708 9196 49748
rect 9236 49708 9237 49748
rect 9195 49699 9237 49708
rect 11403 49748 11445 49757
rect 11403 49708 11404 49748
rect 11444 49708 11445 49748
rect 11403 49699 11445 49708
rect 15819 49748 15861 49757
rect 15819 49708 15820 49748
rect 15860 49708 15861 49748
rect 15819 49699 15861 49708
rect 17451 49748 17493 49757
rect 17451 49708 17452 49748
rect 17492 49708 17493 49748
rect 17451 49699 17493 49708
rect 20379 49748 20421 49757
rect 20379 49708 20380 49748
rect 20420 49708 20421 49748
rect 20379 49699 20421 49708
rect 11835 49664 11877 49673
rect 11835 49624 11836 49664
rect 11876 49624 11877 49664
rect 11835 49615 11877 49624
rect 1995 49580 2037 49589
rect 5451 49580 5493 49589
rect 7563 49580 7605 49589
rect 1995 49540 1996 49580
rect 2036 49540 2037 49580
rect 1995 49531 2037 49540
rect 3243 49571 3285 49580
rect 3243 49531 3244 49571
rect 3284 49531 3285 49571
rect 3243 49522 3285 49531
rect 4203 49571 4245 49580
rect 4203 49531 4204 49571
rect 4244 49531 4245 49571
rect 5451 49540 5452 49580
rect 5492 49540 5493 49580
rect 5451 49531 5493 49540
rect 6315 49571 6357 49580
rect 6315 49531 6316 49571
rect 6356 49531 6357 49571
rect 7563 49540 7564 49580
rect 7604 49540 7605 49580
rect 7563 49531 7605 49540
rect 7755 49580 7797 49589
rect 9658 49580 9716 49581
rect 7755 49540 7756 49580
rect 7796 49540 7797 49580
rect 7755 49531 7797 49540
rect 9003 49571 9045 49580
rect 9003 49531 9004 49571
rect 9044 49531 9045 49571
rect 9658 49540 9667 49580
rect 9707 49540 9716 49580
rect 9658 49539 9716 49540
rect 9771 49580 9813 49589
rect 9771 49540 9772 49580
rect 9812 49540 9813 49580
rect 9771 49531 9813 49540
rect 10155 49580 10197 49589
rect 11979 49580 12021 49589
rect 14379 49580 14421 49589
rect 16011 49580 16053 49589
rect 10155 49540 10156 49580
rect 10196 49540 10197 49580
rect 10155 49531 10197 49540
rect 10731 49571 10773 49580
rect 10731 49531 10732 49571
rect 10772 49531 10773 49571
rect 4203 49522 4245 49531
rect 6315 49522 6357 49531
rect 9003 49522 9045 49531
rect 10731 49522 10773 49531
rect 11211 49571 11253 49580
rect 11211 49531 11212 49571
rect 11252 49531 11253 49571
rect 11979 49540 11980 49580
rect 12020 49540 12021 49580
rect 11979 49531 12021 49540
rect 13227 49571 13269 49580
rect 13227 49531 13228 49571
rect 13268 49531 13269 49571
rect 14379 49540 14380 49580
rect 14420 49540 14421 49580
rect 14379 49531 14421 49540
rect 15627 49571 15669 49580
rect 15627 49531 15628 49571
rect 15668 49531 15669 49571
rect 16011 49540 16012 49580
rect 16052 49540 16053 49580
rect 16011 49531 16053 49540
rect 17259 49571 17301 49580
rect 17259 49531 17260 49571
rect 17300 49531 17301 49571
rect 11211 49522 11253 49531
rect 13227 49522 13269 49531
rect 15627 49522 15669 49531
rect 17259 49522 17301 49531
rect 10251 49496 10293 49505
rect 10251 49456 10252 49496
rect 10292 49456 10293 49496
rect 10251 49447 10293 49456
rect 11595 49496 11637 49505
rect 11595 49456 11596 49496
rect 11636 49456 11637 49496
rect 11595 49447 11637 49456
rect 17835 49496 17877 49505
rect 17835 49456 17836 49496
rect 17876 49456 17877 49496
rect 17835 49447 17877 49456
rect 19371 49496 19413 49505
rect 19371 49456 19372 49496
rect 19412 49456 19413 49496
rect 19371 49447 19413 49456
rect 19755 49496 19797 49505
rect 19755 49456 19756 49496
rect 19796 49456 19797 49496
rect 19755 49447 19797 49456
rect 20139 49496 20181 49505
rect 20139 49456 20140 49496
rect 20180 49456 20181 49496
rect 20139 49447 20181 49456
rect 3435 49412 3477 49421
rect 3435 49372 3436 49412
rect 3476 49372 3477 49412
rect 3435 49363 3477 49372
rect 19995 49412 20037 49421
rect 19995 49372 19996 49412
rect 20036 49372 20037 49412
rect 19995 49363 20037 49372
rect 4011 49328 4053 49337
rect 4011 49288 4012 49328
rect 4052 49288 4053 49328
rect 4011 49279 4053 49288
rect 6123 49328 6165 49337
rect 6123 49288 6124 49328
rect 6164 49288 6165 49328
rect 6123 49279 6165 49288
rect 13419 49328 13461 49337
rect 13419 49288 13420 49328
rect 13460 49288 13461 49328
rect 13419 49279 13461 49288
rect 17595 49328 17637 49337
rect 17595 49288 17596 49328
rect 17636 49288 17637 49328
rect 17595 49279 17637 49288
rect 19611 49328 19653 49337
rect 19611 49288 19612 49328
rect 19652 49288 19653 49328
rect 19611 49279 19653 49288
rect 1152 49160 20448 49184
rect 1152 49120 3688 49160
rect 3728 49120 3770 49160
rect 3810 49120 3852 49160
rect 3892 49120 3934 49160
rect 3974 49120 4016 49160
rect 4056 49120 18808 49160
rect 18848 49120 18890 49160
rect 18930 49120 18972 49160
rect 19012 49120 19054 49160
rect 19094 49120 19136 49160
rect 19176 49120 20448 49160
rect 1152 49096 20448 49120
rect 11403 48992 11445 49001
rect 11403 48952 11404 48992
rect 11444 48952 11445 48992
rect 11403 48943 11445 48952
rect 4539 48908 4581 48917
rect 4539 48868 4540 48908
rect 4580 48868 4581 48908
rect 4539 48859 4581 48868
rect 6987 48908 7029 48917
rect 6987 48868 6988 48908
rect 7028 48868 7029 48908
rect 6987 48859 7029 48868
rect 8571 48908 8613 48917
rect 8571 48868 8572 48908
rect 8612 48868 8613 48908
rect 8571 48859 8613 48868
rect 14715 48908 14757 48917
rect 14715 48868 14716 48908
rect 14756 48868 14757 48908
rect 14715 48859 14757 48868
rect 3819 48824 3861 48833
rect 3819 48784 3820 48824
rect 3860 48784 3861 48824
rect 3819 48775 3861 48784
rect 4779 48824 4821 48833
rect 4779 48784 4780 48824
rect 4820 48784 4821 48824
rect 4779 48775 4821 48784
rect 5547 48824 5589 48833
rect 5547 48784 5548 48824
rect 5588 48784 5589 48824
rect 5547 48775 5589 48784
rect 8811 48824 8853 48833
rect 8811 48784 8812 48824
rect 8852 48784 8853 48824
rect 8811 48775 8853 48784
rect 8955 48824 8997 48833
rect 8955 48784 8956 48824
rect 8996 48784 8997 48824
rect 8955 48775 8997 48784
rect 9195 48824 9237 48833
rect 9195 48784 9196 48824
rect 9236 48784 9237 48824
rect 9195 48775 9237 48784
rect 9675 48824 9717 48833
rect 9675 48784 9676 48824
rect 9716 48784 9717 48824
rect 9675 48775 9717 48784
rect 12171 48824 12213 48833
rect 12171 48784 12172 48824
rect 12212 48784 12213 48824
rect 12171 48775 12213 48784
rect 14955 48824 14997 48833
rect 14955 48784 14956 48824
rect 14996 48784 14997 48824
rect 14955 48775 14997 48784
rect 16299 48824 16341 48833
rect 16299 48784 16300 48824
rect 16340 48784 16341 48824
rect 16299 48775 16341 48784
rect 18603 48824 18645 48833
rect 18603 48784 18604 48824
rect 18644 48784 18645 48824
rect 18603 48775 18645 48784
rect 19995 48824 20037 48833
rect 19995 48784 19996 48824
rect 20036 48784 20037 48824
rect 19995 48775 20037 48784
rect 20235 48824 20277 48833
rect 20235 48784 20236 48824
rect 20276 48784 20277 48824
rect 20235 48775 20277 48784
rect 16892 48759 16934 48768
rect 5050 48740 5108 48741
rect 5050 48700 5059 48740
rect 5099 48700 5108 48740
rect 5050 48699 5108 48700
rect 5163 48740 5205 48749
rect 5163 48700 5164 48740
rect 5204 48700 5205 48740
rect 5163 48691 5205 48700
rect 5643 48740 5685 48749
rect 5643 48700 5644 48740
rect 5684 48700 5685 48740
rect 5643 48691 5685 48700
rect 6115 48740 6173 48741
rect 6115 48700 6124 48740
rect 6164 48700 6173 48740
rect 6115 48699 6173 48700
rect 6603 48740 6661 48741
rect 6603 48700 6612 48740
rect 6652 48700 6661 48740
rect 6603 48699 6661 48700
rect 7171 48740 7229 48741
rect 7171 48700 7180 48740
rect 7220 48700 7229 48740
rect 7171 48699 7229 48700
rect 8427 48740 8469 48749
rect 8427 48700 8428 48740
rect 8468 48700 8469 48740
rect 8427 48691 8469 48700
rect 9963 48740 10005 48749
rect 9963 48700 9964 48740
rect 10004 48700 10005 48740
rect 9963 48691 10005 48700
rect 11203 48740 11261 48741
rect 11203 48700 11212 48740
rect 11252 48700 11261 48740
rect 11203 48699 11261 48700
rect 11674 48740 11732 48741
rect 11674 48700 11683 48740
rect 11723 48700 11732 48740
rect 11674 48699 11732 48700
rect 11787 48740 11829 48749
rect 11787 48700 11788 48740
rect 11828 48700 11829 48740
rect 11787 48691 11829 48700
rect 12267 48740 12309 48749
rect 12267 48700 12268 48740
rect 12308 48700 12309 48740
rect 12267 48691 12309 48700
rect 12739 48740 12797 48741
rect 12739 48700 12748 48740
rect 12788 48700 12797 48740
rect 12739 48699 12797 48700
rect 13258 48740 13316 48741
rect 13258 48700 13267 48740
rect 13307 48700 13316 48740
rect 13258 48699 13316 48700
rect 15322 48740 15380 48741
rect 15322 48700 15331 48740
rect 15371 48700 15380 48740
rect 15322 48699 15380 48700
rect 15811 48740 15869 48741
rect 15811 48700 15820 48740
rect 15860 48700 15869 48740
rect 15811 48699 15869 48700
rect 16395 48740 16437 48749
rect 16395 48700 16396 48740
rect 16436 48700 16437 48740
rect 16395 48691 16437 48700
rect 16779 48740 16821 48749
rect 16779 48700 16780 48740
rect 16820 48700 16821 48740
rect 16892 48719 16893 48759
rect 16933 48719 16934 48759
rect 16892 48710 16934 48719
rect 18106 48740 18164 48741
rect 16779 48691 16821 48700
rect 18106 48700 18115 48740
rect 18155 48700 18164 48740
rect 18106 48699 18164 48700
rect 18219 48740 18261 48749
rect 18219 48700 18220 48740
rect 18260 48700 18261 48740
rect 18219 48691 18261 48700
rect 18699 48740 18741 48749
rect 18699 48700 18700 48740
rect 18740 48700 18741 48740
rect 18699 48691 18741 48700
rect 19171 48740 19229 48741
rect 19171 48700 19180 48740
rect 19220 48700 19229 48740
rect 19171 48699 19229 48700
rect 19659 48740 19717 48741
rect 19659 48700 19668 48740
rect 19708 48700 19717 48740
rect 19659 48699 19717 48700
rect 4059 48572 4101 48581
rect 4059 48532 4060 48572
rect 4100 48532 4101 48572
rect 4059 48523 4101 48532
rect 6795 48572 6837 48581
rect 6795 48532 6796 48572
rect 6836 48532 6837 48572
rect 6795 48523 6837 48532
rect 9435 48572 9477 48581
rect 9435 48532 9436 48572
rect 9476 48532 9477 48572
rect 9435 48523 9477 48532
rect 13419 48572 13461 48581
rect 13419 48532 13420 48572
rect 13460 48532 13461 48572
rect 13419 48523 13461 48532
rect 15147 48572 15189 48581
rect 15147 48532 15148 48572
rect 15188 48532 15189 48572
rect 15147 48523 15189 48532
rect 19851 48572 19893 48581
rect 19851 48532 19852 48572
rect 19892 48532 19893 48572
rect 19851 48523 19893 48532
rect 1152 48404 20452 48428
rect 1152 48364 4928 48404
rect 4968 48364 5010 48404
rect 5050 48364 5092 48404
rect 5132 48364 5174 48404
rect 5214 48364 5256 48404
rect 5296 48364 20048 48404
rect 20088 48364 20130 48404
rect 20170 48364 20212 48404
rect 20252 48364 20294 48404
rect 20334 48364 20376 48404
rect 20416 48364 20452 48404
rect 1152 48340 20452 48364
rect 3915 48236 3957 48245
rect 3915 48196 3916 48236
rect 3956 48196 3957 48236
rect 3915 48187 3957 48196
rect 5931 48236 5973 48245
rect 5931 48196 5932 48236
rect 5972 48196 5973 48236
rect 5931 48187 5973 48196
rect 17451 48236 17493 48245
rect 17451 48196 17452 48236
rect 17492 48196 17493 48236
rect 17451 48187 17493 48196
rect 19083 48236 19125 48245
rect 19083 48196 19084 48236
rect 19124 48196 19125 48236
rect 19083 48187 19125 48196
rect 20379 48236 20421 48245
rect 20379 48196 20380 48236
rect 20420 48196 20421 48236
rect 20379 48187 20421 48196
rect 2170 48068 2228 48069
rect 2170 48028 2179 48068
rect 2219 48028 2228 48068
rect 2170 48027 2228 48028
rect 2283 48068 2325 48077
rect 2283 48028 2284 48068
rect 2324 48028 2325 48068
rect 2283 48019 2325 48028
rect 2667 48068 2709 48077
rect 4173 48068 4215 48077
rect 2667 48028 2668 48068
rect 2708 48028 2709 48068
rect 2667 48019 2709 48028
rect 3243 48059 3285 48068
rect 3243 48019 3244 48059
rect 3284 48019 3285 48059
rect 3243 48010 3285 48019
rect 3723 48059 3765 48068
rect 3723 48019 3724 48059
rect 3764 48019 3765 48059
rect 4173 48028 4174 48068
rect 4214 48028 4215 48068
rect 4173 48019 4215 48028
rect 4297 48068 4339 48077
rect 4297 48028 4298 48068
rect 4338 48028 4339 48068
rect 4297 48019 4339 48028
rect 4683 48068 4725 48077
rect 12939 48068 12981 48077
rect 15706 48068 15764 48069
rect 4683 48028 4684 48068
rect 4724 48028 4725 48068
rect 4683 48019 4725 48028
rect 5259 48059 5301 48068
rect 5259 48019 5260 48059
rect 5300 48019 5301 48059
rect 3723 48010 3765 48019
rect 5259 48010 5301 48019
rect 5739 48059 5781 48068
rect 5739 48019 5740 48059
rect 5780 48019 5781 48059
rect 12939 48028 12940 48068
rect 12980 48028 12981 48068
rect 12939 48019 12981 48028
rect 14187 48059 14229 48068
rect 14187 48019 14188 48059
rect 14228 48019 14229 48059
rect 15706 48028 15715 48068
rect 15755 48028 15764 48068
rect 15706 48027 15764 48028
rect 15819 48068 15861 48077
rect 15819 48028 15820 48068
rect 15860 48028 15861 48068
rect 15819 48019 15861 48028
rect 16203 48068 16245 48077
rect 17643 48068 17685 48077
rect 16203 48028 16204 48068
rect 16244 48028 16245 48068
rect 16203 48019 16245 48028
rect 16779 48059 16821 48068
rect 16779 48019 16780 48059
rect 16820 48019 16821 48059
rect 5739 48010 5781 48019
rect 14187 48010 14229 48019
rect 16779 48010 16821 48019
rect 17259 48059 17301 48068
rect 17259 48019 17260 48059
rect 17300 48019 17301 48059
rect 17643 48028 17644 48068
rect 17684 48028 17685 48068
rect 17643 48019 17685 48028
rect 18891 48059 18933 48068
rect 18891 48019 18892 48059
rect 18932 48019 18933 48059
rect 17259 48010 17301 48019
rect 18891 48010 18933 48019
rect 2763 47984 2805 47993
rect 2763 47944 2764 47984
rect 2804 47944 2805 47984
rect 2763 47935 2805 47944
rect 4779 47984 4821 47993
rect 4779 47944 4780 47984
rect 4820 47944 4821 47984
rect 4779 47935 4821 47944
rect 7947 47984 7989 47993
rect 7947 47944 7948 47984
rect 7988 47944 7989 47984
rect 7947 47935 7989 47944
rect 9291 47984 9333 47993
rect 9291 47944 9292 47984
rect 9332 47944 9333 47984
rect 9291 47935 9333 47944
rect 9675 47984 9717 47993
rect 9675 47944 9676 47984
rect 9716 47944 9717 47984
rect 9675 47935 9717 47944
rect 10347 47984 10389 47993
rect 10347 47944 10348 47984
rect 10388 47944 10389 47984
rect 10347 47935 10389 47944
rect 10923 47984 10965 47993
rect 10923 47944 10924 47984
rect 10964 47944 10965 47984
rect 10923 47935 10965 47944
rect 16299 47984 16341 47993
rect 16299 47944 16300 47984
rect 16340 47944 16341 47984
rect 16299 47935 16341 47944
rect 19755 47984 19797 47993
rect 19755 47944 19756 47984
rect 19796 47944 19797 47984
rect 19755 47935 19797 47944
rect 20139 47984 20181 47993
rect 20139 47944 20140 47984
rect 20180 47944 20181 47984
rect 20139 47935 20181 47944
rect 10587 47900 10629 47909
rect 10587 47860 10588 47900
rect 10628 47860 10629 47900
rect 10587 47851 10629 47860
rect 19995 47900 20037 47909
rect 19995 47860 19996 47900
rect 20036 47860 20037 47900
rect 19995 47851 20037 47860
rect 8187 47816 8229 47825
rect 8187 47776 8188 47816
rect 8228 47776 8229 47816
rect 8187 47767 8229 47776
rect 9051 47816 9093 47825
rect 9051 47776 9052 47816
rect 9092 47776 9093 47816
rect 9051 47767 9093 47776
rect 9915 47816 9957 47825
rect 9915 47776 9916 47816
rect 9956 47776 9957 47816
rect 9915 47767 9957 47776
rect 10683 47816 10725 47825
rect 10683 47776 10684 47816
rect 10724 47776 10725 47816
rect 10683 47767 10725 47776
rect 14379 47816 14421 47825
rect 14379 47776 14380 47816
rect 14420 47776 14421 47816
rect 14379 47767 14421 47776
rect 1152 47648 20448 47672
rect 1152 47608 3688 47648
rect 3728 47608 3770 47648
rect 3810 47608 3852 47648
rect 3892 47608 3934 47648
rect 3974 47608 4016 47648
rect 4056 47608 18808 47648
rect 18848 47608 18890 47648
rect 18930 47608 18972 47648
rect 19012 47608 19054 47648
rect 19094 47608 19136 47648
rect 19176 47608 20448 47648
rect 1152 47584 20448 47608
rect 3051 47480 3093 47489
rect 3051 47440 3052 47480
rect 3092 47440 3093 47480
rect 3051 47431 3093 47440
rect 9802 47480 9860 47481
rect 9802 47440 9811 47480
rect 9851 47440 9860 47480
rect 9802 47439 9860 47440
rect 15819 47480 15861 47489
rect 15819 47440 15820 47480
rect 15860 47440 15861 47480
rect 15819 47431 15861 47440
rect 17451 47480 17493 47489
rect 17451 47440 17452 47480
rect 17492 47440 17493 47480
rect 17451 47431 17493 47440
rect 19467 47480 19509 47489
rect 19467 47440 19468 47480
rect 19508 47440 19509 47480
rect 19467 47431 19509 47440
rect 3819 47312 3861 47321
rect 3819 47272 3820 47312
rect 3860 47272 3861 47312
rect 3819 47263 3861 47272
rect 8523 47312 8565 47321
rect 8523 47272 8524 47312
rect 8564 47272 8565 47312
rect 8523 47263 8565 47272
rect 19755 47312 19797 47321
rect 19755 47272 19756 47312
rect 19796 47272 19797 47312
rect 19755 47263 19797 47272
rect 20139 47312 20181 47321
rect 20139 47272 20140 47312
rect 20180 47272 20181 47312
rect 20139 47263 20181 47272
rect 20379 47312 20421 47321
rect 20379 47272 20380 47312
rect 20420 47272 20421 47312
rect 20379 47263 20421 47272
rect 1611 47228 1653 47237
rect 1611 47188 1612 47228
rect 1652 47188 1653 47228
rect 1611 47179 1653 47188
rect 2851 47228 2909 47229
rect 2851 47188 2860 47228
rect 2900 47188 2909 47228
rect 2851 47187 2909 47188
rect 3322 47228 3380 47229
rect 3322 47188 3331 47228
rect 3371 47188 3380 47228
rect 3322 47187 3380 47188
rect 3435 47228 3477 47237
rect 3435 47188 3436 47228
rect 3476 47188 3477 47228
rect 3435 47179 3477 47188
rect 3915 47228 3957 47237
rect 3915 47188 3916 47228
rect 3956 47188 3957 47228
rect 3915 47179 3957 47188
rect 4387 47228 4445 47229
rect 4387 47188 4396 47228
rect 4436 47188 4445 47228
rect 4387 47187 4445 47188
rect 4875 47228 4933 47229
rect 4875 47188 4884 47228
rect 4924 47188 4933 47228
rect 4875 47187 4933 47188
rect 6123 47228 6165 47237
rect 6123 47188 6124 47228
rect 6164 47188 6165 47228
rect 6123 47179 6165 47188
rect 6315 47228 6357 47237
rect 6315 47188 6316 47228
rect 6356 47188 6357 47228
rect 6315 47179 6357 47188
rect 7555 47228 7613 47229
rect 7555 47188 7564 47228
rect 7604 47188 7613 47228
rect 7555 47187 7613 47188
rect 8026 47228 8084 47229
rect 8026 47188 8035 47228
rect 8075 47188 8084 47228
rect 8026 47187 8084 47188
rect 8139 47228 8181 47237
rect 8139 47188 8140 47228
rect 8180 47188 8181 47228
rect 8139 47179 8181 47188
rect 8619 47228 8661 47237
rect 8619 47188 8620 47228
rect 8660 47188 8661 47228
rect 8619 47179 8661 47188
rect 9091 47228 9149 47229
rect 9091 47188 9100 47228
rect 9140 47188 9149 47228
rect 9091 47187 9149 47188
rect 9579 47228 9637 47229
rect 9579 47188 9588 47228
rect 9628 47188 9637 47228
rect 9579 47187 9637 47188
rect 10443 47228 10485 47237
rect 10443 47188 10444 47228
rect 10484 47188 10485 47228
rect 10443 47179 10485 47188
rect 10827 47228 10869 47237
rect 10827 47188 10828 47228
rect 10868 47188 10869 47228
rect 10827 47179 10869 47188
rect 12067 47228 12125 47229
rect 12067 47188 12076 47228
rect 12116 47188 12125 47228
rect 12067 47187 12125 47188
rect 12747 47228 12789 47237
rect 12747 47188 12748 47228
rect 12788 47188 12789 47228
rect 12747 47179 12789 47188
rect 13987 47228 14045 47229
rect 13987 47188 13996 47228
rect 14036 47188 14045 47228
rect 13987 47187 14045 47188
rect 14379 47228 14421 47237
rect 14379 47188 14380 47228
rect 14420 47188 14421 47228
rect 14379 47179 14421 47188
rect 15619 47228 15677 47229
rect 15619 47188 15628 47228
rect 15668 47188 15677 47228
rect 15619 47187 15677 47188
rect 16011 47228 16053 47237
rect 16011 47188 16012 47228
rect 16052 47188 16053 47228
rect 16011 47179 16053 47188
rect 17251 47228 17309 47229
rect 17251 47188 17260 47228
rect 17300 47188 17309 47228
rect 17251 47187 17309 47188
rect 18027 47228 18069 47237
rect 18027 47188 18028 47228
rect 18068 47188 18069 47228
rect 18027 47179 18069 47188
rect 19267 47228 19325 47229
rect 19267 47188 19276 47228
rect 19316 47188 19325 47228
rect 19267 47187 19325 47188
rect 7755 47144 7797 47153
rect 7755 47104 7756 47144
rect 7796 47104 7797 47144
rect 7755 47095 7797 47104
rect 5067 47060 5109 47069
rect 5067 47020 5068 47060
rect 5108 47020 5109 47060
rect 5067 47011 5109 47020
rect 5979 47060 6021 47069
rect 5979 47020 5980 47060
rect 6020 47020 6021 47060
rect 5979 47011 6021 47020
rect 10587 47060 10629 47069
rect 10587 47020 10588 47060
rect 10628 47020 10629 47060
rect 10587 47011 10629 47020
rect 12267 47060 12309 47069
rect 12267 47020 12268 47060
rect 12308 47020 12309 47060
rect 12267 47011 12309 47020
rect 14187 47060 14229 47069
rect 14187 47020 14188 47060
rect 14228 47020 14229 47060
rect 14187 47011 14229 47020
rect 19995 47060 20037 47069
rect 19995 47020 19996 47060
rect 20036 47020 20037 47060
rect 19995 47011 20037 47020
rect 1152 46892 20452 46916
rect 1152 46852 4928 46892
rect 4968 46852 5010 46892
rect 5050 46852 5092 46892
rect 5132 46852 5174 46892
rect 5214 46852 5256 46892
rect 5296 46852 20048 46892
rect 20088 46852 20130 46892
rect 20170 46852 20212 46892
rect 20252 46852 20294 46892
rect 20334 46852 20376 46892
rect 20416 46852 20452 46892
rect 1152 46828 20452 46852
rect 2763 46724 2805 46733
rect 2763 46684 2764 46724
rect 2804 46684 2805 46724
rect 2763 46675 2805 46684
rect 3867 46724 3909 46733
rect 3867 46684 3868 46724
rect 3908 46684 3909 46724
rect 3867 46675 3909 46684
rect 4347 46724 4389 46733
rect 4347 46684 4348 46724
rect 4388 46684 4389 46724
rect 4347 46675 4389 46684
rect 5355 46724 5397 46733
rect 5355 46684 5356 46724
rect 5396 46684 5397 46724
rect 5355 46675 5397 46684
rect 9387 46724 9429 46733
rect 9387 46684 9388 46724
rect 9428 46684 9429 46724
rect 9387 46675 9429 46684
rect 10347 46724 10389 46733
rect 10347 46684 10348 46724
rect 10388 46684 10389 46724
rect 10347 46675 10389 46684
rect 15147 46724 15189 46733
rect 15147 46684 15148 46724
rect 15188 46684 15189 46724
rect 15147 46675 15189 46684
rect 1323 46556 1365 46565
rect 4954 46556 5012 46557
rect 6755 46556 6797 46565
rect 1323 46516 1324 46556
rect 1364 46516 1365 46556
rect 1323 46507 1365 46516
rect 2571 46547 2613 46556
rect 2571 46507 2572 46547
rect 2612 46507 2613 46547
rect 4954 46516 4963 46556
rect 5003 46516 5012 46556
rect 4954 46515 5012 46516
rect 5547 46547 5589 46556
rect 2571 46498 2613 46507
rect 5547 46507 5548 46547
rect 5588 46507 5589 46547
rect 6755 46516 6756 46556
rect 6796 46516 6797 46556
rect 6755 46507 6797 46516
rect 6987 46556 7029 46565
rect 6987 46516 6988 46556
rect 7028 46516 7029 46556
rect 6987 46507 7029 46516
rect 7179 46556 7221 46565
rect 7179 46516 7180 46556
rect 7220 46516 7221 46556
rect 7179 46507 7221 46516
rect 7323 46556 7365 46565
rect 7323 46516 7324 46556
rect 7364 46516 7365 46556
rect 7323 46507 7365 46516
rect 7467 46556 7509 46565
rect 7467 46516 7468 46556
rect 7508 46516 7509 46556
rect 7467 46507 7509 46516
rect 7947 46556 7989 46565
rect 9579 46556 9621 46565
rect 7947 46516 7948 46556
rect 7988 46516 7989 46556
rect 7947 46507 7989 46516
rect 9195 46547 9237 46556
rect 9195 46507 9196 46547
rect 9236 46507 9237 46547
rect 9579 46516 9580 46556
rect 9620 46516 9621 46556
rect 9579 46507 9621 46516
rect 9754 46556 9812 46557
rect 9754 46516 9763 46556
rect 9803 46516 9812 46556
rect 9754 46515 9812 46516
rect 9867 46556 9909 46565
rect 9867 46516 9868 46556
rect 9908 46516 9909 46556
rect 9867 46507 9909 46516
rect 10059 46556 10101 46565
rect 10059 46516 10060 46556
rect 10100 46516 10101 46556
rect 10059 46507 10101 46516
rect 10193 46556 10251 46557
rect 10193 46516 10202 46556
rect 10242 46516 10251 46556
rect 10193 46515 10251 46516
rect 10618 46556 10676 46557
rect 10618 46516 10627 46556
rect 10667 46516 10676 46556
rect 10618 46515 10676 46516
rect 10731 46556 10773 46565
rect 10731 46516 10732 46556
rect 10772 46516 10773 46556
rect 10731 46507 10773 46516
rect 11115 46556 11157 46565
rect 13402 46556 13460 46557
rect 11115 46516 11116 46556
rect 11156 46516 11157 46556
rect 11115 46507 11157 46516
rect 11691 46547 11733 46556
rect 11691 46507 11692 46547
rect 11732 46507 11733 46547
rect 5547 46498 5589 46507
rect 9195 46498 9237 46507
rect 11691 46498 11733 46507
rect 12171 46547 12213 46556
rect 12171 46507 12172 46547
rect 12212 46507 12213 46547
rect 13402 46516 13411 46556
rect 13451 46516 13460 46556
rect 13402 46515 13460 46516
rect 13515 46556 13557 46565
rect 13515 46516 13516 46556
rect 13556 46516 13557 46556
rect 13515 46507 13557 46516
rect 13899 46556 13941 46565
rect 16779 46556 16821 46565
rect 13899 46516 13900 46556
rect 13940 46516 13941 46556
rect 13899 46507 13941 46516
rect 14475 46547 14517 46556
rect 14475 46507 14476 46547
rect 14516 46507 14517 46547
rect 12171 46498 12213 46507
rect 14475 46498 14517 46507
rect 14955 46547 14997 46556
rect 14955 46507 14956 46547
rect 14996 46507 14997 46547
rect 14955 46498 14997 46507
rect 15531 46547 15573 46556
rect 15531 46507 15532 46547
rect 15572 46507 15573 46547
rect 16779 46516 16780 46556
rect 16820 46516 16821 46556
rect 16779 46507 16821 46516
rect 17835 46556 17877 46565
rect 17835 46516 17836 46556
rect 17876 46516 17877 46556
rect 17835 46507 17877 46516
rect 19083 46547 19125 46556
rect 19083 46507 19084 46547
rect 19124 46507 19125 46547
rect 15531 46498 15573 46507
rect 19083 46498 19125 46507
rect 3627 46472 3669 46481
rect 3627 46432 3628 46472
rect 3668 46432 3669 46472
rect 3627 46423 3669 46432
rect 4107 46472 4149 46481
rect 4107 46432 4108 46472
rect 4148 46432 4149 46472
rect 4107 46423 4149 46432
rect 4491 46472 4533 46481
rect 4491 46432 4492 46472
rect 4532 46432 4533 46472
rect 4491 46423 4533 46432
rect 11211 46472 11253 46481
rect 11211 46432 11212 46472
rect 11252 46432 11253 46472
rect 11211 46423 11253 46432
rect 12394 46472 12452 46473
rect 12394 46432 12403 46472
rect 12443 46432 12452 46472
rect 12394 46431 12452 46432
rect 12747 46472 12789 46481
rect 12747 46432 12748 46472
rect 12788 46432 12789 46472
rect 12747 46423 12789 46432
rect 13995 46472 14037 46481
rect 13995 46432 13996 46472
rect 14036 46432 14037 46472
rect 13995 46423 14037 46432
rect 19755 46472 19797 46481
rect 19755 46432 19756 46472
rect 19796 46432 19797 46472
rect 19755 46423 19797 46432
rect 20139 46472 20181 46481
rect 20139 46432 20140 46472
rect 20180 46432 20181 46472
rect 20139 46423 20181 46432
rect 4934 46388 4976 46397
rect 4934 46348 4935 46388
rect 4975 46348 4976 46388
rect 4934 46339 4976 46348
rect 5146 46388 5204 46389
rect 5146 46348 5155 46388
rect 5195 46348 5204 46388
rect 5146 46347 5204 46348
rect 19995 46388 20037 46397
rect 19995 46348 19996 46388
rect 20036 46348 20037 46388
rect 19995 46339 20037 46348
rect 4731 46304 4773 46313
rect 4731 46264 4732 46304
rect 4772 46264 4773 46304
rect 4731 46255 4773 46264
rect 7083 46304 7125 46313
rect 7083 46264 7084 46304
rect 7124 46264 7125 46304
rect 7083 46255 7125 46264
rect 9867 46304 9909 46313
rect 9867 46264 9868 46304
rect 9908 46264 9909 46304
rect 9867 46255 9909 46264
rect 12507 46304 12549 46313
rect 12507 46264 12508 46304
rect 12548 46264 12549 46304
rect 12507 46255 12549 46264
rect 15339 46304 15381 46313
rect 15339 46264 15340 46304
rect 15380 46264 15381 46304
rect 15339 46255 15381 46264
rect 19275 46304 19317 46313
rect 19275 46264 19276 46304
rect 19316 46264 19317 46304
rect 19275 46255 19317 46264
rect 20379 46304 20421 46313
rect 20379 46264 20380 46304
rect 20420 46264 20421 46304
rect 20379 46255 20421 46264
rect 1152 46136 20448 46160
rect 1152 46096 3688 46136
rect 3728 46096 3770 46136
rect 3810 46096 3852 46136
rect 3892 46096 3934 46136
rect 3974 46096 4016 46136
rect 4056 46096 18808 46136
rect 18848 46096 18890 46136
rect 18930 46096 18972 46136
rect 19012 46096 19054 46136
rect 19094 46096 19136 46136
rect 19176 46096 20448 46136
rect 1152 46072 20448 46096
rect 1851 45968 1893 45977
rect 1851 45928 1852 45968
rect 1892 45928 1893 45968
rect 1851 45919 1893 45928
rect 4683 45968 4725 45977
rect 4683 45928 4684 45968
rect 4724 45928 4725 45968
rect 4683 45919 4725 45928
rect 9771 45968 9813 45977
rect 9771 45928 9772 45968
rect 9812 45928 9813 45968
rect 9771 45919 9813 45928
rect 11403 45968 11445 45977
rect 11403 45928 11404 45968
rect 11444 45928 11445 45968
rect 11403 45919 11445 45928
rect 13419 45968 13461 45977
rect 13419 45928 13420 45968
rect 13460 45928 13461 45968
rect 13419 45919 13461 45928
rect 1467 45884 1509 45893
rect 1467 45844 1468 45884
rect 1508 45844 1509 45884
rect 1467 45835 1509 45844
rect 5067 45884 5109 45893
rect 5067 45844 5068 45884
rect 5108 45844 5109 45884
rect 5067 45835 5109 45844
rect 7467 45884 7509 45893
rect 7467 45844 7468 45884
rect 7508 45844 7509 45884
rect 7467 45835 7509 45844
rect 11835 45884 11877 45893
rect 11835 45844 11836 45884
rect 11876 45844 11877 45884
rect 11835 45835 11877 45844
rect 1227 45800 1269 45809
rect 1227 45760 1228 45800
rect 1268 45760 1269 45800
rect 1227 45751 1269 45760
rect 1611 45800 1653 45809
rect 1611 45760 1612 45800
rect 1652 45760 1653 45800
rect 5163 45800 5205 45809
rect 1611 45751 1653 45760
rect 4999 45758 5041 45767
rect 3915 45716 3957 45725
rect 3915 45676 3916 45716
rect 3956 45676 3957 45716
rect 3915 45667 3957 45676
rect 4049 45716 4107 45717
rect 4049 45676 4058 45716
rect 4098 45676 4107 45716
rect 4049 45675 4107 45676
rect 4395 45716 4437 45725
rect 4395 45676 4396 45716
rect 4436 45676 4437 45716
rect 4395 45667 4437 45676
rect 4550 45716 4592 45725
rect 4550 45676 4551 45716
rect 4591 45676 4592 45716
rect 4550 45667 4592 45676
rect 4673 45716 4715 45725
rect 4673 45676 4674 45716
rect 4714 45676 4715 45716
rect 4673 45667 4715 45676
rect 4851 45716 4893 45725
rect 4851 45676 4852 45716
rect 4892 45676 4893 45716
rect 4999 45718 5000 45758
rect 5040 45718 5041 45758
rect 5163 45760 5164 45800
rect 5204 45760 5205 45800
rect 5163 45751 5205 45760
rect 6914 45800 6956 45809
rect 6914 45760 6915 45800
rect 6955 45760 6956 45800
rect 6914 45751 6956 45760
rect 11595 45800 11637 45809
rect 11595 45760 11596 45800
rect 11636 45760 11637 45800
rect 11595 45751 11637 45760
rect 14667 45800 14709 45809
rect 14667 45760 14668 45800
rect 14708 45760 14709 45800
rect 14667 45751 14709 45760
rect 17547 45800 17589 45809
rect 17547 45760 17548 45800
rect 17588 45760 17589 45800
rect 17547 45751 17589 45760
rect 18315 45800 18357 45809
rect 18315 45760 18316 45800
rect 18356 45760 18357 45800
rect 18315 45751 18357 45760
rect 19755 45800 19797 45809
rect 19755 45760 19756 45800
rect 19796 45760 19797 45800
rect 19755 45751 19797 45760
rect 20139 45800 20181 45809
rect 20139 45760 20140 45800
rect 20180 45760 20181 45800
rect 20139 45751 20181 45760
rect 4999 45709 5041 45718
rect 5284 45716 5326 45725
rect 4851 45667 4893 45676
rect 5284 45676 5285 45716
rect 5325 45676 5326 45716
rect 5284 45667 5326 45676
rect 5434 45716 5492 45717
rect 5434 45676 5443 45716
rect 5483 45676 5492 45716
rect 5434 45675 5492 45676
rect 5578 45716 5636 45717
rect 5578 45676 5587 45716
rect 5627 45676 5636 45716
rect 5578 45675 5636 45676
rect 5692 45716 5750 45717
rect 5692 45676 5701 45716
rect 5741 45676 5750 45716
rect 5692 45675 5750 45676
rect 5818 45716 5876 45717
rect 5818 45676 5827 45716
rect 5867 45676 5876 45716
rect 5818 45675 5876 45676
rect 5995 45716 6053 45717
rect 5995 45676 6004 45716
rect 6044 45676 6053 45716
rect 5995 45675 6053 45676
rect 6219 45716 6261 45725
rect 6219 45676 6220 45716
rect 6260 45676 6261 45716
rect 6219 45667 6261 45676
rect 6353 45716 6411 45717
rect 6353 45676 6362 45716
rect 6402 45676 6411 45716
rect 6353 45675 6411 45676
rect 6795 45716 6837 45725
rect 6795 45676 6796 45716
rect 6836 45676 6837 45716
rect 6795 45667 6837 45676
rect 7024 45716 7082 45717
rect 7024 45676 7033 45716
rect 7073 45676 7082 45716
rect 7024 45675 7082 45676
rect 7176 45716 7218 45725
rect 7176 45676 7177 45716
rect 7217 45676 7218 45716
rect 7176 45667 7218 45676
rect 7306 45716 7364 45717
rect 7306 45676 7315 45716
rect 7355 45676 7364 45716
rect 7306 45675 7364 45676
rect 7420 45716 7478 45717
rect 7420 45676 7429 45716
rect 7469 45676 7478 45716
rect 7420 45675 7478 45676
rect 7755 45716 7797 45725
rect 7755 45676 7756 45716
rect 7796 45676 7797 45716
rect 7755 45667 7797 45676
rect 7874 45716 7916 45725
rect 7874 45676 7875 45716
rect 7915 45676 7916 45716
rect 7874 45667 7916 45676
rect 7984 45716 8042 45717
rect 7984 45676 7993 45716
rect 8033 45676 8042 45716
rect 7984 45675 8042 45676
rect 8331 45716 8373 45725
rect 8331 45676 8332 45716
rect 8372 45676 8373 45716
rect 8331 45667 8373 45676
rect 9571 45716 9629 45717
rect 9571 45676 9580 45716
rect 9620 45676 9629 45716
rect 9571 45675 9629 45676
rect 9963 45716 10005 45725
rect 9963 45676 9964 45716
rect 10004 45676 10005 45716
rect 9963 45667 10005 45676
rect 11203 45716 11261 45717
rect 11203 45676 11212 45716
rect 11252 45676 11261 45716
rect 11203 45675 11261 45676
rect 11979 45716 12021 45725
rect 11979 45676 11980 45716
rect 12020 45676 12021 45716
rect 11979 45667 12021 45676
rect 13219 45716 13277 45717
rect 13219 45676 13228 45716
rect 13268 45676 13277 45716
rect 13219 45675 13277 45676
rect 14170 45716 14228 45717
rect 14170 45676 14179 45716
rect 14219 45676 14228 45716
rect 14170 45675 14228 45676
rect 14283 45716 14325 45725
rect 14283 45676 14284 45716
rect 14324 45676 14325 45716
rect 14283 45667 14325 45676
rect 14763 45716 14805 45725
rect 14763 45676 14764 45716
rect 14804 45676 14805 45716
rect 14763 45667 14805 45676
rect 15235 45716 15293 45717
rect 15235 45676 15244 45716
rect 15284 45676 15293 45716
rect 15235 45675 15293 45676
rect 15723 45716 15781 45717
rect 15723 45676 15732 45716
rect 15772 45676 15781 45716
rect 15723 45675 15781 45676
rect 17818 45716 17876 45717
rect 17818 45676 17827 45716
rect 17867 45676 17876 45716
rect 17818 45675 17876 45676
rect 17931 45716 17973 45725
rect 17931 45676 17932 45716
rect 17972 45676 17973 45716
rect 17931 45667 17973 45676
rect 18411 45716 18453 45725
rect 18411 45676 18412 45716
rect 18452 45676 18453 45716
rect 18411 45667 18453 45676
rect 18883 45716 18941 45717
rect 18883 45676 18892 45716
rect 18932 45676 18941 45716
rect 18883 45675 18941 45676
rect 19371 45716 19429 45717
rect 19371 45676 19380 45716
rect 19420 45676 19429 45716
rect 19371 45675 19429 45676
rect 6699 45632 6741 45641
rect 6699 45592 6700 45632
rect 6740 45592 6741 45632
rect 6699 45583 6741 45592
rect 7659 45632 7701 45641
rect 7659 45592 7660 45632
rect 7700 45592 7701 45632
rect 7659 45583 7701 45592
rect 19995 45632 20037 45641
rect 19995 45592 19996 45632
rect 20036 45592 20037 45632
rect 19995 45583 20037 45592
rect 4203 45548 4245 45557
rect 4203 45508 4204 45548
rect 4244 45508 4245 45548
rect 4203 45499 4245 45508
rect 5914 45548 5972 45549
rect 5914 45508 5923 45548
rect 5963 45508 5972 45548
rect 5914 45507 5972 45508
rect 6507 45548 6549 45557
rect 6507 45508 6508 45548
rect 6548 45508 6549 45548
rect 6507 45499 6549 45508
rect 9771 45548 9813 45557
rect 9771 45508 9772 45548
rect 9812 45508 9813 45548
rect 9771 45499 9813 45508
rect 15915 45548 15957 45557
rect 15915 45508 15916 45548
rect 15956 45508 15957 45548
rect 15915 45499 15957 45508
rect 17307 45548 17349 45557
rect 17307 45508 17308 45548
rect 17348 45508 17349 45548
rect 17307 45499 17349 45508
rect 19563 45548 19605 45557
rect 19563 45508 19564 45548
rect 19604 45508 19605 45548
rect 19563 45499 19605 45508
rect 20379 45548 20421 45557
rect 20379 45508 20380 45548
rect 20420 45508 20421 45548
rect 20379 45499 20421 45508
rect 1152 45380 20452 45404
rect 1152 45340 4928 45380
rect 4968 45340 5010 45380
rect 5050 45340 5092 45380
rect 5132 45340 5174 45380
rect 5214 45340 5256 45380
rect 5296 45340 20048 45380
rect 20088 45340 20130 45380
rect 20170 45340 20212 45380
rect 20252 45340 20294 45380
rect 20334 45340 20376 45380
rect 20416 45340 20452 45380
rect 1152 45316 20452 45340
rect 4203 45212 4245 45221
rect 4203 45172 4204 45212
rect 4244 45172 4245 45212
rect 4203 45163 4245 45172
rect 5451 45212 5493 45221
rect 5451 45172 5452 45212
rect 5492 45172 5493 45212
rect 5451 45163 5493 45172
rect 5722 45212 5780 45213
rect 5722 45172 5731 45212
rect 5771 45172 5780 45212
rect 5722 45171 5780 45172
rect 8139 45212 8181 45221
rect 8139 45172 8140 45212
rect 8180 45172 8181 45212
rect 8139 45163 8181 45172
rect 10635 45212 10677 45221
rect 10635 45172 10636 45212
rect 10676 45172 10677 45212
rect 10635 45163 10677 45172
rect 11931 45212 11973 45221
rect 11931 45172 11932 45212
rect 11972 45172 11973 45212
rect 11931 45163 11973 45172
rect 15243 45212 15285 45221
rect 15243 45172 15244 45212
rect 15284 45172 15285 45212
rect 15243 45163 15285 45172
rect 17451 45212 17493 45221
rect 17451 45172 17452 45212
rect 17492 45172 17493 45212
rect 17451 45163 17493 45172
rect 19755 45212 19797 45221
rect 19755 45172 19756 45212
rect 19796 45172 19797 45212
rect 19755 45163 19797 45172
rect 5632 45128 5674 45137
rect 5632 45088 5633 45128
rect 5673 45088 5674 45128
rect 5632 45079 5674 45088
rect 6315 45128 6357 45137
rect 6315 45088 6316 45128
rect 6356 45088 6357 45128
rect 6315 45079 6357 45088
rect 11106 45119 11152 45128
rect 11106 45079 11107 45119
rect 11147 45079 11152 45119
rect 11106 45070 11152 45079
rect 2763 45044 2805 45053
rect 4395 45044 4437 45053
rect 2763 45004 2764 45044
rect 2804 45004 2805 45044
rect 2763 44995 2805 45004
rect 4011 45035 4053 45044
rect 4011 44995 4012 45035
rect 4052 44995 4053 45035
rect 4395 45004 4396 45044
rect 4436 45004 4437 45044
rect 4395 44995 4437 45004
rect 4564 45044 4606 45053
rect 4564 45004 4565 45044
rect 4605 45004 4606 45044
rect 4564 44995 4606 45004
rect 4683 45044 4725 45053
rect 4683 45004 4684 45044
rect 4724 45004 4725 45044
rect 4683 44995 4725 45004
rect 5067 45044 5109 45053
rect 5067 45004 5068 45044
rect 5108 45004 5109 45044
rect 5067 44995 5109 45004
rect 5181 45044 5239 45045
rect 5835 45044 5877 45053
rect 6109 45044 6151 45053
rect 6747 45044 6789 45053
rect 5181 45004 5190 45044
rect 5230 45004 5239 45044
rect 5181 45003 5239 45004
rect 5406 45035 5448 45044
rect 5296 45002 5354 45003
rect 4011 44986 4053 44995
rect 1227 44960 1269 44969
rect 1227 44920 1228 44960
rect 1268 44920 1269 44960
rect 1227 44911 1269 44920
rect 1611 44960 1653 44969
rect 5296 44962 5305 45002
rect 5345 44962 5354 45002
rect 5406 44995 5407 45035
rect 5447 44995 5448 45035
rect 5835 45004 5836 45044
rect 5876 45004 5877 45044
rect 5835 44995 5877 45004
rect 5931 45035 5973 45044
rect 5931 44995 5932 45035
rect 5972 44995 5973 45035
rect 6109 45004 6110 45044
rect 6150 45004 6151 45044
rect 6109 44995 6151 45004
rect 6411 45035 6453 45044
rect 6411 44995 6412 45035
rect 6452 44995 6453 45035
rect 6747 45004 6748 45044
rect 6788 45004 6789 45044
rect 6747 44995 6789 45004
rect 7048 45044 7090 45053
rect 7048 45004 7049 45044
rect 7089 45004 7090 45044
rect 7048 44995 7090 45004
rect 7210 45044 7268 45045
rect 8235 45044 8277 45053
rect 7210 45004 7219 45044
rect 7259 45004 7268 45044
rect 7210 45003 7268 45004
rect 7563 45035 7605 45044
rect 7563 44995 7564 45035
rect 7604 44995 7605 45035
rect 5406 44986 5448 44995
rect 5931 44986 5973 44995
rect 6411 44986 6453 44995
rect 7563 44986 7605 44995
rect 7674 45035 7716 45044
rect 7674 44995 7675 45035
rect 7715 44995 7716 45035
rect 7674 44986 7716 44995
rect 7794 45035 7840 45044
rect 7794 44995 7795 45035
rect 7835 44995 7840 45035
rect 8235 45004 8236 45044
rect 8276 45004 8277 45044
rect 8235 44995 8277 45004
rect 8452 45044 8494 45053
rect 8452 45004 8453 45044
rect 8493 45004 8494 45044
rect 8452 44995 8494 45004
rect 8715 45044 8757 45053
rect 8715 45004 8716 45044
rect 8756 45004 8757 45044
rect 8715 44995 8757 45004
rect 8834 45044 8876 45053
rect 8834 45004 8835 45044
rect 8875 45004 8876 45044
rect 8834 44995 8876 45004
rect 8944 45044 9002 45045
rect 8944 45004 8953 45044
rect 8993 45004 9002 45044
rect 8944 45003 9002 45004
rect 9195 45044 9237 45053
rect 10810 45044 10868 45045
rect 11190 45044 11248 45045
rect 9195 45004 9196 45044
rect 9236 45004 9237 45044
rect 9195 44995 9237 45004
rect 10443 45035 10485 45044
rect 10443 44995 10444 45035
rect 10484 44995 10485 45035
rect 10810 45004 10819 45044
rect 10859 45004 10868 45044
rect 10810 45003 10868 45004
rect 10923 45035 10965 45044
rect 7794 44986 7840 44995
rect 10443 44986 10485 44995
rect 10923 44995 10924 45035
rect 10964 44995 10965 45035
rect 11190 45004 11199 45044
rect 11239 45004 11248 45044
rect 11190 45003 11248 45004
rect 11371 45044 11429 45045
rect 11371 45004 11380 45044
rect 11420 45004 11429 45044
rect 11371 45003 11429 45004
rect 13485 45044 13527 45053
rect 13485 45004 13486 45044
rect 13526 45004 13527 45044
rect 13485 44995 13527 45004
rect 13616 45044 13658 45053
rect 13616 45004 13617 45044
rect 13657 45004 13658 45044
rect 13616 44995 13658 45004
rect 13995 45044 14037 45053
rect 16011 45044 16053 45053
rect 18010 45044 18068 45045
rect 13995 45004 13996 45044
rect 14036 45004 14037 45044
rect 13995 44995 14037 45004
rect 14571 45035 14613 45044
rect 14571 44995 14572 45035
rect 14612 44995 14613 45035
rect 10923 44986 10965 44995
rect 14571 44986 14613 44995
rect 15051 45035 15093 45044
rect 15051 44995 15052 45035
rect 15092 44995 15093 45035
rect 16011 45004 16012 45044
rect 16052 45004 16053 45044
rect 16011 44995 16053 45004
rect 17259 45035 17301 45044
rect 17259 44995 17260 45035
rect 17300 44995 17301 45035
rect 18010 45004 18019 45044
rect 18059 45004 18068 45044
rect 18010 45003 18068 45004
rect 18123 45044 18165 45053
rect 18123 45004 18124 45044
rect 18164 45004 18165 45044
rect 18123 44995 18165 45004
rect 18507 45044 18549 45053
rect 18507 45004 18508 45044
rect 18548 45004 18549 45044
rect 18507 44995 18549 45004
rect 19083 45035 19125 45044
rect 19083 44995 19084 45035
rect 19124 44995 19125 45035
rect 15051 44986 15093 44995
rect 17259 44986 17301 44995
rect 19083 44986 19125 44995
rect 19563 45035 19605 45044
rect 19563 44995 19564 45035
rect 19604 44995 19605 45035
rect 19563 44986 19605 44995
rect 5296 44961 5354 44962
rect 1611 44920 1612 44960
rect 1652 44920 1653 44960
rect 1611 44911 1653 44920
rect 6891 44960 6933 44969
rect 8619 44960 8661 44969
rect 6891 44920 6892 44960
rect 6932 44920 6933 44960
rect 6891 44911 6933 44920
rect 8370 44951 8416 44960
rect 8370 44911 8371 44951
rect 8411 44911 8416 44951
rect 8619 44920 8620 44960
rect 8660 44920 8661 44960
rect 8619 44911 8661 44920
rect 11691 44960 11733 44969
rect 11691 44920 11692 44960
rect 11732 44920 11733 44960
rect 11691 44911 11733 44920
rect 12651 44960 12693 44969
rect 12651 44920 12652 44960
rect 12692 44920 12693 44960
rect 12651 44911 12693 44920
rect 14091 44960 14133 44969
rect 14091 44920 14092 44960
rect 14132 44920 14133 44960
rect 14091 44911 14133 44920
rect 15723 44960 15765 44969
rect 15723 44920 15724 44960
rect 15764 44920 15765 44960
rect 15723 44911 15765 44920
rect 18603 44960 18645 44969
rect 18603 44920 18604 44960
rect 18644 44920 18645 44960
rect 18603 44911 18645 44920
rect 20139 44960 20181 44969
rect 20139 44920 20140 44960
rect 20180 44920 20181 44960
rect 20139 44911 20181 44920
rect 8370 44902 8416 44911
rect 4203 44876 4245 44885
rect 4203 44836 4204 44876
rect 4244 44836 4245 44876
rect 4203 44827 4245 44836
rect 4875 44876 4917 44885
rect 4875 44836 4876 44876
rect 4916 44836 4917 44876
rect 4875 44827 4917 44836
rect 6987 44876 7029 44885
rect 6987 44836 6988 44876
rect 7028 44836 7029 44876
rect 6987 44827 7029 44836
rect 1467 44792 1509 44801
rect 1467 44752 1468 44792
rect 1508 44752 1509 44792
rect 1467 44743 1509 44752
rect 1851 44792 1893 44801
rect 1851 44752 1852 44792
rect 1892 44752 1893 44792
rect 1851 44743 1893 44752
rect 6106 44792 6164 44793
rect 6106 44752 6115 44792
rect 6155 44752 6164 44792
rect 6106 44751 6164 44752
rect 7947 44792 7989 44801
rect 7947 44752 7948 44792
rect 7988 44752 7989 44792
rect 7947 44743 7989 44752
rect 10810 44792 10868 44793
rect 10810 44752 10819 44792
rect 10859 44752 10868 44792
rect 10810 44751 10868 44752
rect 12411 44792 12453 44801
rect 12411 44752 12412 44792
rect 12452 44752 12453 44792
rect 12411 44743 12453 44752
rect 15483 44792 15525 44801
rect 15483 44752 15484 44792
rect 15524 44752 15525 44792
rect 15483 44743 15525 44752
rect 20379 44792 20421 44801
rect 20379 44752 20380 44792
rect 20420 44752 20421 44792
rect 20379 44743 20421 44752
rect 1152 44624 20448 44648
rect 1152 44584 3688 44624
rect 3728 44584 3770 44624
rect 3810 44584 3852 44624
rect 3892 44584 3934 44624
rect 3974 44584 4016 44624
rect 4056 44584 18808 44624
rect 18848 44584 18890 44624
rect 18930 44584 18972 44624
rect 19012 44584 19054 44624
rect 19094 44584 19136 44624
rect 19176 44584 20448 44624
rect 1152 44560 20448 44584
rect 1851 44456 1893 44465
rect 1851 44416 1852 44456
rect 1892 44416 1893 44456
rect 1851 44407 1893 44416
rect 4666 44456 4724 44457
rect 4666 44416 4675 44456
rect 4715 44416 4724 44456
rect 4666 44415 4724 44416
rect 5451 44456 5493 44465
rect 5451 44416 5452 44456
rect 5492 44416 5493 44456
rect 5451 44407 5493 44416
rect 6603 44456 6645 44465
rect 6603 44416 6604 44456
rect 6644 44416 6645 44456
rect 6603 44407 6645 44416
rect 6843 44456 6885 44465
rect 6843 44416 6844 44456
rect 6884 44416 6885 44456
rect 6843 44407 6885 44416
rect 7179 44456 7221 44465
rect 7179 44416 7180 44456
rect 7220 44416 7221 44456
rect 7179 44407 7221 44416
rect 11163 44456 11205 44465
rect 11163 44416 11164 44456
rect 11204 44416 11205 44456
rect 11163 44407 11205 44416
rect 13419 44456 13461 44465
rect 13419 44416 13420 44456
rect 13460 44416 13461 44456
rect 13419 44407 13461 44416
rect 15051 44456 15093 44465
rect 15051 44416 15052 44456
rect 15092 44416 15093 44456
rect 15051 44407 15093 44416
rect 17643 44456 17685 44465
rect 17643 44416 17644 44456
rect 17684 44416 17685 44456
rect 17643 44407 17685 44416
rect 18171 44456 18213 44465
rect 18171 44416 18172 44456
rect 18212 44416 18213 44456
rect 18171 44407 18213 44416
rect 20139 44456 20181 44465
rect 20139 44416 20140 44456
rect 20180 44416 20181 44456
rect 20139 44407 20181 44416
rect 1467 44372 1509 44381
rect 6123 44372 6165 44381
rect 1467 44332 1468 44372
rect 1508 44332 1509 44372
rect 1467 44323 1509 44332
rect 4459 44363 4501 44372
rect 4459 44323 4460 44363
rect 4500 44323 4501 44363
rect 6123 44332 6124 44372
rect 6164 44332 6165 44372
rect 6123 44323 6165 44332
rect 11547 44372 11589 44381
rect 11547 44332 11548 44372
rect 11588 44332 11589 44372
rect 11547 44323 11589 44332
rect 16011 44372 16053 44381
rect 16011 44332 16012 44372
rect 16052 44332 16053 44372
rect 16011 44323 16053 44332
rect 4459 44314 4501 44323
rect 1227 44288 1269 44297
rect 1227 44248 1228 44288
rect 1268 44248 1269 44288
rect 1227 44239 1269 44248
rect 1611 44288 1653 44297
rect 1611 44248 1612 44288
rect 1652 44248 1653 44288
rect 1611 44239 1653 44248
rect 2859 44288 2901 44297
rect 2859 44248 2860 44288
rect 2900 44248 2901 44288
rect 2859 44239 2901 44248
rect 6219 44288 6261 44297
rect 6219 44248 6220 44288
rect 6260 44248 6261 44288
rect 5470 44246 5528 44247
rect 5014 44237 5056 44246
rect 2362 44204 2420 44205
rect 2362 44164 2371 44204
rect 2411 44164 2420 44204
rect 2362 44163 2420 44164
rect 2475 44204 2517 44213
rect 2475 44164 2476 44204
rect 2516 44164 2517 44204
rect 2475 44155 2517 44164
rect 2955 44204 2997 44213
rect 2955 44164 2956 44204
rect 2996 44164 2997 44204
rect 2955 44155 2997 44164
rect 3427 44204 3485 44205
rect 3427 44164 3436 44204
rect 3476 44164 3485 44204
rect 3427 44163 3485 44164
rect 3915 44204 3973 44205
rect 3915 44164 3924 44204
rect 3964 44164 3973 44204
rect 3915 44163 3973 44164
rect 4474 44204 4532 44205
rect 4474 44164 4483 44204
rect 4523 44164 4532 44204
rect 4474 44163 4532 44164
rect 4906 44204 4964 44205
rect 4906 44164 4915 44204
rect 4955 44164 4964 44204
rect 5014 44197 5015 44237
rect 5055 44197 5056 44237
rect 5014 44188 5056 44197
rect 5355 44204 5397 44213
rect 5470 44206 5479 44246
rect 5519 44206 5528 44246
rect 5694 44237 5736 44246
rect 6219 44239 6261 44248
rect 9754 44288 9812 44289
rect 9754 44248 9763 44288
rect 9803 44248 9812 44288
rect 9754 44247 9812 44248
rect 10539 44288 10581 44297
rect 10539 44248 10540 44288
rect 10580 44248 10581 44288
rect 10539 44239 10581 44248
rect 11403 44288 11445 44297
rect 11403 44248 11404 44288
rect 11444 44248 11445 44288
rect 11403 44239 11445 44248
rect 11787 44288 11829 44297
rect 11787 44248 11788 44288
rect 11828 44248 11829 44288
rect 11787 44239 11829 44248
rect 17835 44288 17877 44297
rect 17835 44248 17836 44288
rect 17876 44248 17877 44288
rect 17835 44239 17877 44248
rect 18411 44288 18453 44297
rect 18411 44248 18412 44288
rect 18452 44248 18453 44288
rect 18411 44239 18453 44248
rect 5470 44205 5528 44206
rect 4906 44163 4964 44164
rect 5355 44164 5356 44204
rect 5396 44164 5397 44204
rect 5355 44155 5397 44164
rect 5592 44204 5634 44213
rect 5592 44164 5593 44204
rect 5633 44164 5634 44204
rect 5694 44197 5695 44237
rect 5735 44197 5736 44237
rect 5694 44188 5736 44197
rect 5883 44204 5925 44213
rect 5592 44155 5634 44164
rect 5883 44164 5884 44204
rect 5924 44164 5925 44204
rect 6340 44204 6382 44213
rect 5883 44155 5925 44164
rect 6055 44162 6097 44171
rect 6055 44122 6056 44162
rect 6096 44122 6097 44162
rect 6340 44164 6341 44204
rect 6381 44164 6382 44204
rect 6700 44204 6758 44205
rect 6340 44155 6382 44164
rect 6496 44177 6554 44178
rect 6496 44137 6505 44177
rect 6545 44137 6554 44177
rect 6700 44164 6709 44204
rect 6749 44164 6758 44204
rect 6700 44163 6758 44164
rect 6939 44204 6981 44213
rect 6939 44164 6940 44204
rect 6980 44164 6981 44204
rect 6939 44155 6981 44164
rect 7179 44204 7221 44213
rect 7179 44164 7180 44204
rect 7220 44164 7221 44204
rect 7179 44155 7221 44164
rect 7371 44204 7413 44213
rect 7371 44164 7372 44204
rect 7412 44164 7413 44204
rect 7371 44155 7413 44164
rect 7563 44204 7605 44213
rect 7563 44164 7564 44204
rect 7604 44164 7605 44204
rect 7563 44155 7605 44164
rect 8803 44204 8861 44205
rect 8803 44164 8812 44204
rect 8852 44164 8861 44204
rect 8803 44163 8861 44164
rect 9178 44204 9236 44205
rect 9178 44164 9187 44204
rect 9227 44164 9236 44204
rect 9178 44163 9236 44164
rect 9634 44204 9692 44205
rect 9634 44164 9643 44204
rect 9683 44164 9692 44204
rect 9634 44163 9692 44164
rect 9867 44204 9909 44213
rect 9867 44164 9868 44204
rect 9908 44164 9909 44204
rect 9867 44155 9909 44164
rect 11979 44204 12021 44213
rect 11979 44164 11980 44204
rect 12020 44164 12021 44204
rect 11979 44155 12021 44164
rect 13219 44204 13277 44205
rect 13219 44164 13228 44204
rect 13268 44164 13277 44204
rect 13219 44163 13277 44164
rect 13611 44204 13653 44213
rect 13611 44164 13612 44204
rect 13652 44164 13653 44204
rect 13611 44155 13653 44164
rect 14851 44204 14909 44205
rect 14851 44164 14860 44204
rect 14900 44164 14909 44204
rect 14851 44163 14909 44164
rect 15339 44204 15381 44213
rect 15339 44164 15340 44204
rect 15380 44164 15381 44204
rect 15339 44155 15381 44164
rect 15610 44204 15668 44205
rect 15610 44164 15619 44204
rect 15659 44164 15668 44204
rect 15610 44163 15668 44164
rect 16203 44204 16245 44213
rect 16203 44164 16204 44204
rect 16244 44164 16245 44204
rect 16203 44155 16245 44164
rect 17443 44204 17501 44205
rect 17443 44164 17452 44204
rect 17492 44164 17501 44204
rect 17443 44163 17501 44164
rect 18699 44204 18741 44213
rect 18699 44164 18700 44204
rect 18740 44164 18741 44204
rect 18699 44155 18741 44164
rect 19939 44204 19997 44205
rect 19939 44164 19948 44204
rect 19988 44164 19997 44204
rect 19939 44163 19997 44164
rect 6496 44136 6554 44137
rect 6055 44113 6097 44122
rect 9387 44120 9429 44129
rect 9387 44080 9388 44120
rect 9428 44080 9429 44120
rect 9387 44071 9429 44080
rect 9497 44120 9539 44129
rect 9497 44080 9498 44120
rect 9538 44080 9539 44120
rect 9497 44071 9539 44080
rect 11163 44120 11205 44129
rect 11163 44080 11164 44120
rect 11204 44080 11205 44120
rect 11163 44071 11205 44080
rect 15723 44120 15765 44129
rect 15723 44080 15724 44120
rect 15764 44080 15765 44120
rect 15723 44071 15765 44080
rect 4107 44036 4149 44045
rect 4107 43996 4108 44036
rect 4148 43996 4149 44036
rect 4107 43987 4149 43996
rect 5163 44036 5205 44045
rect 5163 43996 5164 44036
rect 5204 43996 5205 44036
rect 5163 43987 5205 43996
rect 9003 44036 9045 44045
rect 9003 43996 9004 44036
rect 9044 43996 9045 44036
rect 9003 43987 9045 43996
rect 9274 44036 9332 44037
rect 9274 43996 9283 44036
rect 9323 43996 9332 44036
rect 9274 43995 9332 43996
rect 9946 44036 10004 44037
rect 9946 43996 9955 44036
rect 9995 43996 10004 44036
rect 9946 43995 10004 43996
rect 10299 44036 10341 44045
rect 10299 43996 10300 44036
rect 10340 43996 10341 44036
rect 10299 43987 10341 43996
rect 18075 44036 18117 44045
rect 18075 43996 18076 44036
rect 18116 43996 18117 44036
rect 18075 43987 18117 43996
rect 1152 43868 20452 43892
rect 1152 43828 4928 43868
rect 4968 43828 5010 43868
rect 5050 43828 5092 43868
rect 5132 43828 5174 43868
rect 5214 43828 5256 43868
rect 5296 43828 20048 43868
rect 20088 43828 20130 43868
rect 20170 43828 20212 43868
rect 20252 43828 20294 43868
rect 20334 43828 20376 43868
rect 20416 43828 20452 43868
rect 1152 43804 20452 43828
rect 1467 43700 1509 43709
rect 1467 43660 1468 43700
rect 1508 43660 1509 43700
rect 1467 43651 1509 43660
rect 3915 43700 3957 43709
rect 3915 43660 3916 43700
rect 3956 43660 3957 43700
rect 3915 43651 3957 43660
rect 5067 43700 5109 43709
rect 5067 43660 5068 43700
rect 5108 43660 5109 43700
rect 5067 43651 5109 43660
rect 5914 43700 5972 43701
rect 5914 43660 5923 43700
rect 5963 43660 5972 43700
rect 5914 43659 5972 43660
rect 8235 43700 8277 43709
rect 8235 43660 8236 43700
rect 8276 43660 8277 43700
rect 8235 43651 8277 43660
rect 10347 43700 10389 43709
rect 10347 43660 10348 43700
rect 10388 43660 10389 43700
rect 10347 43651 10389 43660
rect 12651 43700 12693 43709
rect 12651 43660 12652 43700
rect 12692 43660 12693 43700
rect 12651 43651 12693 43660
rect 13083 43700 13125 43709
rect 13083 43660 13084 43700
rect 13124 43660 13125 43700
rect 13083 43651 13125 43660
rect 16155 43700 16197 43709
rect 16155 43660 16156 43700
rect 16196 43660 16197 43700
rect 16155 43651 16197 43660
rect 19755 43700 19797 43709
rect 19755 43660 19756 43700
rect 19796 43660 19797 43700
rect 19755 43651 19797 43660
rect 20379 43700 20421 43709
rect 20379 43660 20380 43700
rect 20420 43660 20421 43700
rect 20379 43651 20421 43660
rect 5824 43616 5866 43625
rect 5824 43576 5825 43616
rect 5865 43576 5866 43616
rect 5824 43567 5866 43576
rect 14331 43616 14373 43625
rect 14331 43576 14332 43616
rect 14372 43576 14373 43616
rect 14331 43567 14373 43576
rect 15435 43616 15477 43625
rect 15435 43576 15436 43616
rect 15476 43576 15477 43616
rect 15435 43567 15477 43576
rect 17739 43616 17781 43625
rect 17739 43576 17740 43616
rect 17780 43576 17781 43616
rect 17739 43567 17781 43576
rect 2475 43532 2517 43541
rect 4585 43532 4627 43541
rect 2475 43492 2476 43532
rect 2516 43492 2517 43532
rect 2475 43483 2517 43492
rect 3723 43523 3765 43532
rect 3723 43483 3724 43523
rect 3764 43483 3765 43523
rect 3723 43474 3765 43483
rect 4347 43490 4389 43499
rect 1227 43448 1269 43457
rect 1227 43408 1228 43448
rect 1268 43408 1269 43448
rect 1227 43399 1269 43408
rect 1611 43448 1653 43457
rect 1611 43408 1612 43448
rect 1652 43408 1653 43448
rect 1611 43399 1653 43408
rect 2091 43448 2133 43457
rect 2091 43408 2092 43448
rect 2132 43408 2133 43448
rect 4347 43450 4348 43490
rect 4388 43450 4389 43490
rect 4585 43492 4586 43532
rect 4626 43492 4627 43532
rect 4585 43483 4627 43492
rect 4858 43532 4916 43533
rect 4858 43492 4867 43532
rect 4907 43492 4916 43532
rect 4858 43491 4916 43492
rect 5163 43532 5205 43541
rect 5163 43492 5164 43532
rect 5204 43492 5205 43532
rect 5163 43483 5205 43492
rect 5398 43532 5440 43541
rect 5398 43492 5399 43532
rect 5439 43492 5440 43532
rect 5398 43483 5440 43492
rect 5499 43532 5541 43541
rect 5499 43492 5500 43532
rect 5540 43492 5541 43532
rect 5499 43483 5541 43492
rect 5643 43532 5685 43541
rect 5643 43492 5644 43532
rect 5684 43492 5685 43532
rect 5643 43483 5685 43492
rect 6027 43532 6069 43541
rect 6490 43532 6548 43533
rect 6027 43492 6028 43532
rect 6068 43492 6069 43532
rect 6027 43483 6069 43492
rect 6123 43523 6165 43532
rect 6123 43483 6124 43523
rect 6164 43483 6165 43523
rect 6490 43492 6499 43532
rect 6539 43492 6548 43532
rect 6490 43491 6548 43492
rect 6603 43532 6645 43541
rect 6603 43492 6604 43532
rect 6644 43492 6645 43532
rect 6603 43483 6645 43492
rect 6987 43532 7029 43541
rect 8907 43532 8949 43541
rect 10906 43532 10964 43533
rect 6987 43492 6988 43532
rect 7028 43492 7029 43532
rect 6987 43483 7029 43492
rect 7563 43523 7605 43532
rect 7563 43483 7564 43523
rect 7604 43483 7605 43523
rect 6123 43474 6165 43483
rect 7563 43474 7605 43483
rect 8043 43523 8085 43532
rect 8043 43483 8044 43523
rect 8084 43483 8085 43523
rect 8907 43492 8908 43532
rect 8948 43492 8949 43532
rect 8907 43483 8949 43492
rect 10155 43523 10197 43532
rect 10155 43483 10156 43523
rect 10196 43483 10197 43523
rect 10906 43492 10915 43532
rect 10955 43492 10964 43532
rect 10906 43491 10964 43492
rect 11019 43532 11061 43541
rect 11019 43492 11020 43532
rect 11060 43492 11061 43532
rect 11019 43483 11061 43492
rect 11403 43532 11445 43541
rect 14187 43532 14229 43541
rect 11403 43492 11404 43532
rect 11444 43492 11445 43532
rect 11403 43483 11445 43492
rect 11979 43523 12021 43532
rect 11979 43483 11980 43523
rect 12020 43483 12021 43523
rect 8043 43474 8085 43483
rect 10155 43474 10197 43483
rect 11979 43474 12021 43483
rect 12459 43523 12501 43532
rect 12459 43483 12460 43523
rect 12500 43483 12501 43523
rect 14187 43492 14188 43532
rect 14228 43492 14229 43532
rect 14187 43483 14229 43492
rect 14571 43532 14613 43541
rect 14571 43492 14572 43532
rect 14612 43492 14613 43532
rect 14571 43483 14613 43492
rect 14800 43532 14858 43533
rect 14800 43492 14809 43532
rect 14849 43492 14858 43532
rect 14800 43491 14858 43492
rect 15051 43532 15093 43541
rect 15051 43492 15052 43532
rect 15092 43492 15093 43532
rect 15051 43483 15093 43492
rect 15322 43532 15380 43533
rect 15322 43492 15331 43532
rect 15371 43492 15380 43532
rect 15322 43491 15380 43492
rect 16299 43532 16341 43541
rect 18010 43532 18068 43533
rect 16299 43492 16300 43532
rect 16340 43492 16341 43532
rect 16299 43483 16341 43492
rect 17547 43523 17589 43532
rect 17547 43483 17548 43523
rect 17588 43483 17589 43523
rect 18010 43492 18019 43532
rect 18059 43492 18068 43532
rect 18010 43491 18068 43492
rect 18123 43532 18165 43541
rect 18123 43492 18124 43532
rect 18164 43492 18165 43532
rect 18123 43483 18165 43492
rect 18507 43532 18549 43541
rect 18507 43492 18508 43532
rect 18548 43492 18549 43532
rect 18507 43483 18549 43492
rect 19083 43523 19125 43532
rect 19083 43483 19084 43523
rect 19124 43483 19125 43523
rect 12459 43474 12501 43483
rect 17547 43474 17589 43483
rect 19083 43474 19125 43483
rect 19563 43523 19605 43532
rect 19563 43483 19564 43523
rect 19604 43483 19605 43523
rect 19563 43474 19605 43483
rect 4347 43441 4389 43450
rect 4474 43448 4532 43449
rect 2091 43399 2133 43408
rect 4474 43408 4483 43448
rect 4523 43408 4532 43448
rect 4474 43407 4532 43408
rect 4683 43448 4725 43457
rect 4683 43408 4684 43448
rect 4724 43408 4725 43448
rect 4683 43399 4725 43408
rect 7083 43448 7125 43457
rect 7083 43408 7084 43448
rect 7124 43408 7125 43448
rect 7083 43399 7125 43408
rect 11499 43448 11541 43457
rect 11499 43408 11500 43448
rect 11540 43408 11541 43448
rect 11499 43399 11541 43408
rect 12843 43448 12885 43457
rect 12843 43408 12844 43448
rect 12884 43408 12885 43448
rect 12843 43399 12885 43408
rect 13419 43448 13461 43457
rect 13419 43408 13420 43448
rect 13460 43408 13461 43448
rect 13419 43399 13461 43408
rect 14475 43448 14517 43457
rect 14475 43408 14476 43448
rect 14516 43408 14517 43448
rect 14475 43399 14517 43408
rect 14690 43448 14732 43457
rect 14690 43408 14691 43448
rect 14731 43408 14732 43448
rect 14690 43399 14732 43408
rect 15915 43448 15957 43457
rect 15915 43408 15916 43448
rect 15956 43408 15957 43448
rect 15915 43399 15957 43408
rect 18603 43448 18645 43457
rect 18603 43408 18604 43448
rect 18644 43408 18645 43448
rect 18603 43399 18645 43408
rect 20139 43448 20181 43457
rect 20139 43408 20140 43448
rect 20180 43408 20181 43448
rect 20139 43399 20181 43408
rect 2331 43364 2373 43373
rect 2331 43324 2332 43364
rect 2372 43324 2373 43364
rect 2331 43315 2373 43324
rect 13179 43364 13221 43373
rect 13179 43324 13180 43364
rect 13220 43324 13221 43364
rect 13179 43315 13221 43324
rect 15723 43364 15765 43373
rect 15723 43324 15724 43364
rect 15764 43324 15765 43364
rect 15723 43315 15765 43324
rect 1851 43280 1893 43289
rect 1851 43240 1852 43280
rect 1892 43240 1893 43280
rect 1851 43231 1893 43240
rect 5355 43280 5397 43289
rect 5355 43240 5356 43280
rect 5396 43240 5397 43280
rect 5355 43231 5397 43240
rect 1152 43112 20448 43136
rect 1152 43072 3688 43112
rect 3728 43072 3770 43112
rect 3810 43072 3852 43112
rect 3892 43072 3934 43112
rect 3974 43072 4016 43112
rect 4056 43072 18808 43112
rect 18848 43072 18890 43112
rect 18930 43072 18972 43112
rect 19012 43072 19054 43112
rect 19094 43072 19136 43112
rect 19176 43072 20448 43112
rect 1152 43048 20448 43072
rect 4587 42944 4629 42953
rect 4587 42904 4588 42944
rect 4628 42904 4629 42944
rect 4587 42895 4629 42904
rect 5338 42944 5396 42945
rect 5338 42904 5347 42944
rect 5387 42904 5396 42944
rect 5338 42903 5396 42904
rect 5931 42944 5973 42953
rect 5931 42904 5932 42944
rect 5972 42904 5973 42944
rect 5931 42895 5973 42904
rect 9003 42944 9045 42953
rect 9003 42904 9004 42944
rect 9044 42904 9045 42944
rect 9003 42895 9045 42904
rect 12891 42944 12933 42953
rect 12891 42904 12892 42944
rect 12932 42904 12933 42944
rect 12891 42895 12933 42904
rect 20379 42944 20421 42953
rect 20379 42904 20380 42944
rect 20420 42904 20421 42944
rect 20379 42895 20421 42904
rect 2235 42860 2277 42869
rect 2235 42820 2236 42860
rect 2276 42820 2277 42860
rect 2235 42811 2277 42820
rect 4011 42860 4053 42869
rect 4011 42820 4012 42860
rect 4052 42820 4053 42860
rect 4011 42811 4053 42820
rect 5163 42860 5205 42869
rect 5163 42820 5164 42860
rect 5204 42820 5205 42860
rect 5163 42811 5205 42820
rect 1227 42776 1269 42785
rect 1227 42736 1228 42776
rect 1268 42736 1269 42776
rect 1227 42727 1269 42736
rect 1611 42776 1653 42785
rect 1611 42736 1612 42776
rect 1652 42736 1653 42776
rect 1611 42727 1653 42736
rect 1995 42776 2037 42785
rect 1995 42736 1996 42776
rect 2036 42736 2037 42776
rect 1995 42727 2037 42736
rect 6795 42776 6837 42785
rect 6795 42736 6796 42776
rect 6836 42736 6837 42776
rect 6795 42727 6837 42736
rect 13131 42776 13173 42785
rect 13131 42736 13132 42776
rect 13172 42736 13173 42776
rect 13131 42727 13173 42736
rect 15514 42776 15572 42777
rect 15514 42736 15523 42776
rect 15563 42736 15572 42776
rect 15514 42735 15572 42736
rect 18507 42776 18549 42785
rect 18507 42736 18508 42776
rect 18548 42736 18549 42776
rect 18507 42727 18549 42736
rect 20139 42776 20181 42785
rect 20139 42736 20140 42776
rect 20180 42736 20181 42776
rect 20139 42727 20181 42736
rect 2571 42692 2613 42701
rect 2571 42652 2572 42692
rect 2612 42652 2613 42692
rect 2571 42643 2613 42652
rect 3811 42692 3869 42693
rect 3811 42652 3820 42692
rect 3860 42652 3869 42692
rect 3811 42651 3869 42652
rect 4203 42692 4245 42701
rect 4203 42652 4204 42692
rect 4244 42652 4245 42692
rect 4203 42643 4245 42652
rect 4491 42692 4533 42701
rect 4491 42652 4492 42692
rect 4532 42652 4533 42692
rect 4491 42643 4533 42652
rect 4683 42692 4725 42701
rect 4683 42652 4684 42692
rect 4724 42652 4725 42692
rect 4683 42643 4725 42652
rect 4971 42692 5013 42701
rect 4971 42652 4972 42692
rect 5012 42652 5013 42692
rect 4971 42643 5013 42652
rect 5344 42692 5386 42701
rect 5344 42652 5345 42692
rect 5385 42652 5386 42692
rect 5344 42643 5386 42652
rect 5635 42692 5693 42693
rect 5635 42652 5644 42692
rect 5684 42652 5693 42692
rect 5635 42651 5693 42652
rect 5835 42692 5877 42701
rect 5835 42652 5836 42692
rect 5876 42652 5877 42692
rect 5835 42643 5877 42652
rect 6027 42692 6069 42701
rect 6027 42652 6028 42692
rect 6068 42652 6069 42692
rect 6027 42643 6069 42652
rect 6298 42692 6356 42693
rect 6298 42652 6307 42692
rect 6347 42652 6356 42692
rect 6298 42651 6356 42652
rect 6411 42692 6453 42701
rect 6411 42652 6412 42692
rect 6452 42652 6453 42692
rect 6411 42643 6453 42652
rect 6891 42692 6933 42701
rect 6891 42652 6892 42692
rect 6932 42652 6933 42692
rect 6891 42643 6933 42652
rect 7363 42692 7421 42693
rect 7363 42652 7372 42692
rect 7412 42652 7421 42692
rect 7363 42651 7421 42652
rect 7882 42692 7940 42693
rect 7882 42652 7891 42692
rect 7931 42652 7940 42692
rect 7882 42651 7940 42652
rect 8331 42692 8373 42701
rect 8331 42652 8332 42692
rect 8372 42652 8373 42692
rect 8331 42643 8373 42652
rect 8578 42692 8636 42693
rect 8578 42652 8587 42692
rect 8627 42652 8636 42692
rect 8578 42651 8636 42652
rect 8698 42692 8756 42693
rect 8698 42652 8707 42692
rect 8747 42652 8756 42692
rect 8698 42651 8756 42652
rect 9675 42692 9717 42701
rect 9675 42652 9676 42692
rect 9716 42652 9717 42692
rect 9675 42643 9717 42652
rect 10915 42692 10973 42693
rect 10915 42652 10924 42692
rect 10964 42652 10973 42692
rect 10915 42651 10973 42652
rect 11307 42692 11349 42701
rect 11307 42652 11308 42692
rect 11348 42652 11349 42692
rect 11307 42643 11349 42652
rect 12547 42692 12605 42693
rect 12547 42652 12556 42692
rect 12596 42652 12605 42692
rect 12547 42651 12605 42652
rect 13306 42692 13364 42693
rect 13306 42652 13315 42692
rect 13355 42652 13364 42692
rect 13306 42651 13364 42652
rect 13803 42692 13845 42701
rect 13803 42652 13804 42692
rect 13844 42652 13845 42692
rect 13803 42643 13845 42652
rect 15043 42692 15101 42693
rect 15043 42652 15052 42692
rect 15092 42652 15101 42692
rect 15043 42651 15101 42652
rect 15382 42692 15424 42701
rect 15382 42652 15383 42692
rect 15423 42652 15424 42692
rect 15382 42643 15424 42652
rect 15627 42692 15669 42701
rect 15627 42652 15628 42692
rect 15668 42652 15669 42692
rect 15627 42643 15669 42652
rect 15915 42692 15957 42701
rect 15915 42652 15916 42692
rect 15956 42652 15957 42692
rect 15915 42643 15957 42652
rect 16107 42692 16149 42701
rect 16107 42652 16108 42692
rect 16148 42652 16149 42692
rect 16107 42643 16149 42652
rect 16299 42692 16341 42701
rect 16299 42652 16300 42692
rect 16340 42652 16341 42692
rect 16299 42643 16341 42652
rect 17539 42692 17597 42693
rect 17539 42652 17548 42692
rect 17588 42652 17597 42692
rect 17539 42651 17597 42652
rect 18010 42692 18068 42693
rect 18010 42652 18019 42692
rect 18059 42652 18068 42692
rect 18010 42651 18068 42652
rect 18123 42692 18165 42701
rect 18123 42652 18124 42692
rect 18164 42652 18165 42692
rect 18123 42643 18165 42652
rect 18603 42692 18645 42701
rect 18603 42652 18604 42692
rect 18644 42652 18645 42692
rect 18603 42643 18645 42652
rect 19075 42692 19133 42693
rect 19075 42652 19084 42692
rect 19124 42652 19133 42692
rect 19075 42651 19133 42652
rect 19563 42692 19621 42693
rect 19563 42652 19572 42692
rect 19612 42652 19621 42692
rect 19563 42651 19621 42652
rect 1851 42608 1893 42617
rect 1851 42568 1852 42608
rect 1892 42568 1893 42608
rect 1851 42559 1893 42568
rect 12747 42608 12789 42617
rect 12747 42568 12748 42608
rect 12788 42568 12789 42608
rect 12747 42559 12789 42568
rect 13625 42608 13667 42617
rect 13625 42568 13626 42608
rect 13666 42568 13667 42608
rect 13625 42559 13667 42568
rect 17739 42608 17781 42617
rect 17739 42568 17740 42608
rect 17780 42568 17781 42608
rect 17739 42559 17781 42568
rect 1467 42524 1509 42533
rect 1467 42484 1468 42524
rect 1508 42484 1509 42524
rect 1467 42475 1509 42484
rect 4347 42524 4389 42533
rect 4347 42484 4348 42524
rect 4388 42484 4389 42524
rect 4347 42475 4389 42484
rect 4858 42524 4916 42525
rect 4858 42484 4867 42524
rect 4907 42484 4916 42524
rect 4858 42483 4916 42484
rect 5547 42524 5589 42533
rect 5547 42484 5548 42524
rect 5588 42484 5589 42524
rect 5547 42475 5589 42484
rect 8043 42524 8085 42533
rect 8043 42484 8044 42524
rect 8084 42484 8085 42524
rect 8043 42475 8085 42484
rect 11115 42524 11157 42533
rect 11115 42484 11116 42524
rect 11156 42484 11157 42524
rect 11115 42475 11157 42484
rect 13402 42524 13460 42525
rect 13402 42484 13411 42524
rect 13451 42484 13460 42524
rect 13402 42483 13460 42484
rect 13515 42524 13557 42533
rect 13515 42484 13516 42524
rect 13556 42484 13557 42524
rect 13515 42475 13557 42484
rect 15243 42524 15285 42533
rect 15243 42484 15244 42524
rect 15284 42484 15285 42524
rect 15243 42475 15285 42484
rect 15706 42524 15764 42525
rect 15706 42484 15715 42524
rect 15755 42484 15764 42524
rect 15706 42483 15764 42484
rect 16011 42524 16053 42533
rect 16011 42484 16012 42524
rect 16052 42484 16053 42524
rect 16011 42475 16053 42484
rect 19755 42524 19797 42533
rect 19755 42484 19756 42524
rect 19796 42484 19797 42524
rect 19755 42475 19797 42484
rect 1152 42356 20452 42380
rect 1152 42316 4928 42356
rect 4968 42316 5010 42356
rect 5050 42316 5092 42356
rect 5132 42316 5174 42356
rect 5214 42316 5256 42356
rect 5296 42316 20048 42356
rect 20088 42316 20130 42356
rect 20170 42316 20212 42356
rect 20252 42316 20294 42356
rect 20334 42316 20376 42356
rect 20416 42316 20452 42356
rect 1152 42292 20452 42316
rect 3291 42188 3333 42197
rect 3291 42148 3292 42188
rect 3332 42148 3333 42188
rect 3291 42139 3333 42148
rect 6987 42188 7029 42197
rect 6987 42148 6988 42188
rect 7028 42148 7029 42188
rect 6987 42139 7029 42148
rect 9099 42188 9141 42197
rect 9099 42148 9100 42188
rect 9140 42148 9141 42188
rect 9099 42139 9141 42148
rect 10731 42188 10773 42197
rect 10731 42148 10732 42188
rect 10772 42148 10773 42188
rect 10731 42139 10773 42148
rect 13227 42188 13269 42197
rect 13227 42148 13228 42188
rect 13268 42148 13269 42188
rect 13227 42139 13269 42148
rect 15051 42188 15093 42197
rect 15051 42148 15052 42188
rect 15092 42148 15093 42188
rect 15051 42139 15093 42148
rect 16203 42188 16245 42197
rect 16203 42148 16204 42188
rect 16244 42148 16245 42188
rect 16203 42139 16245 42148
rect 18027 42188 18069 42197
rect 18027 42148 18028 42188
rect 18068 42148 18069 42188
rect 18027 42139 18069 42148
rect 19659 42188 19701 42197
rect 19659 42148 19660 42188
rect 19700 42148 19701 42188
rect 19659 42139 19701 42148
rect 20379 42188 20421 42197
rect 20379 42148 20380 42188
rect 20420 42148 20421 42188
rect 20379 42139 20421 42148
rect 2859 42104 2901 42113
rect 2859 42064 2860 42104
rect 2900 42064 2901 42104
rect 2859 42055 2901 42064
rect 4971 42104 5013 42113
rect 4971 42064 4972 42104
rect 5012 42064 5013 42104
rect 4971 42055 5013 42064
rect 16000 42104 16042 42113
rect 16000 42064 16001 42104
rect 16041 42064 16042 42104
rect 16000 42055 16042 42064
rect 1419 42020 1461 42029
rect 3531 42020 3573 42029
rect 5242 42020 5300 42021
rect 1419 41980 1420 42020
rect 1460 41980 1461 42020
rect 1419 41971 1461 41980
rect 2667 42011 2709 42020
rect 2667 41971 2668 42011
rect 2708 41971 2709 42011
rect 3531 41980 3532 42020
rect 3572 41980 3573 42020
rect 3531 41971 3573 41980
rect 4779 42011 4821 42020
rect 4779 41971 4780 42011
rect 4820 41971 4821 42011
rect 5242 41980 5251 42020
rect 5291 41980 5300 42020
rect 5242 41979 5300 41980
rect 5355 42020 5397 42029
rect 5355 41980 5356 42020
rect 5396 41980 5397 42020
rect 5355 41971 5397 41980
rect 5739 42020 5781 42029
rect 7659 42020 7701 42029
rect 9291 42020 9333 42029
rect 11482 42020 11540 42021
rect 5739 41980 5740 42020
rect 5780 41980 5781 42020
rect 5739 41971 5781 41980
rect 6315 42011 6357 42020
rect 6315 41971 6316 42011
rect 6356 41971 6357 42011
rect 2667 41962 2709 41971
rect 4779 41962 4821 41971
rect 6315 41962 6357 41971
rect 6795 42011 6837 42020
rect 6795 41971 6796 42011
rect 6836 41971 6837 42011
rect 7659 41980 7660 42020
rect 7700 41980 7701 42020
rect 7659 41971 7701 41980
rect 8907 42011 8949 42020
rect 8907 41971 8908 42011
rect 8948 41971 8949 42011
rect 9291 41980 9292 42020
rect 9332 41980 9333 42020
rect 9291 41971 9333 41980
rect 10539 42011 10581 42020
rect 10539 41971 10540 42011
rect 10580 41971 10581 42011
rect 11482 41980 11491 42020
rect 11531 41980 11540 42020
rect 11482 41979 11540 41980
rect 11595 42020 11637 42029
rect 11595 41980 11596 42020
rect 11636 41980 11637 42020
rect 11595 41971 11637 41980
rect 11979 42020 12021 42029
rect 13419 42020 13461 42029
rect 15147 42020 15189 42029
rect 15376 42020 15434 42021
rect 11979 41980 11980 42020
rect 12020 41980 12021 42020
rect 11979 41971 12021 41980
rect 12555 42011 12597 42020
rect 12555 41971 12556 42011
rect 12596 41971 12597 42011
rect 6795 41962 6837 41971
rect 8907 41962 8949 41971
rect 10539 41962 10581 41971
rect 12555 41962 12597 41971
rect 13035 42011 13077 42020
rect 13035 41971 13036 42011
rect 13076 41971 13077 42011
rect 13419 41980 13420 42020
rect 13460 41980 13461 42020
rect 13419 41971 13461 41980
rect 14667 42011 14709 42020
rect 14667 41971 14668 42011
rect 14708 41971 14709 42011
rect 15147 41980 15148 42020
rect 15188 41980 15189 42020
rect 15147 41971 15189 41980
rect 15282 42011 15328 42020
rect 15282 41971 15283 42011
rect 15323 41971 15328 42011
rect 15376 41980 15385 42020
rect 15425 41980 15434 42020
rect 15376 41979 15434 41980
rect 15626 42020 15668 42029
rect 15626 41980 15627 42020
rect 15667 41980 15668 42020
rect 15626 41971 15668 41980
rect 15844 42020 15886 42029
rect 16587 42020 16629 42029
rect 18219 42020 18261 42029
rect 15844 41980 15845 42020
rect 15885 41980 15886 42020
rect 15844 41971 15886 41980
rect 16301 42011 16343 42020
rect 16301 41971 16302 42011
rect 16342 41971 16343 42011
rect 16587 41980 16588 42020
rect 16628 41980 16629 42020
rect 16587 41971 16629 41980
rect 17835 42011 17877 42020
rect 17835 41971 17836 42011
rect 17876 41971 17877 42011
rect 18219 41980 18220 42020
rect 18260 41980 18261 42020
rect 18219 41971 18261 41980
rect 19467 42011 19509 42020
rect 19467 41971 19468 42011
rect 19508 41971 19509 42011
rect 13035 41962 13077 41971
rect 14667 41962 14709 41971
rect 15282 41962 15328 41971
rect 16301 41962 16343 41971
rect 17835 41962 17877 41971
rect 19467 41962 19509 41971
rect 3051 41936 3093 41945
rect 3051 41896 3052 41936
rect 3092 41896 3093 41936
rect 3051 41887 3093 41896
rect 5835 41936 5877 41945
rect 5835 41896 5836 41936
rect 5876 41896 5877 41936
rect 5835 41887 5877 41896
rect 12075 41936 12117 41945
rect 12075 41896 12076 41936
rect 12116 41896 12117 41936
rect 12075 41887 12117 41896
rect 15531 41936 15573 41945
rect 20139 41936 20181 41945
rect 15531 41896 15532 41936
rect 15572 41896 15573 41936
rect 15531 41887 15573 41896
rect 15762 41927 15808 41936
rect 15762 41887 15763 41927
rect 15803 41887 15808 41927
rect 20139 41896 20140 41936
rect 20180 41896 20181 41936
rect 20139 41887 20181 41896
rect 15762 41878 15808 41887
rect 14859 41768 14901 41777
rect 14859 41728 14860 41768
rect 14900 41728 14901 41768
rect 14859 41719 14901 41728
rect 15994 41768 16052 41769
rect 15994 41728 16003 41768
rect 16043 41728 16052 41768
rect 15994 41727 16052 41728
rect 1152 41600 20448 41624
rect 1152 41560 3688 41600
rect 3728 41560 3770 41600
rect 3810 41560 3852 41600
rect 3892 41560 3934 41600
rect 3974 41560 4016 41600
rect 4056 41560 18808 41600
rect 18848 41560 18890 41600
rect 18930 41560 18972 41600
rect 19012 41560 19054 41600
rect 19094 41560 19136 41600
rect 19176 41560 20448 41600
rect 1152 41536 20448 41560
rect 2667 41432 2709 41441
rect 2667 41392 2668 41432
rect 2708 41392 2709 41432
rect 2667 41383 2709 41392
rect 4539 41432 4581 41441
rect 4539 41392 4540 41432
rect 4580 41392 4581 41432
rect 4539 41383 4581 41392
rect 8907 41432 8949 41441
rect 8907 41392 8908 41432
rect 8948 41392 8949 41432
rect 8907 41383 8949 41392
rect 10539 41432 10581 41441
rect 10539 41392 10540 41432
rect 10580 41392 10581 41432
rect 10539 41383 10581 41392
rect 15610 41432 15668 41433
rect 15610 41392 15619 41432
rect 15659 41392 15668 41432
rect 15610 41391 15668 41392
rect 16251 41432 16293 41441
rect 16251 41392 16252 41432
rect 16292 41392 16293 41432
rect 16251 41383 16293 41392
rect 15147 41348 15189 41357
rect 15147 41308 15148 41348
rect 15188 41308 15189 41348
rect 15147 41299 15189 41308
rect 20379 41348 20421 41357
rect 20379 41308 20380 41348
rect 20420 41308 20421 41348
rect 20379 41299 20421 41308
rect 4779 41264 4821 41273
rect 4779 41224 4780 41264
rect 4820 41224 4821 41264
rect 4779 41215 4821 41224
rect 11307 41264 11349 41273
rect 11307 41224 11308 41264
rect 11348 41224 11349 41264
rect 11307 41215 11349 41224
rect 15291 41264 15333 41273
rect 15291 41224 15292 41264
rect 15332 41224 15333 41264
rect 15291 41215 15333 41224
rect 18603 41264 18645 41273
rect 18603 41224 18604 41264
rect 18644 41224 18645 41264
rect 18603 41215 18645 41224
rect 20139 41264 20181 41273
rect 20139 41224 20140 41264
rect 20180 41224 20181 41264
rect 20139 41215 20181 41224
rect 1227 41180 1269 41189
rect 1227 41140 1228 41180
rect 1268 41140 1269 41180
rect 1227 41131 1269 41140
rect 2467 41180 2525 41181
rect 2467 41140 2476 41180
rect 2516 41140 2525 41180
rect 2467 41139 2525 41140
rect 2859 41180 2901 41189
rect 2859 41140 2860 41180
rect 2900 41140 2901 41180
rect 2859 41131 2901 41140
rect 4099 41180 4157 41181
rect 4099 41140 4108 41180
rect 4148 41140 4157 41180
rect 4099 41139 4157 41140
rect 5163 41180 5205 41189
rect 5163 41140 5164 41180
rect 5204 41140 5205 41180
rect 5163 41131 5205 41140
rect 5355 41180 5397 41189
rect 5355 41140 5356 41180
rect 5396 41140 5397 41180
rect 5355 41131 5397 41140
rect 5547 41180 5589 41189
rect 5547 41140 5548 41180
rect 5588 41140 5589 41180
rect 5547 41131 5589 41140
rect 5686 41180 5728 41189
rect 5686 41140 5687 41180
rect 5727 41140 5728 41180
rect 5686 41131 5728 41140
rect 6010 41180 6068 41181
rect 6010 41140 6019 41180
rect 6059 41140 6068 41180
rect 6010 41139 6068 41140
rect 6315 41180 6357 41189
rect 6315 41140 6316 41180
rect 6356 41140 6357 41180
rect 6315 41131 6357 41140
rect 6496 41180 6538 41189
rect 6496 41140 6497 41180
rect 6537 41140 6538 41180
rect 6496 41131 6538 41140
rect 6787 41180 6845 41181
rect 6787 41140 6796 41180
rect 6836 41140 6845 41180
rect 6787 41139 6845 41140
rect 7083 41180 7125 41189
rect 7083 41140 7084 41180
rect 7124 41140 7125 41180
rect 7083 41131 7125 41140
rect 7467 41180 7509 41189
rect 7467 41140 7468 41180
rect 7508 41140 7509 41180
rect 7467 41131 7509 41140
rect 8707 41180 8765 41181
rect 8707 41140 8716 41180
rect 8756 41140 8765 41180
rect 8707 41139 8765 41140
rect 9099 41180 9141 41189
rect 9099 41140 9100 41180
rect 9140 41140 9141 41180
rect 9099 41131 9141 41140
rect 10339 41180 10397 41181
rect 10339 41140 10348 41180
rect 10388 41140 10397 41180
rect 10339 41139 10397 41140
rect 10797 41180 10839 41189
rect 10797 41140 10798 41180
rect 10838 41140 10839 41180
rect 10797 41131 10839 41140
rect 10904 41180 10946 41189
rect 10904 41140 10905 41180
rect 10945 41140 10946 41180
rect 10904 41131 10946 41140
rect 11403 41180 11445 41189
rect 11403 41140 11404 41180
rect 11444 41140 11445 41180
rect 11403 41131 11445 41140
rect 11875 41180 11933 41181
rect 11875 41140 11884 41180
rect 11924 41140 11933 41180
rect 11875 41139 11933 41140
rect 12363 41180 12421 41181
rect 12363 41140 12372 41180
rect 12412 41140 12421 41180
rect 12363 41139 12421 41140
rect 13707 41180 13749 41189
rect 13707 41140 13708 41180
rect 13748 41140 13749 41180
rect 13707 41131 13749 41140
rect 14947 41180 15005 41181
rect 14947 41140 14956 41180
rect 14996 41140 15005 41180
rect 14947 41139 15005 41140
rect 15435 41180 15477 41189
rect 15435 41140 15436 41180
rect 15476 41140 15477 41180
rect 15435 41131 15477 41140
rect 15907 41180 15965 41181
rect 15907 41140 15916 41180
rect 15956 41140 15965 41180
rect 15907 41139 15965 41140
rect 16107 41180 16149 41189
rect 16107 41140 16108 41180
rect 16148 41140 16149 41180
rect 16107 41131 16149 41140
rect 16395 41180 16437 41189
rect 16395 41140 16396 41180
rect 16436 41140 16437 41180
rect 16395 41131 16437 41140
rect 17635 41180 17693 41181
rect 17635 41140 17644 41180
rect 17684 41140 17693 41180
rect 17635 41139 17693 41140
rect 18106 41180 18164 41181
rect 18106 41140 18115 41180
rect 18155 41140 18164 41180
rect 18106 41139 18164 41140
rect 18219 41180 18261 41189
rect 18219 41140 18220 41180
rect 18260 41140 18261 41180
rect 18219 41131 18261 41140
rect 18699 41180 18741 41189
rect 18699 41140 18700 41180
rect 18740 41140 18741 41180
rect 18699 41131 18741 41140
rect 19171 41180 19229 41181
rect 19171 41140 19180 41180
rect 19220 41140 19229 41180
rect 19171 41139 19229 41140
rect 19659 41180 19717 41181
rect 19659 41140 19668 41180
rect 19708 41140 19717 41180
rect 19659 41139 19717 41140
rect 6699 41096 6741 41105
rect 6699 41056 6700 41096
rect 6740 41056 6741 41096
rect 6699 41047 6741 41056
rect 15613 41096 15655 41105
rect 15613 41056 15614 41096
rect 15654 41056 15655 41096
rect 15613 41047 15655 41056
rect 4299 41012 4341 41021
rect 4299 40972 4300 41012
rect 4340 40972 4341 41012
rect 4299 40963 4341 40972
rect 5338 41012 5396 41013
rect 5338 40972 5347 41012
rect 5387 40972 5396 41012
rect 5338 40971 5396 40972
rect 5866 41012 5924 41013
rect 5866 40972 5875 41012
rect 5915 40972 5924 41012
rect 5866 40971 5924 40972
rect 6219 41012 6261 41021
rect 6219 40972 6220 41012
rect 6260 40972 6261 41012
rect 6219 40963 6261 40972
rect 6586 41012 6644 41013
rect 6586 40972 6595 41012
rect 6635 40972 6644 41012
rect 6586 40971 6644 40972
rect 6939 41012 6981 41021
rect 6939 40972 6940 41012
rect 6980 40972 6981 41012
rect 6939 40963 6981 40972
rect 12555 41012 12597 41021
rect 12555 40972 12556 41012
rect 12596 40972 12597 41012
rect 12555 40963 12597 40972
rect 15819 41012 15861 41021
rect 15819 40972 15820 41012
rect 15860 40972 15861 41012
rect 15819 40963 15861 40972
rect 17835 41012 17877 41021
rect 17835 40972 17836 41012
rect 17876 40972 17877 41012
rect 17835 40963 17877 40972
rect 19851 41012 19893 41021
rect 19851 40972 19852 41012
rect 19892 40972 19893 41012
rect 19851 40963 19893 40972
rect 1152 40844 20452 40868
rect 1152 40804 4928 40844
rect 4968 40804 5010 40844
rect 5050 40804 5092 40844
rect 5132 40804 5174 40844
rect 5214 40804 5256 40844
rect 5296 40804 20048 40844
rect 20088 40804 20130 40844
rect 20170 40804 20212 40844
rect 20252 40804 20294 40844
rect 20334 40804 20376 40844
rect 20416 40804 20452 40844
rect 1152 40780 20452 40804
rect 1851 40676 1893 40685
rect 1851 40636 1852 40676
rect 1892 40636 1893 40676
rect 1851 40627 1893 40636
rect 2235 40676 2277 40685
rect 2235 40636 2236 40676
rect 2276 40636 2277 40676
rect 2235 40627 2277 40636
rect 4395 40676 4437 40685
rect 4395 40636 4396 40676
rect 4436 40636 4437 40676
rect 4395 40627 4437 40636
rect 6795 40676 6837 40685
rect 6795 40636 6796 40676
rect 6836 40636 6837 40676
rect 6795 40627 6837 40636
rect 9627 40676 9669 40685
rect 9627 40636 9628 40676
rect 9668 40636 9669 40676
rect 9627 40627 9669 40636
rect 11211 40676 11253 40685
rect 11211 40636 11212 40676
rect 11252 40636 11253 40676
rect 11211 40627 11253 40636
rect 13498 40676 13556 40677
rect 13498 40636 13507 40676
rect 13547 40636 13556 40676
rect 13498 40635 13556 40636
rect 13611 40676 13653 40685
rect 13611 40636 13612 40676
rect 13652 40636 13653 40676
rect 13611 40627 13653 40636
rect 14091 40676 14133 40685
rect 14091 40636 14092 40676
rect 14132 40636 14133 40676
rect 14091 40627 14133 40636
rect 17643 40676 17685 40685
rect 17643 40636 17644 40676
rect 17684 40636 17685 40676
rect 17643 40627 17685 40636
rect 18363 40676 18405 40685
rect 18363 40636 18364 40676
rect 18404 40636 18405 40676
rect 18363 40627 18405 40636
rect 20331 40676 20373 40685
rect 20331 40636 20332 40676
rect 20372 40636 20373 40676
rect 20331 40627 20373 40636
rect 1467 40592 1509 40601
rect 1467 40552 1468 40592
rect 1508 40552 1509 40592
rect 1467 40543 1509 40552
rect 7738 40592 7796 40593
rect 7738 40552 7747 40592
rect 7787 40552 7796 40592
rect 7738 40551 7796 40552
rect 8475 40592 8517 40601
rect 8475 40552 8476 40592
rect 8516 40552 8517 40592
rect 8475 40543 8517 40552
rect 12925 40592 12967 40601
rect 12925 40552 12926 40592
rect 12966 40552 12967 40592
rect 12925 40543 12967 40552
rect 13018 40592 13076 40593
rect 13018 40552 13027 40592
rect 13067 40552 13076 40592
rect 13018 40551 13076 40552
rect 13131 40592 13173 40601
rect 13131 40552 13132 40592
rect 13172 40552 13173 40592
rect 13131 40543 13173 40552
rect 13978 40592 14036 40593
rect 13978 40552 13987 40592
rect 14027 40552 14036 40592
rect 13978 40551 14036 40552
rect 15675 40592 15717 40601
rect 15675 40552 15676 40592
rect 15716 40552 15717 40592
rect 15675 40543 15717 40552
rect 2650 40508 2708 40509
rect 2650 40468 2659 40508
rect 2699 40468 2708 40508
rect 2650 40467 2708 40468
rect 2768 40508 2810 40517
rect 2768 40468 2769 40508
rect 2809 40468 2810 40508
rect 2768 40459 2810 40468
rect 3147 40508 3189 40517
rect 4207 40508 4265 40509
rect 3147 40468 3148 40508
rect 3188 40468 3189 40508
rect 3147 40459 3189 40468
rect 3723 40499 3765 40508
rect 3723 40459 3724 40499
rect 3764 40459 3765 40499
rect 4207 40468 4216 40508
rect 4256 40468 4265 40508
rect 4207 40467 4265 40468
rect 5050 40508 5108 40509
rect 5050 40468 5059 40508
rect 5099 40468 5108 40508
rect 5050 40467 5108 40468
rect 5163 40508 5205 40517
rect 5163 40468 5164 40508
rect 5204 40468 5205 40508
rect 5163 40459 5205 40468
rect 5547 40508 5589 40517
rect 6973 40508 7015 40517
rect 5547 40468 5548 40508
rect 5588 40468 5589 40508
rect 5547 40459 5589 40468
rect 6123 40499 6165 40508
rect 6123 40459 6124 40499
rect 6164 40459 6165 40499
rect 3723 40450 3765 40459
rect 6123 40450 6165 40459
rect 6603 40499 6645 40508
rect 6603 40459 6604 40499
rect 6644 40459 6645 40499
rect 6973 40468 6974 40508
rect 7014 40468 7015 40508
rect 6973 40459 7015 40468
rect 7083 40508 7125 40517
rect 7083 40468 7084 40508
rect 7124 40468 7125 40508
rect 7083 40459 7125 40468
rect 7275 40508 7317 40517
rect 7275 40468 7276 40508
rect 7316 40468 7317 40508
rect 7275 40459 7317 40468
rect 7414 40508 7456 40517
rect 7414 40468 7415 40508
rect 7455 40468 7456 40508
rect 7414 40459 7456 40468
rect 7657 40508 7699 40517
rect 7657 40468 7658 40508
rect 7698 40468 7699 40508
rect 7657 40459 7699 40468
rect 9771 40508 9813 40517
rect 13405 40508 13447 40517
rect 13885 40508 13927 40517
rect 16203 40508 16245 40517
rect 18586 40508 18644 40509
rect 9771 40468 9772 40508
rect 9812 40468 9813 40508
rect 9771 40459 9813 40468
rect 11019 40499 11061 40508
rect 11019 40459 11020 40499
rect 11060 40459 11061 40499
rect 6603 40450 6645 40459
rect 11019 40450 11061 40459
rect 13227 40499 13269 40508
rect 13227 40459 13228 40499
rect 13268 40459 13269 40499
rect 13405 40468 13406 40508
rect 13446 40468 13447 40508
rect 13405 40459 13447 40468
rect 13707 40499 13749 40508
rect 13707 40459 13708 40499
rect 13748 40459 13749 40499
rect 13885 40468 13886 40508
rect 13926 40468 13927 40508
rect 13885 40459 13927 40468
rect 14187 40499 14229 40508
rect 14187 40459 14188 40499
rect 14228 40459 14229 40499
rect 16203 40468 16204 40508
rect 16244 40468 16245 40508
rect 16203 40459 16245 40468
rect 17451 40499 17493 40508
rect 17451 40459 17452 40499
rect 17492 40459 17493 40499
rect 18586 40468 18595 40508
rect 18635 40468 18644 40508
rect 18586 40467 18644 40468
rect 18699 40508 18741 40517
rect 18699 40468 18700 40508
rect 18740 40468 18741 40508
rect 18699 40459 18741 40468
rect 19083 40508 19125 40517
rect 19083 40468 19084 40508
rect 19124 40468 19125 40508
rect 19083 40459 19125 40468
rect 19659 40499 19701 40508
rect 19659 40459 19660 40499
rect 19700 40459 19701 40499
rect 13227 40450 13269 40459
rect 13707 40450 13749 40459
rect 14187 40450 14229 40459
rect 17451 40450 17493 40459
rect 19659 40450 19701 40459
rect 20139 40499 20181 40508
rect 20139 40459 20140 40499
rect 20180 40459 20181 40499
rect 20139 40450 20181 40459
rect 1227 40424 1269 40433
rect 1227 40384 1228 40424
rect 1268 40384 1269 40424
rect 1227 40375 1269 40384
rect 1611 40424 1653 40433
rect 1611 40384 1612 40424
rect 1652 40384 1653 40424
rect 1611 40375 1653 40384
rect 1995 40424 2037 40433
rect 1995 40384 1996 40424
rect 2036 40384 2037 40424
rect 1995 40375 2037 40384
rect 3243 40424 3285 40433
rect 3243 40384 3244 40424
rect 3284 40384 3285 40424
rect 3243 40375 3285 40384
rect 5643 40424 5685 40433
rect 5643 40384 5644 40424
rect 5684 40384 5685 40424
rect 5643 40375 5685 40384
rect 7546 40424 7604 40425
rect 7546 40384 7555 40424
rect 7595 40384 7604 40424
rect 7546 40383 7604 40384
rect 8235 40424 8277 40433
rect 8235 40384 8236 40424
rect 8276 40384 8277 40424
rect 8235 40375 8277 40384
rect 8619 40424 8661 40433
rect 8619 40384 8620 40424
rect 8660 40384 8661 40424
rect 8619 40375 8661 40384
rect 9195 40424 9237 40433
rect 9195 40384 9196 40424
rect 9236 40384 9237 40424
rect 9195 40375 9237 40384
rect 9387 40424 9429 40433
rect 9387 40384 9388 40424
rect 9428 40384 9429 40424
rect 9387 40375 9429 40384
rect 12555 40424 12597 40433
rect 12555 40384 12556 40424
rect 12596 40384 12597 40424
rect 12555 40375 12597 40384
rect 14667 40424 14709 40433
rect 14667 40384 14668 40424
rect 14708 40384 14709 40424
rect 14667 40375 14709 40384
rect 15051 40424 15093 40433
rect 15051 40384 15052 40424
rect 15092 40384 15093 40424
rect 15051 40375 15093 40384
rect 15435 40424 15477 40433
rect 15435 40384 15436 40424
rect 15476 40384 15477 40424
rect 15435 40375 15477 40384
rect 15819 40424 15861 40433
rect 15819 40384 15820 40424
rect 15860 40384 15861 40424
rect 15819 40375 15861 40384
rect 16059 40424 16101 40433
rect 16059 40384 16060 40424
rect 16100 40384 16101 40424
rect 16059 40375 16101 40384
rect 18123 40424 18165 40433
rect 18123 40384 18124 40424
rect 18164 40384 18165 40424
rect 18123 40375 18165 40384
rect 19179 40424 19221 40433
rect 19179 40384 19180 40424
rect 19220 40384 19221 40424
rect 19179 40375 19221 40384
rect 8859 40340 8901 40349
rect 8859 40300 8860 40340
rect 8900 40300 8901 40340
rect 8859 40291 8901 40300
rect 12795 40340 12837 40349
rect 12795 40300 12796 40340
rect 12836 40300 12837 40340
rect 12795 40291 12837 40300
rect 15291 40340 15333 40349
rect 15291 40300 15292 40340
rect 15332 40300 15333 40340
rect 15291 40291 15333 40300
rect 6987 40256 7029 40265
rect 6987 40216 6988 40256
rect 7028 40216 7029 40256
rect 6987 40207 7029 40216
rect 8955 40256 8997 40265
rect 8955 40216 8956 40256
rect 8996 40216 8997 40256
rect 8955 40207 8997 40216
rect 14907 40256 14949 40265
rect 14907 40216 14908 40256
rect 14948 40216 14949 40256
rect 14907 40207 14949 40216
rect 1152 40088 20448 40112
rect 1152 40048 3688 40088
rect 3728 40048 3770 40088
rect 3810 40048 3852 40088
rect 3892 40048 3934 40088
rect 3974 40048 4016 40088
rect 4056 40048 18808 40088
rect 18848 40048 18890 40088
rect 18930 40048 18972 40088
rect 19012 40048 19054 40088
rect 19094 40048 19136 40088
rect 19176 40048 20448 40088
rect 1152 40024 20448 40048
rect 1467 39920 1509 39929
rect 1467 39880 1468 39920
rect 1508 39880 1509 39920
rect 1467 39871 1509 39880
rect 1851 39920 1893 39929
rect 1851 39880 1852 39920
rect 1892 39880 1893 39920
rect 1851 39871 1893 39880
rect 6394 39920 6452 39921
rect 6394 39880 6403 39920
rect 6443 39880 6452 39920
rect 6394 39879 6452 39880
rect 6874 39920 6932 39921
rect 6874 39880 6883 39920
rect 6923 39880 6932 39920
rect 6874 39879 6932 39880
rect 17739 39920 17781 39929
rect 17739 39880 17740 39920
rect 17780 39880 17781 39920
rect 17739 39871 17781 39880
rect 18747 39920 18789 39929
rect 18747 39880 18748 39920
rect 18788 39880 18789 39920
rect 18747 39871 18789 39880
rect 20331 39920 20373 39929
rect 20331 39880 20332 39920
rect 20372 39880 20373 39920
rect 20331 39871 20373 39880
rect 4731 39836 4773 39845
rect 4731 39796 4732 39836
rect 4772 39796 4773 39836
rect 4731 39787 4773 39796
rect 6027 39836 6069 39845
rect 6027 39796 6028 39836
rect 6068 39796 6069 39836
rect 6027 39787 6069 39796
rect 11067 39836 11109 39845
rect 11067 39796 11068 39836
rect 11108 39796 11109 39836
rect 11067 39787 11109 39796
rect 12027 39836 12069 39845
rect 12027 39796 12028 39836
rect 12068 39796 12069 39836
rect 12027 39787 12069 39796
rect 18363 39836 18405 39845
rect 18363 39796 18364 39836
rect 18404 39796 18405 39836
rect 18363 39787 18405 39796
rect 1227 39752 1269 39761
rect 1227 39712 1228 39752
rect 1268 39712 1269 39752
rect 1227 39703 1269 39712
rect 1611 39752 1653 39761
rect 1611 39712 1612 39752
rect 1652 39712 1653 39752
rect 1611 39703 1653 39712
rect 1995 39752 2037 39761
rect 1995 39712 1996 39752
rect 2036 39712 2037 39752
rect 1995 39703 2037 39712
rect 3147 39752 3189 39761
rect 3147 39712 3148 39752
rect 3188 39712 3189 39752
rect 3147 39703 3189 39712
rect 6118 39752 6176 39753
rect 6118 39712 6127 39752
rect 6167 39712 6176 39752
rect 6118 39711 6176 39712
rect 10827 39752 10869 39761
rect 10827 39712 10828 39752
rect 10868 39712 10869 39752
rect 10827 39703 10869 39712
rect 12386 39752 12428 39761
rect 12386 39712 12387 39752
rect 12427 39712 12428 39752
rect 12386 39703 12428 39712
rect 13690 39752 13748 39753
rect 13690 39712 13699 39752
rect 13739 39712 13748 39752
rect 13690 39711 13748 39712
rect 14667 39752 14709 39761
rect 14667 39712 14668 39752
rect 14708 39712 14709 39752
rect 14667 39703 14709 39712
rect 18123 39752 18165 39761
rect 18123 39712 18124 39752
rect 18164 39712 18165 39752
rect 18123 39703 18165 39712
rect 18507 39752 18549 39761
rect 18507 39712 18508 39752
rect 18548 39712 18549 39752
rect 18507 39703 18549 39712
rect 2650 39668 2708 39669
rect 2650 39628 2659 39668
rect 2699 39628 2708 39668
rect 2650 39627 2708 39628
rect 2763 39668 2805 39677
rect 2763 39628 2764 39668
rect 2804 39628 2805 39668
rect 2763 39619 2805 39628
rect 3243 39668 3285 39677
rect 3243 39628 3244 39668
rect 3284 39628 3285 39668
rect 3243 39619 3285 39628
rect 3715 39668 3773 39669
rect 3715 39628 3724 39668
rect 3764 39628 3773 39668
rect 3715 39627 3773 39628
rect 4203 39668 4261 39669
rect 4203 39628 4212 39668
rect 4252 39628 4261 39668
rect 4203 39627 4261 39628
rect 4587 39668 4629 39677
rect 4587 39628 4588 39668
rect 4628 39628 4629 39668
rect 4587 39619 4629 39628
rect 4731 39668 4773 39677
rect 4731 39628 4732 39668
rect 4772 39628 4773 39668
rect 4731 39619 4773 39628
rect 4875 39668 4917 39677
rect 4875 39628 4876 39668
rect 4916 39628 4917 39668
rect 4875 39619 4917 39628
rect 5050 39668 5108 39669
rect 5050 39628 5059 39668
rect 5099 39628 5108 39668
rect 5050 39627 5108 39628
rect 5163 39668 5205 39677
rect 5163 39628 5164 39668
rect 5204 39628 5205 39668
rect 5163 39619 5205 39628
rect 5302 39668 5344 39677
rect 5302 39628 5303 39668
rect 5343 39628 5344 39668
rect 5302 39619 5344 39628
rect 5434 39668 5492 39669
rect 5434 39628 5443 39668
rect 5483 39628 5492 39668
rect 5434 39627 5492 39628
rect 5547 39668 5589 39677
rect 5547 39628 5548 39668
rect 5588 39628 5589 39668
rect 5547 39619 5589 39628
rect 5787 39668 5829 39677
rect 5787 39628 5788 39668
rect 5828 39628 5829 39668
rect 5787 39619 5829 39628
rect 5952 39668 5994 39677
rect 5952 39628 5953 39668
rect 5993 39628 5994 39668
rect 5952 39619 5994 39628
rect 6250 39668 6308 39669
rect 6250 39628 6259 39668
rect 6299 39628 6308 39668
rect 6250 39627 6308 39628
rect 6691 39668 6749 39669
rect 6691 39628 6700 39668
rect 6740 39628 6749 39668
rect 6691 39627 6749 39628
rect 7171 39668 7229 39669
rect 7171 39628 7180 39668
rect 7220 39628 7229 39668
rect 7171 39627 7229 39628
rect 7563 39668 7605 39677
rect 7563 39628 7564 39668
rect 7604 39628 7605 39668
rect 7563 39619 7605 39628
rect 8811 39668 8869 39669
rect 8811 39628 8820 39668
rect 8860 39628 8869 39668
rect 8811 39627 8869 39628
rect 9195 39668 9237 39677
rect 9195 39628 9196 39668
rect 9236 39628 9237 39668
rect 9195 39619 9237 39628
rect 10443 39668 10501 39669
rect 10443 39628 10452 39668
rect 10492 39628 10501 39668
rect 10443 39627 10501 39628
rect 11883 39668 11925 39677
rect 11883 39628 11884 39668
rect 11924 39628 11925 39668
rect 11883 39619 11925 39628
rect 12267 39668 12309 39677
rect 12267 39628 12268 39668
rect 12308 39628 12309 39668
rect 12267 39619 12309 39628
rect 12496 39668 12554 39669
rect 12496 39628 12505 39668
rect 12545 39628 12554 39668
rect 12496 39627 12554 39628
rect 12747 39668 12789 39677
rect 12747 39628 12748 39668
rect 12788 39628 12789 39668
rect 12747 39619 12789 39628
rect 13018 39668 13076 39669
rect 13018 39628 13027 39668
rect 13067 39628 13076 39668
rect 13018 39627 13076 39628
rect 13558 39668 13600 39677
rect 13558 39628 13559 39668
rect 13599 39628 13600 39668
rect 13558 39619 13600 39628
rect 13803 39668 13845 39677
rect 13803 39628 13804 39668
rect 13844 39628 13845 39668
rect 13803 39619 13845 39628
rect 14170 39668 14228 39669
rect 14170 39628 14179 39668
rect 14219 39628 14228 39668
rect 14170 39627 14228 39628
rect 14283 39668 14325 39677
rect 14283 39628 14284 39668
rect 14324 39628 14325 39668
rect 14283 39619 14325 39628
rect 14763 39668 14805 39677
rect 14763 39628 14764 39668
rect 14804 39628 14805 39668
rect 14763 39619 14805 39628
rect 15235 39668 15293 39669
rect 15235 39628 15244 39668
rect 15284 39628 15293 39668
rect 15235 39627 15293 39628
rect 15754 39668 15812 39669
rect 15754 39628 15763 39668
rect 15803 39628 15812 39668
rect 15754 39627 15812 39628
rect 16299 39668 16341 39677
rect 16299 39628 16300 39668
rect 16340 39628 16341 39668
rect 16299 39619 16341 39628
rect 17539 39668 17597 39669
rect 17539 39628 17548 39668
rect 17588 39628 17597 39668
rect 17539 39627 17597 39628
rect 18891 39668 18933 39677
rect 18891 39628 18892 39668
rect 18932 39628 18933 39668
rect 18891 39619 18933 39628
rect 20131 39668 20189 39669
rect 20131 39628 20140 39668
rect 20180 39628 20189 39668
rect 20131 39627 20189 39628
rect 2235 39584 2277 39593
rect 2235 39544 2236 39584
rect 2276 39544 2277 39584
rect 2235 39535 2277 39544
rect 4954 39584 5012 39585
rect 4954 39544 4963 39584
rect 5003 39544 5012 39584
rect 4954 39543 5012 39544
rect 6400 39584 6442 39593
rect 6400 39544 6401 39584
rect 6441 39544 6442 39584
rect 6400 39535 6442 39544
rect 6603 39584 6645 39593
rect 6603 39544 6604 39584
rect 6644 39544 6645 39584
rect 6603 39535 6645 39544
rect 6877 39584 6919 39593
rect 6877 39544 6878 39584
rect 6918 39544 6919 39584
rect 6877 39535 6919 39544
rect 12171 39584 12213 39593
rect 12171 39544 12172 39584
rect 12212 39544 12213 39584
rect 12171 39535 12213 39544
rect 13131 39584 13173 39593
rect 13131 39544 13132 39584
rect 13172 39544 13173 39584
rect 13131 39535 13173 39544
rect 13467 39584 13509 39593
rect 13467 39544 13468 39584
rect 13508 39544 13509 39584
rect 13467 39535 13509 39544
rect 4395 39500 4437 39509
rect 4395 39460 4396 39500
rect 4436 39460 4437 39500
rect 4395 39451 4437 39460
rect 5626 39500 5684 39501
rect 5626 39460 5635 39500
rect 5675 39460 5684 39500
rect 5626 39459 5684 39460
rect 7083 39500 7125 39509
rect 7083 39460 7084 39500
rect 7124 39460 7125 39500
rect 7083 39451 7125 39460
rect 9003 39500 9045 39509
rect 9003 39460 9004 39500
rect 9044 39460 9045 39500
rect 9003 39451 9045 39460
rect 10635 39500 10677 39509
rect 10635 39460 10636 39500
rect 10676 39460 10677 39500
rect 10635 39451 10677 39460
rect 13882 39500 13940 39501
rect 13882 39460 13891 39500
rect 13931 39460 13940 39500
rect 13882 39459 13940 39460
rect 15915 39500 15957 39509
rect 15915 39460 15916 39500
rect 15956 39460 15957 39500
rect 15915 39451 15957 39460
rect 1152 39332 20452 39356
rect 1152 39292 4928 39332
rect 4968 39292 5010 39332
rect 5050 39292 5092 39332
rect 5132 39292 5174 39332
rect 5214 39292 5256 39332
rect 5296 39292 20048 39332
rect 20088 39292 20130 39332
rect 20170 39292 20212 39332
rect 20252 39292 20294 39332
rect 20334 39292 20376 39332
rect 20416 39292 20452 39332
rect 1152 39268 20452 39292
rect 1467 39164 1509 39173
rect 1467 39124 1468 39164
rect 1508 39124 1509 39164
rect 1467 39115 1509 39124
rect 3915 39164 3957 39173
rect 3915 39124 3916 39164
rect 3956 39124 3957 39164
rect 3915 39115 3957 39124
rect 5931 39164 5973 39173
rect 5931 39124 5932 39164
rect 5972 39124 5973 39164
rect 5931 39115 5973 39124
rect 6603 39164 6645 39173
rect 6603 39124 6604 39164
rect 6644 39124 6645 39164
rect 6603 39115 6645 39124
rect 8811 39164 8853 39173
rect 8811 39124 8812 39164
rect 8852 39124 8853 39164
rect 8811 39115 8853 39124
rect 12555 39164 12597 39173
rect 12555 39124 12556 39164
rect 12596 39124 12597 39164
rect 12555 39115 12597 39124
rect 13947 39164 13989 39173
rect 13947 39124 13948 39164
rect 13988 39124 13989 39164
rect 13947 39115 13989 39124
rect 15915 39164 15957 39173
rect 15915 39124 15916 39164
rect 15956 39124 15957 39164
rect 15915 39115 15957 39124
rect 16731 39164 16773 39173
rect 16731 39124 16732 39164
rect 16772 39124 16773 39164
rect 16731 39115 16773 39124
rect 13611 39080 13653 39089
rect 13611 39040 13612 39080
rect 13652 39040 13653 39080
rect 7162 39029 7220 39034
rect 13611 39031 13653 39040
rect 14331 39080 14373 39089
rect 14331 39040 14332 39080
rect 14372 39040 14373 39080
rect 14331 39031 14373 39040
rect 2475 38996 2517 39005
rect 4186 38996 4244 38997
rect 2475 38956 2476 38996
rect 2516 38956 2517 38996
rect 2475 38947 2517 38956
rect 3723 38987 3765 38996
rect 3723 38947 3724 38987
rect 3764 38947 3765 38987
rect 4186 38956 4195 38996
rect 4235 38956 4244 38996
rect 4186 38955 4244 38956
rect 4299 38996 4341 39005
rect 4299 38956 4300 38996
rect 4340 38956 4341 38996
rect 4299 38947 4341 38956
rect 4683 38996 4725 39005
rect 6123 38996 6165 39005
rect 4683 38956 4684 38996
rect 4724 38956 4725 38996
rect 4683 38947 4725 38956
rect 5259 38987 5301 38996
rect 5259 38947 5260 38987
rect 5300 38947 5301 38987
rect 3723 38938 3765 38947
rect 5259 38938 5301 38947
rect 5739 38987 5781 38996
rect 5739 38947 5740 38987
rect 5780 38947 5781 38987
rect 6123 38956 6124 38996
rect 6164 38956 6165 38996
rect 6123 38947 6165 38956
rect 6238 38996 6280 39005
rect 6238 38956 6239 38996
rect 6279 38956 6280 38996
rect 6238 38947 6280 38956
rect 6411 38996 6453 39005
rect 6411 38956 6412 38996
rect 6452 38956 6453 38996
rect 6411 38947 6453 38956
rect 6603 38996 6645 39005
rect 6603 38956 6604 38996
rect 6644 38956 6645 38996
rect 6603 38947 6645 38956
rect 6795 38996 6837 39005
rect 6795 38956 6796 38996
rect 6836 38956 6837 38996
rect 6795 38947 6837 38956
rect 7053 38996 7095 39005
rect 7053 38956 7054 38996
rect 7094 38956 7095 38996
rect 7162 38989 7171 39029
rect 7211 38989 7220 39029
rect 7162 38988 7220 38989
rect 7563 38996 7605 39005
rect 9003 38996 9045 39005
rect 11115 38996 11157 39005
rect 12747 38996 12789 39005
rect 7053 38947 7095 38956
rect 7563 38956 7564 38996
rect 7604 38956 7605 38996
rect 7563 38947 7605 38956
rect 8139 38987 8181 38996
rect 8139 38947 8140 38987
rect 8180 38947 8181 38987
rect 5739 38938 5781 38947
rect 8139 38938 8181 38947
rect 8619 38987 8661 38996
rect 8619 38947 8620 38987
rect 8660 38947 8661 38987
rect 9003 38956 9004 38996
rect 9044 38956 9045 38996
rect 9003 38947 9045 38956
rect 10251 38987 10293 38996
rect 10251 38947 10252 38987
rect 10292 38947 10293 38987
rect 11115 38956 11116 38996
rect 11156 38956 11157 38996
rect 11115 38947 11157 38956
rect 12363 38987 12405 38996
rect 12363 38947 12364 38987
rect 12404 38947 12405 38987
rect 12747 38956 12748 38996
rect 12788 38956 12789 38996
rect 12747 38947 12789 38956
rect 12939 38996 12981 39005
rect 12939 38956 12940 38996
rect 12980 38956 12981 38996
rect 12939 38947 12981 38956
rect 13227 38996 13269 39005
rect 13227 38956 13228 38996
rect 13268 38956 13269 38996
rect 13227 38947 13269 38956
rect 13498 38996 13556 38997
rect 13498 38956 13507 38996
rect 13547 38956 13556 38996
rect 13498 38955 13556 38956
rect 14475 38996 14517 39005
rect 16971 38996 17013 39005
rect 18699 38996 18741 39005
rect 14475 38956 14476 38996
rect 14516 38956 14517 38996
rect 14475 38947 14517 38956
rect 15723 38987 15765 38996
rect 15723 38947 15724 38987
rect 15764 38947 15765 38987
rect 16971 38956 16972 38996
rect 17012 38956 17013 38996
rect 16971 38947 17013 38956
rect 18219 38987 18261 38996
rect 18219 38947 18220 38987
rect 18260 38947 18261 38987
rect 18699 38956 18700 38996
rect 18740 38956 18741 38996
rect 18699 38947 18741 38956
rect 19947 38987 19989 38996
rect 19947 38947 19948 38987
rect 19988 38947 19989 38987
rect 8619 38938 8661 38947
rect 10251 38938 10293 38947
rect 12363 38938 12405 38947
rect 15723 38938 15765 38947
rect 18219 38938 18261 38947
rect 19947 38938 19989 38947
rect 1227 38912 1269 38921
rect 1227 38872 1228 38912
rect 1268 38872 1269 38912
rect 1227 38863 1269 38872
rect 1611 38912 1653 38921
rect 1611 38872 1612 38912
rect 1652 38872 1653 38912
rect 1611 38863 1653 38872
rect 1995 38912 2037 38921
rect 1995 38872 1996 38912
rect 2036 38872 2037 38912
rect 1995 38863 2037 38872
rect 2235 38912 2277 38921
rect 2235 38872 2236 38912
rect 2276 38872 2277 38912
rect 2235 38863 2277 38872
rect 4779 38912 4821 38921
rect 4779 38872 4780 38912
rect 4820 38872 4821 38912
rect 4779 38863 4821 38872
rect 7659 38912 7701 38921
rect 7659 38872 7660 38912
rect 7700 38872 7701 38912
rect 7659 38863 7701 38872
rect 14091 38912 14133 38921
rect 14091 38872 14092 38912
rect 14132 38872 14133 38912
rect 14091 38863 14133 38872
rect 16299 38912 16341 38921
rect 16299 38872 16300 38912
rect 16340 38872 16341 38912
rect 16299 38863 16341 38872
rect 16491 38912 16533 38921
rect 16491 38872 16492 38912
rect 16532 38872 16533 38912
rect 16491 38863 16533 38872
rect 1851 38744 1893 38753
rect 1851 38704 1852 38744
rect 1892 38704 1893 38744
rect 1851 38695 1893 38704
rect 6123 38744 6165 38753
rect 6123 38704 6124 38744
rect 6164 38704 6165 38744
rect 6123 38695 6165 38704
rect 10443 38744 10485 38753
rect 10443 38704 10444 38744
rect 10484 38704 10485 38744
rect 10443 38695 10485 38704
rect 12747 38744 12789 38753
rect 12747 38704 12748 38744
rect 12788 38704 12789 38744
rect 12747 38695 12789 38704
rect 16059 38744 16101 38753
rect 16059 38704 16060 38744
rect 16100 38704 16101 38744
rect 16059 38695 16101 38704
rect 18411 38744 18453 38753
rect 18411 38704 18412 38744
rect 18452 38704 18453 38744
rect 18411 38695 18453 38704
rect 20139 38744 20181 38753
rect 20139 38704 20140 38744
rect 20180 38704 20181 38744
rect 20139 38695 20181 38704
rect 1152 38576 20448 38600
rect 1152 38536 3688 38576
rect 3728 38536 3770 38576
rect 3810 38536 3852 38576
rect 3892 38536 3934 38576
rect 3974 38536 4016 38576
rect 4056 38536 18808 38576
rect 18848 38536 18890 38576
rect 18930 38536 18972 38576
rect 19012 38536 19054 38576
rect 19094 38536 19136 38576
rect 19176 38536 20448 38576
rect 1152 38512 20448 38536
rect 2667 38408 2709 38417
rect 2667 38368 2668 38408
rect 2708 38368 2709 38408
rect 2667 38359 2709 38368
rect 4299 38408 4341 38417
rect 4299 38368 4300 38408
rect 4340 38368 4341 38408
rect 4299 38359 4341 38368
rect 12075 38408 12117 38417
rect 12075 38368 12076 38408
rect 12116 38368 12117 38408
rect 12075 38359 12117 38368
rect 12411 38408 12453 38417
rect 12411 38368 12412 38408
rect 12452 38368 12453 38408
rect 12411 38359 12453 38368
rect 14667 38408 14709 38417
rect 14667 38368 14668 38408
rect 14708 38368 14709 38408
rect 14667 38359 14709 38368
rect 15675 38408 15717 38417
rect 15675 38368 15676 38408
rect 15716 38368 15717 38408
rect 15675 38359 15717 38368
rect 6123 38324 6165 38333
rect 6123 38284 6124 38324
rect 6164 38284 6165 38324
rect 6123 38275 6165 38284
rect 6987 38324 7029 38333
rect 6987 38284 6988 38324
rect 7028 38284 7029 38324
rect 6987 38275 7029 38284
rect 4491 38240 4533 38249
rect 4491 38200 4492 38240
rect 4532 38200 4533 38240
rect 4491 38191 4533 38200
rect 5282 38240 5324 38249
rect 5282 38200 5283 38240
rect 5323 38200 5324 38240
rect 5282 38191 5324 38200
rect 6586 38240 6644 38241
rect 6586 38200 6595 38240
rect 6635 38200 6644 38240
rect 6586 38199 6644 38200
rect 8427 38240 8469 38249
rect 8427 38200 8428 38240
rect 8468 38200 8469 38240
rect 8427 38191 8469 38200
rect 8811 38240 8853 38249
rect 8811 38200 8812 38240
rect 8852 38200 8853 38240
rect 8811 38191 8853 38200
rect 9675 38240 9717 38249
rect 9675 38200 9676 38240
rect 9716 38200 9717 38240
rect 9675 38191 9717 38200
rect 12634 38240 12692 38241
rect 12634 38200 12643 38240
rect 12683 38200 12692 38240
rect 12634 38199 12692 38200
rect 15051 38240 15093 38249
rect 15051 38200 15052 38240
rect 15092 38200 15093 38240
rect 15051 38191 15093 38200
rect 15435 38240 15477 38249
rect 15435 38200 15436 38240
rect 15476 38200 15477 38240
rect 15435 38191 15477 38200
rect 15819 38240 15861 38249
rect 15819 38200 15820 38240
rect 15860 38200 15861 38240
rect 15819 38191 15861 38200
rect 16491 38240 16533 38249
rect 16491 38200 16492 38240
rect 16532 38200 16533 38240
rect 16491 38191 16533 38200
rect 18987 38240 19029 38249
rect 18987 38200 18988 38240
rect 19028 38200 19029 38240
rect 18987 38191 19029 38200
rect 18498 38174 18544 38183
rect 1227 38156 1269 38165
rect 1227 38116 1228 38156
rect 1268 38116 1269 38156
rect 1227 38107 1269 38116
rect 2467 38156 2525 38157
rect 2467 38116 2476 38156
rect 2516 38116 2525 38156
rect 2467 38115 2525 38116
rect 2859 38156 2901 38165
rect 2859 38116 2860 38156
rect 2900 38116 2901 38156
rect 2859 38107 2901 38116
rect 4099 38156 4157 38157
rect 4099 38116 4108 38156
rect 4148 38116 4157 38156
rect 4099 38115 4157 38116
rect 5163 38156 5205 38165
rect 5163 38116 5164 38156
rect 5204 38116 5205 38156
rect 5163 38107 5205 38116
rect 5392 38156 5450 38157
rect 5392 38116 5401 38156
rect 5441 38116 5450 38156
rect 5392 38115 5450 38116
rect 5547 38156 5589 38165
rect 5547 38116 5548 38156
rect 5588 38116 5589 38156
rect 5547 38107 5589 38116
rect 5722 38156 5780 38157
rect 5722 38116 5731 38156
rect 5771 38116 5780 38156
rect 5722 38115 5780 38116
rect 5835 38156 5877 38165
rect 5835 38116 5836 38156
rect 5876 38116 5877 38156
rect 5835 38107 5877 38116
rect 6027 38156 6069 38165
rect 6027 38116 6028 38156
rect 6068 38116 6069 38156
rect 6027 38107 6069 38116
rect 6144 38156 6202 38157
rect 6144 38116 6153 38156
rect 6193 38116 6202 38156
rect 6144 38115 6202 38116
rect 6315 38156 6357 38165
rect 6315 38116 6316 38156
rect 6356 38116 6357 38156
rect 6315 38107 6357 38116
rect 6466 38156 6524 38157
rect 6466 38116 6475 38156
rect 6515 38116 6524 38156
rect 6466 38115 6524 38116
rect 6699 38156 6741 38165
rect 6699 38116 6700 38156
rect 6740 38116 6741 38156
rect 6699 38107 6741 38116
rect 6987 38156 7029 38165
rect 6987 38116 6988 38156
rect 7028 38116 7029 38156
rect 6987 38107 7029 38116
rect 7102 38156 7144 38165
rect 7102 38116 7103 38156
rect 7143 38116 7144 38156
rect 7102 38107 7144 38116
rect 7275 38156 7317 38165
rect 7275 38116 7276 38156
rect 7316 38116 7317 38156
rect 7275 38107 7317 38116
rect 10635 38156 10677 38165
rect 10635 38116 10636 38156
rect 10676 38116 10677 38156
rect 10635 38107 10677 38116
rect 11875 38156 11933 38157
rect 11875 38116 11884 38156
rect 11924 38116 11933 38156
rect 11875 38115 11933 38116
rect 12267 38156 12309 38165
rect 12267 38116 12268 38156
rect 12308 38116 12309 38156
rect 12267 38107 12309 38116
rect 12502 38156 12544 38165
rect 12502 38116 12503 38156
rect 12543 38116 12544 38156
rect 12502 38107 12544 38116
rect 12747 38156 12789 38165
rect 12747 38116 12748 38156
rect 12788 38116 12789 38156
rect 12747 38107 12789 38116
rect 13227 38156 13269 38165
rect 13227 38116 13228 38156
rect 13268 38116 13269 38156
rect 13227 38107 13269 38116
rect 14467 38156 14525 38157
rect 14467 38116 14476 38156
rect 14516 38116 14525 38156
rect 14467 38115 14525 38116
rect 16779 38156 16821 38165
rect 16779 38116 16780 38156
rect 16820 38116 16821 38156
rect 16779 38107 16821 38116
rect 18019 38156 18077 38157
rect 18019 38116 18028 38156
rect 18068 38116 18077 38156
rect 18498 38134 18499 38174
rect 18539 38134 18544 38174
rect 18498 38125 18544 38134
rect 18592 38156 18650 38157
rect 18019 38115 18077 38116
rect 18592 38116 18601 38156
rect 18641 38116 18650 38156
rect 18592 38115 18650 38116
rect 19083 38156 19125 38165
rect 19083 38116 19084 38156
rect 19124 38116 19125 38156
rect 19083 38107 19125 38116
rect 19555 38156 19613 38157
rect 19555 38116 19564 38156
rect 19604 38116 19613 38156
rect 19555 38115 19613 38116
rect 20074 38156 20132 38157
rect 20074 38116 20083 38156
rect 20123 38116 20132 38156
rect 20074 38115 20132 38116
rect 5626 38072 5684 38073
rect 5626 38032 5635 38072
rect 5675 38032 5684 38072
rect 5626 38031 5684 38032
rect 16059 38072 16101 38081
rect 16059 38032 16060 38072
rect 16100 38032 16101 38072
rect 16059 38023 16101 38032
rect 4731 37988 4773 37997
rect 4731 37948 4732 37988
rect 4772 37948 4773 37988
rect 4731 37939 4773 37948
rect 5067 37988 5109 37997
rect 5067 37948 5068 37988
rect 5108 37948 5109 37988
rect 5067 37939 5109 37948
rect 6778 37988 6836 37989
rect 6778 37948 6787 37988
rect 6827 37948 6836 37988
rect 6778 37947 6836 37948
rect 8187 37988 8229 37997
rect 8187 37948 8188 37988
rect 8228 37948 8229 37988
rect 8187 37939 8229 37948
rect 8571 37988 8613 37997
rect 8571 37948 8572 37988
rect 8612 37948 8613 37988
rect 8571 37939 8613 37948
rect 9435 37988 9477 37997
rect 9435 37948 9436 37988
rect 9476 37948 9477 37988
rect 9435 37939 9477 37948
rect 12826 37988 12884 37989
rect 12826 37948 12835 37988
rect 12875 37948 12884 37988
rect 12826 37947 12884 37948
rect 14811 37988 14853 37997
rect 14811 37948 14812 37988
rect 14852 37948 14853 37988
rect 14811 37939 14853 37948
rect 16251 37988 16293 37997
rect 16251 37948 16252 37988
rect 16292 37948 16293 37988
rect 16251 37939 16293 37948
rect 18219 37988 18261 37997
rect 18219 37948 18220 37988
rect 18260 37948 18261 37988
rect 18219 37939 18261 37948
rect 20235 37988 20277 37997
rect 20235 37948 20236 37988
rect 20276 37948 20277 37988
rect 20235 37939 20277 37948
rect 1152 37820 20452 37844
rect 1152 37780 4928 37820
rect 4968 37780 5010 37820
rect 5050 37780 5092 37820
rect 5132 37780 5174 37820
rect 5214 37780 5256 37820
rect 5296 37780 20048 37820
rect 20088 37780 20130 37820
rect 20170 37780 20212 37820
rect 20252 37780 20294 37820
rect 20334 37780 20376 37820
rect 20416 37780 20452 37820
rect 1152 37756 20452 37780
rect 5451 37652 5493 37661
rect 5451 37612 5452 37652
rect 5492 37612 5493 37652
rect 5451 37603 5493 37612
rect 8026 37652 8084 37653
rect 8026 37612 8035 37652
rect 8075 37612 8084 37652
rect 8026 37611 8084 37612
rect 12171 37652 12213 37661
rect 12171 37612 12172 37652
rect 12212 37612 12213 37652
rect 12171 37603 12213 37612
rect 13371 37652 13413 37661
rect 13371 37612 13372 37652
rect 13412 37612 13413 37652
rect 13371 37603 13413 37612
rect 7083 37568 7125 37577
rect 7083 37528 7084 37568
rect 7124 37528 7125 37568
rect 7083 37519 7125 37528
rect 8246 37568 8288 37577
rect 8246 37528 8247 37568
rect 8287 37528 8288 37568
rect 8246 37519 8288 37528
rect 17883 37568 17925 37577
rect 17883 37528 17884 37568
rect 17924 37528 17925 37568
rect 17883 37519 17925 37528
rect 1227 37484 1269 37493
rect 4011 37484 4053 37493
rect 5643 37484 5685 37493
rect 7930 37484 7988 37485
rect 10539 37484 10581 37493
rect 1227 37444 1228 37484
rect 1268 37444 1269 37484
rect 1227 37435 1269 37444
rect 2475 37475 2517 37484
rect 2475 37435 2476 37475
rect 2516 37435 2517 37475
rect 4011 37444 4012 37484
rect 4052 37444 4053 37484
rect 4011 37435 4053 37444
rect 5259 37475 5301 37484
rect 5259 37435 5260 37475
rect 5300 37435 5301 37475
rect 5643 37444 5644 37484
rect 5684 37444 5685 37484
rect 5643 37435 5685 37444
rect 6891 37475 6933 37484
rect 6891 37435 6892 37475
rect 6932 37435 6933 37475
rect 2475 37426 2517 37435
rect 5259 37426 5301 37435
rect 6891 37426 6933 37435
rect 7371 37475 7413 37484
rect 7371 37435 7372 37475
rect 7412 37435 7413 37475
rect 7602 37475 7648 37484
rect 7371 37426 7413 37435
rect 7470 37464 7512 37473
rect 7470 37424 7471 37464
rect 7511 37424 7512 37464
rect 7602 37435 7603 37475
rect 7643 37435 7648 37475
rect 7930 37444 7939 37484
rect 7979 37444 7988 37484
rect 7930 37443 7988 37444
rect 9291 37475 9333 37484
rect 7602 37426 7648 37435
rect 9291 37435 9292 37475
rect 9332 37435 9333 37475
rect 10539 37444 10540 37484
rect 10580 37444 10581 37484
rect 10539 37435 10581 37444
rect 10731 37484 10773 37493
rect 12610 37484 12668 37485
rect 10731 37444 10732 37484
rect 10772 37444 10773 37484
rect 10731 37435 10773 37444
rect 11979 37475 12021 37484
rect 11979 37435 11980 37475
rect 12020 37435 12021 37475
rect 12610 37444 12619 37484
rect 12659 37444 12668 37484
rect 12610 37443 12668 37444
rect 12843 37484 12885 37493
rect 12843 37444 12844 37484
rect 12884 37444 12885 37484
rect 12843 37435 12885 37444
rect 13515 37484 13557 37493
rect 13515 37444 13516 37484
rect 13556 37444 13557 37484
rect 13515 37435 13557 37444
rect 13803 37484 13845 37493
rect 16875 37484 16917 37493
rect 13803 37444 13804 37484
rect 13844 37444 13845 37484
rect 13803 37435 13845 37444
rect 15051 37475 15093 37484
rect 15051 37435 15052 37475
rect 15092 37435 15093 37475
rect 9291 37426 9333 37435
rect 11979 37426 12021 37435
rect 15051 37426 15093 37435
rect 15627 37475 15669 37484
rect 15627 37435 15628 37475
rect 15668 37435 15669 37475
rect 16875 37444 16876 37484
rect 16916 37444 16917 37484
rect 16875 37435 16917 37444
rect 18490 37484 18548 37485
rect 18490 37444 18499 37484
rect 18539 37444 18548 37484
rect 18490 37443 18548 37444
rect 18603 37484 18645 37493
rect 18603 37444 18604 37484
rect 18644 37444 18645 37484
rect 18603 37435 18645 37444
rect 18987 37484 19029 37493
rect 18987 37444 18988 37484
rect 19028 37444 19029 37484
rect 18987 37435 19029 37444
rect 19563 37475 19605 37484
rect 19563 37435 19564 37475
rect 19604 37435 19605 37475
rect 15627 37426 15669 37435
rect 19563 37426 19605 37435
rect 20043 37475 20085 37484
rect 20043 37435 20044 37475
rect 20084 37435 20085 37475
rect 20043 37426 20085 37435
rect 7470 37415 7512 37424
rect 2859 37400 2901 37409
rect 2859 37360 2860 37400
rect 2900 37360 2901 37400
rect 2859 37351 2901 37360
rect 3099 37400 3141 37409
rect 3099 37360 3100 37400
rect 3140 37360 3141 37400
rect 3099 37351 3141 37360
rect 3243 37400 3285 37409
rect 3243 37360 3244 37400
rect 3284 37360 3285 37400
rect 3243 37351 3285 37360
rect 3627 37400 3669 37409
rect 3627 37360 3628 37400
rect 3668 37360 3669 37400
rect 3627 37351 3669 37360
rect 8715 37400 8757 37409
rect 8715 37360 8716 37400
rect 8756 37360 8757 37400
rect 8715 37351 8757 37360
rect 12730 37400 12788 37401
rect 12730 37360 12739 37400
rect 12779 37360 12788 37400
rect 12730 37359 12788 37360
rect 12939 37400 12981 37409
rect 12939 37360 12940 37400
rect 12980 37360 12981 37400
rect 12939 37351 12981 37360
rect 13131 37400 13173 37409
rect 13131 37360 13132 37400
rect 13172 37360 13173 37400
rect 13131 37351 13173 37360
rect 13659 37400 13701 37409
rect 13659 37360 13660 37400
rect 13700 37360 13701 37400
rect 13659 37351 13701 37360
rect 17067 37400 17109 37409
rect 17067 37360 17068 37400
rect 17108 37360 17109 37400
rect 17067 37351 17109 37360
rect 17307 37400 17349 37409
rect 17307 37360 17308 37400
rect 17348 37360 17349 37400
rect 17307 37351 17349 37360
rect 17643 37400 17685 37409
rect 17643 37360 17644 37400
rect 17684 37360 17685 37400
rect 17643 37351 17685 37360
rect 18123 37400 18165 37409
rect 18123 37360 18124 37400
rect 18164 37360 18165 37400
rect 18123 37351 18165 37360
rect 19083 37400 19125 37409
rect 19083 37360 19084 37400
rect 19124 37360 19125 37400
rect 19083 37351 19125 37360
rect 2667 37316 2709 37325
rect 2667 37276 2668 37316
rect 2708 37276 2709 37316
rect 2667 37267 2709 37276
rect 8955 37316 8997 37325
rect 8955 37276 8956 37316
rect 8996 37276 8997 37316
rect 8955 37267 8997 37276
rect 15243 37316 15285 37325
rect 15243 37276 15244 37316
rect 15284 37276 15285 37316
rect 15243 37267 15285 37276
rect 3483 37232 3525 37241
rect 3483 37192 3484 37232
rect 3524 37192 3525 37232
rect 3483 37183 3525 37192
rect 3867 37232 3909 37241
rect 3867 37192 3868 37232
rect 3908 37192 3909 37232
rect 3867 37183 3909 37192
rect 7083 37232 7125 37241
rect 7083 37192 7084 37232
rect 7124 37192 7125 37232
rect 7083 37183 7125 37192
rect 7755 37232 7797 37241
rect 7755 37192 7756 37232
rect 7796 37192 7797 37232
rect 7755 37183 7797 37192
rect 8235 37232 8277 37241
rect 8235 37192 8236 37232
rect 8276 37192 8277 37232
rect 8235 37183 8277 37192
rect 9099 37232 9141 37241
rect 9099 37192 9100 37232
rect 9140 37192 9141 37232
rect 9099 37183 9141 37192
rect 15435 37232 15477 37241
rect 15435 37192 15436 37232
rect 15476 37192 15477 37232
rect 15435 37183 15477 37192
rect 17403 37232 17445 37241
rect 17403 37192 17404 37232
rect 17444 37192 17445 37232
rect 17403 37183 17445 37192
rect 20266 37232 20324 37233
rect 20266 37192 20275 37232
rect 20315 37192 20324 37232
rect 20266 37191 20324 37192
rect 1152 37064 20448 37088
rect 1152 37024 3688 37064
rect 3728 37024 3770 37064
rect 3810 37024 3852 37064
rect 3892 37024 3934 37064
rect 3974 37024 4016 37064
rect 4056 37024 18808 37064
rect 18848 37024 18890 37064
rect 18930 37024 18972 37064
rect 19012 37024 19054 37064
rect 19094 37024 19136 37064
rect 19176 37024 20448 37064
rect 1152 37000 20448 37024
rect 1851 36896 1893 36905
rect 1851 36856 1852 36896
rect 1892 36856 1893 36896
rect 1851 36847 1893 36856
rect 7947 36896 7989 36905
rect 7947 36856 7948 36896
rect 7988 36856 7989 36896
rect 7947 36847 7989 36856
rect 18363 36896 18405 36905
rect 18363 36856 18364 36896
rect 18404 36856 18405 36896
rect 18363 36847 18405 36856
rect 20139 36896 20181 36905
rect 20139 36856 20140 36896
rect 20180 36856 20181 36896
rect 20139 36847 20181 36856
rect 12363 36812 12405 36821
rect 12363 36772 12364 36812
rect 12404 36772 12405 36812
rect 12363 36763 12405 36772
rect 1227 36728 1269 36737
rect 1227 36688 1228 36728
rect 1268 36688 1269 36728
rect 1227 36679 1269 36688
rect 1611 36728 1653 36737
rect 1611 36688 1612 36728
rect 1652 36688 1653 36728
rect 1611 36679 1653 36688
rect 2763 36728 2805 36737
rect 2763 36688 2764 36728
rect 2804 36688 2805 36728
rect 2763 36679 2805 36688
rect 4203 36728 4245 36737
rect 4203 36688 4204 36728
rect 4244 36688 4245 36728
rect 4203 36679 4245 36688
rect 8218 36728 8276 36729
rect 8218 36688 8227 36728
rect 8267 36688 8276 36728
rect 8218 36687 8276 36688
rect 9771 36728 9813 36737
rect 9771 36688 9772 36728
rect 9812 36688 9813 36728
rect 9771 36679 9813 36688
rect 13707 36728 13749 36737
rect 13707 36688 13708 36728
rect 13748 36688 13749 36728
rect 13707 36679 13749 36688
rect 14859 36728 14901 36737
rect 14859 36688 14860 36728
rect 14900 36688 14901 36728
rect 14859 36679 14901 36688
rect 16011 36728 16053 36737
rect 16011 36688 16012 36728
rect 16052 36688 16053 36728
rect 16011 36679 16053 36688
rect 17739 36728 17781 36737
rect 17739 36688 17740 36728
rect 17780 36688 17781 36728
rect 17739 36679 17781 36688
rect 14300 36663 14342 36672
rect 2266 36644 2324 36645
rect 2266 36604 2275 36644
rect 2315 36604 2324 36644
rect 2266 36603 2324 36604
rect 2379 36644 2421 36653
rect 2379 36604 2380 36644
rect 2420 36604 2421 36644
rect 2379 36595 2421 36604
rect 2859 36644 2901 36653
rect 2859 36604 2860 36644
rect 2900 36604 2901 36644
rect 2859 36595 2901 36604
rect 3331 36644 3389 36645
rect 3331 36604 3340 36644
rect 3380 36604 3389 36644
rect 3331 36603 3389 36604
rect 3819 36644 3877 36645
rect 3819 36604 3828 36644
rect 3868 36604 3877 36644
rect 3819 36603 3877 36604
rect 4875 36644 4917 36653
rect 4875 36604 4876 36644
rect 4916 36604 4917 36644
rect 4875 36595 4917 36604
rect 6115 36644 6173 36645
rect 6115 36604 6124 36644
rect 6164 36604 6173 36644
rect 6115 36603 6173 36604
rect 6507 36644 6549 36653
rect 6507 36604 6508 36644
rect 6548 36604 6549 36644
rect 6507 36595 6549 36604
rect 7747 36644 7805 36645
rect 7747 36604 7756 36644
rect 7796 36604 7805 36644
rect 7747 36603 7805 36604
rect 8086 36644 8128 36653
rect 8086 36604 8087 36644
rect 8127 36604 8128 36644
rect 8086 36595 8128 36604
rect 8331 36644 8373 36653
rect 8331 36604 8332 36644
rect 8372 36604 8373 36644
rect 8331 36595 8373 36604
rect 8794 36644 8852 36645
rect 8794 36604 8803 36644
rect 8843 36604 8852 36644
rect 8794 36603 8852 36604
rect 9283 36644 9341 36645
rect 9283 36604 9292 36644
rect 9332 36604 9341 36644
rect 9283 36603 9341 36604
rect 9867 36644 9909 36653
rect 9867 36604 9868 36644
rect 9908 36604 9909 36644
rect 9867 36595 9909 36604
rect 10251 36644 10293 36653
rect 10251 36604 10252 36644
rect 10292 36604 10293 36644
rect 10251 36595 10293 36604
rect 10361 36644 10419 36645
rect 10361 36604 10370 36644
rect 10410 36604 10419 36644
rect 10361 36603 10419 36604
rect 10923 36644 10965 36653
rect 10923 36604 10924 36644
rect 10964 36604 10965 36644
rect 10923 36595 10965 36604
rect 12163 36644 12221 36645
rect 12163 36604 12172 36644
rect 12212 36604 12221 36644
rect 12163 36603 12221 36604
rect 12730 36644 12788 36645
rect 12730 36604 12739 36644
rect 12779 36604 12788 36644
rect 12730 36603 12788 36604
rect 13219 36644 13277 36645
rect 13219 36604 13228 36644
rect 13268 36604 13277 36644
rect 13219 36603 13277 36604
rect 13803 36644 13845 36653
rect 13803 36604 13804 36644
rect 13844 36604 13845 36644
rect 13803 36595 13845 36604
rect 14187 36644 14229 36653
rect 14187 36604 14188 36644
rect 14228 36604 14229 36644
rect 14300 36623 14301 36663
rect 14341 36623 14342 36663
rect 14300 36614 14342 36623
rect 14667 36644 14709 36653
rect 14187 36595 14229 36604
rect 14667 36604 14668 36644
rect 14708 36604 14709 36644
rect 14667 36595 14709 36604
rect 15514 36644 15572 36645
rect 15514 36604 15523 36644
rect 15563 36604 15572 36644
rect 15514 36603 15572 36604
rect 15627 36644 15669 36653
rect 15627 36604 15628 36644
rect 15668 36604 15669 36644
rect 15627 36595 15669 36604
rect 16107 36644 16149 36653
rect 16107 36604 16108 36644
rect 16148 36604 16149 36644
rect 16107 36595 16149 36604
rect 16579 36644 16637 36645
rect 16579 36604 16588 36644
rect 16628 36604 16637 36644
rect 16579 36603 16637 36604
rect 17098 36644 17156 36645
rect 17098 36604 17107 36644
rect 17147 36604 17156 36644
rect 17098 36603 17156 36604
rect 17398 36644 17440 36653
rect 17398 36604 17399 36644
rect 17439 36604 17440 36644
rect 17398 36595 17440 36604
rect 17530 36644 17588 36645
rect 17530 36604 17539 36644
rect 17579 36604 17588 36644
rect 17530 36603 17588 36604
rect 17643 36644 17685 36653
rect 17643 36604 17644 36644
rect 17684 36604 17685 36644
rect 17643 36595 17685 36604
rect 18211 36644 18269 36645
rect 18211 36604 18220 36644
rect 18260 36604 18269 36644
rect 18211 36603 18269 36604
rect 18507 36644 18549 36653
rect 18507 36604 18508 36644
rect 18548 36604 18549 36644
rect 18507 36595 18549 36604
rect 18699 36644 18741 36653
rect 18699 36604 18700 36644
rect 18740 36604 18741 36644
rect 18699 36595 18741 36604
rect 19939 36644 19997 36645
rect 19939 36604 19948 36644
rect 19988 36604 19997 36644
rect 19939 36603 19997 36604
rect 1467 36560 1509 36569
rect 1467 36520 1468 36560
rect 1508 36520 1509 36560
rect 1467 36511 1509 36520
rect 4443 36560 4485 36569
rect 4443 36520 4444 36560
rect 4484 36520 4485 36560
rect 4443 36511 4485 36520
rect 8602 36560 8660 36561
rect 8602 36520 8611 36560
rect 8651 36520 8660 36560
rect 8602 36519 8660 36520
rect 17917 36560 17959 36569
rect 17917 36520 17918 36560
rect 17958 36520 17959 36560
rect 17917 36511 17959 36520
rect 4011 36476 4053 36485
rect 4011 36436 4012 36476
rect 4052 36436 4053 36476
rect 4011 36427 4053 36436
rect 6315 36476 6357 36485
rect 6315 36436 6316 36476
rect 6356 36436 6357 36476
rect 6315 36427 6357 36436
rect 8410 36476 8468 36477
rect 8410 36436 8419 36476
rect 8459 36436 8468 36476
rect 8410 36435 8468 36436
rect 12555 36476 12597 36485
rect 12555 36436 12556 36476
rect 12596 36436 12597 36476
rect 12555 36427 12597 36436
rect 14523 36476 14565 36485
rect 14523 36436 14524 36476
rect 14564 36436 14565 36476
rect 14523 36427 14565 36436
rect 15099 36476 15141 36485
rect 15099 36436 15100 36476
rect 15140 36436 15141 36476
rect 15099 36427 15141 36436
rect 17259 36476 17301 36485
rect 17259 36436 17260 36476
rect 17300 36436 17301 36476
rect 17259 36427 17301 36436
rect 18010 36476 18068 36477
rect 18010 36436 18019 36476
rect 18059 36436 18068 36476
rect 18010 36435 18068 36436
rect 18123 36476 18165 36485
rect 18123 36436 18124 36476
rect 18164 36436 18165 36476
rect 18123 36427 18165 36436
rect 1152 36308 20452 36332
rect 1152 36268 4928 36308
rect 4968 36268 5010 36308
rect 5050 36268 5092 36308
rect 5132 36268 5174 36308
rect 5214 36268 5256 36308
rect 5296 36268 20048 36308
rect 20088 36268 20130 36308
rect 20170 36268 20212 36308
rect 20252 36268 20294 36308
rect 20334 36268 20376 36308
rect 20416 36268 20452 36308
rect 1152 36244 20452 36268
rect 4011 36140 4053 36149
rect 4011 36100 4012 36140
rect 4052 36100 4053 36140
rect 4011 36091 4053 36100
rect 11595 36140 11637 36149
rect 11595 36100 11596 36140
rect 11636 36100 11637 36140
rect 11595 36091 11637 36100
rect 12730 36140 12788 36141
rect 12730 36100 12739 36140
rect 12779 36100 12788 36140
rect 12730 36099 12788 36100
rect 17818 36140 17876 36141
rect 17818 36100 17827 36140
rect 17867 36100 17876 36140
rect 17818 36099 17876 36100
rect 11866 36056 11924 36057
rect 11866 36016 11875 36056
rect 11915 36016 11924 36056
rect 11866 36015 11924 36016
rect 17931 36056 17973 36065
rect 17931 36016 17932 36056
rect 17972 36016 17973 36056
rect 17931 36007 17973 36016
rect 2266 35972 2324 35973
rect 2266 35932 2275 35972
rect 2315 35932 2324 35972
rect 2266 35931 2324 35932
rect 2384 35972 2426 35981
rect 2384 35932 2385 35972
rect 2425 35932 2426 35972
rect 2384 35923 2426 35932
rect 2763 35972 2805 35981
rect 4491 35972 4533 35981
rect 6123 35972 6165 35981
rect 2763 35932 2764 35972
rect 2804 35932 2805 35972
rect 2763 35923 2805 35932
rect 3339 35963 3381 35972
rect 3339 35923 3340 35963
rect 3380 35923 3381 35963
rect 3339 35914 3381 35923
rect 3819 35963 3861 35972
rect 3819 35923 3820 35963
rect 3860 35923 3861 35963
rect 4491 35932 4492 35972
rect 4532 35932 4533 35972
rect 4491 35923 4533 35932
rect 5739 35963 5781 35972
rect 5739 35923 5740 35963
rect 5780 35923 5781 35963
rect 6123 35932 6124 35972
rect 6164 35932 6165 35972
rect 6123 35923 6165 35932
rect 6298 35972 6356 35973
rect 6298 35932 6307 35972
rect 6347 35932 6356 35972
rect 6298 35931 6356 35932
rect 6891 35972 6933 35981
rect 8523 35972 8565 35981
rect 10155 35972 10197 35981
rect 11787 35972 11829 35981
rect 6891 35932 6892 35972
rect 6932 35932 6933 35972
rect 6891 35923 6933 35932
rect 8139 35963 8181 35972
rect 8139 35923 8140 35963
rect 8180 35923 8181 35963
rect 8523 35932 8524 35972
rect 8564 35932 8565 35972
rect 8523 35923 8565 35932
rect 9771 35963 9813 35972
rect 9771 35923 9772 35963
rect 9812 35923 9813 35963
rect 10155 35932 10156 35972
rect 10196 35932 10197 35972
rect 10155 35923 10197 35932
rect 11403 35963 11445 35972
rect 11403 35923 11404 35963
rect 11444 35923 11445 35963
rect 11787 35932 11788 35972
rect 11828 35932 11829 35972
rect 11787 35923 11829 35932
rect 11962 35972 12020 35973
rect 11962 35932 11971 35972
rect 12011 35932 12020 35972
rect 12250 35972 12308 35973
rect 12630 35972 12688 35973
rect 11962 35931 12020 35932
rect 12082 35940 12124 35949
rect 3819 35914 3861 35923
rect 5739 35914 5781 35923
rect 8139 35914 8181 35923
rect 9771 35914 9813 35923
rect 11403 35914 11445 35923
rect 12082 35900 12083 35940
rect 12123 35900 12124 35940
rect 12250 35932 12259 35972
rect 12299 35932 12308 35972
rect 12250 35931 12308 35932
rect 12363 35963 12405 35972
rect 12363 35923 12364 35963
rect 12404 35923 12405 35963
rect 12363 35914 12405 35923
rect 12507 35963 12549 35972
rect 12507 35923 12508 35963
rect 12548 35923 12549 35963
rect 12630 35932 12639 35972
rect 12679 35932 12688 35972
rect 12630 35931 12688 35932
rect 12768 35972 12826 35973
rect 12768 35932 12777 35972
rect 12817 35932 12826 35972
rect 12768 35931 12826 35932
rect 13035 35972 13077 35981
rect 15723 35972 15765 35981
rect 13035 35932 13036 35972
rect 13076 35932 13077 35972
rect 13035 35923 13077 35932
rect 14283 35963 14325 35972
rect 14283 35923 14284 35963
rect 14324 35923 14325 35963
rect 15723 35932 15724 35972
rect 15764 35932 15765 35972
rect 16107 35972 16149 35981
rect 17725 35972 17767 35981
rect 18315 35972 18357 35981
rect 15723 35923 15765 35932
rect 15963 35930 16005 35939
rect 12507 35914 12549 35923
rect 14283 35914 14325 35923
rect 1227 35888 1269 35897
rect 1227 35848 1228 35888
rect 1268 35848 1269 35888
rect 1227 35839 1269 35848
rect 1611 35888 1653 35897
rect 1611 35848 1612 35888
rect 1652 35848 1653 35888
rect 1611 35839 1653 35848
rect 2859 35888 2901 35897
rect 2859 35848 2860 35888
rect 2900 35848 2901 35888
rect 2859 35839 2901 35848
rect 6699 35888 6741 35897
rect 12082 35891 12124 35900
rect 6699 35848 6700 35888
rect 6740 35848 6741 35888
rect 6699 35839 6741 35848
rect 14859 35888 14901 35897
rect 14859 35848 14860 35888
rect 14900 35848 14901 35888
rect 14859 35839 14901 35848
rect 15099 35888 15141 35897
rect 15099 35848 15100 35888
rect 15140 35848 15141 35888
rect 15099 35839 15141 35848
rect 15435 35888 15477 35897
rect 15435 35848 15436 35888
rect 15476 35848 15477 35888
rect 15435 35839 15477 35848
rect 15627 35888 15669 35897
rect 15627 35848 15628 35888
rect 15668 35848 15669 35888
rect 15627 35839 15669 35848
rect 15842 35888 15884 35897
rect 15842 35848 15843 35888
rect 15883 35848 15884 35888
rect 15963 35890 15964 35930
rect 16004 35890 16005 35930
rect 16107 35932 16108 35972
rect 16148 35932 16149 35972
rect 16107 35923 16149 35932
rect 17355 35963 17397 35972
rect 17355 35923 17356 35963
rect 17396 35923 17397 35963
rect 17725 35932 17726 35972
rect 17766 35932 17767 35972
rect 17725 35923 17767 35932
rect 18027 35963 18069 35972
rect 18027 35923 18028 35963
rect 18068 35923 18069 35963
rect 18315 35932 18316 35972
rect 18356 35932 18357 35972
rect 18315 35923 18357 35932
rect 18586 35972 18644 35973
rect 18586 35932 18595 35972
rect 18635 35932 18644 35972
rect 18586 35931 18644 35932
rect 18699 35972 18741 35981
rect 18699 35932 18700 35972
rect 18740 35932 18741 35972
rect 18699 35923 18741 35932
rect 19083 35972 19125 35981
rect 20362 35972 20420 35973
rect 19083 35932 19084 35972
rect 19124 35932 19125 35972
rect 19083 35923 19125 35932
rect 19659 35963 19701 35972
rect 19659 35923 19660 35963
rect 19700 35923 19701 35963
rect 17355 35914 17397 35923
rect 18027 35914 18069 35923
rect 19659 35914 19701 35923
rect 20139 35963 20181 35972
rect 20139 35923 20140 35963
rect 20180 35923 20181 35963
rect 20362 35932 20371 35972
rect 20411 35932 20420 35972
rect 20362 35931 20420 35932
rect 20139 35914 20181 35923
rect 15963 35881 16005 35890
rect 19179 35888 19221 35897
rect 15842 35839 15884 35848
rect 19179 35848 19180 35888
rect 19220 35848 19221 35888
rect 19179 35839 19221 35848
rect 5931 35804 5973 35813
rect 5931 35764 5932 35804
rect 5972 35764 5973 35804
rect 5931 35755 5973 35764
rect 6298 35804 6356 35805
rect 6298 35764 6307 35804
rect 6347 35764 6356 35804
rect 6298 35763 6356 35764
rect 17547 35804 17589 35813
rect 17547 35764 17548 35804
rect 17588 35764 17589 35804
rect 17547 35755 17589 35764
rect 1467 35720 1509 35729
rect 1467 35680 1468 35720
rect 1508 35680 1509 35720
rect 1467 35671 1509 35680
rect 1851 35720 1893 35729
rect 1851 35680 1852 35720
rect 1892 35680 1893 35720
rect 1851 35671 1893 35680
rect 6459 35720 6501 35729
rect 6459 35680 6460 35720
rect 6500 35680 6501 35720
rect 6459 35671 6501 35680
rect 8331 35720 8373 35729
rect 8331 35680 8332 35720
rect 8372 35680 8373 35720
rect 8331 35671 8373 35680
rect 9963 35720 10005 35729
rect 9963 35680 9964 35720
rect 10004 35680 10005 35720
rect 9963 35671 10005 35680
rect 14475 35720 14517 35729
rect 14475 35680 14476 35720
rect 14516 35680 14517 35720
rect 14475 35671 14517 35680
rect 15195 35720 15237 35729
rect 15195 35680 15196 35720
rect 15236 35680 15237 35720
rect 15195 35671 15237 35680
rect 18171 35720 18213 35729
rect 18171 35680 18172 35720
rect 18212 35680 18213 35720
rect 18171 35671 18213 35680
rect 1152 35552 20448 35576
rect 1152 35512 3688 35552
rect 3728 35512 3770 35552
rect 3810 35512 3852 35552
rect 3892 35512 3934 35552
rect 3974 35512 4016 35552
rect 4056 35512 18808 35552
rect 18848 35512 18890 35552
rect 18930 35512 18972 35552
rect 19012 35512 19054 35552
rect 19094 35512 19136 35552
rect 19176 35512 20448 35552
rect 1152 35488 20448 35512
rect 3531 35384 3573 35393
rect 3531 35344 3532 35384
rect 3572 35344 3573 35384
rect 3531 35335 3573 35344
rect 5355 35384 5397 35393
rect 5355 35344 5356 35384
rect 5396 35344 5397 35384
rect 5355 35335 5397 35344
rect 6987 35384 7029 35393
rect 6987 35344 6988 35384
rect 7028 35344 7029 35384
rect 6987 35335 7029 35344
rect 8043 35384 8085 35393
rect 8043 35344 8044 35384
rect 8084 35344 8085 35384
rect 8043 35335 8085 35344
rect 9675 35384 9717 35393
rect 9675 35344 9676 35384
rect 9716 35344 9717 35384
rect 9675 35335 9717 35344
rect 11403 35384 11445 35393
rect 11403 35344 11404 35384
rect 11444 35344 11445 35384
rect 11403 35335 11445 35344
rect 17931 35384 17973 35393
rect 17931 35344 17932 35384
rect 17972 35344 17973 35384
rect 17931 35335 17973 35344
rect 20235 35384 20277 35393
rect 20235 35344 20236 35384
rect 20276 35344 20277 35384
rect 20235 35335 20277 35344
rect 13035 35300 13077 35309
rect 13035 35260 13036 35300
rect 13076 35260 13077 35300
rect 13035 35251 13077 35260
rect 1227 35216 1269 35225
rect 1227 35176 1228 35216
rect 1268 35176 1269 35216
rect 1227 35167 1269 35176
rect 1611 35216 1653 35225
rect 1611 35176 1612 35216
rect 1652 35176 1653 35216
rect 1611 35167 1653 35176
rect 7323 35216 7365 35225
rect 7323 35176 7324 35216
rect 7364 35176 7365 35216
rect 7323 35167 7365 35176
rect 14283 35216 14325 35225
rect 14283 35176 14284 35216
rect 14324 35176 14325 35216
rect 14283 35167 14325 35176
rect 16491 35216 16533 35225
rect 16491 35176 16492 35216
rect 16532 35176 16533 35216
rect 16491 35167 16533 35176
rect 16762 35216 16820 35217
rect 16762 35176 16771 35216
rect 16811 35176 16820 35216
rect 16762 35175 16820 35176
rect 18315 35216 18357 35225
rect 18315 35176 18316 35216
rect 18356 35176 18357 35216
rect 18315 35167 18357 35176
rect 2091 35132 2133 35141
rect 2091 35092 2092 35132
rect 2132 35092 2133 35132
rect 2091 35083 2133 35092
rect 3331 35132 3389 35133
rect 3331 35092 3340 35132
rect 3380 35092 3389 35132
rect 3331 35091 3389 35092
rect 3915 35132 3957 35141
rect 3915 35092 3916 35132
rect 3956 35092 3957 35132
rect 3915 35083 3957 35092
rect 5155 35132 5213 35133
rect 5155 35092 5164 35132
rect 5204 35092 5213 35132
rect 5155 35091 5213 35092
rect 5547 35132 5589 35141
rect 5547 35092 5548 35132
rect 5588 35092 5589 35132
rect 5547 35083 5589 35092
rect 6787 35132 6845 35133
rect 6787 35092 6796 35132
rect 6836 35092 6845 35132
rect 6787 35091 6845 35092
rect 7179 35132 7221 35141
rect 7179 35092 7180 35132
rect 7220 35092 7221 35132
rect 7179 35083 7221 35092
rect 7483 35132 7541 35133
rect 7483 35092 7492 35132
rect 7532 35092 7541 35132
rect 7483 35091 7541 35092
rect 7642 35132 7700 35133
rect 7642 35092 7651 35132
rect 7691 35092 7700 35132
rect 7642 35091 7700 35092
rect 7767 35132 7809 35141
rect 7767 35092 7768 35132
rect 7808 35092 7809 35132
rect 7767 35083 7809 35092
rect 7930 35132 7988 35133
rect 7930 35092 7939 35132
rect 7979 35092 7988 35132
rect 7930 35091 7988 35092
rect 8032 35132 8090 35133
rect 8032 35092 8041 35132
rect 8081 35092 8090 35132
rect 8032 35091 8090 35092
rect 8259 35132 8317 35133
rect 8259 35092 8268 35132
rect 8308 35092 8317 35132
rect 8259 35091 8317 35092
rect 9475 35132 9533 35133
rect 9475 35092 9484 35132
rect 9524 35092 9533 35132
rect 9475 35091 9533 35092
rect 9963 35132 10005 35141
rect 9963 35092 9964 35132
rect 10004 35092 10005 35132
rect 9963 35083 10005 35092
rect 11203 35132 11261 35133
rect 11203 35092 11212 35132
rect 11252 35092 11261 35132
rect 11203 35091 11261 35092
rect 11595 35132 11637 35141
rect 11595 35092 11596 35132
rect 11636 35092 11637 35132
rect 11595 35083 11637 35092
rect 12835 35132 12893 35133
rect 12835 35092 12844 35132
rect 12884 35092 12893 35132
rect 12835 35091 12893 35092
rect 13227 35132 13269 35141
rect 13227 35092 13228 35132
rect 13268 35092 13269 35132
rect 13227 35083 13269 35092
rect 13366 35132 13408 35141
rect 13366 35092 13367 35132
rect 13407 35092 13408 35132
rect 13366 35083 13408 35092
rect 13786 35132 13844 35133
rect 13786 35092 13795 35132
rect 13835 35092 13844 35132
rect 13786 35091 13844 35092
rect 13899 35132 13941 35141
rect 13899 35092 13900 35132
rect 13940 35092 13941 35132
rect 13899 35083 13941 35092
rect 14379 35132 14421 35141
rect 14379 35092 14380 35132
rect 14420 35092 14421 35132
rect 14379 35083 14421 35092
rect 14851 35132 14909 35133
rect 14851 35092 14860 35132
rect 14900 35092 14909 35132
rect 14851 35091 14909 35092
rect 15339 35132 15397 35133
rect 15339 35092 15348 35132
rect 15388 35092 15397 35132
rect 15339 35091 15397 35092
rect 15819 35132 15861 35141
rect 15819 35092 15820 35132
rect 15860 35092 15861 35132
rect 15819 35083 15861 35092
rect 16011 35132 16053 35141
rect 16011 35092 16012 35132
rect 16052 35092 16053 35132
rect 16011 35083 16053 35092
rect 16155 35132 16197 35141
rect 16155 35092 16156 35132
rect 16196 35092 16197 35132
rect 16155 35083 16197 35092
rect 16282 35132 16340 35133
rect 16282 35092 16291 35132
rect 16331 35092 16340 35132
rect 16282 35091 16340 35092
rect 16395 35132 16437 35141
rect 16395 35092 16396 35132
rect 16436 35092 16437 35132
rect 16395 35083 16437 35092
rect 16630 35132 16672 35141
rect 16630 35092 16631 35132
rect 16671 35092 16672 35132
rect 16630 35083 16672 35092
rect 16875 35132 16917 35141
rect 16875 35092 16876 35132
rect 16916 35092 16917 35132
rect 16875 35083 16917 35092
rect 17259 35132 17301 35141
rect 17259 35092 17260 35132
rect 17300 35092 17301 35132
rect 17259 35083 17301 35092
rect 17530 35132 17588 35133
rect 17530 35092 17539 35132
rect 17579 35092 17588 35132
rect 17530 35091 17588 35092
rect 18603 35132 18645 35141
rect 18603 35092 18604 35132
rect 18644 35092 18645 35132
rect 18603 35083 18645 35092
rect 18795 35132 18837 35141
rect 18795 35092 18796 35132
rect 18836 35092 18837 35132
rect 18795 35083 18837 35092
rect 20035 35132 20093 35133
rect 20035 35092 20044 35132
rect 20084 35092 20093 35132
rect 20035 35091 20093 35092
rect 1467 35048 1509 35057
rect 1467 35008 1468 35048
rect 1508 35008 1509 35048
rect 1467 34999 1509 35008
rect 15915 35048 15957 35057
rect 15915 35008 15916 35048
rect 15956 35008 15957 35048
rect 15915 34999 15957 35008
rect 17643 35048 17685 35057
rect 17643 35008 17644 35048
rect 17684 35008 17685 35048
rect 17643 34999 17685 35008
rect 18075 35048 18117 35057
rect 18075 35008 18076 35048
rect 18116 35008 18117 35048
rect 18075 34999 18117 35008
rect 1851 34964 1893 34973
rect 1851 34924 1852 34964
rect 1892 34924 1893 34964
rect 1851 34915 1893 34924
rect 7546 34964 7604 34965
rect 7546 34924 7555 34964
rect 7595 34924 7604 34964
rect 7546 34923 7604 34924
rect 13515 34964 13557 34973
rect 13515 34924 13516 34964
rect 13556 34924 13557 34964
rect 13515 34915 13557 34924
rect 15531 34964 15573 34973
rect 15531 34924 15532 34964
rect 15572 34924 15573 34964
rect 15531 34915 15573 34924
rect 16954 34964 17012 34965
rect 16954 34924 16963 34964
rect 17003 34924 17012 34964
rect 16954 34923 17012 34924
rect 18459 34964 18501 34973
rect 18459 34924 18460 34964
rect 18500 34924 18501 34964
rect 18459 34915 18501 34924
rect 1152 34796 20452 34820
rect 1152 34756 4928 34796
rect 4968 34756 5010 34796
rect 5050 34756 5092 34796
rect 5132 34756 5174 34796
rect 5214 34756 5256 34796
rect 5296 34756 20048 34796
rect 20088 34756 20130 34796
rect 20170 34756 20212 34796
rect 20252 34756 20294 34796
rect 20334 34756 20376 34796
rect 20416 34756 20452 34796
rect 1152 34732 20452 34756
rect 17242 34628 17300 34629
rect 17242 34588 17251 34628
rect 17291 34588 17300 34628
rect 17242 34587 17300 34588
rect 11146 34544 11204 34545
rect 11146 34504 11155 34544
rect 11195 34504 11204 34544
rect 11146 34503 11204 34504
rect 12315 34544 12357 34553
rect 12315 34504 12316 34544
rect 12356 34504 12357 34544
rect 12315 34495 12357 34504
rect 13899 34544 13941 34553
rect 13899 34504 13900 34544
rect 13940 34504 13941 34544
rect 13899 34495 13941 34504
rect 16635 34544 16677 34553
rect 16635 34504 16636 34544
rect 16676 34504 16677 34544
rect 16635 34495 16677 34504
rect 17462 34544 17504 34553
rect 17462 34504 17463 34544
rect 17503 34504 17504 34544
rect 17462 34495 17504 34504
rect 19083 34544 19125 34553
rect 19083 34504 19084 34544
rect 19124 34504 19125 34544
rect 19083 34495 19125 34504
rect 19611 34544 19653 34553
rect 19611 34504 19612 34544
rect 19652 34504 19653 34544
rect 19611 34495 19653 34504
rect 19995 34544 20037 34553
rect 19995 34504 19996 34544
rect 20036 34504 20037 34544
rect 19995 34495 20037 34504
rect 20379 34544 20421 34553
rect 20379 34504 20380 34544
rect 20420 34504 20421 34544
rect 20379 34495 20421 34504
rect 2266 34460 2324 34461
rect 2266 34420 2275 34460
rect 2315 34420 2324 34460
rect 2266 34419 2324 34420
rect 2571 34460 2613 34469
rect 2571 34420 2572 34460
rect 2612 34420 2613 34460
rect 2571 34411 2613 34420
rect 2842 34460 2900 34461
rect 2842 34420 2851 34460
rect 2891 34420 2900 34460
rect 2842 34419 2900 34420
rect 2955 34460 2997 34469
rect 2955 34420 2956 34460
rect 2996 34420 2997 34460
rect 2955 34411 2997 34420
rect 3339 34460 3381 34469
rect 6027 34460 6069 34469
rect 7659 34460 7701 34469
rect 9370 34460 9428 34461
rect 3339 34420 3340 34460
rect 3380 34420 3381 34460
rect 3339 34411 3381 34420
rect 3915 34451 3957 34460
rect 3915 34411 3916 34451
rect 3956 34411 3957 34451
rect 3915 34402 3957 34411
rect 4395 34451 4437 34460
rect 4395 34411 4396 34451
rect 4436 34411 4437 34451
rect 6027 34420 6028 34460
rect 6068 34420 6069 34460
rect 6027 34411 6069 34420
rect 7275 34451 7317 34460
rect 7275 34411 7276 34451
rect 7316 34411 7317 34451
rect 7659 34420 7660 34460
rect 7700 34420 7701 34460
rect 7659 34411 7701 34420
rect 8907 34451 8949 34460
rect 8907 34411 8908 34451
rect 8948 34411 8949 34451
rect 9370 34420 9379 34460
rect 9419 34420 9428 34460
rect 9370 34419 9428 34420
rect 9483 34460 9525 34469
rect 9483 34420 9484 34460
rect 9524 34420 9525 34460
rect 9483 34411 9525 34420
rect 9867 34460 9909 34469
rect 12459 34460 12501 34469
rect 14266 34460 14324 34461
rect 9867 34420 9868 34460
rect 9908 34420 9909 34460
rect 9867 34411 9909 34420
rect 10443 34451 10485 34460
rect 10443 34411 10444 34451
rect 10484 34411 10485 34451
rect 4395 34402 4437 34411
rect 7275 34402 7317 34411
rect 8907 34402 8949 34411
rect 10443 34402 10485 34411
rect 10923 34451 10965 34460
rect 10923 34411 10924 34451
rect 10964 34411 10965 34451
rect 12459 34420 12460 34460
rect 12500 34420 12501 34460
rect 12459 34411 12501 34420
rect 13707 34451 13749 34460
rect 13707 34411 13708 34451
rect 13748 34411 13749 34451
rect 14266 34420 14275 34460
rect 14315 34420 14324 34460
rect 14266 34419 14324 34420
rect 14379 34460 14421 34469
rect 14379 34420 14380 34460
rect 14420 34420 14421 34460
rect 14379 34411 14421 34420
rect 14763 34460 14805 34469
rect 17146 34460 17204 34461
rect 14763 34420 14764 34460
rect 14804 34420 14805 34460
rect 14763 34411 14805 34420
rect 15339 34451 15381 34460
rect 15339 34411 15340 34451
rect 15380 34411 15381 34451
rect 10923 34402 10965 34411
rect 13707 34402 13749 34411
rect 15339 34402 15381 34411
rect 15819 34451 15861 34460
rect 15819 34411 15820 34451
rect 15860 34411 15861 34451
rect 17146 34420 17155 34460
rect 17195 34420 17204 34460
rect 17146 34419 17204 34420
rect 17643 34460 17685 34469
rect 17643 34420 17644 34460
rect 17684 34420 17685 34460
rect 17643 34411 17685 34420
rect 18891 34451 18933 34460
rect 18891 34411 18892 34451
rect 18932 34411 18933 34451
rect 15819 34402 15861 34411
rect 18891 34402 18933 34411
rect 1227 34376 1269 34385
rect 1227 34336 1228 34376
rect 1268 34336 1269 34376
rect 1227 34327 1269 34336
rect 1611 34376 1653 34385
rect 1611 34336 1612 34376
rect 1652 34336 1653 34376
rect 1611 34327 1653 34336
rect 1851 34376 1893 34385
rect 1851 34336 1852 34376
rect 1892 34336 1893 34376
rect 1851 34327 1893 34336
rect 3435 34376 3477 34385
rect 3435 34336 3436 34376
rect 3476 34336 3477 34376
rect 3435 34327 3477 34336
rect 4618 34376 4676 34377
rect 4618 34336 4627 34376
rect 4667 34336 4676 34376
rect 4618 34335 4676 34336
rect 4779 34376 4821 34385
rect 4779 34336 4780 34376
rect 4820 34336 4821 34376
rect 4779 34327 4821 34336
rect 5163 34376 5205 34385
rect 5163 34336 5164 34376
rect 5204 34336 5205 34376
rect 5163 34327 5205 34336
rect 5403 34376 5445 34385
rect 5403 34336 5404 34376
rect 5444 34336 5445 34376
rect 5403 34327 5445 34336
rect 5835 34376 5877 34385
rect 5835 34336 5836 34376
rect 5876 34336 5877 34376
rect 5835 34327 5877 34336
rect 9963 34376 10005 34385
rect 9963 34336 9964 34376
rect 10004 34336 10005 34376
rect 9963 34327 10005 34336
rect 12075 34376 12117 34385
rect 12075 34336 12076 34376
rect 12116 34336 12117 34376
rect 12075 34327 12117 34336
rect 14859 34376 14901 34385
rect 14859 34336 14860 34376
rect 14900 34336 14901 34376
rect 14859 34327 14901 34336
rect 16395 34376 16437 34385
rect 16395 34336 16396 34376
rect 16436 34336 16437 34376
rect 16395 34327 16437 34336
rect 16779 34376 16821 34385
rect 16779 34336 16780 34376
rect 16820 34336 16821 34376
rect 16779 34327 16821 34336
rect 17019 34376 17061 34385
rect 17019 34336 17020 34376
rect 17060 34336 17061 34376
rect 17019 34327 17061 34336
rect 19371 34376 19413 34385
rect 19371 34336 19372 34376
rect 19412 34336 19413 34376
rect 19371 34327 19413 34336
rect 19755 34376 19797 34385
rect 19755 34336 19756 34376
rect 19796 34336 19797 34376
rect 19755 34327 19797 34336
rect 20139 34376 20181 34385
rect 20139 34336 20140 34376
rect 20180 34336 20181 34376
rect 20139 34327 20181 34336
rect 5019 34292 5061 34301
rect 5019 34252 5020 34292
rect 5060 34252 5061 34292
rect 5019 34243 5061 34252
rect 1467 34208 1509 34217
rect 1467 34168 1468 34208
rect 1508 34168 1509 34208
rect 1467 34159 1509 34168
rect 2571 34208 2613 34217
rect 2571 34168 2572 34208
rect 2612 34168 2613 34208
rect 2571 34159 2613 34168
rect 5595 34208 5637 34217
rect 5595 34168 5596 34208
rect 5636 34168 5637 34208
rect 5595 34159 5637 34168
rect 7467 34208 7509 34217
rect 7467 34168 7468 34208
rect 7508 34168 7509 34208
rect 7467 34159 7509 34168
rect 9099 34208 9141 34217
rect 9099 34168 9100 34208
rect 9140 34168 9141 34208
rect 9099 34159 9141 34168
rect 16042 34208 16100 34209
rect 16042 34168 16051 34208
rect 16091 34168 16100 34208
rect 16042 34167 16100 34168
rect 17451 34208 17493 34217
rect 17451 34168 17452 34208
rect 17492 34168 17493 34208
rect 17451 34159 17493 34168
rect 1152 34040 20448 34064
rect 1152 34000 3688 34040
rect 3728 34000 3770 34040
rect 3810 34000 3852 34040
rect 3892 34000 3934 34040
rect 3974 34000 4016 34040
rect 4056 34000 18808 34040
rect 18848 34000 18890 34040
rect 18930 34000 18972 34040
rect 19012 34000 19054 34040
rect 19094 34000 19136 34040
rect 19176 34000 20448 34040
rect 1152 33976 20448 34000
rect 2667 33872 2709 33881
rect 2667 33832 2668 33872
rect 2708 33832 2709 33872
rect 2667 33823 2709 33832
rect 5835 33872 5877 33881
rect 5835 33832 5836 33872
rect 5876 33832 5877 33872
rect 5835 33823 5877 33832
rect 7467 33872 7509 33881
rect 7467 33832 7468 33872
rect 7508 33832 7509 33872
rect 7467 33823 7509 33832
rect 15627 33872 15669 33881
rect 15627 33832 15628 33872
rect 15668 33832 15669 33872
rect 15627 33823 15669 33832
rect 16875 33872 16917 33881
rect 16875 33832 16876 33872
rect 16916 33832 16917 33872
rect 16875 33823 16917 33832
rect 11163 33788 11205 33797
rect 11163 33748 11164 33788
rect 11204 33748 11205 33788
rect 11163 33739 11205 33748
rect 4011 33704 4053 33713
rect 4011 33664 4012 33704
rect 4052 33664 4053 33704
rect 3128 33653 3186 33658
rect 4011 33655 4053 33664
rect 9867 33704 9909 33713
rect 9867 33664 9868 33704
rect 9908 33664 9909 33704
rect 9867 33655 9909 33664
rect 1227 33620 1269 33629
rect 1227 33580 1228 33620
rect 1268 33580 1269 33620
rect 1227 33571 1269 33580
rect 2467 33620 2525 33621
rect 2467 33580 2476 33620
rect 2516 33580 2525 33620
rect 2467 33579 2525 33580
rect 3018 33620 3076 33621
rect 3018 33580 3027 33620
rect 3067 33580 3076 33620
rect 3128 33613 3137 33653
rect 3177 33613 3186 33653
rect 3128 33612 3186 33613
rect 3239 33620 3297 33621
rect 3018 33579 3076 33580
rect 3239 33580 3248 33620
rect 3288 33580 3297 33620
rect 3239 33579 3297 33580
rect 3811 33620 3869 33621
rect 3811 33580 3820 33620
rect 3860 33580 3869 33620
rect 3811 33579 3869 33580
rect 4395 33620 4437 33629
rect 4395 33580 4396 33620
rect 4436 33580 4437 33620
rect 4395 33571 4437 33580
rect 5635 33620 5693 33621
rect 5635 33580 5644 33620
rect 5684 33580 5693 33620
rect 5635 33579 5693 33580
rect 6027 33620 6069 33629
rect 6027 33580 6028 33620
rect 6068 33580 6069 33620
rect 6027 33571 6069 33580
rect 7267 33620 7325 33621
rect 7267 33580 7276 33620
rect 7316 33580 7325 33620
rect 7267 33579 7325 33580
rect 7659 33620 7701 33629
rect 7659 33580 7660 33620
rect 7700 33580 7701 33620
rect 7659 33571 7701 33580
rect 8899 33620 8957 33621
rect 8899 33580 8908 33620
rect 8948 33580 8957 33620
rect 8899 33579 8957 33580
rect 9370 33620 9428 33621
rect 9370 33580 9379 33620
rect 9419 33580 9428 33620
rect 9370 33579 9428 33580
rect 9483 33620 9525 33629
rect 9483 33580 9484 33620
rect 9524 33580 9525 33620
rect 9483 33571 9525 33580
rect 9963 33620 10005 33629
rect 9963 33580 9964 33620
rect 10004 33580 10005 33620
rect 9963 33571 10005 33580
rect 10435 33620 10493 33621
rect 10435 33580 10444 33620
rect 10484 33580 10493 33620
rect 10435 33579 10493 33580
rect 10923 33620 10981 33621
rect 10923 33580 10932 33620
rect 10972 33580 10981 33620
rect 10923 33579 10981 33580
rect 12555 33620 12597 33629
rect 12555 33580 12556 33620
rect 12596 33580 12597 33620
rect 12555 33571 12597 33580
rect 13795 33620 13853 33621
rect 13795 33580 13804 33620
rect 13844 33580 13853 33620
rect 13795 33579 13853 33580
rect 14187 33620 14229 33629
rect 14187 33580 14188 33620
rect 14228 33580 14229 33620
rect 14187 33571 14229 33580
rect 15427 33620 15485 33621
rect 15427 33580 15436 33620
rect 15476 33580 15485 33620
rect 15427 33579 15485 33580
rect 16203 33620 16245 33629
rect 16203 33580 16204 33620
rect 16244 33580 16245 33620
rect 16203 33571 16245 33580
rect 16474 33620 16532 33621
rect 16474 33580 16483 33620
rect 16523 33580 16532 33620
rect 16474 33579 16532 33580
rect 17067 33620 17109 33629
rect 17067 33580 17068 33620
rect 17108 33580 17109 33620
rect 17067 33571 17109 33580
rect 18307 33620 18365 33621
rect 18307 33580 18316 33620
rect 18356 33580 18365 33620
rect 18307 33579 18365 33580
rect 18699 33620 18741 33629
rect 18699 33580 18700 33620
rect 18740 33580 18741 33620
rect 18699 33571 18741 33580
rect 19939 33620 19997 33621
rect 19939 33580 19948 33620
rect 19988 33580 19997 33620
rect 19939 33579 19997 33580
rect 3517 33536 3559 33545
rect 3517 33496 3518 33536
rect 3558 33496 3559 33536
rect 3517 33487 3559 33496
rect 9099 33536 9141 33545
rect 9099 33496 9100 33536
rect 9140 33496 9141 33536
rect 9099 33487 9141 33496
rect 16587 33536 16629 33545
rect 16587 33496 16588 33536
rect 16628 33496 16629 33536
rect 16587 33487 16629 33496
rect 2859 33452 2901 33461
rect 2859 33412 2860 33452
rect 2900 33412 2901 33452
rect 2859 33403 2901 33412
rect 3610 33452 3668 33453
rect 3610 33412 3619 33452
rect 3659 33412 3668 33452
rect 3610 33411 3668 33412
rect 3723 33452 3765 33461
rect 3723 33412 3724 33452
rect 3764 33412 3765 33452
rect 3723 33403 3765 33412
rect 4251 33452 4293 33461
rect 4251 33412 4252 33452
rect 4292 33412 4293 33452
rect 4251 33403 4293 33412
rect 11115 33452 11157 33461
rect 11115 33412 11116 33452
rect 11156 33412 11157 33452
rect 11115 33403 11157 33412
rect 13995 33452 14037 33461
rect 13995 33412 13996 33452
rect 14036 33412 14037 33452
rect 13995 33403 14037 33412
rect 18507 33452 18549 33461
rect 18507 33412 18508 33452
rect 18548 33412 18549 33452
rect 18507 33403 18549 33412
rect 20139 33452 20181 33461
rect 20139 33412 20140 33452
rect 20180 33412 20181 33452
rect 20139 33403 20181 33412
rect 1152 33284 20452 33308
rect 1152 33244 4928 33284
rect 4968 33244 5010 33284
rect 5050 33244 5092 33284
rect 5132 33244 5174 33284
rect 5214 33244 5256 33284
rect 5296 33244 20048 33284
rect 20088 33244 20130 33284
rect 20170 33244 20212 33284
rect 20252 33244 20294 33284
rect 20334 33244 20376 33284
rect 20416 33244 20452 33284
rect 1152 33220 20452 33244
rect 3051 33116 3093 33125
rect 3051 33076 3052 33116
rect 3092 33076 3093 33116
rect 3051 33067 3093 33076
rect 4683 33116 4725 33125
rect 4683 33076 4684 33116
rect 4724 33076 4725 33116
rect 4683 33067 4725 33076
rect 7947 33116 7989 33125
rect 7947 33076 7948 33116
rect 7988 33076 7989 33116
rect 7947 33067 7989 33076
rect 10155 33116 10197 33125
rect 10155 33076 10156 33116
rect 10196 33076 10197 33116
rect 10155 33067 10197 33076
rect 15435 33116 15477 33125
rect 15435 33076 15436 33116
rect 15476 33076 15477 33116
rect 15435 33067 15477 33076
rect 17163 33116 17205 33125
rect 17163 33076 17164 33116
rect 17204 33076 17205 33116
rect 17163 33067 17205 33076
rect 20139 33116 20181 33125
rect 20139 33076 20140 33116
rect 20180 33076 20181 33116
rect 20139 33067 20181 33076
rect 13419 33032 13461 33041
rect 13419 32992 13420 33032
rect 13460 32992 13461 33032
rect 13419 32983 13461 32992
rect 1611 32948 1653 32957
rect 3243 32948 3285 32957
rect 4971 32948 5013 32957
rect 1611 32908 1612 32948
rect 1652 32908 1653 32948
rect 1611 32899 1653 32908
rect 2859 32939 2901 32948
rect 2859 32899 2860 32939
rect 2900 32899 2901 32939
rect 3243 32908 3244 32948
rect 3284 32908 3285 32948
rect 3243 32899 3285 32908
rect 4491 32939 4533 32948
rect 4491 32899 4492 32939
rect 4532 32899 4533 32939
rect 4971 32908 4972 32948
rect 5012 32908 5013 32948
rect 4971 32899 5013 32908
rect 5242 32948 5300 32949
rect 5242 32908 5251 32948
rect 5291 32908 5300 32948
rect 5242 32907 5300 32908
rect 5360 32948 5402 32957
rect 5360 32908 5361 32948
rect 5401 32908 5402 32948
rect 5360 32899 5402 32908
rect 5739 32948 5781 32957
rect 7659 32948 7701 32957
rect 5739 32908 5740 32948
rect 5780 32908 5781 32948
rect 5739 32899 5781 32908
rect 6315 32939 6357 32948
rect 6315 32899 6316 32939
rect 6356 32899 6357 32939
rect 2859 32890 2901 32899
rect 4491 32890 4533 32899
rect 6315 32890 6357 32899
rect 6795 32939 6837 32948
rect 6795 32899 6796 32939
rect 6836 32899 6837 32939
rect 7659 32908 7660 32948
rect 7700 32908 7701 32948
rect 7659 32899 7701 32908
rect 7793 32948 7851 32949
rect 7793 32908 7802 32948
rect 7842 32908 7851 32948
rect 7793 32907 7851 32908
rect 8139 32948 8181 32957
rect 8139 32908 8140 32948
rect 8180 32908 8181 32948
rect 8139 32899 8181 32908
rect 8254 32948 8296 32957
rect 8254 32908 8255 32948
rect 8295 32908 8296 32948
rect 8254 32899 8296 32908
rect 8427 32948 8469 32957
rect 8427 32908 8428 32948
rect 8468 32908 8469 32948
rect 8427 32899 8469 32908
rect 8715 32948 8757 32957
rect 11787 32948 11829 32957
rect 8715 32908 8716 32948
rect 8756 32908 8757 32948
rect 8715 32899 8757 32908
rect 9963 32939 10005 32948
rect 9963 32899 9964 32939
rect 10004 32899 10005 32939
rect 6795 32890 6837 32899
rect 9963 32890 10005 32899
rect 10539 32939 10581 32948
rect 10539 32899 10540 32939
rect 10580 32899 10581 32939
rect 11787 32908 11788 32948
rect 11828 32908 11829 32948
rect 11787 32899 11829 32908
rect 11979 32948 12021 32957
rect 13690 32948 13748 32949
rect 11979 32908 11980 32948
rect 12020 32908 12021 32948
rect 11979 32899 12021 32908
rect 13227 32939 13269 32948
rect 13227 32899 13228 32939
rect 13268 32899 13269 32939
rect 13690 32908 13699 32948
rect 13739 32908 13748 32948
rect 13690 32907 13748 32908
rect 13803 32948 13845 32957
rect 13803 32908 13804 32948
rect 13844 32908 13845 32948
rect 13803 32899 13845 32908
rect 14187 32948 14229 32957
rect 15723 32948 15765 32957
rect 18394 32948 18452 32949
rect 14187 32908 14188 32948
rect 14228 32908 14229 32948
rect 14187 32899 14229 32908
rect 14763 32939 14805 32948
rect 14763 32899 14764 32939
rect 14804 32899 14805 32939
rect 10539 32890 10581 32899
rect 13227 32890 13269 32899
rect 14763 32890 14805 32899
rect 15243 32939 15285 32948
rect 15243 32899 15244 32939
rect 15284 32899 15285 32939
rect 15723 32908 15724 32948
rect 15764 32908 15765 32948
rect 15723 32899 15765 32908
rect 16971 32939 17013 32948
rect 16971 32899 16972 32939
rect 17012 32899 17013 32939
rect 18394 32908 18403 32948
rect 18443 32908 18452 32948
rect 18394 32907 18452 32908
rect 18507 32948 18549 32957
rect 18507 32908 18508 32948
rect 18548 32908 18549 32948
rect 18507 32899 18549 32908
rect 18891 32948 18933 32957
rect 18891 32908 18892 32948
rect 18932 32908 18933 32948
rect 18891 32899 18933 32908
rect 19467 32939 19509 32948
rect 19467 32899 19468 32939
rect 19508 32899 19509 32939
rect 15243 32890 15285 32899
rect 16971 32890 17013 32899
rect 19467 32890 19509 32899
rect 19947 32939 19989 32948
rect 19947 32899 19948 32939
rect 19988 32899 19989 32939
rect 19947 32890 19989 32899
rect 1227 32864 1269 32873
rect 1227 32824 1228 32864
rect 1268 32824 1269 32864
rect 1227 32815 1269 32824
rect 5835 32864 5877 32873
rect 5835 32824 5836 32864
rect 5876 32824 5877 32864
rect 5835 32815 5877 32824
rect 7275 32864 7317 32873
rect 7275 32824 7276 32864
rect 7316 32824 7317 32864
rect 7275 32815 7317 32824
rect 14283 32864 14325 32873
rect 14283 32824 14284 32864
rect 14324 32824 14325 32864
rect 14283 32815 14325 32824
rect 17547 32864 17589 32873
rect 17547 32824 17548 32864
rect 17588 32824 17589 32864
rect 17547 32815 17589 32824
rect 17931 32864 17973 32873
rect 17931 32824 17932 32864
rect 17972 32824 17973 32864
rect 17931 32815 17973 32824
rect 18987 32864 19029 32873
rect 18987 32824 18988 32864
rect 19028 32824 19029 32864
rect 18987 32815 19029 32824
rect 8139 32780 8181 32789
rect 8139 32740 8140 32780
rect 8180 32740 8181 32780
rect 8139 32731 8181 32740
rect 1467 32696 1509 32705
rect 1467 32656 1468 32696
rect 1508 32656 1509 32696
rect 1467 32647 1509 32656
rect 4827 32696 4869 32705
rect 4827 32656 4828 32696
rect 4868 32656 4869 32696
rect 4827 32647 4869 32656
rect 7018 32696 7076 32697
rect 7018 32656 7027 32696
rect 7067 32656 7076 32696
rect 7018 32655 7076 32656
rect 7515 32696 7557 32705
rect 7515 32656 7516 32696
rect 7556 32656 7557 32696
rect 7515 32647 7557 32656
rect 10347 32696 10389 32705
rect 10347 32656 10348 32696
rect 10388 32656 10389 32696
rect 10347 32647 10389 32656
rect 17307 32696 17349 32705
rect 17307 32656 17308 32696
rect 17348 32656 17349 32696
rect 17307 32647 17349 32656
rect 17691 32696 17733 32705
rect 17691 32656 17692 32696
rect 17732 32656 17733 32696
rect 17691 32647 17733 32656
rect 1152 32528 20448 32552
rect 1152 32488 3688 32528
rect 3728 32488 3770 32528
rect 3810 32488 3852 32528
rect 3892 32488 3934 32528
rect 3974 32488 4016 32528
rect 4056 32488 18808 32528
rect 18848 32488 18890 32528
rect 18930 32488 18972 32528
rect 19012 32488 19054 32528
rect 19094 32488 19136 32528
rect 19176 32488 20448 32528
rect 1152 32464 20448 32488
rect 4779 32360 4821 32369
rect 4779 32320 4780 32360
rect 4820 32320 4821 32360
rect 4779 32311 4821 32320
rect 6411 32360 6453 32369
rect 6411 32320 6412 32360
rect 6452 32320 6453 32360
rect 6411 32311 6453 32320
rect 7899 32360 7941 32369
rect 7899 32320 7900 32360
rect 7940 32320 7941 32360
rect 7899 32311 7941 32320
rect 12027 32360 12069 32369
rect 12027 32320 12028 32360
rect 12068 32320 12069 32360
rect 12027 32311 12069 32320
rect 17067 32360 17109 32369
rect 17067 32320 17068 32360
rect 17108 32320 17109 32360
rect 17067 32311 17109 32320
rect 18171 32360 18213 32369
rect 18171 32320 18172 32360
rect 18212 32320 18213 32360
rect 18171 32311 18213 32320
rect 2667 32276 2709 32285
rect 2667 32236 2668 32276
rect 2708 32236 2709 32276
rect 2667 32227 2709 32236
rect 6603 32192 6645 32201
rect 3090 32183 3136 32192
rect 3090 32143 3091 32183
rect 3131 32143 3136 32183
rect 6603 32152 6604 32192
rect 6644 32152 6645 32192
rect 6603 32143 6645 32152
rect 6987 32192 7029 32201
rect 6987 32152 6988 32192
rect 7028 32152 7029 32192
rect 6987 32143 7029 32152
rect 7371 32192 7413 32201
rect 7371 32152 7372 32192
rect 7412 32152 7413 32192
rect 7371 32143 7413 32152
rect 8139 32192 8181 32201
rect 8139 32152 8140 32192
rect 8180 32152 8181 32192
rect 8139 32143 8181 32152
rect 8331 32192 8373 32201
rect 8331 32152 8332 32192
rect 8372 32152 8373 32192
rect 8331 32143 8373 32152
rect 8715 32192 8757 32201
rect 8715 32152 8716 32192
rect 8756 32152 8757 32192
rect 8715 32143 8757 32152
rect 8955 32192 8997 32201
rect 8955 32152 8956 32192
rect 8996 32152 8997 32192
rect 8955 32143 8997 32152
rect 9195 32192 9237 32201
rect 9195 32152 9196 32192
rect 9236 32152 9237 32192
rect 9195 32143 9237 32152
rect 10251 32192 10293 32201
rect 10251 32152 10252 32192
rect 10292 32152 10293 32192
rect 10251 32143 10293 32152
rect 11787 32192 11829 32201
rect 11787 32152 11788 32192
rect 11828 32152 11829 32192
rect 11787 32143 11829 32152
rect 12363 32192 12405 32201
rect 12363 32152 12364 32192
rect 12404 32152 12405 32192
rect 12363 32143 12405 32152
rect 14187 32192 14229 32201
rect 14187 32152 14188 32192
rect 14228 32152 14229 32192
rect 14187 32143 14229 32152
rect 17259 32192 17301 32201
rect 17259 32152 17260 32192
rect 17300 32152 17301 32192
rect 17259 32143 17301 32152
rect 17931 32192 17973 32201
rect 17931 32152 17932 32192
rect 17972 32152 17973 32192
rect 17931 32143 17973 32152
rect 18891 32192 18933 32201
rect 18891 32152 18892 32192
rect 18932 32152 18933 32192
rect 18891 32143 18933 32152
rect 3090 32134 3136 32143
rect 1227 32108 1269 32117
rect 1227 32068 1228 32108
rect 1268 32068 1269 32108
rect 1227 32059 1269 32068
rect 2467 32108 2525 32109
rect 2467 32068 2476 32108
rect 2516 32068 2525 32108
rect 2467 32067 2525 32068
rect 2954 32108 2996 32117
rect 2954 32068 2955 32108
rect 2995 32068 2996 32108
rect 2954 32059 2996 32068
rect 3184 32108 3242 32109
rect 3184 32068 3193 32108
rect 3233 32068 3242 32108
rect 3184 32067 3242 32068
rect 3339 32108 3381 32117
rect 3339 32068 3340 32108
rect 3380 32068 3381 32108
rect 3339 32059 3381 32068
rect 4579 32108 4637 32109
rect 4579 32068 4588 32108
rect 4628 32068 4637 32108
rect 4579 32067 4637 32068
rect 4971 32108 5013 32117
rect 4971 32068 4972 32108
rect 5012 32068 5013 32108
rect 4971 32059 5013 32068
rect 6211 32108 6269 32109
rect 6211 32068 6220 32108
rect 6260 32068 6269 32108
rect 6211 32067 6269 32068
rect 9754 32108 9812 32109
rect 9754 32068 9763 32108
rect 9803 32068 9812 32108
rect 9754 32067 9812 32068
rect 9867 32108 9909 32117
rect 9867 32068 9868 32108
rect 9908 32068 9909 32108
rect 9867 32059 9909 32068
rect 10347 32108 10389 32117
rect 10347 32068 10348 32108
rect 10388 32068 10389 32108
rect 10347 32059 10389 32068
rect 10819 32108 10877 32109
rect 10819 32068 10828 32108
rect 10868 32068 10877 32108
rect 10819 32067 10877 32068
rect 11338 32108 11396 32109
rect 11338 32068 11347 32108
rect 11387 32068 11396 32108
rect 11338 32067 11396 32068
rect 13690 32108 13748 32109
rect 13690 32068 13699 32108
rect 13739 32068 13748 32108
rect 13690 32067 13748 32068
rect 13803 32108 13845 32117
rect 13803 32068 13804 32108
rect 13844 32068 13845 32108
rect 13803 32059 13845 32068
rect 14283 32108 14325 32117
rect 14283 32068 14284 32108
rect 14324 32068 14325 32108
rect 14283 32059 14325 32068
rect 14755 32108 14813 32109
rect 14755 32068 14764 32108
rect 14804 32068 14813 32108
rect 14755 32067 14813 32068
rect 15243 32108 15301 32109
rect 15243 32068 15252 32108
rect 15292 32068 15301 32108
rect 15243 32067 15301 32068
rect 15627 32108 15669 32117
rect 15627 32068 15628 32108
rect 15668 32068 15669 32108
rect 15627 32059 15669 32068
rect 16867 32108 16925 32109
rect 16867 32068 16876 32108
rect 16916 32068 16925 32108
rect 16867 32067 16925 32068
rect 18394 32108 18452 32109
rect 18394 32068 18403 32108
rect 18443 32068 18452 32108
rect 18394 32067 18452 32068
rect 18507 32108 18549 32117
rect 18507 32068 18508 32108
rect 18548 32068 18549 32108
rect 18507 32059 18549 32068
rect 18987 32108 19029 32117
rect 18987 32068 18988 32108
rect 19028 32068 19029 32108
rect 18987 32059 19029 32068
rect 19459 32108 19517 32109
rect 19459 32068 19468 32108
rect 19508 32068 19517 32108
rect 19459 32067 19517 32068
rect 19947 32108 20005 32109
rect 19947 32068 19956 32108
rect 19996 32068 20005 32108
rect 19947 32067 20005 32068
rect 2859 31940 2901 31949
rect 2859 31900 2860 31940
rect 2900 31900 2901 31940
rect 2859 31891 2901 31900
rect 6843 31940 6885 31949
rect 6843 31900 6844 31940
rect 6884 31900 6885 31940
rect 6843 31891 6885 31900
rect 7227 31940 7269 31949
rect 7227 31900 7228 31940
rect 7268 31900 7269 31940
rect 7227 31891 7269 31900
rect 7611 31940 7653 31949
rect 7611 31900 7612 31940
rect 7652 31900 7653 31940
rect 7611 31891 7653 31900
rect 8571 31940 8613 31949
rect 8571 31900 8572 31940
rect 8612 31900 8613 31940
rect 8571 31891 8613 31900
rect 9435 31940 9477 31949
rect 9435 31900 9436 31940
rect 9476 31900 9477 31940
rect 9435 31891 9477 31900
rect 11499 31940 11541 31949
rect 11499 31900 11500 31940
rect 11540 31900 11541 31940
rect 11499 31891 11541 31900
rect 12123 31940 12165 31949
rect 12123 31900 12124 31940
rect 12164 31900 12165 31940
rect 12123 31891 12165 31900
rect 15435 31940 15477 31949
rect 15435 31900 15436 31940
rect 15476 31900 15477 31940
rect 15435 31891 15477 31900
rect 17499 31940 17541 31949
rect 17499 31900 17500 31940
rect 17540 31900 17541 31940
rect 17499 31891 17541 31900
rect 20139 31940 20181 31949
rect 20139 31900 20140 31940
rect 20180 31900 20181 31940
rect 20139 31891 20181 31900
rect 1152 31772 20452 31796
rect 1152 31732 4928 31772
rect 4968 31732 5010 31772
rect 5050 31732 5092 31772
rect 5132 31732 5174 31772
rect 5214 31732 5256 31772
rect 5296 31732 20048 31772
rect 20088 31732 20130 31772
rect 20170 31732 20212 31772
rect 20252 31732 20294 31772
rect 20334 31732 20376 31772
rect 20416 31732 20452 31772
rect 1152 31708 20452 31732
rect 6394 31604 6452 31605
rect 6394 31564 6403 31604
rect 6443 31564 6452 31604
rect 6394 31563 6452 31564
rect 9963 31604 10005 31613
rect 9963 31564 9964 31604
rect 10004 31564 10005 31604
rect 9963 31555 10005 31564
rect 11595 31604 11637 31613
rect 11595 31564 11596 31604
rect 11636 31564 11637 31604
rect 11595 31555 11637 31564
rect 18507 31604 18549 31613
rect 18507 31564 18508 31604
rect 18548 31564 18549 31604
rect 18507 31555 18549 31564
rect 20235 31604 20277 31613
rect 20235 31564 20236 31604
rect 20276 31564 20277 31604
rect 20235 31555 20277 31564
rect 3051 31520 3093 31529
rect 3051 31480 3052 31520
rect 3092 31480 3093 31520
rect 3051 31471 3093 31480
rect 4970 31520 5012 31529
rect 4970 31480 4971 31520
rect 5011 31480 5012 31520
rect 4970 31471 5012 31480
rect 5835 31520 5877 31529
rect 5835 31480 5836 31520
rect 5876 31480 5877 31520
rect 5835 31471 5877 31480
rect 13419 31520 13461 31529
rect 13419 31480 13420 31520
rect 13460 31480 13461 31520
rect 13419 31471 13461 31480
rect 14571 31520 14613 31529
rect 14571 31480 14572 31520
rect 14612 31480 14613 31520
rect 14571 31471 14613 31480
rect 15243 31520 15285 31529
rect 15243 31480 15244 31520
rect 15284 31480 15285 31520
rect 15243 31471 15285 31480
rect 16539 31520 16581 31529
rect 16539 31480 16540 31520
rect 16580 31480 16581 31520
rect 16539 31471 16581 31480
rect 1419 31436 1461 31445
rect 4491 31436 4533 31445
rect 1419 31396 1420 31436
rect 1460 31396 1461 31436
rect 1419 31387 1461 31396
rect 2667 31427 2709 31436
rect 2667 31387 2668 31427
rect 2708 31387 2709 31427
rect 2667 31378 2709 31387
rect 3243 31427 3285 31436
rect 3243 31387 3244 31427
rect 3284 31387 3285 31427
rect 4491 31396 4492 31436
rect 4532 31396 4533 31436
rect 4491 31387 4533 31396
rect 5092 31436 5150 31437
rect 5092 31396 5101 31436
rect 5141 31396 5150 31436
rect 5092 31395 5150 31396
rect 5355 31436 5397 31445
rect 5355 31396 5356 31436
rect 5396 31396 5397 31436
rect 5355 31387 5397 31396
rect 5632 31436 5674 31445
rect 5632 31396 5633 31436
rect 5673 31396 5674 31436
rect 6070 31436 6112 31445
rect 5632 31387 5674 31396
rect 5921 31403 5979 31404
rect 3243 31378 3285 31387
rect 5921 31363 5930 31403
rect 5970 31363 5979 31403
rect 6070 31396 6071 31436
rect 6111 31396 6112 31436
rect 6070 31387 6112 31396
rect 6315 31436 6357 31445
rect 6315 31396 6316 31436
rect 6356 31396 6357 31436
rect 6315 31387 6357 31396
rect 6795 31436 6837 31445
rect 8523 31436 8565 31445
rect 10155 31436 10197 31445
rect 11979 31436 12021 31445
rect 13899 31436 13941 31445
rect 6795 31396 6796 31436
rect 6836 31396 6837 31436
rect 6795 31387 6837 31396
rect 8043 31427 8085 31436
rect 8043 31387 8044 31427
rect 8084 31387 8085 31427
rect 8523 31396 8524 31436
rect 8564 31396 8565 31436
rect 8523 31387 8565 31396
rect 9771 31427 9813 31436
rect 9771 31387 9772 31427
rect 9812 31387 9813 31427
rect 10155 31396 10156 31436
rect 10196 31396 10197 31436
rect 10155 31387 10197 31396
rect 11403 31427 11445 31436
rect 11403 31387 11404 31427
rect 11444 31387 11445 31427
rect 11979 31396 11980 31436
rect 12020 31396 12021 31436
rect 11979 31387 12021 31396
rect 13227 31427 13269 31436
rect 13227 31387 13228 31427
rect 13268 31387 13269 31427
rect 13899 31396 13900 31436
rect 13940 31396 13941 31436
rect 13899 31387 13941 31396
rect 14187 31436 14229 31445
rect 14187 31396 14188 31436
rect 14228 31396 14229 31436
rect 14187 31387 14229 31396
rect 14458 31436 14516 31437
rect 14458 31396 14467 31436
rect 14507 31396 14516 31436
rect 14458 31395 14516 31396
rect 15037 31436 15079 31445
rect 17067 31436 17109 31445
rect 18795 31436 18837 31445
rect 15037 31396 15038 31436
rect 15078 31396 15079 31436
rect 15037 31387 15079 31396
rect 15339 31427 15381 31436
rect 15339 31387 15340 31427
rect 15380 31387 15381 31427
rect 17067 31396 17068 31436
rect 17108 31396 17109 31436
rect 17067 31387 17109 31396
rect 18315 31427 18357 31436
rect 18315 31387 18316 31427
rect 18356 31387 18357 31427
rect 18795 31396 18796 31436
rect 18836 31396 18837 31436
rect 18795 31387 18837 31396
rect 20043 31427 20085 31436
rect 20043 31387 20044 31427
rect 20084 31387 20085 31427
rect 8043 31378 8085 31387
rect 9771 31378 9813 31387
rect 11403 31378 11445 31387
rect 13227 31378 13269 31387
rect 15339 31378 15381 31387
rect 18315 31378 18357 31387
rect 20043 31378 20085 31387
rect 5921 31362 5979 31363
rect 6202 31352 6260 31353
rect 6202 31312 6211 31352
rect 6251 31312 6260 31352
rect 6202 31311 6260 31312
rect 15531 31352 15573 31361
rect 15531 31312 15532 31352
rect 15572 31312 15573 31352
rect 15531 31303 15573 31312
rect 15915 31352 15957 31361
rect 15915 31312 15916 31352
rect 15956 31312 15957 31352
rect 15915 31303 15957 31312
rect 16299 31352 16341 31361
rect 16299 31312 16300 31352
rect 16340 31312 16341 31352
rect 16299 31303 16341 31312
rect 16875 31352 16917 31361
rect 16875 31312 16876 31352
rect 16916 31312 16917 31352
rect 16875 31303 16917 31312
rect 2859 31184 2901 31193
rect 2859 31144 2860 31184
rect 2900 31144 2901 31184
rect 2859 31135 2901 31144
rect 4683 31184 4725 31193
rect 4683 31144 4684 31184
rect 4724 31144 4725 31184
rect 4683 31135 4725 31144
rect 5626 31184 5684 31185
rect 5626 31144 5635 31184
rect 5675 31144 5684 31184
rect 5626 31143 5684 31144
rect 8235 31184 8277 31193
rect 8235 31144 8236 31184
rect 8276 31144 8277 31184
rect 8235 31135 8277 31144
rect 13755 31184 13797 31193
rect 13755 31144 13756 31184
rect 13796 31144 13797 31184
rect 13755 31135 13797 31144
rect 14859 31184 14901 31193
rect 14859 31144 14860 31184
rect 14900 31144 14901 31184
rect 14859 31135 14901 31144
rect 15034 31184 15092 31185
rect 15034 31144 15043 31184
rect 15083 31144 15092 31184
rect 15034 31143 15092 31144
rect 15771 31184 15813 31193
rect 15771 31144 15772 31184
rect 15812 31144 15813 31184
rect 15771 31135 15813 31144
rect 16155 31184 16197 31193
rect 16155 31144 16156 31184
rect 16196 31144 16197 31184
rect 16155 31135 16197 31144
rect 16635 31184 16677 31193
rect 16635 31144 16636 31184
rect 16676 31144 16677 31184
rect 16635 31135 16677 31144
rect 1152 31016 20448 31040
rect 1152 30976 3688 31016
rect 3728 30976 3770 31016
rect 3810 30976 3852 31016
rect 3892 30976 3934 31016
rect 3974 30976 4016 31016
rect 4056 30976 18808 31016
rect 18848 30976 18890 31016
rect 18930 30976 18972 31016
rect 19012 30976 19054 31016
rect 19094 30976 19136 31016
rect 19176 30976 20448 31016
rect 1152 30952 20448 30976
rect 2667 30848 2709 30857
rect 2667 30808 2668 30848
rect 2708 30808 2709 30848
rect 2667 30799 2709 30808
rect 4474 30848 4532 30849
rect 4474 30808 4483 30848
rect 4523 30808 4532 30848
rect 4474 30807 4532 30808
rect 10779 30848 10821 30857
rect 10779 30808 10780 30848
rect 10820 30808 10821 30848
rect 10779 30799 10821 30808
rect 11163 30848 11205 30857
rect 11163 30808 11164 30848
rect 11204 30808 11205 30848
rect 11163 30799 11205 30808
rect 14571 30848 14613 30857
rect 14571 30808 14572 30848
rect 14612 30808 14613 30848
rect 14571 30799 14613 30808
rect 18843 30848 18885 30857
rect 18843 30808 18844 30848
rect 18884 30808 18885 30848
rect 18843 30799 18885 30808
rect 19995 30848 20037 30857
rect 19995 30808 19996 30848
rect 20036 30808 20037 30848
rect 19995 30799 20037 30808
rect 20379 30848 20421 30857
rect 20379 30808 20380 30848
rect 20420 30808 20421 30848
rect 20379 30799 20421 30808
rect 4299 30764 4341 30773
rect 4299 30724 4300 30764
rect 4340 30724 4341 30764
rect 4299 30715 4341 30724
rect 19611 30764 19653 30773
rect 19611 30724 19612 30764
rect 19652 30724 19653 30764
rect 19611 30715 19653 30724
rect 7467 30680 7509 30689
rect 7467 30640 7468 30680
rect 7508 30640 7509 30680
rect 7467 30631 7509 30640
rect 10539 30680 10581 30689
rect 10539 30640 10540 30680
rect 10580 30640 10581 30680
rect 10539 30631 10581 30640
rect 10923 30680 10965 30689
rect 16971 30680 17013 30689
rect 10923 30640 10924 30680
rect 10964 30640 10965 30680
rect 10923 30631 10965 30640
rect 13554 30671 13600 30680
rect 13554 30631 13555 30671
rect 13595 30631 13600 30671
rect 16971 30640 16972 30680
rect 17012 30640 17013 30680
rect 16971 30631 17013 30640
rect 18603 30680 18645 30689
rect 18603 30640 18604 30680
rect 18644 30640 18645 30680
rect 18603 30631 18645 30640
rect 18987 30680 19029 30689
rect 18987 30640 18988 30680
rect 19028 30640 19029 30680
rect 18987 30631 19029 30640
rect 19371 30680 19413 30689
rect 19371 30640 19372 30680
rect 19412 30640 19413 30680
rect 19371 30631 19413 30640
rect 19755 30680 19797 30689
rect 19755 30640 19756 30680
rect 19796 30640 19797 30680
rect 19755 30631 19797 30640
rect 20139 30680 20181 30689
rect 20139 30640 20140 30680
rect 20180 30640 20181 30680
rect 20139 30631 20181 30640
rect 13554 30622 13600 30631
rect 1227 30596 1269 30605
rect 1227 30556 1228 30596
rect 1268 30556 1269 30596
rect 1227 30547 1269 30556
rect 2467 30596 2525 30597
rect 2467 30556 2476 30596
rect 2516 30556 2525 30596
rect 2467 30555 2525 30556
rect 2859 30596 2901 30605
rect 2859 30556 2860 30596
rect 2900 30556 2901 30596
rect 2859 30547 2901 30556
rect 4099 30596 4157 30597
rect 4099 30556 4108 30596
rect 4148 30556 4157 30596
rect 4099 30555 4157 30556
rect 4771 30596 4829 30597
rect 4771 30556 4780 30596
rect 4820 30556 4829 30596
rect 4771 30555 4829 30556
rect 5067 30596 5109 30605
rect 5067 30556 5068 30596
rect 5108 30556 5109 30596
rect 5067 30547 5109 30556
rect 5259 30596 5301 30605
rect 5259 30556 5260 30596
rect 5300 30556 5301 30596
rect 5259 30547 5301 30556
rect 6499 30596 6557 30597
rect 6499 30556 6508 30596
rect 6548 30556 6557 30596
rect 6499 30555 6557 30556
rect 6970 30596 7028 30597
rect 6970 30556 6979 30596
rect 7019 30556 7028 30596
rect 6970 30555 7028 30556
rect 7083 30596 7125 30605
rect 7083 30556 7084 30596
rect 7124 30556 7125 30596
rect 7083 30547 7125 30556
rect 7563 30596 7605 30605
rect 7563 30556 7564 30596
rect 7604 30556 7605 30596
rect 7563 30547 7605 30556
rect 8035 30596 8093 30597
rect 8035 30556 8044 30596
rect 8084 30556 8093 30596
rect 8035 30555 8093 30556
rect 8554 30596 8612 30597
rect 8554 30556 8563 30596
rect 8603 30556 8612 30596
rect 8554 30555 8612 30556
rect 9091 30596 9149 30597
rect 9091 30556 9100 30596
rect 9140 30556 9149 30596
rect 9091 30555 9149 30556
rect 10347 30596 10389 30605
rect 10347 30556 10348 30596
rect 10388 30556 10389 30596
rect 10347 30547 10389 30556
rect 11307 30596 11349 30605
rect 11307 30556 11308 30596
rect 11348 30556 11349 30596
rect 11307 30547 11349 30556
rect 12547 30596 12605 30597
rect 12547 30556 12556 30596
rect 12596 30556 12605 30596
rect 12547 30555 12605 30556
rect 13035 30596 13077 30605
rect 13035 30556 13036 30596
rect 13076 30556 13077 30596
rect 13035 30547 13077 30556
rect 13323 30596 13365 30605
rect 13323 30556 13324 30596
rect 13364 30556 13365 30596
rect 13323 30547 13365 30556
rect 13428 30596 13470 30605
rect 13428 30556 13429 30596
rect 13469 30556 13470 30596
rect 13428 30547 13470 30556
rect 13648 30596 13706 30597
rect 13648 30556 13657 30596
rect 13697 30556 13706 30596
rect 13648 30555 13706 30556
rect 13899 30596 13941 30605
rect 13899 30556 13900 30596
rect 13940 30556 13941 30596
rect 13899 30547 13941 30556
rect 14170 30596 14228 30597
rect 14170 30556 14179 30596
rect 14219 30556 14228 30596
rect 14170 30555 14228 30556
rect 14763 30596 14805 30605
rect 14763 30556 14764 30596
rect 14804 30556 14805 30596
rect 14763 30547 14805 30556
rect 16003 30596 16061 30597
rect 16003 30556 16012 30596
rect 16052 30556 16061 30596
rect 16003 30555 16061 30556
rect 16474 30596 16532 30597
rect 16474 30556 16483 30596
rect 16523 30556 16532 30596
rect 16474 30555 16532 30556
rect 16587 30596 16629 30605
rect 16587 30556 16588 30596
rect 16628 30556 16629 30596
rect 16587 30547 16629 30556
rect 17067 30596 17109 30605
rect 17067 30556 17068 30596
rect 17108 30556 17109 30596
rect 17067 30547 17109 30556
rect 17539 30596 17597 30597
rect 17539 30556 17548 30596
rect 17588 30556 17597 30596
rect 17539 30555 17597 30556
rect 18027 30596 18085 30597
rect 18027 30556 18036 30596
rect 18076 30556 18085 30596
rect 18027 30555 18085 30556
rect 4477 30512 4519 30521
rect 4477 30472 4478 30512
rect 4518 30472 4519 30512
rect 4477 30463 4519 30472
rect 6699 30512 6741 30521
rect 6699 30472 6700 30512
rect 6740 30472 6741 30512
rect 6699 30463 6741 30472
rect 8907 30512 8949 30521
rect 8907 30472 8908 30512
rect 8948 30472 8949 30512
rect 8907 30463 8949 30472
rect 12747 30512 12789 30521
rect 12747 30472 12748 30512
rect 12788 30472 12789 30512
rect 12747 30463 12789 30472
rect 13179 30512 13221 30521
rect 13179 30472 13180 30512
rect 13220 30472 13221 30512
rect 13179 30463 13221 30472
rect 14283 30512 14325 30521
rect 14283 30472 14284 30512
rect 14324 30472 14325 30512
rect 14283 30463 14325 30472
rect 16203 30512 16245 30521
rect 16203 30472 16204 30512
rect 16244 30472 16245 30512
rect 16203 30463 16245 30472
rect 19227 30512 19269 30521
rect 19227 30472 19228 30512
rect 19268 30472 19269 30512
rect 19227 30463 19269 30472
rect 4683 30428 4725 30437
rect 4683 30388 4684 30428
rect 4724 30388 4725 30428
rect 4683 30379 4725 30388
rect 4923 30428 4965 30437
rect 4923 30388 4924 30428
rect 4964 30388 4965 30428
rect 4923 30379 4965 30388
rect 8715 30428 8757 30437
rect 8715 30388 8716 30428
rect 8756 30388 8757 30428
rect 8715 30379 8757 30388
rect 18219 30428 18261 30437
rect 18219 30388 18220 30428
rect 18260 30388 18261 30428
rect 18219 30379 18261 30388
rect 1152 30260 20452 30284
rect 1152 30220 4928 30260
rect 4968 30220 5010 30260
rect 5050 30220 5092 30260
rect 5132 30220 5174 30260
rect 5214 30220 5256 30260
rect 5296 30220 20048 30260
rect 20088 30220 20130 30260
rect 20170 30220 20212 30260
rect 20252 30220 20294 30260
rect 20334 30220 20376 30260
rect 20416 30220 20452 30260
rect 1152 30196 20452 30220
rect 2859 30092 2901 30101
rect 2859 30052 2860 30092
rect 2900 30052 2901 30092
rect 2859 30043 2901 30052
rect 3051 30092 3093 30101
rect 3051 30052 3052 30092
rect 3092 30052 3093 30092
rect 3051 30043 3093 30052
rect 13978 30092 14036 30093
rect 13978 30052 13987 30092
rect 14027 30052 14036 30092
rect 13978 30051 14036 30052
rect 14458 30092 14516 30093
rect 14458 30052 14467 30092
rect 14507 30052 14516 30092
rect 14458 30051 14516 30052
rect 14938 30092 14996 30093
rect 14938 30052 14947 30092
rect 14987 30052 14996 30092
rect 14938 30051 14996 30052
rect 15339 30092 15381 30101
rect 15339 30052 15340 30092
rect 15380 30052 15381 30092
rect 15339 30043 15381 30052
rect 18891 30092 18933 30101
rect 18891 30052 18892 30092
rect 18932 30052 18933 30092
rect 18891 30043 18933 30052
rect 19995 30092 20037 30101
rect 19995 30052 19996 30092
rect 20036 30052 20037 30092
rect 19995 30043 20037 30052
rect 20379 30092 20421 30101
rect 20379 30052 20380 30092
rect 20420 30052 20421 30092
rect 20379 30043 20421 30052
rect 6411 30008 6453 30017
rect 6411 29968 6412 30008
rect 6452 29968 6453 30008
rect 6411 29959 6453 29968
rect 8859 30008 8901 30017
rect 8859 29968 8860 30008
rect 8900 29968 8901 30008
rect 8859 29959 8901 29968
rect 19179 30008 19221 30017
rect 19179 29968 19180 30008
rect 19220 29968 19221 30008
rect 19179 29959 19221 29968
rect 1419 29924 1461 29933
rect 4491 29924 4533 29933
rect 1419 29884 1420 29924
rect 1460 29884 1461 29924
rect 1419 29875 1461 29884
rect 2667 29915 2709 29924
rect 2667 29875 2668 29915
rect 2708 29875 2709 29915
rect 2667 29866 2709 29875
rect 3243 29915 3285 29924
rect 3243 29875 3244 29915
rect 3284 29875 3285 29915
rect 4491 29884 4492 29924
rect 4532 29884 4533 29924
rect 4491 29875 4533 29884
rect 4779 29924 4821 29933
rect 4779 29884 4780 29924
rect 4820 29884 4821 29924
rect 4779 29875 4821 29884
rect 4971 29924 5013 29933
rect 6682 29924 6740 29925
rect 4971 29884 4972 29924
rect 5012 29884 5013 29924
rect 4971 29875 5013 29884
rect 6219 29915 6261 29924
rect 6219 29875 6220 29915
rect 6260 29875 6261 29915
rect 6682 29884 6691 29924
rect 6731 29884 6740 29924
rect 6682 29883 6740 29884
rect 6795 29924 6837 29933
rect 6795 29884 6796 29924
rect 6836 29884 6837 29924
rect 6795 29875 6837 29884
rect 7179 29924 7221 29933
rect 9003 29924 9045 29933
rect 7179 29884 7180 29924
rect 7220 29884 7221 29924
rect 7179 29875 7221 29884
rect 7755 29915 7797 29924
rect 7755 29875 7756 29915
rect 7796 29875 7797 29915
rect 3243 29866 3285 29875
rect 6219 29866 6261 29875
rect 7755 29866 7797 29875
rect 8235 29915 8277 29924
rect 8235 29875 8236 29915
rect 8276 29875 8277 29915
rect 9003 29884 9004 29924
rect 9044 29884 9045 29924
rect 9003 29875 9045 29884
rect 9195 29924 9237 29933
rect 9195 29884 9196 29924
rect 9236 29884 9237 29924
rect 9195 29875 9237 29884
rect 9658 29924 9716 29925
rect 9658 29884 9667 29924
rect 9707 29884 9716 29924
rect 9658 29883 9716 29884
rect 9771 29924 9813 29933
rect 9771 29884 9772 29924
rect 9812 29884 9813 29924
rect 9771 29875 9813 29884
rect 10155 29924 10197 29933
rect 13035 29924 13077 29933
rect 10155 29884 10156 29924
rect 10196 29884 10197 29924
rect 10155 29875 10197 29884
rect 10731 29915 10773 29924
rect 10731 29875 10732 29915
rect 10772 29875 10773 29915
rect 8235 29866 8277 29875
rect 10731 29866 10773 29875
rect 11211 29915 11253 29924
rect 11211 29875 11212 29915
rect 11252 29875 11253 29915
rect 13035 29884 13036 29924
rect 13076 29884 13077 29924
rect 13035 29875 13077 29884
rect 13323 29924 13365 29933
rect 13323 29884 13324 29924
rect 13364 29884 13365 29924
rect 13323 29875 13365 29884
rect 13498 29924 13556 29925
rect 13498 29884 13507 29924
rect 13547 29884 13556 29924
rect 13498 29883 13556 29884
rect 13654 29924 13696 29933
rect 13654 29884 13655 29924
rect 13695 29884 13696 29924
rect 13654 29875 13696 29884
rect 13897 29924 13939 29933
rect 13897 29884 13898 29924
rect 13938 29884 13939 29924
rect 13897 29875 13939 29884
rect 14146 29924 14204 29925
rect 14146 29884 14155 29924
rect 14195 29884 14204 29924
rect 14146 29883 14204 29884
rect 14360 29924 14402 29933
rect 14360 29884 14361 29924
rect 14401 29884 14402 29924
rect 14360 29875 14402 29884
rect 14619 29924 14661 29933
rect 14619 29884 14620 29924
rect 14660 29884 14661 29924
rect 14619 29875 14661 29884
rect 14746 29924 14804 29925
rect 14746 29884 14755 29924
rect 14795 29884 14804 29924
rect 14746 29883 14804 29884
rect 14859 29924 14901 29933
rect 14859 29884 14860 29924
rect 14900 29884 14901 29924
rect 14859 29875 14901 29884
rect 15133 29924 15175 29933
rect 16378 29924 16436 29925
rect 15133 29884 15134 29924
rect 15174 29884 15175 29924
rect 15133 29875 15175 29884
rect 15435 29915 15477 29924
rect 15435 29875 15436 29915
rect 15476 29875 15477 29915
rect 16378 29884 16387 29924
rect 16427 29884 16436 29924
rect 16378 29883 16436 29884
rect 16683 29924 16725 29933
rect 16683 29884 16684 29924
rect 16724 29884 16725 29924
rect 16683 29875 16725 29884
rect 17146 29924 17204 29925
rect 17146 29884 17155 29924
rect 17195 29884 17204 29924
rect 17146 29883 17204 29884
rect 17259 29924 17301 29933
rect 17259 29884 17260 29924
rect 17300 29884 17301 29924
rect 17259 29875 17301 29884
rect 17643 29924 17685 29933
rect 19066 29924 19124 29925
rect 17643 29884 17644 29924
rect 17684 29884 17685 29924
rect 17643 29875 17685 29884
rect 18219 29915 18261 29924
rect 18219 29875 18220 29915
rect 18260 29875 18261 29915
rect 11211 29866 11253 29875
rect 15435 29866 15477 29875
rect 18219 29866 18261 29875
rect 18699 29915 18741 29924
rect 18699 29875 18700 29915
rect 18740 29875 18741 29915
rect 19066 29884 19075 29924
rect 19115 29884 19124 29924
rect 19066 29883 19124 29884
rect 19385 29924 19427 29933
rect 19385 29884 19386 29924
rect 19426 29884 19427 29924
rect 19385 29875 19427 29884
rect 18699 29866 18741 29875
rect 7275 29840 7317 29849
rect 7275 29800 7276 29840
rect 7316 29800 7317 29840
rect 7275 29791 7317 29800
rect 8619 29840 8661 29849
rect 8619 29800 8620 29840
rect 8660 29800 8661 29840
rect 8619 29791 8661 29800
rect 10251 29840 10293 29849
rect 10251 29800 10252 29840
rect 10292 29800 10293 29840
rect 10251 29791 10293 29800
rect 11434 29840 11492 29841
rect 11434 29800 11443 29840
rect 11483 29800 11492 29840
rect 11434 29799 11492 29800
rect 11787 29840 11829 29849
rect 11787 29800 11788 29840
rect 11828 29800 11829 29840
rect 11787 29791 11829 29800
rect 12267 29840 12309 29849
rect 12267 29800 12268 29840
rect 12308 29800 12309 29840
rect 12267 29791 12309 29800
rect 13786 29840 13844 29841
rect 13786 29800 13795 29840
rect 13835 29800 13844 29840
rect 13786 29799 13844 29800
rect 14266 29840 14324 29841
rect 14266 29800 14275 29840
rect 14315 29800 14324 29840
rect 14266 29799 14324 29800
rect 15819 29840 15861 29849
rect 15819 29800 15820 29840
rect 15860 29800 15861 29840
rect 15819 29791 15861 29800
rect 16203 29840 16245 29849
rect 16203 29800 16204 29840
rect 16244 29800 16245 29840
rect 16203 29791 16245 29800
rect 17739 29840 17781 29849
rect 17739 29800 17740 29840
rect 17780 29800 17781 29840
rect 17739 29791 17781 29800
rect 19755 29840 19797 29849
rect 19755 29800 19756 29840
rect 19796 29800 19797 29840
rect 19755 29791 19797 29800
rect 20139 29840 20181 29849
rect 20139 29800 20140 29840
rect 20180 29800 20181 29840
rect 20139 29791 20181 29800
rect 8475 29756 8517 29765
rect 8475 29716 8476 29756
rect 8516 29716 8517 29756
rect 8475 29707 8517 29716
rect 2859 29672 2901 29681
rect 2859 29632 2860 29672
rect 2900 29632 2901 29672
rect 2859 29623 2901 29632
rect 4635 29672 4677 29681
rect 4635 29632 4636 29672
rect 4676 29632 4677 29672
rect 4635 29623 4677 29632
rect 9003 29672 9045 29681
rect 9003 29632 9004 29672
rect 9044 29632 9045 29672
rect 9003 29623 9045 29632
rect 11547 29672 11589 29681
rect 11547 29632 11548 29672
rect 11588 29632 11589 29672
rect 11547 29623 11589 29632
rect 12507 29672 12549 29681
rect 12507 29632 12508 29672
rect 12548 29632 12549 29672
rect 12507 29623 12549 29632
rect 13179 29672 13221 29681
rect 13179 29632 13180 29672
rect 13220 29632 13221 29672
rect 13179 29623 13221 29632
rect 13498 29672 13556 29673
rect 13498 29632 13507 29672
rect 13547 29632 13556 29672
rect 13498 29631 13556 29632
rect 15130 29672 15188 29673
rect 15130 29632 15139 29672
rect 15179 29632 15188 29672
rect 15130 29631 15188 29632
rect 15579 29672 15621 29681
rect 15579 29632 15580 29672
rect 15620 29632 15621 29672
rect 15579 29623 15621 29632
rect 15963 29672 16005 29681
rect 15963 29632 15964 29672
rect 16004 29632 16005 29672
rect 15963 29623 16005 29632
rect 16683 29672 16725 29681
rect 16683 29632 16684 29672
rect 16724 29632 16725 29672
rect 16683 29623 16725 29632
rect 19371 29672 19413 29681
rect 19371 29632 19372 29672
rect 19412 29632 19413 29672
rect 19371 29623 19413 29632
rect 1152 29504 20448 29528
rect 1152 29464 3688 29504
rect 3728 29464 3770 29504
rect 3810 29464 3852 29504
rect 3892 29464 3934 29504
rect 3974 29464 4016 29504
rect 4056 29464 18808 29504
rect 18848 29464 18890 29504
rect 18930 29464 18972 29504
rect 19012 29464 19054 29504
rect 19094 29464 19136 29504
rect 19176 29464 20448 29504
rect 1152 29440 20448 29464
rect 1467 29336 1509 29345
rect 1467 29296 1468 29336
rect 1508 29296 1509 29336
rect 1467 29287 1509 29296
rect 2235 29336 2277 29345
rect 2235 29296 2236 29336
rect 2276 29296 2277 29336
rect 2235 29287 2277 29296
rect 4443 29336 4485 29345
rect 4443 29296 4444 29336
rect 4484 29296 4485 29336
rect 4443 29287 4485 29296
rect 6315 29336 6357 29345
rect 6315 29296 6316 29336
rect 6356 29296 6357 29336
rect 6315 29287 6357 29296
rect 13515 29336 13557 29345
rect 13515 29296 13516 29336
rect 13556 29296 13557 29336
rect 13515 29287 13557 29296
rect 14475 29336 14517 29345
rect 14475 29296 14476 29336
rect 14516 29296 14517 29336
rect 14475 29287 14517 29296
rect 15195 29336 15237 29345
rect 15195 29296 15196 29336
rect 15236 29296 15237 29336
rect 15195 29287 15237 29296
rect 17739 29336 17781 29345
rect 17739 29296 17740 29336
rect 17780 29296 17781 29336
rect 17739 29287 17781 29296
rect 19851 29336 19893 29345
rect 19851 29296 19852 29336
rect 19892 29296 19893 29336
rect 19851 29287 19893 29296
rect 20379 29336 20421 29345
rect 20379 29296 20380 29336
rect 20420 29296 20421 29336
rect 20379 29287 20421 29296
rect 9243 29252 9285 29261
rect 9243 29212 9244 29252
rect 9284 29212 9285 29252
rect 9243 29203 9285 29212
rect 1227 29168 1269 29177
rect 1227 29128 1228 29168
rect 1268 29128 1269 29168
rect 1227 29119 1269 29128
rect 1611 29168 1653 29177
rect 1611 29128 1612 29168
rect 1652 29128 1653 29168
rect 1611 29119 1653 29128
rect 1995 29168 2037 29177
rect 1995 29128 1996 29168
rect 2036 29128 2037 29168
rect 1995 29119 2037 29128
rect 2786 29168 2828 29177
rect 4683 29168 4725 29177
rect 2786 29128 2787 29168
rect 2827 29128 2828 29168
rect 2786 29119 2828 29128
rect 3282 29159 3328 29168
rect 3282 29119 3283 29159
rect 3323 29119 3328 29159
rect 3282 29110 3328 29119
rect 3387 29126 3429 29135
rect 2667 29084 2709 29093
rect 2667 29044 2668 29084
rect 2708 29044 2709 29084
rect 2667 29035 2709 29044
rect 2884 29084 2926 29093
rect 2884 29044 2885 29084
rect 2925 29044 2926 29084
rect 2884 29035 2926 29044
rect 3156 29084 3198 29093
rect 3156 29044 3157 29084
rect 3197 29044 3198 29084
rect 3387 29086 3388 29126
rect 3428 29086 3429 29126
rect 4683 29128 4684 29168
rect 4724 29128 4725 29168
rect 4683 29119 4725 29128
rect 7275 29168 7317 29177
rect 7275 29128 7276 29168
rect 7316 29128 7317 29168
rect 7275 29119 7317 29128
rect 9003 29168 9045 29177
rect 9003 29128 9004 29168
rect 9044 29128 9045 29168
rect 9003 29119 9045 29128
rect 9387 29168 9429 29177
rect 9387 29128 9388 29168
rect 9428 29128 9429 29168
rect 9387 29119 9429 29128
rect 10347 29168 10389 29177
rect 10347 29128 10348 29168
rect 10388 29128 10389 29168
rect 10347 29119 10389 29128
rect 14667 29168 14709 29177
rect 14667 29128 14668 29168
rect 14708 29128 14709 29168
rect 14667 29119 14709 29128
rect 15435 29168 15477 29177
rect 15435 29128 15436 29168
rect 15476 29128 15477 29168
rect 15435 29119 15477 29128
rect 20139 29168 20181 29177
rect 20139 29128 20140 29168
rect 20180 29128 20181 29168
rect 15723 29117 15765 29126
rect 20139 29119 20181 29128
rect 3387 29077 3429 29086
rect 3627 29084 3669 29093
rect 3156 29035 3198 29044
rect 3627 29044 3628 29084
rect 3668 29044 3669 29084
rect 3627 29035 3669 29044
rect 3898 29084 3956 29085
rect 3898 29044 3907 29084
rect 3947 29044 3956 29084
rect 3898 29043 3956 29044
rect 4875 29084 4917 29093
rect 4875 29044 4876 29084
rect 4916 29044 4917 29084
rect 4875 29035 4917 29044
rect 6115 29084 6173 29085
rect 6115 29044 6124 29084
rect 6164 29044 6173 29084
rect 6115 29043 6173 29044
rect 6778 29084 6836 29085
rect 6778 29044 6787 29084
rect 6827 29044 6836 29084
rect 6778 29043 6836 29044
rect 6891 29084 6933 29093
rect 6891 29044 6892 29084
rect 6932 29044 6933 29084
rect 6891 29035 6933 29044
rect 7371 29084 7413 29093
rect 7371 29044 7372 29084
rect 7412 29044 7413 29084
rect 7371 29035 7413 29044
rect 7843 29084 7901 29085
rect 7843 29044 7852 29084
rect 7892 29044 7901 29084
rect 7843 29043 7901 29044
rect 8362 29084 8420 29085
rect 8362 29044 8371 29084
rect 8411 29044 8420 29084
rect 8362 29043 8420 29044
rect 9850 29084 9908 29085
rect 9850 29044 9859 29084
rect 9899 29044 9908 29084
rect 9850 29043 9908 29044
rect 9963 29084 10005 29093
rect 9963 29044 9964 29084
rect 10004 29044 10005 29084
rect 9963 29035 10005 29044
rect 10443 29084 10485 29093
rect 10443 29044 10444 29084
rect 10484 29044 10485 29084
rect 10443 29035 10485 29044
rect 10915 29084 10973 29085
rect 10915 29044 10924 29084
rect 10964 29044 10973 29084
rect 10915 29043 10973 29044
rect 11403 29084 11461 29085
rect 11403 29044 11412 29084
rect 11452 29044 11461 29084
rect 11403 29043 11461 29044
rect 12075 29084 12117 29093
rect 12075 29044 12076 29084
rect 12116 29044 12117 29084
rect 12075 29035 12117 29044
rect 13315 29084 13373 29085
rect 13315 29044 13324 29084
rect 13364 29044 13373 29084
rect 13315 29043 13373 29044
rect 14170 29084 14228 29085
rect 14170 29044 14179 29084
rect 14219 29044 14228 29084
rect 15723 29077 15724 29117
rect 15764 29077 15765 29117
rect 15723 29068 15765 29077
rect 15826 29084 15884 29085
rect 14170 29043 14228 29044
rect 15826 29044 15835 29084
rect 15875 29044 15884 29084
rect 15826 29043 15884 29044
rect 15944 29084 16002 29085
rect 15944 29044 15953 29084
rect 15993 29044 16002 29084
rect 15944 29043 16002 29044
rect 16299 29084 16341 29093
rect 16299 29044 16300 29084
rect 16340 29044 16341 29084
rect 16299 29035 16341 29044
rect 17539 29084 17597 29085
rect 17539 29044 17548 29084
rect 17588 29044 17597 29084
rect 17539 29043 17597 29044
rect 17917 29084 17959 29093
rect 17917 29044 17918 29084
rect 17958 29044 17959 29084
rect 17917 29035 17959 29044
rect 18123 29084 18165 29093
rect 18123 29044 18124 29084
rect 18164 29044 18165 29084
rect 18123 29035 18165 29044
rect 18211 29084 18269 29085
rect 18211 29044 18220 29084
rect 18260 29044 18269 29084
rect 18211 29043 18269 29044
rect 18411 29084 18453 29093
rect 18411 29044 18412 29084
rect 18452 29044 18453 29084
rect 18411 29035 18453 29044
rect 19651 29084 19709 29085
rect 19651 29044 19660 29084
rect 19700 29044 19709 29084
rect 19651 29043 19709 29044
rect 4011 29000 4053 29009
rect 4011 28960 4012 29000
rect 4052 28960 4053 29000
rect 4011 28951 4053 28960
rect 4347 29000 4389 29009
rect 4347 28960 4348 29000
rect 4388 28960 4389 29000
rect 4347 28951 4389 28960
rect 14283 29000 14325 29009
rect 14283 28960 14284 29000
rect 14324 28960 14325 29000
rect 14283 28951 14325 28960
rect 14489 29000 14531 29009
rect 14489 28960 14490 29000
rect 14530 28960 14531 29000
rect 14489 28951 14531 28960
rect 1851 28916 1893 28925
rect 1851 28876 1852 28916
rect 1892 28876 1893 28916
rect 1851 28867 1893 28876
rect 2571 28916 2613 28925
rect 2571 28876 2572 28916
rect 2612 28876 2613 28916
rect 2571 28867 2613 28876
rect 3051 28916 3093 28925
rect 3051 28876 3052 28916
rect 3092 28876 3093 28916
rect 3051 28867 3093 28876
rect 8523 28916 8565 28925
rect 8523 28876 8524 28916
rect 8564 28876 8565 28916
rect 8523 28867 8565 28876
rect 9627 28916 9669 28925
rect 9627 28876 9628 28916
rect 9668 28876 9669 28916
rect 9627 28867 9669 28876
rect 11595 28916 11637 28925
rect 11595 28876 11596 28916
rect 11636 28876 11637 28916
rect 11595 28867 11637 28876
rect 14907 28916 14949 28925
rect 14907 28876 14908 28916
rect 14948 28876 14949 28916
rect 14907 28867 14949 28876
rect 16107 28916 16149 28925
rect 16107 28876 16108 28916
rect 16148 28876 16149 28916
rect 16107 28867 16149 28876
rect 18010 28916 18068 28917
rect 18010 28876 18019 28916
rect 18059 28876 18068 28916
rect 18010 28875 18068 28876
rect 1152 28748 20452 28772
rect 1152 28708 4928 28748
rect 4968 28708 5010 28748
rect 5050 28708 5092 28748
rect 5132 28708 5174 28748
rect 5214 28708 5256 28748
rect 5296 28708 20048 28748
rect 20088 28708 20130 28748
rect 20170 28708 20212 28748
rect 20252 28708 20294 28748
rect 20334 28708 20376 28748
rect 20416 28708 20452 28748
rect 1152 28684 20452 28708
rect 3610 28580 3668 28581
rect 3610 28540 3619 28580
rect 3659 28540 3668 28580
rect 3610 28539 3668 28540
rect 4203 28580 4245 28589
rect 4203 28540 4204 28580
rect 4244 28540 4245 28580
rect 4203 28531 4245 28540
rect 5211 28580 5253 28589
rect 5211 28540 5212 28580
rect 5252 28540 5253 28580
rect 5211 28531 5253 28540
rect 6795 28580 6837 28589
rect 6795 28540 6796 28580
rect 6836 28540 6837 28580
rect 6795 28531 6837 28540
rect 8811 28580 8853 28589
rect 8811 28540 8812 28580
rect 8852 28540 8853 28580
rect 8811 28531 8853 28540
rect 9243 28580 9285 28589
rect 9243 28540 9244 28580
rect 9284 28540 9285 28580
rect 9243 28531 9285 28540
rect 9627 28580 9669 28589
rect 9627 28540 9628 28580
rect 9668 28540 9669 28580
rect 9627 28531 9669 28540
rect 10395 28580 10437 28589
rect 10395 28540 10396 28580
rect 10436 28540 10437 28580
rect 10395 28531 10437 28540
rect 10539 28580 10581 28589
rect 10539 28540 10540 28580
rect 10580 28540 10581 28580
rect 10539 28531 10581 28540
rect 13995 28580 14037 28589
rect 13995 28540 13996 28580
rect 14036 28540 14037 28580
rect 13995 28531 14037 28540
rect 15819 28580 15861 28589
rect 15819 28540 15820 28580
rect 15860 28540 15861 28580
rect 15819 28531 15861 28540
rect 17451 28580 17493 28589
rect 17451 28540 17452 28580
rect 17492 28540 17493 28580
rect 17451 28531 17493 28540
rect 19083 28580 19125 28589
rect 19083 28540 19084 28580
rect 19124 28540 19125 28580
rect 19083 28531 19125 28540
rect 20026 28580 20084 28581
rect 20026 28540 20035 28580
rect 20075 28540 20084 28580
rect 20026 28539 20084 28540
rect 3997 28496 4039 28505
rect 3997 28456 3998 28496
rect 4038 28456 4039 28496
rect 3997 28447 4039 28456
rect 1515 28412 1557 28421
rect 3286 28412 3328 28421
rect 1515 28372 1516 28412
rect 1556 28372 1557 28412
rect 1515 28363 1557 28372
rect 2763 28403 2805 28412
rect 2763 28363 2764 28403
rect 2804 28363 2805 28403
rect 3286 28372 3287 28412
rect 3327 28372 3328 28412
rect 3286 28363 3328 28372
rect 3531 28412 3573 28421
rect 4587 28412 4629 28421
rect 3531 28372 3532 28412
rect 3572 28372 3573 28412
rect 3531 28363 3573 28372
rect 4299 28403 4341 28412
rect 4299 28363 4300 28403
rect 4340 28363 4341 28403
rect 4587 28372 4588 28412
rect 4628 28372 4629 28412
rect 4587 28363 4629 28372
rect 4804 28412 4846 28421
rect 4804 28372 4805 28412
rect 4845 28372 4846 28412
rect 4804 28363 4846 28372
rect 5355 28412 5397 28421
rect 7066 28412 7124 28413
rect 5355 28372 5356 28412
rect 5396 28372 5397 28412
rect 5355 28363 5397 28372
rect 6603 28403 6645 28412
rect 6603 28363 6604 28403
rect 6644 28363 6645 28403
rect 7066 28372 7075 28412
rect 7115 28372 7124 28412
rect 7066 28371 7124 28372
rect 7179 28412 7221 28421
rect 7179 28372 7180 28412
rect 7220 28372 7221 28412
rect 7179 28363 7221 28372
rect 7563 28412 7605 28421
rect 11979 28412 12021 28421
rect 7563 28372 7564 28412
rect 7604 28372 7605 28412
rect 7563 28363 7605 28372
rect 8139 28403 8181 28412
rect 8139 28363 8140 28403
rect 8180 28363 8181 28403
rect 2763 28354 2805 28363
rect 4299 28354 4341 28363
rect 6603 28354 6645 28363
rect 8139 28354 8181 28363
rect 8619 28403 8661 28412
rect 8619 28363 8620 28403
rect 8660 28363 8661 28403
rect 8619 28354 8661 28363
rect 10731 28403 10773 28412
rect 10731 28363 10732 28403
rect 10772 28363 10773 28403
rect 11979 28372 11980 28412
rect 12020 28372 12021 28412
rect 11979 28363 12021 28372
rect 12555 28412 12597 28421
rect 14379 28412 14421 28421
rect 16011 28412 16053 28421
rect 17643 28412 17685 28421
rect 19947 28412 19989 28421
rect 12555 28372 12556 28412
rect 12596 28372 12597 28412
rect 12555 28363 12597 28372
rect 13803 28403 13845 28412
rect 13803 28363 13804 28403
rect 13844 28363 13845 28403
rect 14379 28372 14380 28412
rect 14420 28372 14421 28412
rect 14379 28363 14421 28372
rect 15627 28403 15669 28412
rect 15627 28363 15628 28403
rect 15668 28363 15669 28403
rect 16011 28372 16012 28412
rect 16052 28372 16053 28412
rect 16011 28363 16053 28372
rect 17259 28403 17301 28412
rect 17259 28363 17260 28403
rect 17300 28363 17301 28403
rect 17643 28372 17644 28412
rect 17684 28372 17685 28412
rect 17643 28363 17685 28372
rect 18891 28403 18933 28412
rect 18891 28363 18892 28403
rect 18932 28363 18933 28403
rect 10731 28354 10773 28363
rect 13803 28354 13845 28363
rect 15627 28354 15669 28363
rect 17259 28354 17301 28363
rect 18891 28354 18933 28363
rect 19371 28403 19413 28412
rect 19371 28363 19372 28403
rect 19412 28363 19413 28403
rect 19371 28354 19413 28363
rect 19470 28392 19512 28401
rect 19470 28352 19471 28392
rect 19511 28352 19512 28392
rect 19947 28372 19948 28412
rect 19988 28372 19989 28412
rect 19470 28343 19512 28352
rect 19592 28370 19650 28371
rect 3418 28328 3476 28329
rect 3418 28288 3427 28328
rect 3467 28288 3476 28328
rect 3418 28287 3476 28288
rect 4491 28328 4533 28337
rect 4491 28288 4492 28328
rect 4532 28288 4533 28328
rect 4491 28279 4533 28288
rect 4706 28328 4748 28337
rect 4706 28288 4707 28328
rect 4747 28288 4748 28328
rect 4706 28279 4748 28288
rect 4971 28328 5013 28337
rect 4971 28288 4972 28328
rect 5012 28288 5013 28328
rect 4971 28279 5013 28288
rect 7659 28328 7701 28337
rect 7659 28288 7660 28328
rect 7700 28288 7701 28328
rect 7659 28279 7701 28288
rect 9003 28328 9045 28337
rect 9003 28288 9004 28328
rect 9044 28288 9045 28328
rect 9003 28279 9045 28288
rect 9387 28328 9429 28337
rect 9387 28288 9388 28328
rect 9428 28288 9429 28328
rect 9387 28279 9429 28288
rect 9771 28328 9813 28337
rect 9771 28288 9772 28328
rect 9812 28288 9813 28328
rect 9771 28279 9813 28288
rect 10155 28328 10197 28337
rect 10155 28288 10156 28328
rect 10196 28288 10197 28328
rect 10155 28279 10197 28288
rect 12363 28328 12405 28337
rect 19592 28330 19601 28370
rect 19641 28330 19650 28370
rect 19947 28363 19989 28372
rect 20235 28412 20277 28421
rect 20235 28372 20236 28412
rect 20276 28372 20277 28412
rect 20235 28363 20277 28372
rect 19592 28329 19650 28330
rect 12363 28288 12364 28328
rect 12404 28288 12405 28328
rect 12363 28279 12405 28288
rect 2955 28244 2997 28253
rect 2955 28204 2956 28244
rect 2996 28204 2997 28244
rect 2955 28195 2997 28204
rect 10011 28244 10053 28253
rect 10011 28204 10012 28244
rect 10052 28204 10053 28244
rect 10011 28195 10053 28204
rect 3994 28160 4052 28161
rect 3994 28120 4003 28160
rect 4043 28120 4052 28160
rect 3994 28119 4052 28120
rect 12123 28160 12165 28169
rect 12123 28120 12124 28160
rect 12164 28120 12165 28160
rect 12123 28111 12165 28120
rect 19755 28160 19797 28169
rect 19755 28120 19756 28160
rect 19796 28120 19797 28160
rect 19755 28111 19797 28120
rect 1152 27992 20448 28016
rect 1152 27952 3688 27992
rect 3728 27952 3770 27992
rect 3810 27952 3852 27992
rect 3892 27952 3934 27992
rect 3974 27952 4016 27992
rect 4056 27952 18808 27992
rect 18848 27952 18890 27992
rect 18930 27952 18972 27992
rect 19012 27952 19054 27992
rect 19094 27952 19136 27992
rect 19176 27952 20448 27992
rect 1152 27928 20448 27952
rect 1467 27824 1509 27833
rect 1467 27784 1468 27824
rect 1508 27784 1509 27824
rect 1467 27775 1509 27784
rect 3051 27824 3093 27833
rect 3051 27784 3052 27824
rect 3092 27784 3093 27824
rect 3051 27775 3093 27784
rect 7563 27824 7605 27833
rect 7563 27784 7564 27824
rect 7604 27784 7605 27824
rect 7563 27775 7605 27784
rect 11019 27824 11061 27833
rect 11019 27784 11020 27824
rect 11060 27784 11061 27824
rect 11019 27775 11061 27784
rect 14571 27824 14613 27833
rect 14571 27784 14572 27824
rect 14612 27784 14613 27824
rect 14571 27775 14613 27784
rect 16491 27824 16533 27833
rect 16491 27784 16492 27824
rect 16532 27784 16533 27824
rect 16491 27775 16533 27784
rect 19851 27824 19893 27833
rect 19851 27784 19852 27824
rect 19892 27784 19893 27824
rect 19851 27775 19893 27784
rect 4299 27740 4341 27749
rect 4299 27700 4300 27740
rect 4340 27700 4341 27740
rect 4299 27691 4341 27700
rect 11211 27740 11253 27749
rect 11211 27700 11212 27740
rect 11252 27700 11253 27740
rect 11211 27691 11253 27700
rect 1227 27656 1269 27665
rect 1227 27616 1228 27656
rect 1268 27616 1269 27656
rect 1227 27607 1269 27616
rect 5050 27656 5108 27657
rect 5050 27616 5059 27656
rect 5099 27616 5108 27656
rect 5050 27615 5108 27616
rect 5259 27656 5301 27665
rect 5259 27616 5260 27656
rect 5300 27616 5301 27656
rect 5259 27607 5301 27616
rect 5530 27656 5588 27657
rect 5530 27616 5539 27656
rect 5579 27616 5588 27656
rect 5530 27615 5588 27616
rect 5739 27656 5781 27665
rect 5739 27616 5740 27656
rect 5780 27616 5781 27656
rect 5739 27607 5781 27616
rect 1611 27572 1653 27581
rect 1611 27532 1612 27572
rect 1652 27532 1653 27572
rect 1611 27523 1653 27532
rect 2851 27572 2909 27573
rect 2851 27532 2860 27572
rect 2900 27532 2909 27572
rect 2851 27531 2909 27532
rect 3243 27572 3285 27581
rect 3243 27532 3244 27572
rect 3284 27532 3285 27572
rect 3243 27523 3285 27532
rect 3627 27572 3669 27581
rect 3627 27532 3628 27572
rect 3668 27532 3669 27572
rect 3627 27523 3669 27532
rect 3898 27572 3956 27573
rect 3898 27532 3907 27572
rect 3947 27532 3956 27572
rect 3898 27531 3956 27532
rect 4474 27572 4532 27573
rect 4474 27532 4483 27572
rect 4523 27532 4532 27572
rect 4474 27531 4532 27532
rect 4918 27572 4960 27581
rect 4918 27532 4919 27572
rect 4959 27532 4960 27572
rect 4918 27523 4960 27532
rect 5163 27572 5205 27581
rect 5163 27532 5164 27572
rect 5204 27532 5205 27572
rect 5163 27523 5205 27532
rect 5410 27572 5468 27573
rect 5410 27532 5419 27572
rect 5459 27532 5468 27572
rect 5410 27531 5468 27532
rect 5643 27572 5685 27581
rect 5643 27532 5644 27572
rect 5684 27532 5685 27572
rect 5643 27523 5685 27532
rect 6123 27572 6165 27581
rect 6123 27532 6124 27572
rect 6164 27532 6165 27572
rect 6123 27523 6165 27532
rect 7363 27572 7421 27573
rect 7363 27532 7372 27572
rect 7412 27532 7421 27572
rect 7363 27531 7421 27532
rect 7939 27572 7997 27573
rect 7939 27532 7948 27572
rect 7988 27532 7997 27572
rect 7939 27531 7997 27532
rect 9195 27572 9237 27581
rect 9195 27532 9196 27572
rect 9236 27532 9237 27572
rect 9195 27523 9237 27532
rect 9579 27572 9621 27581
rect 9579 27532 9580 27572
rect 9620 27532 9621 27572
rect 9579 27523 9621 27532
rect 10827 27572 10885 27573
rect 10827 27532 10836 27572
rect 10876 27532 10885 27572
rect 10827 27531 10885 27532
rect 11395 27572 11453 27573
rect 11395 27532 11404 27572
rect 11444 27532 11453 27572
rect 11395 27531 11453 27532
rect 12651 27572 12693 27581
rect 12651 27532 12652 27572
rect 12692 27532 12693 27572
rect 12651 27523 12693 27532
rect 13131 27572 13173 27581
rect 13131 27532 13132 27572
rect 13172 27532 13173 27572
rect 13131 27523 13173 27532
rect 14371 27572 14429 27573
rect 14371 27532 14380 27572
rect 14420 27532 14429 27572
rect 14371 27531 14429 27532
rect 15051 27572 15093 27581
rect 15051 27532 15052 27572
rect 15092 27532 15093 27572
rect 15051 27523 15093 27532
rect 16291 27572 16349 27573
rect 16291 27532 16300 27572
rect 16340 27532 16349 27572
rect 16291 27531 16349 27532
rect 16779 27572 16821 27581
rect 16779 27532 16780 27572
rect 16820 27532 16821 27572
rect 16779 27523 16821 27532
rect 18019 27572 18077 27573
rect 18019 27532 18028 27572
rect 18068 27532 18077 27572
rect 18019 27531 18077 27532
rect 18411 27572 18453 27581
rect 18411 27532 18412 27572
rect 18452 27532 18453 27572
rect 18411 27523 18453 27532
rect 19651 27572 19709 27573
rect 19651 27532 19660 27572
rect 19700 27532 19709 27572
rect 19651 27531 19709 27532
rect 19990 27572 20032 27581
rect 19990 27532 19991 27572
rect 20031 27532 20032 27572
rect 19990 27523 20032 27532
rect 20122 27572 20180 27573
rect 20122 27532 20131 27572
rect 20171 27532 20180 27572
rect 20122 27531 20180 27532
rect 20235 27572 20277 27581
rect 20235 27532 20236 27572
rect 20276 27532 20277 27572
rect 20235 27523 20277 27532
rect 4011 27488 4053 27497
rect 4011 27448 4012 27488
rect 4052 27448 4053 27488
rect 4011 27439 4053 27448
rect 4793 27488 4835 27497
rect 4793 27448 4794 27488
rect 4834 27448 4835 27488
rect 4793 27439 4835 27448
rect 19851 27488 19893 27497
rect 19851 27448 19852 27488
rect 19892 27448 19893 27488
rect 19851 27439 19893 27448
rect 3387 27404 3429 27413
rect 3387 27364 3388 27404
rect 3428 27364 3429 27404
rect 3387 27355 3429 27364
rect 4570 27404 4628 27405
rect 4570 27364 4579 27404
rect 4619 27364 4628 27404
rect 4570 27363 4628 27364
rect 4683 27404 4725 27413
rect 4683 27364 4684 27404
rect 4724 27364 4725 27404
rect 4683 27355 4725 27364
rect 7755 27404 7797 27413
rect 7755 27364 7756 27404
rect 7796 27364 7797 27404
rect 7755 27355 7797 27364
rect 16491 27404 16533 27413
rect 16491 27364 16492 27404
rect 16532 27364 16533 27404
rect 16491 27355 16533 27364
rect 18219 27404 18261 27413
rect 18219 27364 18220 27404
rect 18260 27364 18261 27404
rect 18219 27355 18261 27364
rect 20314 27404 20372 27405
rect 20314 27364 20323 27404
rect 20363 27364 20372 27404
rect 20314 27363 20372 27364
rect 1152 27236 20452 27260
rect 1152 27196 4928 27236
rect 4968 27196 5010 27236
rect 5050 27196 5092 27236
rect 5132 27196 5174 27236
rect 5214 27196 5256 27236
rect 5296 27196 20048 27236
rect 20088 27196 20130 27236
rect 20170 27196 20212 27236
rect 20252 27196 20294 27236
rect 20334 27196 20376 27236
rect 20416 27196 20452 27236
rect 1152 27172 20452 27196
rect 2955 27068 2997 27077
rect 2955 27028 2956 27068
rect 2996 27028 2997 27068
rect 2955 27019 2997 27028
rect 7467 27068 7509 27077
rect 7467 27028 7468 27068
rect 7508 27028 7509 27068
rect 7467 27019 7509 27028
rect 7899 27068 7941 27077
rect 7899 27028 7900 27068
rect 7940 27028 7941 27068
rect 7899 27019 7941 27028
rect 10587 27068 10629 27077
rect 10587 27028 10588 27068
rect 10628 27028 10629 27068
rect 10587 27019 10629 27028
rect 11259 27068 11301 27077
rect 11259 27028 11260 27068
rect 11300 27028 11301 27068
rect 11259 27019 11301 27028
rect 20139 27068 20181 27077
rect 20139 27028 20140 27068
rect 20180 27028 20181 27068
rect 20139 27019 20181 27028
rect 3915 26984 3957 26993
rect 3915 26944 3916 26984
rect 3956 26944 3957 26984
rect 3915 26935 3957 26944
rect 17883 26984 17925 26993
rect 17883 26944 17884 26984
rect 17924 26944 17925 26984
rect 17883 26935 17925 26944
rect 1515 26900 1557 26909
rect 3147 26900 3189 26909
rect 1515 26860 1516 26900
rect 1556 26860 1557 26900
rect 1515 26851 1557 26860
rect 2763 26891 2805 26900
rect 2763 26851 2764 26891
rect 2804 26851 2805 26891
rect 3147 26860 3148 26900
rect 3188 26860 3189 26900
rect 3147 26851 3189 26860
rect 3531 26900 3573 26909
rect 3531 26860 3532 26900
rect 3572 26860 3573 26900
rect 3531 26851 3573 26860
rect 3802 26900 3860 26901
rect 3802 26860 3811 26900
rect 3851 26860 3860 26900
rect 3802 26859 3860 26860
rect 4395 26900 4437 26909
rect 6027 26900 6069 26909
rect 8218 26900 8276 26901
rect 4395 26860 4396 26900
rect 4436 26860 4437 26900
rect 4395 26851 4437 26860
rect 5643 26891 5685 26900
rect 5643 26851 5644 26891
rect 5684 26851 5685 26891
rect 6027 26860 6028 26900
rect 6068 26860 6069 26900
rect 6027 26851 6069 26860
rect 7275 26891 7317 26900
rect 7275 26851 7276 26891
rect 7316 26851 7317 26891
rect 8218 26860 8227 26900
rect 8267 26860 8276 26900
rect 8218 26859 8276 26860
rect 8331 26900 8373 26909
rect 8331 26860 8332 26900
rect 8372 26860 8373 26900
rect 8331 26851 8373 26860
rect 8715 26900 8757 26909
rect 9994 26900 10052 26901
rect 12843 26900 12885 26909
rect 8715 26860 8716 26900
rect 8756 26860 8757 26900
rect 8715 26851 8757 26860
rect 9291 26891 9333 26900
rect 9291 26851 9292 26891
rect 9332 26851 9333 26891
rect 2763 26842 2805 26851
rect 5643 26842 5685 26851
rect 7275 26842 7317 26851
rect 9291 26842 9333 26851
rect 9771 26891 9813 26900
rect 9771 26851 9772 26891
rect 9812 26851 9813 26891
rect 9994 26860 10003 26900
rect 10043 26860 10052 26900
rect 9994 26859 10052 26860
rect 11595 26891 11637 26900
rect 9771 26842 9813 26851
rect 11595 26851 11596 26891
rect 11636 26851 11637 26891
rect 12843 26860 12844 26900
rect 12884 26860 12885 26900
rect 12843 26851 12885 26860
rect 13611 26900 13653 26909
rect 15243 26900 15285 26909
rect 16822 26900 16864 26909
rect 13611 26860 13612 26900
rect 13652 26860 13653 26900
rect 13611 26851 13653 26860
rect 14859 26891 14901 26900
rect 14859 26851 14860 26891
rect 14900 26851 14901 26891
rect 15243 26860 15244 26900
rect 15284 26860 15285 26900
rect 15243 26851 15285 26860
rect 16491 26891 16533 26900
rect 16491 26851 16492 26891
rect 16532 26851 16533 26891
rect 16822 26860 16823 26900
rect 16863 26860 16864 26900
rect 16822 26851 16864 26860
rect 17067 26900 17109 26909
rect 17067 26860 17068 26900
rect 17108 26860 17109 26900
rect 17067 26851 17109 26860
rect 18394 26900 18452 26901
rect 18394 26860 18403 26900
rect 18443 26860 18452 26900
rect 18394 26859 18452 26860
rect 18507 26900 18549 26909
rect 18507 26860 18508 26900
rect 18548 26860 18549 26900
rect 18507 26851 18549 26860
rect 18891 26900 18933 26909
rect 18891 26860 18892 26900
rect 18932 26860 18933 26900
rect 18891 26851 18933 26860
rect 19467 26891 19509 26900
rect 19467 26851 19468 26891
rect 19508 26851 19509 26891
rect 11595 26842 11637 26851
rect 14859 26842 14901 26851
rect 16491 26842 16533 26851
rect 19467 26842 19509 26851
rect 19947 26891 19989 26900
rect 19947 26851 19948 26891
rect 19988 26851 19989 26891
rect 19947 26842 19989 26851
rect 7659 26816 7701 26825
rect 7659 26776 7660 26816
rect 7700 26776 7701 26816
rect 7659 26767 7701 26776
rect 8811 26816 8853 26825
rect 8811 26776 8812 26816
rect 8852 26776 8853 26816
rect 8811 26767 8853 26776
rect 10155 26816 10197 26825
rect 10155 26776 10156 26816
rect 10196 26776 10197 26816
rect 10155 26767 10197 26776
rect 10827 26816 10869 26825
rect 10827 26776 10828 26816
rect 10868 26776 10869 26816
rect 10827 26767 10869 26776
rect 11019 26816 11061 26825
rect 11019 26776 11020 26816
rect 11060 26776 11061 26816
rect 11019 26767 11061 26776
rect 13035 26816 13077 26825
rect 13035 26776 13036 26816
rect 13076 26776 13077 26816
rect 13035 26767 13077 26776
rect 16954 26816 17012 26817
rect 16954 26776 16963 26816
rect 17003 26776 17012 26816
rect 16954 26775 17012 26776
rect 17163 26816 17205 26825
rect 17163 26776 17164 26816
rect 17204 26776 17205 26816
rect 17163 26767 17205 26776
rect 17739 26816 17781 26825
rect 17739 26776 17740 26816
rect 17780 26776 17781 26816
rect 17739 26767 17781 26776
rect 18123 26816 18165 26825
rect 18123 26776 18124 26816
rect 18164 26776 18165 26816
rect 18123 26767 18165 26776
rect 18987 26816 19029 26825
rect 18987 26776 18988 26816
rect 19028 26776 19029 26816
rect 18987 26767 19029 26776
rect 10395 26732 10437 26741
rect 10395 26692 10396 26732
rect 10436 26692 10437 26732
rect 10395 26683 10437 26692
rect 3291 26648 3333 26657
rect 3291 26608 3292 26648
rect 3332 26608 3333 26648
rect 3291 26599 3333 26608
rect 4203 26648 4245 26657
rect 4203 26608 4204 26648
rect 4244 26608 4245 26648
rect 4203 26599 4245 26608
rect 5835 26648 5877 26657
rect 5835 26608 5836 26648
rect 5876 26608 5877 26648
rect 5835 26599 5877 26608
rect 11403 26648 11445 26657
rect 11403 26608 11404 26648
rect 11444 26608 11445 26648
rect 11403 26599 11445 26608
rect 13275 26648 13317 26657
rect 13275 26608 13276 26648
rect 13316 26608 13317 26648
rect 13275 26599 13317 26608
rect 15051 26648 15093 26657
rect 15051 26608 15052 26648
rect 15092 26608 15093 26648
rect 15051 26599 15093 26608
rect 16683 26648 16725 26657
rect 16683 26608 16684 26648
rect 16724 26608 16725 26648
rect 16683 26599 16725 26608
rect 17499 26648 17541 26657
rect 17499 26608 17500 26648
rect 17540 26608 17541 26648
rect 17499 26599 17541 26608
rect 1152 26480 20448 26504
rect 1152 26440 3688 26480
rect 3728 26440 3770 26480
rect 3810 26440 3852 26480
rect 3892 26440 3934 26480
rect 3974 26440 4016 26480
rect 4056 26440 18808 26480
rect 18848 26440 18890 26480
rect 18930 26440 18972 26480
rect 19012 26440 19054 26480
rect 19094 26440 19136 26480
rect 19176 26440 20448 26480
rect 1152 26416 20448 26440
rect 4587 26312 4629 26321
rect 4587 26272 4588 26312
rect 4628 26272 4629 26312
rect 4587 26263 4629 26272
rect 5019 26312 5061 26321
rect 5019 26272 5020 26312
rect 5060 26272 5061 26312
rect 5019 26263 5061 26272
rect 5307 26312 5349 26321
rect 5307 26272 5308 26312
rect 5348 26272 5349 26312
rect 5307 26263 5349 26272
rect 7275 26312 7317 26321
rect 7275 26272 7276 26312
rect 7316 26272 7317 26312
rect 7275 26263 7317 26272
rect 9322 26312 9380 26313
rect 9322 26272 9331 26312
rect 9371 26272 9380 26312
rect 9322 26271 9380 26272
rect 13947 26312 13989 26321
rect 13947 26272 13948 26312
rect 13988 26272 13989 26312
rect 13947 26263 13989 26272
rect 20235 26312 20277 26321
rect 20235 26272 20236 26312
rect 20276 26272 20277 26312
rect 20235 26263 20277 26272
rect 15003 26228 15045 26237
rect 15003 26188 15004 26228
rect 15044 26188 15045 26228
rect 15003 26179 15045 26188
rect 3418 26144 3476 26145
rect 3418 26104 3427 26144
rect 3467 26104 3476 26144
rect 3418 26103 3476 26104
rect 4779 26144 4821 26153
rect 4779 26104 4780 26144
rect 4820 26104 4821 26144
rect 4779 26095 4821 26104
rect 5547 26144 5589 26153
rect 5547 26104 5548 26144
rect 5588 26104 5589 26144
rect 5547 26095 5589 26104
rect 8043 26144 8085 26153
rect 8043 26104 8044 26144
rect 8084 26104 8085 26144
rect 8043 26095 8085 26104
rect 10059 26144 10101 26153
rect 10059 26104 10060 26144
rect 10100 26104 10101 26144
rect 10059 26095 10101 26104
rect 11338 26144 11396 26145
rect 11338 26104 11347 26144
rect 11387 26104 11396 26144
rect 11338 26103 11396 26104
rect 11691 26144 11733 26153
rect 11691 26104 11692 26144
rect 11732 26104 11733 26144
rect 11691 26095 11733 26104
rect 11931 26144 11973 26153
rect 11931 26104 11932 26144
rect 11972 26104 11973 26144
rect 11931 26095 11973 26104
rect 13707 26144 13749 26153
rect 13707 26104 13708 26144
rect 13748 26104 13749 26144
rect 13707 26095 13749 26104
rect 14283 26144 14325 26153
rect 14283 26104 14284 26144
rect 14324 26104 14325 26144
rect 14283 26095 14325 26104
rect 14763 26144 14805 26153
rect 14763 26104 14764 26144
rect 14804 26104 14805 26144
rect 14763 26095 14805 26104
rect 15723 26144 15765 26153
rect 15723 26104 15724 26144
rect 15764 26104 15765 26144
rect 15723 26095 15765 26104
rect 1419 26060 1461 26069
rect 1419 26020 1420 26060
rect 1460 26020 1461 26060
rect 1419 26011 1461 26020
rect 2659 26060 2717 26061
rect 2659 26020 2668 26060
rect 2708 26020 2717 26060
rect 2659 26019 2717 26020
rect 3051 26060 3093 26069
rect 3051 26020 3052 26060
rect 3092 26020 3093 26060
rect 3051 26011 3093 26020
rect 3286 26060 3328 26069
rect 3286 26020 3287 26060
rect 3327 26020 3328 26060
rect 3286 26011 3328 26020
rect 3531 26060 3573 26069
rect 3531 26020 3532 26060
rect 3572 26020 3573 26060
rect 3531 26011 3573 26020
rect 3805 26060 3847 26069
rect 3805 26020 3806 26060
rect 3846 26020 3847 26060
rect 3805 26011 3847 26020
rect 4101 26060 4159 26061
rect 4101 26020 4110 26060
rect 4150 26020 4159 26060
rect 4101 26019 4159 26020
rect 4280 26060 4338 26061
rect 4280 26020 4289 26060
rect 4329 26020 4338 26060
rect 4280 26019 4338 26020
rect 4395 26060 4437 26069
rect 4395 26020 4396 26060
rect 4436 26020 4437 26060
rect 4395 26011 4437 26020
rect 5835 26060 5877 26069
rect 5835 26020 5836 26060
rect 5876 26020 5877 26060
rect 5835 26011 5877 26020
rect 7075 26060 7133 26061
rect 7075 26020 7084 26060
rect 7124 26020 7133 26060
rect 7075 26019 7133 26020
rect 7546 26060 7604 26061
rect 7546 26020 7555 26060
rect 7595 26020 7604 26060
rect 7546 26019 7604 26020
rect 7659 26060 7701 26069
rect 7659 26020 7660 26060
rect 7700 26020 7701 26060
rect 7659 26011 7701 26020
rect 8139 26060 8181 26069
rect 8139 26020 8140 26060
rect 8180 26020 8181 26060
rect 8139 26011 8181 26020
rect 8614 26060 8672 26061
rect 8614 26020 8623 26060
rect 8663 26020 8672 26060
rect 8614 26019 8672 26020
rect 9130 26060 9188 26061
rect 9130 26020 9139 26060
rect 9179 26020 9188 26060
rect 9130 26019 9188 26020
rect 9562 26060 9620 26061
rect 9562 26020 9571 26060
rect 9611 26020 9620 26060
rect 9562 26019 9620 26020
rect 9675 26060 9717 26069
rect 9675 26020 9676 26060
rect 9716 26020 9717 26060
rect 9675 26011 9717 26020
rect 10155 26060 10197 26069
rect 10155 26020 10156 26060
rect 10196 26020 10197 26060
rect 10155 26011 10197 26020
rect 10627 26060 10685 26061
rect 10627 26020 10636 26060
rect 10676 26020 10685 26060
rect 10627 26019 10685 26020
rect 11146 26060 11204 26061
rect 11146 26020 11155 26060
rect 11195 26020 11204 26060
rect 11146 26019 11204 26020
rect 12259 26060 12317 26061
rect 12259 26020 12268 26060
rect 12308 26020 12317 26060
rect 12259 26019 12317 26020
rect 13515 26060 13557 26069
rect 13515 26020 13516 26060
rect 13556 26020 13557 26060
rect 13515 26011 13557 26020
rect 15213 26060 15255 26069
rect 15213 26020 15214 26060
rect 15254 26020 15255 26060
rect 15213 26011 15255 26020
rect 15337 26060 15379 26069
rect 15337 26020 15338 26060
rect 15378 26020 15379 26060
rect 15337 26011 15379 26020
rect 15819 26060 15861 26069
rect 15819 26020 15820 26060
rect 15860 26020 15861 26060
rect 15819 26011 15861 26020
rect 16291 26060 16349 26061
rect 16291 26020 16300 26060
rect 16340 26020 16349 26060
rect 16291 26019 16349 26020
rect 16779 26060 16837 26061
rect 16779 26020 16788 26060
rect 16828 26020 16837 26060
rect 16779 26019 16837 26020
rect 17347 26060 17405 26061
rect 17347 26020 17356 26060
rect 17396 26020 17405 26060
rect 17347 26019 17405 26020
rect 18603 26060 18645 26069
rect 18603 26020 18604 26060
rect 18644 26020 18645 26060
rect 18603 26011 18645 26020
rect 18795 26060 18837 26069
rect 18795 26020 18796 26060
rect 18836 26020 18837 26060
rect 18795 26011 18837 26020
rect 20035 26060 20093 26061
rect 20035 26020 20044 26060
rect 20084 26020 20093 26060
rect 20035 26019 20093 26020
rect 3195 25976 3237 25985
rect 3195 25936 3196 25976
rect 3236 25936 3237 25976
rect 3195 25927 3237 25936
rect 4601 25976 4643 25985
rect 4601 25936 4602 25976
rect 4642 25936 4643 25976
rect 4601 25927 4643 25936
rect 12075 25976 12117 25985
rect 12075 25936 12076 25976
rect 12116 25936 12117 25976
rect 12075 25927 12117 25936
rect 14043 25976 14085 25985
rect 14043 25936 14044 25976
rect 14084 25936 14085 25976
rect 14043 25927 14085 25936
rect 17163 25976 17205 25985
rect 17163 25936 17164 25976
rect 17204 25936 17205 25976
rect 17163 25927 17205 25936
rect 2859 25892 2901 25901
rect 2859 25852 2860 25892
rect 2900 25852 2901 25892
rect 2859 25843 2901 25852
rect 3610 25892 3668 25893
rect 3610 25852 3619 25892
rect 3659 25852 3668 25892
rect 3610 25851 3668 25852
rect 3898 25892 3956 25893
rect 3898 25852 3907 25892
rect 3947 25852 3956 25892
rect 3898 25851 3956 25852
rect 4011 25892 4053 25901
rect 4011 25852 4012 25892
rect 4052 25852 4053 25892
rect 4011 25843 4053 25852
rect 16971 25892 17013 25901
rect 16971 25852 16972 25892
rect 17012 25852 17013 25892
rect 16971 25843 17013 25852
rect 1152 25724 20452 25748
rect 1152 25684 4928 25724
rect 4968 25684 5010 25724
rect 5050 25684 5092 25724
rect 5132 25684 5174 25724
rect 5214 25684 5256 25724
rect 5296 25684 20048 25724
rect 20088 25684 20130 25724
rect 20170 25684 20212 25724
rect 20252 25684 20294 25724
rect 20334 25684 20376 25724
rect 20416 25684 20452 25724
rect 1152 25660 20452 25684
rect 3339 25556 3381 25565
rect 3339 25516 3340 25556
rect 3380 25516 3381 25556
rect 3339 25507 3381 25516
rect 5211 25556 5253 25565
rect 5211 25516 5212 25556
rect 5252 25516 5253 25556
rect 5211 25507 5253 25516
rect 9099 25556 9141 25565
rect 9099 25516 9100 25556
rect 9140 25516 9141 25556
rect 9099 25507 9141 25516
rect 11115 25556 11157 25565
rect 11115 25516 11116 25556
rect 11156 25516 11157 25556
rect 11115 25507 11157 25516
rect 11403 25556 11445 25565
rect 11403 25516 11404 25556
rect 11444 25516 11445 25556
rect 11403 25507 11445 25516
rect 20379 25556 20421 25565
rect 20379 25516 20380 25556
rect 20420 25516 20421 25556
rect 20379 25507 20421 25516
rect 1467 25472 1509 25481
rect 1467 25432 1468 25472
rect 1508 25432 1509 25472
rect 1467 25423 1509 25432
rect 3771 25472 3813 25481
rect 3771 25432 3772 25472
rect 3812 25432 3813 25472
rect 3771 25423 3813 25432
rect 4155 25472 4197 25481
rect 4155 25432 4156 25472
rect 4196 25432 4197 25472
rect 4155 25423 4197 25432
rect 15915 25472 15957 25481
rect 15915 25432 15916 25472
rect 15956 25432 15957 25472
rect 15915 25423 15957 25432
rect 19995 25472 20037 25481
rect 19995 25432 19996 25472
rect 20036 25432 20037 25472
rect 19995 25423 20037 25432
rect 1899 25388 1941 25397
rect 5355 25388 5397 25397
rect 7659 25388 7701 25397
rect 9357 25388 9399 25397
rect 1899 25348 1900 25388
rect 1940 25348 1941 25388
rect 1899 25339 1941 25348
rect 3147 25379 3189 25388
rect 3147 25339 3148 25379
rect 3188 25339 3189 25379
rect 5355 25348 5356 25388
rect 5396 25348 5397 25388
rect 5355 25339 5397 25348
rect 6603 25379 6645 25388
rect 6603 25339 6604 25379
rect 6644 25339 6645 25379
rect 7659 25348 7660 25388
rect 7700 25348 7701 25388
rect 7659 25339 7701 25348
rect 8907 25379 8949 25388
rect 8907 25339 8908 25379
rect 8948 25339 8949 25379
rect 9357 25348 9358 25388
rect 9398 25348 9399 25388
rect 9357 25339 9399 25348
rect 9472 25388 9530 25389
rect 9472 25348 9481 25388
rect 9521 25348 9530 25388
rect 9472 25347 9530 25348
rect 9860 25388 9902 25397
rect 9860 25348 9861 25388
rect 9901 25348 9902 25388
rect 9860 25339 9902 25348
rect 9963 25388 10005 25397
rect 12843 25388 12885 25397
rect 9963 25348 9964 25388
rect 10004 25348 10005 25388
rect 9963 25339 10005 25348
rect 10443 25379 10485 25388
rect 10443 25339 10444 25379
rect 10484 25339 10485 25379
rect 3147 25330 3189 25339
rect 6603 25330 6645 25339
rect 8907 25330 8949 25339
rect 10443 25330 10485 25339
rect 10923 25379 10965 25388
rect 10923 25339 10924 25379
rect 10964 25339 10965 25379
rect 10923 25330 10965 25339
rect 11595 25379 11637 25388
rect 11595 25339 11596 25379
rect 11636 25339 11637 25379
rect 12843 25348 12844 25388
rect 12884 25348 12885 25388
rect 12843 25339 12885 25348
rect 14187 25388 14229 25397
rect 14187 25348 14188 25388
rect 14228 25348 14229 25388
rect 14187 25339 14229 25348
rect 14475 25388 14517 25397
rect 16186 25388 16244 25389
rect 14475 25348 14476 25388
rect 14516 25348 14517 25388
rect 14475 25339 14517 25348
rect 15723 25379 15765 25388
rect 15723 25339 15724 25379
rect 15764 25339 15765 25379
rect 16186 25348 16195 25388
rect 16235 25348 16244 25388
rect 16186 25347 16244 25348
rect 16299 25388 16341 25397
rect 16299 25348 16300 25388
rect 16340 25348 16341 25388
rect 16299 25339 16341 25348
rect 16683 25388 16725 25397
rect 18123 25388 18165 25397
rect 16683 25348 16684 25388
rect 16724 25348 16725 25388
rect 16683 25339 16725 25348
rect 17259 25379 17301 25388
rect 17259 25339 17260 25379
rect 17300 25339 17301 25379
rect 11595 25330 11637 25339
rect 15723 25330 15765 25339
rect 17259 25330 17301 25339
rect 17739 25379 17781 25388
rect 17739 25339 17740 25379
rect 17780 25339 17781 25379
rect 18123 25348 18124 25388
rect 18164 25348 18165 25388
rect 18123 25339 18165 25348
rect 19371 25379 19413 25388
rect 19371 25339 19372 25379
rect 19412 25339 19413 25379
rect 17739 25330 17781 25339
rect 19371 25330 19413 25339
rect 1227 25304 1269 25313
rect 1227 25264 1228 25304
rect 1268 25264 1269 25304
rect 1227 25255 1269 25264
rect 3531 25304 3573 25313
rect 3531 25264 3532 25304
rect 3572 25264 3573 25304
rect 3531 25255 3573 25264
rect 3915 25304 3957 25313
rect 3915 25264 3916 25304
rect 3956 25264 3957 25304
rect 3915 25255 3957 25264
rect 4587 25304 4629 25313
rect 4587 25264 4588 25304
rect 4628 25264 4629 25304
rect 4587 25255 4629 25264
rect 4971 25304 5013 25313
rect 4971 25264 4972 25304
rect 5012 25264 5013 25304
rect 4971 25255 5013 25264
rect 5211 25304 5253 25313
rect 5211 25264 5212 25304
rect 5252 25264 5253 25304
rect 5211 25255 5253 25264
rect 7179 25304 7221 25313
rect 7179 25264 7180 25304
rect 7220 25264 7221 25304
rect 7179 25255 7221 25264
rect 13803 25304 13845 25313
rect 13803 25264 13804 25304
rect 13844 25264 13845 25304
rect 13803 25255 13845 25264
rect 16779 25304 16821 25313
rect 16779 25264 16780 25304
rect 16820 25264 16821 25304
rect 16779 25255 16821 25264
rect 19755 25304 19797 25313
rect 19755 25264 19756 25304
rect 19796 25264 19797 25304
rect 19755 25255 19797 25264
rect 20139 25304 20181 25313
rect 20139 25264 20140 25304
rect 20180 25264 20181 25304
rect 20139 25255 20181 25264
rect 6939 25220 6981 25229
rect 6939 25180 6940 25220
rect 6980 25180 6981 25220
rect 6939 25171 6981 25180
rect 17979 25220 18021 25229
rect 17979 25180 17980 25220
rect 18020 25180 18021 25220
rect 17979 25171 18021 25180
rect 4347 25136 4389 25145
rect 4347 25096 4348 25136
rect 4388 25096 4389 25136
rect 4347 25087 4389 25096
rect 6795 25136 6837 25145
rect 6795 25096 6796 25136
rect 6836 25096 6837 25136
rect 6795 25087 6837 25096
rect 13563 25136 13605 25145
rect 13563 25096 13564 25136
rect 13604 25096 13605 25136
rect 13563 25087 13605 25096
rect 14331 25136 14373 25145
rect 14331 25096 14332 25136
rect 14372 25096 14373 25136
rect 14331 25087 14373 25096
rect 19563 25136 19605 25145
rect 19563 25096 19564 25136
rect 19604 25096 19605 25136
rect 19563 25087 19605 25096
rect 1152 24968 20448 24992
rect 1152 24928 3688 24968
rect 3728 24928 3770 24968
rect 3810 24928 3852 24968
rect 3892 24928 3934 24968
rect 3974 24928 4016 24968
rect 4056 24928 18808 24968
rect 18848 24928 18890 24968
rect 18930 24928 18972 24968
rect 19012 24928 19054 24968
rect 19094 24928 19136 24968
rect 19176 24928 20448 24968
rect 1152 24904 20448 24928
rect 5211 24800 5253 24809
rect 5211 24760 5212 24800
rect 5252 24760 5253 24800
rect 5211 24751 5253 24760
rect 5979 24800 6021 24809
rect 5979 24760 5980 24800
rect 6020 24760 6021 24800
rect 5979 24751 6021 24760
rect 9723 24800 9765 24809
rect 9723 24760 9724 24800
rect 9764 24760 9765 24800
rect 9723 24751 9765 24760
rect 11307 24800 11349 24809
rect 11307 24760 11308 24800
rect 11348 24760 11349 24800
rect 11307 24751 11349 24760
rect 15195 24800 15237 24809
rect 15195 24760 15196 24800
rect 15236 24760 15237 24800
rect 15195 24751 15237 24760
rect 19227 24800 19269 24809
rect 19227 24760 19228 24800
rect 19268 24760 19269 24800
rect 19227 24751 19269 24760
rect 19995 24800 20037 24809
rect 19995 24760 19996 24800
rect 20036 24760 20037 24800
rect 19995 24751 20037 24760
rect 20379 24800 20421 24809
rect 20379 24760 20380 24800
rect 20420 24760 20421 24800
rect 20379 24751 20421 24760
rect 2763 24716 2805 24725
rect 2763 24676 2764 24716
rect 2804 24676 2805 24716
rect 2763 24667 2805 24676
rect 5307 24716 5349 24725
rect 5307 24676 5308 24716
rect 5348 24676 5349 24716
rect 5307 24667 5349 24676
rect 8955 24716 8997 24725
rect 8955 24676 8956 24716
rect 8996 24676 8997 24716
rect 8955 24667 8997 24676
rect 9339 24716 9381 24725
rect 9339 24676 9340 24716
rect 9380 24676 9381 24716
rect 9339 24667 9381 24676
rect 14763 24716 14805 24725
rect 14763 24676 14764 24716
rect 14804 24676 14805 24716
rect 14763 24667 14805 24676
rect 16779 24716 16821 24725
rect 16779 24676 16780 24716
rect 16820 24676 16821 24716
rect 16779 24667 16821 24676
rect 3531 24632 3573 24641
rect 3531 24592 3532 24632
rect 3572 24592 3573 24632
rect 3531 24583 3573 24592
rect 4971 24632 5013 24641
rect 4971 24592 4972 24632
rect 5012 24592 5013 24632
rect 4971 24583 5013 24592
rect 5547 24632 5589 24641
rect 5547 24592 5548 24632
rect 5588 24592 5589 24632
rect 5547 24583 5589 24592
rect 5739 24632 5781 24641
rect 5739 24592 5740 24632
rect 5780 24592 5781 24632
rect 5739 24583 5781 24592
rect 6891 24632 6933 24641
rect 6891 24592 6892 24632
rect 6932 24592 6933 24632
rect 6891 24583 6933 24592
rect 8170 24632 8228 24633
rect 8170 24592 8179 24632
rect 8219 24592 8228 24632
rect 8170 24591 8228 24592
rect 8331 24632 8373 24641
rect 8331 24592 8332 24632
rect 8372 24592 8373 24632
rect 8331 24583 8373 24592
rect 8571 24632 8613 24641
rect 8571 24592 8572 24632
rect 8612 24592 8613 24632
rect 8571 24583 8613 24592
rect 8715 24632 8757 24641
rect 8715 24592 8716 24632
rect 8756 24592 8757 24632
rect 8715 24583 8757 24592
rect 9099 24632 9141 24641
rect 9099 24592 9100 24632
rect 9140 24592 9141 24632
rect 9099 24583 9141 24592
rect 9483 24632 9525 24641
rect 9483 24592 9484 24632
rect 9524 24592 9525 24632
rect 9483 24583 9525 24592
rect 14955 24632 14997 24641
rect 14955 24592 14956 24632
rect 14996 24592 14997 24632
rect 14955 24583 14997 24592
rect 17547 24632 17589 24641
rect 17547 24592 17548 24632
rect 17588 24592 17589 24632
rect 17547 24583 17589 24592
rect 18987 24632 19029 24641
rect 18987 24592 18988 24632
rect 19028 24592 19029 24632
rect 18603 24581 18645 24590
rect 18987 24583 19029 24592
rect 19371 24632 19413 24641
rect 19371 24592 19372 24632
rect 19412 24592 19413 24632
rect 19371 24583 19413 24592
rect 19611 24632 19653 24641
rect 19611 24592 19612 24632
rect 19652 24592 19653 24632
rect 19611 24583 19653 24592
rect 19755 24632 19797 24641
rect 19755 24592 19756 24632
rect 19796 24592 19797 24632
rect 19755 24583 19797 24592
rect 20139 24632 20181 24641
rect 20139 24592 20140 24632
rect 20180 24592 20181 24632
rect 20139 24583 20181 24592
rect 1323 24548 1365 24557
rect 1323 24508 1324 24548
rect 1364 24508 1365 24548
rect 1323 24499 1365 24508
rect 2563 24548 2621 24549
rect 2563 24508 2572 24548
rect 2612 24508 2621 24548
rect 2563 24507 2621 24508
rect 3034 24548 3092 24549
rect 3034 24508 3043 24548
rect 3083 24508 3092 24548
rect 3034 24507 3092 24508
rect 3147 24548 3189 24557
rect 3147 24508 3148 24548
rect 3188 24508 3189 24548
rect 3147 24499 3189 24508
rect 3627 24548 3669 24557
rect 3627 24508 3628 24548
rect 3668 24508 3669 24548
rect 3627 24499 3669 24508
rect 4099 24548 4157 24549
rect 4099 24508 4108 24548
rect 4148 24508 4157 24548
rect 4099 24507 4157 24508
rect 4587 24548 4645 24549
rect 4587 24508 4596 24548
rect 4636 24508 4645 24548
rect 4587 24507 4645 24508
rect 6394 24548 6452 24549
rect 6394 24508 6403 24548
rect 6443 24508 6452 24548
rect 6394 24507 6452 24508
rect 6507 24548 6549 24557
rect 6507 24508 6508 24548
rect 6548 24508 6549 24548
rect 6507 24499 6549 24508
rect 6987 24548 7029 24557
rect 6987 24508 6988 24548
rect 7028 24508 7029 24548
rect 6987 24499 7029 24508
rect 7459 24548 7517 24549
rect 7459 24508 7468 24548
rect 7508 24508 7517 24548
rect 7459 24507 7517 24508
rect 7947 24548 8005 24549
rect 7947 24508 7956 24548
rect 7996 24508 8005 24548
rect 7947 24507 8005 24508
rect 9867 24548 9909 24557
rect 9867 24508 9868 24548
rect 9908 24508 9909 24548
rect 9867 24499 9909 24508
rect 11107 24548 11165 24549
rect 11107 24508 11116 24548
rect 11156 24508 11165 24548
rect 11107 24507 11165 24508
rect 11499 24548 11541 24557
rect 11499 24508 11500 24548
rect 11540 24508 11541 24548
rect 11499 24499 11541 24508
rect 12739 24548 12797 24549
rect 12739 24508 12748 24548
rect 12788 24508 12797 24548
rect 12739 24507 12797 24508
rect 13323 24548 13365 24557
rect 13323 24508 13324 24548
rect 13364 24508 13365 24548
rect 13323 24499 13365 24508
rect 14563 24548 14621 24549
rect 14563 24508 14572 24548
rect 14612 24508 14621 24548
rect 14563 24507 14621 24508
rect 15339 24548 15381 24557
rect 15339 24508 15340 24548
rect 15380 24508 15381 24548
rect 15339 24499 15381 24508
rect 16579 24548 16637 24549
rect 16579 24508 16588 24548
rect 16628 24508 16637 24548
rect 16579 24507 16637 24508
rect 17050 24548 17108 24549
rect 17050 24508 17059 24548
rect 17099 24508 17108 24548
rect 17050 24507 17108 24508
rect 17163 24548 17205 24557
rect 17163 24508 17164 24548
rect 17204 24508 17205 24548
rect 17163 24499 17205 24508
rect 17643 24548 17685 24557
rect 17643 24508 17644 24548
rect 17684 24508 17685 24548
rect 17643 24499 17685 24508
rect 18115 24548 18173 24549
rect 18115 24508 18124 24548
rect 18164 24508 18173 24548
rect 18603 24541 18604 24581
rect 18644 24541 18645 24581
rect 18603 24532 18645 24541
rect 18115 24507 18173 24508
rect 4779 24380 4821 24389
rect 4779 24340 4780 24380
rect 4820 24340 4821 24380
rect 4779 24331 4821 24340
rect 12939 24380 12981 24389
rect 12939 24340 12940 24380
rect 12980 24340 12981 24380
rect 12939 24331 12981 24340
rect 18795 24380 18837 24389
rect 18795 24340 18796 24380
rect 18836 24340 18837 24380
rect 18795 24331 18837 24340
rect 1152 24212 20452 24236
rect 1152 24172 4928 24212
rect 4968 24172 5010 24212
rect 5050 24172 5092 24212
rect 5132 24172 5174 24212
rect 5214 24172 5256 24212
rect 5296 24172 20048 24212
rect 20088 24172 20130 24212
rect 20170 24172 20212 24212
rect 20252 24172 20294 24212
rect 20334 24172 20376 24212
rect 20416 24172 20452 24212
rect 1152 24148 20452 24172
rect 4779 24044 4821 24053
rect 4779 24004 4780 24044
rect 4820 24004 4821 24044
rect 4779 23995 4821 24004
rect 7467 24044 7509 24053
rect 7467 24004 7468 24044
rect 7508 24004 7509 24044
rect 7467 23995 7509 24004
rect 9291 24044 9333 24053
rect 9291 24004 9292 24044
rect 9332 24004 9333 24044
rect 9291 23995 9333 24004
rect 9723 24044 9765 24053
rect 9723 24004 9724 24044
rect 9764 24004 9765 24044
rect 9723 23995 9765 24004
rect 15723 24044 15765 24053
rect 15723 24004 15724 24044
rect 15764 24004 15765 24044
rect 15723 23995 15765 24004
rect 16731 24044 16773 24053
rect 16731 24004 16732 24044
rect 16772 24004 16773 24044
rect 16731 23995 16773 24004
rect 17499 24044 17541 24053
rect 17499 24004 17500 24044
rect 17540 24004 17541 24044
rect 17499 23995 17541 24004
rect 19546 24044 19604 24045
rect 19546 24004 19555 24044
rect 19595 24004 19604 24044
rect 19546 24003 19604 24004
rect 2763 23960 2805 23969
rect 2763 23920 2764 23960
rect 2804 23920 2805 23960
rect 2763 23911 2805 23920
rect 9819 23960 9861 23969
rect 9819 23920 9820 23960
rect 9860 23920 9861 23960
rect 9819 23911 9861 23920
rect 11979 23960 12021 23969
rect 11979 23920 11980 23960
rect 12020 23920 12021 23960
rect 11979 23911 12021 23920
rect 18843 23960 18885 23969
rect 18843 23920 18844 23960
rect 18884 23920 18885 23960
rect 18843 23911 18885 23920
rect 19258 23960 19316 23961
rect 19258 23920 19267 23960
rect 19307 23920 19316 23960
rect 19258 23919 19316 23920
rect 19766 23960 19808 23969
rect 19766 23920 19767 23960
rect 19807 23920 19808 23960
rect 19766 23911 19808 23920
rect 20139 23960 20181 23969
rect 20139 23920 20140 23960
rect 20180 23920 20181 23960
rect 20139 23911 20181 23920
rect 1323 23876 1365 23885
rect 3034 23876 3092 23877
rect 1323 23836 1324 23876
rect 1364 23836 1365 23876
rect 1323 23827 1365 23836
rect 2571 23867 2613 23876
rect 2571 23827 2572 23867
rect 2612 23827 2613 23867
rect 3034 23836 3043 23876
rect 3083 23836 3092 23876
rect 3034 23835 3092 23836
rect 3147 23876 3189 23885
rect 3147 23836 3148 23876
rect 3188 23836 3189 23876
rect 3147 23827 3189 23836
rect 3531 23876 3573 23885
rect 6027 23876 6069 23885
rect 7851 23876 7893 23885
rect 10539 23876 10581 23885
rect 12171 23876 12213 23885
rect 13978 23876 14036 23877
rect 3531 23836 3532 23876
rect 3572 23836 3573 23876
rect 3531 23827 3573 23836
rect 4107 23867 4149 23876
rect 4107 23827 4108 23867
rect 4148 23827 4149 23867
rect 2571 23818 2613 23827
rect 4107 23818 4149 23827
rect 4587 23867 4629 23876
rect 4587 23827 4588 23867
rect 4628 23827 4629 23867
rect 6027 23836 6028 23876
rect 6068 23836 6069 23876
rect 6027 23827 6069 23836
rect 7275 23867 7317 23876
rect 7275 23827 7276 23867
rect 7316 23827 7317 23867
rect 7851 23836 7852 23876
rect 7892 23836 7893 23876
rect 7851 23827 7893 23836
rect 9099 23867 9141 23876
rect 9099 23827 9100 23867
rect 9140 23827 9141 23867
rect 10539 23836 10540 23876
rect 10580 23836 10581 23876
rect 10539 23827 10581 23836
rect 11787 23867 11829 23876
rect 11787 23827 11788 23867
rect 11828 23827 11829 23867
rect 12171 23836 12172 23876
rect 12212 23836 12213 23876
rect 12171 23827 12213 23836
rect 13419 23867 13461 23876
rect 13419 23827 13420 23867
rect 13460 23827 13461 23867
rect 13978 23836 13987 23876
rect 14027 23836 14036 23876
rect 13978 23835 14036 23836
rect 14091 23876 14133 23885
rect 14091 23836 14092 23876
rect 14132 23836 14133 23876
rect 14091 23827 14133 23836
rect 14475 23876 14517 23885
rect 18946 23876 19004 23877
rect 14475 23836 14476 23876
rect 14516 23836 14517 23876
rect 14475 23827 14517 23836
rect 15051 23867 15093 23876
rect 15051 23827 15052 23867
rect 15092 23827 15093 23867
rect 4587 23818 4629 23827
rect 7275 23818 7317 23827
rect 9099 23818 9141 23827
rect 11787 23818 11829 23827
rect 13419 23818 13461 23827
rect 15051 23818 15093 23827
rect 15531 23867 15573 23876
rect 15531 23827 15532 23867
rect 15572 23827 15573 23867
rect 18946 23836 18955 23876
rect 18995 23836 19004 23876
rect 18946 23835 19004 23836
rect 19177 23876 19219 23885
rect 19177 23836 19178 23876
rect 19218 23836 19219 23876
rect 19177 23827 19219 23836
rect 19450 23876 19508 23877
rect 19450 23836 19459 23876
rect 19499 23836 19508 23876
rect 19450 23835 19508 23836
rect 19933 23876 19975 23885
rect 19933 23836 19934 23876
rect 19974 23836 19975 23876
rect 19933 23827 19975 23836
rect 20235 23867 20277 23876
rect 20235 23827 20236 23867
rect 20276 23827 20277 23867
rect 15531 23818 15573 23827
rect 20235 23818 20277 23827
rect 3627 23792 3669 23801
rect 3627 23752 3628 23792
rect 3668 23752 3669 23792
rect 3627 23743 3669 23752
rect 4971 23792 5013 23801
rect 4971 23752 4972 23792
rect 5012 23752 5013 23792
rect 4971 23743 5013 23752
rect 5355 23792 5397 23801
rect 5355 23752 5356 23792
rect 5396 23752 5397 23792
rect 5355 23743 5397 23752
rect 9483 23792 9525 23801
rect 9483 23752 9484 23792
rect 9524 23752 9525 23792
rect 9483 23743 9525 23752
rect 10059 23792 10101 23801
rect 10059 23752 10060 23792
rect 10100 23752 10101 23792
rect 10059 23743 10101 23752
rect 14571 23792 14613 23801
rect 14571 23752 14572 23792
rect 14612 23752 14613 23792
rect 14571 23743 14613 23752
rect 16107 23792 16149 23801
rect 16107 23752 16108 23792
rect 16148 23752 16149 23792
rect 16107 23743 16149 23752
rect 16491 23792 16533 23801
rect 16491 23752 16492 23792
rect 16532 23752 16533 23792
rect 16491 23743 16533 23752
rect 16875 23792 16917 23801
rect 16875 23752 16876 23792
rect 16916 23752 16917 23792
rect 16875 23743 16917 23752
rect 17259 23792 17301 23801
rect 17259 23752 17260 23792
rect 17300 23752 17301 23792
rect 17259 23743 17301 23752
rect 17835 23792 17877 23801
rect 17835 23752 17836 23792
rect 17876 23752 17877 23792
rect 17835 23743 17877 23752
rect 17979 23792 18021 23801
rect 17979 23752 17980 23792
rect 18020 23752 18021 23792
rect 17979 23743 18021 23752
rect 18219 23792 18261 23801
rect 18219 23752 18220 23792
rect 18260 23752 18261 23792
rect 18219 23743 18261 23752
rect 18603 23792 18645 23801
rect 18603 23752 18604 23792
rect 18644 23752 18645 23792
rect 18603 23743 18645 23752
rect 19066 23792 19124 23793
rect 19066 23752 19075 23792
rect 19115 23752 19124 23792
rect 19066 23751 19124 23752
rect 5211 23624 5253 23633
rect 5211 23584 5212 23624
rect 5252 23584 5253 23624
rect 5211 23575 5253 23584
rect 5595 23624 5637 23633
rect 5595 23584 5596 23624
rect 5636 23584 5637 23624
rect 5595 23575 5637 23584
rect 13611 23624 13653 23633
rect 13611 23584 13612 23624
rect 13652 23584 13653 23624
rect 13611 23575 13653 23584
rect 15867 23624 15909 23633
rect 15867 23584 15868 23624
rect 15908 23584 15909 23624
rect 15867 23575 15909 23584
rect 17115 23624 17157 23633
rect 17115 23584 17116 23624
rect 17156 23584 17157 23624
rect 17115 23575 17157 23584
rect 17595 23624 17637 23633
rect 17595 23584 17596 23624
rect 17636 23584 17637 23624
rect 17595 23575 17637 23584
rect 19755 23624 19797 23633
rect 19755 23584 19756 23624
rect 19796 23584 19797 23624
rect 19755 23575 19797 23584
rect 19930 23624 19988 23625
rect 19930 23584 19939 23624
rect 19979 23584 19988 23624
rect 19930 23583 19988 23584
rect 1152 23456 20448 23480
rect 1152 23416 3688 23456
rect 3728 23416 3770 23456
rect 3810 23416 3852 23456
rect 3892 23416 3934 23456
rect 3974 23416 4016 23456
rect 4056 23416 18808 23456
rect 18848 23416 18890 23456
rect 18930 23416 18972 23456
rect 19012 23416 19054 23456
rect 19094 23416 19136 23456
rect 19176 23416 20448 23456
rect 1152 23392 20448 23416
rect 3339 23288 3381 23297
rect 3339 23248 3340 23288
rect 3380 23248 3381 23288
rect 3339 23239 3381 23248
rect 4155 23288 4197 23297
rect 4155 23248 4156 23288
rect 4196 23248 4197 23288
rect 4155 23239 4197 23248
rect 10474 23288 10532 23289
rect 10474 23248 10483 23288
rect 10523 23248 10532 23288
rect 10474 23247 10532 23248
rect 10971 23288 11013 23297
rect 10971 23248 10972 23288
rect 11012 23248 11013 23288
rect 10971 23239 11013 23248
rect 11643 23288 11685 23297
rect 11643 23248 11644 23288
rect 11684 23248 11685 23288
rect 11643 23239 11685 23248
rect 15562 23288 15620 23289
rect 15562 23248 15571 23288
rect 15611 23248 15620 23288
rect 15562 23247 15620 23248
rect 17674 23288 17732 23289
rect 17674 23248 17683 23288
rect 17723 23248 17732 23288
rect 17674 23247 17732 23248
rect 18459 23288 18501 23297
rect 18459 23248 18460 23288
rect 18500 23248 18501 23288
rect 18459 23239 18501 23248
rect 1467 23204 1509 23213
rect 1467 23164 1468 23204
rect 1508 23164 1509 23204
rect 1467 23155 1509 23164
rect 3706 23204 3764 23205
rect 3706 23164 3715 23204
rect 3755 23164 3764 23204
rect 3706 23163 3764 23164
rect 4539 23204 4581 23213
rect 4539 23164 4540 23204
rect 4580 23164 4581 23204
rect 4539 23155 4581 23164
rect 10875 23204 10917 23213
rect 10875 23164 10876 23204
rect 10916 23164 10917 23204
rect 10875 23155 10917 23164
rect 20187 23204 20229 23213
rect 20187 23164 20188 23204
rect 20228 23164 20229 23204
rect 20187 23155 20229 23164
rect 1227 23120 1269 23129
rect 1227 23080 1228 23120
rect 1268 23080 1269 23120
rect 1227 23071 1269 23080
rect 3915 23120 3957 23129
rect 3915 23080 3916 23120
rect 3956 23080 3957 23120
rect 3915 23071 3957 23080
rect 4299 23120 4341 23129
rect 4299 23080 4300 23120
rect 4340 23080 4341 23120
rect 4299 23071 4341 23080
rect 7179 23120 7221 23129
rect 7179 23080 7180 23120
rect 7220 23080 7221 23120
rect 7179 23071 7221 23080
rect 9195 23120 9237 23129
rect 9195 23080 9196 23120
rect 9236 23080 9237 23120
rect 9195 23071 9237 23080
rect 10635 23120 10677 23129
rect 10635 23080 10636 23120
rect 10676 23080 10677 23120
rect 10635 23071 10677 23080
rect 11211 23120 11253 23129
rect 11211 23080 11212 23120
rect 11252 23080 11253 23120
rect 11211 23071 11253 23080
rect 11883 23120 11925 23129
rect 11883 23080 11884 23120
rect 11924 23080 11925 23120
rect 11883 23071 11925 23080
rect 14283 23120 14325 23129
rect 14283 23080 14284 23120
rect 14324 23080 14325 23120
rect 14283 23071 14325 23080
rect 16395 23120 16437 23129
rect 16395 23080 16396 23120
rect 16436 23080 16437 23120
rect 16395 23071 16437 23080
rect 17787 23120 17829 23129
rect 17787 23080 17788 23120
rect 17828 23080 17829 23120
rect 17787 23071 17829 23080
rect 18027 23120 18069 23129
rect 18027 23080 18028 23120
rect 18068 23080 18069 23120
rect 18027 23071 18069 23080
rect 18219 23120 18261 23129
rect 18219 23080 18220 23120
rect 18260 23080 18261 23120
rect 18219 23071 18261 23080
rect 1899 23036 1941 23045
rect 1899 22996 1900 23036
rect 1940 22996 1941 23036
rect 1899 22987 1941 22996
rect 3139 23036 3197 23037
rect 3139 22996 3148 23036
rect 3188 22996 3197 23036
rect 3139 22995 3197 22996
rect 3531 23036 3573 23045
rect 3531 22996 3532 23036
rect 3572 22996 3573 23036
rect 3531 22987 3573 22996
rect 3706 23036 3764 23037
rect 3706 22996 3715 23036
rect 3755 22996 3764 23036
rect 3706 22995 3764 22996
rect 4683 23036 4725 23045
rect 4683 22996 4684 23036
rect 4724 22996 4725 23036
rect 4683 22987 4725 22996
rect 5923 23036 5981 23037
rect 5923 22996 5932 23036
rect 5972 22996 5981 23036
rect 5923 22995 5981 22996
rect 6682 23036 6740 23037
rect 6682 22996 6691 23036
rect 6731 22996 6740 23036
rect 6682 22995 6740 22996
rect 6795 23036 6837 23045
rect 6795 22996 6796 23036
rect 6836 22996 6837 23036
rect 6795 22987 6837 22996
rect 7275 23036 7317 23045
rect 7275 22996 7276 23036
rect 7316 22996 7317 23036
rect 7275 22987 7317 22996
rect 7747 23036 7805 23037
rect 7747 22996 7756 23036
rect 7796 22996 7805 23036
rect 7747 22995 7805 22996
rect 8235 23036 8293 23037
rect 8235 22996 8244 23036
rect 8284 22996 8293 23036
rect 8235 22995 8293 22996
rect 8698 23036 8756 23037
rect 8698 22996 8707 23036
rect 8747 22996 8756 23036
rect 8698 22995 8756 22996
rect 8811 23036 8853 23045
rect 8811 22996 8812 23036
rect 8852 22996 8853 23036
rect 8811 22987 8853 22996
rect 9291 23036 9333 23045
rect 9291 22996 9292 23036
rect 9332 22996 9333 23036
rect 9291 22987 9333 22996
rect 9763 23036 9821 23037
rect 9763 22996 9772 23036
rect 9812 22996 9821 23036
rect 9763 22995 9821 22996
rect 10282 23036 10340 23037
rect 10282 22996 10291 23036
rect 10331 22996 10340 23036
rect 10282 22995 10340 22996
rect 12075 23036 12117 23045
rect 12075 22996 12076 23036
rect 12116 22996 12117 23036
rect 12075 22987 12117 22996
rect 13315 23036 13373 23037
rect 13315 22996 13324 23036
rect 13364 22996 13373 23036
rect 13315 22995 13373 22996
rect 13786 23036 13844 23037
rect 13786 22996 13795 23036
rect 13835 22996 13844 23036
rect 13786 22995 13844 22996
rect 13899 23036 13941 23045
rect 13899 22996 13900 23036
rect 13940 22996 13941 23036
rect 13899 22987 13941 22996
rect 14379 23036 14421 23045
rect 14379 22996 14380 23036
rect 14420 22996 14421 23036
rect 14379 22987 14421 22996
rect 14851 23036 14909 23037
rect 14851 22996 14860 23036
rect 14900 22996 14909 23036
rect 14851 22995 14909 22996
rect 15339 23036 15397 23037
rect 15339 22996 15348 23036
rect 15388 22996 15397 23036
rect 15339 22995 15397 22996
rect 15898 23036 15956 23037
rect 15898 22996 15907 23036
rect 15947 22996 15956 23036
rect 15898 22995 15956 22996
rect 16011 23036 16053 23045
rect 16011 22996 16012 23036
rect 16052 22996 16053 23036
rect 16011 22987 16053 22996
rect 16491 23036 16533 23045
rect 16491 22996 16492 23036
rect 16532 22996 16533 23036
rect 16491 22987 16533 22996
rect 16963 23036 17021 23037
rect 16963 22996 16972 23036
rect 17012 22996 17021 23036
rect 16963 22995 17021 22996
rect 17482 23036 17540 23037
rect 17482 22996 17491 23036
rect 17531 22996 17540 23036
rect 17482 22995 17540 22996
rect 18603 23036 18645 23045
rect 18603 22996 18604 23036
rect 18644 22996 18645 23036
rect 18603 22987 18645 22996
rect 19843 23036 19901 23037
rect 19843 22996 19852 23036
rect 19892 22996 19901 23036
rect 19843 22995 19901 22996
rect 20331 23036 20373 23045
rect 20331 22996 20332 23036
rect 20372 22996 20373 23036
rect 20331 22987 20373 22996
rect 6123 22952 6165 22961
rect 6123 22912 6124 22952
rect 6164 22912 6165 22952
rect 6123 22903 6165 22912
rect 8427 22868 8469 22877
rect 8427 22828 8428 22868
rect 8468 22828 8469 22868
rect 8427 22819 8469 22828
rect 13515 22868 13557 22877
rect 13515 22828 13516 22868
rect 13556 22828 13557 22868
rect 13515 22819 13557 22828
rect 20043 22868 20085 22877
rect 20043 22828 20044 22868
rect 20084 22828 20085 22868
rect 20043 22819 20085 22828
rect 1152 22700 20452 22724
rect 1152 22660 4928 22700
rect 4968 22660 5010 22700
rect 5050 22660 5092 22700
rect 5132 22660 5174 22700
rect 5214 22660 5256 22700
rect 5296 22660 20048 22700
rect 20088 22660 20130 22700
rect 20170 22660 20212 22700
rect 20252 22660 20294 22700
rect 20334 22660 20376 22700
rect 20416 22660 20452 22700
rect 1152 22636 20452 22660
rect 5355 22532 5397 22541
rect 5355 22492 5356 22532
rect 5396 22492 5397 22532
rect 5355 22483 5397 22492
rect 5787 22532 5829 22541
rect 5787 22492 5788 22532
rect 5828 22492 5829 22532
rect 5787 22483 5829 22492
rect 8043 22532 8085 22541
rect 8043 22492 8044 22532
rect 8084 22492 8085 22532
rect 8043 22483 8085 22492
rect 10827 22532 10869 22541
rect 10827 22492 10828 22532
rect 10868 22492 10869 22532
rect 10827 22483 10869 22492
rect 14650 22532 14708 22533
rect 14650 22492 14659 22532
rect 14699 22492 14708 22532
rect 14650 22491 14708 22492
rect 16491 22532 16533 22541
rect 16491 22492 16492 22532
rect 16532 22492 16533 22532
rect 16491 22483 16533 22492
rect 18123 22532 18165 22541
rect 18123 22492 18124 22532
rect 18164 22492 18165 22532
rect 18123 22483 18165 22492
rect 18778 22532 18836 22533
rect 18778 22492 18787 22532
rect 18827 22492 18836 22532
rect 18778 22491 18836 22492
rect 19258 22532 19316 22533
rect 19258 22492 19267 22532
rect 19307 22492 19316 22532
rect 19258 22491 19316 22492
rect 19738 22532 19796 22533
rect 19738 22492 19747 22532
rect 19787 22492 19796 22532
rect 19738 22491 19796 22492
rect 20139 22532 20181 22541
rect 20139 22492 20140 22532
rect 20180 22492 20181 22532
rect 20139 22483 20181 22492
rect 3339 22448 3381 22457
rect 3339 22408 3340 22448
rect 3380 22408 3381 22448
rect 3339 22399 3381 22408
rect 8331 22448 8373 22457
rect 8331 22408 8332 22448
rect 8372 22408 8373 22448
rect 8331 22399 8373 22408
rect 8986 22448 9044 22449
rect 8986 22408 8995 22448
rect 9035 22408 9044 22448
rect 8986 22407 9044 22408
rect 13786 22448 13844 22449
rect 13786 22408 13795 22448
rect 13835 22408 13844 22448
rect 13786 22407 13844 22408
rect 14466 22439 14512 22448
rect 14466 22399 14467 22439
rect 14507 22399 14512 22439
rect 14466 22390 14512 22399
rect 1899 22364 1941 22373
rect 3610 22364 3668 22365
rect 1899 22324 1900 22364
rect 1940 22324 1941 22364
rect 1899 22315 1941 22324
rect 3147 22355 3189 22364
rect 3147 22315 3148 22355
rect 3188 22315 3189 22355
rect 3610 22324 3619 22364
rect 3659 22324 3668 22364
rect 3610 22323 3668 22324
rect 3723 22364 3765 22373
rect 3723 22324 3724 22364
rect 3764 22324 3765 22364
rect 3723 22315 3765 22324
rect 4107 22364 4149 22373
rect 6603 22364 6645 22373
rect 8218 22364 8276 22365
rect 4107 22324 4108 22364
rect 4148 22324 4149 22364
rect 4107 22315 4149 22324
rect 4683 22355 4725 22364
rect 4683 22315 4684 22355
rect 4724 22315 4725 22355
rect 3147 22306 3189 22315
rect 4683 22306 4725 22315
rect 5163 22355 5205 22364
rect 5163 22315 5164 22355
rect 5204 22315 5205 22355
rect 5163 22306 5205 22315
rect 6027 22355 6069 22364
rect 6027 22315 6028 22355
rect 6068 22315 6069 22355
rect 6258 22355 6304 22364
rect 6027 22306 6069 22315
rect 6126 22344 6168 22353
rect 6126 22304 6127 22344
rect 6167 22304 6168 22344
rect 6258 22315 6259 22355
rect 6299 22315 6304 22355
rect 6603 22324 6604 22364
rect 6644 22324 6645 22364
rect 6603 22315 6645 22324
rect 7851 22355 7893 22364
rect 7851 22315 7852 22355
rect 7892 22315 7893 22355
rect 8218 22324 8227 22364
rect 8267 22324 8276 22364
rect 8218 22323 8276 22324
rect 8534 22364 8576 22373
rect 8534 22324 8535 22364
rect 8575 22324 8576 22364
rect 8534 22315 8576 22324
rect 8662 22364 8704 22373
rect 8662 22324 8663 22364
rect 8703 22324 8704 22364
rect 8662 22315 8704 22324
rect 8907 22364 8949 22373
rect 8907 22324 8908 22364
rect 8948 22324 8949 22364
rect 8907 22315 8949 22324
rect 9387 22364 9429 22373
rect 11691 22364 11733 22373
rect 13707 22364 13749 22373
rect 9387 22324 9388 22364
rect 9428 22324 9429 22364
rect 9387 22315 9429 22324
rect 10635 22355 10677 22364
rect 10635 22315 10636 22355
rect 10676 22315 10677 22355
rect 11691 22324 11692 22364
rect 11732 22324 11733 22364
rect 11691 22315 11733 22324
rect 12939 22355 12981 22364
rect 12939 22315 12940 22355
rect 12980 22315 12981 22355
rect 13707 22324 13708 22364
rect 13748 22324 13749 22364
rect 13707 22315 13749 22324
rect 13882 22364 13940 22365
rect 13882 22324 13891 22364
rect 13931 22324 13940 22364
rect 13882 22323 13940 22324
rect 13995 22364 14037 22373
rect 13995 22324 13996 22364
rect 14036 22324 14037 22364
rect 13995 22315 14037 22324
rect 14170 22364 14228 22365
rect 14562 22364 14620 22365
rect 14170 22324 14179 22364
rect 14219 22324 14228 22364
rect 14170 22323 14228 22324
rect 14283 22355 14325 22364
rect 14283 22315 14284 22355
rect 14324 22315 14325 22355
rect 14562 22324 14571 22364
rect 14611 22324 14620 22364
rect 15051 22364 15093 22373
rect 16683 22364 16725 22373
rect 18466 22364 18524 22365
rect 14562 22323 14620 22324
rect 14688 22353 14730 22362
rect 6258 22306 6304 22315
rect 7851 22306 7893 22315
rect 10635 22306 10677 22315
rect 12939 22306 12981 22315
rect 14283 22306 14325 22315
rect 14688 22313 14689 22353
rect 14729 22313 14730 22353
rect 15051 22324 15052 22364
rect 15092 22324 15093 22364
rect 15051 22315 15093 22324
rect 16299 22355 16341 22364
rect 16299 22315 16300 22355
rect 16340 22315 16341 22355
rect 16683 22324 16684 22364
rect 16724 22324 16725 22364
rect 16683 22315 16725 22324
rect 17931 22355 17973 22364
rect 17931 22315 17932 22355
rect 17972 22315 17973 22355
rect 18466 22324 18475 22364
rect 18515 22324 18524 22364
rect 18466 22323 18524 22324
rect 18699 22364 18741 22373
rect 18699 22324 18700 22364
rect 18740 22324 18741 22364
rect 18699 22315 18741 22324
rect 18934 22364 18976 22373
rect 18934 22324 18935 22364
rect 18975 22324 18976 22364
rect 18934 22315 18976 22324
rect 19179 22364 19221 22373
rect 19179 22324 19180 22364
rect 19220 22324 19221 22364
rect 19546 22364 19604 22365
rect 19179 22315 19221 22324
rect 19419 22322 19461 22331
rect 19546 22324 19555 22364
rect 19595 22324 19604 22364
rect 19546 22323 19604 22324
rect 19659 22364 19701 22373
rect 19659 22324 19660 22364
rect 19700 22324 19701 22364
rect 14688 22304 14730 22313
rect 16299 22306 16341 22315
rect 17931 22306 17973 22315
rect 6126 22295 6168 22304
rect 1227 22280 1269 22289
rect 1227 22240 1228 22280
rect 1268 22240 1269 22280
rect 1227 22231 1269 22240
rect 4203 22280 4245 22289
rect 4203 22240 4204 22280
rect 4244 22240 4245 22280
rect 4203 22231 4245 22240
rect 5547 22280 5589 22289
rect 5547 22240 5548 22280
rect 5588 22240 5589 22280
rect 5547 22231 5589 22240
rect 8794 22280 8852 22281
rect 8794 22240 8803 22280
rect 8843 22240 8852 22280
rect 8794 22239 8852 22240
rect 11019 22280 11061 22289
rect 19419 22282 19420 22322
rect 19460 22282 19461 22322
rect 19659 22315 19701 22324
rect 19933 22364 19975 22373
rect 19933 22324 19934 22364
rect 19974 22324 19975 22364
rect 19933 22315 19975 22324
rect 20235 22355 20277 22364
rect 20235 22315 20236 22355
rect 20276 22315 20277 22355
rect 20235 22306 20277 22315
rect 11019 22240 11020 22280
rect 11060 22240 11061 22280
rect 11019 22231 11061 22240
rect 18586 22280 18644 22281
rect 18586 22240 18595 22280
rect 18635 22240 18644 22280
rect 18586 22239 18644 22240
rect 19066 22280 19124 22281
rect 19066 22240 19075 22280
rect 19115 22240 19124 22280
rect 19419 22273 19461 22282
rect 19066 22239 19124 22240
rect 6411 22196 6453 22205
rect 6411 22156 6412 22196
rect 6452 22156 6453 22196
rect 6411 22147 6453 22156
rect 13131 22196 13173 22205
rect 13131 22156 13132 22196
rect 13172 22156 13173 22196
rect 13131 22147 13173 22156
rect 1467 22112 1509 22121
rect 1467 22072 1468 22112
rect 1508 22072 1509 22112
rect 1467 22063 1509 22072
rect 8523 22112 8565 22121
rect 8523 22072 8524 22112
rect 8564 22072 8565 22112
rect 8523 22063 8565 22072
rect 11259 22112 11301 22121
rect 11259 22072 11260 22112
rect 11300 22072 11301 22112
rect 11259 22063 11301 22072
rect 19930 22112 19988 22113
rect 19930 22072 19939 22112
rect 19979 22072 19988 22112
rect 19930 22071 19988 22072
rect 1152 21944 20448 21968
rect 1152 21904 3688 21944
rect 3728 21904 3770 21944
rect 3810 21904 3852 21944
rect 3892 21904 3934 21944
rect 3974 21904 4016 21944
rect 4056 21904 18808 21944
rect 18848 21904 18890 21944
rect 18930 21904 18972 21944
rect 19012 21904 19054 21944
rect 19094 21904 19136 21944
rect 19176 21904 20448 21944
rect 1152 21880 20448 21904
rect 1851 21776 1893 21785
rect 1851 21736 1852 21776
rect 1892 21736 1893 21776
rect 1851 21727 1893 21736
rect 4347 21776 4389 21785
rect 4347 21736 4348 21776
rect 4388 21736 4389 21776
rect 4347 21727 4389 21736
rect 5259 21776 5301 21785
rect 5259 21736 5260 21776
rect 5300 21736 5301 21776
rect 5259 21727 5301 21736
rect 6891 21776 6933 21785
rect 6891 21736 6892 21776
rect 6932 21736 6933 21776
rect 6891 21727 6933 21736
rect 9003 21776 9045 21785
rect 9003 21736 9004 21776
rect 9044 21736 9045 21776
rect 9003 21727 9045 21736
rect 18123 21776 18165 21785
rect 18123 21736 18124 21776
rect 18164 21736 18165 21776
rect 18123 21727 18165 21736
rect 19371 21776 19413 21785
rect 19371 21736 19372 21776
rect 19412 21736 19413 21776
rect 19371 21727 19413 21736
rect 20331 21776 20373 21785
rect 20331 21736 20332 21776
rect 20372 21736 20373 21776
rect 20331 21727 20373 21736
rect 1227 21608 1269 21617
rect 1227 21568 1228 21608
rect 1268 21568 1269 21608
rect 1227 21559 1269 21568
rect 1611 21608 1653 21617
rect 1611 21568 1612 21608
rect 1652 21568 1653 21608
rect 1611 21559 1653 21568
rect 1995 21608 2037 21617
rect 1995 21568 1996 21608
rect 2036 21568 2037 21608
rect 1995 21559 2037 21568
rect 2955 21608 2997 21617
rect 2955 21568 2956 21608
rect 2996 21568 2997 21608
rect 2955 21559 2997 21568
rect 4587 21608 4629 21617
rect 15339 21608 15381 21617
rect 4587 21568 4588 21608
rect 4628 21568 4629 21608
rect 4587 21559 4629 21568
rect 14802 21599 14848 21608
rect 14802 21559 14803 21599
rect 14843 21559 14848 21599
rect 15339 21568 15340 21608
rect 15380 21568 15381 21608
rect 15339 21559 15381 21568
rect 15610 21608 15668 21609
rect 15610 21568 15619 21608
rect 15659 21568 15668 21608
rect 15610 21567 15668 21568
rect 14802 21550 14848 21559
rect 2458 21524 2516 21525
rect 2458 21484 2467 21524
rect 2507 21484 2516 21524
rect 2458 21483 2516 21484
rect 2571 21524 2613 21533
rect 2571 21484 2572 21524
rect 2612 21484 2613 21524
rect 2571 21475 2613 21484
rect 3051 21524 3093 21533
rect 3051 21484 3052 21524
rect 3092 21484 3093 21524
rect 3051 21475 3093 21484
rect 3523 21524 3581 21525
rect 3523 21484 3532 21524
rect 3572 21484 3581 21524
rect 3523 21483 3581 21484
rect 4011 21524 4069 21525
rect 4011 21484 4020 21524
rect 4060 21484 4069 21524
rect 4011 21483 4069 21484
rect 4234 21524 4292 21525
rect 4234 21484 4243 21524
rect 4283 21484 4292 21524
rect 4234 21483 4292 21484
rect 4954 21524 5012 21525
rect 4954 21484 4963 21524
rect 5003 21484 5012 21524
rect 4954 21483 5012 21484
rect 5259 21524 5301 21533
rect 5259 21484 5260 21524
rect 5300 21484 5301 21524
rect 5259 21475 5301 21484
rect 5451 21524 5493 21533
rect 5451 21484 5452 21524
rect 5492 21484 5493 21524
rect 5451 21475 5493 21484
rect 6691 21524 6749 21525
rect 6691 21484 6700 21524
rect 6740 21484 6749 21524
rect 6691 21483 6749 21484
rect 7371 21524 7413 21533
rect 7371 21484 7372 21524
rect 7412 21484 7413 21524
rect 7371 21475 7413 21484
rect 8611 21524 8669 21525
rect 8611 21484 8620 21524
rect 8660 21484 8669 21524
rect 8611 21483 8669 21484
rect 9187 21524 9245 21525
rect 9187 21484 9196 21524
rect 9236 21484 9245 21524
rect 9187 21483 9245 21484
rect 10403 21524 10445 21533
rect 10403 21484 10404 21524
rect 10444 21484 10445 21524
rect 10403 21475 10445 21484
rect 10819 21524 10877 21525
rect 10819 21484 10828 21524
rect 10868 21484 10877 21524
rect 10819 21483 10877 21484
rect 12075 21524 12117 21533
rect 12075 21484 12076 21524
rect 12116 21484 12117 21524
rect 12075 21475 12117 21484
rect 12459 21524 12501 21533
rect 12459 21484 12460 21524
rect 12500 21484 12501 21524
rect 12459 21475 12501 21484
rect 13699 21524 13757 21525
rect 13699 21484 13708 21524
rect 13748 21484 13757 21524
rect 13699 21483 13757 21484
rect 14091 21524 14133 21533
rect 14091 21484 14092 21524
rect 14132 21484 14133 21524
rect 14091 21475 14133 21484
rect 14225 21524 14283 21525
rect 14225 21484 14234 21524
rect 14274 21484 14283 21524
rect 14225 21483 14283 21484
rect 14666 21524 14708 21533
rect 14666 21484 14667 21524
rect 14707 21484 14708 21524
rect 14666 21475 14708 21484
rect 14907 21524 14949 21533
rect 14907 21484 14908 21524
rect 14948 21484 14949 21524
rect 14907 21475 14949 21484
rect 15012 21524 15054 21533
rect 15012 21484 15013 21524
rect 15053 21484 15054 21524
rect 15012 21475 15054 21484
rect 15130 21524 15188 21525
rect 15130 21484 15139 21524
rect 15179 21484 15188 21524
rect 15130 21483 15188 21484
rect 15243 21524 15285 21533
rect 15243 21484 15244 21524
rect 15284 21484 15285 21524
rect 15243 21475 15285 21484
rect 15478 21524 15520 21533
rect 15478 21484 15479 21524
rect 15519 21484 15520 21524
rect 15478 21475 15520 21484
rect 15723 21524 15765 21533
rect 15723 21484 15724 21524
rect 15764 21484 15765 21524
rect 15723 21475 15765 21484
rect 16291 21524 16349 21525
rect 16291 21484 16300 21524
rect 16340 21484 16349 21524
rect 16291 21483 16349 21484
rect 16683 21524 16725 21533
rect 16683 21484 16684 21524
rect 16724 21484 16725 21524
rect 16683 21475 16725 21484
rect 17923 21524 17981 21525
rect 17923 21484 17932 21524
rect 17972 21484 17981 21524
rect 17923 21483 17981 21484
rect 18411 21524 18453 21533
rect 18411 21484 18412 21524
rect 18452 21484 18453 21524
rect 18411 21475 18453 21484
rect 18699 21524 18741 21533
rect 18699 21484 18700 21524
rect 18740 21484 18741 21524
rect 18699 21475 18741 21484
rect 18970 21524 19028 21525
rect 18970 21484 18979 21524
rect 19019 21484 19028 21524
rect 18970 21483 19028 21484
rect 19659 21524 19701 21533
rect 19659 21484 19660 21524
rect 19700 21484 19701 21524
rect 19659 21475 19701 21484
rect 19906 21524 19964 21525
rect 19906 21484 19915 21524
rect 19955 21484 19964 21524
rect 19906 21483 19964 21484
rect 20026 21524 20084 21525
rect 20026 21484 20035 21524
rect 20075 21484 20084 21524
rect 20026 21483 20084 21484
rect 8811 21440 8853 21449
rect 8811 21400 8812 21440
rect 8852 21400 8853 21440
rect 8811 21391 8853 21400
rect 15802 21440 15860 21441
rect 15802 21400 15811 21440
rect 15851 21400 15860 21440
rect 15802 21399 15860 21400
rect 15997 21440 16039 21449
rect 15997 21400 15998 21440
rect 16038 21400 16039 21440
rect 15997 21391 16039 21400
rect 16203 21440 16245 21449
rect 16203 21400 16204 21440
rect 16244 21400 16245 21440
rect 16203 21391 16245 21400
rect 19083 21440 19125 21449
rect 19083 21400 19084 21440
rect 19124 21400 19125 21440
rect 19083 21391 19125 21400
rect 1467 21356 1509 21365
rect 1467 21316 1468 21356
rect 1508 21316 1509 21356
rect 1467 21307 1509 21316
rect 2235 21356 2277 21365
rect 2235 21316 2236 21356
rect 2276 21316 2277 21356
rect 2235 21307 2277 21316
rect 10635 21356 10677 21365
rect 10635 21316 10636 21356
rect 10676 21316 10677 21356
rect 10635 21307 10677 21316
rect 13899 21356 13941 21365
rect 13899 21316 13900 21356
rect 13940 21316 13941 21356
rect 13899 21307 13941 21316
rect 14379 21356 14421 21365
rect 14379 21316 14380 21356
rect 14420 21316 14421 21356
rect 14379 21307 14421 21316
rect 14571 21356 14613 21365
rect 14571 21316 14572 21356
rect 14612 21316 14613 21356
rect 14571 21307 14613 21316
rect 16090 21356 16148 21357
rect 16090 21316 16099 21356
rect 16139 21316 16148 21356
rect 16090 21315 16148 21316
rect 18267 21356 18309 21365
rect 18267 21316 18268 21356
rect 18308 21316 18309 21356
rect 18267 21307 18309 21316
rect 1152 21188 20452 21212
rect 1152 21148 4928 21188
rect 4968 21148 5010 21188
rect 5050 21148 5092 21188
rect 5132 21148 5174 21188
rect 5214 21148 5256 21188
rect 5296 21148 20048 21188
rect 20088 21148 20130 21188
rect 20170 21148 20212 21188
rect 20252 21148 20294 21188
rect 20334 21148 20376 21188
rect 20416 21148 20452 21188
rect 1152 21124 20452 21148
rect 2667 21020 2709 21029
rect 2667 20980 2668 21020
rect 2708 20980 2709 21020
rect 2667 20971 2709 20980
rect 3483 21020 3525 21029
rect 3483 20980 3484 21020
rect 3524 20980 3525 21020
rect 3483 20971 3525 20980
rect 5355 21020 5397 21029
rect 5355 20980 5356 21020
rect 5396 20980 5397 21020
rect 5355 20971 5397 20980
rect 9099 21020 9141 21029
rect 9099 20980 9100 21020
rect 9140 20980 9141 21020
rect 9099 20971 9141 20980
rect 15147 21020 15189 21029
rect 15147 20980 15148 21020
rect 15188 20980 15189 21020
rect 15147 20971 15189 20980
rect 20379 21020 20421 21029
rect 20379 20980 20380 21020
rect 20420 20980 20421 21020
rect 20379 20971 20421 20980
rect 7083 20936 7125 20945
rect 7083 20896 7084 20936
rect 7124 20896 7125 20936
rect 7083 20887 7125 20896
rect 13515 20936 13557 20945
rect 13515 20896 13516 20936
rect 13556 20896 13557 20936
rect 13515 20887 13557 20896
rect 16251 20936 16293 20945
rect 16251 20896 16252 20936
rect 16292 20896 16293 20936
rect 16251 20887 16293 20896
rect 1227 20852 1269 20861
rect 3915 20852 3957 20861
rect 5643 20852 5685 20861
rect 7354 20852 7412 20853
rect 1227 20812 1228 20852
rect 1268 20812 1269 20852
rect 1227 20803 1269 20812
rect 2475 20843 2517 20852
rect 2475 20803 2476 20843
rect 2516 20803 2517 20843
rect 3915 20812 3916 20852
rect 3956 20812 3957 20852
rect 3915 20803 3957 20812
rect 5163 20843 5205 20852
rect 5163 20803 5164 20843
rect 5204 20803 5205 20843
rect 5643 20812 5644 20852
rect 5684 20812 5685 20852
rect 5643 20803 5685 20812
rect 6891 20843 6933 20852
rect 6891 20803 6892 20843
rect 6932 20803 6933 20843
rect 7354 20812 7363 20852
rect 7403 20812 7412 20852
rect 7354 20811 7412 20812
rect 7467 20852 7509 20861
rect 7467 20812 7468 20852
rect 7508 20812 7509 20852
rect 7467 20803 7509 20812
rect 7851 20852 7893 20861
rect 9370 20852 9428 20853
rect 7851 20812 7852 20852
rect 7892 20812 7893 20852
rect 7851 20803 7893 20812
rect 8427 20843 8469 20852
rect 8427 20803 8428 20843
rect 8468 20803 8469 20843
rect 2475 20794 2517 20803
rect 5163 20794 5205 20803
rect 6891 20794 6933 20803
rect 8427 20794 8469 20803
rect 8907 20843 8949 20852
rect 8907 20803 8908 20843
rect 8948 20803 8949 20843
rect 9370 20812 9379 20852
rect 9419 20812 9428 20852
rect 9370 20811 9428 20812
rect 9483 20852 9525 20861
rect 9483 20812 9484 20852
rect 9524 20812 9525 20852
rect 9483 20803 9525 20812
rect 9867 20852 9909 20861
rect 12075 20852 12117 20861
rect 9867 20812 9868 20852
rect 9908 20812 9909 20852
rect 9867 20803 9909 20812
rect 10443 20843 10485 20852
rect 10443 20803 10444 20843
rect 10484 20803 10485 20843
rect 8907 20794 8949 20803
rect 10443 20794 10485 20803
rect 10923 20843 10965 20852
rect 10923 20803 10924 20843
rect 10964 20803 10965 20843
rect 12075 20812 12076 20852
rect 12116 20812 12117 20852
rect 12075 20803 12117 20812
rect 13707 20852 13749 20861
rect 13707 20812 13708 20852
rect 13748 20812 13749 20852
rect 13319 20810 13377 20811
rect 10923 20794 10965 20803
rect 2859 20768 2901 20777
rect 2859 20728 2860 20768
rect 2900 20728 2901 20768
rect 2859 20719 2901 20728
rect 3243 20768 3285 20777
rect 3243 20728 3244 20768
rect 3284 20728 3285 20768
rect 3243 20719 3285 20728
rect 7947 20768 7989 20777
rect 7947 20728 7948 20768
rect 7988 20728 7989 20768
rect 7947 20719 7989 20728
rect 9963 20768 10005 20777
rect 9963 20728 9964 20768
rect 10004 20728 10005 20768
rect 9963 20719 10005 20728
rect 11146 20768 11204 20769
rect 11146 20728 11155 20768
rect 11195 20728 11204 20768
rect 11146 20727 11204 20728
rect 11499 20768 11541 20777
rect 13319 20770 13328 20810
rect 13368 20770 13377 20810
rect 13707 20803 13749 20812
rect 15627 20852 15669 20861
rect 15627 20812 15628 20852
rect 15668 20812 15669 20852
rect 14951 20810 15009 20811
rect 13319 20769 13377 20770
rect 14951 20770 14960 20810
rect 15000 20770 15009 20810
rect 15627 20803 15669 20812
rect 15748 20852 15806 20853
rect 15748 20812 15757 20852
rect 15797 20812 15806 20852
rect 15748 20811 15806 20812
rect 16011 20852 16053 20861
rect 16011 20812 16012 20852
rect 16052 20812 16053 20852
rect 16011 20803 16053 20812
rect 16683 20852 16725 20861
rect 18507 20852 18549 20861
rect 16683 20812 16684 20852
rect 16724 20812 16725 20852
rect 16683 20803 16725 20812
rect 17931 20843 17973 20852
rect 17931 20803 17932 20843
rect 17972 20803 17973 20843
rect 18507 20812 18508 20852
rect 18548 20812 18549 20852
rect 18507 20803 18549 20812
rect 19755 20843 19797 20852
rect 19755 20803 19756 20843
rect 19796 20803 19797 20843
rect 17931 20794 17973 20803
rect 19755 20794 19797 20803
rect 14951 20769 15009 20770
rect 11499 20728 11500 20768
rect 11540 20728 11541 20768
rect 11499 20719 11541 20728
rect 16491 20768 16533 20777
rect 16491 20728 16492 20768
rect 16532 20728 16533 20768
rect 16491 20719 16533 20728
rect 20139 20768 20181 20777
rect 20139 20728 20140 20768
rect 20180 20728 20181 20768
rect 20139 20719 20181 20728
rect 18123 20684 18165 20693
rect 18123 20644 18124 20684
rect 18164 20644 18165 20684
rect 18123 20635 18165 20644
rect 3099 20600 3141 20609
rect 3099 20560 3100 20600
rect 3140 20560 3141 20600
rect 3099 20551 3141 20560
rect 11259 20600 11301 20609
rect 11259 20560 11260 20600
rect 11300 20560 11301 20600
rect 11259 20551 11301 20560
rect 15339 20600 15381 20609
rect 15339 20560 15340 20600
rect 15380 20560 15381 20600
rect 15339 20551 15381 20560
rect 19947 20600 19989 20609
rect 19947 20560 19948 20600
rect 19988 20560 19989 20600
rect 19947 20551 19989 20560
rect 1152 20432 20448 20456
rect 1152 20392 3688 20432
rect 3728 20392 3770 20432
rect 3810 20392 3852 20432
rect 3892 20392 3934 20432
rect 3974 20392 4016 20432
rect 4056 20392 18808 20432
rect 18848 20392 18890 20432
rect 18930 20392 18972 20432
rect 19012 20392 19054 20432
rect 19094 20392 19136 20432
rect 19176 20392 20448 20432
rect 1152 20368 20448 20392
rect 6603 20264 6645 20273
rect 6603 20224 6604 20264
rect 6644 20224 6645 20264
rect 6603 20215 6645 20224
rect 15915 20264 15957 20273
rect 15915 20224 15916 20264
rect 15956 20224 15957 20264
rect 15915 20215 15957 20224
rect 14043 20180 14085 20189
rect 14043 20140 14044 20180
rect 14084 20140 14085 20180
rect 14043 20131 14085 20140
rect 15435 20180 15477 20189
rect 15435 20140 15436 20180
rect 15476 20140 15477 20180
rect 15435 20131 15477 20140
rect 20187 20180 20229 20189
rect 20187 20140 20188 20180
rect 20228 20140 20229 20180
rect 20187 20131 20229 20140
rect 2859 20096 2901 20105
rect 2859 20056 2860 20096
rect 2900 20056 2901 20096
rect 2859 20047 2901 20056
rect 3099 20096 3141 20105
rect 3099 20056 3100 20096
rect 3140 20056 3141 20096
rect 3099 20047 3141 20056
rect 6987 20096 7029 20105
rect 6987 20056 6988 20096
rect 7028 20056 7029 20096
rect 6987 20047 7029 20056
rect 11115 20096 11157 20105
rect 11115 20056 11116 20096
rect 11156 20056 11157 20096
rect 11115 20047 11157 20056
rect 12394 20096 12452 20097
rect 12394 20056 12403 20096
rect 12443 20056 12452 20096
rect 12394 20055 12452 20056
rect 12747 20096 12789 20105
rect 12747 20056 12748 20096
rect 12788 20056 12789 20096
rect 12747 20047 12789 20056
rect 12939 20096 12981 20105
rect 12939 20056 12940 20096
rect 12980 20056 12981 20096
rect 12939 20047 12981 20056
rect 13179 20096 13221 20105
rect 13179 20056 13180 20096
rect 13220 20056 13221 20096
rect 13179 20047 13221 20056
rect 13803 20096 13845 20105
rect 13803 20056 13804 20096
rect 13844 20056 13845 20096
rect 13803 20047 13845 20056
rect 16395 20096 16437 20105
rect 16395 20056 16396 20096
rect 16436 20056 16437 20096
rect 16395 20047 16437 20056
rect 18795 20096 18837 20105
rect 18795 20056 18796 20096
rect 18836 20056 18837 20096
rect 18795 20047 18837 20056
rect 1227 20012 1269 20021
rect 1227 19972 1228 20012
rect 1268 19972 1269 20012
rect 1227 19963 1269 19972
rect 2475 20012 2533 20013
rect 2475 19972 2484 20012
rect 2524 19972 2533 20012
rect 2475 19971 2533 19972
rect 3531 20012 3573 20021
rect 3531 19972 3532 20012
rect 3572 19972 3573 20012
rect 3531 19963 3573 19972
rect 4771 20012 4829 20013
rect 4771 19972 4780 20012
rect 4820 19972 4829 20012
rect 4771 19971 4829 19972
rect 5163 20012 5205 20021
rect 5163 19972 5164 20012
rect 5204 19972 5205 20012
rect 5163 19963 5205 19972
rect 6403 20012 6461 20013
rect 6403 19972 6412 20012
rect 6452 19972 6461 20012
rect 6403 19971 6461 19972
rect 7275 20012 7317 20021
rect 7275 19972 7276 20012
rect 7316 19972 7317 20012
rect 7275 19963 7317 19972
rect 8515 20012 8573 20013
rect 8515 19972 8524 20012
rect 8564 19972 8573 20012
rect 8515 19971 8573 19972
rect 8907 20012 8949 20021
rect 8907 19972 8908 20012
rect 8948 19972 8949 20012
rect 8907 19963 8949 19972
rect 10147 20012 10205 20013
rect 10147 19972 10156 20012
rect 10196 19972 10205 20012
rect 10147 19971 10205 19972
rect 10618 20012 10676 20013
rect 10618 19972 10627 20012
rect 10667 19972 10676 20012
rect 10618 19971 10676 19972
rect 10731 20012 10773 20021
rect 10731 19972 10732 20012
rect 10772 19972 10773 20012
rect 10731 19963 10773 19972
rect 11211 20012 11253 20021
rect 11211 19972 11212 20012
rect 11252 19972 11253 20012
rect 11211 19963 11253 19972
rect 11683 20012 11741 20013
rect 11683 19972 11692 20012
rect 11732 19972 11741 20012
rect 11683 19971 11741 19972
rect 12171 20012 12229 20013
rect 12171 19972 12180 20012
rect 12220 19972 12229 20012
rect 12171 19971 12229 19972
rect 13515 20012 13557 20021
rect 13515 19972 13516 20012
rect 13556 19972 13557 20012
rect 13515 19963 13557 19972
rect 13659 20012 13701 20021
rect 13659 19972 13660 20012
rect 13700 19972 13701 20012
rect 13659 19963 13701 19972
rect 14134 20012 14176 20021
rect 14134 19972 14135 20012
rect 14175 19972 14176 20012
rect 14134 19963 14176 19972
rect 14266 20012 14324 20013
rect 14266 19972 14275 20012
rect 14315 19972 14324 20012
rect 14266 19971 14324 19972
rect 14379 20012 14421 20021
rect 14379 19972 14380 20012
rect 14420 19972 14421 20012
rect 14379 19963 14421 19972
rect 14763 20012 14805 20021
rect 14763 19972 14764 20012
rect 14804 19972 14805 20012
rect 14763 19963 14805 19972
rect 15034 20012 15092 20013
rect 15034 19972 15043 20012
rect 15083 19972 15092 20012
rect 15034 19971 15092 19972
rect 15610 20012 15668 20013
rect 15610 19972 15619 20012
rect 15659 19972 15668 20012
rect 15610 19971 15668 19972
rect 15929 20012 15971 20021
rect 15929 19972 15930 20012
rect 15970 19972 15971 20012
rect 15929 19963 15971 19972
rect 16587 20012 16629 20021
rect 16587 19972 16588 20012
rect 16628 19972 16629 20012
rect 16587 19963 16629 19972
rect 17827 20012 17885 20013
rect 17827 19972 17836 20012
rect 17876 19972 17885 20012
rect 17827 19971 17885 19972
rect 18298 20012 18356 20013
rect 18298 19972 18307 20012
rect 18347 19972 18356 20012
rect 18298 19971 18356 19972
rect 18411 20012 18453 20021
rect 18411 19972 18412 20012
rect 18452 19972 18453 20012
rect 18411 19963 18453 19972
rect 18891 20012 18933 20021
rect 18891 19972 18892 20012
rect 18932 19972 18933 20012
rect 18891 19963 18933 19972
rect 19362 20012 19420 20013
rect 19362 19972 19371 20012
rect 19411 19972 19420 20012
rect 19362 19971 19420 19972
rect 19882 20012 19940 20013
rect 19882 19972 19891 20012
rect 19931 19972 19940 20012
rect 19882 19971 19940 19972
rect 20331 20012 20373 20021
rect 20331 19972 20332 20012
rect 20372 19972 20373 20012
rect 20331 19963 20373 19972
rect 8715 19928 8757 19937
rect 8715 19888 8716 19928
rect 8756 19888 8757 19928
rect 8715 19879 8757 19888
rect 10347 19928 10389 19937
rect 10347 19888 10348 19928
rect 10388 19888 10389 19928
rect 10347 19879 10389 19888
rect 15147 19928 15189 19937
rect 15147 19888 15148 19928
rect 15188 19888 15189 19928
rect 15147 19879 15189 19888
rect 18027 19928 18069 19937
rect 18027 19888 18028 19928
rect 18068 19888 18069 19928
rect 18027 19879 18069 19888
rect 2667 19844 2709 19853
rect 2667 19804 2668 19844
rect 2708 19804 2709 19844
rect 2667 19795 2709 19804
rect 4971 19844 5013 19853
rect 4971 19804 4972 19844
rect 5012 19804 5013 19844
rect 4971 19795 5013 19804
rect 6747 19844 6789 19853
rect 6747 19804 6748 19844
rect 6788 19804 6789 19844
rect 6747 19795 6789 19804
rect 12507 19844 12549 19853
rect 12507 19804 12508 19844
rect 12548 19804 12549 19844
rect 12507 19795 12549 19804
rect 14458 19844 14516 19845
rect 14458 19804 14467 19844
rect 14507 19804 14516 19844
rect 14458 19803 14516 19804
rect 15706 19844 15764 19845
rect 15706 19804 15715 19844
rect 15755 19804 15764 19844
rect 15706 19803 15764 19804
rect 16155 19844 16197 19853
rect 16155 19804 16156 19844
rect 16196 19804 16197 19844
rect 16155 19795 16197 19804
rect 20043 19844 20085 19853
rect 20043 19804 20044 19844
rect 20084 19804 20085 19844
rect 20043 19795 20085 19804
rect 1152 19676 20452 19700
rect 1152 19636 4928 19676
rect 4968 19636 5010 19676
rect 5050 19636 5092 19676
rect 5132 19636 5174 19676
rect 5214 19636 5256 19676
rect 5296 19636 20048 19676
rect 20088 19636 20130 19676
rect 20170 19636 20212 19676
rect 20252 19636 20294 19676
rect 20334 19636 20376 19676
rect 20416 19636 20452 19676
rect 1152 19612 20452 19636
rect 4779 19508 4821 19517
rect 4779 19468 4780 19508
rect 4820 19468 4821 19508
rect 4779 19459 4821 19468
rect 7371 19508 7413 19517
rect 7371 19468 7372 19508
rect 7412 19468 7413 19508
rect 7371 19459 7413 19468
rect 7899 19508 7941 19517
rect 7899 19468 7900 19508
rect 7940 19468 7941 19508
rect 7899 19459 7941 19468
rect 8667 19508 8709 19517
rect 8667 19468 8668 19508
rect 8708 19468 8709 19508
rect 8667 19459 8709 19468
rect 10107 19508 10149 19517
rect 10107 19468 10108 19508
rect 10148 19468 10149 19508
rect 10107 19459 10149 19468
rect 12267 19508 12309 19517
rect 12267 19468 12268 19508
rect 12308 19468 12309 19508
rect 12267 19459 12309 19468
rect 14235 19508 14277 19517
rect 14235 19468 14236 19508
rect 14276 19468 14277 19508
rect 14235 19459 14277 19468
rect 14667 19508 14709 19517
rect 14667 19468 14668 19508
rect 14708 19468 14709 19508
rect 14667 19459 14709 19468
rect 15243 19508 15285 19517
rect 15243 19468 15244 19508
rect 15284 19468 15285 19508
rect 15243 19459 15285 19468
rect 15963 19508 16005 19517
rect 15963 19468 15964 19508
rect 16004 19468 16005 19508
rect 15963 19459 16005 19468
rect 20139 19508 20181 19517
rect 20139 19468 20140 19508
rect 20180 19468 20181 19508
rect 20139 19459 20181 19468
rect 2763 19424 2805 19433
rect 2763 19384 2764 19424
rect 2804 19384 2805 19424
rect 2763 19375 2805 19384
rect 15147 19424 15189 19433
rect 15147 19384 15148 19424
rect 15188 19384 15189 19424
rect 15147 19375 15189 19384
rect 17931 19424 17973 19433
rect 17931 19384 17932 19424
rect 17972 19384 17973 19424
rect 17931 19375 17973 19384
rect 1323 19340 1365 19349
rect 3034 19340 3092 19341
rect 1323 19300 1324 19340
rect 1364 19300 1365 19340
rect 1323 19291 1365 19300
rect 2571 19331 2613 19340
rect 2571 19291 2572 19331
rect 2612 19291 2613 19331
rect 3034 19300 3043 19340
rect 3083 19300 3092 19340
rect 3034 19299 3092 19300
rect 3147 19340 3189 19349
rect 3147 19300 3148 19340
rect 3188 19300 3189 19340
rect 3147 19291 3189 19300
rect 3531 19340 3573 19349
rect 5626 19340 5684 19341
rect 3531 19300 3532 19340
rect 3572 19300 3573 19340
rect 3531 19291 3573 19300
rect 4107 19331 4149 19340
rect 4107 19291 4108 19331
rect 4148 19291 4149 19331
rect 2571 19282 2613 19291
rect 4107 19282 4149 19291
rect 4587 19331 4629 19340
rect 4587 19291 4588 19331
rect 4628 19291 4629 19331
rect 5626 19300 5635 19340
rect 5675 19300 5684 19340
rect 5626 19299 5684 19300
rect 5739 19340 5781 19349
rect 10827 19340 10869 19349
rect 13995 19340 14037 19349
rect 5739 19300 5740 19340
rect 5780 19300 5781 19340
rect 5739 19291 5781 19300
rect 6699 19331 6741 19340
rect 6699 19291 6700 19331
rect 6740 19291 6741 19331
rect 4587 19282 4629 19291
rect 6699 19282 6741 19291
rect 7179 19331 7221 19340
rect 7179 19291 7180 19331
rect 7220 19291 7221 19331
rect 10827 19300 10828 19340
rect 10868 19300 10869 19340
rect 10827 19291 10869 19300
rect 12075 19331 12117 19340
rect 12075 19291 12076 19331
rect 12116 19291 12117 19331
rect 13995 19300 13996 19340
rect 14036 19300 14037 19340
rect 13995 19291 14037 19300
rect 14379 19340 14421 19349
rect 14379 19300 14380 19340
rect 14420 19300 14421 19340
rect 14379 19291 14421 19300
rect 14571 19340 14613 19349
rect 14571 19300 14572 19340
rect 14612 19300 14613 19340
rect 14571 19291 14613 19300
rect 14746 19340 14804 19341
rect 14746 19300 14755 19340
rect 14795 19300 14804 19340
rect 14746 19299 14804 19300
rect 15034 19340 15092 19341
rect 15034 19300 15043 19340
rect 15083 19300 15092 19340
rect 15034 19299 15092 19300
rect 15353 19340 15395 19349
rect 15353 19300 15354 19340
rect 15394 19300 15395 19340
rect 15353 19291 15395 19300
rect 16491 19340 16533 19349
rect 18394 19340 18452 19341
rect 16491 19300 16492 19340
rect 16532 19300 16533 19340
rect 16491 19291 16533 19300
rect 17739 19331 17781 19340
rect 17739 19291 17740 19331
rect 17780 19291 17781 19331
rect 18394 19300 18403 19340
rect 18443 19300 18452 19340
rect 18394 19299 18452 19300
rect 18507 19340 18549 19349
rect 18507 19300 18508 19340
rect 18548 19300 18549 19340
rect 18507 19291 18549 19300
rect 18891 19340 18933 19349
rect 18891 19300 18892 19340
rect 18932 19300 18933 19340
rect 18891 19291 18933 19300
rect 19467 19331 19509 19340
rect 19467 19291 19468 19331
rect 19508 19291 19509 19331
rect 7179 19282 7221 19291
rect 12075 19282 12117 19291
rect 17739 19282 17781 19291
rect 19467 19282 19509 19291
rect 19947 19331 19989 19340
rect 19947 19291 19948 19331
rect 19988 19291 19989 19331
rect 19947 19282 19989 19291
rect 3627 19256 3669 19265
rect 3627 19216 3628 19256
rect 3668 19216 3669 19256
rect 3627 19207 3669 19216
rect 4971 19256 5013 19265
rect 4971 19216 4972 19256
rect 5012 19216 5013 19256
rect 4971 19207 5013 19216
rect 6123 19256 6165 19265
rect 6123 19216 6124 19256
rect 6164 19216 6165 19256
rect 6123 19207 6165 19216
rect 6250 19256 6308 19257
rect 6250 19216 6259 19256
rect 6299 19216 6308 19256
rect 6250 19215 6308 19216
rect 7755 19256 7797 19265
rect 7755 19216 7756 19256
rect 7796 19216 7797 19256
rect 7755 19207 7797 19216
rect 8139 19256 8181 19265
rect 8139 19216 8140 19256
rect 8180 19216 8181 19256
rect 8139 19207 8181 19216
rect 8523 19256 8565 19265
rect 8523 19216 8524 19256
rect 8564 19216 8565 19256
rect 8523 19207 8565 19216
rect 8907 19256 8949 19265
rect 8907 19216 8908 19256
rect 8948 19216 8949 19256
rect 8907 19207 8949 19216
rect 9099 19256 9141 19265
rect 9099 19216 9100 19256
rect 9140 19216 9141 19256
rect 9099 19207 9141 19216
rect 9675 19256 9717 19265
rect 9675 19216 9676 19256
rect 9716 19216 9717 19256
rect 9675 19207 9717 19216
rect 9867 19256 9909 19265
rect 9867 19216 9868 19256
rect 9908 19216 9909 19256
rect 9867 19207 9909 19216
rect 10443 19256 10485 19265
rect 10443 19216 10444 19256
rect 10484 19216 10485 19256
rect 10443 19207 10485 19216
rect 15675 19256 15717 19265
rect 15675 19216 15676 19256
rect 15716 19216 15717 19256
rect 15675 19207 15717 19216
rect 16299 19256 16341 19265
rect 16299 19216 16300 19256
rect 16340 19216 16341 19256
rect 16299 19207 16341 19216
rect 18987 19256 19029 19265
rect 18987 19216 18988 19256
rect 19028 19216 19029 19256
rect 18987 19207 19029 19216
rect 9339 19172 9381 19181
rect 9339 19132 9340 19172
rect 9380 19132 9381 19172
rect 9339 19123 9381 19132
rect 14139 19172 14181 19181
rect 14139 19132 14140 19172
rect 14180 19132 14181 19172
rect 14139 19123 14181 19132
rect 5211 19088 5253 19097
rect 5211 19048 5212 19088
rect 5252 19048 5253 19088
rect 5211 19039 5253 19048
rect 7515 19088 7557 19097
rect 7515 19048 7516 19088
rect 7556 19048 7557 19088
rect 7515 19039 7557 19048
rect 8283 19088 8325 19097
rect 8283 19048 8284 19088
rect 8324 19048 8325 19088
rect 8283 19039 8325 19048
rect 9435 19088 9477 19097
rect 9435 19048 9436 19088
rect 9476 19048 9477 19088
rect 9435 19039 9477 19048
rect 10203 19088 10245 19097
rect 10203 19048 10204 19088
rect 10244 19048 10245 19088
rect 10203 19039 10245 19048
rect 16059 19088 16101 19097
rect 16059 19048 16060 19088
rect 16100 19048 16101 19088
rect 16059 19039 16101 19048
rect 1152 18920 20448 18944
rect 1152 18880 3688 18920
rect 3728 18880 3770 18920
rect 3810 18880 3852 18920
rect 3892 18880 3934 18920
rect 3974 18880 4016 18920
rect 4056 18880 18808 18920
rect 18848 18880 18890 18920
rect 18930 18880 18972 18920
rect 19012 18880 19054 18920
rect 19094 18880 19136 18920
rect 19176 18880 20448 18920
rect 1152 18856 20448 18880
rect 1467 18752 1509 18761
rect 1467 18712 1468 18752
rect 1508 18712 1509 18752
rect 1467 18703 1509 18712
rect 19947 18752 19989 18761
rect 19947 18712 19948 18752
rect 19988 18712 19989 18752
rect 19947 18703 19989 18712
rect 18123 18668 18165 18677
rect 18123 18628 18124 18668
rect 18164 18628 18165 18668
rect 18123 18619 18165 18628
rect 20379 18668 20421 18677
rect 20379 18628 20380 18668
rect 20420 18628 20421 18668
rect 20379 18619 20421 18628
rect 1227 18584 1269 18593
rect 1227 18544 1228 18584
rect 1268 18544 1269 18584
rect 1227 18535 1269 18544
rect 1611 18584 1653 18593
rect 1611 18544 1612 18584
rect 1652 18544 1653 18584
rect 1611 18535 1653 18544
rect 1995 18584 2037 18593
rect 1995 18544 1996 18584
rect 2036 18544 2037 18584
rect 1995 18535 2037 18544
rect 2955 18584 2997 18593
rect 2955 18544 2956 18584
rect 2996 18544 2997 18584
rect 2955 18535 2997 18544
rect 4234 18584 4292 18585
rect 4234 18544 4243 18584
rect 4283 18544 4292 18584
rect 4234 18543 4292 18544
rect 4587 18584 4629 18593
rect 4587 18544 4588 18584
rect 4628 18544 4629 18584
rect 4587 18535 4629 18544
rect 4779 18584 4821 18593
rect 4779 18544 4780 18584
rect 4820 18544 4821 18584
rect 4779 18535 4821 18544
rect 5163 18584 5205 18593
rect 5163 18544 5164 18584
rect 5204 18544 5205 18584
rect 5163 18535 5205 18544
rect 5403 18584 5445 18593
rect 5403 18544 5404 18584
rect 5444 18544 5445 18584
rect 5403 18535 5445 18544
rect 8043 18584 8085 18593
rect 8043 18544 8044 18584
rect 8084 18544 8085 18584
rect 8043 18535 8085 18544
rect 9322 18584 9380 18585
rect 9322 18544 9331 18584
rect 9371 18544 9380 18584
rect 9322 18543 9380 18544
rect 9675 18584 9717 18593
rect 9675 18544 9676 18584
rect 9716 18544 9717 18584
rect 9675 18535 9717 18544
rect 12939 18584 12981 18593
rect 12939 18544 12940 18584
rect 12980 18544 12981 18584
rect 12939 18535 12981 18544
rect 17739 18584 17781 18593
rect 17739 18544 17740 18584
rect 17780 18544 17781 18584
rect 17739 18535 17781 18544
rect 20139 18584 20181 18593
rect 20139 18544 20140 18584
rect 20180 18544 20181 18584
rect 20139 18535 20181 18544
rect 2445 18500 2487 18509
rect 2445 18460 2446 18500
rect 2486 18460 2487 18500
rect 2445 18451 2487 18460
rect 2571 18500 2613 18509
rect 2571 18460 2572 18500
rect 2612 18460 2613 18500
rect 2571 18451 2613 18460
rect 3051 18500 3093 18509
rect 3051 18460 3052 18500
rect 3092 18460 3093 18500
rect 3051 18451 3093 18460
rect 3523 18500 3581 18501
rect 3523 18460 3532 18500
rect 3572 18460 3581 18500
rect 3523 18459 3581 18460
rect 4011 18500 4069 18501
rect 4011 18460 4020 18500
rect 4060 18460 4069 18500
rect 4011 18459 4069 18460
rect 5739 18500 5781 18509
rect 5739 18460 5740 18500
rect 5780 18460 5781 18500
rect 5739 18451 5781 18460
rect 6979 18500 7037 18501
rect 6979 18460 6988 18500
rect 7028 18460 7037 18500
rect 6979 18459 7037 18460
rect 7546 18500 7604 18501
rect 7546 18460 7555 18500
rect 7595 18460 7604 18500
rect 7546 18459 7604 18460
rect 7659 18500 7701 18509
rect 7659 18460 7660 18500
rect 7700 18460 7701 18500
rect 7659 18451 7701 18460
rect 8139 18500 8181 18509
rect 8139 18460 8140 18500
rect 8180 18460 8181 18500
rect 8139 18451 8181 18460
rect 8614 18500 8672 18501
rect 8614 18460 8623 18500
rect 8663 18460 8672 18500
rect 8614 18459 8672 18460
rect 9099 18500 9157 18501
rect 9099 18460 9108 18500
rect 9148 18460 9157 18500
rect 9099 18459 9157 18460
rect 10731 18500 10773 18509
rect 10731 18460 10732 18500
rect 10772 18460 10773 18500
rect 10731 18451 10773 18460
rect 11971 18500 12029 18501
rect 11971 18460 11980 18500
rect 12020 18460 12029 18500
rect 11971 18459 12029 18460
rect 12442 18500 12500 18501
rect 12442 18460 12451 18500
rect 12491 18460 12500 18500
rect 12442 18459 12500 18460
rect 12555 18500 12597 18509
rect 12555 18460 12556 18500
rect 12596 18460 12597 18500
rect 12555 18451 12597 18460
rect 13035 18500 13077 18509
rect 13035 18460 13036 18500
rect 13076 18460 13077 18500
rect 13035 18451 13077 18460
rect 13507 18500 13565 18501
rect 13507 18460 13516 18500
rect 13556 18460 13565 18500
rect 13507 18459 13565 18460
rect 13995 18500 14053 18501
rect 13995 18460 14004 18500
rect 14044 18460 14053 18500
rect 13995 18459 14053 18460
rect 14379 18500 14421 18509
rect 14379 18460 14380 18500
rect 14420 18460 14421 18500
rect 14379 18451 14421 18460
rect 15619 18500 15677 18501
rect 15619 18460 15628 18500
rect 15668 18460 15677 18500
rect 15619 18459 15677 18460
rect 16011 18500 16053 18509
rect 16011 18460 16012 18500
rect 16052 18460 16053 18500
rect 16011 18451 16053 18460
rect 17251 18500 17309 18501
rect 17251 18460 17260 18500
rect 17300 18460 17309 18500
rect 17251 18459 17309 18460
rect 18123 18500 18165 18509
rect 18123 18460 18124 18500
rect 18164 18460 18165 18500
rect 18123 18451 18165 18460
rect 18315 18500 18357 18509
rect 18315 18460 18316 18500
rect 18356 18460 18357 18500
rect 18315 18451 18357 18460
rect 18507 18500 18549 18509
rect 18507 18460 18508 18500
rect 18548 18460 18549 18500
rect 18507 18451 18549 18460
rect 19747 18500 19805 18501
rect 19747 18460 19756 18500
rect 19796 18460 19805 18500
rect 19747 18459 19805 18460
rect 1851 18416 1893 18425
rect 1851 18376 1852 18416
rect 1892 18376 1893 18416
rect 1851 18367 1893 18376
rect 4347 18416 4389 18425
rect 4347 18376 4348 18416
rect 4388 18376 4389 18416
rect 4347 18367 4389 18376
rect 5019 18416 5061 18425
rect 5019 18376 5020 18416
rect 5060 18376 5061 18416
rect 5019 18367 5061 18376
rect 7179 18416 7221 18425
rect 7179 18376 7180 18416
rect 7220 18376 7221 18416
rect 7179 18367 7221 18376
rect 12171 18416 12213 18425
rect 12171 18376 12172 18416
rect 12212 18376 12213 18416
rect 12171 18367 12213 18376
rect 2235 18332 2277 18341
rect 2235 18292 2236 18332
rect 2276 18292 2277 18332
rect 2235 18283 2277 18292
rect 9435 18332 9477 18341
rect 9435 18292 9436 18332
rect 9476 18292 9477 18332
rect 9435 18283 9477 18292
rect 14187 18332 14229 18341
rect 14187 18292 14188 18332
rect 14228 18292 14229 18332
rect 14187 18283 14229 18292
rect 15819 18332 15861 18341
rect 15819 18292 15820 18332
rect 15860 18292 15861 18332
rect 15819 18283 15861 18292
rect 17451 18332 17493 18341
rect 17451 18292 17452 18332
rect 17492 18292 17493 18332
rect 17451 18283 17493 18292
rect 17979 18332 18021 18341
rect 17979 18292 17980 18332
rect 18020 18292 18021 18332
rect 17979 18283 18021 18292
rect 1152 18164 20452 18188
rect 1152 18124 4928 18164
rect 4968 18124 5010 18164
rect 5050 18124 5092 18164
rect 5132 18124 5174 18164
rect 5214 18124 5256 18164
rect 5296 18124 20048 18164
rect 20088 18124 20130 18164
rect 20170 18124 20212 18164
rect 20252 18124 20294 18164
rect 20334 18124 20376 18164
rect 20416 18124 20452 18164
rect 1152 18100 20452 18124
rect 1467 17996 1509 18005
rect 1467 17956 1468 17996
rect 1508 17956 1509 17996
rect 1467 17947 1509 17956
rect 3051 17996 3093 18005
rect 3051 17956 3052 17996
rect 3092 17956 3093 17996
rect 3051 17947 3093 17956
rect 5163 17996 5205 18005
rect 5163 17956 5164 17996
rect 5204 17956 5205 17996
rect 5163 17947 5205 17956
rect 8139 17996 8181 18005
rect 8139 17956 8140 17996
rect 8180 17956 8181 17996
rect 8139 17947 8181 17956
rect 13323 17996 13365 18005
rect 13323 17956 13324 17996
rect 13364 17956 13365 17996
rect 13323 17947 13365 17956
rect 20379 17996 20421 18005
rect 20379 17956 20380 17996
rect 20420 17956 20421 17996
rect 20379 17947 20421 17956
rect 5691 17912 5733 17921
rect 5691 17872 5692 17912
rect 5732 17872 5733 17912
rect 5691 17863 5733 17872
rect 1611 17828 1653 17837
rect 3418 17828 3476 17829
rect 1611 17788 1612 17828
rect 1652 17788 1653 17828
rect 1611 17779 1653 17788
rect 2859 17819 2901 17828
rect 2859 17779 2860 17819
rect 2900 17779 2901 17819
rect 3418 17788 3427 17828
rect 3467 17788 3476 17828
rect 3418 17787 3476 17788
rect 3531 17828 3573 17837
rect 3531 17788 3532 17828
rect 3572 17788 3573 17828
rect 3531 17779 3573 17788
rect 3915 17828 3957 17837
rect 6699 17828 6741 17837
rect 8410 17828 8468 17829
rect 3915 17788 3916 17828
rect 3956 17788 3957 17828
rect 3915 17779 3957 17788
rect 4491 17819 4533 17828
rect 4491 17779 4492 17819
rect 4532 17779 4533 17819
rect 2859 17770 2901 17779
rect 4491 17770 4533 17779
rect 4971 17819 5013 17828
rect 4971 17779 4972 17819
rect 5012 17779 5013 17819
rect 6699 17788 6700 17828
rect 6740 17788 6741 17828
rect 6699 17779 6741 17788
rect 7947 17819 7989 17828
rect 7947 17779 7948 17819
rect 7988 17779 7989 17819
rect 8410 17788 8419 17828
rect 8459 17788 8468 17828
rect 8410 17787 8468 17788
rect 8523 17828 8565 17837
rect 8523 17788 8524 17828
rect 8564 17788 8565 17828
rect 8523 17779 8565 17788
rect 8907 17828 8949 17837
rect 11883 17828 11925 17837
rect 15130 17828 15188 17829
rect 8907 17788 8908 17828
rect 8948 17788 8949 17828
rect 8907 17779 8949 17788
rect 9483 17819 9525 17828
rect 9483 17779 9484 17819
rect 9524 17779 9525 17819
rect 4971 17770 5013 17779
rect 7947 17770 7989 17779
rect 9483 17770 9525 17779
rect 9963 17819 10005 17828
rect 9963 17779 9964 17819
rect 10004 17779 10005 17819
rect 11883 17788 11884 17828
rect 11924 17788 11925 17828
rect 11883 17779 11925 17788
rect 13131 17819 13173 17828
rect 13131 17779 13132 17819
rect 13172 17779 13173 17819
rect 15130 17788 15139 17828
rect 15179 17788 15188 17828
rect 15130 17787 15188 17788
rect 15243 17828 15285 17837
rect 15243 17788 15244 17828
rect 15284 17788 15285 17828
rect 15243 17779 15285 17788
rect 15723 17828 15765 17837
rect 17530 17828 17588 17829
rect 15723 17788 15724 17828
rect 15764 17788 15765 17828
rect 15723 17779 15765 17788
rect 16203 17819 16245 17828
rect 16203 17779 16204 17819
rect 16244 17779 16245 17819
rect 9963 17770 10005 17779
rect 13131 17770 13173 17779
rect 16203 17770 16245 17779
rect 16683 17819 16725 17828
rect 16683 17779 16684 17819
rect 16724 17779 16725 17819
rect 17530 17788 17539 17828
rect 17579 17788 17588 17828
rect 17530 17787 17588 17788
rect 17643 17828 17685 17837
rect 17643 17788 17644 17828
rect 17684 17788 17685 17828
rect 17643 17779 17685 17788
rect 18027 17828 18069 17837
rect 18027 17788 18028 17828
rect 18068 17788 18069 17828
rect 18027 17779 18069 17788
rect 18603 17819 18645 17828
rect 18603 17779 18604 17819
rect 18644 17779 18645 17819
rect 16683 17770 16725 17779
rect 18603 17770 18645 17779
rect 19083 17819 19125 17828
rect 19083 17779 19084 17819
rect 19124 17779 19125 17819
rect 19083 17770 19125 17779
rect 1227 17744 1269 17753
rect 1227 17704 1228 17744
rect 1268 17704 1269 17744
rect 1227 17695 1269 17704
rect 4011 17744 4053 17753
rect 4011 17704 4012 17744
rect 4052 17704 4053 17744
rect 4011 17695 4053 17704
rect 5355 17744 5397 17753
rect 5355 17704 5356 17744
rect 5396 17704 5397 17744
rect 5355 17695 5397 17704
rect 5931 17744 5973 17753
rect 5931 17704 5932 17744
rect 5972 17704 5973 17744
rect 5931 17695 5973 17704
rect 6123 17744 6165 17753
rect 6123 17704 6124 17744
rect 6164 17704 6165 17744
rect 6123 17695 6165 17704
rect 9003 17744 9045 17753
rect 9003 17704 9004 17744
rect 9044 17704 9045 17744
rect 9003 17695 9045 17704
rect 10186 17744 10244 17745
rect 10186 17704 10195 17744
rect 10235 17704 10244 17744
rect 10186 17703 10244 17704
rect 10635 17744 10677 17753
rect 10635 17704 10636 17744
rect 10676 17704 10677 17744
rect 10635 17695 10677 17704
rect 14379 17744 14421 17753
rect 14379 17704 14380 17744
rect 14420 17704 14421 17744
rect 14379 17695 14421 17704
rect 14859 17744 14901 17753
rect 14859 17704 14860 17744
rect 14900 17704 14901 17744
rect 14859 17695 14901 17704
rect 15627 17744 15669 17753
rect 15627 17704 15628 17744
rect 15668 17704 15669 17744
rect 15627 17695 15669 17704
rect 16906 17744 16964 17745
rect 16906 17704 16915 17744
rect 16955 17704 16964 17744
rect 16906 17703 16964 17704
rect 17259 17744 17301 17753
rect 17259 17704 17260 17744
rect 17300 17704 17301 17744
rect 17259 17695 17301 17704
rect 18123 17744 18165 17753
rect 18123 17704 18124 17744
rect 18164 17704 18165 17744
rect 18123 17695 18165 17704
rect 19659 17744 19701 17753
rect 19659 17704 19660 17744
rect 19700 17704 19701 17744
rect 19659 17695 19701 17704
rect 20139 17744 20181 17753
rect 20139 17704 20140 17744
rect 20180 17704 20181 17744
rect 20139 17695 20181 17704
rect 5595 17576 5637 17585
rect 5595 17536 5596 17576
rect 5636 17536 5637 17576
rect 5595 17527 5637 17536
rect 6363 17576 6405 17585
rect 6363 17536 6364 17576
rect 6404 17536 6405 17576
rect 6363 17527 6405 17536
rect 10395 17576 10437 17585
rect 10395 17536 10396 17576
rect 10436 17536 10437 17576
rect 10395 17527 10437 17536
rect 14139 17576 14181 17585
rect 14139 17536 14140 17576
rect 14180 17536 14181 17576
rect 14139 17527 14181 17536
rect 14619 17576 14661 17585
rect 14619 17536 14620 17576
rect 14660 17536 14661 17576
rect 14619 17527 14661 17536
rect 17019 17576 17061 17585
rect 17019 17536 17020 17576
rect 17060 17536 17061 17576
rect 17019 17527 17061 17536
rect 19306 17576 19364 17577
rect 19306 17536 19315 17576
rect 19355 17536 19364 17576
rect 19306 17535 19364 17536
rect 19419 17576 19461 17585
rect 19419 17536 19420 17576
rect 19460 17536 19461 17576
rect 19419 17527 19461 17536
rect 1152 17408 20448 17432
rect 1152 17368 3688 17408
rect 3728 17368 3770 17408
rect 3810 17368 3852 17408
rect 3892 17368 3934 17408
rect 3974 17368 4016 17408
rect 4056 17368 18808 17408
rect 18848 17368 18890 17408
rect 18930 17368 18972 17408
rect 19012 17368 19054 17408
rect 19094 17368 19136 17408
rect 19176 17368 20448 17408
rect 1152 17344 20448 17368
rect 6507 17240 6549 17249
rect 6507 17200 6508 17240
rect 6548 17200 6549 17240
rect 6507 17191 6549 17200
rect 8139 17240 8181 17249
rect 8139 17200 8140 17240
rect 8180 17200 8181 17240
rect 8139 17191 8181 17200
rect 16971 17240 17013 17249
rect 16971 17200 16972 17240
rect 17012 17200 17013 17240
rect 16971 17191 17013 17200
rect 17307 17240 17349 17249
rect 17307 17200 17308 17240
rect 17348 17200 17349 17240
rect 17307 17191 17349 17200
rect 19179 17240 19221 17249
rect 19179 17200 19180 17240
rect 19220 17200 19221 17240
rect 19179 17191 19221 17200
rect 19611 17240 19653 17249
rect 19611 17200 19612 17240
rect 19652 17200 19653 17240
rect 19611 17191 19653 17200
rect 20379 17240 20421 17249
rect 20379 17200 20380 17240
rect 20420 17200 20421 17240
rect 20379 17191 20421 17200
rect 2667 17156 2709 17165
rect 2667 17116 2668 17156
rect 2708 17116 2709 17156
rect 2667 17107 2709 17116
rect 8283 17156 8325 17165
rect 8283 17116 8284 17156
rect 8324 17116 8325 17156
rect 8283 17107 8325 17116
rect 19995 17156 20037 17165
rect 19995 17116 19996 17156
rect 20036 17116 20037 17156
rect 19995 17107 20037 17116
rect 3531 17072 3573 17081
rect 3531 17032 3532 17072
rect 3572 17032 3573 17072
rect 3531 17023 3573 17032
rect 8523 17072 8565 17081
rect 8523 17032 8524 17072
rect 8564 17032 8565 17072
rect 8523 17023 8565 17032
rect 9483 17072 9525 17081
rect 9483 17032 9484 17072
rect 9524 17032 9525 17072
rect 9483 17023 9525 17032
rect 10762 17072 10820 17073
rect 10762 17032 10771 17072
rect 10811 17032 10820 17072
rect 10762 17031 10820 17032
rect 11115 17072 11157 17081
rect 11115 17032 11116 17072
rect 11156 17032 11157 17072
rect 11115 17023 11157 17032
rect 14091 17072 14133 17081
rect 14091 17032 14092 17072
rect 14132 17032 14133 17072
rect 14091 17023 14133 17032
rect 17547 17072 17589 17081
rect 17547 17032 17548 17072
rect 17588 17032 17589 17072
rect 17547 17023 17589 17032
rect 19371 17072 19413 17081
rect 19371 17032 19372 17072
rect 19412 17032 19413 17072
rect 19371 17023 19413 17032
rect 19755 17072 19797 17081
rect 19755 17032 19756 17072
rect 19796 17032 19797 17072
rect 19755 17023 19797 17032
rect 20139 17072 20181 17081
rect 20139 17032 20140 17072
rect 20180 17032 20181 17072
rect 20139 17023 20181 17032
rect 1227 16988 1269 16997
rect 1227 16948 1228 16988
rect 1268 16948 1269 16988
rect 1227 16939 1269 16948
rect 2467 16988 2525 16989
rect 2467 16948 2476 16988
rect 2516 16948 2525 16988
rect 2467 16947 2525 16948
rect 3034 16988 3092 16989
rect 3034 16948 3043 16988
rect 3083 16948 3092 16988
rect 3034 16947 3092 16948
rect 3147 16988 3189 16997
rect 3147 16948 3148 16988
rect 3188 16948 3189 16988
rect 3147 16939 3189 16948
rect 3627 16988 3669 16997
rect 3627 16948 3628 16988
rect 3668 16948 3669 16988
rect 3627 16939 3669 16948
rect 4099 16988 4157 16989
rect 4099 16948 4108 16988
rect 4148 16948 4157 16988
rect 4099 16947 4157 16948
rect 4587 16988 4645 16989
rect 4587 16948 4596 16988
rect 4636 16948 4645 16988
rect 4587 16947 4645 16948
rect 5067 16988 5109 16997
rect 5067 16948 5068 16988
rect 5108 16948 5109 16988
rect 5067 16939 5109 16948
rect 6307 16988 6365 16989
rect 6307 16948 6316 16988
rect 6356 16948 6365 16988
rect 6307 16947 6365 16948
rect 6699 16988 6741 16997
rect 6699 16948 6700 16988
rect 6740 16948 6741 16988
rect 6699 16939 6741 16948
rect 7939 16988 7997 16989
rect 7939 16948 7948 16988
rect 7988 16948 7997 16988
rect 7939 16947 7997 16948
rect 8986 16988 9044 16989
rect 8986 16948 8995 16988
rect 9035 16948 9044 16988
rect 8986 16947 9044 16948
rect 9099 16988 9141 16997
rect 9099 16948 9100 16988
rect 9140 16948 9141 16988
rect 9099 16939 9141 16948
rect 9579 16988 9621 16997
rect 9579 16948 9580 16988
rect 9620 16948 9621 16988
rect 9579 16939 9621 16948
rect 10051 16988 10109 16989
rect 10051 16948 10060 16988
rect 10100 16948 10109 16988
rect 10051 16947 10109 16948
rect 10570 16988 10628 16989
rect 10570 16948 10579 16988
rect 10619 16948 10628 16988
rect 10570 16947 10628 16948
rect 11499 16988 11541 16997
rect 11499 16948 11500 16988
rect 11540 16948 11541 16988
rect 11499 16939 11541 16948
rect 12739 16988 12797 16989
rect 12739 16948 12748 16988
rect 12788 16948 12797 16988
rect 12739 16947 12797 16948
rect 13594 16988 13652 16989
rect 13594 16948 13603 16988
rect 13643 16948 13652 16988
rect 13594 16947 13652 16948
rect 13707 16988 13749 16997
rect 13707 16948 13708 16988
rect 13748 16948 13749 16988
rect 13707 16939 13749 16948
rect 14187 16988 14229 16997
rect 14187 16948 14188 16988
rect 14228 16948 14229 16988
rect 14187 16939 14229 16948
rect 14659 16988 14717 16989
rect 14659 16948 14668 16988
rect 14708 16948 14717 16988
rect 14659 16947 14717 16948
rect 15178 16988 15236 16989
rect 15178 16948 15187 16988
rect 15227 16948 15236 16988
rect 15178 16947 15236 16948
rect 15531 16988 15573 16997
rect 15531 16948 15532 16988
rect 15572 16948 15573 16988
rect 15531 16939 15573 16948
rect 16771 16988 16829 16989
rect 16771 16948 16780 16988
rect 16820 16948 16829 16988
rect 16771 16947 16829 16948
rect 17739 16988 17781 16997
rect 17739 16948 17740 16988
rect 17780 16948 17781 16988
rect 17739 16939 17781 16948
rect 18979 16988 19037 16989
rect 18979 16948 18988 16988
rect 19028 16948 19037 16988
rect 18979 16947 19037 16948
rect 12939 16904 12981 16913
rect 12939 16864 12940 16904
rect 12980 16864 12981 16904
rect 12939 16855 12981 16864
rect 4779 16820 4821 16829
rect 4779 16780 4780 16820
rect 4820 16780 4821 16820
rect 4779 16771 4821 16780
rect 10875 16820 10917 16829
rect 10875 16780 10876 16820
rect 10916 16780 10917 16820
rect 10875 16771 10917 16780
rect 15339 16820 15381 16829
rect 15339 16780 15340 16820
rect 15380 16780 15381 16820
rect 15339 16771 15381 16780
rect 1152 16652 20452 16676
rect 1152 16612 4928 16652
rect 4968 16612 5010 16652
rect 5050 16612 5092 16652
rect 5132 16612 5174 16652
rect 5214 16612 5256 16652
rect 5296 16612 20048 16652
rect 20088 16612 20130 16652
rect 20170 16612 20212 16652
rect 20252 16612 20294 16652
rect 20334 16612 20376 16652
rect 20416 16612 20452 16652
rect 1152 16588 20452 16612
rect 1467 16484 1509 16493
rect 1467 16444 1468 16484
rect 1508 16444 1509 16484
rect 1467 16435 1509 16444
rect 5451 16484 5493 16493
rect 5451 16444 5452 16484
rect 5492 16444 5493 16484
rect 5451 16435 5493 16444
rect 7131 16484 7173 16493
rect 7131 16444 7132 16484
rect 7172 16444 7173 16484
rect 7131 16435 7173 16444
rect 8907 16484 8949 16493
rect 8907 16444 8908 16484
rect 8948 16444 8949 16484
rect 8907 16435 8949 16444
rect 10635 16484 10677 16493
rect 10635 16444 10636 16484
rect 10676 16444 10677 16484
rect 10635 16435 10677 16444
rect 15051 16484 15093 16493
rect 15051 16444 15052 16484
rect 15092 16444 15093 16484
rect 15051 16435 15093 16444
rect 15243 16484 15285 16493
rect 15243 16444 15244 16484
rect 15284 16444 15285 16484
rect 15243 16435 15285 16444
rect 17115 16484 17157 16493
rect 17115 16444 17116 16484
rect 17156 16444 17157 16484
rect 17115 16435 17157 16444
rect 17883 16484 17925 16493
rect 17883 16444 17884 16484
rect 17924 16444 17925 16484
rect 17883 16435 17925 16444
rect 20139 16484 20181 16493
rect 20139 16444 20140 16484
rect 20180 16444 20181 16484
rect 20139 16435 20181 16444
rect 12651 16400 12693 16409
rect 12651 16360 12652 16400
rect 12692 16360 12693 16400
rect 12651 16351 12693 16360
rect 1707 16316 1749 16325
rect 3706 16316 3764 16317
rect 1707 16276 1708 16316
rect 1748 16276 1749 16316
rect 1707 16267 1749 16276
rect 2955 16307 2997 16316
rect 2955 16267 2956 16307
rect 2996 16267 2997 16307
rect 3706 16276 3715 16316
rect 3755 16276 3764 16316
rect 3706 16275 3764 16276
rect 3819 16316 3861 16325
rect 3819 16276 3820 16316
rect 3860 16276 3861 16316
rect 3819 16267 3861 16276
rect 4203 16316 4245 16325
rect 7467 16316 7509 16325
rect 9195 16316 9237 16325
rect 11211 16316 11253 16325
rect 13306 16316 13364 16317
rect 4203 16276 4204 16316
rect 4244 16276 4245 16316
rect 4203 16267 4245 16276
rect 4779 16307 4821 16316
rect 4779 16267 4780 16307
rect 4820 16267 4821 16307
rect 2955 16258 2997 16267
rect 4779 16258 4821 16267
rect 5259 16307 5301 16316
rect 5259 16267 5260 16307
rect 5300 16267 5301 16307
rect 7467 16276 7468 16316
rect 7508 16276 7509 16316
rect 7467 16267 7509 16276
rect 8715 16307 8757 16316
rect 8715 16267 8716 16307
rect 8756 16267 8757 16307
rect 9195 16276 9196 16316
rect 9236 16276 9237 16316
rect 9195 16267 9237 16276
rect 10443 16307 10485 16316
rect 10443 16267 10444 16307
rect 10484 16267 10485 16307
rect 11211 16276 11212 16316
rect 11252 16276 11253 16316
rect 11211 16267 11253 16276
rect 12459 16307 12501 16316
rect 12459 16267 12460 16307
rect 12500 16267 12501 16307
rect 13306 16276 13315 16316
rect 13355 16276 13364 16316
rect 13306 16275 13364 16276
rect 13419 16316 13461 16325
rect 13419 16276 13420 16316
rect 13460 16276 13461 16316
rect 13419 16267 13461 16276
rect 13803 16316 13845 16325
rect 16683 16316 16725 16325
rect 13803 16276 13804 16316
rect 13844 16276 13845 16316
rect 13803 16267 13845 16276
rect 14379 16307 14421 16316
rect 14379 16267 14380 16307
rect 14420 16267 14421 16307
rect 5259 16258 5301 16267
rect 8715 16258 8757 16267
rect 10443 16258 10485 16267
rect 12459 16258 12501 16267
rect 14379 16258 14421 16267
rect 14859 16307 14901 16316
rect 14859 16267 14860 16307
rect 14900 16267 14901 16307
rect 14859 16258 14901 16267
rect 15435 16307 15477 16316
rect 15435 16267 15436 16307
rect 15476 16267 15477 16307
rect 16683 16276 16684 16316
rect 16724 16276 16725 16316
rect 16683 16267 16725 16276
rect 18394 16316 18452 16317
rect 18394 16276 18403 16316
rect 18443 16276 18452 16316
rect 18394 16275 18452 16276
rect 18507 16316 18549 16325
rect 18507 16276 18508 16316
rect 18548 16276 18549 16316
rect 18507 16267 18549 16276
rect 18891 16316 18933 16325
rect 18891 16276 18892 16316
rect 18932 16276 18933 16316
rect 18891 16267 18933 16276
rect 19467 16307 19509 16316
rect 19467 16267 19468 16307
rect 19508 16267 19509 16307
rect 15435 16258 15477 16267
rect 19467 16258 19509 16267
rect 19947 16307 19989 16316
rect 19947 16267 19948 16307
rect 19988 16267 19989 16307
rect 19947 16258 19989 16267
rect 1227 16232 1269 16241
rect 1227 16192 1228 16232
rect 1268 16192 1269 16232
rect 1227 16183 1269 16192
rect 4299 16232 4341 16241
rect 4299 16192 4300 16232
rect 4340 16192 4341 16232
rect 4299 16183 4341 16192
rect 5835 16232 5877 16241
rect 5835 16192 5836 16232
rect 5876 16192 5877 16232
rect 5835 16183 5877 16192
rect 6219 16232 6261 16241
rect 6219 16192 6220 16232
rect 6260 16192 6261 16232
rect 6219 16183 6261 16192
rect 6411 16232 6453 16241
rect 6411 16192 6412 16232
rect 6452 16192 6453 16232
rect 6411 16183 6453 16192
rect 6891 16232 6933 16241
rect 6891 16192 6892 16232
rect 6932 16192 6933 16232
rect 6891 16183 6933 16192
rect 10827 16232 10869 16241
rect 10827 16192 10828 16232
rect 10868 16192 10869 16232
rect 10827 16183 10869 16192
rect 13899 16232 13941 16241
rect 13899 16192 13900 16232
rect 13940 16192 13941 16232
rect 13899 16183 13941 16192
rect 17355 16232 17397 16241
rect 17355 16192 17356 16232
rect 17396 16192 17397 16232
rect 17355 16183 17397 16192
rect 17739 16232 17781 16241
rect 17739 16192 17740 16232
rect 17780 16192 17781 16232
rect 17739 16183 17781 16192
rect 18123 16232 18165 16241
rect 18123 16192 18124 16232
rect 18164 16192 18165 16232
rect 18123 16183 18165 16192
rect 18987 16232 19029 16241
rect 18987 16192 18988 16232
rect 19028 16192 19029 16232
rect 18987 16183 19029 16192
rect 3147 16148 3189 16157
rect 3147 16108 3148 16148
rect 3188 16108 3189 16148
rect 3147 16099 3189 16108
rect 17499 16148 17541 16157
rect 17499 16108 17500 16148
rect 17540 16108 17541 16148
rect 17499 16099 17541 16108
rect 5595 16064 5637 16073
rect 5595 16024 5596 16064
rect 5636 16024 5637 16064
rect 5595 16015 5637 16024
rect 5979 16064 6021 16073
rect 5979 16024 5980 16064
rect 6020 16024 6021 16064
rect 5979 16015 6021 16024
rect 6651 16064 6693 16073
rect 6651 16024 6652 16064
rect 6692 16024 6693 16064
rect 6651 16015 6693 16024
rect 11067 16064 11109 16073
rect 11067 16024 11068 16064
rect 11108 16024 11109 16064
rect 11067 16015 11109 16024
rect 15082 16064 15140 16065
rect 15082 16024 15091 16064
rect 15131 16024 15140 16064
rect 15082 16023 15140 16024
rect 1152 15896 20448 15920
rect 1152 15856 3688 15896
rect 3728 15856 3770 15896
rect 3810 15856 3852 15896
rect 3892 15856 3934 15896
rect 3974 15856 4016 15896
rect 4056 15856 18808 15896
rect 18848 15856 18890 15896
rect 18930 15856 18972 15896
rect 19012 15856 19054 15896
rect 19094 15856 19136 15896
rect 19176 15856 20448 15896
rect 1152 15832 20448 15856
rect 2763 15728 2805 15737
rect 2763 15688 2764 15728
rect 2804 15688 2805 15728
rect 2763 15679 2805 15688
rect 4683 15728 4725 15737
rect 4683 15688 4684 15728
rect 4724 15688 4725 15728
rect 4683 15679 4725 15688
rect 6651 15728 6693 15737
rect 6651 15688 6652 15728
rect 6692 15688 6693 15728
rect 6651 15679 6693 15688
rect 10731 15728 10773 15737
rect 10731 15688 10732 15728
rect 10772 15688 10773 15728
rect 10731 15679 10773 15688
rect 14571 15728 14613 15737
rect 14571 15688 14572 15728
rect 14612 15688 14613 15728
rect 14571 15679 14613 15688
rect 18123 15728 18165 15737
rect 18123 15688 18124 15728
rect 18164 15688 18165 15728
rect 18123 15679 18165 15688
rect 4491 15644 4533 15653
rect 4491 15604 4492 15644
rect 4532 15604 4533 15644
rect 4491 15595 4533 15604
rect 12459 15644 12501 15653
rect 12459 15604 12460 15644
rect 12500 15604 12501 15644
rect 12459 15595 12501 15604
rect 6507 15560 6549 15569
rect 6507 15520 6508 15560
rect 6548 15520 6549 15560
rect 6507 15511 6549 15520
rect 6891 15560 6933 15569
rect 6891 15520 6892 15560
rect 6932 15520 6933 15560
rect 6891 15511 6933 15520
rect 7179 15560 7221 15569
rect 7179 15520 7180 15560
rect 7220 15520 7221 15560
rect 7179 15511 7221 15520
rect 12651 15560 12693 15569
rect 12651 15520 12652 15560
rect 12692 15520 12693 15560
rect 12651 15511 12693 15520
rect 18891 15560 18933 15569
rect 18891 15520 18892 15560
rect 18932 15520 18933 15560
rect 18891 15511 18933 15520
rect 1323 15476 1365 15485
rect 1323 15436 1324 15476
rect 1364 15436 1365 15476
rect 1323 15427 1365 15436
rect 2563 15476 2621 15477
rect 2563 15436 2572 15476
rect 2612 15436 2621 15476
rect 2563 15435 2621 15436
rect 3051 15476 3093 15485
rect 3051 15436 3052 15476
rect 3092 15436 3093 15476
rect 3051 15427 3093 15436
rect 4291 15476 4349 15477
rect 4291 15436 4300 15476
rect 4340 15436 4349 15476
rect 4291 15435 4349 15436
rect 4867 15476 4925 15477
rect 4867 15436 4876 15476
rect 4916 15436 4925 15476
rect 4867 15435 4925 15436
rect 6123 15476 6165 15485
rect 6123 15436 6124 15476
rect 6164 15436 6165 15476
rect 6123 15427 6165 15436
rect 7659 15476 7701 15485
rect 7659 15436 7660 15476
rect 7700 15436 7701 15476
rect 7659 15427 7701 15436
rect 8899 15476 8957 15477
rect 8899 15436 8908 15476
rect 8948 15436 8957 15476
rect 8899 15435 8957 15436
rect 9291 15476 9333 15485
rect 9291 15436 9292 15476
rect 9332 15436 9333 15476
rect 9291 15427 9333 15436
rect 10531 15476 10589 15477
rect 10531 15436 10540 15476
rect 10580 15436 10589 15476
rect 10531 15435 10589 15436
rect 11019 15476 11061 15485
rect 11019 15436 11020 15476
rect 11060 15436 11061 15476
rect 11019 15427 11061 15436
rect 12259 15476 12317 15477
rect 12259 15436 12268 15476
rect 12308 15436 12317 15476
rect 12259 15435 12317 15436
rect 13131 15476 13173 15485
rect 13131 15436 13132 15476
rect 13172 15436 13173 15476
rect 13131 15427 13173 15436
rect 14371 15476 14429 15477
rect 14371 15436 14380 15476
rect 14420 15436 14429 15476
rect 14371 15435 14429 15436
rect 15051 15476 15093 15485
rect 15051 15436 15052 15476
rect 15092 15436 15093 15476
rect 15051 15427 15093 15436
rect 16291 15476 16349 15477
rect 16291 15436 16300 15476
rect 16340 15436 16349 15476
rect 16291 15435 16349 15436
rect 16683 15476 16725 15485
rect 16683 15436 16684 15476
rect 16724 15436 16725 15476
rect 16683 15427 16725 15436
rect 17923 15476 17981 15477
rect 17923 15436 17932 15476
rect 17972 15436 17981 15476
rect 17923 15435 17981 15436
rect 18394 15476 18452 15477
rect 18394 15436 18403 15476
rect 18443 15436 18452 15476
rect 18394 15435 18452 15436
rect 18507 15476 18549 15485
rect 18507 15436 18508 15476
rect 18548 15436 18549 15476
rect 18507 15427 18549 15436
rect 18987 15476 19029 15485
rect 18987 15436 18988 15476
rect 19028 15436 19029 15476
rect 18987 15427 19029 15436
rect 19459 15476 19517 15477
rect 19459 15436 19468 15476
rect 19508 15436 19517 15476
rect 19459 15435 19517 15436
rect 19978 15476 20036 15477
rect 19978 15436 19987 15476
rect 20027 15436 20036 15476
rect 19978 15435 20036 15436
rect 12891 15392 12933 15401
rect 12891 15352 12892 15392
rect 12932 15352 12933 15392
rect 12891 15343 12933 15352
rect 6267 15308 6309 15317
rect 6267 15268 6268 15308
rect 6308 15268 6309 15308
rect 6267 15259 6309 15268
rect 7419 15308 7461 15317
rect 7419 15268 7420 15308
rect 7460 15268 7461 15308
rect 7419 15259 7461 15268
rect 9099 15308 9141 15317
rect 9099 15268 9100 15308
rect 9140 15268 9141 15308
rect 9099 15259 9141 15268
rect 16491 15308 16533 15317
rect 16491 15268 16492 15308
rect 16532 15268 16533 15308
rect 16491 15259 16533 15268
rect 20139 15308 20181 15317
rect 20139 15268 20140 15308
rect 20180 15268 20181 15308
rect 20139 15259 20181 15268
rect 1152 15140 20452 15164
rect 1152 15100 4928 15140
rect 4968 15100 5010 15140
rect 5050 15100 5092 15140
rect 5132 15100 5174 15140
rect 5214 15100 5256 15140
rect 5296 15100 20048 15140
rect 20088 15100 20130 15140
rect 20170 15100 20212 15140
rect 20252 15100 20294 15140
rect 20334 15100 20376 15140
rect 20416 15100 20452 15140
rect 1152 15076 20452 15100
rect 2859 14972 2901 14981
rect 2859 14932 2860 14972
rect 2900 14932 2901 14972
rect 2859 14923 2901 14932
rect 14571 14972 14613 14981
rect 14571 14932 14572 14972
rect 14612 14932 14613 14972
rect 14571 14923 14613 14932
rect 15291 14972 15333 14981
rect 15291 14932 15292 14972
rect 15332 14932 15333 14972
rect 15291 14923 15333 14932
rect 18267 14972 18309 14981
rect 18267 14932 18268 14972
rect 18308 14932 18309 14972
rect 18267 14923 18309 14932
rect 20139 14972 20181 14981
rect 20139 14932 20140 14972
rect 20180 14932 20181 14972
rect 20139 14923 20181 14932
rect 7755 14888 7797 14897
rect 7755 14848 7756 14888
rect 7796 14848 7797 14888
rect 7755 14839 7797 14848
rect 16090 14888 16148 14889
rect 16090 14848 16099 14888
rect 16139 14848 16148 14888
rect 16090 14847 16148 14848
rect 17852 14824 17894 14833
rect 1419 14804 1461 14813
rect 3051 14804 3093 14813
rect 4683 14804 4725 14813
rect 6315 14804 6357 14813
rect 8410 14804 8468 14805
rect 1419 14764 1420 14804
rect 1460 14764 1461 14804
rect 1419 14755 1461 14764
rect 2667 14795 2709 14804
rect 2667 14755 2668 14795
rect 2708 14755 2709 14795
rect 3051 14764 3052 14804
rect 3092 14764 3093 14804
rect 3051 14755 3093 14764
rect 4299 14795 4341 14804
rect 4299 14755 4300 14795
rect 4340 14755 4341 14795
rect 4683 14764 4684 14804
rect 4724 14764 4725 14804
rect 4683 14755 4725 14764
rect 5931 14795 5973 14804
rect 5931 14755 5932 14795
rect 5972 14755 5973 14795
rect 6315 14764 6316 14804
rect 6356 14764 6357 14804
rect 6315 14755 6357 14764
rect 7563 14795 7605 14804
rect 7563 14755 7564 14795
rect 7604 14755 7605 14795
rect 8410 14764 8419 14804
rect 8459 14764 8468 14804
rect 8410 14763 8468 14764
rect 8523 14804 8565 14813
rect 8523 14764 8524 14804
rect 8564 14764 8565 14804
rect 8523 14755 8565 14764
rect 8907 14804 8949 14813
rect 11019 14804 11061 14813
rect 12826 14804 12884 14805
rect 8907 14764 8908 14804
rect 8948 14764 8949 14804
rect 8907 14755 8949 14764
rect 9483 14795 9525 14804
rect 9483 14755 9484 14795
rect 9524 14755 9525 14795
rect 2667 14746 2709 14755
rect 4299 14746 4341 14755
rect 5931 14746 5973 14755
rect 7563 14746 7605 14755
rect 9483 14746 9525 14755
rect 9963 14795 10005 14804
rect 9963 14755 9964 14795
rect 10004 14755 10005 14795
rect 11019 14764 11020 14804
rect 11060 14764 11061 14804
rect 11019 14755 11061 14764
rect 12267 14795 12309 14804
rect 12267 14755 12268 14795
rect 12308 14755 12309 14795
rect 12826 14764 12835 14804
rect 12875 14764 12884 14804
rect 12826 14763 12884 14764
rect 12939 14804 12981 14813
rect 12939 14764 12940 14804
rect 12980 14764 12981 14804
rect 12939 14755 12981 14764
rect 13323 14804 13365 14813
rect 16282 14804 16340 14805
rect 17259 14804 17301 14813
rect 13323 14764 13324 14804
rect 13364 14764 13365 14804
rect 13323 14755 13365 14764
rect 13899 14795 13941 14804
rect 13899 14755 13900 14795
rect 13940 14755 13941 14795
rect 9963 14746 10005 14755
rect 12267 14746 12309 14755
rect 13899 14746 13941 14755
rect 14379 14795 14421 14804
rect 14379 14755 14380 14795
rect 14420 14755 14421 14795
rect 16282 14764 16291 14804
rect 16331 14764 16340 14804
rect 16282 14763 16340 14764
rect 16779 14795 16821 14804
rect 14379 14746 14421 14755
rect 16779 14755 16780 14795
rect 16820 14755 16821 14795
rect 17259 14764 17260 14804
rect 17300 14764 17301 14804
rect 17259 14755 17301 14764
rect 17739 14804 17781 14813
rect 17739 14764 17740 14804
rect 17780 14764 17781 14804
rect 17852 14784 17853 14824
rect 17893 14784 17894 14824
rect 17852 14775 17894 14784
rect 18699 14804 18741 14813
rect 17739 14755 17781 14764
rect 18699 14764 18700 14804
rect 18740 14764 18741 14804
rect 18699 14755 18741 14764
rect 19947 14795 19989 14804
rect 19947 14755 19948 14795
rect 19988 14755 19989 14795
rect 16779 14746 16821 14755
rect 19947 14746 19989 14755
rect 8139 14720 8181 14729
rect 8139 14680 8140 14720
rect 8180 14680 8181 14720
rect 8139 14671 8181 14680
rect 9003 14720 9045 14729
rect 9003 14680 9004 14720
rect 9044 14680 9045 14720
rect 9003 14671 9045 14680
rect 10635 14720 10677 14729
rect 10635 14680 10636 14720
rect 10676 14680 10677 14720
rect 10635 14671 10677 14680
rect 13419 14720 13461 14729
rect 13419 14680 13420 14720
rect 13460 14680 13461 14720
rect 13419 14671 13461 14680
rect 15531 14720 15573 14729
rect 15531 14680 15532 14720
rect 15572 14680 15573 14720
rect 15531 14671 15573 14680
rect 15915 14720 15957 14729
rect 15915 14680 15916 14720
rect 15956 14680 15957 14720
rect 15915 14671 15957 14680
rect 17355 14720 17397 14729
rect 17355 14680 17356 14720
rect 17396 14680 17397 14720
rect 17355 14671 17397 14680
rect 18507 14720 18549 14729
rect 18507 14680 18508 14720
rect 18548 14680 18549 14720
rect 18507 14671 18549 14680
rect 10203 14636 10245 14645
rect 10203 14596 10204 14636
rect 10244 14596 10245 14636
rect 10203 14587 10245 14596
rect 10875 14636 10917 14645
rect 10875 14596 10876 14636
rect 10916 14596 10917 14636
rect 10875 14587 10917 14596
rect 4491 14552 4533 14561
rect 4491 14512 4492 14552
rect 4532 14512 4533 14552
rect 4491 14503 4533 14512
rect 6123 14552 6165 14561
rect 6123 14512 6124 14552
rect 6164 14512 6165 14552
rect 6123 14503 6165 14512
rect 7899 14552 7941 14561
rect 7899 14512 7900 14552
rect 7940 14512 7941 14552
rect 7899 14503 7941 14512
rect 12459 14552 12501 14561
rect 12459 14512 12460 14552
rect 12500 14512 12501 14552
rect 12459 14503 12501 14512
rect 15675 14552 15717 14561
rect 15675 14512 15676 14552
rect 15716 14512 15717 14552
rect 15675 14503 15717 14512
rect 1152 14384 20448 14408
rect 1152 14344 3688 14384
rect 3728 14344 3770 14384
rect 3810 14344 3852 14384
rect 3892 14344 3934 14384
rect 3974 14344 4016 14384
rect 4056 14344 18808 14384
rect 18848 14344 18890 14384
rect 18930 14344 18972 14384
rect 19012 14344 19054 14384
rect 19094 14344 19136 14384
rect 19176 14344 20448 14384
rect 1152 14320 20448 14344
rect 9435 14216 9477 14225
rect 9435 14176 9436 14216
rect 9476 14176 9477 14216
rect 9435 14167 9477 14176
rect 10011 14216 10053 14225
rect 10011 14176 10012 14216
rect 10052 14176 10053 14216
rect 10011 14167 10053 14176
rect 12363 14216 12405 14225
rect 12363 14176 12364 14216
rect 12404 14176 12405 14216
rect 12363 14167 12405 14176
rect 18507 14216 18549 14225
rect 18507 14176 18508 14216
rect 18548 14176 18549 14216
rect 18507 14167 18549 14176
rect 20235 14216 20277 14225
rect 20235 14176 20236 14216
rect 20276 14176 20277 14216
rect 20235 14167 20277 14176
rect 1851 14132 1893 14141
rect 1851 14092 1852 14132
rect 1892 14092 1893 14132
rect 1851 14083 1893 14092
rect 2235 14132 2277 14141
rect 2235 14092 2236 14132
rect 2276 14092 2277 14132
rect 2235 14083 2277 14092
rect 4731 14132 4773 14141
rect 4731 14092 4732 14132
rect 4772 14092 4773 14132
rect 4731 14083 4773 14092
rect 1227 14048 1269 14057
rect 1227 14008 1228 14048
rect 1268 14008 1269 14048
rect 1227 13999 1269 14008
rect 1611 14048 1653 14057
rect 1611 14008 1612 14048
rect 1652 14008 1653 14048
rect 1611 13999 1653 14008
rect 1995 14048 2037 14057
rect 1995 14008 1996 14048
rect 2036 14008 2037 14048
rect 1995 13999 2037 14008
rect 3051 14048 3093 14057
rect 3051 14008 3052 14048
rect 3092 14008 3093 14048
rect 3051 13999 3093 14008
rect 4491 14048 4533 14057
rect 4491 14008 4492 14048
rect 4532 14008 4533 14048
rect 4491 13999 4533 14008
rect 5067 14048 5109 14057
rect 5067 14008 5068 14048
rect 5108 14008 5109 14048
rect 5067 13999 5109 14008
rect 6027 14048 6069 14057
rect 6027 14008 6028 14048
rect 6068 14008 6069 14048
rect 6027 13999 6069 14008
rect 8043 14048 8085 14057
rect 8043 14008 8044 14048
rect 8084 14008 8085 14048
rect 8043 13999 8085 14008
rect 9322 14048 9380 14049
rect 9322 14008 9331 14048
rect 9371 14008 9380 14048
rect 9322 14007 9380 14008
rect 9675 14048 9717 14057
rect 9675 14008 9676 14048
rect 9716 14008 9717 14048
rect 9675 13999 9717 14008
rect 10251 14048 10293 14057
rect 10251 14008 10252 14048
rect 10292 14008 10293 14048
rect 10251 13999 10293 14008
rect 10539 14048 10581 14057
rect 10539 14008 10540 14048
rect 10580 14008 10581 14048
rect 10539 13999 10581 14008
rect 13611 14048 13653 14057
rect 13611 14008 13612 14048
rect 13652 14008 13653 14048
rect 13611 13999 13653 14008
rect 15627 14048 15669 14057
rect 15627 14008 15628 14048
rect 15668 14008 15669 14048
rect 15627 13999 15669 14008
rect 2554 13964 2612 13965
rect 2554 13924 2563 13964
rect 2603 13924 2612 13964
rect 2554 13923 2612 13924
rect 2667 13964 2709 13973
rect 2667 13924 2668 13964
rect 2708 13924 2709 13964
rect 2667 13915 2709 13924
rect 3147 13964 3189 13973
rect 3147 13924 3148 13964
rect 3188 13924 3189 13964
rect 3147 13915 3189 13924
rect 3619 13964 3677 13965
rect 3619 13924 3628 13964
rect 3668 13924 3677 13964
rect 3619 13923 3677 13924
rect 4107 13964 4165 13965
rect 4107 13924 4116 13964
rect 4156 13924 4165 13964
rect 4107 13923 4165 13924
rect 5530 13964 5588 13965
rect 5530 13924 5539 13964
rect 5579 13924 5588 13964
rect 5530 13923 5588 13924
rect 5643 13964 5685 13973
rect 5643 13924 5644 13964
rect 5684 13924 5685 13964
rect 5643 13915 5685 13924
rect 6123 13964 6165 13973
rect 6123 13924 6124 13964
rect 6164 13924 6165 13964
rect 6123 13915 6165 13924
rect 6595 13964 6653 13965
rect 6595 13924 6604 13964
rect 6644 13924 6653 13964
rect 6595 13923 6653 13924
rect 7083 13964 7141 13965
rect 7083 13924 7092 13964
rect 7132 13924 7141 13964
rect 7083 13923 7141 13924
rect 7546 13964 7604 13965
rect 7546 13924 7555 13964
rect 7595 13924 7604 13964
rect 7546 13923 7604 13924
rect 7659 13964 7701 13973
rect 7659 13924 7660 13964
rect 7700 13924 7701 13964
rect 7659 13915 7701 13924
rect 8139 13964 8181 13973
rect 8139 13924 8140 13964
rect 8180 13924 8181 13964
rect 8139 13915 8181 13924
rect 8611 13964 8669 13965
rect 8611 13924 8620 13964
rect 8660 13924 8669 13964
rect 8611 13923 8669 13924
rect 9099 13964 9157 13965
rect 9099 13924 9108 13964
rect 9148 13924 9157 13964
rect 9099 13923 9157 13924
rect 10923 13964 10965 13973
rect 10923 13924 10924 13964
rect 10964 13924 10965 13964
rect 10923 13915 10965 13924
rect 12163 13964 12221 13965
rect 12163 13924 12172 13964
rect 12212 13924 12221 13964
rect 12163 13923 12221 13924
rect 13114 13964 13172 13965
rect 13114 13924 13123 13964
rect 13163 13924 13172 13964
rect 13114 13923 13172 13924
rect 13227 13964 13269 13973
rect 13227 13924 13228 13964
rect 13268 13924 13269 13964
rect 13227 13915 13269 13924
rect 13707 13964 13749 13973
rect 13707 13924 13708 13964
rect 13748 13924 13749 13964
rect 13707 13915 13749 13924
rect 14179 13964 14237 13965
rect 14179 13924 14188 13964
rect 14228 13924 14237 13964
rect 14179 13923 14237 13924
rect 14667 13964 14725 13965
rect 14667 13924 14676 13964
rect 14716 13924 14725 13964
rect 14667 13923 14725 13924
rect 15130 13964 15188 13965
rect 15130 13924 15139 13964
rect 15179 13924 15188 13964
rect 15130 13923 15188 13924
rect 15243 13964 15285 13973
rect 15243 13924 15244 13964
rect 15284 13924 15285 13964
rect 15243 13915 15285 13924
rect 15723 13964 15765 13973
rect 15723 13924 15724 13964
rect 15764 13924 15765 13964
rect 15723 13915 15765 13924
rect 16195 13964 16253 13965
rect 16195 13924 16204 13964
rect 16244 13924 16253 13964
rect 16195 13923 16253 13924
rect 16714 13964 16772 13965
rect 16714 13924 16723 13964
rect 16763 13924 16772 13964
rect 16714 13923 16772 13924
rect 17067 13964 17109 13973
rect 17067 13924 17068 13964
rect 17108 13924 17109 13964
rect 17067 13915 17109 13924
rect 18307 13964 18365 13965
rect 18307 13924 18316 13964
rect 18356 13924 18365 13964
rect 18307 13923 18365 13924
rect 18795 13964 18837 13973
rect 18795 13924 18796 13964
rect 18836 13924 18837 13964
rect 18795 13915 18837 13924
rect 20035 13964 20093 13965
rect 20035 13924 20044 13964
rect 20084 13924 20093 13964
rect 20035 13923 20093 13924
rect 1467 13880 1509 13889
rect 1467 13840 1468 13880
rect 1508 13840 1509 13880
rect 1467 13831 1509 13840
rect 4827 13880 4869 13889
rect 4827 13840 4828 13880
rect 4868 13840 4869 13880
rect 4827 13831 4869 13840
rect 4299 13796 4341 13805
rect 4299 13756 4300 13796
rect 4340 13756 4341 13796
rect 4299 13747 4341 13756
rect 7275 13796 7317 13805
rect 7275 13756 7276 13796
rect 7316 13756 7317 13796
rect 7275 13747 7317 13756
rect 10779 13796 10821 13805
rect 10779 13756 10780 13796
rect 10820 13756 10821 13796
rect 10779 13747 10821 13756
rect 14859 13796 14901 13805
rect 14859 13756 14860 13796
rect 14900 13756 14901 13796
rect 14859 13747 14901 13756
rect 16875 13796 16917 13805
rect 16875 13756 16876 13796
rect 16916 13756 16917 13796
rect 16875 13747 16917 13756
rect 1152 13628 20452 13652
rect 1152 13588 4928 13628
rect 4968 13588 5010 13628
rect 5050 13588 5092 13628
rect 5132 13588 5174 13628
rect 5214 13588 5256 13628
rect 5296 13588 20048 13628
rect 20088 13588 20130 13628
rect 20170 13588 20212 13628
rect 20252 13588 20294 13628
rect 20334 13588 20376 13628
rect 20416 13588 20452 13628
rect 1152 13564 20452 13588
rect 1467 13460 1509 13469
rect 1467 13420 1468 13460
rect 1508 13420 1509 13460
rect 1467 13411 1509 13420
rect 3051 13460 3093 13469
rect 3051 13420 3052 13460
rect 3092 13420 3093 13460
rect 3051 13411 3093 13420
rect 3579 13460 3621 13469
rect 3579 13420 3580 13460
rect 3620 13420 3621 13460
rect 3579 13411 3621 13420
rect 14379 13460 14421 13469
rect 14379 13420 14380 13460
rect 14420 13420 14421 13460
rect 14379 13411 14421 13420
rect 15483 13460 15525 13469
rect 15483 13420 15484 13460
rect 15524 13420 15525 13460
rect 15483 13411 15525 13420
rect 17355 13460 17397 13469
rect 17355 13420 17356 13460
rect 17396 13420 17397 13460
rect 17355 13411 17397 13420
rect 19851 13460 19893 13469
rect 19851 13420 19852 13460
rect 19892 13420 19893 13460
rect 19851 13411 19893 13420
rect 20091 13460 20133 13469
rect 20091 13420 20092 13460
rect 20132 13420 20133 13460
rect 20091 13411 20133 13420
rect 1611 13292 1653 13301
rect 4107 13292 4149 13301
rect 5835 13292 5877 13301
rect 9579 13292 9621 13301
rect 11211 13292 11253 13301
rect 12939 13292 12981 13301
rect 15915 13292 15957 13301
rect 18106 13292 18164 13293
rect 1611 13252 1612 13292
rect 1652 13252 1653 13292
rect 1611 13243 1653 13252
rect 2859 13283 2901 13292
rect 2859 13243 2860 13283
rect 2900 13243 2901 13283
rect 4107 13252 4108 13292
rect 4148 13252 4149 13292
rect 4107 13243 4149 13252
rect 5355 13283 5397 13292
rect 5355 13243 5356 13283
rect 5396 13243 5397 13283
rect 5835 13252 5836 13292
rect 5876 13252 5877 13292
rect 5835 13243 5877 13252
rect 7083 13283 7125 13292
rect 7083 13243 7084 13283
rect 7124 13243 7125 13283
rect 9579 13252 9580 13292
rect 9620 13252 9621 13292
rect 9579 13243 9621 13252
rect 10827 13283 10869 13292
rect 10827 13243 10828 13283
rect 10868 13243 10869 13283
rect 11211 13252 11212 13292
rect 11252 13252 11253 13292
rect 11211 13243 11253 13252
rect 12459 13283 12501 13292
rect 12459 13243 12460 13283
rect 12500 13243 12501 13283
rect 12939 13252 12940 13292
rect 12980 13252 12981 13292
rect 12939 13243 12981 13252
rect 14187 13283 14229 13292
rect 14187 13243 14188 13283
rect 14228 13243 14229 13283
rect 15915 13252 15916 13292
rect 15956 13252 15957 13292
rect 15915 13243 15957 13252
rect 17163 13283 17205 13292
rect 17163 13243 17164 13283
rect 17204 13243 17205 13283
rect 18106 13252 18115 13292
rect 18155 13252 18164 13292
rect 18106 13251 18164 13252
rect 18219 13292 18261 13301
rect 18219 13252 18220 13292
rect 18260 13252 18261 13292
rect 18219 13243 18261 13252
rect 18603 13292 18645 13301
rect 18603 13252 18604 13292
rect 18644 13252 18645 13292
rect 18603 13243 18645 13252
rect 19179 13283 19221 13292
rect 19179 13243 19180 13283
rect 19220 13243 19221 13283
rect 2859 13234 2901 13243
rect 5355 13234 5397 13243
rect 7083 13234 7125 13243
rect 10827 13234 10869 13243
rect 12459 13234 12501 13243
rect 14187 13234 14229 13243
rect 17163 13234 17205 13243
rect 19179 13234 19221 13243
rect 19659 13283 19701 13292
rect 19659 13243 19660 13283
rect 19700 13243 19701 13283
rect 19659 13234 19701 13243
rect 1227 13208 1269 13217
rect 1227 13168 1228 13208
rect 1268 13168 1269 13208
rect 1227 13159 1269 13168
rect 3243 13208 3285 13217
rect 3243 13168 3244 13208
rect 3284 13168 3285 13208
rect 3243 13159 3285 13168
rect 3819 13208 3861 13217
rect 3819 13168 3820 13208
rect 3860 13168 3861 13208
rect 3819 13159 3861 13168
rect 7947 13208 7989 13217
rect 7947 13168 7948 13208
rect 7988 13168 7989 13208
rect 7947 13159 7989 13168
rect 8331 13208 8373 13217
rect 8331 13168 8332 13208
rect 8372 13168 8373 13208
rect 8331 13159 8373 13168
rect 8715 13208 8757 13217
rect 8715 13168 8716 13208
rect 8756 13168 8757 13208
rect 8715 13159 8757 13168
rect 15723 13208 15765 13217
rect 15723 13168 15724 13208
rect 15764 13168 15765 13208
rect 15723 13159 15765 13168
rect 17739 13208 17781 13217
rect 17739 13168 17740 13208
rect 17780 13168 17781 13208
rect 17739 13159 17781 13168
rect 18699 13208 18741 13217
rect 18699 13168 18700 13208
rect 18740 13168 18741 13208
rect 18699 13159 18741 13168
rect 20331 13208 20373 13217
rect 20331 13168 20332 13208
rect 20372 13168 20373 13208
rect 20331 13159 20373 13168
rect 7275 13124 7317 13133
rect 7275 13084 7276 13124
rect 7316 13084 7317 13124
rect 7275 13075 7317 13084
rect 8091 13124 8133 13133
rect 8091 13084 8092 13124
rect 8132 13084 8133 13124
rect 8091 13075 8133 13084
rect 17499 13124 17541 13133
rect 17499 13084 17500 13124
rect 17540 13084 17541 13124
rect 17499 13075 17541 13084
rect 3483 13040 3525 13049
rect 3483 13000 3484 13040
rect 3524 13000 3525 13040
rect 3483 12991 3525 13000
rect 5547 13040 5589 13049
rect 5547 13000 5548 13040
rect 5588 13000 5589 13040
rect 5547 12991 5589 13000
rect 7707 13040 7749 13049
rect 7707 13000 7708 13040
rect 7748 13000 7749 13040
rect 7707 12991 7749 13000
rect 8475 13040 8517 13049
rect 8475 13000 8476 13040
rect 8516 13000 8517 13040
rect 8475 12991 8517 13000
rect 11019 13040 11061 13049
rect 11019 13000 11020 13040
rect 11060 13000 11061 13040
rect 11019 12991 11061 13000
rect 12651 13040 12693 13049
rect 12651 13000 12652 13040
rect 12692 13000 12693 13040
rect 12651 12991 12693 13000
rect 1152 12872 20448 12896
rect 1152 12832 3688 12872
rect 3728 12832 3770 12872
rect 3810 12832 3852 12872
rect 3892 12832 3934 12872
rect 3974 12832 4016 12872
rect 4056 12832 18808 12872
rect 18848 12832 18890 12872
rect 18930 12832 18972 12872
rect 19012 12832 19054 12872
rect 19094 12832 19136 12872
rect 19176 12832 20448 12872
rect 1152 12808 20448 12832
rect 2235 12704 2277 12713
rect 2235 12664 2236 12704
rect 2276 12664 2277 12704
rect 2235 12655 2277 12664
rect 7227 12704 7269 12713
rect 7227 12664 7228 12704
rect 7268 12664 7269 12704
rect 7227 12655 7269 12664
rect 15243 12704 15285 12713
rect 15243 12664 15244 12704
rect 15284 12664 15285 12704
rect 15243 12655 15285 12664
rect 16875 12704 16917 12713
rect 16875 12664 16876 12704
rect 16916 12664 16917 12704
rect 16875 12655 16917 12664
rect 17403 12704 17445 12713
rect 17403 12664 17404 12704
rect 17444 12664 17445 12704
rect 17403 12655 17445 12664
rect 7611 12620 7653 12629
rect 7611 12580 7612 12620
rect 7652 12580 7653 12620
rect 7611 12571 7653 12580
rect 17019 12620 17061 12629
rect 17019 12580 17020 12620
rect 17060 12580 17061 12620
rect 17019 12571 17061 12580
rect 1227 12536 1269 12545
rect 1227 12496 1228 12536
rect 1268 12496 1269 12536
rect 1227 12487 1269 12496
rect 1611 12536 1653 12545
rect 1611 12496 1612 12536
rect 1652 12496 1653 12536
rect 1611 12487 1653 12496
rect 1995 12536 2037 12545
rect 1995 12496 1996 12536
rect 2036 12496 2037 12536
rect 1995 12487 2037 12496
rect 2955 12536 2997 12545
rect 2955 12496 2956 12536
rect 2996 12496 2997 12536
rect 2955 12487 2997 12496
rect 4395 12536 4437 12545
rect 4395 12496 4396 12536
rect 4436 12496 4437 12536
rect 4395 12487 4437 12496
rect 4635 12536 4677 12545
rect 4635 12496 4636 12536
rect 4676 12496 4677 12536
rect 4635 12487 4677 12496
rect 4875 12536 4917 12545
rect 4875 12496 4876 12536
rect 4916 12496 4917 12536
rect 4875 12487 4917 12496
rect 5115 12536 5157 12545
rect 5115 12496 5116 12536
rect 5156 12496 5157 12536
rect 5115 12487 5157 12496
rect 5835 12536 5877 12545
rect 5835 12496 5836 12536
rect 5876 12496 5877 12536
rect 5835 12487 5877 12496
rect 7114 12536 7172 12537
rect 7114 12496 7123 12536
rect 7163 12496 7172 12536
rect 7114 12495 7172 12496
rect 7467 12536 7509 12545
rect 7467 12496 7468 12536
rect 7508 12496 7509 12536
rect 7467 12487 7509 12496
rect 7851 12536 7893 12545
rect 7851 12496 7852 12536
rect 7892 12496 7893 12536
rect 7851 12487 7893 12496
rect 8427 12536 8469 12545
rect 8427 12496 8428 12536
rect 8468 12496 8469 12536
rect 8427 12487 8469 12496
rect 12363 12536 12405 12545
rect 12363 12496 12364 12536
rect 12404 12496 12405 12536
rect 12363 12487 12405 12496
rect 17259 12536 17301 12545
rect 17259 12496 17260 12536
rect 17300 12496 17301 12536
rect 17259 12487 17301 12496
rect 17643 12536 17685 12545
rect 17643 12496 17644 12536
rect 17684 12496 17685 12536
rect 17643 12487 17685 12496
rect 18411 12536 18453 12545
rect 18411 12496 18412 12536
rect 18452 12496 18453 12536
rect 18411 12487 18453 12496
rect 20331 12536 20373 12545
rect 20331 12496 20332 12536
rect 20372 12496 20373 12536
rect 20331 12487 20373 12496
rect 2458 12452 2516 12453
rect 2458 12412 2467 12452
rect 2507 12412 2516 12452
rect 2458 12411 2516 12412
rect 2571 12452 2613 12461
rect 2571 12412 2572 12452
rect 2612 12412 2613 12452
rect 2571 12403 2613 12412
rect 3051 12452 3093 12461
rect 3051 12412 3052 12452
rect 3092 12412 3093 12452
rect 3051 12403 3093 12412
rect 3523 12452 3581 12453
rect 3523 12412 3532 12452
rect 3572 12412 3581 12452
rect 3523 12411 3581 12412
rect 4011 12452 4069 12453
rect 4011 12412 4020 12452
rect 4060 12412 4069 12452
rect 4011 12411 4069 12412
rect 5338 12452 5396 12453
rect 5338 12412 5347 12452
rect 5387 12412 5396 12452
rect 5338 12411 5396 12412
rect 5451 12452 5493 12461
rect 5451 12412 5452 12452
rect 5492 12412 5493 12452
rect 5451 12403 5493 12412
rect 5931 12452 5973 12461
rect 5931 12412 5932 12452
rect 5972 12412 5973 12452
rect 5931 12403 5973 12412
rect 6403 12452 6461 12453
rect 6403 12412 6412 12452
rect 6452 12412 6461 12452
rect 6403 12411 6461 12412
rect 6895 12452 6953 12453
rect 6895 12412 6904 12452
rect 6944 12412 6953 12452
rect 6895 12411 6953 12412
rect 8619 12452 8661 12461
rect 8619 12412 8620 12452
rect 8660 12412 8661 12452
rect 8619 12403 8661 12412
rect 9859 12452 9917 12453
rect 9859 12412 9868 12452
rect 9908 12412 9917 12452
rect 9859 12411 9917 12412
rect 11853 12452 11895 12461
rect 11853 12412 11854 12452
rect 11894 12412 11895 12452
rect 11853 12403 11895 12412
rect 11968 12452 12026 12453
rect 11968 12412 11977 12452
rect 12017 12412 12026 12452
rect 11968 12411 12026 12412
rect 12459 12452 12501 12461
rect 12459 12412 12460 12452
rect 12500 12412 12501 12452
rect 12459 12403 12501 12412
rect 12931 12452 12989 12453
rect 12931 12412 12940 12452
rect 12980 12412 12989 12452
rect 12931 12411 12989 12412
rect 13419 12452 13477 12453
rect 13419 12412 13428 12452
rect 13468 12412 13477 12452
rect 13419 12411 13477 12412
rect 13803 12452 13845 12461
rect 13803 12412 13804 12452
rect 13844 12412 13845 12452
rect 13803 12403 13845 12412
rect 15043 12452 15101 12453
rect 15043 12412 15052 12452
rect 15092 12412 15101 12452
rect 15043 12411 15101 12412
rect 15435 12452 15477 12461
rect 15435 12412 15436 12452
rect 15476 12412 15477 12452
rect 15435 12403 15477 12412
rect 16675 12452 16733 12453
rect 16675 12412 16684 12452
rect 16724 12412 16733 12452
rect 16675 12411 16733 12412
rect 17901 12452 17943 12461
rect 17901 12412 17902 12452
rect 17942 12412 17943 12452
rect 17901 12403 17943 12412
rect 18027 12452 18069 12461
rect 18027 12412 18028 12452
rect 18068 12412 18069 12452
rect 18027 12403 18069 12412
rect 18507 12452 18549 12461
rect 18507 12412 18508 12452
rect 18548 12412 18549 12452
rect 18507 12403 18549 12412
rect 18979 12452 19037 12453
rect 18979 12412 18988 12452
rect 19028 12412 19037 12452
rect 18979 12411 19037 12412
rect 19467 12452 19525 12453
rect 19467 12412 19476 12452
rect 19516 12412 19525 12452
rect 19467 12411 19525 12412
rect 20091 12368 20133 12377
rect 20091 12328 20092 12368
rect 20132 12328 20133 12368
rect 20091 12319 20133 12328
rect 1467 12284 1509 12293
rect 1467 12244 1468 12284
rect 1508 12244 1509 12284
rect 1467 12235 1509 12244
rect 1851 12284 1893 12293
rect 1851 12244 1852 12284
rect 1892 12244 1893 12284
rect 1851 12235 1893 12244
rect 4203 12284 4245 12293
rect 4203 12244 4204 12284
rect 4244 12244 4245 12284
rect 4203 12235 4245 12244
rect 8187 12284 8229 12293
rect 8187 12244 8188 12284
rect 8228 12244 8229 12284
rect 8187 12235 8229 12244
rect 10059 12284 10101 12293
rect 10059 12244 10060 12284
rect 10100 12244 10101 12284
rect 10059 12235 10101 12244
rect 13611 12284 13653 12293
rect 13611 12244 13612 12284
rect 13652 12244 13653 12284
rect 13611 12235 13653 12244
rect 19659 12284 19701 12293
rect 19659 12244 19660 12284
rect 19700 12244 19701 12284
rect 19659 12235 19701 12244
rect 1152 12116 20452 12140
rect 1152 12076 4928 12116
rect 4968 12076 5010 12116
rect 5050 12076 5092 12116
rect 5132 12076 5174 12116
rect 5214 12076 5256 12116
rect 5296 12076 20048 12116
rect 20088 12076 20130 12116
rect 20170 12076 20212 12116
rect 20252 12076 20294 12116
rect 20334 12076 20376 12116
rect 20416 12076 20452 12116
rect 1152 12052 20452 12076
rect 1179 11948 1221 11957
rect 1179 11908 1180 11948
rect 1220 11908 1221 11948
rect 1179 11899 1221 11908
rect 1563 11948 1605 11957
rect 1563 11908 1564 11948
rect 1604 11908 1605 11948
rect 1563 11899 1605 11908
rect 3627 11948 3669 11957
rect 3627 11908 3628 11948
rect 3668 11908 3669 11948
rect 3627 11899 3669 11908
rect 6507 11948 6549 11957
rect 6507 11908 6508 11948
rect 6548 11908 6549 11948
rect 6507 11899 6549 11908
rect 8427 11948 8469 11957
rect 8427 11908 8428 11948
rect 8468 11908 8469 11948
rect 8427 11899 8469 11908
rect 16443 11948 16485 11957
rect 16443 11908 16444 11948
rect 16484 11908 16485 11948
rect 16443 11899 16485 11908
rect 18315 11948 18357 11957
rect 18315 11908 18316 11948
rect 18356 11908 18357 11948
rect 18315 11899 18357 11908
rect 3771 11864 3813 11873
rect 3771 11824 3772 11864
rect 3812 11824 3813 11864
rect 3771 11815 3813 11824
rect 13131 11864 13173 11873
rect 13131 11824 13132 11864
rect 13172 11824 13173 11864
rect 13131 11815 13173 11824
rect 16347 11864 16389 11873
rect 16347 11824 16348 11864
rect 16388 11824 16389 11864
rect 16347 11815 16389 11824
rect 20091 11864 20133 11873
rect 20091 11824 20092 11864
rect 20132 11824 20133 11864
rect 20091 11815 20133 11824
rect 2187 11780 2229 11789
rect 5067 11780 5109 11789
rect 6987 11780 7029 11789
rect 8698 11780 8756 11781
rect 2187 11740 2188 11780
rect 2228 11740 2229 11780
rect 2187 11731 2229 11740
rect 3439 11771 3481 11780
rect 3439 11731 3440 11771
rect 3480 11731 3481 11771
rect 5067 11740 5068 11780
rect 5108 11740 5109 11780
rect 5067 11731 5109 11740
rect 6315 11771 6357 11780
rect 6315 11731 6316 11771
rect 6356 11731 6357 11771
rect 6987 11740 6988 11780
rect 7028 11740 7029 11780
rect 6987 11731 7029 11740
rect 8235 11771 8277 11780
rect 8235 11731 8236 11771
rect 8276 11731 8277 11771
rect 8698 11740 8707 11780
rect 8747 11740 8756 11780
rect 8698 11739 8756 11740
rect 8811 11780 8853 11789
rect 8811 11740 8812 11780
rect 8852 11740 8853 11780
rect 8811 11731 8853 11740
rect 9195 11780 9237 11789
rect 11691 11780 11733 11789
rect 13402 11780 13460 11781
rect 9195 11740 9196 11780
rect 9236 11740 9237 11780
rect 9195 11731 9237 11740
rect 9771 11771 9813 11780
rect 9771 11731 9772 11771
rect 9812 11731 9813 11771
rect 3439 11722 3481 11731
rect 6315 11722 6357 11731
rect 8235 11722 8277 11731
rect 9771 11722 9813 11731
rect 10251 11771 10293 11780
rect 10251 11731 10252 11771
rect 10292 11731 10293 11771
rect 11691 11740 11692 11780
rect 11732 11740 11733 11780
rect 11691 11731 11733 11740
rect 12939 11771 12981 11780
rect 12939 11731 12940 11771
rect 12980 11731 12981 11771
rect 13402 11740 13411 11780
rect 13451 11740 13460 11780
rect 13402 11739 13460 11740
rect 13515 11780 13557 11789
rect 13515 11740 13516 11780
rect 13556 11740 13557 11780
rect 13515 11731 13557 11740
rect 13899 11780 13941 11789
rect 16875 11780 16917 11789
rect 18507 11780 18549 11789
rect 13899 11740 13900 11780
rect 13940 11740 13941 11780
rect 13899 11731 13941 11740
rect 14475 11771 14517 11780
rect 14475 11731 14476 11771
rect 14516 11731 14517 11771
rect 10251 11722 10293 11731
rect 12939 11722 12981 11731
rect 14475 11722 14517 11731
rect 14955 11771 14997 11780
rect 14955 11731 14956 11771
rect 14996 11731 14997 11771
rect 16875 11740 16876 11780
rect 16916 11740 16917 11780
rect 16875 11731 16917 11740
rect 18123 11771 18165 11780
rect 18123 11731 18124 11771
rect 18164 11731 18165 11771
rect 18507 11740 18508 11780
rect 18548 11740 18549 11780
rect 18507 11731 18549 11740
rect 19755 11771 19797 11780
rect 19755 11731 19756 11771
rect 19796 11731 19797 11771
rect 14955 11722 14997 11731
rect 18123 11722 18165 11731
rect 19755 11722 19797 11731
rect 1419 11696 1461 11705
rect 1419 11656 1420 11696
rect 1460 11656 1461 11696
rect 1419 11647 1461 11656
rect 1803 11696 1845 11705
rect 1803 11656 1804 11696
rect 1844 11656 1845 11696
rect 1803 11647 1845 11656
rect 4011 11696 4053 11705
rect 4011 11656 4012 11696
rect 4052 11656 4053 11696
rect 4011 11647 4053 11656
rect 4491 11696 4533 11705
rect 4491 11656 4492 11696
rect 4532 11656 4533 11696
rect 4491 11647 4533 11656
rect 4875 11696 4917 11705
rect 4875 11656 4876 11696
rect 4916 11656 4917 11696
rect 4875 11647 4917 11656
rect 9291 11696 9333 11705
rect 9291 11656 9292 11696
rect 9332 11656 9333 11696
rect 9291 11647 9333 11656
rect 10474 11696 10532 11697
rect 10474 11656 10483 11696
rect 10523 11656 10532 11696
rect 10474 11655 10532 11656
rect 10827 11696 10869 11705
rect 10827 11656 10828 11696
rect 10868 11656 10869 11696
rect 10827 11647 10869 11656
rect 13995 11696 14037 11705
rect 13995 11656 13996 11696
rect 14036 11656 14037 11696
rect 13995 11647 14037 11656
rect 15178 11696 15236 11697
rect 15178 11656 15187 11696
rect 15227 11656 15236 11696
rect 15178 11655 15236 11656
rect 15531 11696 15573 11705
rect 15531 11656 15532 11696
rect 15572 11656 15573 11696
rect 15531 11647 15573 11656
rect 16107 11696 16149 11705
rect 16107 11656 16108 11696
rect 16148 11656 16149 11696
rect 16107 11647 16149 11656
rect 16683 11696 16725 11705
rect 16683 11656 16684 11696
rect 16724 11656 16725 11696
rect 16683 11647 16725 11656
rect 20331 11696 20373 11705
rect 20331 11656 20332 11696
rect 20372 11656 20373 11696
rect 20331 11647 20373 11656
rect 4251 11612 4293 11621
rect 4251 11572 4252 11612
rect 4292 11572 4293 11612
rect 4251 11563 4293 11572
rect 4635 11612 4677 11621
rect 4635 11572 4636 11612
rect 4676 11572 4677 11612
rect 4635 11563 4677 11572
rect 15291 11612 15333 11621
rect 15291 11572 15292 11612
rect 15332 11572 15333 11612
rect 15291 11563 15333 11572
rect 19947 11612 19989 11621
rect 19947 11572 19948 11612
rect 19988 11572 19989 11612
rect 19947 11563 19989 11572
rect 10587 11528 10629 11537
rect 10587 11488 10588 11528
rect 10628 11488 10629 11528
rect 10587 11479 10629 11488
rect 1152 11360 20448 11384
rect 1152 11320 3688 11360
rect 3728 11320 3770 11360
rect 3810 11320 3852 11360
rect 3892 11320 3934 11360
rect 3974 11320 4016 11360
rect 4056 11320 18808 11360
rect 18848 11320 18890 11360
rect 18930 11320 18972 11360
rect 19012 11320 19054 11360
rect 19094 11320 19136 11360
rect 19176 11320 20448 11360
rect 1152 11296 20448 11320
rect 2667 11192 2709 11201
rect 2667 11152 2668 11192
rect 2708 11152 2709 11192
rect 2667 11143 2709 11152
rect 3483 11192 3525 11201
rect 3483 11152 3484 11192
rect 3524 11152 3525 11192
rect 3483 11143 3525 11152
rect 8043 11192 8085 11201
rect 8043 11152 8044 11192
rect 8084 11152 8085 11192
rect 8043 11143 8085 11152
rect 15051 11192 15093 11201
rect 15051 11152 15052 11192
rect 15092 11152 15093 11192
rect 15051 11143 15093 11152
rect 19371 11192 19413 11201
rect 19371 11152 19372 11192
rect 19412 11152 19413 11192
rect 19371 11143 19413 11152
rect 19707 11192 19749 11201
rect 19707 11152 19708 11192
rect 19748 11152 19749 11192
rect 19707 11143 19749 11152
rect 20091 11192 20133 11201
rect 20091 11152 20092 11192
rect 20132 11152 20133 11192
rect 20091 11143 20133 11152
rect 2811 11108 2853 11117
rect 2811 11068 2812 11108
rect 2852 11068 2853 11108
rect 2811 11059 2853 11068
rect 3051 11024 3093 11033
rect 3051 10984 3052 11024
rect 3092 10984 3093 11024
rect 3051 10975 3093 10984
rect 3243 11024 3285 11033
rect 3243 10984 3244 11024
rect 3284 10984 3285 11024
rect 3243 10975 3285 10984
rect 3819 11024 3861 11033
rect 3819 10984 3820 11024
rect 3860 10984 3861 11024
rect 3819 10975 3861 10984
rect 4011 11024 4053 11033
rect 4011 10984 4012 11024
rect 4052 10984 4053 11024
rect 4011 10975 4053 10984
rect 6603 11024 6645 11033
rect 6603 10984 6604 11024
rect 6644 10984 6645 11024
rect 6603 10975 6645 10984
rect 11979 11024 12021 11033
rect 11979 10984 11980 11024
rect 12020 10984 12021 11024
rect 11979 10975 12021 10984
rect 15915 11024 15957 11033
rect 15915 10984 15916 11024
rect 15956 10984 15957 11024
rect 15915 10975 15957 10984
rect 17194 11024 17252 11025
rect 17194 10984 17203 11024
rect 17243 10984 17252 11024
rect 17194 10983 17252 10984
rect 17547 11024 17589 11033
rect 17547 10984 17548 11024
rect 17588 10984 17589 11024
rect 17547 10975 17589 10984
rect 19947 11024 19989 11033
rect 19947 10984 19948 11024
rect 19988 10984 19989 11024
rect 19947 10975 19989 10984
rect 20331 11024 20373 11033
rect 20331 10984 20332 11024
rect 20372 10984 20373 11024
rect 20331 10975 20373 10984
rect 1227 10940 1269 10949
rect 1227 10900 1228 10940
rect 1268 10900 1269 10940
rect 1227 10891 1269 10900
rect 2467 10940 2525 10941
rect 2467 10900 2476 10940
rect 2516 10900 2525 10940
rect 2467 10899 2525 10900
rect 4395 10940 4437 10949
rect 4395 10900 4396 10940
rect 4436 10900 4437 10940
rect 4395 10891 4437 10900
rect 5635 10940 5693 10941
rect 5635 10900 5644 10940
rect 5684 10900 5693 10940
rect 5635 10899 5693 10900
rect 6106 10940 6164 10941
rect 6106 10900 6115 10940
rect 6155 10900 6164 10940
rect 6106 10899 6164 10900
rect 6219 10940 6261 10949
rect 6219 10900 6220 10940
rect 6260 10900 6261 10940
rect 6219 10891 6261 10900
rect 6699 10940 6741 10949
rect 6699 10900 6700 10940
rect 6740 10900 6741 10940
rect 6699 10891 6741 10900
rect 7171 10940 7229 10941
rect 7171 10900 7180 10940
rect 7220 10900 7229 10940
rect 7171 10899 7229 10900
rect 7690 10940 7748 10941
rect 7690 10900 7699 10940
rect 7739 10900 7748 10940
rect 7690 10899 7748 10900
rect 8227 10940 8285 10941
rect 8227 10900 8236 10940
rect 8276 10900 8285 10940
rect 8227 10899 8285 10900
rect 9483 10940 9525 10949
rect 9483 10900 9484 10940
rect 9524 10900 9525 10940
rect 9483 10891 9525 10900
rect 9771 10940 9813 10949
rect 9771 10900 9772 10940
rect 9812 10900 9813 10940
rect 9771 10891 9813 10900
rect 11011 10940 11069 10941
rect 11011 10900 11020 10940
rect 11060 10900 11069 10940
rect 11011 10899 11069 10900
rect 11482 10940 11540 10941
rect 11482 10900 11491 10940
rect 11531 10900 11540 10940
rect 11482 10899 11540 10900
rect 11595 10940 11637 10949
rect 11595 10900 11596 10940
rect 11636 10900 11637 10940
rect 11595 10891 11637 10900
rect 12075 10940 12117 10949
rect 12075 10900 12076 10940
rect 12116 10900 12117 10940
rect 12075 10891 12117 10900
rect 12547 10940 12605 10941
rect 12547 10900 12556 10940
rect 12596 10900 12605 10940
rect 12547 10899 12605 10900
rect 13035 10940 13093 10941
rect 13035 10900 13044 10940
rect 13084 10900 13093 10940
rect 13035 10899 13093 10900
rect 13611 10940 13653 10949
rect 13611 10900 13612 10940
rect 13652 10900 13653 10940
rect 13611 10891 13653 10900
rect 14851 10940 14909 10941
rect 14851 10900 14860 10940
rect 14900 10900 14909 10940
rect 14851 10899 14909 10900
rect 15418 10940 15476 10941
rect 15418 10900 15427 10940
rect 15467 10900 15476 10940
rect 15418 10899 15476 10900
rect 15531 10940 15573 10949
rect 15531 10900 15532 10940
rect 15572 10900 15573 10940
rect 15531 10891 15573 10900
rect 16011 10940 16053 10949
rect 16011 10900 16012 10940
rect 16052 10900 16053 10940
rect 16011 10891 16053 10900
rect 16483 10940 16541 10941
rect 16483 10900 16492 10940
rect 16532 10900 16541 10940
rect 16483 10899 16541 10900
rect 16971 10940 17029 10941
rect 16971 10900 16980 10940
rect 17020 10900 17029 10940
rect 16971 10899 17029 10900
rect 17931 10940 17973 10949
rect 17931 10900 17932 10940
rect 17972 10900 17973 10940
rect 17931 10891 17973 10900
rect 19171 10940 19229 10941
rect 19171 10900 19180 10940
rect 19220 10900 19229 10940
rect 19171 10899 19229 10900
rect 5835 10856 5877 10865
rect 5835 10816 5836 10856
rect 5876 10816 5877 10856
rect 5835 10807 5877 10816
rect 11211 10856 11253 10865
rect 11211 10816 11212 10856
rect 11252 10816 11253 10856
rect 11211 10807 11253 10816
rect 3579 10772 3621 10781
rect 3579 10732 3580 10772
rect 3620 10732 3621 10772
rect 3579 10723 3621 10732
rect 4251 10772 4293 10781
rect 4251 10732 4252 10772
rect 4292 10732 4293 10772
rect 4251 10723 4293 10732
rect 7851 10772 7893 10781
rect 7851 10732 7852 10772
rect 7892 10732 7893 10772
rect 7851 10723 7893 10732
rect 13227 10772 13269 10781
rect 13227 10732 13228 10772
rect 13268 10732 13269 10772
rect 13227 10723 13269 10732
rect 17307 10772 17349 10781
rect 17307 10732 17308 10772
rect 17348 10732 17349 10772
rect 17307 10723 17349 10732
rect 1152 10604 20452 10628
rect 1152 10564 4928 10604
rect 4968 10564 5010 10604
rect 5050 10564 5092 10604
rect 5132 10564 5174 10604
rect 5214 10564 5256 10604
rect 5296 10564 20048 10604
rect 20088 10564 20130 10604
rect 20170 10564 20212 10604
rect 20252 10564 20294 10604
rect 20334 10564 20376 10604
rect 20416 10564 20452 10604
rect 1152 10540 20452 10564
rect 1179 10436 1221 10445
rect 1179 10396 1180 10436
rect 1220 10396 1221 10436
rect 1179 10387 1221 10396
rect 2235 10436 2277 10445
rect 2235 10396 2236 10436
rect 2276 10396 2277 10436
rect 2235 10387 2277 10396
rect 4587 10436 4629 10445
rect 4587 10396 4588 10436
rect 4628 10396 4629 10436
rect 4587 10387 4629 10396
rect 7947 10436 7989 10445
rect 7947 10396 7948 10436
rect 7988 10396 7989 10436
rect 7947 10387 7989 10396
rect 12171 10436 12213 10445
rect 12171 10396 12172 10436
rect 12212 10396 12213 10436
rect 12171 10387 12213 10396
rect 14187 10436 14229 10445
rect 14187 10396 14188 10436
rect 14228 10396 14229 10436
rect 14187 10387 14229 10396
rect 15819 10436 15861 10445
rect 15819 10396 15820 10436
rect 15860 10396 15861 10436
rect 15819 10387 15861 10396
rect 17643 10436 17685 10445
rect 17643 10396 17644 10436
rect 17684 10396 17685 10436
rect 17643 10387 17685 10396
rect 20091 10436 20133 10445
rect 20091 10396 20092 10436
rect 20132 10396 20133 10436
rect 20091 10387 20133 10396
rect 17914 10352 17972 10353
rect 17914 10312 17923 10352
rect 17963 10312 17972 10352
rect 17914 10311 17972 10312
rect 2938 10301 2996 10306
rect 2829 10268 2871 10277
rect 2829 10228 2830 10268
rect 2870 10228 2871 10268
rect 2938 10261 2947 10301
rect 2987 10261 2996 10301
rect 2938 10260 2996 10261
rect 3339 10268 3381 10277
rect 4779 10268 4821 10277
rect 6507 10268 6549 10277
rect 10731 10268 10773 10277
rect 12442 10268 12500 10269
rect 2829 10219 2871 10228
rect 3339 10228 3340 10268
rect 3380 10228 3381 10268
rect 3339 10219 3381 10228
rect 3915 10259 3957 10268
rect 3915 10219 3916 10259
rect 3956 10219 3957 10259
rect 3915 10210 3957 10219
rect 4395 10259 4437 10268
rect 4395 10219 4396 10259
rect 4436 10219 4437 10259
rect 4779 10228 4780 10268
rect 4820 10228 4821 10268
rect 4779 10219 4821 10228
rect 6027 10259 6069 10268
rect 6027 10219 6028 10259
rect 6068 10219 6069 10259
rect 6507 10228 6508 10268
rect 6548 10228 6549 10268
rect 6507 10219 6549 10228
rect 7755 10259 7797 10268
rect 7755 10219 7756 10259
rect 7796 10219 7797 10259
rect 10731 10228 10732 10268
rect 10772 10228 10773 10268
rect 10731 10219 10773 10228
rect 11979 10259 12021 10268
rect 11979 10219 11980 10259
rect 12020 10219 12021 10259
rect 12442 10228 12451 10268
rect 12491 10228 12500 10268
rect 12442 10227 12500 10228
rect 12555 10268 12597 10277
rect 12555 10228 12556 10268
rect 12596 10228 12597 10268
rect 12555 10219 12597 10228
rect 12939 10268 12981 10277
rect 14379 10268 14421 10277
rect 16203 10268 16245 10277
rect 18106 10268 18164 10269
rect 19083 10268 19125 10277
rect 12939 10228 12940 10268
rect 12980 10228 12981 10268
rect 12939 10219 12981 10228
rect 13515 10259 13557 10268
rect 13515 10219 13516 10259
rect 13556 10219 13557 10259
rect 4395 10210 4437 10219
rect 6027 10210 6069 10219
rect 7755 10210 7797 10219
rect 11979 10210 12021 10219
rect 13515 10210 13557 10219
rect 13995 10259 14037 10268
rect 13995 10219 13996 10259
rect 14036 10219 14037 10259
rect 14379 10228 14380 10268
rect 14420 10228 14421 10268
rect 14379 10219 14421 10228
rect 15627 10259 15669 10268
rect 15627 10219 15628 10259
rect 15668 10219 15669 10259
rect 16203 10228 16204 10268
rect 16244 10228 16245 10268
rect 16203 10219 16245 10228
rect 17451 10259 17493 10268
rect 17451 10219 17452 10259
rect 17492 10219 17493 10259
rect 18106 10228 18115 10268
rect 18155 10228 18164 10268
rect 18106 10227 18164 10228
rect 18603 10259 18645 10268
rect 13995 10210 14037 10219
rect 15627 10210 15669 10219
rect 17451 10210 17493 10219
rect 18603 10219 18604 10259
rect 18644 10219 18645 10259
rect 19083 10228 19084 10268
rect 19124 10228 19125 10268
rect 19083 10219 19125 10228
rect 19563 10268 19605 10277
rect 19563 10228 19564 10268
rect 19604 10228 19605 10268
rect 19563 10219 19605 10228
rect 19676 10249 19718 10258
rect 18603 10210 18645 10219
rect 19676 10209 19677 10249
rect 19717 10209 19718 10249
rect 19676 10200 19718 10209
rect 1419 10184 1461 10193
rect 1419 10144 1420 10184
rect 1460 10144 1461 10184
rect 1419 10135 1461 10144
rect 1899 10184 1941 10193
rect 1899 10144 1900 10184
rect 1940 10144 1941 10184
rect 1899 10135 1941 10144
rect 2139 10184 2181 10193
rect 2139 10144 2140 10184
rect 2180 10144 2181 10184
rect 2139 10135 2181 10144
rect 2475 10184 2517 10193
rect 2475 10144 2476 10184
rect 2516 10144 2517 10184
rect 2475 10135 2517 10144
rect 3435 10184 3477 10193
rect 3435 10144 3436 10184
rect 3476 10144 3477 10184
rect 3435 10135 3477 10144
rect 8331 10184 8373 10193
rect 8331 10144 8332 10184
rect 8372 10144 8373 10184
rect 8331 10135 8373 10144
rect 13035 10184 13077 10193
rect 13035 10144 13036 10184
rect 13076 10144 13077 10184
rect 13035 10135 13077 10144
rect 19179 10184 19221 10193
rect 19179 10144 19180 10184
rect 19220 10144 19221 10184
rect 19179 10135 19221 10144
rect 20331 10184 20373 10193
rect 20331 10144 20332 10184
rect 20372 10144 20373 10184
rect 20331 10135 20373 10144
rect 8091 10100 8133 10109
rect 8091 10060 8092 10100
rect 8132 10060 8133 10100
rect 8091 10051 8133 10060
rect 6219 10016 6261 10025
rect 6219 9976 6220 10016
rect 6260 9976 6261 10016
rect 6219 9967 6261 9976
rect 1152 9848 20448 9872
rect 1152 9808 3688 9848
rect 3728 9808 3770 9848
rect 3810 9808 3852 9848
rect 3892 9808 3934 9848
rect 3974 9808 4016 9848
rect 4056 9808 18808 9848
rect 18848 9808 18890 9848
rect 18930 9808 18972 9848
rect 19012 9808 19054 9848
rect 19094 9808 19136 9848
rect 19176 9808 20448 9848
rect 1152 9784 20448 9808
rect 1179 9680 1221 9689
rect 1179 9640 1180 9680
rect 1220 9640 1221 9680
rect 1179 9631 1221 9640
rect 3483 9680 3525 9689
rect 3483 9640 3484 9680
rect 3524 9640 3525 9680
rect 3483 9631 3525 9640
rect 6075 9680 6117 9689
rect 6075 9640 6076 9680
rect 6116 9640 6117 9680
rect 6075 9631 6117 9640
rect 14218 9680 14276 9681
rect 14218 9640 14227 9680
rect 14267 9640 14276 9680
rect 14218 9639 14276 9640
rect 15291 9680 15333 9689
rect 15291 9640 15292 9680
rect 15332 9640 15333 9680
rect 15291 9631 15333 9640
rect 16875 9680 16917 9689
rect 16875 9640 16876 9680
rect 16916 9640 16917 9680
rect 16875 9631 16917 9640
rect 20091 9680 20133 9689
rect 20091 9640 20092 9680
rect 20132 9640 20133 9680
rect 20091 9631 20133 9640
rect 3339 9596 3381 9605
rect 3339 9556 3340 9596
rect 3380 9556 3381 9596
rect 3339 9547 3381 9556
rect 11163 9596 11205 9605
rect 11163 9556 11164 9596
rect 11204 9556 11205 9596
rect 11163 9547 11205 9556
rect 1419 9512 1461 9521
rect 1419 9472 1420 9512
rect 1460 9472 1461 9512
rect 1419 9463 1461 9472
rect 3723 9512 3765 9521
rect 3723 9472 3724 9512
rect 3764 9472 3765 9512
rect 3723 9463 3765 9472
rect 4683 9512 4725 9521
rect 4683 9472 4684 9512
rect 4724 9472 4725 9512
rect 4683 9463 4725 9472
rect 5962 9512 6020 9513
rect 5962 9472 5971 9512
rect 6011 9472 6020 9512
rect 5962 9471 6020 9472
rect 6315 9512 6357 9521
rect 6315 9472 6316 9512
rect 6356 9472 6357 9512
rect 6315 9463 6357 9472
rect 6891 9512 6933 9521
rect 6891 9472 6892 9512
rect 6932 9472 6933 9512
rect 6891 9463 6933 9472
rect 9771 9512 9813 9521
rect 9771 9472 9772 9512
rect 9812 9472 9813 9512
rect 9771 9463 9813 9472
rect 11050 9512 11108 9513
rect 11050 9472 11059 9512
rect 11099 9472 11108 9512
rect 11050 9471 11108 9472
rect 11403 9512 11445 9521
rect 11403 9472 11404 9512
rect 11444 9472 11445 9512
rect 11403 9463 11445 9472
rect 12939 9512 12981 9521
rect 12939 9472 12940 9512
rect 12980 9472 12981 9512
rect 12939 9463 12981 9472
rect 14571 9512 14613 9521
rect 14571 9472 14572 9512
rect 14612 9472 14613 9512
rect 14571 9463 14613 9472
rect 15051 9512 15093 9521
rect 15051 9472 15052 9512
rect 15092 9472 15093 9512
rect 15051 9463 15093 9472
rect 17259 9512 17301 9521
rect 17259 9472 17260 9512
rect 17300 9472 17301 9512
rect 17259 9463 17301 9472
rect 17643 9512 17685 9521
rect 17643 9472 17644 9512
rect 17684 9472 17685 9512
rect 17643 9463 17685 9472
rect 18411 9512 18453 9521
rect 18411 9472 18412 9512
rect 18452 9472 18453 9512
rect 18411 9463 18453 9472
rect 20331 9512 20373 9521
rect 20331 9472 20332 9512
rect 20372 9472 20373 9512
rect 20331 9463 20373 9472
rect 1899 9428 1941 9437
rect 1899 9388 1900 9428
rect 1940 9388 1941 9428
rect 1899 9379 1941 9388
rect 3139 9428 3197 9429
rect 3139 9388 3148 9428
rect 3188 9388 3197 9428
rect 3139 9387 3197 9388
rect 4186 9428 4244 9429
rect 4186 9388 4195 9428
rect 4235 9388 4244 9428
rect 4186 9387 4244 9388
rect 4299 9428 4341 9437
rect 4299 9388 4300 9428
rect 4340 9388 4341 9428
rect 4299 9379 4341 9388
rect 4779 9428 4821 9437
rect 4779 9388 4780 9428
rect 4820 9388 4821 9428
rect 4779 9379 4821 9388
rect 5251 9428 5309 9429
rect 5251 9388 5260 9428
rect 5300 9388 5309 9428
rect 5251 9387 5309 9388
rect 5770 9428 5828 9429
rect 5770 9388 5779 9428
rect 5819 9388 5828 9428
rect 5770 9387 5828 9388
rect 7563 9428 7605 9437
rect 7563 9388 7564 9428
rect 7604 9388 7605 9428
rect 7563 9379 7605 9388
rect 8803 9428 8861 9429
rect 8803 9388 8812 9428
rect 8852 9388 8861 9428
rect 8803 9387 8861 9388
rect 9274 9428 9332 9429
rect 9274 9388 9283 9428
rect 9323 9388 9332 9428
rect 9274 9387 9332 9388
rect 9387 9428 9429 9437
rect 9387 9388 9388 9428
rect 9428 9388 9429 9428
rect 9387 9379 9429 9388
rect 9867 9428 9909 9437
rect 9867 9388 9868 9428
rect 9908 9388 9909 9428
rect 9867 9379 9909 9388
rect 10339 9428 10397 9429
rect 10339 9388 10348 9428
rect 10388 9388 10397 9428
rect 10339 9387 10397 9388
rect 10827 9428 10885 9429
rect 10827 9388 10836 9428
rect 10876 9388 10885 9428
rect 10827 9387 10885 9388
rect 12442 9428 12500 9429
rect 12442 9388 12451 9428
rect 12491 9388 12500 9428
rect 12442 9387 12500 9388
rect 12555 9428 12597 9437
rect 12555 9388 12556 9428
rect 12596 9388 12597 9428
rect 12555 9379 12597 9388
rect 13035 9428 13077 9437
rect 13035 9388 13036 9428
rect 13076 9388 13077 9428
rect 13035 9379 13077 9388
rect 13507 9428 13565 9429
rect 13507 9388 13516 9428
rect 13556 9388 13565 9428
rect 13507 9387 13565 9388
rect 14026 9428 14084 9429
rect 14026 9388 14035 9428
rect 14075 9388 14084 9428
rect 14026 9387 14084 9388
rect 15435 9428 15477 9437
rect 15435 9388 15436 9428
rect 15476 9388 15477 9428
rect 15435 9379 15477 9388
rect 16675 9428 16733 9429
rect 16675 9388 16684 9428
rect 16724 9388 16733 9428
rect 16675 9387 16733 9388
rect 17914 9428 17972 9429
rect 17914 9388 17923 9428
rect 17963 9388 17972 9428
rect 17914 9387 17972 9388
rect 18027 9428 18069 9437
rect 18027 9388 18028 9428
rect 18068 9388 18069 9428
rect 18027 9379 18069 9388
rect 18507 9428 18549 9437
rect 18507 9388 18508 9428
rect 18548 9388 18549 9428
rect 18507 9379 18549 9388
rect 18979 9428 19037 9429
rect 18979 9388 18988 9428
rect 19028 9388 19037 9428
rect 18979 9387 19037 9388
rect 19498 9428 19556 9429
rect 19498 9388 19507 9428
rect 19547 9388 19556 9428
rect 19498 9387 19556 9388
rect 9003 9344 9045 9353
rect 9003 9304 9004 9344
rect 9044 9304 9045 9344
rect 9003 9295 9045 9304
rect 6651 9260 6693 9269
rect 6651 9220 6652 9260
rect 6692 9220 6693 9260
rect 6651 9211 6693 9220
rect 14331 9260 14373 9269
rect 14331 9220 14332 9260
rect 14372 9220 14373 9260
rect 14331 9211 14373 9220
rect 17019 9260 17061 9269
rect 17019 9220 17020 9260
rect 17060 9220 17061 9260
rect 17019 9211 17061 9220
rect 17403 9260 17445 9269
rect 17403 9220 17404 9260
rect 17444 9220 17445 9260
rect 17403 9211 17445 9220
rect 19659 9260 19701 9269
rect 19659 9220 19660 9260
rect 19700 9220 19701 9260
rect 19659 9211 19701 9220
rect 1152 9092 20452 9116
rect 1152 9052 4928 9092
rect 4968 9052 5010 9092
rect 5050 9052 5092 9092
rect 5132 9052 5174 9092
rect 5214 9052 5256 9092
rect 5296 9052 20048 9092
rect 20088 9052 20130 9092
rect 20170 9052 20212 9092
rect 20252 9052 20294 9092
rect 20334 9052 20376 9092
rect 20416 9052 20452 9092
rect 1152 9028 20452 9052
rect 2667 8924 2709 8933
rect 2667 8884 2668 8924
rect 2708 8884 2709 8924
rect 2667 8875 2709 8884
rect 11883 8924 11925 8933
rect 11883 8884 11884 8924
rect 11924 8884 11925 8924
rect 11883 8875 11925 8884
rect 13995 8924 14037 8933
rect 13995 8884 13996 8924
rect 14036 8884 14037 8924
rect 13995 8875 14037 8884
rect 15291 8924 15333 8933
rect 15291 8884 15292 8924
rect 15332 8884 15333 8924
rect 15291 8875 15333 8884
rect 17547 8924 17589 8933
rect 17547 8884 17548 8924
rect 17588 8884 17589 8924
rect 17547 8875 17589 8884
rect 19179 8924 19221 8933
rect 19179 8884 19180 8924
rect 19220 8884 19221 8924
rect 19179 8875 19221 8884
rect 20091 8924 20133 8933
rect 20091 8884 20092 8924
rect 20132 8884 20133 8924
rect 20091 8875 20133 8884
rect 2811 8840 2853 8849
rect 2811 8800 2812 8840
rect 2852 8800 2853 8840
rect 2811 8791 2853 8800
rect 3771 8840 3813 8849
rect 3771 8800 3772 8840
rect 3812 8800 3813 8840
rect 3771 8791 3813 8800
rect 8187 8840 8229 8849
rect 8187 8800 8188 8840
rect 8228 8800 8229 8840
rect 8187 8791 8229 8800
rect 15099 8840 15141 8849
rect 15099 8800 15100 8840
rect 15140 8800 15141 8840
rect 15099 8791 15141 8800
rect 19707 8840 19749 8849
rect 19707 8800 19708 8840
rect 19748 8800 19749 8840
rect 19707 8791 19749 8800
rect 1227 8756 1269 8765
rect 4282 8756 4340 8757
rect 1227 8716 1228 8756
rect 1268 8716 1269 8756
rect 1227 8707 1269 8716
rect 2475 8747 2517 8756
rect 2475 8707 2476 8747
rect 2516 8707 2517 8747
rect 4282 8716 4291 8756
rect 4331 8716 4340 8756
rect 4282 8715 4340 8716
rect 4395 8756 4437 8765
rect 4395 8716 4396 8756
rect 4436 8716 4437 8756
rect 4395 8707 4437 8716
rect 4779 8756 4821 8765
rect 6298 8756 6356 8757
rect 4779 8716 4780 8756
rect 4820 8716 4821 8756
rect 4779 8707 4821 8716
rect 5355 8747 5397 8756
rect 5355 8707 5356 8747
rect 5396 8707 5397 8747
rect 2475 8698 2517 8707
rect 5355 8698 5397 8707
rect 5835 8747 5877 8756
rect 5835 8707 5836 8747
rect 5876 8707 5877 8747
rect 6298 8716 6307 8756
rect 6347 8716 6356 8756
rect 6298 8715 6356 8716
rect 6411 8756 6453 8765
rect 6411 8716 6412 8756
rect 6452 8716 6453 8756
rect 6411 8707 6453 8716
rect 6795 8756 6837 8765
rect 8619 8756 8661 8765
rect 10443 8756 10485 8765
rect 12250 8756 12308 8757
rect 6795 8716 6796 8756
rect 6836 8716 6837 8756
rect 6795 8707 6837 8716
rect 7371 8747 7413 8756
rect 7371 8707 7372 8747
rect 7412 8707 7413 8747
rect 5835 8698 5877 8707
rect 7371 8698 7413 8707
rect 7851 8747 7893 8756
rect 7851 8707 7852 8747
rect 7892 8707 7893 8747
rect 8619 8716 8620 8756
rect 8660 8716 8661 8756
rect 8619 8707 8661 8716
rect 9867 8747 9909 8756
rect 9867 8707 9868 8747
rect 9908 8707 9909 8747
rect 10443 8716 10444 8756
rect 10484 8716 10485 8756
rect 10443 8707 10485 8716
rect 11691 8747 11733 8756
rect 11691 8707 11692 8747
rect 11732 8707 11733 8747
rect 12250 8716 12259 8756
rect 12299 8716 12308 8756
rect 12250 8715 12308 8716
rect 12363 8756 12405 8765
rect 12363 8716 12364 8756
rect 12404 8716 12405 8756
rect 12363 8707 12405 8716
rect 12747 8756 12789 8765
rect 15802 8756 15860 8757
rect 12747 8716 12748 8756
rect 12788 8716 12789 8756
rect 12747 8707 12789 8716
rect 13323 8747 13365 8756
rect 13323 8707 13324 8747
rect 13364 8707 13365 8747
rect 7851 8698 7893 8707
rect 9867 8698 9909 8707
rect 11691 8698 11733 8707
rect 13323 8698 13365 8707
rect 13803 8747 13845 8756
rect 13803 8707 13804 8747
rect 13844 8707 13845 8747
rect 15802 8716 15811 8756
rect 15851 8716 15860 8756
rect 15802 8715 15860 8716
rect 15915 8756 15957 8765
rect 15915 8716 15916 8756
rect 15956 8716 15957 8756
rect 15915 8707 15957 8716
rect 16299 8756 16341 8765
rect 17739 8756 17781 8765
rect 16299 8716 16300 8756
rect 16340 8716 16341 8756
rect 16299 8707 16341 8716
rect 16875 8747 16917 8756
rect 16875 8707 16876 8747
rect 16916 8707 16917 8747
rect 13803 8698 13845 8707
rect 16875 8698 16917 8707
rect 17355 8747 17397 8756
rect 17355 8707 17356 8747
rect 17396 8707 17397 8747
rect 17739 8716 17740 8756
rect 17780 8716 17781 8756
rect 17739 8707 17781 8716
rect 18987 8747 19029 8756
rect 18987 8707 18988 8747
rect 19028 8707 19029 8747
rect 17355 8698 17397 8707
rect 18987 8698 19029 8707
rect 3051 8672 3093 8681
rect 3051 8632 3052 8672
rect 3092 8632 3093 8672
rect 3051 8623 3093 8632
rect 3243 8672 3285 8681
rect 3243 8632 3244 8672
rect 3284 8632 3285 8672
rect 3243 8623 3285 8632
rect 3483 8672 3525 8681
rect 3483 8632 3484 8672
rect 3524 8632 3525 8672
rect 3483 8623 3525 8632
rect 4011 8672 4053 8681
rect 4011 8632 4012 8672
rect 4052 8632 4053 8672
rect 4011 8623 4053 8632
rect 4875 8672 4917 8681
rect 4875 8632 4876 8672
rect 4916 8632 4917 8672
rect 4875 8623 4917 8632
rect 6058 8672 6116 8673
rect 6058 8632 6067 8672
rect 6107 8632 6116 8672
rect 6058 8631 6116 8632
rect 6891 8672 6933 8681
rect 6891 8632 6892 8672
rect 6932 8632 6933 8672
rect 6891 8623 6933 8632
rect 8074 8672 8132 8673
rect 8074 8632 8083 8672
rect 8123 8632 8132 8672
rect 8074 8631 8132 8632
rect 8427 8672 8469 8681
rect 8427 8632 8428 8672
rect 8468 8632 8469 8672
rect 8427 8623 8469 8632
rect 12843 8672 12885 8681
rect 12843 8632 12844 8672
rect 12884 8632 12885 8672
rect 12843 8623 12885 8632
rect 14859 8672 14901 8681
rect 14859 8632 14860 8672
rect 14900 8632 14901 8672
rect 14859 8623 14901 8632
rect 15531 8672 15573 8681
rect 15531 8632 15532 8672
rect 15572 8632 15573 8672
rect 15531 8623 15573 8632
rect 16395 8672 16437 8681
rect 16395 8632 16396 8672
rect 16436 8632 16437 8672
rect 16395 8623 16437 8632
rect 19323 8672 19365 8681
rect 19323 8632 19324 8672
rect 19364 8632 19365 8672
rect 19323 8623 19365 8632
rect 19563 8672 19605 8681
rect 19563 8632 19564 8672
rect 19604 8632 19605 8672
rect 19563 8623 19605 8632
rect 19947 8672 19989 8681
rect 19947 8632 19948 8672
rect 19988 8632 19989 8672
rect 19947 8623 19989 8632
rect 20331 8672 20373 8681
rect 20331 8632 20332 8672
rect 20372 8632 20373 8672
rect 20331 8623 20373 8632
rect 10059 8504 10101 8513
rect 10059 8464 10060 8504
rect 10100 8464 10101 8504
rect 10059 8455 10101 8464
rect 1152 8336 20448 8360
rect 1152 8296 3688 8336
rect 3728 8296 3770 8336
rect 3810 8296 3852 8336
rect 3892 8296 3934 8336
rect 3974 8296 4016 8336
rect 4056 8296 18808 8336
rect 18848 8296 18890 8336
rect 18930 8296 18972 8336
rect 19012 8296 19054 8336
rect 19094 8296 19136 8336
rect 19176 8296 20448 8336
rect 1152 8272 20448 8296
rect 2859 8168 2901 8177
rect 2859 8128 2860 8168
rect 2900 8128 2901 8168
rect 2859 8119 2901 8128
rect 4491 8168 4533 8177
rect 4491 8128 4492 8168
rect 4532 8128 4533 8168
rect 4491 8119 4533 8128
rect 6219 8168 6261 8177
rect 6219 8128 6220 8168
rect 6260 8128 6261 8168
rect 6219 8119 6261 8128
rect 7947 8168 7989 8177
rect 7947 8128 7948 8168
rect 7988 8128 7989 8168
rect 7947 8119 7989 8128
rect 11787 8168 11829 8177
rect 11787 8128 11788 8168
rect 11828 8128 11829 8168
rect 11787 8119 11829 8128
rect 13803 8168 13845 8177
rect 13803 8128 13804 8168
rect 13844 8128 13845 8168
rect 13803 8119 13845 8128
rect 13995 8168 14037 8177
rect 13995 8128 13996 8168
rect 14036 8128 14037 8168
rect 13995 8119 14037 8128
rect 16155 8168 16197 8177
rect 16155 8128 16156 8168
rect 16196 8128 16197 8168
rect 16155 8119 16197 8128
rect 17739 8168 17781 8177
rect 17739 8128 17740 8168
rect 17780 8128 17781 8168
rect 17739 8119 17781 8128
rect 19947 8168 19989 8177
rect 19947 8128 19948 8168
rect 19988 8128 19989 8168
rect 19947 8119 19989 8128
rect 20091 8084 20133 8093
rect 20091 8044 20092 8084
rect 20132 8044 20133 8084
rect 20091 8035 20133 8044
rect 15915 8000 15957 8009
rect 15915 7960 15916 8000
rect 15956 7960 15957 8000
rect 15915 7951 15957 7960
rect 18123 8000 18165 8009
rect 18123 7960 18124 8000
rect 18164 7960 18165 8000
rect 18123 7951 18165 7960
rect 20331 8000 20373 8009
rect 20331 7960 20332 8000
rect 20372 7960 20373 8000
rect 20331 7951 20373 7960
rect 1419 7916 1461 7925
rect 1419 7876 1420 7916
rect 1460 7876 1461 7916
rect 1419 7867 1461 7876
rect 2659 7916 2717 7917
rect 2659 7876 2668 7916
rect 2708 7876 2717 7916
rect 2659 7875 2717 7876
rect 3051 7916 3093 7925
rect 3051 7876 3052 7916
rect 3092 7876 3093 7916
rect 3051 7867 3093 7876
rect 4291 7916 4349 7917
rect 4291 7876 4300 7916
rect 4340 7876 4349 7916
rect 4291 7875 4349 7876
rect 4779 7916 4821 7925
rect 4779 7876 4780 7916
rect 4820 7876 4821 7916
rect 4779 7867 4821 7876
rect 6019 7916 6077 7917
rect 6019 7876 6028 7916
rect 6068 7876 6077 7916
rect 6019 7875 6077 7876
rect 6507 7916 6549 7925
rect 6507 7876 6508 7916
rect 6548 7876 6549 7916
rect 6507 7867 6549 7876
rect 7747 7916 7805 7917
rect 7747 7876 7756 7916
rect 7796 7876 7805 7916
rect 7747 7875 7805 7876
rect 8619 7916 8661 7925
rect 8619 7876 8620 7916
rect 8660 7876 8661 7916
rect 8619 7867 8661 7876
rect 9859 7916 9917 7917
rect 9859 7876 9868 7916
rect 9908 7876 9917 7916
rect 9859 7875 9917 7876
rect 10347 7916 10389 7925
rect 10347 7876 10348 7916
rect 10388 7876 10389 7916
rect 10347 7867 10389 7876
rect 11587 7916 11645 7917
rect 11587 7876 11596 7916
rect 11636 7876 11645 7916
rect 11587 7875 11645 7876
rect 12363 7916 12405 7925
rect 12363 7876 12364 7916
rect 12404 7876 12405 7916
rect 12363 7867 12405 7876
rect 13603 7916 13661 7917
rect 13603 7876 13612 7916
rect 13652 7876 13661 7916
rect 13603 7875 13661 7876
rect 14179 7916 14237 7917
rect 14179 7876 14188 7916
rect 14228 7876 14237 7916
rect 14179 7875 14237 7876
rect 15435 7916 15477 7925
rect 15435 7876 15436 7916
rect 15476 7876 15477 7916
rect 15435 7867 15477 7876
rect 16299 7916 16341 7925
rect 16299 7876 16300 7916
rect 16340 7876 16341 7916
rect 16299 7867 16341 7876
rect 17539 7916 17597 7917
rect 17539 7876 17548 7916
rect 17588 7876 17597 7916
rect 17539 7875 17597 7876
rect 18507 7916 18549 7925
rect 18507 7876 18508 7916
rect 18548 7876 18549 7916
rect 18507 7867 18549 7876
rect 19747 7916 19805 7917
rect 19747 7876 19756 7916
rect 19796 7876 19805 7916
rect 19747 7875 19805 7876
rect 10059 7748 10101 7757
rect 10059 7708 10060 7748
rect 10100 7708 10101 7748
rect 10059 7699 10101 7708
rect 17883 7748 17925 7757
rect 17883 7708 17884 7748
rect 17924 7708 17925 7748
rect 17883 7699 17925 7708
rect 1152 7580 20452 7604
rect 1152 7540 4928 7580
rect 4968 7540 5010 7580
rect 5050 7540 5092 7580
rect 5132 7540 5174 7580
rect 5214 7540 5256 7580
rect 5296 7540 20048 7580
rect 20088 7540 20130 7580
rect 20170 7540 20212 7580
rect 20252 7540 20294 7580
rect 20334 7540 20376 7580
rect 20416 7540 20452 7580
rect 1152 7516 20452 7540
rect 3819 7412 3861 7421
rect 3819 7372 3820 7412
rect 3860 7372 3861 7412
rect 3819 7363 3861 7372
rect 6699 7412 6741 7421
rect 6699 7372 6700 7412
rect 6740 7372 6741 7412
rect 6699 7363 6741 7372
rect 2379 7244 2421 7253
rect 5259 7244 5301 7253
rect 6987 7244 7029 7253
rect 8698 7244 8756 7245
rect 2379 7204 2380 7244
rect 2420 7204 2421 7244
rect 2379 7195 2421 7204
rect 3627 7235 3669 7244
rect 3627 7195 3628 7235
rect 3668 7195 3669 7235
rect 5259 7204 5260 7244
rect 5300 7204 5301 7244
rect 5259 7195 5301 7204
rect 6507 7235 6549 7244
rect 6507 7195 6508 7235
rect 6548 7195 6549 7235
rect 6987 7204 6988 7244
rect 7028 7204 7029 7244
rect 6987 7195 7029 7204
rect 8235 7235 8277 7244
rect 8235 7195 8236 7235
rect 8276 7195 8277 7235
rect 8698 7204 8707 7244
rect 8747 7204 8756 7244
rect 8698 7203 8756 7204
rect 8811 7244 8853 7253
rect 8811 7204 8812 7244
rect 8852 7204 8853 7244
rect 8811 7195 8853 7204
rect 9195 7244 9237 7253
rect 10635 7244 10677 7253
rect 12843 7244 12885 7253
rect 15915 7244 15957 7253
rect 17547 7244 17589 7253
rect 19179 7244 19221 7253
rect 9195 7204 9196 7244
rect 9236 7204 9237 7244
rect 9195 7195 9237 7204
rect 9771 7235 9813 7244
rect 9771 7195 9772 7235
rect 9812 7195 9813 7235
rect 3627 7186 3669 7195
rect 6507 7186 6549 7195
rect 8235 7186 8277 7195
rect 9771 7186 9813 7195
rect 10251 7235 10293 7244
rect 10251 7195 10252 7235
rect 10292 7195 10293 7235
rect 10635 7204 10636 7244
rect 10676 7204 10677 7244
rect 10635 7195 10677 7204
rect 11883 7235 11925 7244
rect 11883 7195 11884 7235
rect 11924 7195 11925 7235
rect 12843 7204 12844 7244
rect 12884 7204 12885 7244
rect 12843 7195 12885 7204
rect 14091 7235 14133 7244
rect 14091 7195 14092 7235
rect 14132 7195 14133 7235
rect 10251 7186 10293 7195
rect 11883 7186 11925 7195
rect 14091 7186 14133 7195
rect 14667 7235 14709 7244
rect 14667 7195 14668 7235
rect 14708 7195 14709 7235
rect 15915 7204 15916 7244
rect 15956 7204 15957 7244
rect 15915 7195 15957 7204
rect 16299 7235 16341 7244
rect 16299 7195 16300 7235
rect 16340 7195 16341 7235
rect 17547 7204 17548 7244
rect 17588 7204 17589 7244
rect 17547 7195 17589 7204
rect 17931 7235 17973 7244
rect 17931 7195 17932 7235
rect 17972 7195 17973 7235
rect 19179 7204 19180 7244
rect 19220 7204 19221 7244
rect 19179 7195 19221 7204
rect 14667 7186 14709 7195
rect 16299 7186 16341 7195
rect 17931 7186 17973 7195
rect 1179 7160 1221 7169
rect 1179 7120 1180 7160
rect 1220 7120 1221 7160
rect 1179 7111 1221 7120
rect 1419 7160 1461 7169
rect 1419 7120 1420 7160
rect 1460 7120 1461 7160
rect 1419 7111 1461 7120
rect 1803 7160 1845 7169
rect 1803 7120 1804 7160
rect 1844 7120 1845 7160
rect 1803 7111 1845 7120
rect 1947 7160 1989 7169
rect 1947 7120 1948 7160
rect 1988 7120 1989 7160
rect 1947 7111 1989 7120
rect 2187 7160 2229 7169
rect 2187 7120 2188 7160
rect 2228 7120 2229 7160
rect 2187 7111 2229 7120
rect 4203 7160 4245 7169
rect 4203 7120 4204 7160
rect 4244 7120 4245 7160
rect 4203 7111 4245 7120
rect 4587 7160 4629 7169
rect 4587 7120 4588 7160
rect 4628 7120 4629 7160
rect 4587 7111 4629 7120
rect 4971 7160 5013 7169
rect 4971 7120 4972 7160
rect 5012 7120 5013 7160
rect 4971 7111 5013 7120
rect 9291 7160 9333 7169
rect 9291 7120 9292 7160
rect 9332 7120 9333 7160
rect 9291 7111 9333 7120
rect 16090 7160 16148 7161
rect 16090 7120 16099 7160
rect 16139 7120 16148 7160
rect 16090 7119 16148 7120
rect 17722 7160 17780 7161
rect 17722 7120 17731 7160
rect 17771 7120 17780 7160
rect 17722 7119 17780 7120
rect 19659 7160 19701 7169
rect 19659 7120 19660 7160
rect 19700 7120 19701 7160
rect 19659 7111 19701 7120
rect 20331 7160 20373 7169
rect 20331 7120 20332 7160
rect 20372 7120 20373 7160
rect 20331 7111 20373 7120
rect 4347 7076 4389 7085
rect 4347 7036 4348 7076
rect 4388 7036 4389 7076
rect 4347 7027 4389 7036
rect 8427 7076 8469 7085
rect 8427 7036 8428 7076
rect 8468 7036 8469 7076
rect 8427 7027 8469 7036
rect 10491 7076 10533 7085
rect 10491 7036 10492 7076
rect 10532 7036 10533 7076
rect 10491 7027 10533 7036
rect 12075 7076 12117 7085
rect 12075 7036 12076 7076
rect 12116 7036 12117 7076
rect 12075 7027 12117 7036
rect 14283 7076 14325 7085
rect 14283 7036 14284 7076
rect 14324 7036 14325 7076
rect 14283 7027 14325 7036
rect 20091 7076 20133 7085
rect 20091 7036 20092 7076
rect 20132 7036 20133 7076
rect 20091 7027 20133 7036
rect 1563 6992 1605 7001
rect 1563 6952 1564 6992
rect 1604 6952 1605 6992
rect 1563 6943 1605 6952
rect 3963 6992 4005 7001
rect 3963 6952 3964 6992
rect 4004 6952 4005 6992
rect 3963 6943 4005 6952
rect 4731 6992 4773 7001
rect 4731 6952 4732 6992
rect 4772 6952 4773 6992
rect 4731 6943 4773 6952
rect 14475 6992 14517 7001
rect 14475 6952 14476 6992
rect 14516 6952 14517 6992
rect 14475 6943 14517 6952
rect 19419 6992 19461 7001
rect 19419 6952 19420 6992
rect 19460 6952 19461 6992
rect 19419 6943 19461 6952
rect 1152 6824 20448 6848
rect 1152 6784 3688 6824
rect 3728 6784 3770 6824
rect 3810 6784 3852 6824
rect 3892 6784 3934 6824
rect 3974 6784 4016 6824
rect 4056 6784 18808 6824
rect 18848 6784 18890 6824
rect 18930 6784 18972 6824
rect 19012 6784 19054 6824
rect 19094 6784 19136 6824
rect 19176 6784 20448 6824
rect 1152 6760 20448 6784
rect 1179 6656 1221 6665
rect 1179 6616 1180 6656
rect 1220 6616 1221 6656
rect 1179 6607 1221 6616
rect 1563 6656 1605 6665
rect 1563 6616 1564 6656
rect 1604 6616 1605 6656
rect 1563 6607 1605 6616
rect 2811 6656 2853 6665
rect 2811 6616 2812 6656
rect 2852 6616 2853 6656
rect 2811 6607 2853 6616
rect 3195 6656 3237 6665
rect 3195 6616 3196 6656
rect 3236 6616 3237 6656
rect 3195 6607 3237 6616
rect 3915 6656 3957 6665
rect 3915 6616 3916 6656
rect 3956 6616 3957 6656
rect 3915 6607 3957 6616
rect 19755 6656 19797 6665
rect 19755 6616 19756 6656
rect 19796 6616 19797 6656
rect 19755 6607 19797 6616
rect 2331 6572 2373 6581
rect 2331 6532 2332 6572
rect 2372 6532 2373 6572
rect 2331 6523 2373 6532
rect 10299 6572 10341 6581
rect 10299 6532 10300 6572
rect 10340 6532 10341 6572
rect 10299 6523 10341 6532
rect 20091 6572 20133 6581
rect 20091 6532 20092 6572
rect 20132 6532 20133 6572
rect 20091 6523 20133 6532
rect 1419 6488 1461 6497
rect 1419 6448 1420 6488
rect 1460 6448 1461 6488
rect 1419 6439 1461 6448
rect 1803 6488 1845 6497
rect 1803 6448 1804 6488
rect 1844 6448 1845 6488
rect 1803 6439 1845 6448
rect 1995 6488 2037 6497
rect 1995 6448 1996 6488
rect 2036 6448 2037 6488
rect 1995 6439 2037 6448
rect 2571 6488 2613 6497
rect 2571 6448 2572 6488
rect 2612 6448 2613 6488
rect 2571 6439 2613 6448
rect 3051 6488 3093 6497
rect 3051 6448 3052 6488
rect 3092 6448 3093 6488
rect 3051 6439 3093 6448
rect 3435 6488 3477 6497
rect 3435 6448 3436 6488
rect 3476 6448 3477 6488
rect 3435 6439 3477 6448
rect 8907 6488 8949 6497
rect 8907 6448 8908 6488
rect 8948 6448 8949 6488
rect 8907 6439 8949 6448
rect 10539 6488 10581 6497
rect 10539 6448 10540 6488
rect 10580 6448 10581 6488
rect 10539 6439 10581 6448
rect 15051 6488 15093 6497
rect 15051 6448 15052 6488
rect 15092 6448 15093 6488
rect 15051 6439 15093 6448
rect 15915 6488 15957 6497
rect 15915 6448 15916 6488
rect 15956 6448 15957 6488
rect 15915 6439 15957 6448
rect 17194 6488 17252 6489
rect 17194 6448 17203 6488
rect 17243 6448 17252 6488
rect 17194 6447 17252 6448
rect 17547 6488 17589 6497
rect 17547 6448 17548 6488
rect 17588 6448 17589 6488
rect 17547 6439 17589 6448
rect 20331 6488 20373 6497
rect 20331 6448 20332 6488
rect 20372 6448 20373 6488
rect 20331 6439 20373 6448
rect 4099 6404 4157 6405
rect 4099 6364 4108 6404
rect 4148 6364 4157 6404
rect 4099 6363 4157 6364
rect 5355 6404 5397 6413
rect 5355 6364 5356 6404
rect 5396 6364 5397 6404
rect 5355 6355 5397 6364
rect 6507 6404 6549 6413
rect 6507 6364 6508 6404
rect 6548 6364 6549 6404
rect 6507 6355 6549 6364
rect 7747 6404 7805 6405
rect 7747 6364 7756 6404
rect 7796 6364 7805 6404
rect 7747 6363 7805 6364
rect 8410 6404 8468 6405
rect 8410 6364 8419 6404
rect 8459 6364 8468 6404
rect 8410 6363 8468 6364
rect 8523 6404 8565 6413
rect 8523 6364 8524 6404
rect 8564 6364 8565 6404
rect 8523 6355 8565 6364
rect 9003 6404 9045 6413
rect 9003 6364 9004 6404
rect 9044 6364 9045 6404
rect 9003 6355 9045 6364
rect 9478 6404 9536 6405
rect 9478 6364 9487 6404
rect 9527 6364 9536 6404
rect 9478 6363 9536 6364
rect 9963 6404 10021 6405
rect 9963 6364 9972 6404
rect 10012 6364 10021 6404
rect 9963 6363 10021 6364
rect 11115 6404 11157 6413
rect 11115 6364 11116 6404
rect 11156 6364 11157 6404
rect 11115 6355 11157 6364
rect 12355 6404 12413 6405
rect 12355 6364 12364 6404
rect 12404 6364 12413 6404
rect 12355 6363 12413 6364
rect 13227 6404 13269 6413
rect 13227 6364 13228 6404
rect 13268 6364 13269 6404
rect 13227 6355 13269 6364
rect 14467 6404 14525 6405
rect 14467 6364 14476 6404
rect 14516 6364 14525 6404
rect 14467 6363 14525 6364
rect 15405 6404 15447 6413
rect 15405 6364 15406 6404
rect 15446 6364 15447 6404
rect 15405 6355 15447 6364
rect 15531 6404 15573 6413
rect 15531 6364 15532 6404
rect 15572 6364 15573 6404
rect 15531 6355 15573 6364
rect 16011 6404 16053 6413
rect 16011 6364 16012 6404
rect 16052 6364 16053 6404
rect 16011 6355 16053 6364
rect 16483 6404 16541 6405
rect 16483 6364 16492 6404
rect 16532 6364 16541 6404
rect 16483 6363 16541 6364
rect 16971 6404 17029 6405
rect 16971 6364 16980 6404
rect 17020 6364 17029 6404
rect 16971 6363 17029 6364
rect 18315 6404 18357 6413
rect 18315 6364 18316 6404
rect 18356 6364 18357 6404
rect 18315 6355 18357 6364
rect 19555 6404 19613 6405
rect 19555 6364 19564 6404
rect 19604 6364 19613 6404
rect 19555 6363 19613 6364
rect 2235 6320 2277 6329
rect 2235 6280 2236 6320
rect 2276 6280 2277 6320
rect 2235 6271 2277 6280
rect 7947 6236 7989 6245
rect 7947 6196 7948 6236
rect 7988 6196 7989 6236
rect 7947 6187 7989 6196
rect 10155 6236 10197 6245
rect 10155 6196 10156 6236
rect 10196 6196 10197 6236
rect 10155 6187 10197 6196
rect 12555 6236 12597 6245
rect 12555 6196 12556 6236
rect 12596 6196 12597 6236
rect 12555 6187 12597 6196
rect 14667 6236 14709 6245
rect 14667 6196 14668 6236
rect 14708 6196 14709 6236
rect 14667 6187 14709 6196
rect 14811 6236 14853 6245
rect 14811 6196 14812 6236
rect 14852 6196 14853 6236
rect 14811 6187 14853 6196
rect 17307 6236 17349 6245
rect 17307 6196 17308 6236
rect 17348 6196 17349 6236
rect 17307 6187 17349 6196
rect 1152 6068 20452 6092
rect 1152 6028 4928 6068
rect 4968 6028 5010 6068
rect 5050 6028 5092 6068
rect 5132 6028 5174 6068
rect 5214 6028 5256 6068
rect 5296 6028 20048 6068
rect 20088 6028 20130 6068
rect 20170 6028 20212 6068
rect 20252 6028 20294 6068
rect 20334 6028 20376 6068
rect 20416 6028 20452 6068
rect 1152 6004 20452 6028
rect 14667 5900 14709 5909
rect 14667 5860 14668 5900
rect 14708 5860 14709 5900
rect 14667 5851 14709 5860
rect 16299 5900 16341 5909
rect 16299 5860 16300 5900
rect 16340 5860 16341 5900
rect 16299 5851 16341 5860
rect 16491 5900 16533 5909
rect 16491 5860 16492 5900
rect 16532 5860 16533 5900
rect 16491 5851 16533 5860
rect 2331 5816 2373 5825
rect 2331 5776 2332 5816
rect 2372 5776 2373 5816
rect 2331 5767 2373 5776
rect 5259 5732 5301 5741
rect 6891 5732 6933 5741
rect 8523 5732 8565 5741
rect 10906 5732 10964 5733
rect 5259 5692 5260 5732
rect 5300 5692 5301 5732
rect 5259 5683 5301 5692
rect 6507 5723 6549 5732
rect 6507 5683 6508 5723
rect 6548 5683 6549 5723
rect 6891 5692 6892 5732
rect 6932 5692 6933 5732
rect 6891 5683 6933 5692
rect 8139 5723 8181 5732
rect 8139 5683 8140 5723
rect 8180 5683 8181 5723
rect 8523 5692 8524 5732
rect 8564 5692 8565 5732
rect 8523 5683 8565 5692
rect 9771 5723 9813 5732
rect 9771 5683 9772 5723
rect 9812 5683 9813 5723
rect 10906 5692 10915 5732
rect 10955 5692 10964 5732
rect 10906 5691 10964 5692
rect 11019 5732 11061 5741
rect 11019 5692 11020 5732
rect 11060 5692 11061 5732
rect 11019 5683 11061 5692
rect 11403 5732 11445 5741
rect 12922 5732 12980 5733
rect 11403 5692 11404 5732
rect 11444 5692 11445 5732
rect 11403 5683 11445 5692
rect 11979 5723 12021 5732
rect 11979 5683 11980 5723
rect 12020 5683 12021 5723
rect 6507 5674 6549 5683
rect 8139 5674 8181 5683
rect 9771 5674 9813 5683
rect 11979 5674 12021 5683
rect 12459 5723 12501 5732
rect 12459 5683 12460 5723
rect 12500 5683 12501 5723
rect 12922 5692 12931 5732
rect 12971 5692 12980 5732
rect 12922 5691 12980 5692
rect 13035 5732 13077 5741
rect 13035 5692 13036 5732
rect 13076 5692 13077 5732
rect 13035 5683 13077 5692
rect 13419 5732 13461 5741
rect 14859 5732 14901 5741
rect 17931 5732 17973 5741
rect 13419 5692 13420 5732
rect 13460 5692 13461 5732
rect 13419 5683 13461 5692
rect 13995 5723 14037 5732
rect 13995 5683 13996 5723
rect 14036 5683 14037 5723
rect 12459 5674 12501 5683
rect 13995 5674 14037 5683
rect 14475 5723 14517 5732
rect 14475 5683 14476 5723
rect 14516 5683 14517 5723
rect 14859 5692 14860 5732
rect 14900 5692 14901 5732
rect 14859 5683 14901 5692
rect 16107 5723 16149 5732
rect 16107 5683 16108 5723
rect 16148 5683 16149 5723
rect 14475 5674 14517 5683
rect 16107 5674 16149 5683
rect 16683 5723 16725 5732
rect 16683 5683 16684 5723
rect 16724 5683 16725 5723
rect 17931 5692 17932 5732
rect 17972 5692 17973 5732
rect 17931 5683 17973 5692
rect 16683 5674 16725 5683
rect 1179 5648 1221 5657
rect 1179 5608 1180 5648
rect 1220 5608 1221 5648
rect 1179 5599 1221 5608
rect 1419 5648 1461 5657
rect 1419 5608 1420 5648
rect 1460 5608 1461 5648
rect 1419 5599 1461 5608
rect 1803 5648 1845 5657
rect 1803 5608 1804 5648
rect 1844 5608 1845 5648
rect 1803 5599 1845 5608
rect 2187 5648 2229 5657
rect 2187 5608 2188 5648
rect 2228 5608 2229 5648
rect 2187 5599 2229 5608
rect 2571 5648 2613 5657
rect 2571 5608 2572 5648
rect 2612 5608 2613 5648
rect 2571 5599 2613 5608
rect 2763 5648 2805 5657
rect 2763 5608 2764 5648
rect 2804 5608 2805 5648
rect 2763 5599 2805 5608
rect 3339 5648 3381 5657
rect 3339 5608 3340 5648
rect 3380 5608 3381 5648
rect 3339 5599 3381 5608
rect 4299 5648 4341 5657
rect 4299 5608 4300 5648
rect 4340 5608 4341 5648
rect 4299 5599 4341 5608
rect 4683 5648 4725 5657
rect 4683 5608 4684 5648
rect 4724 5608 4725 5648
rect 4683 5599 4725 5608
rect 4923 5648 4965 5657
rect 4923 5608 4924 5648
rect 4964 5608 4965 5648
rect 4923 5599 4965 5608
rect 10347 5648 10389 5657
rect 10347 5608 10348 5648
rect 10388 5608 10389 5648
rect 10347 5599 10389 5608
rect 11499 5648 11541 5657
rect 11499 5608 11500 5648
rect 11540 5608 11541 5648
rect 11499 5599 11541 5608
rect 13515 5648 13557 5657
rect 13515 5608 13516 5648
rect 13556 5608 13557 5648
rect 13515 5599 13557 5608
rect 18939 5648 18981 5657
rect 18939 5608 18940 5648
rect 18980 5608 18981 5648
rect 18939 5599 18981 5608
rect 19179 5648 19221 5657
rect 19179 5608 19180 5648
rect 19220 5608 19221 5648
rect 19179 5599 19221 5608
rect 19563 5648 19605 5657
rect 19563 5608 19564 5648
rect 19604 5608 19605 5648
rect 19563 5599 19605 5608
rect 19947 5648 19989 5657
rect 19947 5608 19948 5648
rect 19988 5608 19989 5648
rect 19947 5599 19989 5608
rect 20331 5648 20373 5657
rect 20331 5608 20332 5648
rect 20372 5608 20373 5648
rect 20331 5599 20373 5608
rect 3003 5564 3045 5573
rect 3003 5524 3004 5564
rect 3044 5524 3045 5564
rect 3003 5515 3045 5524
rect 8331 5564 8373 5573
rect 8331 5524 8332 5564
rect 8372 5524 8373 5564
rect 8331 5515 8373 5524
rect 19707 5564 19749 5573
rect 19707 5524 19708 5564
rect 19748 5524 19749 5564
rect 19707 5515 19749 5524
rect 1563 5480 1605 5489
rect 1563 5440 1564 5480
rect 1604 5440 1605 5480
rect 1563 5431 1605 5440
rect 1947 5480 1989 5489
rect 1947 5440 1948 5480
rect 1988 5440 1989 5480
rect 1947 5431 1989 5440
rect 3099 5480 3141 5489
rect 3099 5440 3100 5480
rect 3140 5440 3141 5480
rect 3099 5431 3141 5440
rect 4539 5480 4581 5489
rect 4539 5440 4540 5480
rect 4580 5440 4581 5480
rect 4539 5431 4581 5440
rect 6699 5480 6741 5489
rect 6699 5440 6700 5480
rect 6740 5440 6741 5480
rect 6699 5431 6741 5440
rect 9963 5480 10005 5489
rect 9963 5440 9964 5480
rect 10004 5440 10005 5480
rect 9963 5431 10005 5440
rect 10107 5480 10149 5489
rect 10107 5440 10108 5480
rect 10148 5440 10149 5480
rect 10107 5431 10149 5440
rect 12682 5480 12740 5481
rect 12682 5440 12691 5480
rect 12731 5440 12740 5480
rect 12682 5439 12740 5440
rect 19323 5480 19365 5489
rect 19323 5440 19324 5480
rect 19364 5440 19365 5480
rect 19323 5431 19365 5440
rect 20091 5480 20133 5489
rect 20091 5440 20092 5480
rect 20132 5440 20133 5480
rect 20091 5431 20133 5440
rect 1152 5312 20448 5336
rect 1152 5272 3688 5312
rect 3728 5272 3770 5312
rect 3810 5272 3852 5312
rect 3892 5272 3934 5312
rect 3974 5272 4016 5312
rect 4056 5272 18808 5312
rect 18848 5272 18890 5312
rect 18930 5272 18972 5312
rect 19012 5272 19054 5312
rect 19094 5272 19136 5312
rect 19176 5272 20448 5312
rect 1152 5248 20448 5272
rect 1179 5144 1221 5153
rect 1179 5104 1180 5144
rect 1220 5104 1221 5144
rect 1179 5095 1221 5104
rect 1563 5144 1605 5153
rect 1563 5104 1564 5144
rect 1604 5104 1605 5144
rect 1563 5095 1605 5104
rect 8043 5144 8085 5153
rect 8043 5104 8044 5144
rect 8084 5104 8085 5144
rect 8043 5095 8085 5104
rect 10539 5144 10581 5153
rect 10539 5104 10540 5144
rect 10580 5104 10581 5144
rect 10539 5095 10581 5104
rect 13083 5144 13125 5153
rect 13083 5104 13084 5144
rect 13124 5104 13125 5144
rect 13083 5095 13125 5104
rect 15867 5144 15909 5153
rect 15867 5104 15868 5144
rect 15908 5104 15909 5144
rect 15867 5095 15909 5104
rect 19323 5144 19365 5153
rect 19323 5104 19324 5144
rect 19364 5104 19365 5144
rect 19323 5095 19365 5104
rect 20091 5144 20133 5153
rect 20091 5104 20092 5144
rect 20132 5104 20133 5144
rect 20091 5095 20133 5104
rect 2331 5060 2373 5069
rect 2331 5020 2332 5060
rect 2372 5020 2373 5060
rect 2331 5011 2373 5020
rect 19707 5060 19749 5069
rect 19707 5020 19708 5060
rect 19748 5020 19749 5060
rect 19707 5011 19749 5020
rect 1419 4976 1461 4985
rect 1419 4936 1420 4976
rect 1460 4936 1461 4976
rect 1419 4927 1461 4936
rect 1803 4976 1845 4985
rect 1803 4936 1804 4976
rect 1844 4936 1845 4976
rect 1803 4927 1845 4936
rect 2187 4976 2229 4985
rect 2187 4936 2188 4976
rect 2228 4936 2229 4976
rect 2187 4927 2229 4936
rect 2571 4976 2613 4985
rect 2571 4936 2572 4976
rect 2612 4936 2613 4976
rect 2571 4927 2613 4936
rect 2955 4976 2997 4985
rect 2955 4936 2956 4976
rect 2996 4936 2997 4976
rect 2955 4927 2997 4936
rect 11307 4976 11349 4985
rect 11307 4936 11308 4976
rect 11348 4936 11349 4976
rect 11307 4927 11349 4936
rect 12586 4976 12644 4977
rect 12586 4936 12595 4976
rect 12635 4936 12644 4976
rect 12586 4935 12644 4936
rect 12939 4976 12981 4985
rect 12939 4936 12940 4976
rect 12980 4936 12981 4976
rect 12939 4927 12981 4936
rect 13323 4976 13365 4985
rect 13323 4936 13324 4976
rect 13364 4936 13365 4976
rect 13323 4927 13365 4936
rect 14475 4976 14517 4985
rect 14475 4936 14476 4976
rect 14516 4936 14517 4976
rect 14475 4927 14517 4936
rect 15754 4976 15812 4977
rect 15754 4936 15763 4976
rect 15803 4936 15812 4976
rect 15754 4935 15812 4936
rect 16107 4976 16149 4985
rect 16107 4936 16108 4976
rect 16148 4936 16149 4976
rect 16107 4927 16149 4936
rect 19563 4976 19605 4985
rect 19563 4936 19564 4976
rect 19604 4936 19605 4976
rect 19563 4927 19605 4936
rect 19947 4976 19989 4985
rect 19947 4936 19948 4976
rect 19988 4936 19989 4976
rect 19947 4927 19989 4936
rect 20331 4976 20373 4985
rect 20331 4936 20332 4976
rect 20372 4936 20373 4976
rect 20331 4927 20373 4936
rect 6603 4892 6645 4901
rect 6603 4852 6604 4892
rect 6644 4852 6645 4892
rect 6603 4843 6645 4852
rect 7843 4892 7901 4893
rect 7843 4852 7852 4892
rect 7892 4852 7901 4892
rect 7843 4851 7901 4852
rect 9099 4892 9141 4901
rect 9099 4852 9100 4892
rect 9140 4852 9141 4892
rect 9099 4843 9141 4852
rect 10339 4892 10397 4893
rect 10339 4852 10348 4892
rect 10388 4852 10397 4892
rect 10339 4851 10397 4852
rect 10810 4892 10868 4893
rect 10810 4852 10819 4892
rect 10859 4852 10868 4892
rect 10810 4851 10868 4852
rect 10923 4892 10965 4901
rect 10923 4852 10924 4892
rect 10964 4852 10965 4892
rect 10923 4843 10965 4852
rect 11403 4892 11445 4901
rect 11403 4852 11404 4892
rect 11444 4852 11445 4892
rect 11403 4843 11445 4852
rect 11875 4892 11933 4893
rect 11875 4852 11884 4892
rect 11924 4852 11933 4892
rect 11875 4851 11933 4852
rect 12363 4892 12421 4893
rect 12363 4852 12372 4892
rect 12412 4852 12421 4892
rect 12363 4851 12421 4852
rect 13978 4892 14036 4893
rect 13978 4852 13987 4892
rect 14027 4852 14036 4892
rect 13978 4851 14036 4852
rect 14091 4892 14133 4901
rect 14091 4852 14092 4892
rect 14132 4852 14133 4892
rect 14091 4843 14133 4852
rect 14571 4892 14613 4901
rect 14571 4852 14572 4892
rect 14612 4852 14613 4892
rect 14571 4843 14613 4852
rect 15043 4892 15101 4893
rect 15043 4852 15052 4892
rect 15092 4852 15101 4892
rect 15043 4851 15101 4852
rect 15562 4892 15620 4893
rect 15562 4852 15571 4892
rect 15611 4852 15620 4892
rect 15562 4851 15620 4852
rect 2715 4808 2757 4817
rect 2715 4768 2716 4808
rect 2756 4768 2757 4808
rect 2715 4759 2757 4768
rect 1947 4724 1989 4733
rect 1947 4684 1948 4724
rect 1988 4684 1989 4724
rect 1947 4675 1989 4684
rect 12699 4724 12741 4733
rect 12699 4684 12700 4724
rect 12740 4684 12741 4724
rect 12699 4675 12741 4684
rect 1152 4556 20452 4580
rect 1152 4516 4928 4556
rect 4968 4516 5010 4556
rect 5050 4516 5092 4556
rect 5132 4516 5174 4556
rect 5214 4516 5256 4556
rect 5296 4516 20048 4556
rect 20088 4516 20130 4556
rect 20170 4516 20212 4556
rect 20252 4516 20294 4556
rect 20334 4516 20376 4556
rect 20416 4516 20452 4556
rect 1152 4492 20452 4516
rect 1179 4304 1221 4313
rect 1179 4264 1180 4304
rect 1220 4264 1221 4304
rect 1179 4255 1221 4264
rect 1563 4304 1605 4313
rect 1563 4264 1564 4304
rect 1604 4264 1605 4304
rect 1563 4255 1605 4264
rect 19707 4304 19749 4313
rect 19707 4264 19708 4304
rect 19748 4264 19749 4304
rect 19707 4255 19749 4264
rect 10923 4220 10965 4229
rect 10923 4180 10924 4220
rect 10964 4180 10965 4220
rect 10923 4171 10965 4180
rect 12171 4211 12213 4220
rect 12171 4171 12172 4211
rect 12212 4171 12213 4211
rect 12171 4162 12213 4171
rect 1419 4136 1461 4145
rect 1419 4096 1420 4136
rect 1460 4096 1461 4136
rect 1419 4087 1461 4096
rect 1803 4136 1845 4145
rect 1803 4096 1804 4136
rect 1844 4096 1845 4136
rect 1803 4087 1845 4096
rect 2187 4136 2229 4145
rect 2187 4096 2188 4136
rect 2228 4096 2229 4136
rect 2187 4087 2229 4096
rect 2571 4136 2613 4145
rect 2571 4096 2572 4136
rect 2612 4096 2613 4136
rect 2571 4087 2613 4096
rect 2763 4136 2805 4145
rect 2763 4096 2764 4136
rect 2804 4096 2805 4136
rect 2763 4087 2805 4096
rect 19947 4136 19989 4145
rect 19947 4096 19948 4136
rect 19988 4096 19989 4136
rect 19947 4087 19989 4096
rect 20331 4136 20373 4145
rect 20331 4096 20332 4136
rect 20372 4096 20373 4136
rect 20331 4087 20373 4096
rect 3003 4052 3045 4061
rect 3003 4012 3004 4052
rect 3044 4012 3045 4052
rect 3003 4003 3045 4012
rect 20091 4052 20133 4061
rect 20091 4012 20092 4052
rect 20132 4012 20133 4052
rect 20091 4003 20133 4012
rect 1947 3968 1989 3977
rect 1947 3928 1948 3968
rect 1988 3928 1989 3968
rect 1947 3919 1989 3928
rect 2331 3968 2373 3977
rect 2331 3928 2332 3968
rect 2372 3928 2373 3968
rect 2331 3919 2373 3928
rect 12363 3968 12405 3977
rect 12363 3928 12364 3968
rect 12404 3928 12405 3968
rect 12363 3919 12405 3928
rect 1152 3800 20448 3824
rect 1152 3760 3688 3800
rect 3728 3760 3770 3800
rect 3810 3760 3852 3800
rect 3892 3760 3934 3800
rect 3974 3760 4016 3800
rect 4056 3760 18808 3800
rect 18848 3760 18890 3800
rect 18930 3760 18972 3800
rect 19012 3760 19054 3800
rect 19094 3760 19136 3800
rect 19176 3760 20448 3800
rect 1152 3736 20448 3760
rect 1179 3632 1221 3641
rect 1179 3592 1180 3632
rect 1220 3592 1221 3632
rect 1179 3583 1221 3592
rect 1563 3632 1605 3641
rect 1563 3592 1564 3632
rect 1604 3592 1605 3632
rect 1563 3583 1605 3592
rect 3771 3632 3813 3641
rect 3771 3592 3772 3632
rect 3812 3592 3813 3632
rect 3771 3583 3813 3592
rect 3387 3548 3429 3557
rect 3387 3508 3388 3548
rect 3428 3508 3429 3548
rect 3387 3499 3429 3508
rect 1419 3464 1461 3473
rect 1419 3424 1420 3464
rect 1460 3424 1461 3464
rect 1419 3415 1461 3424
rect 1803 3464 1845 3473
rect 1803 3424 1804 3464
rect 1844 3424 1845 3464
rect 1803 3415 1845 3424
rect 2187 3464 2229 3473
rect 2187 3424 2188 3464
rect 2228 3424 2229 3464
rect 2187 3415 2229 3424
rect 2379 3464 2421 3473
rect 2379 3424 2380 3464
rect 2420 3424 2421 3464
rect 2379 3415 2421 3424
rect 2955 3464 2997 3473
rect 2955 3424 2956 3464
rect 2996 3424 2997 3464
rect 2955 3415 2997 3424
rect 3147 3464 3189 3473
rect 3147 3424 3148 3464
rect 3188 3424 3189 3464
rect 3147 3415 3189 3424
rect 3531 3464 3573 3473
rect 3531 3424 3532 3464
rect 3572 3424 3573 3464
rect 3531 3415 3573 3424
rect 20331 3464 20373 3473
rect 20331 3424 20332 3464
rect 20372 3424 20373 3464
rect 20331 3415 20373 3424
rect 1947 3296 1989 3305
rect 1947 3256 1948 3296
rect 1988 3256 1989 3296
rect 1947 3247 1989 3256
rect 2619 3296 2661 3305
rect 2619 3256 2620 3296
rect 2660 3256 2661 3296
rect 2619 3247 2661 3256
rect 2715 3212 2757 3221
rect 2715 3172 2716 3212
rect 2756 3172 2757 3212
rect 2715 3163 2757 3172
rect 20091 3212 20133 3221
rect 20091 3172 20092 3212
rect 20132 3172 20133 3212
rect 20091 3163 20133 3172
rect 1152 3044 20452 3068
rect 1152 3004 4928 3044
rect 4968 3004 5010 3044
rect 5050 3004 5092 3044
rect 5132 3004 5174 3044
rect 5214 3004 5256 3044
rect 5296 3004 20048 3044
rect 20088 3004 20130 3044
rect 20170 3004 20212 3044
rect 20252 3004 20294 3044
rect 20334 3004 20376 3044
rect 20416 3004 20452 3044
rect 1152 2980 20452 3004
rect 1179 2876 1221 2885
rect 1179 2836 1180 2876
rect 1220 2836 1221 2876
rect 1179 2827 1221 2836
rect 3867 2876 3909 2885
rect 3867 2836 3868 2876
rect 3908 2836 3909 2876
rect 3867 2827 3909 2836
rect 4251 2876 4293 2885
rect 4251 2836 4252 2876
rect 4292 2836 4293 2876
rect 4251 2827 4293 2836
rect 4635 2876 4677 2885
rect 4635 2836 4636 2876
rect 4676 2836 4677 2876
rect 4635 2827 4677 2836
rect 5787 2876 5829 2885
rect 5787 2836 5788 2876
rect 5828 2836 5829 2876
rect 5787 2827 5829 2836
rect 6171 2876 6213 2885
rect 6171 2836 6172 2876
rect 6212 2836 6213 2876
rect 6171 2827 6213 2836
rect 8475 2876 8517 2885
rect 8475 2836 8476 2876
rect 8516 2836 8517 2876
rect 8475 2827 8517 2836
rect 3483 2792 3525 2801
rect 3483 2752 3484 2792
rect 3524 2752 3525 2792
rect 3483 2743 3525 2752
rect 5019 2792 5061 2801
rect 5019 2752 5020 2792
rect 5060 2752 5061 2792
rect 5019 2743 5061 2752
rect 1419 2624 1461 2633
rect 1419 2584 1420 2624
rect 1460 2584 1461 2624
rect 1419 2575 1461 2584
rect 1707 2624 1749 2633
rect 1707 2584 1708 2624
rect 1748 2584 1749 2624
rect 1707 2575 1749 2584
rect 2091 2624 2133 2633
rect 2091 2584 2092 2624
rect 2132 2584 2133 2624
rect 2091 2575 2133 2584
rect 2571 2624 2613 2633
rect 2571 2584 2572 2624
rect 2612 2584 2613 2624
rect 2571 2575 2613 2584
rect 2811 2624 2853 2633
rect 2811 2584 2812 2624
rect 2852 2584 2853 2624
rect 2811 2575 2853 2584
rect 3243 2624 3285 2633
rect 3243 2584 3244 2624
rect 3284 2584 3285 2624
rect 3243 2575 3285 2584
rect 3627 2624 3669 2633
rect 3627 2584 3628 2624
rect 3668 2584 3669 2624
rect 3627 2575 3669 2584
rect 4011 2624 4053 2633
rect 4011 2584 4012 2624
rect 4052 2584 4053 2624
rect 4011 2575 4053 2584
rect 4395 2624 4437 2633
rect 4395 2584 4396 2624
rect 4436 2584 4437 2624
rect 4395 2575 4437 2584
rect 4779 2624 4821 2633
rect 4779 2584 4780 2624
rect 4820 2584 4821 2624
rect 4779 2575 4821 2584
rect 5163 2624 5205 2633
rect 5163 2584 5164 2624
rect 5204 2584 5205 2624
rect 5163 2575 5205 2584
rect 5547 2624 5589 2633
rect 5547 2584 5548 2624
rect 5588 2584 5589 2624
rect 5547 2575 5589 2584
rect 5931 2624 5973 2633
rect 5931 2584 5932 2624
rect 5972 2584 5973 2624
rect 5931 2575 5973 2584
rect 8235 2624 8277 2633
rect 8235 2584 8236 2624
rect 8276 2584 8277 2624
rect 8235 2575 8277 2584
rect 9195 2624 9237 2633
rect 9195 2584 9196 2624
rect 9236 2584 9237 2624
rect 9195 2575 9237 2584
rect 9579 2624 9621 2633
rect 9579 2584 9580 2624
rect 9620 2584 9621 2624
rect 9579 2575 9621 2584
rect 9963 2624 10005 2633
rect 9963 2584 9964 2624
rect 10004 2584 10005 2624
rect 9963 2575 10005 2584
rect 10347 2624 10389 2633
rect 10347 2584 10348 2624
rect 10388 2584 10389 2624
rect 10347 2575 10389 2584
rect 10731 2624 10773 2633
rect 10731 2584 10732 2624
rect 10772 2584 10773 2624
rect 10731 2575 10773 2584
rect 11115 2624 11157 2633
rect 11115 2584 11116 2624
rect 11156 2584 11157 2624
rect 11115 2575 11157 2584
rect 12843 2624 12885 2633
rect 12843 2584 12844 2624
rect 12884 2584 12885 2624
rect 12843 2575 12885 2584
rect 13227 2624 13269 2633
rect 13227 2584 13228 2624
rect 13268 2584 13269 2624
rect 13227 2575 13269 2584
rect 13611 2624 13653 2633
rect 13611 2584 13612 2624
rect 13652 2584 13653 2624
rect 13611 2575 13653 2584
rect 13995 2624 14037 2633
rect 13995 2584 13996 2624
rect 14036 2584 14037 2624
rect 13995 2575 14037 2584
rect 14379 2624 14421 2633
rect 14379 2584 14380 2624
rect 14420 2584 14421 2624
rect 14379 2575 14421 2584
rect 14763 2624 14805 2633
rect 14763 2584 14764 2624
rect 14804 2584 14805 2624
rect 14763 2575 14805 2584
rect 15147 2624 15189 2633
rect 15147 2584 15148 2624
rect 15188 2584 15189 2624
rect 15147 2575 15189 2584
rect 15531 2624 15573 2633
rect 15531 2584 15532 2624
rect 15572 2584 15573 2624
rect 15531 2575 15573 2584
rect 1947 2540 1989 2549
rect 1947 2500 1948 2540
rect 1988 2500 1989 2540
rect 1947 2491 1989 2500
rect 2331 2456 2373 2465
rect 2331 2416 2332 2456
rect 2372 2416 2373 2456
rect 2331 2407 2373 2416
rect 5403 2456 5445 2465
rect 5403 2416 5404 2456
rect 5444 2416 5445 2456
rect 5403 2407 5445 2416
rect 8955 2456 8997 2465
rect 8955 2416 8956 2456
rect 8996 2416 8997 2456
rect 8955 2407 8997 2416
rect 9339 2456 9381 2465
rect 9339 2416 9340 2456
rect 9380 2416 9381 2456
rect 9339 2407 9381 2416
rect 9723 2456 9765 2465
rect 9723 2416 9724 2456
rect 9764 2416 9765 2456
rect 9723 2407 9765 2416
rect 10107 2456 10149 2465
rect 10107 2416 10108 2456
rect 10148 2416 10149 2456
rect 10107 2407 10149 2416
rect 10491 2456 10533 2465
rect 10491 2416 10492 2456
rect 10532 2416 10533 2456
rect 10491 2407 10533 2416
rect 10875 2456 10917 2465
rect 10875 2416 10876 2456
rect 10916 2416 10917 2456
rect 10875 2407 10917 2416
rect 12603 2456 12645 2465
rect 12603 2416 12604 2456
rect 12644 2416 12645 2456
rect 12603 2407 12645 2416
rect 12987 2456 13029 2465
rect 12987 2416 12988 2456
rect 13028 2416 13029 2456
rect 12987 2407 13029 2416
rect 13371 2456 13413 2465
rect 13371 2416 13372 2456
rect 13412 2416 13413 2456
rect 13371 2407 13413 2416
rect 13755 2456 13797 2465
rect 13755 2416 13756 2456
rect 13796 2416 13797 2456
rect 13755 2407 13797 2416
rect 14139 2456 14181 2465
rect 14139 2416 14140 2456
rect 14180 2416 14181 2456
rect 14139 2407 14181 2416
rect 14523 2456 14565 2465
rect 14523 2416 14524 2456
rect 14564 2416 14565 2456
rect 14523 2407 14565 2416
rect 14907 2456 14949 2465
rect 14907 2416 14908 2456
rect 14948 2416 14949 2456
rect 14907 2407 14949 2416
rect 15291 2456 15333 2465
rect 15291 2416 15292 2456
rect 15332 2416 15333 2456
rect 15291 2407 15333 2416
rect 1152 2288 20448 2312
rect 1152 2248 3688 2288
rect 3728 2248 3770 2288
rect 3810 2248 3852 2288
rect 3892 2248 3934 2288
rect 3974 2248 4016 2288
rect 4056 2248 18808 2288
rect 18848 2248 18890 2288
rect 18930 2248 18972 2288
rect 19012 2248 19054 2288
rect 19094 2248 19136 2288
rect 19176 2248 20448 2288
rect 1152 2224 20448 2248
rect 1947 2120 1989 2129
rect 1947 2080 1948 2120
rect 1988 2080 1989 2120
rect 1947 2071 1989 2080
rect 2811 2120 2853 2129
rect 2811 2080 2812 2120
rect 2852 2080 2853 2120
rect 2811 2071 2853 2080
rect 3867 2120 3909 2129
rect 3867 2080 3868 2120
rect 3908 2080 3909 2120
rect 3867 2071 3909 2080
rect 4251 2120 4293 2129
rect 4251 2080 4252 2120
rect 4292 2080 4293 2120
rect 4251 2071 4293 2080
rect 5019 2120 5061 2129
rect 5019 2080 5020 2120
rect 5060 2080 5061 2120
rect 5019 2071 5061 2080
rect 6171 2120 6213 2129
rect 6171 2080 6172 2120
rect 6212 2080 6213 2120
rect 6171 2071 6213 2080
rect 6555 2120 6597 2129
rect 6555 2080 6556 2120
rect 6596 2080 6597 2120
rect 6555 2071 6597 2080
rect 7035 2120 7077 2129
rect 7035 2080 7036 2120
rect 7076 2080 7077 2120
rect 7035 2071 7077 2080
rect 7707 2120 7749 2129
rect 7707 2080 7708 2120
rect 7748 2080 7749 2120
rect 7707 2071 7749 2080
rect 17403 2120 17445 2129
rect 17403 2080 17404 2120
rect 17444 2080 17445 2120
rect 17403 2071 17445 2080
rect 4347 2036 4389 2045
rect 4347 1996 4348 2036
rect 4388 1996 4389 2036
rect 4347 1987 4389 1996
rect 6939 2036 6981 2045
rect 6939 1996 6940 2036
rect 6980 1996 6981 2036
rect 6939 1987 6981 1996
rect 14715 2036 14757 2045
rect 14715 1996 14716 2036
rect 14756 1996 14757 2036
rect 14715 1987 14757 1996
rect 1323 1952 1365 1961
rect 1323 1912 1324 1952
rect 1364 1912 1365 1952
rect 1323 1903 1365 1912
rect 1707 1952 1749 1961
rect 1707 1912 1708 1952
rect 1748 1912 1749 1952
rect 1707 1903 1749 1912
rect 2091 1952 2133 1961
rect 2091 1912 2092 1952
rect 2132 1912 2133 1952
rect 2091 1903 2133 1912
rect 2475 1952 2517 1961
rect 2475 1912 2476 1952
rect 2516 1912 2517 1952
rect 2475 1903 2517 1912
rect 3051 1952 3093 1961
rect 3051 1912 3052 1952
rect 3092 1912 3093 1952
rect 3051 1903 3093 1912
rect 3243 1952 3285 1961
rect 3243 1912 3244 1952
rect 3284 1912 3285 1952
rect 3243 1903 3285 1912
rect 3627 1952 3669 1961
rect 3627 1912 3628 1952
rect 3668 1912 3669 1952
rect 3627 1903 3669 1912
rect 4011 1952 4053 1961
rect 4011 1912 4012 1952
rect 4052 1912 4053 1952
rect 4011 1903 4053 1912
rect 4587 1952 4629 1961
rect 4587 1912 4588 1952
rect 4628 1912 4629 1952
rect 4587 1903 4629 1912
rect 4779 1952 4821 1961
rect 4779 1912 4780 1952
rect 4820 1912 4821 1952
rect 4779 1903 4821 1912
rect 5163 1952 5205 1961
rect 5163 1912 5164 1952
rect 5204 1912 5205 1952
rect 5163 1903 5205 1912
rect 5547 1952 5589 1961
rect 5547 1912 5548 1952
rect 5588 1912 5589 1952
rect 5547 1903 5589 1912
rect 5931 1952 5973 1961
rect 5931 1912 5932 1952
rect 5972 1912 5973 1952
rect 5931 1903 5973 1912
rect 6315 1952 6357 1961
rect 6315 1912 6316 1952
rect 6356 1912 6357 1952
rect 6315 1903 6357 1912
rect 6699 1952 6741 1961
rect 6699 1912 6700 1952
rect 6740 1912 6741 1952
rect 6699 1903 6741 1912
rect 7275 1952 7317 1961
rect 7275 1912 7276 1952
rect 7316 1912 7317 1952
rect 7275 1903 7317 1912
rect 7467 1952 7509 1961
rect 7467 1912 7468 1952
rect 7508 1912 7509 1952
rect 7467 1903 7509 1912
rect 8235 1952 8277 1961
rect 8235 1912 8236 1952
rect 8276 1912 8277 1952
rect 8235 1903 8277 1912
rect 8619 1952 8661 1961
rect 8619 1912 8620 1952
rect 8660 1912 8661 1952
rect 8619 1903 8661 1912
rect 9003 1952 9045 1961
rect 9003 1912 9004 1952
rect 9044 1912 9045 1952
rect 9003 1903 9045 1912
rect 9387 1952 9429 1961
rect 9387 1912 9388 1952
rect 9428 1912 9429 1952
rect 9387 1903 9429 1912
rect 9771 1952 9813 1961
rect 9771 1912 9772 1952
rect 9812 1912 9813 1952
rect 9771 1903 9813 1912
rect 10155 1952 10197 1961
rect 10155 1912 10156 1952
rect 10196 1912 10197 1952
rect 10155 1903 10197 1912
rect 10539 1952 10581 1961
rect 10539 1912 10540 1952
rect 10580 1912 10581 1952
rect 10539 1903 10581 1912
rect 10923 1952 10965 1961
rect 10923 1912 10924 1952
rect 10964 1912 10965 1952
rect 10923 1903 10965 1912
rect 11499 1952 11541 1961
rect 11499 1912 11500 1952
rect 11540 1912 11541 1952
rect 11499 1903 11541 1912
rect 11883 1952 11925 1961
rect 11883 1912 11884 1952
rect 11924 1912 11925 1952
rect 11883 1903 11925 1912
rect 12267 1952 12309 1961
rect 12267 1912 12268 1952
rect 12308 1912 12309 1952
rect 12267 1903 12309 1912
rect 12651 1952 12693 1961
rect 12651 1912 12652 1952
rect 12692 1912 12693 1952
rect 12651 1903 12693 1912
rect 13035 1952 13077 1961
rect 13035 1912 13036 1952
rect 13076 1912 13077 1952
rect 13035 1903 13077 1912
rect 13419 1952 13461 1961
rect 13419 1912 13420 1952
rect 13460 1912 13461 1952
rect 13419 1903 13461 1912
rect 13803 1952 13845 1961
rect 13803 1912 13804 1952
rect 13844 1912 13845 1952
rect 13803 1903 13845 1912
rect 14187 1952 14229 1961
rect 14187 1912 14188 1952
rect 14228 1912 14229 1952
rect 14187 1903 14229 1912
rect 14571 1952 14613 1961
rect 14571 1912 14572 1952
rect 14612 1912 14613 1952
rect 14571 1903 14613 1912
rect 14955 1952 14997 1961
rect 14955 1912 14956 1952
rect 14996 1912 14997 1952
rect 14955 1903 14997 1912
rect 15339 1952 15381 1961
rect 15339 1912 15340 1952
rect 15380 1912 15381 1952
rect 15339 1903 15381 1912
rect 15723 1952 15765 1961
rect 15723 1912 15724 1952
rect 15764 1912 15765 1952
rect 15723 1903 15765 1912
rect 16107 1952 16149 1961
rect 16107 1912 16108 1952
rect 16148 1912 16149 1952
rect 16107 1903 16149 1912
rect 16491 1952 16533 1961
rect 16491 1912 16492 1952
rect 16532 1912 16533 1952
rect 16491 1903 16533 1912
rect 17643 1952 17685 1961
rect 17643 1912 17644 1952
rect 17684 1912 17685 1952
rect 17643 1903 17685 1912
rect 2715 1784 2757 1793
rect 2715 1744 2716 1784
rect 2756 1744 2757 1784
rect 2715 1735 2757 1744
rect 5403 1784 5445 1793
rect 5403 1744 5404 1784
rect 5444 1744 5445 1784
rect 5403 1735 5445 1744
rect 11163 1784 11205 1793
rect 11163 1744 11164 1784
rect 11204 1744 11205 1784
rect 11163 1735 11205 1744
rect 12411 1784 12453 1793
rect 12411 1744 12412 1784
rect 12452 1744 12453 1784
rect 12411 1735 12453 1744
rect 13563 1784 13605 1793
rect 13563 1744 13564 1784
rect 13604 1744 13605 1784
rect 13563 1735 13605 1744
rect 15483 1784 15525 1793
rect 15483 1744 15484 1784
rect 15524 1744 15525 1784
rect 15483 1735 15525 1744
rect 1563 1700 1605 1709
rect 1563 1660 1564 1700
rect 1604 1660 1605 1700
rect 1563 1651 1605 1660
rect 2331 1700 2373 1709
rect 2331 1660 2332 1700
rect 2372 1660 2373 1700
rect 2331 1651 2373 1660
rect 3483 1700 3525 1709
rect 3483 1660 3484 1700
rect 3524 1660 3525 1700
rect 3483 1651 3525 1660
rect 5787 1700 5829 1709
rect 5787 1660 5788 1700
rect 5828 1660 5829 1700
rect 5787 1651 5829 1660
rect 8475 1700 8517 1709
rect 8475 1660 8476 1700
rect 8516 1660 8517 1700
rect 8475 1651 8517 1660
rect 8859 1700 8901 1709
rect 8859 1660 8860 1700
rect 8900 1660 8901 1700
rect 8859 1651 8901 1660
rect 9243 1700 9285 1709
rect 9243 1660 9244 1700
rect 9284 1660 9285 1700
rect 9243 1651 9285 1660
rect 9627 1700 9669 1709
rect 9627 1660 9628 1700
rect 9668 1660 9669 1700
rect 9627 1651 9669 1660
rect 10011 1700 10053 1709
rect 10011 1660 10012 1700
rect 10052 1660 10053 1700
rect 10011 1651 10053 1660
rect 10395 1700 10437 1709
rect 10395 1660 10396 1700
rect 10436 1660 10437 1700
rect 10395 1651 10437 1660
rect 10779 1700 10821 1709
rect 10779 1660 10780 1700
rect 10820 1660 10821 1700
rect 10779 1651 10821 1660
rect 11259 1700 11301 1709
rect 11259 1660 11260 1700
rect 11300 1660 11301 1700
rect 11259 1651 11301 1660
rect 11643 1700 11685 1709
rect 11643 1660 11644 1700
rect 11684 1660 11685 1700
rect 11643 1651 11685 1660
rect 12027 1700 12069 1709
rect 12027 1660 12028 1700
rect 12068 1660 12069 1700
rect 12027 1651 12069 1660
rect 12795 1700 12837 1709
rect 12795 1660 12796 1700
rect 12836 1660 12837 1700
rect 12795 1651 12837 1660
rect 13179 1700 13221 1709
rect 13179 1660 13180 1700
rect 13220 1660 13221 1700
rect 13179 1651 13221 1660
rect 13947 1700 13989 1709
rect 13947 1660 13948 1700
rect 13988 1660 13989 1700
rect 13947 1651 13989 1660
rect 14331 1700 14373 1709
rect 14331 1660 14332 1700
rect 14372 1660 14373 1700
rect 14331 1651 14373 1660
rect 15099 1700 15141 1709
rect 15099 1660 15100 1700
rect 15140 1660 15141 1700
rect 15099 1651 15141 1660
rect 15867 1700 15909 1709
rect 15867 1660 15868 1700
rect 15908 1660 15909 1700
rect 15867 1651 15909 1660
rect 16251 1700 16293 1709
rect 16251 1660 16252 1700
rect 16292 1660 16293 1700
rect 16251 1651 16293 1660
rect 1152 1532 20452 1556
rect 1152 1492 4928 1532
rect 4968 1492 5010 1532
rect 5050 1492 5092 1532
rect 5132 1492 5174 1532
rect 5214 1492 5256 1532
rect 5296 1492 20048 1532
rect 20088 1492 20130 1532
rect 20170 1492 20212 1532
rect 20252 1492 20294 1532
rect 20334 1492 20376 1532
rect 20416 1492 20452 1532
rect 1152 1468 20452 1492
<< via1 >>
rect 4928 95236 4968 95276
rect 5010 95236 5050 95276
rect 5092 95236 5132 95276
rect 5174 95236 5214 95276
rect 5256 95236 5296 95276
rect 20048 95236 20088 95276
rect 20130 95236 20170 95276
rect 20212 95236 20252 95276
rect 20294 95236 20334 95276
rect 20376 95236 20416 95276
rect 7324 95068 7364 95108
rect 1564 94984 1604 95024
rect 2716 94984 2756 95024
rect 3484 94984 3524 95024
rect 4636 94984 4676 95024
rect 5020 94984 5060 95024
rect 5788 94984 5828 95024
rect 6940 94984 6980 95024
rect 8092 94984 8132 95024
rect 15676 94984 15716 95024
rect 16060 94984 16100 95024
rect 16828 94984 16868 95024
rect 17212 94984 17252 95024
rect 18364 94984 18404 95024
rect 18748 94984 18788 95024
rect 19900 94984 19940 95024
rect 1324 94816 1364 94856
rect 1708 94816 1748 94856
rect 2092 94816 2132 94856
rect 2476 94816 2516 94856
rect 2860 94816 2900 94856
rect 3244 94816 3284 94856
rect 3628 94816 3668 94856
rect 4012 94816 4052 94856
rect 4396 94816 4436 94856
rect 4780 94816 4820 94856
rect 5164 94816 5204 94856
rect 5548 94816 5588 94856
rect 5932 94816 5972 94856
rect 6316 94816 6356 94856
rect 6700 94816 6740 94856
rect 7084 94816 7124 94856
rect 7468 94816 7508 94856
rect 7852 94816 7892 94856
rect 8236 94816 8276 94856
rect 8620 94816 8660 94856
rect 9196 94816 9236 94856
rect 9580 94816 9620 94856
rect 9964 94816 10004 94856
rect 10156 94816 10196 94856
rect 10732 94816 10772 94856
rect 10924 94816 10964 94856
rect 11308 94816 11348 94856
rect 11884 94816 11924 94856
rect 12076 94816 12116 94856
rect 12652 94816 12692 94856
rect 12844 94816 12884 94856
rect 13420 94816 13460 94856
rect 13612 94816 13652 94856
rect 14188 94816 14228 94856
rect 14380 94816 14420 94856
rect 14956 94816 14996 94856
rect 15916 94816 15956 94856
rect 16348 94816 16388 94856
rect 16684 94816 16724 94856
rect 17068 94816 17108 94856
rect 17452 94816 17492 94856
rect 17836 94816 17876 94856
rect 18220 94816 18260 94856
rect 18604 94816 18644 94856
rect 18988 94816 19028 94856
rect 19372 94816 19412 94856
rect 19756 94816 19796 94856
rect 20140 94816 20180 94856
rect 1948 94732 1988 94772
rect 3100 94732 3140 94772
rect 3868 94732 3908 94772
rect 5404 94732 5444 94772
rect 6172 94732 6212 94772
rect 7708 94732 7748 94772
rect 8860 94732 8900 94772
rect 10396 94732 10436 94772
rect 11548 94732 11588 94772
rect 12316 94732 12356 94772
rect 13084 94732 13124 94772
rect 13852 94732 13892 94772
rect 14620 94732 14660 94772
rect 2332 94648 2372 94688
rect 4252 94648 4292 94688
rect 6556 94648 6596 94688
rect 8476 94648 8516 94688
rect 8956 94648 8996 94688
rect 9340 94648 9380 94688
rect 9724 94648 9764 94688
rect 10492 94648 10532 94688
rect 11164 94648 11204 94688
rect 11644 94648 11684 94688
rect 12412 94648 12452 94688
rect 13180 94648 13220 94688
rect 13948 94648 13988 94688
rect 14716 94648 14756 94688
rect 16444 94648 16484 94688
rect 17596 94648 17636 94688
rect 17980 94648 18020 94688
rect 19132 94648 19172 94688
rect 19516 94648 19556 94688
rect 3688 94480 3728 94520
rect 3770 94480 3810 94520
rect 3852 94480 3892 94520
rect 3934 94480 3974 94520
rect 4016 94480 4056 94520
rect 18808 94480 18848 94520
rect 18890 94480 18930 94520
rect 18972 94480 19012 94520
rect 19054 94480 19094 94520
rect 19136 94480 19176 94520
rect 2236 94312 2276 94352
rect 2620 94312 2660 94352
rect 3004 94312 3044 94352
rect 3580 94312 3620 94352
rect 3964 94312 4004 94352
rect 4348 94312 4388 94352
rect 4732 94312 4772 94352
rect 5116 94312 5156 94352
rect 5884 94312 5924 94352
rect 6268 94312 6308 94352
rect 6652 94312 6692 94352
rect 7036 94312 7076 94352
rect 7420 94312 7460 94352
rect 7804 94312 7844 94352
rect 8572 94312 8612 94352
rect 16444 94312 16484 94352
rect 1852 94228 1892 94268
rect 3388 94228 3428 94268
rect 5500 94228 5540 94268
rect 8188 94228 8228 94268
rect 17212 94228 17252 94268
rect 1228 94144 1268 94184
rect 1612 94144 1652 94184
rect 1996 94144 2036 94184
rect 2380 94144 2420 94184
rect 2764 94144 2804 94184
rect 3148 94144 3188 94184
rect 3820 94144 3860 94184
rect 4204 94144 4244 94184
rect 4588 94144 4628 94184
rect 4972 94144 5012 94184
rect 5356 94144 5396 94184
rect 5740 94144 5780 94184
rect 6124 94144 6164 94184
rect 6508 94144 6548 94184
rect 6892 94144 6932 94184
rect 7276 94144 7316 94184
rect 7660 94144 7700 94184
rect 8044 94144 8084 94184
rect 8428 94144 8468 94184
rect 8812 94144 8852 94184
rect 9004 94144 9044 94184
rect 9580 94144 9620 94184
rect 9772 94144 9812 94184
rect 10348 94144 10388 94184
rect 10540 94144 10580 94184
rect 11116 94144 11156 94184
rect 12844 94144 12884 94184
rect 13036 94144 13076 94184
rect 13612 94144 13652 94184
rect 13804 94144 13844 94184
rect 14572 94144 14612 94184
rect 14956 94144 14996 94184
rect 15340 94144 15380 94184
rect 16204 94144 16244 94184
rect 16780 94144 16820 94184
rect 16972 94144 17012 94184
rect 17356 94144 17396 94184
rect 17596 94144 17636 94184
rect 17932 94144 17972 94184
rect 18124 94144 18164 94184
rect 18700 94144 18740 94184
rect 18844 94144 18884 94184
rect 19084 94144 19124 94184
rect 19468 94144 19508 94184
rect 19852 94144 19892 94184
rect 20236 94144 20276 94184
rect 9244 93976 9284 94016
rect 10012 93976 10052 94016
rect 10780 93976 10820 94016
rect 13276 93976 13316 94016
rect 18364 93976 18404 94016
rect 1468 93892 1508 93932
rect 9340 93892 9380 93932
rect 10108 93892 10148 93932
rect 10876 93892 10916 93932
rect 12604 93892 12644 93932
rect 13372 93892 13412 93932
rect 14044 93892 14084 93932
rect 14332 93892 14372 93932
rect 14716 93892 14756 93932
rect 15100 93892 15140 93932
rect 16540 93892 16580 93932
rect 17692 93892 17732 93932
rect 18460 93892 18500 93932
rect 19228 93892 19268 93932
rect 19612 93892 19652 93932
rect 19996 93892 20036 93932
rect 4928 93724 4968 93764
rect 5010 93724 5050 93764
rect 5092 93724 5132 93764
rect 5174 93724 5214 93764
rect 5256 93724 5296 93764
rect 20048 93724 20088 93764
rect 20130 93724 20170 93764
rect 20212 93724 20252 93764
rect 20294 93724 20334 93764
rect 20376 93724 20416 93764
rect 2716 93556 2756 93596
rect 18556 93556 18596 93596
rect 19708 93556 19748 93596
rect 2620 93472 2660 93512
rect 18460 93472 18500 93512
rect 1228 93304 1268 93344
rect 1612 93304 1652 93344
rect 1996 93304 2036 93344
rect 2380 93304 2420 93344
rect 2956 93304 2996 93344
rect 3148 93304 3188 93344
rect 17836 93304 17876 93344
rect 18220 93304 18260 93344
rect 18796 93304 18836 93344
rect 18988 93304 19028 93344
rect 19564 93304 19604 93344
rect 19948 93304 19988 93344
rect 20140 93304 20180 93344
rect 18076 93220 18116 93260
rect 19228 93220 19268 93260
rect 1468 93136 1508 93176
rect 1852 93136 1892 93176
rect 2236 93136 2276 93176
rect 3388 93136 3428 93176
rect 19324 93136 19364 93176
rect 20380 93136 20420 93176
rect 3688 92968 3728 93008
rect 3770 92968 3810 93008
rect 3852 92968 3892 93008
rect 3934 92968 3974 93008
rect 4016 92968 4056 93008
rect 18808 92968 18848 93008
rect 18890 92968 18930 93008
rect 18972 92968 19012 93008
rect 19054 92968 19094 93008
rect 19136 92968 19176 93008
rect 2716 92800 2756 92840
rect 18940 92800 18980 92840
rect 18844 92716 18884 92756
rect 1228 92632 1268 92672
rect 1612 92632 1652 92672
rect 1996 92632 2036 92672
rect 2236 92632 2276 92672
rect 2380 92632 2420 92672
rect 2956 92632 2996 92672
rect 18604 92632 18644 92672
rect 19180 92632 19220 92672
rect 19564 92632 19604 92672
rect 19756 92632 19796 92672
rect 20140 92632 20180 92672
rect 2620 92464 2660 92504
rect 19324 92464 19364 92504
rect 1468 92380 1508 92420
rect 1852 92380 1892 92420
rect 19996 92380 20036 92420
rect 20380 92380 20420 92420
rect 4928 92212 4968 92252
rect 5010 92212 5050 92252
rect 5092 92212 5132 92252
rect 5174 92212 5214 92252
rect 5256 92212 5296 92252
rect 20048 92212 20088 92252
rect 20130 92212 20170 92252
rect 20212 92212 20252 92252
rect 20294 92212 20334 92252
rect 20376 92212 20416 92252
rect 7804 92044 7844 92084
rect 19324 92044 19364 92084
rect 1228 91792 1268 91832
rect 1612 91792 1652 91832
rect 1996 91792 2036 91832
rect 2380 91792 2420 91832
rect 2764 91792 2804 91832
rect 8044 91792 8084 91832
rect 19564 91792 19604 91832
rect 19756 91792 19796 91832
rect 20140 91792 20180 91832
rect 1468 91624 1508 91664
rect 1852 91624 1892 91664
rect 2236 91624 2276 91664
rect 2620 91624 2660 91664
rect 3004 91624 3044 91664
rect 19996 91624 20036 91664
rect 20380 91624 20420 91664
rect 3688 91456 3728 91496
rect 3770 91456 3810 91496
rect 3852 91456 3892 91496
rect 3934 91456 3974 91496
rect 4016 91456 4056 91496
rect 18808 91456 18848 91496
rect 18890 91456 18930 91496
rect 18972 91456 19012 91496
rect 19054 91456 19094 91496
rect 19136 91456 19176 91496
rect 7708 91288 7748 91328
rect 8092 91204 8132 91244
rect 1228 91120 1268 91160
rect 1612 91120 1652 91160
rect 1996 91120 2036 91160
rect 2380 91120 2420 91160
rect 2764 91120 2804 91160
rect 7948 91120 7988 91160
rect 8332 91120 8372 91160
rect 19756 91120 19796 91160
rect 20140 91120 20180 91160
rect 2236 90952 2276 90992
rect 19996 90952 20036 90992
rect 1468 90868 1508 90908
rect 1852 90868 1892 90908
rect 2620 90868 2660 90908
rect 3004 90868 3044 90908
rect 20380 90868 20420 90908
rect 4928 90700 4968 90740
rect 5010 90700 5050 90740
rect 5092 90700 5132 90740
rect 5174 90700 5214 90740
rect 5256 90700 5296 90740
rect 20048 90700 20088 90740
rect 20130 90700 20170 90740
rect 20212 90700 20252 90740
rect 20294 90700 20334 90740
rect 20376 90700 20416 90740
rect 17020 90532 17060 90572
rect 11404 90364 11444 90404
rect 12652 90355 12692 90395
rect 14380 90364 14420 90404
rect 15628 90355 15668 90395
rect 1228 90280 1268 90320
rect 1468 90280 1508 90320
rect 1612 90280 1652 90320
rect 1996 90280 2036 90320
rect 2380 90280 2420 90320
rect 2764 90280 2804 90320
rect 3340 90280 3380 90320
rect 3532 90280 3572 90320
rect 3916 90280 3956 90320
rect 17260 90280 17300 90320
rect 19372 90280 19412 90320
rect 19756 90280 19796 90320
rect 20140 90280 20180 90320
rect 1852 90196 1892 90236
rect 3004 90196 3044 90236
rect 20380 90196 20420 90236
rect 2236 90112 2276 90152
rect 2620 90112 2660 90152
rect 3100 90112 3140 90152
rect 3772 90112 3812 90152
rect 4156 90112 4196 90152
rect 12844 90112 12884 90152
rect 15820 90112 15860 90152
rect 19612 90112 19652 90152
rect 19996 90112 20036 90152
rect 3688 89944 3728 89984
rect 3770 89944 3810 89984
rect 3852 89944 3892 89984
rect 3934 89944 3974 89984
rect 4016 89944 4056 89984
rect 18808 89944 18848 89984
rect 18890 89944 18930 89984
rect 18972 89944 19012 89984
rect 19054 89944 19094 89984
rect 19136 89944 19176 89984
rect 2620 89776 2660 89816
rect 3772 89776 3812 89816
rect 4156 89776 4196 89816
rect 3004 89692 3044 89732
rect 19996 89692 20036 89732
rect 1228 89608 1268 89648
rect 1612 89608 1652 89648
rect 1996 89608 2036 89648
rect 2380 89608 2420 89648
rect 2764 89608 2804 89648
rect 3148 89608 3188 89648
rect 3532 89608 3572 89648
rect 3916 89608 3956 89648
rect 4300 89608 4340 89648
rect 13612 89608 13652 89648
rect 15043 89608 15083 89648
rect 18988 89608 19028 89648
rect 19372 89608 19412 89648
rect 19756 89608 19796 89648
rect 20140 89608 20180 89648
rect 4684 89524 4724 89564
rect 5932 89524 5972 89564
rect 11404 89524 11444 89564
rect 12652 89524 12692 89564
rect 13123 89524 13163 89564
rect 13228 89524 13268 89564
rect 13708 89524 13748 89564
rect 14188 89524 14228 89564
rect 14707 89524 14747 89564
rect 15244 89524 15284 89564
rect 16492 89524 16532 89564
rect 16876 89524 16916 89564
rect 18124 89524 18164 89564
rect 2236 89440 2276 89480
rect 19228 89440 19268 89480
rect 1468 89356 1508 89396
rect 1852 89356 1892 89396
rect 3388 89356 3428 89396
rect 4540 89356 4580 89396
rect 6124 89356 6164 89396
rect 12844 89356 12884 89396
rect 14860 89356 14900 89396
rect 18316 89356 18356 89396
rect 19612 89356 19652 89396
rect 20380 89356 20420 89396
rect 4928 89188 4968 89228
rect 5010 89188 5050 89228
rect 5092 89188 5132 89228
rect 5174 89188 5214 89228
rect 5256 89188 5296 89228
rect 20048 89188 20088 89228
rect 20130 89188 20170 89228
rect 20212 89188 20252 89228
rect 20294 89188 20334 89228
rect 20376 89188 20416 89228
rect 2620 89020 2660 89060
rect 9436 89020 9476 89060
rect 14284 89020 14324 89060
rect 16300 89020 16340 89060
rect 12268 88936 12308 88976
rect 19996 88936 20036 88976
rect 2764 88852 2804 88892
rect 4012 88843 4052 88883
rect 4492 88852 4532 88892
rect 5740 88843 5780 88883
rect 7276 88843 7316 88883
rect 8524 88852 8564 88892
rect 10828 88852 10868 88892
rect 12076 88843 12116 88883
rect 12547 88852 12587 88892
rect 12652 88852 12692 88892
rect 13036 88852 13076 88892
rect 13612 88843 13652 88883
rect 14092 88843 14132 88883
rect 14563 88852 14603 88892
rect 14668 88852 14708 88892
rect 15052 88852 15092 88892
rect 15628 88843 15668 88883
rect 16108 88843 16148 88883
rect 16876 88852 16916 88892
rect 18124 88843 18164 88883
rect 1228 88768 1268 88808
rect 1612 88768 1652 88808
rect 1996 88768 2036 88808
rect 2380 88768 2420 88808
rect 6124 88768 6164 88808
rect 9196 88768 9236 88808
rect 9532 88768 9572 88808
rect 9772 88768 9812 88808
rect 10156 88768 10196 88808
rect 10636 88768 10676 88808
rect 13132 88768 13172 88808
rect 15148 88768 15188 88808
rect 18604 88768 18644 88808
rect 18988 88768 19028 88808
rect 19372 88768 19412 88808
rect 19756 88768 19796 88808
rect 20140 88768 20180 88808
rect 20380 88768 20420 88808
rect 2236 88684 2276 88724
rect 18844 88684 18884 88724
rect 1468 88600 1508 88640
rect 1852 88600 1892 88640
rect 4204 88600 4244 88640
rect 5932 88600 5972 88640
rect 6364 88600 6404 88640
rect 7084 88600 7124 88640
rect 9916 88600 9956 88640
rect 10396 88600 10436 88640
rect 18316 88600 18356 88640
rect 19228 88600 19268 88640
rect 19612 88600 19652 88640
rect 3688 88432 3728 88472
rect 3770 88432 3810 88472
rect 3852 88432 3892 88472
rect 3934 88432 3974 88472
rect 4016 88432 4056 88472
rect 18808 88432 18848 88472
rect 18890 88432 18930 88472
rect 18972 88432 19012 88472
rect 19054 88432 19094 88472
rect 19136 88432 19176 88472
rect 8668 88264 8708 88304
rect 12172 88264 12212 88304
rect 12796 88264 12836 88304
rect 9100 88180 9140 88220
rect 1228 88096 1268 88136
rect 1900 88096 1940 88136
rect 2284 88096 2324 88136
rect 4396 88096 4436 88136
rect 5356 88096 5396 88136
rect 8908 88096 8948 88136
rect 12556 88096 12596 88136
rect 13516 88096 13556 88136
rect 18220 88096 18260 88136
rect 2764 88012 2804 88052
rect 4012 88012 4052 88052
rect 4867 88012 4907 88052
rect 4972 88012 5012 88052
rect 5452 88012 5492 88052
rect 5932 88012 5972 88052
rect 6420 88012 6460 88052
rect 6988 88012 7028 88052
rect 8236 88012 8276 88052
rect 9292 88012 9332 88052
rect 10540 88012 10580 88052
rect 10732 88012 10772 88052
rect 11988 88012 12028 88052
rect 13027 88012 13067 88052
rect 13132 88012 13172 88052
rect 13612 88012 13652 88052
rect 14092 88012 14132 88052
rect 14611 88012 14651 88052
rect 15148 88012 15188 88052
rect 16396 88012 16436 88052
rect 16588 88012 16628 88052
rect 17836 88012 17876 88052
rect 18604 88012 18644 88052
rect 19852 88012 19892 88052
rect 2140 87928 2180 87968
rect 4204 87928 4244 87968
rect 14956 87928 14996 87968
rect 18028 87928 18068 87968
rect 1468 87844 1508 87884
rect 2524 87844 2564 87884
rect 4636 87844 4676 87884
rect 6604 87844 6644 87884
rect 6796 87844 6836 87884
rect 14764 87844 14804 87884
rect 18460 87844 18500 87884
rect 20044 87844 20084 87884
rect 4928 87676 4968 87716
rect 5010 87676 5050 87716
rect 5092 87676 5132 87716
rect 5174 87676 5214 87716
rect 5256 87676 5296 87716
rect 20048 87676 20088 87716
rect 20130 87676 20170 87716
rect 20212 87676 20252 87716
rect 20294 87676 20334 87716
rect 20376 87676 20416 87716
rect 6604 87508 6644 87548
rect 8716 87508 8756 87548
rect 13516 87508 13556 87548
rect 3868 87424 3908 87464
rect 8908 87424 8948 87464
rect 17443 87424 17483 87464
rect 1612 87340 1652 87380
rect 2860 87331 2900 87371
rect 4846 87340 4886 87380
rect 4972 87340 5012 87380
rect 5356 87340 5396 87380
rect 5932 87331 5972 87371
rect 6412 87331 6452 87371
rect 6979 87340 7019 87380
rect 7084 87340 7124 87380
rect 7468 87340 7508 87380
rect 8044 87331 8084 87371
rect 8524 87331 8564 87371
rect 9100 87331 9140 87371
rect 10348 87340 10388 87380
rect 11116 87340 11156 87380
rect 12364 87331 12404 87371
rect 12748 87340 12788 87380
rect 12863 87340 12903 87380
rect 13036 87340 13076 87380
rect 13267 87340 13307 87380
rect 13369 87308 13409 87348
rect 15724 87340 15764 87380
rect 16972 87331 17012 87371
rect 17635 87340 17675 87380
rect 18124 87331 18164 87371
rect 18604 87340 18644 87380
rect 19084 87340 19124 87380
rect 19202 87340 19242 87380
rect 1228 87256 1268 87296
rect 3436 87256 3476 87296
rect 3628 87256 3668 87296
rect 4012 87256 4052 87296
rect 4588 87256 4628 87296
rect 5452 87256 5492 87296
rect 7564 87256 7604 87296
rect 10732 87256 10772 87296
rect 18700 87256 18740 87296
rect 19756 87256 19796 87296
rect 20140 87256 20180 87296
rect 20380 87256 20420 87296
rect 4252 87172 4292 87212
rect 12556 87172 12596 87212
rect 1468 87088 1508 87128
rect 3052 87088 3092 87128
rect 3196 87088 3236 87128
rect 4348 87088 4388 87128
rect 10972 87088 11012 87128
rect 12748 87088 12788 87128
rect 17164 87088 17204 87128
rect 19996 87088 20036 87128
rect 3688 86920 3728 86960
rect 3770 86920 3810 86960
rect 3852 86920 3892 86960
rect 3934 86920 3974 86960
rect 4016 86920 4056 86960
rect 18808 86920 18848 86960
rect 18890 86920 18930 86960
rect 18972 86920 19012 86960
rect 19054 86920 19094 86960
rect 19136 86920 19176 86960
rect 2764 86752 2804 86792
rect 6844 86752 6884 86792
rect 9235 86752 9275 86792
rect 9628 86752 9668 86792
rect 10300 86752 10340 86792
rect 10684 86752 10724 86792
rect 12268 86752 12308 86792
rect 5164 86584 5204 86624
rect 6604 86584 6644 86624
rect 6988 86584 7028 86624
rect 7948 86584 7988 86624
rect 9388 86584 9428 86624
rect 10060 86584 10100 86624
rect 10444 86584 10484 86624
rect 12460 86584 12500 86624
rect 18028 86584 18068 86624
rect 19756 86584 19796 86624
rect 20140 86584 20180 86624
rect 1324 86500 1364 86540
rect 2572 86500 2612 86540
rect 2956 86500 2996 86540
rect 4204 86500 4244 86540
rect 4675 86500 4715 86540
rect 4780 86500 4820 86540
rect 5260 86500 5300 86540
rect 5740 86500 5780 86540
rect 6228 86500 6268 86540
rect 7438 86500 7478 86540
rect 7564 86500 7604 86540
rect 8044 86500 8084 86540
rect 8523 86500 8563 86540
rect 9012 86500 9052 86540
rect 10828 86500 10868 86540
rect 12076 86500 12116 86540
rect 12835 86500 12875 86540
rect 12953 86500 12993 86540
rect 13085 86500 13125 86540
rect 13219 86500 13259 86540
rect 13363 86500 13403 86540
rect 13900 86500 13940 86540
rect 15148 86500 15188 86540
rect 15532 86500 15572 86540
rect 16780 86500 16820 86540
rect 17539 86500 17579 86540
rect 17644 86500 17684 86540
rect 18124 86500 18164 86540
rect 18604 86500 18644 86540
rect 19092 86500 19132 86540
rect 4396 86416 4436 86456
rect 12268 86416 12308 86456
rect 15340 86416 15380 86456
rect 16972 86416 17012 86456
rect 20380 86416 20420 86456
rect 6412 86332 6452 86372
rect 7228 86332 7268 86372
rect 12700 86332 12740 86372
rect 13036 86332 13076 86372
rect 19276 86332 19316 86372
rect 19996 86332 20036 86372
rect 4928 86164 4968 86204
rect 5010 86164 5050 86204
rect 5092 86164 5132 86204
rect 5174 86164 5214 86204
rect 5256 86164 5296 86204
rect 20048 86164 20088 86204
rect 20130 86164 20170 86204
rect 20212 86164 20252 86204
rect 20294 86164 20334 86204
rect 20376 86164 20416 86204
rect 3964 85996 4004 86036
rect 5836 85996 5876 86036
rect 6748 85996 6788 86036
rect 8620 85996 8660 86036
rect 12508 85996 12548 86036
rect 3580 85912 3620 85952
rect 18172 85912 18212 85952
rect 1708 85828 1748 85868
rect 2956 85819 2996 85859
rect 4396 85828 4436 85868
rect 5644 85819 5684 85859
rect 7180 85828 7220 85868
rect 8428 85819 8468 85859
rect 8812 85828 8852 85868
rect 10060 85819 10100 85859
rect 10444 85828 10484 85868
rect 11692 85819 11732 85859
rect 12364 85828 12404 85868
rect 12652 85828 12692 85868
rect 12835 85828 12875 85868
rect 13132 85828 13172 85868
rect 13369 85828 13409 85868
rect 13516 85828 13556 85868
rect 13804 85828 13844 85868
rect 15052 85819 15092 85859
rect 15436 85828 15476 85868
rect 16684 85819 16724 85859
rect 18604 85828 18644 85868
rect 19852 85819 19892 85859
rect 1228 85744 1268 85784
rect 3340 85744 3380 85784
rect 3724 85744 3764 85784
rect 6076 85744 6116 85784
rect 6316 85744 6356 85784
rect 6508 85744 6548 85784
rect 13036 85744 13076 85784
rect 13267 85735 13307 85775
rect 17260 85744 17300 85784
rect 17452 85744 17492 85784
rect 17836 85744 17876 85784
rect 18412 85744 18452 85784
rect 17020 85660 17060 85700
rect 18076 85660 18116 85700
rect 1468 85576 1508 85616
rect 3148 85576 3188 85616
rect 10252 85576 10292 85616
rect 11884 85576 11924 85616
rect 12835 85576 12875 85616
rect 13660 85576 13700 85616
rect 15244 85576 15284 85616
rect 16876 85576 16916 85616
rect 17692 85576 17732 85616
rect 20044 85576 20084 85616
rect 3688 85408 3728 85448
rect 3770 85408 3810 85448
rect 3852 85408 3892 85448
rect 3934 85408 3974 85448
rect 4016 85408 4056 85448
rect 18808 85408 18848 85448
rect 18890 85408 18930 85448
rect 18972 85408 19012 85448
rect 19054 85408 19094 85448
rect 19136 85408 19176 85448
rect 8188 85240 8228 85280
rect 8860 85240 8900 85280
rect 4876 85156 4916 85196
rect 14284 85156 14324 85196
rect 3052 85072 3092 85112
rect 7468 85072 7508 85112
rect 7708 85072 7748 85112
rect 8428 85072 8468 85112
rect 8620 85072 8660 85112
rect 12844 85072 12884 85112
rect 15628 85072 15668 85112
rect 1420 84988 1460 85028
rect 2668 84988 2708 85028
rect 3436 84988 3476 85028
rect 4684 84988 4724 85028
rect 5260 84988 5300 85028
rect 6508 84988 6548 85028
rect 6883 84988 6923 85028
rect 7852 84988 7892 85028
rect 8044 84988 8084 85028
rect 9004 84988 9044 85028
rect 10252 84988 10292 85028
rect 10636 84988 10676 85028
rect 11884 84988 11924 85028
rect 12355 84988 12395 85028
rect 12460 84988 12500 85028
rect 12940 84988 12980 85028
rect 13420 84988 13460 85028
rect 13908 84988 13948 85028
rect 14284 84988 14324 85028
rect 14572 84988 14612 85028
rect 15139 84988 15179 85028
rect 15244 84988 15284 85028
rect 15724 84988 15764 85028
rect 16204 84988 16244 85028
rect 16723 84988 16763 85028
rect 17068 84988 17108 85028
rect 18316 84988 18356 85028
rect 18700 84988 18740 85028
rect 19948 84988 19988 85028
rect 3292 84904 3332 84944
rect 7084 84904 7124 84944
rect 7194 84904 7234 84944
rect 7948 84904 7988 84944
rect 2860 84820 2900 84860
rect 6700 84820 6740 84860
rect 6979 84820 7019 84860
rect 10444 84820 10484 84860
rect 12076 84820 12116 84860
rect 14092 84820 14132 84860
rect 16876 84820 16916 84860
rect 18508 84820 18548 84860
rect 20140 84820 20180 84860
rect 4928 84652 4968 84692
rect 5010 84652 5050 84692
rect 5092 84652 5132 84692
rect 5174 84652 5214 84692
rect 5256 84652 5296 84692
rect 20048 84652 20088 84692
rect 20130 84652 20170 84692
rect 20212 84652 20252 84692
rect 20294 84652 20334 84692
rect 20376 84652 20416 84692
rect 4492 84484 4532 84524
rect 7660 84484 7700 84524
rect 8428 84484 8468 84524
rect 9148 84484 9188 84524
rect 12364 84484 12404 84524
rect 12748 84484 12788 84524
rect 14380 84484 14420 84524
rect 14764 84484 14804 84524
rect 16876 84484 16916 84524
rect 19564 84484 19604 84524
rect 5692 84400 5732 84440
rect 13708 84400 13748 84440
rect 14174 84400 14214 84440
rect 14275 84400 14315 84440
rect 2755 84316 2795 84356
rect 2860 84316 2900 84356
rect 3244 84316 3284 84356
rect 3820 84307 3860 84347
rect 4300 84307 4340 84347
rect 5923 84316 5963 84356
rect 6028 84316 6068 84356
rect 6412 84316 6452 84356
rect 6988 84307 7028 84347
rect 7468 84307 7508 84347
rect 7948 84316 7988 84356
rect 8179 84316 8219 84356
rect 8333 84316 8373 84356
rect 8524 84316 8564 84356
rect 9292 84316 9332 84356
rect 10540 84307 10580 84347
rect 10924 84316 10964 84356
rect 12172 84307 12212 84347
rect 12844 84316 12884 84356
rect 13081 84316 13121 84356
rect 13324 84316 13364 84356
rect 13603 84316 13643 84356
rect 14482 84291 14522 84331
rect 14668 84316 14708 84356
rect 14860 84316 14900 84356
rect 15139 84316 15179 84356
rect 15244 84316 15284 84356
rect 15628 84316 15668 84356
rect 16204 84307 16244 84347
rect 16684 84307 16724 84347
rect 17827 84316 17867 84356
rect 17932 84316 17972 84356
rect 18316 84316 18356 84356
rect 18892 84307 18932 84347
rect 19372 84307 19412 84347
rect 1228 84232 1268 84272
rect 1612 84232 1652 84272
rect 1996 84232 2036 84272
rect 3340 84232 3380 84272
rect 4684 84232 4724 84272
rect 5068 84232 5108 84272
rect 5452 84232 5492 84272
rect 6508 84232 6548 84272
rect 7852 84232 7892 84272
rect 8067 84232 8107 84272
rect 8908 84232 8948 84272
rect 12979 84223 13019 84263
rect 15724 84232 15764 84272
rect 17068 84232 17108 84272
rect 18412 84232 18452 84272
rect 19756 84232 19796 84272
rect 20140 84232 20180 84272
rect 5308 84148 5348 84188
rect 13996 84148 14036 84188
rect 1468 84064 1508 84104
rect 1852 84064 1892 84104
rect 2236 84064 2276 84104
rect 4924 84064 4964 84104
rect 9148 84064 9188 84104
rect 10732 84064 10772 84104
rect 17308 84064 17348 84104
rect 19996 84064 20036 84104
rect 20380 84064 20420 84104
rect 3688 83896 3728 83936
rect 3770 83896 3810 83936
rect 3852 83896 3892 83936
rect 3934 83896 3974 83936
rect 4016 83896 4056 83936
rect 18808 83896 18848 83936
rect 18890 83896 18930 83936
rect 18972 83896 19012 83936
rect 19054 83896 19094 83936
rect 19136 83896 19176 83936
rect 5308 83728 5348 83768
rect 5884 83728 5924 83768
rect 7660 83728 7700 83768
rect 9340 83728 9380 83768
rect 13075 83728 13115 83768
rect 14812 83728 14852 83768
rect 19603 83728 19643 83768
rect 7468 83644 7508 83684
rect 11020 83644 11060 83684
rect 19756 83644 19796 83684
rect 3916 83560 3956 83600
rect 5548 83560 5588 83600
rect 8908 83560 8948 83600
rect 9100 83560 9140 83600
rect 11788 83560 11828 83600
rect 13612 83560 13652 83600
rect 13852 83560 13892 83600
rect 14188 83560 14228 83600
rect 14524 83560 14564 83600
rect 15676 83560 15716 83600
rect 15916 83560 15956 83600
rect 18316 83560 18356 83600
rect 20140 83560 20180 83600
rect 20380 83560 20420 83600
rect 1516 83476 1556 83516
rect 2764 83476 2804 83516
rect 3427 83476 3467 83516
rect 3532 83476 3572 83516
rect 4012 83476 4052 83516
rect 4492 83476 4532 83516
rect 4980 83476 5020 83516
rect 5740 83476 5780 83516
rect 6028 83476 6068 83516
rect 7276 83476 7316 83516
rect 8044 83467 8084 83507
rect 8332 83476 8372 83516
rect 8567 83476 8607 83516
rect 8707 83476 8747 83516
rect 8812 83476 8852 83516
rect 9580 83476 9620 83516
rect 10828 83476 10868 83516
rect 11278 83476 11318 83516
rect 11404 83476 11444 83516
rect 11884 83476 11924 83516
rect 12364 83476 12404 83516
rect 12852 83476 12892 83516
rect 14947 83476 14987 83516
rect 15258 83476 15298 83516
rect 16108 83476 16148 83516
rect 17356 83476 17396 83516
rect 17827 83476 17867 83516
rect 17932 83476 17972 83516
rect 18412 83476 18452 83516
rect 18892 83476 18932 83516
rect 19411 83476 19451 83516
rect 19756 83476 19796 83516
rect 19948 83476 19988 83516
rect 7948 83392 7988 83432
rect 13948 83392 13988 83432
rect 15052 83392 15092 83432
rect 17548 83392 17588 83432
rect 2956 83308 2996 83348
rect 5164 83308 5204 83348
rect 15148 83308 15188 83348
rect 4928 83140 4968 83180
rect 5010 83140 5050 83180
rect 5092 83140 5132 83180
rect 5174 83140 5214 83180
rect 5256 83140 5296 83180
rect 20048 83140 20088 83180
rect 20130 83140 20170 83180
rect 20212 83140 20252 83180
rect 20294 83140 20334 83180
rect 20376 83140 20416 83180
rect 4972 82972 5012 83012
rect 8428 82972 8468 83012
rect 13132 82972 13172 83012
rect 14476 82972 14516 83012
rect 14908 82972 14948 83012
rect 5164 82888 5204 82928
rect 16012 82888 16052 82928
rect 1516 82804 1556 82844
rect 2764 82795 2804 82835
rect 3235 82804 3275 82844
rect 3340 82804 3380 82844
rect 3724 82804 3764 82844
rect 4300 82795 4340 82835
rect 4780 82795 4820 82835
rect 5356 82795 5396 82835
rect 6604 82804 6644 82844
rect 6988 82804 7028 82844
rect 8236 82795 8276 82835
rect 8620 82804 8660 82844
rect 9868 82795 9908 82835
rect 11395 82804 11435 82844
rect 11500 82804 11540 82844
rect 11884 82804 11924 82844
rect 12460 82795 12500 82835
rect 12940 82795 12980 82835
rect 14572 82804 14612 82844
rect 14809 82804 14849 82844
rect 15244 82804 15284 82844
rect 15353 82804 15393 82844
rect 15628 82804 15668 82844
rect 15916 82804 15956 82844
rect 16108 82804 16148 82844
rect 16300 82804 16340 82844
rect 16492 82804 16532 82844
rect 16876 82804 16916 82844
rect 18124 82795 18164 82835
rect 18700 82795 18740 82835
rect 19948 82804 19988 82844
rect 3859 82720 3899 82760
rect 11980 82720 12020 82760
rect 13420 82720 13460 82760
rect 14092 82720 14132 82760
rect 14691 82720 14731 82760
rect 20140 82720 20180 82760
rect 13660 82636 13700 82676
rect 16300 82636 16340 82676
rect 20380 82636 20420 82676
rect 2956 82552 2996 82592
rect 10060 82552 10100 82592
rect 14332 82552 14372 82592
rect 18316 82552 18356 82592
rect 18508 82552 18548 82592
rect 3688 82384 3728 82424
rect 3770 82384 3810 82424
rect 3852 82384 3892 82424
rect 3934 82384 3974 82424
rect 4016 82384 4056 82424
rect 18808 82384 18848 82424
rect 18890 82384 18930 82424
rect 18972 82384 19012 82424
rect 19054 82384 19094 82424
rect 19136 82384 19176 82424
rect 7276 82216 7316 82256
rect 13660 82216 13700 82256
rect 6604 82132 6644 82172
rect 3724 82048 3764 82088
rect 8428 82048 8468 82088
rect 8620 82048 8660 82088
rect 11692 82048 11732 82088
rect 13420 82048 13460 82088
rect 14380 82048 14420 82088
rect 16252 82048 16292 82088
rect 18892 82048 18932 82088
rect 1516 81964 1556 82004
rect 2764 81964 2804 82004
rect 3235 81964 3275 82004
rect 3340 81964 3380 82004
rect 3820 81964 3860 82004
rect 4300 81964 4340 82004
rect 4788 81964 4828 82004
rect 5164 81964 5204 82004
rect 6412 81964 6452 82004
rect 6743 81964 6783 82004
rect 6883 81964 6923 82004
rect 6988 81964 7028 82004
rect 7276 81964 7316 82004
rect 7564 81964 7604 82004
rect 7756 81964 7796 82004
rect 7939 81964 7979 82004
rect 9100 81964 9140 82004
rect 9292 81964 9332 82004
rect 10540 81964 10580 82004
rect 11203 81964 11243 82004
rect 11308 81964 11348 82004
rect 11788 81964 11828 82004
rect 12268 81964 12308 82004
rect 12756 81964 12796 82004
rect 13891 81964 13931 82004
rect 13996 81964 14036 82004
rect 14476 81964 14516 82004
rect 14956 81964 14996 82004
rect 15444 81964 15484 82004
rect 15811 81964 15851 82004
rect 16108 81964 16148 82004
rect 16396 81964 16436 82004
rect 16588 81964 16628 82004
rect 17836 81964 17876 82004
rect 18382 81964 18422 82004
rect 18513 81964 18553 82004
rect 18988 81964 19028 82004
rect 19468 81964 19508 82004
rect 19956 81964 19996 82004
rect 7852 81880 7892 81920
rect 8860 81880 8900 81920
rect 10732 81880 10772 81920
rect 16012 81880 16052 81920
rect 2956 81796 2996 81836
rect 4972 81796 5012 81836
rect 7075 81796 7115 81836
rect 8188 81796 8228 81836
rect 8956 81796 8996 81836
rect 12940 81796 12980 81836
rect 13660 81796 13700 81836
rect 15628 81796 15668 81836
rect 18028 81796 18068 81836
rect 20140 81796 20180 81836
rect 4928 81628 4968 81668
rect 5010 81628 5050 81668
rect 5092 81628 5132 81668
rect 5174 81628 5214 81668
rect 5256 81628 5296 81668
rect 20048 81628 20088 81668
rect 20130 81628 20170 81668
rect 20212 81628 20252 81668
rect 20294 81628 20334 81668
rect 20376 81628 20416 81668
rect 4636 81460 4676 81500
rect 6604 81460 6644 81500
rect 7843 81460 7883 81500
rect 8860 81460 8900 81500
rect 10972 81460 11012 81500
rect 13036 81460 13076 81500
rect 17059 81460 17099 81500
rect 17500 81460 17540 81500
rect 20140 81460 20180 81500
rect 7276 81376 7316 81416
rect 7948 81376 7988 81416
rect 10540 81376 10580 81416
rect 14956 81376 14996 81416
rect 1612 81292 1652 81332
rect 2860 81283 2900 81323
rect 4867 81292 4907 81332
rect 4972 81292 5012 81332
rect 5356 81292 5396 81332
rect 5932 81283 5972 81323
rect 6412 81283 6452 81323
rect 6892 81292 6932 81332
rect 7171 81292 7211 81332
rect 7747 81292 7787 81332
rect 8055 81292 8095 81332
rect 8236 81292 8276 81332
rect 8419 81292 8459 81332
rect 9100 81292 9140 81332
rect 10348 81283 10388 81323
rect 11299 81292 11339 81332
rect 11404 81292 11444 81332
rect 11788 81292 11828 81332
rect 12364 81283 12404 81323
rect 12844 81283 12884 81323
rect 13516 81292 13556 81332
rect 14764 81283 14804 81323
rect 15340 81283 15380 81323
rect 16588 81292 16628 81332
rect 1228 81208 1268 81248
rect 3244 81208 3284 81248
rect 3628 81208 3668 81248
rect 3964 81208 4004 81248
rect 4204 81208 4244 81248
rect 4396 81208 4436 81248
rect 5452 81208 5492 81248
rect 8620 81208 8660 81248
rect 10732 81208 10772 81248
rect 11884 81208 11924 81248
rect 16732 81250 16772 81290
rect 16972 81292 17012 81332
rect 18403 81292 18443 81332
rect 18508 81292 18548 81332
rect 18892 81292 18932 81332
rect 19468 81283 19508 81323
rect 19948 81283 19988 81323
rect 16867 81208 16907 81248
rect 17740 81208 17780 81248
rect 17932 81208 17972 81248
rect 18988 81208 19028 81248
rect 3868 81124 3908 81164
rect 7564 81124 7604 81164
rect 8419 81124 8459 81164
rect 1468 81040 1508 81080
rect 3052 81040 3092 81080
rect 3484 81040 3524 81080
rect 15148 81040 15188 81080
rect 18172 81040 18212 81080
rect 3688 80872 3728 80912
rect 3770 80872 3810 80912
rect 3852 80872 3892 80912
rect 3934 80872 3974 80912
rect 4016 80872 4056 80912
rect 18808 80872 18848 80912
rect 18890 80872 18930 80912
rect 18972 80872 19012 80912
rect 19054 80872 19094 80912
rect 19136 80872 19176 80912
rect 5932 80704 5972 80744
rect 4348 80620 4388 80660
rect 1228 80536 1268 80576
rect 3340 80536 3380 80576
rect 3724 80536 3764 80576
rect 4108 80536 4148 80576
rect 6691 80536 6731 80576
rect 10348 80536 10388 80576
rect 12460 80536 12500 80576
rect 12844 80536 12884 80576
rect 17164 80536 17204 80576
rect 1708 80452 1748 80492
rect 2956 80452 2996 80492
rect 4492 80452 4532 80492
rect 5740 80452 5780 80492
rect 6115 80452 6155 80492
rect 6412 80452 6452 80492
rect 6551 80452 6591 80492
rect 6796 80452 6836 80492
rect 7084 80452 7124 80492
rect 8332 80452 8372 80492
rect 8908 80452 8948 80492
rect 10156 80452 10196 80492
rect 10732 80452 10772 80492
rect 11980 80452 12020 80492
rect 13228 80452 13268 80492
rect 14476 80452 14516 80492
rect 14956 80452 14996 80492
rect 16204 80452 16244 80492
rect 16675 80452 16715 80492
rect 16780 80452 16820 80492
rect 17260 80452 17300 80492
rect 17740 80452 17780 80492
rect 18228 80452 18268 80492
rect 18604 80452 18644 80492
rect 19852 80452 19892 80492
rect 3580 80368 3620 80408
rect 6316 80368 6356 80408
rect 6883 80368 6923 80408
rect 12172 80368 12212 80408
rect 14668 80368 14708 80408
rect 16396 80368 16436 80408
rect 1468 80284 1508 80324
rect 3148 80284 3188 80324
rect 3964 80284 4004 80324
rect 8524 80284 8564 80324
rect 8716 80284 8756 80324
rect 10588 80284 10628 80324
rect 12700 80284 12740 80324
rect 13084 80284 13124 80324
rect 18412 80284 18452 80324
rect 20044 80284 20084 80324
rect 4928 80116 4968 80156
rect 5010 80116 5050 80156
rect 5092 80116 5132 80156
rect 5174 80116 5214 80156
rect 5256 80116 5296 80156
rect 20048 80116 20088 80156
rect 20130 80116 20170 80156
rect 20212 80116 20252 80156
rect 20294 80116 20334 80156
rect 20376 80116 20416 80156
rect 3619 79948 3659 79988
rect 7468 79948 7508 79988
rect 9484 79948 9524 79988
rect 10300 79948 10340 79988
rect 17020 79948 17060 79988
rect 3427 79855 3467 79895
rect 5836 79864 5876 79904
rect 9916 79864 9956 79904
rect 12508 79864 12548 79904
rect 1516 79780 1556 79820
rect 2764 79771 2804 79811
rect 3139 79780 3179 79820
rect 3244 79771 3284 79811
rect 3523 79780 3563 79820
rect 3657 79780 3697 79820
rect 4396 79780 4436 79820
rect 5644 79771 5684 79811
rect 6028 79780 6068 79820
rect 7276 79771 7316 79811
rect 7747 79780 7787 79820
rect 7852 79780 7892 79820
rect 8236 79780 8276 79820
rect 8812 79771 8852 79811
rect 9292 79771 9332 79811
rect 12172 79780 12212 79820
rect 12300 79756 12340 79796
rect 12638 79780 12678 79820
rect 12748 79780 12788 79820
rect 12940 79780 12980 79820
rect 13132 79780 13172 79820
rect 14380 79771 14420 79811
rect 14764 79780 14804 79820
rect 16012 79771 16052 79811
rect 17452 79780 17492 79820
rect 18700 79771 18740 79811
rect 3916 79696 3956 79736
rect 8332 79696 8372 79736
rect 9676 79696 9716 79736
rect 10060 79696 10100 79736
rect 10636 79696 10676 79736
rect 11116 79696 11156 79736
rect 11788 79696 11828 79736
rect 16684 79696 16724 79736
rect 17260 79696 17300 79736
rect 19372 79696 19412 79736
rect 19756 79696 19796 79736
rect 20140 79696 20180 79736
rect 12748 79612 12788 79652
rect 19612 79612 19652 79652
rect 20380 79612 20420 79652
rect 2956 79528 2996 79568
rect 4156 79528 4196 79568
rect 10396 79528 10436 79568
rect 11356 79528 11396 79568
rect 12028 79528 12068 79568
rect 14572 79528 14612 79568
rect 16204 79528 16244 79568
rect 16924 79528 16964 79568
rect 18892 79528 18932 79568
rect 19996 79528 20036 79568
rect 3688 79360 3728 79400
rect 3770 79360 3810 79400
rect 3852 79360 3892 79400
rect 3934 79360 3974 79400
rect 4016 79360 4056 79400
rect 18808 79360 18848 79400
rect 18890 79360 18930 79400
rect 18972 79360 19012 79400
rect 19054 79360 19094 79400
rect 19136 79360 19176 79400
rect 3244 79192 3284 79232
rect 5500 79108 5540 79148
rect 17932 79108 17972 79148
rect 1228 79024 1268 79064
rect 8140 79024 8180 79064
rect 9772 79024 9812 79064
rect 9964 79024 10004 79064
rect 10732 79024 10772 79064
rect 14284 79024 14324 79064
rect 15571 79024 15611 79064
rect 15916 79024 15956 79064
rect 16108 79024 16148 79064
rect 1612 78940 1652 78980
rect 2860 78940 2900 78980
rect 3244 78940 3284 78980
rect 3359 78940 3399 78980
rect 3532 78940 3572 78980
rect 3916 78940 3956 78980
rect 5164 78940 5204 78980
rect 5644 78940 5684 78980
rect 5836 78940 5876 78980
rect 7084 78940 7124 78980
rect 7651 78940 7691 78980
rect 7756 78940 7796 78980
rect 8236 78940 8276 78980
rect 8719 78940 8759 78980
rect 9204 78940 9244 78980
rect 11116 78940 11156 78980
rect 12364 78940 12404 78980
rect 12739 78940 12779 78980
rect 12844 78951 12884 78991
rect 12989 78940 13029 78980
rect 13123 78940 13163 78980
rect 13257 78940 13297 78980
rect 13795 78940 13835 78980
rect 13900 78940 13940 78980
rect 14380 78940 14420 78980
rect 14860 78940 14900 78980
rect 15348 78940 15388 78980
rect 16492 78940 16532 78980
rect 17740 78940 17780 78980
rect 18124 78940 18164 78980
rect 19372 78940 19412 78980
rect 19703 78940 19743 78980
rect 19843 78940 19883 78980
rect 19948 78940 19988 78980
rect 7276 78856 7316 78896
rect 9532 78856 9572 78896
rect 12556 78856 12596 78896
rect 1468 78772 1508 78812
rect 3052 78772 3092 78812
rect 5356 78772 5396 78812
rect 9388 78772 9428 78812
rect 10204 78772 10244 78812
rect 10492 78772 10532 78812
rect 13219 78772 13259 78812
rect 15676 78772 15716 78812
rect 16348 78772 16388 78812
rect 19564 78772 19604 78812
rect 20035 78772 20075 78812
rect 4928 78604 4968 78644
rect 5010 78604 5050 78644
rect 5092 78604 5132 78644
rect 5174 78604 5214 78644
rect 5256 78604 5296 78644
rect 20048 78604 20088 78644
rect 20130 78604 20170 78644
rect 20212 78604 20252 78644
rect 20294 78604 20334 78644
rect 20376 78604 20416 78644
rect 3043 78436 3083 78476
rect 5356 78436 5396 78476
rect 8716 78436 8756 78476
rect 11980 78436 12020 78476
rect 12316 78436 12356 78476
rect 13900 78436 13940 78476
rect 14860 78436 14900 78476
rect 16972 78436 17012 78476
rect 20323 78436 20363 78476
rect 17539 78352 17579 78392
rect 1228 78268 1268 78308
rect 2476 78259 2516 78299
rect 3204 78254 3244 78294
rect 3340 78268 3380 78308
rect 3598 78268 3638 78308
rect 3724 78268 3764 78308
rect 4108 78268 4148 78308
rect 4684 78259 4724 78299
rect 5164 78259 5204 78299
rect 5740 78259 5780 78299
rect 6988 78268 7028 78308
rect 7276 78268 7316 78308
rect 8524 78247 8564 78287
rect 8908 78268 8948 78308
rect 10156 78259 10196 78299
rect 10540 78268 10580 78308
rect 11788 78259 11828 78299
rect 12172 78268 12212 78308
rect 12460 78268 12500 78308
rect 13708 78259 13748 78299
rect 14764 78268 14804 78308
rect 14947 78268 14987 78308
rect 15235 78268 15275 78308
rect 15340 78268 15380 78308
rect 15724 78268 15764 78308
rect 16300 78259 16340 78299
rect 16780 78259 16820 78299
rect 17731 78268 17771 78308
rect 18220 78248 18260 78288
rect 18700 78268 18740 78308
rect 19180 78268 19220 78308
rect 19298 78268 19338 78308
rect 19564 78268 19604 78308
rect 19852 78268 19892 78308
rect 19991 78268 20031 78308
rect 20236 78268 20276 78308
rect 4204 78184 4244 78224
rect 14092 78184 14132 78224
rect 15820 78184 15860 78224
rect 17164 78184 17204 78224
rect 18796 78184 18836 78224
rect 20131 78184 20171 78224
rect 5548 78100 5588 78140
rect 10348 78100 10388 78140
rect 19564 78100 19604 78140
rect 2668 78016 2708 78056
rect 14332 78016 14372 78056
rect 17404 78016 17444 78056
rect 3688 77848 3728 77888
rect 3770 77848 3810 77888
rect 3852 77848 3892 77888
rect 3934 77848 3974 77888
rect 4016 77848 4056 77888
rect 18808 77848 18848 77888
rect 18890 77848 18930 77888
rect 18972 77848 19012 77888
rect 19054 77848 19094 77888
rect 19136 77848 19176 77888
rect 10540 77680 10580 77720
rect 15292 77680 15332 77720
rect 20035 77680 20075 77720
rect 1468 77596 1508 77636
rect 14572 77596 14612 77636
rect 19852 77596 19892 77636
rect 1228 77512 1268 77552
rect 1612 77512 1652 77552
rect 12556 77512 12596 77552
rect 12748 77512 12788 77552
rect 15052 77512 15092 77552
rect 16012 77512 16052 77552
rect 2188 77428 2228 77468
rect 3436 77428 3476 77468
rect 3820 77428 3860 77468
rect 5068 77428 5108 77468
rect 5740 77428 5780 77468
rect 6988 77428 7028 77468
rect 7564 77428 7604 77468
rect 8812 77428 8852 77468
rect 9100 77428 9140 77468
rect 10348 77428 10388 77468
rect 10732 77428 10772 77468
rect 11980 77428 12020 77468
rect 13132 77428 13172 77468
rect 14380 77428 14420 77468
rect 15523 77428 15563 77468
rect 15628 77428 15668 77468
rect 16108 77428 16148 77468
rect 16588 77428 16628 77468
rect 17107 77428 17147 77468
rect 17644 77428 17684 77468
rect 18892 77428 18932 77468
rect 19180 77428 19220 77468
rect 19459 77428 19499 77468
rect 20030 77428 20070 77468
rect 20332 77428 20372 77468
rect 12316 77344 12356 77384
rect 12988 77344 13028 77384
rect 17452 77344 17492 77384
rect 19564 77344 19604 77384
rect 1852 77260 1892 77300
rect 3628 77260 3668 77300
rect 5260 77260 5300 77300
rect 7180 77260 7220 77300
rect 7372 77260 7412 77300
rect 12172 77260 12212 77300
rect 17260 77260 17300 77300
rect 20236 77260 20276 77300
rect 4928 77092 4968 77132
rect 5010 77092 5050 77132
rect 5092 77092 5132 77132
rect 5174 77092 5214 77132
rect 5256 77092 5296 77132
rect 20048 77092 20088 77132
rect 20130 77092 20170 77132
rect 20212 77092 20252 77132
rect 20294 77092 20334 77132
rect 20376 77092 20416 77132
rect 4876 76924 4916 76964
rect 10204 76924 10244 76964
rect 15244 76924 15284 76964
rect 15772 76924 15812 76964
rect 19996 76924 20036 76964
rect 10972 76840 11012 76880
rect 13036 76840 13076 76880
rect 15676 76840 15716 76880
rect 1420 76756 1460 76796
rect 2668 76747 2708 76787
rect 3139 76756 3179 76796
rect 3244 76756 3284 76796
rect 3628 76756 3668 76796
rect 4204 76747 4244 76787
rect 4684 76747 4724 76787
rect 6124 76756 6164 76796
rect 6307 76756 6347 76796
rect 6412 76756 6452 76796
rect 6604 76756 6644 76796
rect 7852 76747 7892 76787
rect 8323 76756 8363 76796
rect 8428 76756 8468 76796
rect 8812 76756 8852 76796
rect 9388 76747 9428 76787
rect 9868 76747 9908 76787
rect 11596 76756 11636 76796
rect 12844 76747 12884 76787
rect 13507 76756 13547 76796
rect 13612 76756 13652 76796
rect 13996 76756 14036 76796
rect 14572 76747 14612 76787
rect 15052 76747 15092 76787
rect 16204 76756 16244 76796
rect 17452 76747 17492 76787
rect 18220 76756 18260 76796
rect 19468 76747 19508 76787
rect 19852 76756 19892 76796
rect 3724 76672 3764 76712
rect 5068 76672 5108 76712
rect 5644 76672 5684 76712
rect 8908 76672 8948 76712
rect 10099 76672 10139 76712
rect 10444 76672 10484 76712
rect 10588 76672 10628 76712
rect 11212 76672 11252 76712
rect 14092 76672 14132 76712
rect 15436 76672 15476 76712
rect 16012 76672 16052 76712
rect 17836 76672 17876 76712
rect 20140 76672 20180 76712
rect 20380 76672 20420 76712
rect 5404 76588 5444 76628
rect 8044 76588 8084 76628
rect 10876 76588 10916 76628
rect 18076 76588 18116 76628
rect 2860 76504 2900 76544
rect 5308 76504 5348 76544
rect 6412 76504 6452 76544
rect 17644 76504 17684 76544
rect 19660 76504 19700 76544
rect 3688 76336 3728 76376
rect 3770 76336 3810 76376
rect 3852 76336 3892 76376
rect 3934 76336 3974 76376
rect 4016 76336 4056 76376
rect 18808 76336 18848 76376
rect 18890 76336 18930 76376
rect 18972 76336 19012 76376
rect 19054 76336 19094 76376
rect 19136 76336 19176 76376
rect 5980 76168 6020 76208
rect 8332 76168 8372 76208
rect 9964 76168 10004 76208
rect 11932 76168 11972 76208
rect 18364 76168 18404 76208
rect 11692 76084 11732 76124
rect 2860 76000 2900 76040
rect 3916 76000 3956 76040
rect 5548 76000 5588 76040
rect 5740 76000 5780 76040
rect 6124 76000 6164 76040
rect 6508 76000 6548 76040
rect 13132 76000 13172 76040
rect 18124 76000 18164 76040
rect 20140 76000 20180 76040
rect 1228 75916 1268 75956
rect 2476 75916 2516 75956
rect 3406 75916 3446 75956
rect 3532 75916 3572 75956
rect 4012 75916 4052 75956
rect 4492 75916 4532 75956
rect 5011 75916 5051 75956
rect 6892 75916 6932 75956
rect 8140 75916 8180 75956
rect 8524 75916 8564 75956
rect 9772 75916 9812 75956
rect 10252 75916 10292 75956
rect 11500 75916 11540 75956
rect 12163 75916 12203 75956
rect 12657 75916 12697 75956
rect 13228 75916 13268 75956
rect 13612 75916 13652 75956
rect 13725 75916 13765 75956
rect 14092 75916 14132 75956
rect 15340 75916 15380 75956
rect 15724 75916 15764 75956
rect 16972 75916 17012 75956
rect 17347 75916 17387 75956
rect 17491 75916 17531 75956
rect 17631 75916 17671 75956
rect 17731 75916 17771 75956
rect 17865 75916 17905 75956
rect 18508 75916 18548 75956
rect 19756 75916 19796 75956
rect 2668 75748 2708 75788
rect 3100 75748 3140 75788
rect 5164 75748 5204 75788
rect 5308 75748 5348 75788
rect 6364 75748 6404 75788
rect 6748 75748 6788 75788
rect 15532 75748 15572 75788
rect 17164 75748 17204 75788
rect 17548 75748 17588 75788
rect 19948 75748 19988 75788
rect 20380 75748 20420 75788
rect 4928 75580 4968 75620
rect 5010 75580 5050 75620
rect 5092 75580 5132 75620
rect 5174 75580 5214 75620
rect 5256 75580 5296 75620
rect 20048 75580 20088 75620
rect 20130 75580 20170 75620
rect 20212 75580 20252 75620
rect 20294 75580 20334 75620
rect 20376 75580 20416 75620
rect 2236 75412 2276 75452
rect 9004 75412 9044 75452
rect 11164 75412 11204 75452
rect 14044 75412 14084 75452
rect 16684 75412 16724 75452
rect 10732 75328 10772 75368
rect 2668 75244 2708 75284
rect 3916 75235 3956 75275
rect 4684 75244 4724 75284
rect 5932 75235 5972 75275
rect 6316 75244 6356 75284
rect 7564 75235 7604 75275
rect 7939 75244 7979 75284
rect 8044 75235 8084 75275
rect 8188 75235 8228 75275
rect 8362 75244 8402 75284
rect 8500 75244 8540 75284
rect 8716 75244 8756 75284
rect 8858 75244 8898 75284
rect 9292 75244 9332 75284
rect 10540 75235 10580 75275
rect 14947 75244 14987 75284
rect 15052 75244 15092 75284
rect 15436 75244 15476 75284
rect 16012 75235 16052 75275
rect 16492 75235 16532 75275
rect 16876 75244 16916 75284
rect 18124 75235 18164 75275
rect 18892 75244 18932 75284
rect 20140 75235 20180 75275
rect 1228 75160 1268 75200
rect 1612 75160 1652 75200
rect 1996 75160 2036 75200
rect 4492 75160 4532 75200
rect 10924 75160 10964 75200
rect 12748 75160 12788 75200
rect 12940 75160 12980 75200
rect 13180 75160 13220 75200
rect 13324 75160 13364 75200
rect 13708 75160 13748 75200
rect 14284 75160 14324 75200
rect 14476 75160 14516 75200
rect 15532 75160 15572 75200
rect 18508 75160 18548 75200
rect 4252 75076 4292 75116
rect 13564 75076 13604 75116
rect 13948 75076 13988 75116
rect 1468 74992 1508 75032
rect 1852 74992 1892 75032
rect 4108 74992 4148 75032
rect 6124 74992 6164 75032
rect 7756 74992 7796 75032
rect 7939 74992 7979 75032
rect 12508 74992 12548 75032
rect 14716 74992 14756 75032
rect 18316 74992 18356 75032
rect 18748 74992 18788 75032
rect 20332 74992 20372 75032
rect 3688 74824 3728 74864
rect 3770 74824 3810 74864
rect 3852 74824 3892 74864
rect 3934 74824 3974 74864
rect 4016 74824 4056 74864
rect 18808 74824 18848 74864
rect 18890 74824 18930 74864
rect 18972 74824 19012 74864
rect 19054 74824 19094 74864
rect 19136 74824 19176 74864
rect 5500 74656 5540 74696
rect 11692 74656 11732 74696
rect 17356 74656 17396 74696
rect 17692 74656 17732 74696
rect 10060 74572 10100 74612
rect 2860 74488 2900 74528
rect 3916 74488 3956 74528
rect 6220 74488 6260 74528
rect 7852 74488 7892 74528
rect 8428 74488 8468 74528
rect 13612 74488 13652 74528
rect 14860 74488 14900 74528
rect 18412 74488 18452 74528
rect 20140 74488 20180 74528
rect 1228 74404 1268 74444
rect 2476 74404 2516 74444
rect 3427 74404 3467 74444
rect 3532 74404 3572 74444
rect 4012 74404 4052 74444
rect 4492 74404 4532 74444
rect 5011 74404 5051 74444
rect 5356 74404 5396 74444
rect 5731 74404 5771 74444
rect 5836 74404 5876 74444
rect 6316 74404 6356 74444
rect 6796 74404 6836 74444
rect 7284 74404 7324 74444
rect 8620 74404 8660 74444
rect 9868 74404 9908 74444
rect 10252 74404 10292 74444
rect 11500 74404 11540 74444
rect 11980 74404 12020 74444
rect 13228 74404 13268 74444
rect 14371 74404 14411 74444
rect 14476 74404 14516 74444
rect 14956 74404 14996 74444
rect 15436 74404 15476 74444
rect 15924 74404 15964 74444
rect 16732 74404 16772 74444
rect 16876 74404 16916 74444
rect 17059 74430 17099 74470
rect 17251 74404 17291 74444
rect 17356 74404 17396 74444
rect 17548 74404 17588 74444
rect 17923 74404 17963 74444
rect 18028 74404 18068 74444
rect 18508 74404 18548 74444
rect 18988 74404 19028 74444
rect 19507 74404 19547 74444
rect 8092 74320 8132 74360
rect 13852 74320 13892 74360
rect 2668 74236 2708 74276
rect 3100 74236 3140 74276
rect 5164 74236 5204 74276
rect 7468 74236 7508 74276
rect 8188 74236 8228 74276
rect 13420 74236 13460 74276
rect 16108 74236 16148 74276
rect 16579 74236 16619 74276
rect 19660 74236 19700 74276
rect 20380 74236 20420 74276
rect 4928 74068 4968 74108
rect 5010 74068 5050 74108
rect 5092 74068 5132 74108
rect 5174 74068 5214 74108
rect 5256 74068 5296 74108
rect 20048 74068 20088 74108
rect 20130 74068 20170 74108
rect 20212 74068 20252 74108
rect 20294 74068 20334 74108
rect 20376 74068 20416 74108
rect 4780 73900 4820 73940
rect 6604 73900 6644 73940
rect 12220 73900 12260 73940
rect 14476 73900 14516 73940
rect 12076 73816 12116 73856
rect 1324 73732 1364 73772
rect 2572 73723 2612 73763
rect 3043 73732 3083 73772
rect 3148 73732 3188 73772
rect 3532 73732 3572 73772
rect 4108 73723 4148 73763
rect 4588 73723 4628 73763
rect 5164 73732 5204 73772
rect 6412 73723 6452 73763
rect 6979 73732 7019 73772
rect 7468 73723 7508 73763
rect 7948 73732 7988 73772
rect 8428 73732 8468 73772
rect 8529 73732 8569 73772
rect 9004 73732 9044 73772
rect 10252 73732 10292 73772
rect 10636 73732 10676 73772
rect 11884 73723 11924 73763
rect 12739 73732 12779 73772
rect 12844 73732 12884 73772
rect 13228 73732 13268 73772
rect 13804 73723 13844 73763
rect 14284 73723 14324 73763
rect 16396 73732 16436 73772
rect 17644 73723 17684 73763
rect 18604 73732 18644 73772
rect 19852 73723 19892 73763
rect 20332 73732 20372 73772
rect 3628 73648 3668 73688
rect 6748 73648 6788 73688
rect 8044 73648 8084 73688
rect 12460 73648 12500 73688
rect 13324 73648 13364 73688
rect 14860 73648 14900 73688
rect 15100 73648 15140 73688
rect 15484 73648 15524 73688
rect 15724 73648 15764 73688
rect 15916 73648 15956 73688
rect 18220 73648 18260 73688
rect 15388 73564 15428 73604
rect 20188 73564 20228 73604
rect 2764 73480 2804 73520
rect 8812 73480 8852 73520
rect 14620 73480 14660 73520
rect 16156 73480 16196 73520
rect 17836 73480 17876 73520
rect 18460 73480 18500 73520
rect 20044 73480 20084 73520
rect 3688 73312 3728 73352
rect 3770 73312 3810 73352
rect 3852 73312 3892 73352
rect 3934 73312 3974 73352
rect 4016 73312 4056 73352
rect 18808 73312 18848 73352
rect 18890 73312 18930 73352
rect 18972 73312 19012 73352
rect 19054 73312 19094 73352
rect 19136 73312 19176 73352
rect 4828 73144 4868 73184
rect 6940 73144 6980 73184
rect 17452 73144 17492 73184
rect 19267 73144 19307 73184
rect 15484 73060 15524 73100
rect 19084 73060 19124 73100
rect 4588 72976 4628 73016
rect 6700 72976 6740 73016
rect 8188 72976 8228 73016
rect 8331 72976 8371 73016
rect 13420 72976 13460 73016
rect 14860 72976 14900 73016
rect 15244 72976 15284 73016
rect 15628 72976 15668 73016
rect 20140 72976 20180 73016
rect 1324 72892 1364 72932
rect 2572 72892 2612 72932
rect 2956 72892 2996 72932
rect 4204 72892 4244 72932
rect 4972 72892 5012 72932
rect 6220 72892 6260 72932
rect 7267 72892 7307 72932
rect 7756 72892 7796 72932
rect 8716 72892 8756 72932
rect 8834 72892 8874 72932
rect 9580 72892 9620 72932
rect 10828 72892 10868 72932
rect 11020 72892 11060 72932
rect 12268 72892 12308 72932
rect 12931 72892 12971 72932
rect 13036 72892 13076 72932
rect 13516 72892 13556 72932
rect 13996 72892 14036 72932
rect 14515 72892 14555 72932
rect 16012 72892 16052 72932
rect 17260 72892 17300 72932
rect 17644 72892 17684 72932
rect 18892 72892 18932 72932
rect 19267 72892 19307 72932
rect 19372 72903 19412 72943
rect 19517 72892 19557 72932
rect 19647 72892 19687 72932
rect 19777 72903 19817 72943
rect 7075 72808 7115 72848
rect 12460 72808 12500 72848
rect 15100 72808 15140 72848
rect 2764 72724 2804 72764
rect 4396 72724 4436 72764
rect 6412 72724 6452 72764
rect 9388 72724 9428 72764
rect 14668 72724 14708 72764
rect 15868 72724 15908 72764
rect 17452 72724 17492 72764
rect 19084 72724 19124 72764
rect 20380 72724 20420 72764
rect 4928 72556 4968 72596
rect 5010 72556 5050 72596
rect 5092 72556 5132 72596
rect 5174 72556 5214 72596
rect 5256 72556 5296 72596
rect 20048 72556 20088 72596
rect 20130 72556 20170 72596
rect 20212 72556 20252 72596
rect 20294 72556 20334 72596
rect 20376 72556 20416 72596
rect 10492 72388 10532 72428
rect 11260 72388 11300 72428
rect 15052 72388 15092 72428
rect 17155 72388 17195 72428
rect 20140 72388 20180 72428
rect 2332 72304 2372 72344
rect 5116 72304 5156 72344
rect 5500 72304 5540 72344
rect 10108 72304 10148 72344
rect 2851 72220 2891 72260
rect 2956 72220 2996 72260
rect 3340 72220 3380 72260
rect 3916 72211 3956 72251
rect 4396 72211 4436 72251
rect 4627 72220 4667 72260
rect 6286 72220 6326 72260
rect 6412 72220 6452 72260
rect 6796 72220 6836 72260
rect 7372 72211 7412 72251
rect 7852 72211 7892 72251
rect 11980 72220 12020 72260
rect 13228 72211 13268 72251
rect 13612 72220 13652 72260
rect 14860 72211 14900 72251
rect 15244 72220 15284 72260
rect 16492 72211 16532 72251
rect 17308 72220 17348 72260
rect 17452 72220 17492 72260
rect 17644 72220 17684 72260
rect 17827 72220 17867 72260
rect 17932 72220 17972 72260
rect 18382 72220 18422 72260
rect 18513 72220 18553 72260
rect 18892 72220 18932 72260
rect 19468 72211 19508 72251
rect 19948 72211 19988 72251
rect 1420 72136 1460 72176
rect 1804 72136 1844 72176
rect 2188 72136 2228 72176
rect 2572 72136 2612 72176
rect 3436 72136 3476 72176
rect 4732 72136 4772 72176
rect 4972 72136 5012 72176
rect 5356 72136 5396 72176
rect 5740 72136 5780 72176
rect 6892 72136 6932 72176
rect 8083 72136 8123 72176
rect 8428 72136 8468 72176
rect 8620 72136 8660 72176
rect 8956 72136 8996 72176
rect 9196 72136 9236 72176
rect 9388 72136 9428 72176
rect 9964 72136 10004 72176
rect 10348 72136 10388 72176
rect 10732 72136 10772 72176
rect 11500 72136 11540 72176
rect 18988 72136 19028 72176
rect 1180 72052 1220 72092
rect 1564 72052 1604 72092
rect 1948 72052 1988 72092
rect 8188 72052 8228 72092
rect 8860 72052 8900 72092
rect 9628 72052 9668 72092
rect 17932 72052 17972 72092
rect 9724 71968 9764 72008
rect 13420 71968 13460 72008
rect 16684 71968 16724 72008
rect 3688 71800 3728 71840
rect 3770 71800 3810 71840
rect 3852 71800 3892 71840
rect 3934 71800 3974 71840
rect 4016 71800 4056 71840
rect 18808 71800 18848 71840
rect 18890 71800 18930 71840
rect 18972 71800 19012 71840
rect 19054 71800 19094 71840
rect 19136 71800 19176 71840
rect 2140 71632 2180 71672
rect 8140 71632 8180 71672
rect 1420 71464 1460 71504
rect 1900 71464 1940 71504
rect 2284 71464 2324 71504
rect 3340 71464 3380 71504
rect 12460 71464 12500 71504
rect 13747 71464 13787 71504
rect 14092 71464 14132 71504
rect 14764 71464 14804 71504
rect 15532 71464 15572 71504
rect 17260 71464 17300 71504
rect 17644 71464 17684 71504
rect 18604 71464 18644 71504
rect 20140 71464 20180 71504
rect 2830 71380 2870 71420
rect 2956 71380 2996 71420
rect 3436 71380 3476 71420
rect 3916 71380 3956 71420
rect 4404 71380 4444 71420
rect 4780 71380 4820 71420
rect 6028 71380 6068 71420
rect 6700 71380 6740 71420
rect 7948 71380 7988 71420
rect 8620 71380 8660 71420
rect 9868 71380 9908 71420
rect 10252 71380 10292 71420
rect 11500 71380 11540 71420
rect 11971 71380 12011 71420
rect 12076 71380 12116 71420
rect 12556 71380 12596 71420
rect 13036 71380 13076 71420
rect 13524 71380 13564 71420
rect 15043 71380 15083 71420
rect 15148 71380 15188 71420
rect 15628 71380 15668 71420
rect 16108 71380 16148 71420
rect 16627 71380 16667 71420
rect 18115 71380 18155 71420
rect 18220 71380 18260 71420
rect 18700 71380 18740 71420
rect 19180 71380 19220 71420
rect 19699 71380 19739 71420
rect 2524 71296 2564 71336
rect 11692 71296 11732 71336
rect 1180 71212 1220 71252
rect 4588 71212 4628 71252
rect 6220 71212 6260 71252
rect 10060 71212 10100 71252
rect 13852 71212 13892 71252
rect 14524 71212 14564 71252
rect 16780 71212 16820 71252
rect 17500 71212 17540 71252
rect 17884 71212 17924 71252
rect 19852 71212 19892 71252
rect 20380 71212 20420 71252
rect 4928 71044 4968 71084
rect 5010 71044 5050 71084
rect 5092 71044 5132 71084
rect 5174 71044 5214 71084
rect 5256 71044 5296 71084
rect 20048 71044 20088 71084
rect 20130 71044 20170 71084
rect 20212 71044 20252 71084
rect 20294 71044 20334 71084
rect 20376 71044 20416 71084
rect 1564 70876 1604 70916
rect 7468 70876 7508 70916
rect 13420 70876 13460 70916
rect 15244 70876 15284 70916
rect 18364 70876 18404 70916
rect 10924 70792 10964 70832
rect 1996 70708 2036 70748
rect 3244 70699 3284 70739
rect 4387 70708 4427 70748
rect 4492 70708 4532 70748
rect 4876 70708 4916 70748
rect 5452 70699 5492 70739
rect 5932 70699 5972 70739
rect 7180 70708 7220 70748
rect 7322 70708 7362 70748
rect 7852 70699 7892 70739
rect 9100 70708 9140 70748
rect 9484 70708 9524 70748
rect 10732 70699 10772 70739
rect 11683 70708 11723 70748
rect 11788 70708 11828 70748
rect 12172 70708 12212 70748
rect 12748 70699 12788 70739
rect 13228 70699 13268 70739
rect 13804 70708 13844 70748
rect 15052 70699 15092 70739
rect 16108 70708 16148 70748
rect 17356 70699 17396 70739
rect 18796 70708 18836 70748
rect 20044 70699 20084 70739
rect 1420 70624 1460 70664
rect 1804 70624 1844 70664
rect 3820 70624 3860 70664
rect 4972 70624 5012 70664
rect 6316 70624 6356 70664
rect 6892 70624 6932 70664
rect 11068 70624 11108 70664
rect 11308 70624 11348 70664
rect 12268 70624 12308 70664
rect 15916 70624 15956 70664
rect 18028 70624 18068 70664
rect 18604 70624 18644 70664
rect 1180 70540 1220 70580
rect 3580 70540 3620 70580
rect 6172 70540 6212 70580
rect 6652 70540 6692 70580
rect 15676 70540 15716 70580
rect 18268 70540 18308 70580
rect 20236 70540 20276 70580
rect 3436 70456 3476 70496
rect 6556 70456 6596 70496
rect 7660 70456 7700 70496
rect 17548 70456 17588 70496
rect 3688 70288 3728 70328
rect 3770 70288 3810 70328
rect 3852 70288 3892 70328
rect 3934 70288 3974 70328
rect 4016 70288 4056 70328
rect 18808 70288 18848 70328
rect 18890 70288 18930 70328
rect 18972 70288 19012 70328
rect 19054 70288 19094 70328
rect 19136 70288 19176 70328
rect 12604 70120 12644 70160
rect 16060 70120 16100 70160
rect 17404 70120 17444 70160
rect 16732 70036 16772 70076
rect 3532 69952 3572 69992
rect 8140 69952 8180 69992
rect 9196 69952 9236 69992
rect 9571 69952 9611 69992
rect 11212 69952 11252 69992
rect 12364 69952 12404 69992
rect 16300 69952 16340 69992
rect 16972 69952 17012 69992
rect 17164 69952 17204 69992
rect 18124 69952 18164 69992
rect 19756 69952 19796 69992
rect 20140 69952 20180 69992
rect 1516 69868 1556 69908
rect 2764 69868 2804 69908
rect 3916 69868 3956 69908
rect 5164 69868 5204 69908
rect 5356 69868 5396 69908
rect 6604 69868 6644 69908
rect 7171 69868 7211 69908
rect 7660 69868 7700 69908
rect 8236 69868 8276 69908
rect 8620 69868 8660 69908
rect 8738 69868 8778 69908
rect 9772 69868 9812 69908
rect 11020 69868 11060 69908
rect 12748 69868 12788 69908
rect 13996 69868 14036 69908
rect 14476 69868 14516 69908
rect 15724 69868 15764 69908
rect 17614 69868 17654 69908
rect 17740 69868 17780 69908
rect 18220 69868 18260 69908
rect 18700 69868 18740 69908
rect 19219 69868 19259 69908
rect 19996 69784 20036 69824
rect 2956 69700 2996 69740
rect 3292 69700 3332 69740
rect 3724 69700 3764 69740
rect 6796 69700 6836 69740
rect 6988 69700 7028 69740
rect 8956 69700 8996 69740
rect 11452 69700 11492 69740
rect 14188 69700 14228 69740
rect 15916 69700 15956 69740
rect 19372 69700 19412 69740
rect 20380 69700 20420 69740
rect 4928 69532 4968 69572
rect 5010 69532 5050 69572
rect 5092 69532 5132 69572
rect 5174 69532 5214 69572
rect 5256 69532 5296 69572
rect 20048 69532 20088 69572
rect 20130 69532 20170 69572
rect 20212 69532 20252 69572
rect 20294 69532 20334 69572
rect 20376 69532 20416 69572
rect 4876 69364 4916 69404
rect 7555 69364 7595 69404
rect 16012 69364 16052 69404
rect 20044 69364 20084 69404
rect 5020 69280 5060 69320
rect 7843 69271 7883 69311
rect 10684 69280 10724 69320
rect 18028 69280 18068 69320
rect 1420 69196 1460 69236
rect 2668 69187 2708 69227
rect 3118 69196 3158 69236
rect 3244 69196 3284 69236
rect 3628 69196 3668 69236
rect 4204 69187 4244 69227
rect 4684 69187 4724 69227
rect 5452 69196 5492 69236
rect 5635 69196 5675 69236
rect 5740 69196 5780 69236
rect 5932 69196 5972 69236
rect 7180 69187 7220 69227
rect 7555 69196 7595 69236
rect 7660 69187 7700 69227
rect 7939 69196 7979 69236
rect 8073 69196 8113 69236
rect 8428 69196 8468 69236
rect 9676 69187 9716 69227
rect 11500 69196 11540 69236
rect 12748 69187 12788 69227
rect 14275 69196 14315 69236
rect 14380 69196 14420 69236
rect 14860 69196 14900 69236
rect 15340 69187 15380 69227
rect 15820 69187 15860 69227
rect 16588 69196 16628 69236
rect 17836 69187 17876 69227
rect 18307 69196 18347 69236
rect 18412 69196 18452 69236
rect 18796 69196 18836 69236
rect 19372 69187 19412 69227
rect 19852 69187 19892 69227
rect 3724 69112 3764 69152
rect 5260 69112 5300 69152
rect 10252 69112 10292 69152
rect 10444 69112 10484 69152
rect 13324 69112 13364 69152
rect 13804 69112 13844 69152
rect 14044 69112 14084 69152
rect 14764 69112 14804 69152
rect 16156 69112 16196 69152
rect 16396 69112 16436 69152
rect 18892 69112 18932 69152
rect 7372 69028 7412 69068
rect 13564 69028 13604 69068
rect 2860 68944 2900 68984
rect 5740 68944 5780 68984
rect 9868 68944 9908 68984
rect 10012 68944 10052 68984
rect 12940 68944 12980 68984
rect 3688 68776 3728 68816
rect 3770 68776 3810 68816
rect 3852 68776 3892 68816
rect 3934 68776 3974 68816
rect 4016 68776 4056 68816
rect 18808 68776 18848 68816
rect 18890 68776 18930 68816
rect 18972 68776 19012 68816
rect 19054 68776 19094 68816
rect 19136 68776 19176 68816
rect 3196 68608 3236 68648
rect 10012 68608 10052 68648
rect 16828 68608 16868 68648
rect 18988 68608 19028 68648
rect 2812 68524 2852 68564
rect 19420 68524 19460 68564
rect 3052 68440 3092 68480
rect 3436 68440 3476 68480
rect 4300 68440 4340 68480
rect 7372 68440 7412 68480
rect 8332 68440 8372 68480
rect 8467 68440 8507 68480
rect 9772 68440 9812 68480
rect 12748 68440 12788 68480
rect 14035 68440 14075 68480
rect 14380 68440 14420 68480
rect 15340 68440 15380 68480
rect 17068 68440 17108 68480
rect 19660 68440 19700 68480
rect 20140 68440 20180 68480
rect 1228 68356 1268 68396
rect 2476 68356 2516 68396
rect 3811 68356 3851 68396
rect 3916 68356 3956 68396
rect 4396 68356 4436 68396
rect 4876 68356 4916 68396
rect 5395 68356 5435 68396
rect 5932 68356 5972 68396
rect 7180 68356 7220 68396
rect 7843 68356 7883 68396
rect 7948 68356 7988 68396
rect 8908 68356 8948 68396
rect 9427 68356 9467 68396
rect 10444 68356 10484 68396
rect 11692 68356 11732 68396
rect 12259 68356 12299 68396
rect 12364 68356 12404 68396
rect 12844 68356 12884 68396
rect 13324 68356 13364 68396
rect 13812 68356 13852 68396
rect 14851 68356 14891 68396
rect 14956 68356 14996 68396
rect 15436 68356 15476 68396
rect 15916 68356 15956 68396
rect 16404 68356 16444 68396
rect 17548 68356 17588 68396
rect 18796 68356 18836 68396
rect 5740 68272 5780 68312
rect 11884 68272 11924 68312
rect 2668 68188 2708 68228
rect 5548 68188 5588 68228
rect 7612 68188 7652 68228
rect 9580 68188 9620 68228
rect 14140 68188 14180 68228
rect 16588 68188 16628 68228
rect 20380 68188 20420 68228
rect 4928 68020 4968 68060
rect 5010 68020 5050 68060
rect 5092 68020 5132 68060
rect 5174 68020 5214 68060
rect 5256 68020 5296 68060
rect 20048 68020 20088 68060
rect 20130 68020 20170 68060
rect 20212 68020 20252 68060
rect 20294 68020 20334 68060
rect 20376 68020 20416 68060
rect 16204 67852 16244 67892
rect 1324 67684 1364 67724
rect 2572 67675 2612 67715
rect 3043 67684 3083 67724
rect 3148 67684 3188 67724
rect 3532 67684 3572 67724
rect 4108 67675 4148 67715
rect 4588 67675 4628 67715
rect 5356 67684 5396 67724
rect 5644 67684 5684 67724
rect 6892 67675 6932 67715
rect 7372 67684 7412 67724
rect 8620 67675 8660 67715
rect 9484 67684 9524 67724
rect 10732 67675 10772 67715
rect 11116 67684 11156 67724
rect 12364 67675 12404 67715
rect 12748 67684 12788 67724
rect 13996 67675 14036 67715
rect 14764 67684 14804 67724
rect 16012 67675 16052 67715
rect 16972 67684 17012 67724
rect 18220 67675 18260 67715
rect 18604 67684 18644 67724
rect 19852 67675 19892 67715
rect 3628 67600 3668 67640
rect 5164 67600 5204 67640
rect 9004 67600 9044 67640
rect 9244 67600 9284 67640
rect 14380 67600 14420 67640
rect 16588 67600 16628 67640
rect 16828 67600 16868 67640
rect 4828 67516 4868 67556
rect 5500 67516 5540 67556
rect 14188 67516 14228 67556
rect 2764 67432 2804 67472
rect 4924 67432 4964 67472
rect 7084 67432 7124 67472
rect 8812 67432 8852 67472
rect 10924 67432 10964 67472
rect 12556 67432 12596 67472
rect 14620 67432 14660 67472
rect 18412 67432 18452 67472
rect 20044 67432 20084 67472
rect 3688 67264 3728 67304
rect 3770 67264 3810 67304
rect 3852 67264 3892 67304
rect 3934 67264 3974 67304
rect 4016 67264 4056 67304
rect 18808 67264 18848 67304
rect 18890 67264 18930 67304
rect 18972 67264 19012 67304
rect 19054 67264 19094 67304
rect 19136 67264 19176 67304
rect 8956 67096 8996 67136
rect 13372 67096 13412 67136
rect 15484 67096 15524 67136
rect 5212 67012 5252 67052
rect 15868 67012 15908 67052
rect 1420 66928 1460 66968
rect 4972 66928 5012 66968
rect 7564 66928 7604 66968
rect 9196 66928 9236 66968
rect 11692 66928 11732 66968
rect 13132 66928 13172 66968
rect 15244 66928 15284 66968
rect 15628 66928 15668 66968
rect 16012 66928 16052 66968
rect 18604 66928 18644 66968
rect 20236 66928 20276 66968
rect 1708 66844 1748 66884
rect 2956 66844 2996 66884
rect 3532 66844 3572 66884
rect 4780 66844 4820 66884
rect 5356 66844 5396 66884
rect 6604 66844 6644 66884
rect 7075 66844 7115 66884
rect 7180 66844 7220 66884
rect 7660 66844 7700 66884
rect 8140 66844 8180 66884
rect 8659 66844 8699 66884
rect 9484 66844 9524 66884
rect 10732 66844 10772 66884
rect 11203 66844 11243 66884
rect 11308 66844 11348 66884
rect 11788 66844 11828 66884
rect 12268 66844 12308 66884
rect 12756 66844 12796 66884
rect 13612 66844 13652 66884
rect 14860 66844 14900 66884
rect 16396 66844 16436 66884
rect 17644 66844 17684 66884
rect 18115 66844 18155 66884
rect 18220 66844 18260 66884
rect 18700 66844 18740 66884
rect 19180 66844 19220 66884
rect 19699 66844 19739 66884
rect 6796 66760 6836 66800
rect 1180 66676 1220 66716
rect 3148 66676 3188 66716
rect 3340 66676 3380 66716
rect 8812 66676 8852 66716
rect 10924 66676 10964 66716
rect 12940 66676 12980 66716
rect 15052 66676 15092 66716
rect 16252 66676 16292 66716
rect 17836 66676 17876 66716
rect 19852 66676 19892 66716
rect 19996 66676 20036 66716
rect 4928 66508 4968 66548
rect 5010 66508 5050 66548
rect 5092 66508 5132 66548
rect 5174 66508 5214 66548
rect 5256 66508 5296 66548
rect 20048 66508 20088 66548
rect 20130 66508 20170 66548
rect 20212 66508 20252 66548
rect 20294 66508 20334 66548
rect 20376 66508 20416 66548
rect 4396 66340 4436 66380
rect 17116 66340 17156 66380
rect 20332 66340 20372 66380
rect 6844 66256 6884 66296
rect 16732 66256 16772 66296
rect 2638 66172 2678 66212
rect 2764 66172 2804 66212
rect 3148 66172 3188 66212
rect 3724 66163 3764 66203
rect 4204 66163 4244 66203
rect 4780 66172 4820 66212
rect 6028 66163 6068 66203
rect 7948 66172 7988 66212
rect 9196 66163 9236 66203
rect 9868 66172 9908 66212
rect 11116 66163 11156 66203
rect 13036 66172 13076 66212
rect 14284 66163 14324 66203
rect 14851 66172 14891 66212
rect 14956 66172 14996 66212
rect 15340 66172 15380 66212
rect 15916 66163 15956 66203
rect 16396 66163 16436 66203
rect 18211 66172 18251 66212
rect 18316 66172 18356 66212
rect 18700 66172 18740 66212
rect 19276 66163 19316 66203
rect 19756 66163 19796 66203
rect 1420 66088 1460 66128
rect 1804 66088 1844 66128
rect 2188 66088 2228 66128
rect 3244 66088 3284 66128
rect 6643 66088 6683 66128
rect 6988 66088 7028 66128
rect 7564 66088 7604 66128
rect 12844 66088 12884 66128
rect 15436 66088 15476 66128
rect 16627 66088 16667 66128
rect 16972 66088 17012 66128
rect 17356 66088 17396 66128
rect 17740 66088 17780 66128
rect 18796 66088 18836 66128
rect 7228 66004 7268 66044
rect 14476 66004 14516 66044
rect 19996 66004 20036 66044
rect 1180 65920 1220 65960
rect 1564 65920 1604 65960
rect 1948 65920 1988 65960
rect 6220 65920 6260 65960
rect 7324 65920 7364 65960
rect 9388 65920 9428 65960
rect 11308 65920 11348 65960
rect 12604 65920 12644 65960
rect 17980 65920 18020 65960
rect 3688 65752 3728 65792
rect 3770 65752 3810 65792
rect 3852 65752 3892 65792
rect 3934 65752 3974 65792
rect 4016 65752 4056 65792
rect 18808 65752 18848 65792
rect 18890 65752 18930 65792
rect 18972 65752 19012 65792
rect 19054 65752 19094 65792
rect 19136 65752 19176 65792
rect 3100 65584 3140 65624
rect 12028 65584 12068 65624
rect 16915 65584 16955 65624
rect 20140 65584 20180 65624
rect 17068 65500 17108 65540
rect 3340 65416 3380 65456
rect 3724 65416 3764 65456
rect 4300 65416 4340 65456
rect 9964 65416 10004 65456
rect 11788 65416 11828 65456
rect 12124 65416 12164 65456
rect 12364 65416 12404 65456
rect 13132 65416 13172 65456
rect 14419 65416 14459 65456
rect 14764 65416 14804 65456
rect 15628 65416 15668 65456
rect 1516 65332 1556 65372
rect 2772 65332 2812 65372
rect 4492 65332 4532 65372
rect 5740 65332 5780 65372
rect 6124 65332 6164 65372
rect 7372 65332 7412 65372
rect 7756 65332 7796 65372
rect 9004 65332 9044 65372
rect 9475 65332 9515 65372
rect 9580 65332 9620 65372
rect 10060 65332 10100 65372
rect 10540 65332 10580 65372
rect 11028 65332 11068 65372
rect 12643 65332 12683 65372
rect 12748 65332 12788 65372
rect 13228 65332 13268 65372
rect 13708 65332 13748 65372
rect 14196 65332 14236 65372
rect 15118 65332 15158 65372
rect 15244 65331 15284 65371
rect 15724 65332 15764 65372
rect 16204 65332 16244 65372
rect 16692 65332 16732 65372
rect 17260 65332 17300 65372
rect 18508 65332 18548 65372
rect 18700 65332 18740 65372
rect 19948 65332 19988 65372
rect 3484 65248 3524 65288
rect 14524 65248 14564 65288
rect 2956 65164 2996 65204
rect 4060 65164 4100 65204
rect 5932 65164 5972 65204
rect 7564 65164 7604 65204
rect 9196 65164 9236 65204
rect 11212 65164 11252 65204
rect 12028 65164 12068 65204
rect 4928 64996 4968 65036
rect 5010 64996 5050 65036
rect 5092 64996 5132 65036
rect 5174 64996 5214 65036
rect 5256 64996 5296 65036
rect 20048 64996 20088 65036
rect 20130 64996 20170 65036
rect 20212 64996 20252 65036
rect 20294 64996 20334 65036
rect 20376 64996 20416 65036
rect 14092 64828 14132 64868
rect 16108 64828 16148 64868
rect 2179 64744 2219 64784
rect 8332 64744 8372 64784
rect 14524 64744 14564 64784
rect 2371 64660 2411 64700
rect 2860 64651 2900 64691
rect 3340 64660 3380 64700
rect 3820 64660 3860 64700
rect 3938 64660 3978 64700
rect 4291 64660 4331 64700
rect 4396 64660 4436 64700
rect 4780 64660 4820 64700
rect 5356 64651 5396 64691
rect 5836 64651 5876 64691
rect 6892 64660 6932 64700
rect 8140 64651 8180 64691
rect 8515 64660 8555 64700
rect 8812 64660 8852 64700
rect 9100 64660 9140 64700
rect 9571 64660 9611 64700
rect 9681 64660 9721 64700
rect 10060 64660 10100 64700
rect 10636 64651 10676 64691
rect 11116 64651 11156 64691
rect 12652 64660 12692 64700
rect 13900 64651 13940 64691
rect 14668 64660 14708 64700
rect 15916 64651 15956 64691
rect 16588 64660 16628 64700
rect 17836 64651 17876 64691
rect 18316 64660 18356 64700
rect 19564 64651 19604 64691
rect 1420 64576 1460 64616
rect 1804 64576 1844 64616
rect 3436 64576 3476 64616
rect 4876 64576 4916 64616
rect 6067 64576 6107 64616
rect 6412 64576 6452 64616
rect 10156 64576 10196 64616
rect 12268 64576 12308 64616
rect 12508 64576 12548 64616
rect 14284 64576 14324 64616
rect 20140 64576 20180 64616
rect 6172 64492 6212 64532
rect 8956 64492 8996 64532
rect 1180 64408 1220 64448
rect 1564 64408 1604 64448
rect 8812 64408 8852 64448
rect 11347 64408 11387 64448
rect 18028 64408 18068 64448
rect 19756 64408 19796 64448
rect 20380 64408 20420 64448
rect 3688 64240 3728 64280
rect 3770 64240 3810 64280
rect 3852 64240 3892 64280
rect 3934 64240 3974 64280
rect 4016 64240 4056 64280
rect 18808 64240 18848 64280
rect 18890 64240 18930 64280
rect 18972 64240 19012 64280
rect 19054 64240 19094 64280
rect 19136 64240 19176 64280
rect 5692 64072 5732 64112
rect 9436 64072 9476 64112
rect 15004 64072 15044 64112
rect 19996 64072 20036 64112
rect 2956 63988 2996 64028
rect 6076 63988 6116 64028
rect 15484 63988 15524 64028
rect 3340 63904 3380 63944
rect 3724 63904 3764 63944
rect 5932 63904 5972 63944
rect 6316 63904 6356 63944
rect 6700 63904 6740 63944
rect 9091 63904 9131 63944
rect 9676 63904 9716 63944
rect 11692 63904 11732 63944
rect 12556 63904 12596 63944
rect 14572 63904 14612 63944
rect 14764 63904 14804 63944
rect 15148 63904 15188 63944
rect 15724 63904 15764 63944
rect 16204 63904 16244 63944
rect 18604 63904 18644 63944
rect 20236 63904 20276 63944
rect 1516 63820 1556 63860
rect 2764 63820 2804 63860
rect 3916 63820 3956 63860
rect 5164 63820 5204 63860
rect 6892 63820 6932 63860
rect 8140 63820 8180 63860
rect 8515 63820 8555 63860
rect 8951 63820 8991 63860
rect 9196 63820 9236 63860
rect 10060 63820 10100 63860
rect 11308 63820 11348 63860
rect 12748 63820 12788 63860
rect 13996 63820 14036 63860
rect 16396 63820 16436 63860
rect 17644 63820 17684 63860
rect 18115 63820 18155 63860
rect 18220 63820 18260 63860
rect 18700 63820 18740 63860
rect 19180 63820 19220 63860
rect 19672 63820 19712 63860
rect 3100 63736 3140 63776
rect 6460 63736 6500 63776
rect 8826 63736 8866 63776
rect 11932 63736 11972 63776
rect 14332 63736 14372 63776
rect 15388 63736 15428 63776
rect 17836 63736 17876 63776
rect 3484 63652 3524 63692
rect 5356 63652 5396 63692
rect 8332 63652 8372 63692
rect 8611 63652 8651 63692
rect 8716 63652 8756 63692
rect 9283 63652 9323 63692
rect 11500 63652 11540 63692
rect 12316 63652 12356 63692
rect 14188 63652 14228 63692
rect 15964 63652 16004 63692
rect 19852 63652 19892 63692
rect 4928 63484 4968 63524
rect 5010 63484 5050 63524
rect 5092 63484 5132 63524
rect 5174 63484 5214 63524
rect 5256 63484 5296 63524
rect 20048 63484 20088 63524
rect 20130 63484 20170 63524
rect 20212 63484 20252 63524
rect 20294 63484 20334 63524
rect 20376 63484 20416 63524
rect 5548 63316 5588 63356
rect 9187 63316 9227 63356
rect 9484 63316 9524 63356
rect 12412 63316 12452 63356
rect 13564 63316 13604 63356
rect 15532 63316 15572 63356
rect 19852 63316 19892 63356
rect 8428 63232 8468 63272
rect 9868 63232 9908 63272
rect 1708 63148 1748 63188
rect 2956 63139 2996 63179
rect 3916 63148 3956 63188
rect 5164 63139 5204 63179
rect 5740 63139 5780 63179
rect 6988 63148 7028 63188
rect 8044 63148 8084 63188
rect 8299 63148 8339 63188
rect 8855 63148 8895 63188
rect 9100 63148 9140 63188
rect 9388 63148 9428 63188
rect 9571 63148 9611 63188
rect 9772 63148 9812 63188
rect 9964 63148 10004 63188
rect 10348 63148 10388 63188
rect 11596 63139 11636 63179
rect 13795 63148 13835 63188
rect 13900 63148 13940 63188
rect 14284 63148 14324 63188
rect 14860 63139 14900 63179
rect 15340 63139 15380 63179
rect 15916 63139 15956 63179
rect 17164 63148 17204 63188
rect 18094 63148 18134 63188
rect 18218 63148 18258 63188
rect 18604 63148 18644 63188
rect 19180 63139 19220 63179
rect 19660 63139 19700 63179
rect 1420 63064 1460 63104
rect 3532 63064 3572 63104
rect 7372 63064 7412 63104
rect 7756 63064 7796 63104
rect 8995 63064 9035 63104
rect 12172 63064 12212 63104
rect 12940 63064 12980 63104
rect 13324 63064 13364 63104
rect 14380 63064 14420 63104
rect 17644 63064 17684 63104
rect 18700 63064 18740 63104
rect 20140 63064 20180 63104
rect 3292 62980 3332 63020
rect 5356 62980 5396 63020
rect 8716 62980 8756 63020
rect 13180 62980 13220 63020
rect 1180 62896 1220 62936
rect 3148 62896 3188 62936
rect 7132 62896 7172 62936
rect 7516 62896 7556 62936
rect 11788 62896 11828 62936
rect 15724 62896 15764 62936
rect 17884 62896 17924 62936
rect 20380 62896 20420 62936
rect 3688 62728 3728 62768
rect 3770 62728 3810 62768
rect 3852 62728 3892 62768
rect 3934 62728 3974 62768
rect 4016 62728 4056 62768
rect 18808 62728 18848 62768
rect 18890 62728 18930 62768
rect 18972 62728 19012 62768
rect 19054 62728 19094 62768
rect 19136 62728 19176 62768
rect 9523 62560 9563 62600
rect 13516 62560 13556 62600
rect 14332 62560 14372 62600
rect 19852 62560 19892 62600
rect 3052 62392 3092 62432
rect 3916 62392 3956 62432
rect 6220 62392 6260 62432
rect 8236 62392 8276 62432
rect 10444 62392 10484 62432
rect 13708 62392 13748 62432
rect 14092 62392 14132 62432
rect 15244 62392 15284 62432
rect 20140 62392 20180 62432
rect 1228 62308 1268 62348
rect 2476 62308 2516 62348
rect 3427 62308 3467 62348
rect 3532 62308 3572 62348
rect 4012 62308 4052 62348
rect 4492 62308 4532 62348
rect 5011 62308 5051 62348
rect 5727 62308 5767 62348
rect 5836 62308 5876 62348
rect 6316 62308 6356 62348
rect 6796 62308 6836 62348
rect 7315 62308 7355 62348
rect 7747 62308 7787 62348
rect 7852 62308 7892 62348
rect 8332 62308 8372 62348
rect 8812 62308 8852 62348
rect 9331 62308 9371 62348
rect 9955 62308 9995 62348
rect 10060 62308 10100 62348
rect 10540 62308 10580 62348
rect 11020 62308 11060 62348
rect 11539 62308 11579 62348
rect 12076 62308 12116 62348
rect 13324 62308 13364 62348
rect 14755 62308 14795 62348
rect 14860 62308 14900 62348
rect 15340 62308 15380 62348
rect 15820 62308 15860 62348
rect 16308 62308 16348 62348
rect 16684 62308 16724 62348
rect 17932 62308 17972 62348
rect 18412 62308 18452 62348
rect 19660 62308 19700 62348
rect 13948 62224 13988 62264
rect 2668 62140 2708 62180
rect 2812 62140 2852 62180
rect 5164 62140 5204 62180
rect 7468 62140 7508 62180
rect 11692 62140 11732 62180
rect 16492 62140 16532 62180
rect 18124 62140 18164 62180
rect 20380 62140 20420 62180
rect 4928 61972 4968 62012
rect 5010 61972 5050 62012
rect 5092 61972 5132 62012
rect 5174 61972 5214 62012
rect 5256 61972 5296 62012
rect 20048 61972 20088 62012
rect 20130 61972 20170 62012
rect 20212 61972 20252 62012
rect 20294 61972 20334 62012
rect 20376 61972 20416 62012
rect 5308 61804 5348 61844
rect 7372 61804 7412 61844
rect 11404 61804 11444 61844
rect 11740 61804 11780 61844
rect 13612 61804 13652 61844
rect 15244 61804 15284 61844
rect 18124 61804 18164 61844
rect 20140 61804 20180 61844
rect 7516 61720 7556 61760
rect 9388 61720 9428 61760
rect 1708 61636 1748 61676
rect 2956 61627 2996 61667
rect 3406 61636 3446 61676
rect 3532 61636 3572 61676
rect 3916 61636 3956 61676
rect 4492 61627 4532 61667
rect 4972 61627 5012 61667
rect 5932 61636 5972 61676
rect 7180 61627 7220 61667
rect 7948 61636 7988 61676
rect 9196 61627 9236 61667
rect 9667 61636 9707 61676
rect 9772 61636 9812 61676
rect 10156 61636 10196 61676
rect 10732 61627 10772 61667
rect 11212 61627 11252 61667
rect 12172 61636 12212 61676
rect 13420 61627 13460 61667
rect 13804 61636 13844 61676
rect 15052 61627 15092 61667
rect 16387 61636 16427 61676
rect 16492 61636 16532 61676
rect 16876 61636 16916 61676
rect 17452 61627 17492 61667
rect 17932 61627 17972 61667
rect 18403 61636 18443 61676
rect 18508 61636 18548 61676
rect 18892 61636 18932 61676
rect 19468 61627 19508 61667
rect 19948 61627 19988 61667
rect 1420 61552 1460 61592
rect 4012 61552 4052 61592
rect 5548 61552 5588 61592
rect 7756 61552 7796 61592
rect 10252 61552 10292 61592
rect 11980 61552 12020 61592
rect 15724 61552 15764 61592
rect 16108 61552 16148 61592
rect 16972 61552 17012 61592
rect 18988 61552 19028 61592
rect 15868 61468 15908 61508
rect 1180 61384 1220 61424
rect 3148 61384 3188 61424
rect 5203 61384 5243 61424
rect 15484 61384 15524 61424
rect 3688 61216 3728 61256
rect 3770 61216 3810 61256
rect 3852 61216 3892 61256
rect 3934 61216 3974 61256
rect 4016 61216 4056 61256
rect 18808 61216 18848 61256
rect 18890 61216 18930 61256
rect 18972 61216 19012 61256
rect 19054 61216 19094 61256
rect 19136 61216 19176 61256
rect 11500 61048 11540 61088
rect 14140 61048 14180 61088
rect 16492 61048 16532 61088
rect 18124 61048 18164 61088
rect 20044 61048 20084 61088
rect 5500 60964 5540 61004
rect 12556 60964 12596 61004
rect 3052 60880 3092 60920
rect 4108 60880 4148 60920
rect 5395 60880 5435 60920
rect 5740 60880 5780 60920
rect 6124 60880 6164 60920
rect 8524 60880 8564 60920
rect 12172 60880 12212 60920
rect 14380 60880 14420 60920
rect 14668 60880 14708 60920
rect 1228 60796 1268 60836
rect 2476 60796 2516 60836
rect 3619 60796 3659 60836
rect 3724 60796 3764 60836
rect 4204 60796 4244 60836
rect 4684 60796 4724 60836
rect 5203 60796 5243 60836
rect 6316 60796 6356 60836
rect 7564 60796 7604 60836
rect 8035 60796 8075 60836
rect 8140 60796 8180 60836
rect 8620 60796 8660 60836
rect 9100 60796 9140 60836
rect 9619 60796 9659 60836
rect 10060 60796 10100 60836
rect 11308 60796 11348 60836
rect 12748 60796 12788 60836
rect 13996 60796 14036 60836
rect 15052 60796 15092 60836
rect 16300 60796 16340 60836
rect 16684 60796 16724 60836
rect 17932 60796 17972 60836
rect 18604 60796 18644 60836
rect 19852 60796 19892 60836
rect 7756 60712 7796 60752
rect 2668 60628 2708 60668
rect 2812 60628 2852 60668
rect 5884 60628 5924 60668
rect 9772 60628 9812 60668
rect 12412 60628 12452 60668
rect 14908 60628 14948 60668
rect 4928 60460 4968 60500
rect 5010 60460 5050 60500
rect 5092 60460 5132 60500
rect 5174 60460 5214 60500
rect 5256 60460 5296 60500
rect 20048 60460 20088 60500
rect 20130 60460 20170 60500
rect 20212 60460 20252 60500
rect 20294 60460 20334 60500
rect 20376 60460 20416 60500
rect 5548 60292 5588 60332
rect 7900 60292 7940 60332
rect 12604 60292 12644 60332
rect 14140 60292 14180 60332
rect 14908 60292 14948 60332
rect 15436 60292 15476 60332
rect 16012 60208 16052 60248
rect 17164 60208 17204 60248
rect 2179 60124 2219 60164
rect 2284 60124 2324 60164
rect 2668 60124 2708 60164
rect 3244 60115 3284 60155
rect 3724 60115 3764 60155
rect 4108 60124 4148 60164
rect 5356 60115 5396 60155
rect 5836 60124 5876 60164
rect 7084 60115 7124 60155
rect 9100 60124 9140 60164
rect 10348 60115 10388 60155
rect 10732 60124 10772 60164
rect 11980 60115 12020 60155
rect 15532 60124 15572 60164
rect 15769 60124 15809 60164
rect 15915 60124 15955 60164
rect 16207 60124 16247 60164
rect 16396 60124 16436 60164
rect 16780 60124 16820 60164
rect 17059 60124 17099 60164
rect 17644 60124 17684 60164
rect 17827 60124 17867 60164
rect 18700 60124 18740 60164
rect 19948 60115 19988 60155
rect 1180 60040 1220 60080
rect 1420 60040 1460 60080
rect 1804 60040 1844 60080
rect 2764 60040 2804 60080
rect 7660 60040 7700 60080
rect 12364 60040 12404 60080
rect 13036 60040 13076 60080
rect 13420 60040 13460 60080
rect 14380 60040 14420 60080
rect 14668 60040 14708 60080
rect 15052 60040 15092 60080
rect 15667 60031 15707 60071
rect 18316 60040 18356 60080
rect 12796 59956 12836 59996
rect 13996 59956 14036 59996
rect 16540 59956 16580 59996
rect 1564 59872 1604 59912
rect 3955 59872 3995 59912
rect 7276 59872 7316 59912
rect 10540 59872 10580 59912
rect 12172 59872 12212 59912
rect 13180 59872 13220 59912
rect 15292 59872 15332 59912
rect 17452 59872 17492 59912
rect 17827 59872 17867 59912
rect 18556 59872 18596 59912
rect 20140 59872 20180 59912
rect 3688 59704 3728 59744
rect 3770 59704 3810 59744
rect 3852 59704 3892 59744
rect 3934 59704 3974 59744
rect 4016 59704 4056 59744
rect 18808 59704 18848 59744
rect 18890 59704 18930 59744
rect 18972 59704 19012 59744
rect 19054 59704 19094 59744
rect 19136 59704 19176 59744
rect 3676 59536 3716 59576
rect 7804 59536 7844 59576
rect 8188 59536 8228 59576
rect 14668 59536 14708 59576
rect 16300 59452 16340 59492
rect 1420 59368 1460 59408
rect 3532 59368 3572 59408
rect 3916 59368 3956 59408
rect 6316 59368 6356 59408
rect 8044 59368 8084 59408
rect 8428 59368 8468 59408
rect 11212 59368 11252 59408
rect 12499 59368 12539 59408
rect 12844 59368 12884 59408
rect 18892 59368 18932 59408
rect 1612 59284 1652 59324
rect 2860 59284 2900 59324
rect 4108 59284 4148 59324
rect 5356 59284 5396 59324
rect 5827 59284 5867 59324
rect 5932 59284 5972 59324
rect 6412 59284 6452 59324
rect 6892 59284 6932 59324
rect 7380 59284 7420 59324
rect 9004 59284 9044 59324
rect 10252 59284 10292 59324
rect 10723 59284 10763 59324
rect 10828 59284 10868 59324
rect 11308 59284 11348 59324
rect 11791 59284 11831 59324
rect 12307 59284 12347 59324
rect 13228 59284 13268 59324
rect 14476 59284 14516 59324
rect 14860 59284 14900 59324
rect 16108 59284 16148 59324
rect 16684 59284 16724 59324
rect 17932 59284 17972 59324
rect 18403 59284 18443 59324
rect 18508 59284 18548 59324
rect 18988 59284 19028 59324
rect 19468 59284 19508 59324
rect 19987 59284 20027 59324
rect 3052 59200 3092 59240
rect 5548 59200 5588 59240
rect 18124 59200 18164 59240
rect 1180 59116 1220 59156
rect 3292 59116 3332 59156
rect 7564 59116 7604 59156
rect 8812 59116 8852 59156
rect 12604 59116 12644 59156
rect 16300 59116 16340 59156
rect 20140 59116 20180 59156
rect 4928 58948 4968 58988
rect 5010 58948 5050 58988
rect 5092 58948 5132 58988
rect 5174 58948 5214 58988
rect 5256 58948 5296 58988
rect 20048 58948 20088 58988
rect 20130 58948 20170 58988
rect 20212 58948 20252 58988
rect 20294 58948 20334 58988
rect 20376 58948 20416 58988
rect 4012 58780 4052 58820
rect 5788 58780 5828 58820
rect 8236 58780 8276 58820
rect 10723 58780 10763 58820
rect 12988 58780 13028 58820
rect 15052 58780 15092 58820
rect 17164 58780 17204 58820
rect 17932 58780 17972 58820
rect 8419 58696 8459 58736
rect 11260 58696 11300 58736
rect 17342 58696 17382 58736
rect 2275 58612 2315 58652
rect 2380 58612 2420 58652
rect 2764 58612 2804 58652
rect 3340 58603 3380 58643
rect 3820 58603 3860 58643
rect 4204 58612 4244 58652
rect 5452 58603 5492 58643
rect 6796 58612 6836 58652
rect 8044 58603 8084 58643
rect 8611 58612 8651 58652
rect 9100 58603 9140 58643
rect 9580 58612 9620 58652
rect 10060 58612 10100 58652
rect 10173 58632 10213 58672
rect 10564 58612 10604 58652
rect 10723 58612 10763 58652
rect 10867 58612 10907 58652
rect 11011 58601 11051 58641
rect 11113 58612 11153 58652
rect 11404 58612 11444 58652
rect 13612 58612 13652 58652
rect 14860 58603 14900 58643
rect 15427 58612 15467 58652
rect 15532 58612 15572 58652
rect 15916 58612 15956 58652
rect 16492 58603 16532 58643
rect 16972 58603 17012 58643
rect 17548 58612 17588 58652
rect 17644 58603 17684 58643
rect 17836 58612 17876 58652
rect 18028 58612 18068 58652
rect 18700 58612 18740 58652
rect 19948 58603 19988 58643
rect 1420 58528 1460 58568
rect 1804 58528 1844 58568
rect 2860 58528 2900 58568
rect 6028 58528 6068 58568
rect 6412 58528 6452 58568
rect 9676 58528 9716 58568
rect 11788 58528 11828 58568
rect 12748 58528 12788 58568
rect 13132 58528 13172 58568
rect 16012 58528 16052 58568
rect 18412 58528 18452 58568
rect 6172 58444 6212 58484
rect 1180 58360 1220 58400
rect 1564 58360 1604 58400
rect 5644 58360 5684 58400
rect 12028 58360 12068 58400
rect 13372 58360 13412 58400
rect 17347 58360 17387 58400
rect 18172 58360 18212 58400
rect 20140 58360 20180 58400
rect 3688 58192 3728 58232
rect 3770 58192 3810 58232
rect 3852 58192 3892 58232
rect 3934 58192 3974 58232
rect 4016 58192 4056 58232
rect 18808 58192 18848 58232
rect 18890 58192 18930 58232
rect 18972 58192 19012 58232
rect 19054 58192 19094 58232
rect 19136 58192 19176 58232
rect 5299 58024 5339 58064
rect 11308 58024 11348 58064
rect 11500 58024 11540 58064
rect 14332 58024 14372 58064
rect 15004 58024 15044 58064
rect 15388 58024 15428 58064
rect 14908 57940 14948 57980
rect 4012 57856 4052 57896
rect 7084 57856 7124 57896
rect 14092 57856 14132 57896
rect 1516 57772 1556 57812
rect 2764 57772 2804 57812
rect 3523 57772 3563 57812
rect 3628 57772 3668 57812
rect 4108 57772 4148 57812
rect 4588 57772 4628 57812
rect 5068 57805 5108 57845
rect 14668 57856 14708 57896
rect 15244 57856 15284 57896
rect 15628 57856 15668 57896
rect 15820 57856 15860 57896
rect 16051 57847 16091 57887
rect 18796 57856 18836 57896
rect 5636 57772 5676 57812
rect 6892 57772 6932 57812
rect 7468 57772 7508 57812
rect 8716 57772 8756 57812
rect 9868 57772 9908 57812
rect 11116 57772 11156 57812
rect 11500 57772 11540 57812
rect 11615 57772 11655 57812
rect 11788 57772 11828 57812
rect 11980 57772 12020 57812
rect 12119 57805 12159 57845
rect 12460 57772 12500 57812
rect 13708 57772 13748 57812
rect 15916 57772 15956 57812
rect 16153 57772 16193 57812
rect 16588 57772 16628 57812
rect 17836 57772 17876 57812
rect 18307 57772 18347 57812
rect 18412 57772 18452 57812
rect 18892 57772 18932 57812
rect 19372 57772 19412 57812
rect 19891 57772 19931 57812
rect 2956 57688 2996 57728
rect 18028 57688 18068 57728
rect 5452 57604 5492 57644
rect 7324 57604 7364 57644
rect 8908 57604 8948 57644
rect 11308 57604 11348 57644
rect 12268 57604 12308 57644
rect 13900 57604 13940 57644
rect 20044 57604 20084 57644
rect 4928 57436 4968 57476
rect 5010 57436 5050 57476
rect 5092 57436 5132 57476
rect 5174 57436 5214 57476
rect 5256 57436 5296 57476
rect 20048 57436 20088 57476
rect 20130 57436 20170 57476
rect 20212 57436 20252 57476
rect 20294 57436 20334 57476
rect 20376 57436 20416 57476
rect 2236 57268 2276 57308
rect 6748 57268 6788 57308
rect 11308 57268 11348 57308
rect 14956 57268 14996 57308
rect 4204 57184 4244 57224
rect 12940 57184 12980 57224
rect 2764 57100 2804 57140
rect 4012 57091 4052 57131
rect 4867 57100 4907 57140
rect 4972 57100 5012 57140
rect 5356 57100 5396 57140
rect 5932 57091 5972 57131
rect 6412 57091 6452 57131
rect 7747 57100 7787 57140
rect 7852 57100 7892 57140
rect 8236 57100 8276 57140
rect 8812 57091 8852 57131
rect 9292 57091 9332 57131
rect 9868 57100 9908 57140
rect 11116 57091 11156 57131
rect 11500 57100 11540 57140
rect 12748 57091 12788 57131
rect 13219 57100 13259 57140
rect 13324 57100 13364 57140
rect 13708 57100 13748 57140
rect 14284 57091 14324 57131
rect 14764 57091 14804 57131
rect 15340 57100 15380 57140
rect 16588 57091 16628 57131
rect 16972 57100 17012 57140
rect 18220 57091 18260 57131
rect 18604 57100 18644 57140
rect 19852 57091 19892 57131
rect 1420 57016 1460 57056
rect 1804 57016 1844 57056
rect 1996 57016 2036 57056
rect 2572 57016 2612 57056
rect 4588 57016 4628 57056
rect 5452 57016 5492 57056
rect 6643 57016 6683 57056
rect 6988 57016 7028 57056
rect 8332 57016 8372 57056
rect 13804 57016 13844 57056
rect 1180 56848 1220 56888
rect 1564 56848 1604 56888
rect 2332 56848 2372 56888
rect 4348 56848 4388 56888
rect 9523 56848 9563 56888
rect 16780 56848 16820 56888
rect 18412 56848 18452 56888
rect 20044 56848 20084 56888
rect 3688 56680 3728 56720
rect 3770 56680 3810 56720
rect 3852 56680 3892 56720
rect 3934 56680 3974 56720
rect 4016 56680 4056 56720
rect 18808 56680 18848 56720
rect 18890 56680 18930 56720
rect 18972 56680 19012 56720
rect 19054 56680 19094 56720
rect 19136 56680 19176 56720
rect 8044 56512 8084 56552
rect 10108 56512 10148 56552
rect 13036 56512 13076 56552
rect 17980 56512 18020 56552
rect 5404 56428 5444 56468
rect 17308 56428 17348 56468
rect 1420 56344 1460 56384
rect 4012 56344 4052 56384
rect 5299 56344 5339 56384
rect 5644 56344 5684 56384
rect 6412 56344 6452 56384
rect 10348 56344 10388 56384
rect 13804 56344 13844 56384
rect 15820 56344 15860 56384
rect 17548 56344 17588 56384
rect 17740 56344 17780 56384
rect 18700 56344 18740 56384
rect 20140 56344 20180 56384
rect 1708 56260 1748 56300
rect 2956 56260 2996 56300
rect 3523 56260 3563 56300
rect 3628 56260 3668 56300
rect 4108 56260 4148 56300
rect 4588 56260 4628 56300
rect 5107 56260 5147 56300
rect 6609 56260 6649 56300
rect 7852 56260 7892 56300
rect 8524 56260 8564 56300
rect 9772 56260 9812 56300
rect 11596 56260 11636 56300
rect 12844 56260 12884 56300
rect 13315 56260 13355 56300
rect 13420 56260 13460 56300
rect 13900 56260 13940 56300
rect 14380 56260 14420 56300
rect 14868 56260 14908 56300
rect 15331 56260 15371 56300
rect 15436 56260 15476 56300
rect 15916 56260 15956 56300
rect 16396 56260 16436 56300
rect 16884 56260 16924 56300
rect 18211 56260 18251 56300
rect 18316 56260 18356 56300
rect 18796 56260 18836 56300
rect 19276 56260 19316 56300
rect 19756 56293 19796 56333
rect 1180 56176 1220 56216
rect 3148 56176 3188 56216
rect 20380 56176 20420 56216
rect 6172 56092 6212 56132
rect 9964 56092 10004 56132
rect 15052 56092 15092 56132
rect 17068 56092 17108 56132
rect 19948 56092 19988 56132
rect 4928 55924 4968 55964
rect 5010 55924 5050 55964
rect 5092 55924 5132 55964
rect 5174 55924 5214 55964
rect 5256 55924 5296 55964
rect 20048 55924 20088 55964
rect 20130 55924 20170 55964
rect 20212 55924 20252 55964
rect 20294 55924 20334 55964
rect 20376 55924 20416 55964
rect 3292 55756 3332 55796
rect 5356 55756 5396 55796
rect 5500 55756 5540 55796
rect 17068 55756 17108 55796
rect 17212 55756 17252 55796
rect 2860 55672 2900 55712
rect 8044 55672 8084 55712
rect 15052 55672 15092 55712
rect 1420 55588 1460 55628
rect 2668 55579 2708 55619
rect 3916 55588 3956 55628
rect 5164 55579 5204 55619
rect 6604 55588 6644 55628
rect 7852 55579 7892 55619
rect 8419 55588 8459 55628
rect 8524 55588 8564 55628
rect 8908 55588 8948 55628
rect 9484 55579 9524 55619
rect 9964 55579 10004 55619
rect 10828 55579 10868 55619
rect 12076 55588 12116 55628
rect 13612 55588 13652 55628
rect 14860 55579 14900 55619
rect 15331 55588 15371 55628
rect 15436 55588 15476 55628
rect 15820 55588 15860 55628
rect 16396 55579 16436 55619
rect 16876 55579 16916 55619
rect 18028 55588 18068 55628
rect 19276 55579 19316 55619
rect 3052 55504 3092 55544
rect 3628 55504 3668 55544
rect 5740 55504 5780 55544
rect 5932 55504 5972 55544
rect 9004 55504 9044 55544
rect 12268 55504 12308 55544
rect 15916 55504 15956 55544
rect 17452 55504 17492 55544
rect 17644 55504 17684 55544
rect 19756 55504 19796 55544
rect 20140 55504 20180 55544
rect 3388 55420 3428 55460
rect 19996 55420 20036 55460
rect 6172 55336 6212 55376
rect 10195 55336 10235 55376
rect 10636 55336 10676 55376
rect 12508 55336 12548 55376
rect 17884 55336 17924 55376
rect 19468 55336 19508 55376
rect 20380 55336 20420 55376
rect 3688 55168 3728 55208
rect 3770 55168 3810 55208
rect 3852 55168 3892 55208
rect 3934 55168 3974 55208
rect 4016 55168 4056 55208
rect 18808 55168 18848 55208
rect 18890 55168 18930 55208
rect 18972 55168 19012 55208
rect 19054 55168 19094 55208
rect 19136 55168 19176 55208
rect 13420 55000 13460 55040
rect 15052 55000 15092 55040
rect 16780 55000 16820 55040
rect 20332 54916 20372 54956
rect 10060 54832 10100 54872
rect 11347 54832 11387 54872
rect 1420 54748 1460 54788
rect 2668 54748 2708 54788
rect 3052 54748 3092 54788
rect 3191 54748 3231 54788
rect 3532 54748 3572 54788
rect 3715 54748 3755 54788
rect 3820 54748 3860 54788
rect 4012 54748 4052 54788
rect 4300 54748 4340 54788
rect 5548 54748 5588 54788
rect 6220 54748 6260 54788
rect 7468 54748 7508 54788
rect 7852 54748 7892 54788
rect 9100 54748 9140 54788
rect 9571 54748 9611 54788
rect 9676 54748 9716 54788
rect 10156 54748 10196 54788
rect 10636 54748 10676 54788
rect 11155 54748 11195 54788
rect 11980 54748 12020 54788
rect 13228 54748 13268 54788
rect 13612 54748 13652 54788
rect 14860 54748 14900 54788
rect 15340 54748 15380 54788
rect 16588 54748 16628 54788
rect 17068 54748 17108 54788
rect 18316 54748 18356 54788
rect 18892 54748 18932 54788
rect 20140 54748 20180 54788
rect 3619 54664 3659 54704
rect 2860 54580 2900 54620
rect 3340 54580 3380 54620
rect 4156 54580 4196 54620
rect 5740 54580 5780 54620
rect 7660 54580 7700 54620
rect 9292 54580 9332 54620
rect 18508 54580 18548 54620
rect 4928 54412 4968 54452
rect 5010 54412 5050 54452
rect 5092 54412 5132 54452
rect 5174 54412 5214 54452
rect 5256 54412 5296 54452
rect 20048 54412 20088 54452
rect 20130 54412 20170 54452
rect 20212 54412 20252 54452
rect 20294 54412 20334 54452
rect 20376 54412 20416 54452
rect 1948 54244 1988 54284
rect 7948 54244 7988 54284
rect 11308 54244 11348 54284
rect 12892 54244 12932 54284
rect 17020 54244 17060 54284
rect 17692 54244 17732 54284
rect 20044 54244 20084 54284
rect 4003 54151 4043 54191
rect 14860 54160 14900 54200
rect 17788 54160 17828 54200
rect 2092 54076 2132 54116
rect 3340 54067 3380 54107
rect 3699 54065 3739 54105
rect 3820 54067 3860 54107
rect 4099 54076 4139 54116
rect 4233 54076 4273 54116
rect 4492 54076 4532 54116
rect 5740 54067 5780 54107
rect 6211 54076 6251 54116
rect 6316 54076 6356 54116
rect 6700 54076 6740 54116
rect 7276 54067 7316 54107
rect 7756 54067 7796 54107
rect 9379 54076 9419 54116
rect 9489 54076 9529 54116
rect 9868 54076 9908 54116
rect 10444 54067 10484 54107
rect 10924 54067 10964 54107
rect 11500 54067 11540 54107
rect 12748 54076 12788 54116
rect 13420 54076 13460 54116
rect 14668 54067 14708 54107
rect 15139 54076 15179 54116
rect 15244 54076 15284 54116
rect 15628 54076 15668 54116
rect 16204 54067 16244 54107
rect 16684 54067 16724 54107
rect 18307 54076 18347 54116
rect 18412 54076 18452 54116
rect 18796 54076 18836 54116
rect 19372 54067 19412 54107
rect 19852 54067 19892 54107
rect 1420 53992 1460 54032
rect 1708 53992 1748 54032
rect 6796 53992 6836 54032
rect 9964 53992 10004 54032
rect 13132 53992 13172 54032
rect 15724 53992 15764 54032
rect 16915 53992 16955 54032
rect 17260 53992 17300 54032
rect 17452 53992 17492 54032
rect 18028 53992 18068 54032
rect 18892 53992 18932 54032
rect 3532 53908 3572 53948
rect 1180 53824 1220 53864
rect 3715 53824 3755 53864
rect 5932 53824 5972 53864
rect 11155 53824 11195 53864
rect 3688 53656 3728 53696
rect 3770 53656 3810 53696
rect 3852 53656 3892 53696
rect 3934 53656 3974 53696
rect 4016 53656 4056 53696
rect 18808 53656 18848 53696
rect 18890 53656 18930 53696
rect 18972 53656 19012 53696
rect 19054 53656 19094 53696
rect 19136 53656 19176 53696
rect 2140 53488 2180 53528
rect 8467 53488 8507 53528
rect 10492 53488 10532 53528
rect 12412 53488 12452 53528
rect 15244 53488 15284 53528
rect 17788 53488 17828 53528
rect 10060 53404 10100 53444
rect 12508 53404 12548 53444
rect 17308 53404 17348 53444
rect 1180 53320 1220 53360
rect 1420 53320 1460 53360
rect 1900 53320 1940 53360
rect 3148 53320 3188 53360
rect 7180 53320 7220 53360
rect 10252 53320 10292 53360
rect 10588 53320 10628 53360
rect 12172 53320 12212 53360
rect 12748 53320 12788 53360
rect 16012 53320 16052 53360
rect 17404 53320 17444 53360
rect 17644 53320 17684 53360
rect 18028 53320 18068 53360
rect 18988 53320 19028 53360
rect 2659 53236 2699 53276
rect 2764 53236 2804 53276
rect 3244 53236 3284 53276
rect 3724 53236 3764 53276
rect 4212 53236 4252 53276
rect 4876 53236 4916 53276
rect 6124 53236 6164 53276
rect 6670 53236 6710 53276
rect 6796 53236 6836 53276
rect 7276 53236 7316 53276
rect 7756 53236 7796 53276
rect 8244 53236 8284 53276
rect 8716 53236 8756 53276
rect 9004 53236 9044 53276
rect 9388 53236 9428 53276
rect 9643 53236 9683 53276
rect 9763 53236 9803 53276
rect 10732 53236 10772 53276
rect 13804 53236 13844 53276
rect 15052 53236 15092 53276
rect 15523 53236 15563 53276
rect 15628 53236 15668 53276
rect 16108 53236 16148 53276
rect 16588 53236 16628 53276
rect 17107 53236 17147 53276
rect 18499 53236 18539 53276
rect 18604 53236 18644 53276
rect 19084 53236 19124 53276
rect 19564 53236 19604 53276
rect 20052 53236 20092 53276
rect 4396 53068 4436 53108
rect 6316 53068 6356 53108
rect 8803 53068 8843 53108
rect 20236 53068 20276 53108
rect 4928 52900 4968 52940
rect 5010 52900 5050 52940
rect 5092 52900 5132 52940
rect 5174 52900 5214 52940
rect 5256 52900 5296 52940
rect 20048 52900 20088 52940
rect 20130 52900 20170 52940
rect 20212 52900 20252 52940
rect 20294 52900 20334 52940
rect 20376 52900 20416 52940
rect 2668 52732 2708 52772
rect 9868 52732 9908 52772
rect 10636 52732 10676 52772
rect 10924 52732 10964 52772
rect 12556 52732 12596 52772
rect 15628 52732 15668 52772
rect 17260 52732 17300 52772
rect 18892 52732 18932 52772
rect 19036 52732 19076 52772
rect 5068 52648 5108 52688
rect 19420 52648 19460 52688
rect 1228 52564 1268 52604
rect 2476 52555 2516 52595
rect 3628 52564 3668 52604
rect 4876 52555 4916 52595
rect 5347 52564 5387 52604
rect 5452 52564 5492 52604
rect 5836 52564 5876 52604
rect 6412 52555 6452 52595
rect 6892 52555 6932 52595
rect 8131 52564 8171 52604
rect 8236 52564 8276 52604
rect 8620 52564 8660 52604
rect 9196 52555 9236 52595
rect 9676 52555 9716 52595
rect 10007 52564 10047 52604
rect 10252 52564 10292 52604
rect 10540 52564 10580 52604
rect 10723 52564 10763 52604
rect 11116 52555 11156 52595
rect 12364 52564 12404 52604
rect 12748 52555 12788 52595
rect 13996 52564 14036 52604
rect 14188 52564 14228 52604
rect 15436 52555 15476 52595
rect 15820 52564 15860 52604
rect 17068 52555 17108 52595
rect 17452 52564 17492 52604
rect 18700 52555 18740 52595
rect 3052 52480 3092 52520
rect 5932 52480 5972 52520
rect 8716 52480 8756 52520
rect 10147 52480 10187 52520
rect 10348 52480 10388 52520
rect 19276 52480 19316 52520
rect 19660 52480 19700 52520
rect 20140 52480 20180 52520
rect 2812 52312 2852 52352
rect 7123 52312 7163 52352
rect 20380 52312 20420 52352
rect 3688 52144 3728 52184
rect 3770 52144 3810 52184
rect 3852 52144 3892 52184
rect 3934 52144 3974 52184
rect 4016 52144 4056 52184
rect 18808 52144 18848 52184
rect 18890 52144 18930 52184
rect 18972 52144 19012 52184
rect 19054 52144 19094 52184
rect 19136 52144 19176 52184
rect 7852 51976 7892 52016
rect 10348 51976 10388 52016
rect 10540 51976 10580 52016
rect 10924 51976 10964 52016
rect 1420 51808 1460 51848
rect 1804 51808 1844 51848
rect 2092 51808 2132 51848
rect 2476 51808 2516 51848
rect 2716 51808 2756 51848
rect 4012 51808 4052 51848
rect 5068 51808 5108 51848
rect 6412 51808 6452 51848
rect 9868 51808 9908 51848
rect 12556 51808 12596 51848
rect 20140 51808 20180 51848
rect 3043 51724 3083 51764
rect 3532 51724 3572 51764
rect 4108 51724 4148 51764
rect 4492 51724 4532 51764
rect 4610 51724 4650 51764
rect 5923 51724 5963 51764
rect 6028 51724 6068 51764
rect 6508 51724 6548 51764
rect 6988 51724 7028 51764
rect 7480 51724 7520 51764
rect 8044 51724 8084 51764
rect 9292 51724 9332 51764
rect 9527 51724 9567 51764
rect 9667 51724 9707 51764
rect 9772 51724 9812 51764
rect 10051 51724 10091 51764
rect 10359 51724 10399 51764
rect 10540 51724 10580 51764
rect 10729 51724 10769 51764
rect 11116 51724 11156 51764
rect 12364 51724 12404 51764
rect 13420 51724 13460 51764
rect 14668 51724 14708 51764
rect 14860 51724 14900 51764
rect 16108 51724 16148 51764
rect 16684 51724 16724 51764
rect 17932 51724 17972 51764
rect 18220 51724 18260 51764
rect 19468 51724 19508 51764
rect 2332 51640 2372 51680
rect 4828 51640 4868 51680
rect 10156 51640 10196 51680
rect 10924 51640 10964 51680
rect 12796 51640 12836 51680
rect 1180 51556 1220 51596
rect 1564 51556 1604 51596
rect 2860 51556 2900 51596
rect 7660 51556 7700 51596
rect 13228 51556 13268 51596
rect 16300 51556 16340 51596
rect 16492 51556 16532 51596
rect 19660 51556 19700 51596
rect 20380 51556 20420 51596
rect 4928 51388 4968 51428
rect 5010 51388 5050 51428
rect 5092 51388 5132 51428
rect 5174 51388 5214 51428
rect 5256 51388 5296 51428
rect 20048 51388 20088 51428
rect 20130 51388 20170 51428
rect 20212 51388 20252 51428
rect 20294 51388 20334 51428
rect 20376 51388 20416 51428
rect 1180 51220 1220 51260
rect 1564 51220 1604 51260
rect 5932 51220 5972 51260
rect 7564 51220 7604 51260
rect 12124 51220 12164 51260
rect 17452 51220 17492 51260
rect 19612 51220 19652 51260
rect 13324 51136 13364 51176
rect 4492 51052 4532 51092
rect 5740 51043 5780 51083
rect 6124 51052 6164 51092
rect 7372 51043 7412 51083
rect 8908 51052 8948 51092
rect 10156 51043 10196 51083
rect 10540 51052 10580 51092
rect 11788 51043 11828 51083
rect 13516 51043 13556 51083
rect 14764 51052 14804 51092
rect 15715 51052 15755 51092
rect 15820 51052 15860 51092
rect 16204 51052 16244 51092
rect 16780 51043 16820 51083
rect 17260 51043 17300 51083
rect 17644 51052 17684 51092
rect 18892 51043 18932 51083
rect 1420 50968 1460 51008
rect 1804 50968 1844 51008
rect 2764 50968 2804 51008
rect 12364 50968 12404 51008
rect 16300 50968 16340 51008
rect 19372 50968 19412 51008
rect 19756 50968 19796 51008
rect 20140 50968 20180 51008
rect 19996 50884 20036 50924
rect 2524 50800 2564 50840
rect 10348 50800 10388 50840
rect 11980 50800 12020 50840
rect 19084 50800 19124 50840
rect 20380 50800 20420 50840
rect 3688 50632 3728 50672
rect 3770 50632 3810 50672
rect 3852 50632 3892 50672
rect 3934 50632 3974 50672
rect 4016 50632 4056 50672
rect 18808 50632 18848 50672
rect 18890 50632 18930 50672
rect 18972 50632 19012 50672
rect 19054 50632 19094 50672
rect 19136 50632 19176 50672
rect 8908 50380 8948 50420
rect 11932 50380 11972 50420
rect 18460 50380 18500 50420
rect 9676 50296 9716 50336
rect 11404 50296 11444 50336
rect 11692 50296 11732 50336
rect 12268 50296 12308 50336
rect 16396 50296 16436 50336
rect 19660 50296 19700 50336
rect 2092 50212 2132 50252
rect 3340 50212 3380 50252
rect 4012 50212 4052 50252
rect 5260 50212 5300 50252
rect 7468 50212 7508 50252
rect 8716 50212 8756 50252
rect 9187 50212 9227 50252
rect 9292 50212 9332 50252
rect 9772 50212 9812 50252
rect 10252 50212 10292 50252
rect 10740 50212 10780 50252
rect 12556 50212 12596 50252
rect 13804 50212 13844 50252
rect 14188 50212 14228 50252
rect 15436 50212 15476 50252
rect 15907 50212 15947 50252
rect 16012 50212 16052 50252
rect 16492 50212 16532 50252
rect 16972 50212 17012 50252
rect 17460 50212 17500 50252
rect 18691 50212 18731 50252
rect 19180 50212 19220 50252
rect 19756 50212 19796 50252
rect 20140 50212 20180 50252
rect 20241 50212 20281 50252
rect 3532 50044 3572 50084
rect 5452 50044 5492 50084
rect 10924 50044 10964 50084
rect 11164 50044 11204 50084
rect 12028 50044 12068 50084
rect 13996 50044 14036 50084
rect 15628 50044 15668 50084
rect 17644 50044 17684 50084
rect 4928 49876 4968 49916
rect 5010 49876 5050 49916
rect 5092 49876 5132 49916
rect 5174 49876 5214 49916
rect 5256 49876 5296 49916
rect 20048 49876 20088 49916
rect 20130 49876 20170 49916
rect 20212 49876 20252 49916
rect 20294 49876 20334 49916
rect 20376 49876 20416 49916
rect 9196 49708 9236 49748
rect 11404 49708 11444 49748
rect 15820 49708 15860 49748
rect 17452 49708 17492 49748
rect 20380 49708 20420 49748
rect 11836 49624 11876 49664
rect 1996 49540 2036 49580
rect 3244 49531 3284 49571
rect 4204 49531 4244 49571
rect 5452 49540 5492 49580
rect 6316 49531 6356 49571
rect 7564 49540 7604 49580
rect 7756 49540 7796 49580
rect 9004 49531 9044 49571
rect 9667 49540 9707 49580
rect 9772 49540 9812 49580
rect 10156 49540 10196 49580
rect 10732 49531 10772 49571
rect 11212 49531 11252 49571
rect 11980 49540 12020 49580
rect 13228 49531 13268 49571
rect 14380 49540 14420 49580
rect 15628 49531 15668 49571
rect 16012 49540 16052 49580
rect 17260 49531 17300 49571
rect 10252 49456 10292 49496
rect 11596 49456 11636 49496
rect 17836 49456 17876 49496
rect 19372 49456 19412 49496
rect 19756 49456 19796 49496
rect 20140 49456 20180 49496
rect 3436 49372 3476 49412
rect 19996 49372 20036 49412
rect 4012 49288 4052 49328
rect 6124 49288 6164 49328
rect 13420 49288 13460 49328
rect 17596 49288 17636 49328
rect 19612 49288 19652 49328
rect 3688 49120 3728 49160
rect 3770 49120 3810 49160
rect 3852 49120 3892 49160
rect 3934 49120 3974 49160
rect 4016 49120 4056 49160
rect 18808 49120 18848 49160
rect 18890 49120 18930 49160
rect 18972 49120 19012 49160
rect 19054 49120 19094 49160
rect 19136 49120 19176 49160
rect 11404 48952 11444 48992
rect 4540 48868 4580 48908
rect 6988 48868 7028 48908
rect 8572 48868 8612 48908
rect 14716 48868 14756 48908
rect 3820 48784 3860 48824
rect 4780 48784 4820 48824
rect 5548 48784 5588 48824
rect 8812 48784 8852 48824
rect 8956 48784 8996 48824
rect 9196 48784 9236 48824
rect 9676 48784 9716 48824
rect 12172 48784 12212 48824
rect 14956 48784 14996 48824
rect 16300 48784 16340 48824
rect 18604 48784 18644 48824
rect 19996 48784 20036 48824
rect 20236 48784 20276 48824
rect 5059 48700 5099 48740
rect 5164 48700 5204 48740
rect 5644 48700 5684 48740
rect 6124 48700 6164 48740
rect 6612 48700 6652 48740
rect 7180 48700 7220 48740
rect 8428 48700 8468 48740
rect 9964 48700 10004 48740
rect 11212 48700 11252 48740
rect 11683 48700 11723 48740
rect 11788 48700 11828 48740
rect 12268 48700 12308 48740
rect 12748 48700 12788 48740
rect 13267 48700 13307 48740
rect 15331 48700 15371 48740
rect 15820 48700 15860 48740
rect 16396 48700 16436 48740
rect 16780 48700 16820 48740
rect 16893 48719 16933 48759
rect 18115 48700 18155 48740
rect 18220 48700 18260 48740
rect 18700 48700 18740 48740
rect 19180 48700 19220 48740
rect 19668 48700 19708 48740
rect 4060 48532 4100 48572
rect 6796 48532 6836 48572
rect 9436 48532 9476 48572
rect 13420 48532 13460 48572
rect 15148 48532 15188 48572
rect 19852 48532 19892 48572
rect 4928 48364 4968 48404
rect 5010 48364 5050 48404
rect 5092 48364 5132 48404
rect 5174 48364 5214 48404
rect 5256 48364 5296 48404
rect 20048 48364 20088 48404
rect 20130 48364 20170 48404
rect 20212 48364 20252 48404
rect 20294 48364 20334 48404
rect 20376 48364 20416 48404
rect 3916 48196 3956 48236
rect 5932 48196 5972 48236
rect 17452 48196 17492 48236
rect 19084 48196 19124 48236
rect 20380 48196 20420 48236
rect 2179 48028 2219 48068
rect 2284 48028 2324 48068
rect 2668 48028 2708 48068
rect 3244 48019 3284 48059
rect 3724 48019 3764 48059
rect 4174 48028 4214 48068
rect 4298 48028 4338 48068
rect 4684 48028 4724 48068
rect 5260 48019 5300 48059
rect 5740 48019 5780 48059
rect 12940 48028 12980 48068
rect 14188 48019 14228 48059
rect 15715 48028 15755 48068
rect 15820 48028 15860 48068
rect 16204 48028 16244 48068
rect 16780 48019 16820 48059
rect 17260 48019 17300 48059
rect 17644 48028 17684 48068
rect 18892 48019 18932 48059
rect 2764 47944 2804 47984
rect 4780 47944 4820 47984
rect 7948 47944 7988 47984
rect 9292 47944 9332 47984
rect 9676 47944 9716 47984
rect 10348 47944 10388 47984
rect 10924 47944 10964 47984
rect 16300 47944 16340 47984
rect 19756 47944 19796 47984
rect 20140 47944 20180 47984
rect 10588 47860 10628 47900
rect 19996 47860 20036 47900
rect 8188 47776 8228 47816
rect 9052 47776 9092 47816
rect 9916 47776 9956 47816
rect 10684 47776 10724 47816
rect 14380 47776 14420 47816
rect 3688 47608 3728 47648
rect 3770 47608 3810 47648
rect 3852 47608 3892 47648
rect 3934 47608 3974 47648
rect 4016 47608 4056 47648
rect 18808 47608 18848 47648
rect 18890 47608 18930 47648
rect 18972 47608 19012 47648
rect 19054 47608 19094 47648
rect 19136 47608 19176 47648
rect 3052 47440 3092 47480
rect 9811 47440 9851 47480
rect 15820 47440 15860 47480
rect 17452 47440 17492 47480
rect 19468 47440 19508 47480
rect 3820 47272 3860 47312
rect 8524 47272 8564 47312
rect 19756 47272 19796 47312
rect 20140 47272 20180 47312
rect 20380 47272 20420 47312
rect 1612 47188 1652 47228
rect 2860 47188 2900 47228
rect 3331 47188 3371 47228
rect 3436 47188 3476 47228
rect 3916 47188 3956 47228
rect 4396 47188 4436 47228
rect 4884 47188 4924 47228
rect 6124 47188 6164 47228
rect 6316 47188 6356 47228
rect 7564 47188 7604 47228
rect 8035 47188 8075 47228
rect 8140 47188 8180 47228
rect 8620 47188 8660 47228
rect 9100 47188 9140 47228
rect 9588 47188 9628 47228
rect 10444 47188 10484 47228
rect 10828 47188 10868 47228
rect 12076 47188 12116 47228
rect 12748 47188 12788 47228
rect 13996 47188 14036 47228
rect 14380 47188 14420 47228
rect 15628 47188 15668 47228
rect 16012 47188 16052 47228
rect 17260 47188 17300 47228
rect 18028 47188 18068 47228
rect 19276 47188 19316 47228
rect 7756 47104 7796 47144
rect 5068 47020 5108 47060
rect 5980 47020 6020 47060
rect 10588 47020 10628 47060
rect 12268 47020 12308 47060
rect 14188 47020 14228 47060
rect 19996 47020 20036 47060
rect 4928 46852 4968 46892
rect 5010 46852 5050 46892
rect 5092 46852 5132 46892
rect 5174 46852 5214 46892
rect 5256 46852 5296 46892
rect 20048 46852 20088 46892
rect 20130 46852 20170 46892
rect 20212 46852 20252 46892
rect 20294 46852 20334 46892
rect 20376 46852 20416 46892
rect 2764 46684 2804 46724
rect 3868 46684 3908 46724
rect 4348 46684 4388 46724
rect 5356 46684 5396 46724
rect 9388 46684 9428 46724
rect 10348 46684 10388 46724
rect 15148 46684 15188 46724
rect 1324 46516 1364 46556
rect 2572 46507 2612 46547
rect 4963 46516 5003 46556
rect 5548 46507 5588 46547
rect 6756 46516 6796 46556
rect 6988 46516 7028 46556
rect 7180 46516 7220 46556
rect 7324 46516 7364 46556
rect 7468 46516 7508 46556
rect 7948 46516 7988 46556
rect 9196 46507 9236 46547
rect 9580 46516 9620 46556
rect 9763 46516 9803 46556
rect 9868 46516 9908 46556
rect 10060 46516 10100 46556
rect 10202 46516 10242 46556
rect 10627 46516 10667 46556
rect 10732 46516 10772 46556
rect 11116 46516 11156 46556
rect 11692 46507 11732 46547
rect 12172 46507 12212 46547
rect 13411 46516 13451 46556
rect 13516 46516 13556 46556
rect 13900 46516 13940 46556
rect 14476 46507 14516 46547
rect 14956 46507 14996 46547
rect 15532 46507 15572 46547
rect 16780 46516 16820 46556
rect 17836 46516 17876 46556
rect 19084 46507 19124 46547
rect 3628 46432 3668 46472
rect 4108 46432 4148 46472
rect 4492 46432 4532 46472
rect 11212 46432 11252 46472
rect 12403 46432 12443 46472
rect 12748 46432 12788 46472
rect 13996 46432 14036 46472
rect 19756 46432 19796 46472
rect 20140 46432 20180 46472
rect 4935 46348 4975 46388
rect 5155 46348 5195 46388
rect 19996 46348 20036 46388
rect 4732 46264 4772 46304
rect 7084 46264 7124 46304
rect 9868 46264 9908 46304
rect 12508 46264 12548 46304
rect 15340 46264 15380 46304
rect 19276 46264 19316 46304
rect 20380 46264 20420 46304
rect 3688 46096 3728 46136
rect 3770 46096 3810 46136
rect 3852 46096 3892 46136
rect 3934 46096 3974 46136
rect 4016 46096 4056 46136
rect 18808 46096 18848 46136
rect 18890 46096 18930 46136
rect 18972 46096 19012 46136
rect 19054 46096 19094 46136
rect 19136 46096 19176 46136
rect 1852 45928 1892 45968
rect 4684 45928 4724 45968
rect 9772 45928 9812 45968
rect 11404 45928 11444 45968
rect 13420 45928 13460 45968
rect 1468 45844 1508 45884
rect 5068 45844 5108 45884
rect 7468 45844 7508 45884
rect 11836 45844 11876 45884
rect 1228 45760 1268 45800
rect 1612 45760 1652 45800
rect 3916 45676 3956 45716
rect 4058 45676 4098 45716
rect 4396 45676 4436 45716
rect 4551 45676 4591 45716
rect 4674 45676 4714 45716
rect 4852 45676 4892 45716
rect 5000 45718 5040 45758
rect 5164 45760 5204 45800
rect 6915 45760 6955 45800
rect 11596 45760 11636 45800
rect 14668 45760 14708 45800
rect 17548 45760 17588 45800
rect 18316 45760 18356 45800
rect 19756 45760 19796 45800
rect 20140 45760 20180 45800
rect 5285 45676 5325 45716
rect 5443 45676 5483 45716
rect 5587 45676 5627 45716
rect 5701 45676 5741 45716
rect 5827 45676 5867 45716
rect 6004 45676 6044 45716
rect 6220 45676 6260 45716
rect 6362 45676 6402 45716
rect 6796 45676 6836 45716
rect 7033 45676 7073 45716
rect 7177 45676 7217 45716
rect 7315 45676 7355 45716
rect 7429 45676 7469 45716
rect 7756 45676 7796 45716
rect 7875 45676 7915 45716
rect 7993 45676 8033 45716
rect 8332 45676 8372 45716
rect 9580 45676 9620 45716
rect 9964 45676 10004 45716
rect 11212 45676 11252 45716
rect 11980 45676 12020 45716
rect 13228 45676 13268 45716
rect 14179 45676 14219 45716
rect 14284 45676 14324 45716
rect 14764 45676 14804 45716
rect 15244 45676 15284 45716
rect 15732 45676 15772 45716
rect 17827 45676 17867 45716
rect 17932 45676 17972 45716
rect 18412 45676 18452 45716
rect 18892 45676 18932 45716
rect 19380 45676 19420 45716
rect 6700 45592 6740 45632
rect 7660 45592 7700 45632
rect 19996 45592 20036 45632
rect 4204 45508 4244 45548
rect 5923 45508 5963 45548
rect 6508 45508 6548 45548
rect 9772 45508 9812 45548
rect 15916 45508 15956 45548
rect 17308 45508 17348 45548
rect 19564 45508 19604 45548
rect 20380 45508 20420 45548
rect 4928 45340 4968 45380
rect 5010 45340 5050 45380
rect 5092 45340 5132 45380
rect 5174 45340 5214 45380
rect 5256 45340 5296 45380
rect 20048 45340 20088 45380
rect 20130 45340 20170 45380
rect 20212 45340 20252 45380
rect 20294 45340 20334 45380
rect 20376 45340 20416 45380
rect 4204 45172 4244 45212
rect 5452 45172 5492 45212
rect 5731 45172 5771 45212
rect 8140 45172 8180 45212
rect 10636 45172 10676 45212
rect 11932 45172 11972 45212
rect 15244 45172 15284 45212
rect 17452 45172 17492 45212
rect 19756 45172 19796 45212
rect 5633 45088 5673 45128
rect 6316 45088 6356 45128
rect 11107 45079 11147 45119
rect 2764 45004 2804 45044
rect 4012 44995 4052 45035
rect 4396 45004 4436 45044
rect 4565 45004 4605 45044
rect 4684 45004 4724 45044
rect 5068 45004 5108 45044
rect 5190 45004 5230 45044
rect 1228 44920 1268 44960
rect 5305 44962 5345 45002
rect 5407 44995 5447 45035
rect 5836 45004 5876 45044
rect 5932 44995 5972 45035
rect 6110 45004 6150 45044
rect 6412 44995 6452 45035
rect 6748 45004 6788 45044
rect 7049 45004 7089 45044
rect 7219 45004 7259 45044
rect 7564 44995 7604 45035
rect 7675 44995 7715 45035
rect 7795 44995 7835 45035
rect 8236 45004 8276 45044
rect 8453 45004 8493 45044
rect 8716 45004 8756 45044
rect 8835 45004 8875 45044
rect 8953 45004 8993 45044
rect 9196 45004 9236 45044
rect 10444 44995 10484 45035
rect 10819 45004 10859 45044
rect 10924 44995 10964 45035
rect 11199 45004 11239 45044
rect 11380 45004 11420 45044
rect 13486 45004 13526 45044
rect 13617 45004 13657 45044
rect 13996 45004 14036 45044
rect 14572 44995 14612 45035
rect 15052 44995 15092 45035
rect 16012 45004 16052 45044
rect 17260 44995 17300 45035
rect 18019 45004 18059 45044
rect 18124 45004 18164 45044
rect 18508 45004 18548 45044
rect 19084 44995 19124 45035
rect 19564 44995 19604 45035
rect 1612 44920 1652 44960
rect 6892 44920 6932 44960
rect 8371 44911 8411 44951
rect 8620 44920 8660 44960
rect 11692 44920 11732 44960
rect 12652 44920 12692 44960
rect 14092 44920 14132 44960
rect 15724 44920 15764 44960
rect 18604 44920 18644 44960
rect 20140 44920 20180 44960
rect 4204 44836 4244 44876
rect 4876 44836 4916 44876
rect 6988 44836 7028 44876
rect 1468 44752 1508 44792
rect 1852 44752 1892 44792
rect 6115 44752 6155 44792
rect 7948 44752 7988 44792
rect 10819 44752 10859 44792
rect 12412 44752 12452 44792
rect 15484 44752 15524 44792
rect 20380 44752 20420 44792
rect 3688 44584 3728 44624
rect 3770 44584 3810 44624
rect 3852 44584 3892 44624
rect 3934 44584 3974 44624
rect 4016 44584 4056 44624
rect 18808 44584 18848 44624
rect 18890 44584 18930 44624
rect 18972 44584 19012 44624
rect 19054 44584 19094 44624
rect 19136 44584 19176 44624
rect 1852 44416 1892 44456
rect 4675 44416 4715 44456
rect 5452 44416 5492 44456
rect 6604 44416 6644 44456
rect 6844 44416 6884 44456
rect 7180 44416 7220 44456
rect 11164 44416 11204 44456
rect 13420 44416 13460 44456
rect 15052 44416 15092 44456
rect 17644 44416 17684 44456
rect 18172 44416 18212 44456
rect 20140 44416 20180 44456
rect 1468 44332 1508 44372
rect 4460 44323 4500 44363
rect 6124 44332 6164 44372
rect 11548 44332 11588 44372
rect 16012 44332 16052 44372
rect 1228 44248 1268 44288
rect 1612 44248 1652 44288
rect 2860 44248 2900 44288
rect 6220 44248 6260 44288
rect 2371 44164 2411 44204
rect 2476 44164 2516 44204
rect 2956 44164 2996 44204
rect 3436 44164 3476 44204
rect 3924 44164 3964 44204
rect 4483 44164 4523 44204
rect 4915 44164 4955 44204
rect 5015 44197 5055 44237
rect 5479 44206 5519 44246
rect 9763 44248 9803 44288
rect 10540 44248 10580 44288
rect 11404 44248 11444 44288
rect 11788 44248 11828 44288
rect 17836 44248 17876 44288
rect 18412 44248 18452 44288
rect 5356 44164 5396 44204
rect 5593 44164 5633 44204
rect 5695 44197 5735 44237
rect 5884 44164 5924 44204
rect 6056 44122 6096 44162
rect 6341 44164 6381 44204
rect 6505 44137 6545 44177
rect 6709 44164 6749 44204
rect 6940 44164 6980 44204
rect 7180 44164 7220 44204
rect 7372 44164 7412 44204
rect 7564 44164 7604 44204
rect 8812 44164 8852 44204
rect 9187 44164 9227 44204
rect 9643 44164 9683 44204
rect 9868 44164 9908 44204
rect 11980 44164 12020 44204
rect 13228 44164 13268 44204
rect 13612 44164 13652 44204
rect 14860 44164 14900 44204
rect 15340 44164 15380 44204
rect 15619 44164 15659 44204
rect 16204 44164 16244 44204
rect 17452 44164 17492 44204
rect 18700 44164 18740 44204
rect 19948 44164 19988 44204
rect 9388 44080 9428 44120
rect 9498 44080 9538 44120
rect 11164 44080 11204 44120
rect 15724 44080 15764 44120
rect 4108 43996 4148 44036
rect 5164 43996 5204 44036
rect 9004 43996 9044 44036
rect 9283 43996 9323 44036
rect 9955 43996 9995 44036
rect 10300 43996 10340 44036
rect 18076 43996 18116 44036
rect 4928 43828 4968 43868
rect 5010 43828 5050 43868
rect 5092 43828 5132 43868
rect 5174 43828 5214 43868
rect 5256 43828 5296 43868
rect 20048 43828 20088 43868
rect 20130 43828 20170 43868
rect 20212 43828 20252 43868
rect 20294 43828 20334 43868
rect 20376 43828 20416 43868
rect 1468 43660 1508 43700
rect 3916 43660 3956 43700
rect 5068 43660 5108 43700
rect 5923 43660 5963 43700
rect 8236 43660 8276 43700
rect 10348 43660 10388 43700
rect 12652 43660 12692 43700
rect 13084 43660 13124 43700
rect 16156 43660 16196 43700
rect 19756 43660 19796 43700
rect 20380 43660 20420 43700
rect 5825 43576 5865 43616
rect 14332 43576 14372 43616
rect 15436 43576 15476 43616
rect 17740 43576 17780 43616
rect 2476 43492 2516 43532
rect 3724 43483 3764 43523
rect 1228 43408 1268 43448
rect 1612 43408 1652 43448
rect 2092 43408 2132 43448
rect 4348 43450 4388 43490
rect 4586 43492 4626 43532
rect 4867 43492 4907 43532
rect 5164 43492 5204 43532
rect 5399 43492 5439 43532
rect 5500 43492 5540 43532
rect 5644 43492 5684 43532
rect 6028 43492 6068 43532
rect 6124 43483 6164 43523
rect 6499 43492 6539 43532
rect 6604 43492 6644 43532
rect 6988 43492 7028 43532
rect 7564 43483 7604 43523
rect 8044 43483 8084 43523
rect 8908 43492 8948 43532
rect 10156 43483 10196 43523
rect 10915 43492 10955 43532
rect 11020 43492 11060 43532
rect 11404 43492 11444 43532
rect 11980 43483 12020 43523
rect 12460 43483 12500 43523
rect 14188 43492 14228 43532
rect 14572 43492 14612 43532
rect 14809 43492 14849 43532
rect 15052 43492 15092 43532
rect 15331 43492 15371 43532
rect 16300 43492 16340 43532
rect 17548 43483 17588 43523
rect 18019 43492 18059 43532
rect 18124 43492 18164 43532
rect 18508 43492 18548 43532
rect 19084 43483 19124 43523
rect 19564 43483 19604 43523
rect 4483 43408 4523 43448
rect 4684 43408 4724 43448
rect 7084 43408 7124 43448
rect 11500 43408 11540 43448
rect 12844 43408 12884 43448
rect 13420 43408 13460 43448
rect 14476 43408 14516 43448
rect 14691 43408 14731 43448
rect 15916 43408 15956 43448
rect 18604 43408 18644 43448
rect 20140 43408 20180 43448
rect 2332 43324 2372 43364
rect 13180 43324 13220 43364
rect 15724 43324 15764 43364
rect 1852 43240 1892 43280
rect 5356 43240 5396 43280
rect 3688 43072 3728 43112
rect 3770 43072 3810 43112
rect 3852 43072 3892 43112
rect 3934 43072 3974 43112
rect 4016 43072 4056 43112
rect 18808 43072 18848 43112
rect 18890 43072 18930 43112
rect 18972 43072 19012 43112
rect 19054 43072 19094 43112
rect 19136 43072 19176 43112
rect 4588 42904 4628 42944
rect 5347 42904 5387 42944
rect 5932 42904 5972 42944
rect 9004 42904 9044 42944
rect 12892 42904 12932 42944
rect 20380 42904 20420 42944
rect 2236 42820 2276 42860
rect 4012 42820 4052 42860
rect 5164 42820 5204 42860
rect 1228 42736 1268 42776
rect 1612 42736 1652 42776
rect 1996 42736 2036 42776
rect 6796 42736 6836 42776
rect 13132 42736 13172 42776
rect 15523 42736 15563 42776
rect 18508 42736 18548 42776
rect 20140 42736 20180 42776
rect 2572 42652 2612 42692
rect 3820 42652 3860 42692
rect 4204 42652 4244 42692
rect 4492 42652 4532 42692
rect 4684 42652 4724 42692
rect 4972 42652 5012 42692
rect 5345 42652 5385 42692
rect 5644 42652 5684 42692
rect 5836 42652 5876 42692
rect 6028 42652 6068 42692
rect 6307 42652 6347 42692
rect 6412 42652 6452 42692
rect 6892 42652 6932 42692
rect 7372 42652 7412 42692
rect 7891 42652 7931 42692
rect 8332 42652 8372 42692
rect 8587 42652 8627 42692
rect 8707 42652 8747 42692
rect 9676 42652 9716 42692
rect 10924 42652 10964 42692
rect 11308 42652 11348 42692
rect 12556 42652 12596 42692
rect 13315 42652 13355 42692
rect 13804 42652 13844 42692
rect 15052 42652 15092 42692
rect 15383 42652 15423 42692
rect 15628 42652 15668 42692
rect 15916 42652 15956 42692
rect 16108 42652 16148 42692
rect 16300 42652 16340 42692
rect 17548 42652 17588 42692
rect 18019 42652 18059 42692
rect 18124 42652 18164 42692
rect 18604 42652 18644 42692
rect 19084 42652 19124 42692
rect 19572 42652 19612 42692
rect 1852 42568 1892 42608
rect 12748 42568 12788 42608
rect 13626 42568 13666 42608
rect 17740 42568 17780 42608
rect 1468 42484 1508 42524
rect 4348 42484 4388 42524
rect 4867 42484 4907 42524
rect 5548 42484 5588 42524
rect 8044 42484 8084 42524
rect 11116 42484 11156 42524
rect 13411 42484 13451 42524
rect 13516 42484 13556 42524
rect 15244 42484 15284 42524
rect 15715 42484 15755 42524
rect 16012 42484 16052 42524
rect 19756 42484 19796 42524
rect 4928 42316 4968 42356
rect 5010 42316 5050 42356
rect 5092 42316 5132 42356
rect 5174 42316 5214 42356
rect 5256 42316 5296 42356
rect 20048 42316 20088 42356
rect 20130 42316 20170 42356
rect 20212 42316 20252 42356
rect 20294 42316 20334 42356
rect 20376 42316 20416 42356
rect 3292 42148 3332 42188
rect 6988 42148 7028 42188
rect 9100 42148 9140 42188
rect 10732 42148 10772 42188
rect 13228 42148 13268 42188
rect 15052 42148 15092 42188
rect 16204 42148 16244 42188
rect 18028 42148 18068 42188
rect 19660 42148 19700 42188
rect 20380 42148 20420 42188
rect 2860 42064 2900 42104
rect 4972 42064 5012 42104
rect 16001 42064 16041 42104
rect 1420 41980 1460 42020
rect 2668 41971 2708 42011
rect 3532 41980 3572 42020
rect 4780 41971 4820 42011
rect 5251 41980 5291 42020
rect 5356 41980 5396 42020
rect 5740 41980 5780 42020
rect 6316 41971 6356 42011
rect 6796 41971 6836 42011
rect 7660 41980 7700 42020
rect 8908 41971 8948 42011
rect 9292 41980 9332 42020
rect 10540 41971 10580 42011
rect 11491 41980 11531 42020
rect 11596 41980 11636 42020
rect 11980 41980 12020 42020
rect 12556 41971 12596 42011
rect 13036 41971 13076 42011
rect 13420 41980 13460 42020
rect 14668 41971 14708 42011
rect 15148 41980 15188 42020
rect 15283 41971 15323 42011
rect 15385 41980 15425 42020
rect 15627 41980 15667 42020
rect 15845 41980 15885 42020
rect 16302 41971 16342 42011
rect 16588 41980 16628 42020
rect 17836 41971 17876 42011
rect 18220 41980 18260 42020
rect 19468 41971 19508 42011
rect 3052 41896 3092 41936
rect 5836 41896 5876 41936
rect 12076 41896 12116 41936
rect 15532 41896 15572 41936
rect 15763 41887 15803 41927
rect 20140 41896 20180 41936
rect 14860 41728 14900 41768
rect 16003 41728 16043 41768
rect 3688 41560 3728 41600
rect 3770 41560 3810 41600
rect 3852 41560 3892 41600
rect 3934 41560 3974 41600
rect 4016 41560 4056 41600
rect 18808 41560 18848 41600
rect 18890 41560 18930 41600
rect 18972 41560 19012 41600
rect 19054 41560 19094 41600
rect 19136 41560 19176 41600
rect 2668 41392 2708 41432
rect 4540 41392 4580 41432
rect 8908 41392 8948 41432
rect 10540 41392 10580 41432
rect 15619 41392 15659 41432
rect 16252 41392 16292 41432
rect 15148 41308 15188 41348
rect 20380 41308 20420 41348
rect 4780 41224 4820 41264
rect 11308 41224 11348 41264
rect 15292 41224 15332 41264
rect 18604 41224 18644 41264
rect 20140 41224 20180 41264
rect 1228 41140 1268 41180
rect 2476 41140 2516 41180
rect 2860 41140 2900 41180
rect 4108 41140 4148 41180
rect 5164 41140 5204 41180
rect 5356 41140 5396 41180
rect 5548 41140 5588 41180
rect 5687 41140 5727 41180
rect 6019 41140 6059 41180
rect 6316 41140 6356 41180
rect 6497 41140 6537 41180
rect 6796 41140 6836 41180
rect 7084 41140 7124 41180
rect 7468 41140 7508 41180
rect 8716 41140 8756 41180
rect 9100 41140 9140 41180
rect 10348 41140 10388 41180
rect 10798 41140 10838 41180
rect 10905 41140 10945 41180
rect 11404 41140 11444 41180
rect 11884 41140 11924 41180
rect 12372 41140 12412 41180
rect 13708 41140 13748 41180
rect 14956 41140 14996 41180
rect 15436 41140 15476 41180
rect 15916 41140 15956 41180
rect 16108 41140 16148 41180
rect 16396 41140 16436 41180
rect 17644 41140 17684 41180
rect 18115 41140 18155 41180
rect 18220 41140 18260 41180
rect 18700 41140 18740 41180
rect 19180 41140 19220 41180
rect 19668 41140 19708 41180
rect 6700 41056 6740 41096
rect 15614 41056 15654 41096
rect 4300 40972 4340 41012
rect 5347 40972 5387 41012
rect 5875 40972 5915 41012
rect 6220 40972 6260 41012
rect 6595 40972 6635 41012
rect 6940 40972 6980 41012
rect 12556 40972 12596 41012
rect 15820 40972 15860 41012
rect 17836 40972 17876 41012
rect 19852 40972 19892 41012
rect 4928 40804 4968 40844
rect 5010 40804 5050 40844
rect 5092 40804 5132 40844
rect 5174 40804 5214 40844
rect 5256 40804 5296 40844
rect 20048 40804 20088 40844
rect 20130 40804 20170 40844
rect 20212 40804 20252 40844
rect 20294 40804 20334 40844
rect 20376 40804 20416 40844
rect 1852 40636 1892 40676
rect 2236 40636 2276 40676
rect 4396 40636 4436 40676
rect 6796 40636 6836 40676
rect 9628 40636 9668 40676
rect 11212 40636 11252 40676
rect 13507 40636 13547 40676
rect 13612 40636 13652 40676
rect 14092 40636 14132 40676
rect 17644 40636 17684 40676
rect 18364 40636 18404 40676
rect 20332 40636 20372 40676
rect 1468 40552 1508 40592
rect 7747 40552 7787 40592
rect 8476 40552 8516 40592
rect 12926 40552 12966 40592
rect 13027 40552 13067 40592
rect 13132 40552 13172 40592
rect 13987 40552 14027 40592
rect 15676 40552 15716 40592
rect 2659 40468 2699 40508
rect 2769 40468 2809 40508
rect 3148 40468 3188 40508
rect 3724 40459 3764 40499
rect 4216 40468 4256 40508
rect 5059 40468 5099 40508
rect 5164 40468 5204 40508
rect 5548 40468 5588 40508
rect 6124 40459 6164 40499
rect 6604 40459 6644 40499
rect 6974 40468 7014 40508
rect 7084 40468 7124 40508
rect 7276 40468 7316 40508
rect 7415 40468 7455 40508
rect 7658 40468 7698 40508
rect 9772 40468 9812 40508
rect 11020 40459 11060 40499
rect 13228 40459 13268 40499
rect 13406 40468 13446 40508
rect 13708 40459 13748 40499
rect 13886 40468 13926 40508
rect 14188 40459 14228 40499
rect 16204 40468 16244 40508
rect 17452 40459 17492 40499
rect 18595 40468 18635 40508
rect 18700 40468 18740 40508
rect 19084 40468 19124 40508
rect 19660 40459 19700 40499
rect 20140 40459 20180 40499
rect 1228 40384 1268 40424
rect 1612 40384 1652 40424
rect 1996 40384 2036 40424
rect 3244 40384 3284 40424
rect 5644 40384 5684 40424
rect 7555 40384 7595 40424
rect 8236 40384 8276 40424
rect 8620 40384 8660 40424
rect 9196 40384 9236 40424
rect 9388 40384 9428 40424
rect 12556 40384 12596 40424
rect 14668 40384 14708 40424
rect 15052 40384 15092 40424
rect 15436 40384 15476 40424
rect 15820 40384 15860 40424
rect 16060 40384 16100 40424
rect 18124 40384 18164 40424
rect 19180 40384 19220 40424
rect 8860 40300 8900 40340
rect 12796 40300 12836 40340
rect 15292 40300 15332 40340
rect 6988 40216 7028 40256
rect 8956 40216 8996 40256
rect 14908 40216 14948 40256
rect 3688 40048 3728 40088
rect 3770 40048 3810 40088
rect 3852 40048 3892 40088
rect 3934 40048 3974 40088
rect 4016 40048 4056 40088
rect 18808 40048 18848 40088
rect 18890 40048 18930 40088
rect 18972 40048 19012 40088
rect 19054 40048 19094 40088
rect 19136 40048 19176 40088
rect 1468 39880 1508 39920
rect 1852 39880 1892 39920
rect 6403 39880 6443 39920
rect 6883 39880 6923 39920
rect 17740 39880 17780 39920
rect 18748 39880 18788 39920
rect 20332 39880 20372 39920
rect 4732 39796 4772 39836
rect 6028 39796 6068 39836
rect 11068 39796 11108 39836
rect 12028 39796 12068 39836
rect 18364 39796 18404 39836
rect 1228 39712 1268 39752
rect 1612 39712 1652 39752
rect 1996 39712 2036 39752
rect 3148 39712 3188 39752
rect 6127 39712 6167 39752
rect 10828 39712 10868 39752
rect 12387 39712 12427 39752
rect 13699 39712 13739 39752
rect 14668 39712 14708 39752
rect 18124 39712 18164 39752
rect 18508 39712 18548 39752
rect 2659 39628 2699 39668
rect 2764 39628 2804 39668
rect 3244 39628 3284 39668
rect 3724 39628 3764 39668
rect 4212 39628 4252 39668
rect 4588 39628 4628 39668
rect 4732 39628 4772 39668
rect 4876 39628 4916 39668
rect 5059 39628 5099 39668
rect 5164 39628 5204 39668
rect 5303 39628 5343 39668
rect 5443 39628 5483 39668
rect 5548 39628 5588 39668
rect 5788 39628 5828 39668
rect 5953 39628 5993 39668
rect 6259 39628 6299 39668
rect 6700 39628 6740 39668
rect 7180 39628 7220 39668
rect 7564 39628 7604 39668
rect 8820 39628 8860 39668
rect 9196 39628 9236 39668
rect 10452 39628 10492 39668
rect 11884 39628 11924 39668
rect 12268 39628 12308 39668
rect 12505 39628 12545 39668
rect 12748 39628 12788 39668
rect 13027 39628 13067 39668
rect 13559 39628 13599 39668
rect 13804 39628 13844 39668
rect 14179 39628 14219 39668
rect 14284 39628 14324 39668
rect 14764 39628 14804 39668
rect 15244 39628 15284 39668
rect 15763 39628 15803 39668
rect 16300 39628 16340 39668
rect 17548 39628 17588 39668
rect 18892 39628 18932 39668
rect 20140 39628 20180 39668
rect 2236 39544 2276 39584
rect 4963 39544 5003 39584
rect 6401 39544 6441 39584
rect 6604 39544 6644 39584
rect 6878 39544 6918 39584
rect 12172 39544 12212 39584
rect 13132 39544 13172 39584
rect 13468 39544 13508 39584
rect 4396 39460 4436 39500
rect 5635 39460 5675 39500
rect 7084 39460 7124 39500
rect 9004 39460 9044 39500
rect 10636 39460 10676 39500
rect 13891 39460 13931 39500
rect 15916 39460 15956 39500
rect 4928 39292 4968 39332
rect 5010 39292 5050 39332
rect 5092 39292 5132 39332
rect 5174 39292 5214 39332
rect 5256 39292 5296 39332
rect 20048 39292 20088 39332
rect 20130 39292 20170 39332
rect 20212 39292 20252 39332
rect 20294 39292 20334 39332
rect 20376 39292 20416 39332
rect 1468 39124 1508 39164
rect 3916 39124 3956 39164
rect 5932 39124 5972 39164
rect 6604 39124 6644 39164
rect 8812 39124 8852 39164
rect 12556 39124 12596 39164
rect 13948 39124 13988 39164
rect 15916 39124 15956 39164
rect 16732 39124 16772 39164
rect 13612 39040 13652 39080
rect 14332 39040 14372 39080
rect 2476 38956 2516 38996
rect 3724 38947 3764 38987
rect 4195 38956 4235 38996
rect 4300 38956 4340 38996
rect 4684 38956 4724 38996
rect 5260 38947 5300 38987
rect 5740 38947 5780 38987
rect 6124 38956 6164 38996
rect 6239 38956 6279 38996
rect 6412 38956 6452 38996
rect 6604 38956 6644 38996
rect 6796 38956 6836 38996
rect 7054 38956 7094 38996
rect 7171 38989 7211 39029
rect 7564 38956 7604 38996
rect 8140 38947 8180 38987
rect 8620 38947 8660 38987
rect 9004 38956 9044 38996
rect 10252 38947 10292 38987
rect 11116 38956 11156 38996
rect 12364 38947 12404 38987
rect 12748 38956 12788 38996
rect 12940 38956 12980 38996
rect 13228 38956 13268 38996
rect 13507 38956 13547 38996
rect 14476 38956 14516 38996
rect 15724 38947 15764 38987
rect 16972 38956 17012 38996
rect 18220 38947 18260 38987
rect 18700 38956 18740 38996
rect 19948 38947 19988 38987
rect 1228 38872 1268 38912
rect 1612 38872 1652 38912
rect 1996 38872 2036 38912
rect 2236 38872 2276 38912
rect 4780 38872 4820 38912
rect 7660 38872 7700 38912
rect 14092 38872 14132 38912
rect 16300 38872 16340 38912
rect 16492 38872 16532 38912
rect 1852 38704 1892 38744
rect 6124 38704 6164 38744
rect 10444 38704 10484 38744
rect 12748 38704 12788 38744
rect 16060 38704 16100 38744
rect 18412 38704 18452 38744
rect 20140 38704 20180 38744
rect 3688 38536 3728 38576
rect 3770 38536 3810 38576
rect 3852 38536 3892 38576
rect 3934 38536 3974 38576
rect 4016 38536 4056 38576
rect 18808 38536 18848 38576
rect 18890 38536 18930 38576
rect 18972 38536 19012 38576
rect 19054 38536 19094 38576
rect 19136 38536 19176 38576
rect 2668 38368 2708 38408
rect 4300 38368 4340 38408
rect 12076 38368 12116 38408
rect 12412 38368 12452 38408
rect 14668 38368 14708 38408
rect 15676 38368 15716 38408
rect 6124 38284 6164 38324
rect 6988 38284 7028 38324
rect 4492 38200 4532 38240
rect 5283 38200 5323 38240
rect 6595 38200 6635 38240
rect 8428 38200 8468 38240
rect 8812 38200 8852 38240
rect 9676 38200 9716 38240
rect 12643 38200 12683 38240
rect 15052 38200 15092 38240
rect 15436 38200 15476 38240
rect 15820 38200 15860 38240
rect 16492 38200 16532 38240
rect 18988 38200 19028 38240
rect 1228 38116 1268 38156
rect 2476 38116 2516 38156
rect 2860 38116 2900 38156
rect 4108 38116 4148 38156
rect 5164 38116 5204 38156
rect 5401 38116 5441 38156
rect 5548 38116 5588 38156
rect 5731 38116 5771 38156
rect 5836 38116 5876 38156
rect 6028 38116 6068 38156
rect 6153 38116 6193 38156
rect 6316 38116 6356 38156
rect 6475 38116 6515 38156
rect 6700 38116 6740 38156
rect 6988 38116 7028 38156
rect 7103 38116 7143 38156
rect 7276 38116 7316 38156
rect 10636 38116 10676 38156
rect 11884 38116 11924 38156
rect 12268 38116 12308 38156
rect 12503 38116 12543 38156
rect 12748 38116 12788 38156
rect 13228 38116 13268 38156
rect 14476 38116 14516 38156
rect 16780 38116 16820 38156
rect 18028 38116 18068 38156
rect 18499 38134 18539 38174
rect 18601 38116 18641 38156
rect 19084 38116 19124 38156
rect 19564 38116 19604 38156
rect 20083 38116 20123 38156
rect 5635 38032 5675 38072
rect 16060 38032 16100 38072
rect 4732 37948 4772 37988
rect 5068 37948 5108 37988
rect 6787 37948 6827 37988
rect 8188 37948 8228 37988
rect 8572 37948 8612 37988
rect 9436 37948 9476 37988
rect 12835 37948 12875 37988
rect 14812 37948 14852 37988
rect 16252 37948 16292 37988
rect 18220 37948 18260 37988
rect 20236 37948 20276 37988
rect 4928 37780 4968 37820
rect 5010 37780 5050 37820
rect 5092 37780 5132 37820
rect 5174 37780 5214 37820
rect 5256 37780 5296 37820
rect 20048 37780 20088 37820
rect 20130 37780 20170 37820
rect 20212 37780 20252 37820
rect 20294 37780 20334 37820
rect 20376 37780 20416 37820
rect 5452 37612 5492 37652
rect 8035 37612 8075 37652
rect 12172 37612 12212 37652
rect 13372 37612 13412 37652
rect 7084 37528 7124 37568
rect 8247 37528 8287 37568
rect 17884 37528 17924 37568
rect 1228 37444 1268 37484
rect 2476 37435 2516 37475
rect 4012 37444 4052 37484
rect 5260 37435 5300 37475
rect 5644 37444 5684 37484
rect 6892 37435 6932 37475
rect 7372 37435 7412 37475
rect 7471 37424 7511 37464
rect 7603 37435 7643 37475
rect 7939 37444 7979 37484
rect 9292 37435 9332 37475
rect 10540 37444 10580 37484
rect 10732 37444 10772 37484
rect 11980 37435 12020 37475
rect 12619 37444 12659 37484
rect 12844 37444 12884 37484
rect 13516 37444 13556 37484
rect 13804 37444 13844 37484
rect 15052 37435 15092 37475
rect 15628 37435 15668 37475
rect 16876 37444 16916 37484
rect 18499 37444 18539 37484
rect 18604 37444 18644 37484
rect 18988 37444 19028 37484
rect 19564 37435 19604 37475
rect 20044 37435 20084 37475
rect 2860 37360 2900 37400
rect 3100 37360 3140 37400
rect 3244 37360 3284 37400
rect 3628 37360 3668 37400
rect 8716 37360 8756 37400
rect 12739 37360 12779 37400
rect 12940 37360 12980 37400
rect 13132 37360 13172 37400
rect 13660 37360 13700 37400
rect 17068 37360 17108 37400
rect 17308 37360 17348 37400
rect 17644 37360 17684 37400
rect 18124 37360 18164 37400
rect 19084 37360 19124 37400
rect 2668 37276 2708 37316
rect 8956 37276 8996 37316
rect 15244 37276 15284 37316
rect 3484 37192 3524 37232
rect 3868 37192 3908 37232
rect 7084 37192 7124 37232
rect 7756 37192 7796 37232
rect 8236 37192 8276 37232
rect 9100 37192 9140 37232
rect 15436 37192 15476 37232
rect 17404 37192 17444 37232
rect 20275 37192 20315 37232
rect 3688 37024 3728 37064
rect 3770 37024 3810 37064
rect 3852 37024 3892 37064
rect 3934 37024 3974 37064
rect 4016 37024 4056 37064
rect 18808 37024 18848 37064
rect 18890 37024 18930 37064
rect 18972 37024 19012 37064
rect 19054 37024 19094 37064
rect 19136 37024 19176 37064
rect 1852 36856 1892 36896
rect 7948 36856 7988 36896
rect 18364 36856 18404 36896
rect 20140 36856 20180 36896
rect 12364 36772 12404 36812
rect 1228 36688 1268 36728
rect 1612 36688 1652 36728
rect 2764 36688 2804 36728
rect 4204 36688 4244 36728
rect 8227 36688 8267 36728
rect 9772 36688 9812 36728
rect 13708 36688 13748 36728
rect 14860 36688 14900 36728
rect 16012 36688 16052 36728
rect 17740 36688 17780 36728
rect 2275 36604 2315 36644
rect 2380 36604 2420 36644
rect 2860 36604 2900 36644
rect 3340 36604 3380 36644
rect 3828 36604 3868 36644
rect 4876 36604 4916 36644
rect 6124 36604 6164 36644
rect 6508 36604 6548 36644
rect 7756 36604 7796 36644
rect 8087 36604 8127 36644
rect 8332 36604 8372 36644
rect 8803 36604 8843 36644
rect 9292 36604 9332 36644
rect 9868 36604 9908 36644
rect 10252 36604 10292 36644
rect 10370 36604 10410 36644
rect 10924 36604 10964 36644
rect 12172 36604 12212 36644
rect 12739 36604 12779 36644
rect 13228 36604 13268 36644
rect 13804 36604 13844 36644
rect 14188 36604 14228 36644
rect 14301 36623 14341 36663
rect 14668 36604 14708 36644
rect 15523 36604 15563 36644
rect 15628 36604 15668 36644
rect 16108 36604 16148 36644
rect 16588 36604 16628 36644
rect 17107 36604 17147 36644
rect 17399 36604 17439 36644
rect 17539 36604 17579 36644
rect 17644 36604 17684 36644
rect 18220 36604 18260 36644
rect 18508 36604 18548 36644
rect 18700 36604 18740 36644
rect 19948 36604 19988 36644
rect 1468 36520 1508 36560
rect 4444 36520 4484 36560
rect 8611 36520 8651 36560
rect 17918 36520 17958 36560
rect 4012 36436 4052 36476
rect 6316 36436 6356 36476
rect 8419 36436 8459 36476
rect 12556 36436 12596 36476
rect 14524 36436 14564 36476
rect 15100 36436 15140 36476
rect 17260 36436 17300 36476
rect 18019 36436 18059 36476
rect 18124 36436 18164 36476
rect 4928 36268 4968 36308
rect 5010 36268 5050 36308
rect 5092 36268 5132 36308
rect 5174 36268 5214 36308
rect 5256 36268 5296 36308
rect 20048 36268 20088 36308
rect 20130 36268 20170 36308
rect 20212 36268 20252 36308
rect 20294 36268 20334 36308
rect 20376 36268 20416 36308
rect 4012 36100 4052 36140
rect 11596 36100 11636 36140
rect 12739 36100 12779 36140
rect 17827 36100 17867 36140
rect 11875 36016 11915 36056
rect 17932 36016 17972 36056
rect 2275 35932 2315 35972
rect 2385 35932 2425 35972
rect 2764 35932 2804 35972
rect 3340 35923 3380 35963
rect 3820 35923 3860 35963
rect 4492 35932 4532 35972
rect 5740 35923 5780 35963
rect 6124 35932 6164 35972
rect 6307 35932 6347 35972
rect 6892 35932 6932 35972
rect 8140 35923 8180 35963
rect 8524 35932 8564 35972
rect 9772 35923 9812 35963
rect 10156 35932 10196 35972
rect 11404 35923 11444 35963
rect 11788 35932 11828 35972
rect 11971 35932 12011 35972
rect 12083 35900 12123 35940
rect 12259 35932 12299 35972
rect 12364 35923 12404 35963
rect 12508 35923 12548 35963
rect 12639 35932 12679 35972
rect 12777 35932 12817 35972
rect 13036 35932 13076 35972
rect 14284 35923 14324 35963
rect 15724 35932 15764 35972
rect 1228 35848 1268 35888
rect 1612 35848 1652 35888
rect 2860 35848 2900 35888
rect 6700 35848 6740 35888
rect 14860 35848 14900 35888
rect 15100 35848 15140 35888
rect 15436 35848 15476 35888
rect 15628 35848 15668 35888
rect 15843 35848 15883 35888
rect 15964 35890 16004 35930
rect 16108 35932 16148 35972
rect 17356 35923 17396 35963
rect 17726 35932 17766 35972
rect 18028 35923 18068 35963
rect 18316 35932 18356 35972
rect 18595 35932 18635 35972
rect 18700 35932 18740 35972
rect 19084 35932 19124 35972
rect 19660 35923 19700 35963
rect 20140 35923 20180 35963
rect 20371 35932 20411 35972
rect 19180 35848 19220 35888
rect 5932 35764 5972 35804
rect 6307 35764 6347 35804
rect 17548 35764 17588 35804
rect 1468 35680 1508 35720
rect 1852 35680 1892 35720
rect 6460 35680 6500 35720
rect 8332 35680 8372 35720
rect 9964 35680 10004 35720
rect 14476 35680 14516 35720
rect 15196 35680 15236 35720
rect 18172 35680 18212 35720
rect 3688 35512 3728 35552
rect 3770 35512 3810 35552
rect 3852 35512 3892 35552
rect 3934 35512 3974 35552
rect 4016 35512 4056 35552
rect 18808 35512 18848 35552
rect 18890 35512 18930 35552
rect 18972 35512 19012 35552
rect 19054 35512 19094 35552
rect 19136 35512 19176 35552
rect 3532 35344 3572 35384
rect 5356 35344 5396 35384
rect 6988 35344 7028 35384
rect 8044 35344 8084 35384
rect 9676 35344 9716 35384
rect 11404 35344 11444 35384
rect 17932 35344 17972 35384
rect 20236 35344 20276 35384
rect 13036 35260 13076 35300
rect 1228 35176 1268 35216
rect 1612 35176 1652 35216
rect 7324 35176 7364 35216
rect 14284 35176 14324 35216
rect 16492 35176 16532 35216
rect 16771 35176 16811 35216
rect 18316 35176 18356 35216
rect 2092 35092 2132 35132
rect 3340 35092 3380 35132
rect 3916 35092 3956 35132
rect 5164 35092 5204 35132
rect 5548 35092 5588 35132
rect 6796 35092 6836 35132
rect 7180 35092 7220 35132
rect 7492 35092 7532 35132
rect 7651 35092 7691 35132
rect 7768 35092 7808 35132
rect 7939 35092 7979 35132
rect 8041 35092 8081 35132
rect 8268 35092 8308 35132
rect 9484 35092 9524 35132
rect 9964 35092 10004 35132
rect 11212 35092 11252 35132
rect 11596 35092 11636 35132
rect 12844 35092 12884 35132
rect 13228 35092 13268 35132
rect 13367 35092 13407 35132
rect 13795 35092 13835 35132
rect 13900 35092 13940 35132
rect 14380 35092 14420 35132
rect 14860 35092 14900 35132
rect 15348 35092 15388 35132
rect 15820 35092 15860 35132
rect 16012 35092 16052 35132
rect 16156 35092 16196 35132
rect 16291 35092 16331 35132
rect 16396 35092 16436 35132
rect 16631 35092 16671 35132
rect 16876 35092 16916 35132
rect 17260 35092 17300 35132
rect 17539 35092 17579 35132
rect 18604 35092 18644 35132
rect 18796 35092 18836 35132
rect 20044 35092 20084 35132
rect 1468 35008 1508 35048
rect 15916 35008 15956 35048
rect 17644 35008 17684 35048
rect 18076 35008 18116 35048
rect 1852 34924 1892 34964
rect 7555 34924 7595 34964
rect 13516 34924 13556 34964
rect 15532 34924 15572 34964
rect 16963 34924 17003 34964
rect 18460 34924 18500 34964
rect 4928 34756 4968 34796
rect 5010 34756 5050 34796
rect 5092 34756 5132 34796
rect 5174 34756 5214 34796
rect 5256 34756 5296 34796
rect 20048 34756 20088 34796
rect 20130 34756 20170 34796
rect 20212 34756 20252 34796
rect 20294 34756 20334 34796
rect 20376 34756 20416 34796
rect 17251 34588 17291 34628
rect 11155 34504 11195 34544
rect 12316 34504 12356 34544
rect 13900 34504 13940 34544
rect 16636 34504 16676 34544
rect 17463 34504 17503 34544
rect 19084 34504 19124 34544
rect 19612 34504 19652 34544
rect 19996 34504 20036 34544
rect 20380 34504 20420 34544
rect 2275 34420 2315 34460
rect 2572 34420 2612 34460
rect 2851 34420 2891 34460
rect 2956 34420 2996 34460
rect 3340 34420 3380 34460
rect 3916 34411 3956 34451
rect 4396 34411 4436 34451
rect 6028 34420 6068 34460
rect 7276 34411 7316 34451
rect 7660 34420 7700 34460
rect 8908 34411 8948 34451
rect 9379 34420 9419 34460
rect 9484 34420 9524 34460
rect 9868 34420 9908 34460
rect 10444 34411 10484 34451
rect 10924 34411 10964 34451
rect 12460 34420 12500 34460
rect 13708 34411 13748 34451
rect 14275 34420 14315 34460
rect 14380 34420 14420 34460
rect 14764 34420 14804 34460
rect 15340 34411 15380 34451
rect 15820 34411 15860 34451
rect 17155 34420 17195 34460
rect 17644 34420 17684 34460
rect 18892 34411 18932 34451
rect 1228 34336 1268 34376
rect 1612 34336 1652 34376
rect 1852 34336 1892 34376
rect 3436 34336 3476 34376
rect 4627 34336 4667 34376
rect 4780 34336 4820 34376
rect 5164 34336 5204 34376
rect 5404 34336 5444 34376
rect 5836 34336 5876 34376
rect 9964 34336 10004 34376
rect 12076 34336 12116 34376
rect 14860 34336 14900 34376
rect 16396 34336 16436 34376
rect 16780 34336 16820 34376
rect 17020 34336 17060 34376
rect 19372 34336 19412 34376
rect 19756 34336 19796 34376
rect 20140 34336 20180 34376
rect 5020 34252 5060 34292
rect 1468 34168 1508 34208
rect 2572 34168 2612 34208
rect 5596 34168 5636 34208
rect 7468 34168 7508 34208
rect 9100 34168 9140 34208
rect 16051 34168 16091 34208
rect 17452 34168 17492 34208
rect 3688 34000 3728 34040
rect 3770 34000 3810 34040
rect 3852 34000 3892 34040
rect 3934 34000 3974 34040
rect 4016 34000 4056 34040
rect 18808 34000 18848 34040
rect 18890 34000 18930 34040
rect 18972 34000 19012 34040
rect 19054 34000 19094 34040
rect 19136 34000 19176 34040
rect 2668 33832 2708 33872
rect 5836 33832 5876 33872
rect 7468 33832 7508 33872
rect 15628 33832 15668 33872
rect 16876 33832 16916 33872
rect 11164 33748 11204 33788
rect 4012 33664 4052 33704
rect 9868 33664 9908 33704
rect 1228 33580 1268 33620
rect 2476 33580 2516 33620
rect 3027 33580 3067 33620
rect 3137 33613 3177 33653
rect 3248 33580 3288 33620
rect 3820 33580 3860 33620
rect 4396 33580 4436 33620
rect 5644 33580 5684 33620
rect 6028 33580 6068 33620
rect 7276 33580 7316 33620
rect 7660 33580 7700 33620
rect 8908 33580 8948 33620
rect 9379 33580 9419 33620
rect 9484 33580 9524 33620
rect 9964 33580 10004 33620
rect 10444 33580 10484 33620
rect 10932 33580 10972 33620
rect 12556 33580 12596 33620
rect 13804 33580 13844 33620
rect 14188 33580 14228 33620
rect 15436 33580 15476 33620
rect 16204 33580 16244 33620
rect 16483 33580 16523 33620
rect 17068 33580 17108 33620
rect 18316 33580 18356 33620
rect 18700 33580 18740 33620
rect 19948 33580 19988 33620
rect 3518 33496 3558 33536
rect 9100 33496 9140 33536
rect 16588 33496 16628 33536
rect 2860 33412 2900 33452
rect 3619 33412 3659 33452
rect 3724 33412 3764 33452
rect 4252 33412 4292 33452
rect 11116 33412 11156 33452
rect 13996 33412 14036 33452
rect 18508 33412 18548 33452
rect 20140 33412 20180 33452
rect 4928 33244 4968 33284
rect 5010 33244 5050 33284
rect 5092 33244 5132 33284
rect 5174 33244 5214 33284
rect 5256 33244 5296 33284
rect 20048 33244 20088 33284
rect 20130 33244 20170 33284
rect 20212 33244 20252 33284
rect 20294 33244 20334 33284
rect 20376 33244 20416 33284
rect 3052 33076 3092 33116
rect 4684 33076 4724 33116
rect 7948 33076 7988 33116
rect 10156 33076 10196 33116
rect 15436 33076 15476 33116
rect 17164 33076 17204 33116
rect 20140 33076 20180 33116
rect 13420 32992 13460 33032
rect 1612 32908 1652 32948
rect 2860 32899 2900 32939
rect 3244 32908 3284 32948
rect 4492 32899 4532 32939
rect 4972 32908 5012 32948
rect 5251 32908 5291 32948
rect 5361 32908 5401 32948
rect 5740 32908 5780 32948
rect 6316 32899 6356 32939
rect 6796 32899 6836 32939
rect 7660 32908 7700 32948
rect 7802 32908 7842 32948
rect 8140 32908 8180 32948
rect 8255 32908 8295 32948
rect 8428 32908 8468 32948
rect 8716 32908 8756 32948
rect 9964 32899 10004 32939
rect 10540 32899 10580 32939
rect 11788 32908 11828 32948
rect 11980 32908 12020 32948
rect 13228 32899 13268 32939
rect 13699 32908 13739 32948
rect 13804 32908 13844 32948
rect 14188 32908 14228 32948
rect 14764 32899 14804 32939
rect 15244 32899 15284 32939
rect 15724 32908 15764 32948
rect 16972 32899 17012 32939
rect 18403 32908 18443 32948
rect 18508 32908 18548 32948
rect 18892 32908 18932 32948
rect 19468 32899 19508 32939
rect 19948 32899 19988 32939
rect 1228 32824 1268 32864
rect 5836 32824 5876 32864
rect 7276 32824 7316 32864
rect 14284 32824 14324 32864
rect 17548 32824 17588 32864
rect 17932 32824 17972 32864
rect 18988 32824 19028 32864
rect 8140 32740 8180 32780
rect 1468 32656 1508 32696
rect 4828 32656 4868 32696
rect 7027 32656 7067 32696
rect 7516 32656 7556 32696
rect 10348 32656 10388 32696
rect 17308 32656 17348 32696
rect 17692 32656 17732 32696
rect 3688 32488 3728 32528
rect 3770 32488 3810 32528
rect 3852 32488 3892 32528
rect 3934 32488 3974 32528
rect 4016 32488 4056 32528
rect 18808 32488 18848 32528
rect 18890 32488 18930 32528
rect 18972 32488 19012 32528
rect 19054 32488 19094 32528
rect 19136 32488 19176 32528
rect 4780 32320 4820 32360
rect 6412 32320 6452 32360
rect 7900 32320 7940 32360
rect 12028 32320 12068 32360
rect 17068 32320 17108 32360
rect 18172 32320 18212 32360
rect 2668 32236 2708 32276
rect 3091 32143 3131 32183
rect 6604 32152 6644 32192
rect 6988 32152 7028 32192
rect 7372 32152 7412 32192
rect 8140 32152 8180 32192
rect 8332 32152 8372 32192
rect 8716 32152 8756 32192
rect 8956 32152 8996 32192
rect 9196 32152 9236 32192
rect 10252 32152 10292 32192
rect 11788 32152 11828 32192
rect 12364 32152 12404 32192
rect 14188 32152 14228 32192
rect 17260 32152 17300 32192
rect 17932 32152 17972 32192
rect 18892 32152 18932 32192
rect 1228 32068 1268 32108
rect 2476 32068 2516 32108
rect 2955 32068 2995 32108
rect 3193 32068 3233 32108
rect 3340 32068 3380 32108
rect 4588 32068 4628 32108
rect 4972 32068 5012 32108
rect 6220 32068 6260 32108
rect 9763 32068 9803 32108
rect 9868 32068 9908 32108
rect 10348 32068 10388 32108
rect 10828 32068 10868 32108
rect 11347 32068 11387 32108
rect 13699 32068 13739 32108
rect 13804 32068 13844 32108
rect 14284 32068 14324 32108
rect 14764 32068 14804 32108
rect 15252 32068 15292 32108
rect 15628 32068 15668 32108
rect 16876 32068 16916 32108
rect 18403 32068 18443 32108
rect 18508 32068 18548 32108
rect 18988 32068 19028 32108
rect 19468 32068 19508 32108
rect 19956 32068 19996 32108
rect 2860 31900 2900 31940
rect 6844 31900 6884 31940
rect 7228 31900 7268 31940
rect 7612 31900 7652 31940
rect 8572 31900 8612 31940
rect 9436 31900 9476 31940
rect 11500 31900 11540 31940
rect 12124 31900 12164 31940
rect 15436 31900 15476 31940
rect 17500 31900 17540 31940
rect 20140 31900 20180 31940
rect 4928 31732 4968 31772
rect 5010 31732 5050 31772
rect 5092 31732 5132 31772
rect 5174 31732 5214 31772
rect 5256 31732 5296 31772
rect 20048 31732 20088 31772
rect 20130 31732 20170 31772
rect 20212 31732 20252 31772
rect 20294 31732 20334 31772
rect 20376 31732 20416 31772
rect 6403 31564 6443 31604
rect 9964 31564 10004 31604
rect 11596 31564 11636 31604
rect 18508 31564 18548 31604
rect 20236 31564 20276 31604
rect 3052 31480 3092 31520
rect 4971 31480 5011 31520
rect 5836 31480 5876 31520
rect 13420 31480 13460 31520
rect 14572 31480 14612 31520
rect 15244 31480 15284 31520
rect 16540 31480 16580 31520
rect 1420 31396 1460 31436
rect 2668 31387 2708 31427
rect 3244 31387 3284 31427
rect 4492 31396 4532 31436
rect 5101 31396 5141 31436
rect 5356 31396 5396 31436
rect 5633 31396 5673 31436
rect 5930 31363 5970 31403
rect 6071 31396 6111 31436
rect 6316 31396 6356 31436
rect 6796 31396 6836 31436
rect 8044 31387 8084 31427
rect 8524 31396 8564 31436
rect 9772 31387 9812 31427
rect 10156 31396 10196 31436
rect 11404 31387 11444 31427
rect 11980 31396 12020 31436
rect 13228 31387 13268 31427
rect 13900 31396 13940 31436
rect 14188 31396 14228 31436
rect 14467 31396 14507 31436
rect 15038 31396 15078 31436
rect 15340 31387 15380 31427
rect 17068 31396 17108 31436
rect 18316 31387 18356 31427
rect 18796 31396 18836 31436
rect 20044 31387 20084 31427
rect 6211 31312 6251 31352
rect 15532 31312 15572 31352
rect 15916 31312 15956 31352
rect 16300 31312 16340 31352
rect 16876 31312 16916 31352
rect 2860 31144 2900 31184
rect 4684 31144 4724 31184
rect 5635 31144 5675 31184
rect 8236 31144 8276 31184
rect 13756 31144 13796 31184
rect 14860 31144 14900 31184
rect 15043 31144 15083 31184
rect 15772 31144 15812 31184
rect 16156 31144 16196 31184
rect 16636 31144 16676 31184
rect 3688 30976 3728 31016
rect 3770 30976 3810 31016
rect 3852 30976 3892 31016
rect 3934 30976 3974 31016
rect 4016 30976 4056 31016
rect 18808 30976 18848 31016
rect 18890 30976 18930 31016
rect 18972 30976 19012 31016
rect 19054 30976 19094 31016
rect 19136 30976 19176 31016
rect 2668 30808 2708 30848
rect 4483 30808 4523 30848
rect 10780 30808 10820 30848
rect 11164 30808 11204 30848
rect 14572 30808 14612 30848
rect 18844 30808 18884 30848
rect 19996 30808 20036 30848
rect 20380 30808 20420 30848
rect 4300 30724 4340 30764
rect 19612 30724 19652 30764
rect 7468 30640 7508 30680
rect 10540 30640 10580 30680
rect 10924 30640 10964 30680
rect 13555 30631 13595 30671
rect 16972 30640 17012 30680
rect 18604 30640 18644 30680
rect 18988 30640 19028 30680
rect 19372 30640 19412 30680
rect 19756 30640 19796 30680
rect 20140 30640 20180 30680
rect 1228 30556 1268 30596
rect 2476 30556 2516 30596
rect 2860 30556 2900 30596
rect 4108 30556 4148 30596
rect 4780 30556 4820 30596
rect 5068 30556 5108 30596
rect 5260 30556 5300 30596
rect 6508 30556 6548 30596
rect 6979 30556 7019 30596
rect 7084 30556 7124 30596
rect 7564 30556 7604 30596
rect 8044 30556 8084 30596
rect 8563 30556 8603 30596
rect 9100 30556 9140 30596
rect 10348 30556 10388 30596
rect 11308 30556 11348 30596
rect 12556 30556 12596 30596
rect 13036 30556 13076 30596
rect 13324 30556 13364 30596
rect 13429 30556 13469 30596
rect 13657 30556 13697 30596
rect 13900 30556 13940 30596
rect 14179 30556 14219 30596
rect 14764 30556 14804 30596
rect 16012 30556 16052 30596
rect 16483 30556 16523 30596
rect 16588 30556 16628 30596
rect 17068 30556 17108 30596
rect 17548 30556 17588 30596
rect 18036 30556 18076 30596
rect 4478 30472 4518 30512
rect 6700 30472 6740 30512
rect 8908 30472 8948 30512
rect 12748 30472 12788 30512
rect 13180 30472 13220 30512
rect 14284 30472 14324 30512
rect 16204 30472 16244 30512
rect 19228 30472 19268 30512
rect 4684 30388 4724 30428
rect 4924 30388 4964 30428
rect 8716 30388 8756 30428
rect 18220 30388 18260 30428
rect 4928 30220 4968 30260
rect 5010 30220 5050 30260
rect 5092 30220 5132 30260
rect 5174 30220 5214 30260
rect 5256 30220 5296 30260
rect 20048 30220 20088 30260
rect 20130 30220 20170 30260
rect 20212 30220 20252 30260
rect 20294 30220 20334 30260
rect 20376 30220 20416 30260
rect 2860 30052 2900 30092
rect 3052 30052 3092 30092
rect 13987 30052 14027 30092
rect 14467 30052 14507 30092
rect 14947 30052 14987 30092
rect 15340 30052 15380 30092
rect 18892 30052 18932 30092
rect 19996 30052 20036 30092
rect 20380 30052 20420 30092
rect 6412 29968 6452 30008
rect 8860 29968 8900 30008
rect 19180 29968 19220 30008
rect 1420 29884 1460 29924
rect 2668 29875 2708 29915
rect 3244 29875 3284 29915
rect 4492 29884 4532 29924
rect 4780 29884 4820 29924
rect 4972 29884 5012 29924
rect 6220 29875 6260 29915
rect 6691 29884 6731 29924
rect 6796 29884 6836 29924
rect 7180 29884 7220 29924
rect 7756 29875 7796 29915
rect 8236 29875 8276 29915
rect 9004 29884 9044 29924
rect 9196 29884 9236 29924
rect 9667 29884 9707 29924
rect 9772 29884 9812 29924
rect 10156 29884 10196 29924
rect 10732 29875 10772 29915
rect 11212 29875 11252 29915
rect 13036 29884 13076 29924
rect 13324 29884 13364 29924
rect 13507 29884 13547 29924
rect 13655 29884 13695 29924
rect 13898 29884 13938 29924
rect 14155 29884 14195 29924
rect 14361 29884 14401 29924
rect 14620 29884 14660 29924
rect 14755 29884 14795 29924
rect 14860 29884 14900 29924
rect 15134 29884 15174 29924
rect 15436 29875 15476 29915
rect 16387 29884 16427 29924
rect 16684 29884 16724 29924
rect 17155 29884 17195 29924
rect 17260 29884 17300 29924
rect 17644 29884 17684 29924
rect 18220 29875 18260 29915
rect 18700 29875 18740 29915
rect 19075 29884 19115 29924
rect 19386 29884 19426 29924
rect 7276 29800 7316 29840
rect 8620 29800 8660 29840
rect 10252 29800 10292 29840
rect 11443 29800 11483 29840
rect 11788 29800 11828 29840
rect 12268 29800 12308 29840
rect 13795 29800 13835 29840
rect 14275 29800 14315 29840
rect 15820 29800 15860 29840
rect 16204 29800 16244 29840
rect 17740 29800 17780 29840
rect 19756 29800 19796 29840
rect 20140 29800 20180 29840
rect 8476 29716 8516 29756
rect 2860 29632 2900 29672
rect 4636 29632 4676 29672
rect 9004 29632 9044 29672
rect 11548 29632 11588 29672
rect 12508 29632 12548 29672
rect 13180 29632 13220 29672
rect 13507 29632 13547 29672
rect 15139 29632 15179 29672
rect 15580 29632 15620 29672
rect 15964 29632 16004 29672
rect 16684 29632 16724 29672
rect 19372 29632 19412 29672
rect 3688 29464 3728 29504
rect 3770 29464 3810 29504
rect 3852 29464 3892 29504
rect 3934 29464 3974 29504
rect 4016 29464 4056 29504
rect 18808 29464 18848 29504
rect 18890 29464 18930 29504
rect 18972 29464 19012 29504
rect 19054 29464 19094 29504
rect 19136 29464 19176 29504
rect 1468 29296 1508 29336
rect 2236 29296 2276 29336
rect 4444 29296 4484 29336
rect 6316 29296 6356 29336
rect 13516 29296 13556 29336
rect 14476 29296 14516 29336
rect 15196 29296 15236 29336
rect 17740 29296 17780 29336
rect 19852 29296 19892 29336
rect 20380 29296 20420 29336
rect 9244 29212 9284 29252
rect 1228 29128 1268 29168
rect 1612 29128 1652 29168
rect 1996 29128 2036 29168
rect 2787 29128 2827 29168
rect 3283 29119 3323 29159
rect 2668 29044 2708 29084
rect 2885 29044 2925 29084
rect 3157 29044 3197 29084
rect 3388 29086 3428 29126
rect 4684 29128 4724 29168
rect 7276 29128 7316 29168
rect 9004 29128 9044 29168
rect 9388 29128 9428 29168
rect 10348 29128 10388 29168
rect 14668 29128 14708 29168
rect 15436 29128 15476 29168
rect 20140 29128 20180 29168
rect 3628 29044 3668 29084
rect 3907 29044 3947 29084
rect 4876 29044 4916 29084
rect 6124 29044 6164 29084
rect 6787 29044 6827 29084
rect 6892 29044 6932 29084
rect 7372 29044 7412 29084
rect 7852 29044 7892 29084
rect 8371 29044 8411 29084
rect 9859 29044 9899 29084
rect 9964 29044 10004 29084
rect 10444 29044 10484 29084
rect 10924 29044 10964 29084
rect 11412 29044 11452 29084
rect 12076 29044 12116 29084
rect 13324 29044 13364 29084
rect 14179 29044 14219 29084
rect 15724 29077 15764 29117
rect 15835 29044 15875 29084
rect 15953 29044 15993 29084
rect 16300 29044 16340 29084
rect 17548 29044 17588 29084
rect 17918 29044 17958 29084
rect 18124 29044 18164 29084
rect 18220 29044 18260 29084
rect 18412 29044 18452 29084
rect 19660 29044 19700 29084
rect 4012 28960 4052 29000
rect 4348 28960 4388 29000
rect 14284 28960 14324 29000
rect 14490 28960 14530 29000
rect 1852 28876 1892 28916
rect 2572 28876 2612 28916
rect 3052 28876 3092 28916
rect 8524 28876 8564 28916
rect 9628 28876 9668 28916
rect 11596 28876 11636 28916
rect 14908 28876 14948 28916
rect 16108 28876 16148 28916
rect 18019 28876 18059 28916
rect 4928 28708 4968 28748
rect 5010 28708 5050 28748
rect 5092 28708 5132 28748
rect 5174 28708 5214 28748
rect 5256 28708 5296 28748
rect 20048 28708 20088 28748
rect 20130 28708 20170 28748
rect 20212 28708 20252 28748
rect 20294 28708 20334 28748
rect 20376 28708 20416 28748
rect 3619 28540 3659 28580
rect 4204 28540 4244 28580
rect 5212 28540 5252 28580
rect 6796 28540 6836 28580
rect 8812 28540 8852 28580
rect 9244 28540 9284 28580
rect 9628 28540 9668 28580
rect 10396 28540 10436 28580
rect 10540 28540 10580 28580
rect 13996 28540 14036 28580
rect 15820 28540 15860 28580
rect 17452 28540 17492 28580
rect 19084 28540 19124 28580
rect 20035 28540 20075 28580
rect 3998 28456 4038 28496
rect 1516 28372 1556 28412
rect 2764 28363 2804 28403
rect 3287 28372 3327 28412
rect 3532 28372 3572 28412
rect 4300 28363 4340 28403
rect 4588 28372 4628 28412
rect 4805 28372 4845 28412
rect 5356 28372 5396 28412
rect 6604 28363 6644 28403
rect 7075 28372 7115 28412
rect 7180 28372 7220 28412
rect 7564 28372 7604 28412
rect 8140 28363 8180 28403
rect 8620 28363 8660 28403
rect 10732 28363 10772 28403
rect 11980 28372 12020 28412
rect 12556 28372 12596 28412
rect 13804 28363 13844 28403
rect 14380 28372 14420 28412
rect 15628 28363 15668 28403
rect 16012 28372 16052 28412
rect 17260 28363 17300 28403
rect 17644 28372 17684 28412
rect 18892 28363 18932 28403
rect 19372 28363 19412 28403
rect 19471 28352 19511 28392
rect 19948 28372 19988 28412
rect 3427 28288 3467 28328
rect 4492 28288 4532 28328
rect 4707 28288 4747 28328
rect 4972 28288 5012 28328
rect 7660 28288 7700 28328
rect 9004 28288 9044 28328
rect 9388 28288 9428 28328
rect 9772 28288 9812 28328
rect 10156 28288 10196 28328
rect 19601 28330 19641 28370
rect 20236 28372 20276 28412
rect 12364 28288 12404 28328
rect 2956 28204 2996 28244
rect 10012 28204 10052 28244
rect 4003 28120 4043 28160
rect 12124 28120 12164 28160
rect 19756 28120 19796 28160
rect 3688 27952 3728 27992
rect 3770 27952 3810 27992
rect 3852 27952 3892 27992
rect 3934 27952 3974 27992
rect 4016 27952 4056 27992
rect 18808 27952 18848 27992
rect 18890 27952 18930 27992
rect 18972 27952 19012 27992
rect 19054 27952 19094 27992
rect 19136 27952 19176 27992
rect 1468 27784 1508 27824
rect 3052 27784 3092 27824
rect 7564 27784 7604 27824
rect 11020 27784 11060 27824
rect 14572 27784 14612 27824
rect 16492 27784 16532 27824
rect 19852 27784 19892 27824
rect 4300 27700 4340 27740
rect 11212 27700 11252 27740
rect 1228 27616 1268 27656
rect 5059 27616 5099 27656
rect 5260 27616 5300 27656
rect 5539 27616 5579 27656
rect 5740 27616 5780 27656
rect 1612 27532 1652 27572
rect 2860 27532 2900 27572
rect 3244 27532 3284 27572
rect 3628 27532 3668 27572
rect 3907 27532 3947 27572
rect 4483 27532 4523 27572
rect 4919 27532 4959 27572
rect 5164 27532 5204 27572
rect 5419 27532 5459 27572
rect 5644 27532 5684 27572
rect 6124 27532 6164 27572
rect 7372 27532 7412 27572
rect 7948 27532 7988 27572
rect 9196 27532 9236 27572
rect 9580 27532 9620 27572
rect 10836 27532 10876 27572
rect 11404 27532 11444 27572
rect 12652 27532 12692 27572
rect 13132 27532 13172 27572
rect 14380 27532 14420 27572
rect 15052 27532 15092 27572
rect 16300 27532 16340 27572
rect 16780 27532 16820 27572
rect 18028 27532 18068 27572
rect 18412 27532 18452 27572
rect 19660 27532 19700 27572
rect 19991 27532 20031 27572
rect 20131 27532 20171 27572
rect 20236 27532 20276 27572
rect 4012 27448 4052 27488
rect 4794 27448 4834 27488
rect 19852 27448 19892 27488
rect 3388 27364 3428 27404
rect 4579 27364 4619 27404
rect 4684 27364 4724 27404
rect 7756 27364 7796 27404
rect 16492 27364 16532 27404
rect 18220 27364 18260 27404
rect 20323 27364 20363 27404
rect 4928 27196 4968 27236
rect 5010 27196 5050 27236
rect 5092 27196 5132 27236
rect 5174 27196 5214 27236
rect 5256 27196 5296 27236
rect 20048 27196 20088 27236
rect 20130 27196 20170 27236
rect 20212 27196 20252 27236
rect 20294 27196 20334 27236
rect 20376 27196 20416 27236
rect 2956 27028 2996 27068
rect 7468 27028 7508 27068
rect 7900 27028 7940 27068
rect 10588 27028 10628 27068
rect 11260 27028 11300 27068
rect 20140 27028 20180 27068
rect 3916 26944 3956 26984
rect 17884 26944 17924 26984
rect 1516 26860 1556 26900
rect 2764 26851 2804 26891
rect 3148 26860 3188 26900
rect 3532 26860 3572 26900
rect 3811 26860 3851 26900
rect 4396 26860 4436 26900
rect 5644 26851 5684 26891
rect 6028 26860 6068 26900
rect 7276 26851 7316 26891
rect 8227 26860 8267 26900
rect 8332 26860 8372 26900
rect 8716 26860 8756 26900
rect 9292 26851 9332 26891
rect 9772 26851 9812 26891
rect 10003 26860 10043 26900
rect 11596 26851 11636 26891
rect 12844 26860 12884 26900
rect 13612 26860 13652 26900
rect 14860 26851 14900 26891
rect 15244 26860 15284 26900
rect 16492 26851 16532 26891
rect 16823 26860 16863 26900
rect 17068 26860 17108 26900
rect 18403 26860 18443 26900
rect 18508 26860 18548 26900
rect 18892 26860 18932 26900
rect 19468 26851 19508 26891
rect 19948 26851 19988 26891
rect 7660 26776 7700 26816
rect 8812 26776 8852 26816
rect 10156 26776 10196 26816
rect 10828 26776 10868 26816
rect 11020 26776 11060 26816
rect 13036 26776 13076 26816
rect 16963 26776 17003 26816
rect 17164 26776 17204 26816
rect 17740 26776 17780 26816
rect 18124 26776 18164 26816
rect 18988 26776 19028 26816
rect 10396 26692 10436 26732
rect 3292 26608 3332 26648
rect 4204 26608 4244 26648
rect 5836 26608 5876 26648
rect 11404 26608 11444 26648
rect 13276 26608 13316 26648
rect 15052 26608 15092 26648
rect 16684 26608 16724 26648
rect 17500 26608 17540 26648
rect 3688 26440 3728 26480
rect 3770 26440 3810 26480
rect 3852 26440 3892 26480
rect 3934 26440 3974 26480
rect 4016 26440 4056 26480
rect 18808 26440 18848 26480
rect 18890 26440 18930 26480
rect 18972 26440 19012 26480
rect 19054 26440 19094 26480
rect 19136 26440 19176 26480
rect 4588 26272 4628 26312
rect 5020 26272 5060 26312
rect 5308 26272 5348 26312
rect 7276 26272 7316 26312
rect 9331 26272 9371 26312
rect 13948 26272 13988 26312
rect 20236 26272 20276 26312
rect 15004 26188 15044 26228
rect 3427 26104 3467 26144
rect 4780 26104 4820 26144
rect 5548 26104 5588 26144
rect 8044 26104 8084 26144
rect 10060 26104 10100 26144
rect 11347 26104 11387 26144
rect 11692 26104 11732 26144
rect 11932 26104 11972 26144
rect 13708 26104 13748 26144
rect 14284 26104 14324 26144
rect 14764 26104 14804 26144
rect 15724 26104 15764 26144
rect 1420 26020 1460 26060
rect 2668 26020 2708 26060
rect 3052 26020 3092 26060
rect 3287 26020 3327 26060
rect 3532 26020 3572 26060
rect 3806 26020 3846 26060
rect 4110 26020 4150 26060
rect 4289 26020 4329 26060
rect 4396 26020 4436 26060
rect 5836 26020 5876 26060
rect 7084 26020 7124 26060
rect 7555 26020 7595 26060
rect 7660 26020 7700 26060
rect 8140 26020 8180 26060
rect 8623 26020 8663 26060
rect 9139 26020 9179 26060
rect 9571 26020 9611 26060
rect 9676 26020 9716 26060
rect 10156 26020 10196 26060
rect 10636 26020 10676 26060
rect 11155 26020 11195 26060
rect 12268 26020 12308 26060
rect 13516 26020 13556 26060
rect 15214 26020 15254 26060
rect 15338 26020 15378 26060
rect 15820 26020 15860 26060
rect 16300 26020 16340 26060
rect 16788 26020 16828 26060
rect 17356 26020 17396 26060
rect 18604 26020 18644 26060
rect 18796 26020 18836 26060
rect 20044 26020 20084 26060
rect 3196 25936 3236 25976
rect 4602 25936 4642 25976
rect 12076 25936 12116 25976
rect 14044 25936 14084 25976
rect 17164 25936 17204 25976
rect 2860 25852 2900 25892
rect 3619 25852 3659 25892
rect 3907 25852 3947 25892
rect 4012 25852 4052 25892
rect 16972 25852 17012 25892
rect 4928 25684 4968 25724
rect 5010 25684 5050 25724
rect 5092 25684 5132 25724
rect 5174 25684 5214 25724
rect 5256 25684 5296 25724
rect 20048 25684 20088 25724
rect 20130 25684 20170 25724
rect 20212 25684 20252 25724
rect 20294 25684 20334 25724
rect 20376 25684 20416 25724
rect 3340 25516 3380 25556
rect 5212 25516 5252 25556
rect 9100 25516 9140 25556
rect 11116 25516 11156 25556
rect 11404 25516 11444 25556
rect 20380 25516 20420 25556
rect 1468 25432 1508 25472
rect 3772 25432 3812 25472
rect 4156 25432 4196 25472
rect 15916 25432 15956 25472
rect 19996 25432 20036 25472
rect 1900 25348 1940 25388
rect 3148 25339 3188 25379
rect 5356 25348 5396 25388
rect 6604 25339 6644 25379
rect 7660 25348 7700 25388
rect 8908 25339 8948 25379
rect 9358 25348 9398 25388
rect 9481 25348 9521 25388
rect 9861 25348 9901 25388
rect 9964 25348 10004 25388
rect 10444 25339 10484 25379
rect 10924 25339 10964 25379
rect 11596 25339 11636 25379
rect 12844 25348 12884 25388
rect 14188 25348 14228 25388
rect 14476 25348 14516 25388
rect 15724 25339 15764 25379
rect 16195 25348 16235 25388
rect 16300 25348 16340 25388
rect 16684 25348 16724 25388
rect 17260 25339 17300 25379
rect 17740 25339 17780 25379
rect 18124 25348 18164 25388
rect 19372 25339 19412 25379
rect 1228 25264 1268 25304
rect 3532 25264 3572 25304
rect 3916 25264 3956 25304
rect 4588 25264 4628 25304
rect 4972 25264 5012 25304
rect 5212 25264 5252 25304
rect 7180 25264 7220 25304
rect 13804 25264 13844 25304
rect 16780 25264 16820 25304
rect 19756 25264 19796 25304
rect 20140 25264 20180 25304
rect 6940 25180 6980 25220
rect 17980 25180 18020 25220
rect 4348 25096 4388 25136
rect 6796 25096 6836 25136
rect 13564 25096 13604 25136
rect 14332 25096 14372 25136
rect 19564 25096 19604 25136
rect 3688 24928 3728 24968
rect 3770 24928 3810 24968
rect 3852 24928 3892 24968
rect 3934 24928 3974 24968
rect 4016 24928 4056 24968
rect 18808 24928 18848 24968
rect 18890 24928 18930 24968
rect 18972 24928 19012 24968
rect 19054 24928 19094 24968
rect 19136 24928 19176 24968
rect 5212 24760 5252 24800
rect 5980 24760 6020 24800
rect 9724 24760 9764 24800
rect 11308 24760 11348 24800
rect 15196 24760 15236 24800
rect 19228 24760 19268 24800
rect 19996 24760 20036 24800
rect 20380 24760 20420 24800
rect 2764 24676 2804 24716
rect 5308 24676 5348 24716
rect 8956 24676 8996 24716
rect 9340 24676 9380 24716
rect 14764 24676 14804 24716
rect 16780 24676 16820 24716
rect 3532 24592 3572 24632
rect 4972 24592 5012 24632
rect 5548 24592 5588 24632
rect 5740 24592 5780 24632
rect 6892 24592 6932 24632
rect 8179 24592 8219 24632
rect 8332 24592 8372 24632
rect 8572 24592 8612 24632
rect 8716 24592 8756 24632
rect 9100 24592 9140 24632
rect 9484 24592 9524 24632
rect 14956 24592 14996 24632
rect 17548 24592 17588 24632
rect 18988 24592 19028 24632
rect 19372 24592 19412 24632
rect 19612 24592 19652 24632
rect 19756 24592 19796 24632
rect 20140 24592 20180 24632
rect 1324 24508 1364 24548
rect 2572 24508 2612 24548
rect 3043 24508 3083 24548
rect 3148 24508 3188 24548
rect 3628 24508 3668 24548
rect 4108 24508 4148 24548
rect 4596 24508 4636 24548
rect 6403 24508 6443 24548
rect 6508 24508 6548 24548
rect 6988 24508 7028 24548
rect 7468 24508 7508 24548
rect 7956 24508 7996 24548
rect 9868 24508 9908 24548
rect 11116 24508 11156 24548
rect 11500 24508 11540 24548
rect 12748 24508 12788 24548
rect 13324 24508 13364 24548
rect 14572 24508 14612 24548
rect 15340 24508 15380 24548
rect 16588 24508 16628 24548
rect 17059 24508 17099 24548
rect 17164 24508 17204 24548
rect 17644 24508 17684 24548
rect 18124 24508 18164 24548
rect 18604 24541 18644 24581
rect 4780 24340 4820 24380
rect 12940 24340 12980 24380
rect 18796 24340 18836 24380
rect 4928 24172 4968 24212
rect 5010 24172 5050 24212
rect 5092 24172 5132 24212
rect 5174 24172 5214 24212
rect 5256 24172 5296 24212
rect 20048 24172 20088 24212
rect 20130 24172 20170 24212
rect 20212 24172 20252 24212
rect 20294 24172 20334 24212
rect 20376 24172 20416 24212
rect 4780 24004 4820 24044
rect 7468 24004 7508 24044
rect 9292 24004 9332 24044
rect 9724 24004 9764 24044
rect 15724 24004 15764 24044
rect 16732 24004 16772 24044
rect 17500 24004 17540 24044
rect 19555 24004 19595 24044
rect 2764 23920 2804 23960
rect 9820 23920 9860 23960
rect 11980 23920 12020 23960
rect 18844 23920 18884 23960
rect 19267 23920 19307 23960
rect 19767 23920 19807 23960
rect 20140 23920 20180 23960
rect 1324 23836 1364 23876
rect 2572 23827 2612 23867
rect 3043 23836 3083 23876
rect 3148 23836 3188 23876
rect 3532 23836 3572 23876
rect 4108 23827 4148 23867
rect 4588 23827 4628 23867
rect 6028 23836 6068 23876
rect 7276 23827 7316 23867
rect 7852 23836 7892 23876
rect 9100 23827 9140 23867
rect 10540 23836 10580 23876
rect 11788 23827 11828 23867
rect 12172 23836 12212 23876
rect 13420 23827 13460 23867
rect 13987 23836 14027 23876
rect 14092 23836 14132 23876
rect 14476 23836 14516 23876
rect 15052 23827 15092 23867
rect 15532 23827 15572 23867
rect 18955 23836 18995 23876
rect 19178 23836 19218 23876
rect 19459 23836 19499 23876
rect 19934 23836 19974 23876
rect 20236 23827 20276 23867
rect 3628 23752 3668 23792
rect 4972 23752 5012 23792
rect 5356 23752 5396 23792
rect 9484 23752 9524 23792
rect 10060 23752 10100 23792
rect 14572 23752 14612 23792
rect 16108 23752 16148 23792
rect 16492 23752 16532 23792
rect 16876 23752 16916 23792
rect 17260 23752 17300 23792
rect 17836 23752 17876 23792
rect 17980 23752 18020 23792
rect 18220 23752 18260 23792
rect 18604 23752 18644 23792
rect 19075 23752 19115 23792
rect 5212 23584 5252 23624
rect 5596 23584 5636 23624
rect 13612 23584 13652 23624
rect 15868 23584 15908 23624
rect 17116 23584 17156 23624
rect 17596 23584 17636 23624
rect 19756 23584 19796 23624
rect 19939 23584 19979 23624
rect 3688 23416 3728 23456
rect 3770 23416 3810 23456
rect 3852 23416 3892 23456
rect 3934 23416 3974 23456
rect 4016 23416 4056 23456
rect 18808 23416 18848 23456
rect 18890 23416 18930 23456
rect 18972 23416 19012 23456
rect 19054 23416 19094 23456
rect 19136 23416 19176 23456
rect 3340 23248 3380 23288
rect 4156 23248 4196 23288
rect 10483 23248 10523 23288
rect 10972 23248 11012 23288
rect 11644 23248 11684 23288
rect 15571 23248 15611 23288
rect 17683 23248 17723 23288
rect 18460 23248 18500 23288
rect 1468 23164 1508 23204
rect 3715 23164 3755 23204
rect 4540 23164 4580 23204
rect 10876 23164 10916 23204
rect 20188 23164 20228 23204
rect 1228 23080 1268 23120
rect 3916 23080 3956 23120
rect 4300 23080 4340 23120
rect 7180 23080 7220 23120
rect 9196 23080 9236 23120
rect 10636 23080 10676 23120
rect 11212 23080 11252 23120
rect 11884 23080 11924 23120
rect 14284 23080 14324 23120
rect 16396 23080 16436 23120
rect 17788 23080 17828 23120
rect 18028 23080 18068 23120
rect 18220 23080 18260 23120
rect 1900 22996 1940 23036
rect 3148 22996 3188 23036
rect 3532 22996 3572 23036
rect 3715 22996 3755 23036
rect 4684 22996 4724 23036
rect 5932 22996 5972 23036
rect 6691 22996 6731 23036
rect 6796 22996 6836 23036
rect 7276 22996 7316 23036
rect 7756 22996 7796 23036
rect 8244 22996 8284 23036
rect 8707 22996 8747 23036
rect 8812 22996 8852 23036
rect 9292 22996 9332 23036
rect 9772 22996 9812 23036
rect 10291 22996 10331 23036
rect 12076 22996 12116 23036
rect 13324 22996 13364 23036
rect 13795 22996 13835 23036
rect 13900 22996 13940 23036
rect 14380 22996 14420 23036
rect 14860 22996 14900 23036
rect 15348 22996 15388 23036
rect 15907 22996 15947 23036
rect 16012 22996 16052 23036
rect 16492 22996 16532 23036
rect 16972 22996 17012 23036
rect 17491 22996 17531 23036
rect 18604 22996 18644 23036
rect 19852 22996 19892 23036
rect 20332 22996 20372 23036
rect 6124 22912 6164 22952
rect 8428 22828 8468 22868
rect 13516 22828 13556 22868
rect 20044 22828 20084 22868
rect 4928 22660 4968 22700
rect 5010 22660 5050 22700
rect 5092 22660 5132 22700
rect 5174 22660 5214 22700
rect 5256 22660 5296 22700
rect 20048 22660 20088 22700
rect 20130 22660 20170 22700
rect 20212 22660 20252 22700
rect 20294 22660 20334 22700
rect 20376 22660 20416 22700
rect 5356 22492 5396 22532
rect 5788 22492 5828 22532
rect 8044 22492 8084 22532
rect 10828 22492 10868 22532
rect 14659 22492 14699 22532
rect 16492 22492 16532 22532
rect 18124 22492 18164 22532
rect 18787 22492 18827 22532
rect 19267 22492 19307 22532
rect 19747 22492 19787 22532
rect 20140 22492 20180 22532
rect 3340 22408 3380 22448
rect 8332 22408 8372 22448
rect 8995 22408 9035 22448
rect 13795 22408 13835 22448
rect 14467 22399 14507 22439
rect 1900 22324 1940 22364
rect 3148 22315 3188 22355
rect 3619 22324 3659 22364
rect 3724 22324 3764 22364
rect 4108 22324 4148 22364
rect 4684 22315 4724 22355
rect 5164 22315 5204 22355
rect 6028 22315 6068 22355
rect 6127 22304 6167 22344
rect 6259 22315 6299 22355
rect 6604 22324 6644 22364
rect 7852 22315 7892 22355
rect 8227 22324 8267 22364
rect 8535 22324 8575 22364
rect 8663 22324 8703 22364
rect 8908 22324 8948 22364
rect 9388 22324 9428 22364
rect 10636 22315 10676 22355
rect 11692 22324 11732 22364
rect 12940 22315 12980 22355
rect 13708 22324 13748 22364
rect 13891 22324 13931 22364
rect 13996 22324 14036 22364
rect 14179 22324 14219 22364
rect 14284 22315 14324 22355
rect 14571 22324 14611 22364
rect 14689 22313 14729 22353
rect 15052 22324 15092 22364
rect 16300 22315 16340 22355
rect 16684 22324 16724 22364
rect 17932 22315 17972 22355
rect 18475 22324 18515 22364
rect 18700 22324 18740 22364
rect 18935 22324 18975 22364
rect 19180 22324 19220 22364
rect 19555 22324 19595 22364
rect 19660 22324 19700 22364
rect 1228 22240 1268 22280
rect 4204 22240 4244 22280
rect 5548 22240 5588 22280
rect 8803 22240 8843 22280
rect 19420 22282 19460 22322
rect 19934 22324 19974 22364
rect 20236 22315 20276 22355
rect 11020 22240 11060 22280
rect 18595 22240 18635 22280
rect 19075 22240 19115 22280
rect 6412 22156 6452 22196
rect 13132 22156 13172 22196
rect 1468 22072 1508 22112
rect 8524 22072 8564 22112
rect 11260 22072 11300 22112
rect 19939 22072 19979 22112
rect 3688 21904 3728 21944
rect 3770 21904 3810 21944
rect 3852 21904 3892 21944
rect 3934 21904 3974 21944
rect 4016 21904 4056 21944
rect 18808 21904 18848 21944
rect 18890 21904 18930 21944
rect 18972 21904 19012 21944
rect 19054 21904 19094 21944
rect 19136 21904 19176 21944
rect 1852 21736 1892 21776
rect 4348 21736 4388 21776
rect 5260 21736 5300 21776
rect 6892 21736 6932 21776
rect 9004 21736 9044 21776
rect 18124 21736 18164 21776
rect 19372 21736 19412 21776
rect 20332 21736 20372 21776
rect 1228 21568 1268 21608
rect 1612 21568 1652 21608
rect 1996 21568 2036 21608
rect 2956 21568 2996 21608
rect 4588 21568 4628 21608
rect 14803 21559 14843 21599
rect 15340 21568 15380 21608
rect 15619 21568 15659 21608
rect 2467 21484 2507 21524
rect 2572 21484 2612 21524
rect 3052 21484 3092 21524
rect 3532 21484 3572 21524
rect 4020 21484 4060 21524
rect 4243 21484 4283 21524
rect 4963 21484 5003 21524
rect 5260 21484 5300 21524
rect 5452 21484 5492 21524
rect 6700 21484 6740 21524
rect 7372 21484 7412 21524
rect 8620 21484 8660 21524
rect 9196 21484 9236 21524
rect 10404 21484 10444 21524
rect 10828 21484 10868 21524
rect 12076 21484 12116 21524
rect 12460 21484 12500 21524
rect 13708 21484 13748 21524
rect 14092 21484 14132 21524
rect 14234 21484 14274 21524
rect 14667 21484 14707 21524
rect 14908 21484 14948 21524
rect 15013 21484 15053 21524
rect 15139 21484 15179 21524
rect 15244 21484 15284 21524
rect 15479 21484 15519 21524
rect 15724 21484 15764 21524
rect 16300 21484 16340 21524
rect 16684 21484 16724 21524
rect 17932 21484 17972 21524
rect 18412 21484 18452 21524
rect 18700 21484 18740 21524
rect 18979 21484 19019 21524
rect 19660 21484 19700 21524
rect 19915 21484 19955 21524
rect 20035 21484 20075 21524
rect 8812 21400 8852 21440
rect 15811 21400 15851 21440
rect 15998 21400 16038 21440
rect 16204 21400 16244 21440
rect 19084 21400 19124 21440
rect 1468 21316 1508 21356
rect 2236 21316 2276 21356
rect 10636 21316 10676 21356
rect 13900 21316 13940 21356
rect 14380 21316 14420 21356
rect 14572 21316 14612 21356
rect 16099 21316 16139 21356
rect 18268 21316 18308 21356
rect 4928 21148 4968 21188
rect 5010 21148 5050 21188
rect 5092 21148 5132 21188
rect 5174 21148 5214 21188
rect 5256 21148 5296 21188
rect 20048 21148 20088 21188
rect 20130 21148 20170 21188
rect 20212 21148 20252 21188
rect 20294 21148 20334 21188
rect 20376 21148 20416 21188
rect 2668 20980 2708 21020
rect 3484 20980 3524 21020
rect 5356 20980 5396 21020
rect 9100 20980 9140 21020
rect 15148 20980 15188 21020
rect 20380 20980 20420 21020
rect 7084 20896 7124 20936
rect 13516 20896 13556 20936
rect 16252 20896 16292 20936
rect 1228 20812 1268 20852
rect 2476 20803 2516 20843
rect 3916 20812 3956 20852
rect 5164 20803 5204 20843
rect 5644 20812 5684 20852
rect 6892 20803 6932 20843
rect 7363 20812 7403 20852
rect 7468 20812 7508 20852
rect 7852 20812 7892 20852
rect 8428 20803 8468 20843
rect 8908 20803 8948 20843
rect 9379 20812 9419 20852
rect 9484 20812 9524 20852
rect 9868 20812 9908 20852
rect 10444 20803 10484 20843
rect 10924 20803 10964 20843
rect 12076 20812 12116 20852
rect 13708 20812 13748 20852
rect 2860 20728 2900 20768
rect 3244 20728 3284 20768
rect 7948 20728 7988 20768
rect 9964 20728 10004 20768
rect 11155 20728 11195 20768
rect 13328 20770 13368 20810
rect 15628 20812 15668 20852
rect 14960 20770 15000 20810
rect 15757 20812 15797 20852
rect 16012 20812 16052 20852
rect 16684 20812 16724 20852
rect 17932 20803 17972 20843
rect 18508 20812 18548 20852
rect 19756 20803 19796 20843
rect 11500 20728 11540 20768
rect 16492 20728 16532 20768
rect 20140 20728 20180 20768
rect 18124 20644 18164 20684
rect 3100 20560 3140 20600
rect 11260 20560 11300 20600
rect 15340 20560 15380 20600
rect 19948 20560 19988 20600
rect 3688 20392 3728 20432
rect 3770 20392 3810 20432
rect 3852 20392 3892 20432
rect 3934 20392 3974 20432
rect 4016 20392 4056 20432
rect 18808 20392 18848 20432
rect 18890 20392 18930 20432
rect 18972 20392 19012 20432
rect 19054 20392 19094 20432
rect 19136 20392 19176 20432
rect 6604 20224 6644 20264
rect 15916 20224 15956 20264
rect 14044 20140 14084 20180
rect 15436 20140 15476 20180
rect 20188 20140 20228 20180
rect 2860 20056 2900 20096
rect 3100 20056 3140 20096
rect 6988 20056 7028 20096
rect 11116 20056 11156 20096
rect 12403 20056 12443 20096
rect 12748 20056 12788 20096
rect 12940 20056 12980 20096
rect 13180 20056 13220 20096
rect 13804 20056 13844 20096
rect 16396 20056 16436 20096
rect 18796 20056 18836 20096
rect 1228 19972 1268 20012
rect 2484 19972 2524 20012
rect 3532 19972 3572 20012
rect 4780 19972 4820 20012
rect 5164 19972 5204 20012
rect 6412 19972 6452 20012
rect 7276 19972 7316 20012
rect 8524 19972 8564 20012
rect 8908 19972 8948 20012
rect 10156 19972 10196 20012
rect 10627 19972 10667 20012
rect 10732 19972 10772 20012
rect 11212 19972 11252 20012
rect 11692 19972 11732 20012
rect 12180 19972 12220 20012
rect 13516 19972 13556 20012
rect 13660 19972 13700 20012
rect 14135 19972 14175 20012
rect 14275 19972 14315 20012
rect 14380 19972 14420 20012
rect 14764 19972 14804 20012
rect 15043 19972 15083 20012
rect 15619 19972 15659 20012
rect 15930 19972 15970 20012
rect 16588 19972 16628 20012
rect 17836 19972 17876 20012
rect 18307 19972 18347 20012
rect 18412 19972 18452 20012
rect 18892 19972 18932 20012
rect 19371 19972 19411 20012
rect 19891 19972 19931 20012
rect 20332 19972 20372 20012
rect 8716 19888 8756 19928
rect 10348 19888 10388 19928
rect 15148 19888 15188 19928
rect 18028 19888 18068 19928
rect 2668 19804 2708 19844
rect 4972 19804 5012 19844
rect 6748 19804 6788 19844
rect 12508 19804 12548 19844
rect 14467 19804 14507 19844
rect 15715 19804 15755 19844
rect 16156 19804 16196 19844
rect 20044 19804 20084 19844
rect 4928 19636 4968 19676
rect 5010 19636 5050 19676
rect 5092 19636 5132 19676
rect 5174 19636 5214 19676
rect 5256 19636 5296 19676
rect 20048 19636 20088 19676
rect 20130 19636 20170 19676
rect 20212 19636 20252 19676
rect 20294 19636 20334 19676
rect 20376 19636 20416 19676
rect 4780 19468 4820 19508
rect 7372 19468 7412 19508
rect 7900 19468 7940 19508
rect 8668 19468 8708 19508
rect 10108 19468 10148 19508
rect 12268 19468 12308 19508
rect 14236 19468 14276 19508
rect 14668 19468 14708 19508
rect 15244 19468 15284 19508
rect 15964 19468 16004 19508
rect 20140 19468 20180 19508
rect 2764 19384 2804 19424
rect 15148 19384 15188 19424
rect 17932 19384 17972 19424
rect 1324 19300 1364 19340
rect 2572 19291 2612 19331
rect 3043 19300 3083 19340
rect 3148 19300 3188 19340
rect 3532 19300 3572 19340
rect 4108 19291 4148 19331
rect 4588 19291 4628 19331
rect 5635 19300 5675 19340
rect 5740 19300 5780 19340
rect 6700 19291 6740 19331
rect 7180 19291 7220 19331
rect 10828 19300 10868 19340
rect 12076 19291 12116 19331
rect 13996 19300 14036 19340
rect 14380 19300 14420 19340
rect 14572 19300 14612 19340
rect 14755 19300 14795 19340
rect 15043 19300 15083 19340
rect 15354 19300 15394 19340
rect 16492 19300 16532 19340
rect 17740 19291 17780 19331
rect 18403 19300 18443 19340
rect 18508 19300 18548 19340
rect 18892 19300 18932 19340
rect 19468 19291 19508 19331
rect 19948 19291 19988 19331
rect 3628 19216 3668 19256
rect 4972 19216 5012 19256
rect 6124 19216 6164 19256
rect 6259 19216 6299 19256
rect 7756 19216 7796 19256
rect 8140 19216 8180 19256
rect 8524 19216 8564 19256
rect 8908 19216 8948 19256
rect 9100 19216 9140 19256
rect 9676 19216 9716 19256
rect 9868 19216 9908 19256
rect 10444 19216 10484 19256
rect 15676 19216 15716 19256
rect 16300 19216 16340 19256
rect 18988 19216 19028 19256
rect 9340 19132 9380 19172
rect 14140 19132 14180 19172
rect 5212 19048 5252 19088
rect 7516 19048 7556 19088
rect 8284 19048 8324 19088
rect 9436 19048 9476 19088
rect 10204 19048 10244 19088
rect 16060 19048 16100 19088
rect 3688 18880 3728 18920
rect 3770 18880 3810 18920
rect 3852 18880 3892 18920
rect 3934 18880 3974 18920
rect 4016 18880 4056 18920
rect 18808 18880 18848 18920
rect 18890 18880 18930 18920
rect 18972 18880 19012 18920
rect 19054 18880 19094 18920
rect 19136 18880 19176 18920
rect 1468 18712 1508 18752
rect 19948 18712 19988 18752
rect 18124 18628 18164 18668
rect 20380 18628 20420 18668
rect 1228 18544 1268 18584
rect 1612 18544 1652 18584
rect 1996 18544 2036 18584
rect 2956 18544 2996 18584
rect 4243 18544 4283 18584
rect 4588 18544 4628 18584
rect 4780 18544 4820 18584
rect 5164 18544 5204 18584
rect 5404 18544 5444 18584
rect 8044 18544 8084 18584
rect 9331 18544 9371 18584
rect 9676 18544 9716 18584
rect 12940 18544 12980 18584
rect 17740 18544 17780 18584
rect 20140 18544 20180 18584
rect 2446 18460 2486 18500
rect 2572 18460 2612 18500
rect 3052 18460 3092 18500
rect 3532 18460 3572 18500
rect 4020 18460 4060 18500
rect 5740 18460 5780 18500
rect 6988 18460 7028 18500
rect 7555 18460 7595 18500
rect 7660 18460 7700 18500
rect 8140 18460 8180 18500
rect 8623 18460 8663 18500
rect 9108 18460 9148 18500
rect 10732 18460 10772 18500
rect 11980 18460 12020 18500
rect 12451 18460 12491 18500
rect 12556 18460 12596 18500
rect 13036 18460 13076 18500
rect 13516 18460 13556 18500
rect 14004 18460 14044 18500
rect 14380 18460 14420 18500
rect 15628 18460 15668 18500
rect 16012 18460 16052 18500
rect 17260 18460 17300 18500
rect 18124 18460 18164 18500
rect 18316 18460 18356 18500
rect 18508 18460 18548 18500
rect 19756 18460 19796 18500
rect 1852 18376 1892 18416
rect 4348 18376 4388 18416
rect 5020 18376 5060 18416
rect 7180 18376 7220 18416
rect 12172 18376 12212 18416
rect 2236 18292 2276 18332
rect 9436 18292 9476 18332
rect 14188 18292 14228 18332
rect 15820 18292 15860 18332
rect 17452 18292 17492 18332
rect 17980 18292 18020 18332
rect 4928 18124 4968 18164
rect 5010 18124 5050 18164
rect 5092 18124 5132 18164
rect 5174 18124 5214 18164
rect 5256 18124 5296 18164
rect 20048 18124 20088 18164
rect 20130 18124 20170 18164
rect 20212 18124 20252 18164
rect 20294 18124 20334 18164
rect 20376 18124 20416 18164
rect 1468 17956 1508 17996
rect 3052 17956 3092 17996
rect 5164 17956 5204 17996
rect 8140 17956 8180 17996
rect 13324 17956 13364 17996
rect 20380 17956 20420 17996
rect 5692 17872 5732 17912
rect 1612 17788 1652 17828
rect 2860 17779 2900 17819
rect 3427 17788 3467 17828
rect 3532 17788 3572 17828
rect 3916 17788 3956 17828
rect 4492 17779 4532 17819
rect 4972 17779 5012 17819
rect 6700 17788 6740 17828
rect 7948 17779 7988 17819
rect 8419 17788 8459 17828
rect 8524 17788 8564 17828
rect 8908 17788 8948 17828
rect 9484 17779 9524 17819
rect 9964 17779 10004 17819
rect 11884 17788 11924 17828
rect 13132 17779 13172 17819
rect 15139 17788 15179 17828
rect 15244 17788 15284 17828
rect 15724 17788 15764 17828
rect 16204 17779 16244 17819
rect 16684 17779 16724 17819
rect 17539 17788 17579 17828
rect 17644 17788 17684 17828
rect 18028 17788 18068 17828
rect 18604 17779 18644 17819
rect 19084 17779 19124 17819
rect 1228 17704 1268 17744
rect 4012 17704 4052 17744
rect 5356 17704 5396 17744
rect 5932 17704 5972 17744
rect 6124 17704 6164 17744
rect 9004 17704 9044 17744
rect 10195 17704 10235 17744
rect 10636 17704 10676 17744
rect 14380 17704 14420 17744
rect 14860 17704 14900 17744
rect 15628 17704 15668 17744
rect 16915 17704 16955 17744
rect 17260 17704 17300 17744
rect 18124 17704 18164 17744
rect 19660 17704 19700 17744
rect 20140 17704 20180 17744
rect 5596 17536 5636 17576
rect 6364 17536 6404 17576
rect 10396 17536 10436 17576
rect 14140 17536 14180 17576
rect 14620 17536 14660 17576
rect 17020 17536 17060 17576
rect 19315 17536 19355 17576
rect 19420 17536 19460 17576
rect 3688 17368 3728 17408
rect 3770 17368 3810 17408
rect 3852 17368 3892 17408
rect 3934 17368 3974 17408
rect 4016 17368 4056 17408
rect 18808 17368 18848 17408
rect 18890 17368 18930 17408
rect 18972 17368 19012 17408
rect 19054 17368 19094 17408
rect 19136 17368 19176 17408
rect 6508 17200 6548 17240
rect 8140 17200 8180 17240
rect 16972 17200 17012 17240
rect 17308 17200 17348 17240
rect 19180 17200 19220 17240
rect 19612 17200 19652 17240
rect 20380 17200 20420 17240
rect 2668 17116 2708 17156
rect 8284 17116 8324 17156
rect 19996 17116 20036 17156
rect 3532 17032 3572 17072
rect 8524 17032 8564 17072
rect 9484 17032 9524 17072
rect 10771 17032 10811 17072
rect 11116 17032 11156 17072
rect 14092 17032 14132 17072
rect 17548 17032 17588 17072
rect 19372 17032 19412 17072
rect 19756 17032 19796 17072
rect 20140 17032 20180 17072
rect 1228 16948 1268 16988
rect 2476 16948 2516 16988
rect 3043 16948 3083 16988
rect 3148 16948 3188 16988
rect 3628 16948 3668 16988
rect 4108 16948 4148 16988
rect 4596 16948 4636 16988
rect 5068 16948 5108 16988
rect 6316 16948 6356 16988
rect 6700 16948 6740 16988
rect 7948 16948 7988 16988
rect 8995 16948 9035 16988
rect 9100 16948 9140 16988
rect 9580 16948 9620 16988
rect 10060 16948 10100 16988
rect 10579 16948 10619 16988
rect 11500 16948 11540 16988
rect 12748 16948 12788 16988
rect 13603 16948 13643 16988
rect 13708 16948 13748 16988
rect 14188 16948 14228 16988
rect 14668 16948 14708 16988
rect 15187 16948 15227 16988
rect 15532 16948 15572 16988
rect 16780 16948 16820 16988
rect 17740 16948 17780 16988
rect 18988 16948 19028 16988
rect 12940 16864 12980 16904
rect 4780 16780 4820 16820
rect 10876 16780 10916 16820
rect 15340 16780 15380 16820
rect 4928 16612 4968 16652
rect 5010 16612 5050 16652
rect 5092 16612 5132 16652
rect 5174 16612 5214 16652
rect 5256 16612 5296 16652
rect 20048 16612 20088 16652
rect 20130 16612 20170 16652
rect 20212 16612 20252 16652
rect 20294 16612 20334 16652
rect 20376 16612 20416 16652
rect 1468 16444 1508 16484
rect 5452 16444 5492 16484
rect 7132 16444 7172 16484
rect 8908 16444 8948 16484
rect 10636 16444 10676 16484
rect 15052 16444 15092 16484
rect 15244 16444 15284 16484
rect 17116 16444 17156 16484
rect 17884 16444 17924 16484
rect 20140 16444 20180 16484
rect 12652 16360 12692 16400
rect 1708 16276 1748 16316
rect 2956 16267 2996 16307
rect 3715 16276 3755 16316
rect 3820 16276 3860 16316
rect 4204 16276 4244 16316
rect 4780 16267 4820 16307
rect 5260 16267 5300 16307
rect 7468 16276 7508 16316
rect 8716 16267 8756 16307
rect 9196 16276 9236 16316
rect 10444 16267 10484 16307
rect 11212 16276 11252 16316
rect 12460 16267 12500 16307
rect 13315 16276 13355 16316
rect 13420 16276 13460 16316
rect 13804 16276 13844 16316
rect 14380 16267 14420 16307
rect 14860 16267 14900 16307
rect 15436 16267 15476 16307
rect 16684 16276 16724 16316
rect 18403 16276 18443 16316
rect 18508 16276 18548 16316
rect 18892 16276 18932 16316
rect 19468 16267 19508 16307
rect 19948 16267 19988 16307
rect 1228 16192 1268 16232
rect 4300 16192 4340 16232
rect 5836 16192 5876 16232
rect 6220 16192 6260 16232
rect 6412 16192 6452 16232
rect 6892 16192 6932 16232
rect 10828 16192 10868 16232
rect 13900 16192 13940 16232
rect 17356 16192 17396 16232
rect 17740 16192 17780 16232
rect 18124 16192 18164 16232
rect 18988 16192 19028 16232
rect 3148 16108 3188 16148
rect 17500 16108 17540 16148
rect 5596 16024 5636 16064
rect 5980 16024 6020 16064
rect 6652 16024 6692 16064
rect 11068 16024 11108 16064
rect 15091 16024 15131 16064
rect 3688 15856 3728 15896
rect 3770 15856 3810 15896
rect 3852 15856 3892 15896
rect 3934 15856 3974 15896
rect 4016 15856 4056 15896
rect 18808 15856 18848 15896
rect 18890 15856 18930 15896
rect 18972 15856 19012 15896
rect 19054 15856 19094 15896
rect 19136 15856 19176 15896
rect 2764 15688 2804 15728
rect 4684 15688 4724 15728
rect 6652 15688 6692 15728
rect 10732 15688 10772 15728
rect 14572 15688 14612 15728
rect 18124 15688 18164 15728
rect 4492 15604 4532 15644
rect 12460 15604 12500 15644
rect 6508 15520 6548 15560
rect 6892 15520 6932 15560
rect 7180 15520 7220 15560
rect 12652 15520 12692 15560
rect 18892 15520 18932 15560
rect 1324 15436 1364 15476
rect 2572 15436 2612 15476
rect 3052 15436 3092 15476
rect 4300 15436 4340 15476
rect 4876 15436 4916 15476
rect 6124 15436 6164 15476
rect 7660 15436 7700 15476
rect 8908 15436 8948 15476
rect 9292 15436 9332 15476
rect 10540 15436 10580 15476
rect 11020 15436 11060 15476
rect 12268 15436 12308 15476
rect 13132 15436 13172 15476
rect 14380 15436 14420 15476
rect 15052 15436 15092 15476
rect 16300 15436 16340 15476
rect 16684 15436 16724 15476
rect 17932 15436 17972 15476
rect 18403 15436 18443 15476
rect 18508 15436 18548 15476
rect 18988 15436 19028 15476
rect 19468 15436 19508 15476
rect 19987 15436 20027 15476
rect 12892 15352 12932 15392
rect 6268 15268 6308 15308
rect 7420 15268 7460 15308
rect 9100 15268 9140 15308
rect 16492 15268 16532 15308
rect 20140 15268 20180 15308
rect 4928 15100 4968 15140
rect 5010 15100 5050 15140
rect 5092 15100 5132 15140
rect 5174 15100 5214 15140
rect 5256 15100 5296 15140
rect 20048 15100 20088 15140
rect 20130 15100 20170 15140
rect 20212 15100 20252 15140
rect 20294 15100 20334 15140
rect 20376 15100 20416 15140
rect 2860 14932 2900 14972
rect 14572 14932 14612 14972
rect 15292 14932 15332 14972
rect 18268 14932 18308 14972
rect 20140 14932 20180 14972
rect 7756 14848 7796 14888
rect 16099 14848 16139 14888
rect 1420 14764 1460 14804
rect 2668 14755 2708 14795
rect 3052 14764 3092 14804
rect 4300 14755 4340 14795
rect 4684 14764 4724 14804
rect 5932 14755 5972 14795
rect 6316 14764 6356 14804
rect 7564 14755 7604 14795
rect 8419 14764 8459 14804
rect 8524 14764 8564 14804
rect 8908 14764 8948 14804
rect 9484 14755 9524 14795
rect 9964 14755 10004 14795
rect 11020 14764 11060 14804
rect 12268 14755 12308 14795
rect 12835 14764 12875 14804
rect 12940 14764 12980 14804
rect 13324 14764 13364 14804
rect 13900 14755 13940 14795
rect 14380 14755 14420 14795
rect 16291 14764 16331 14804
rect 16780 14755 16820 14795
rect 17260 14764 17300 14804
rect 17740 14764 17780 14804
rect 17853 14784 17893 14824
rect 18700 14764 18740 14804
rect 19948 14755 19988 14795
rect 8140 14680 8180 14720
rect 9004 14680 9044 14720
rect 10636 14680 10676 14720
rect 13420 14680 13460 14720
rect 15532 14680 15572 14720
rect 15916 14680 15956 14720
rect 17356 14680 17396 14720
rect 18508 14680 18548 14720
rect 10204 14596 10244 14636
rect 10876 14596 10916 14636
rect 4492 14512 4532 14552
rect 6124 14512 6164 14552
rect 7900 14512 7940 14552
rect 12460 14512 12500 14552
rect 15676 14512 15716 14552
rect 3688 14344 3728 14384
rect 3770 14344 3810 14384
rect 3852 14344 3892 14384
rect 3934 14344 3974 14384
rect 4016 14344 4056 14384
rect 18808 14344 18848 14384
rect 18890 14344 18930 14384
rect 18972 14344 19012 14384
rect 19054 14344 19094 14384
rect 19136 14344 19176 14384
rect 9436 14176 9476 14216
rect 10012 14176 10052 14216
rect 12364 14176 12404 14216
rect 18508 14176 18548 14216
rect 20236 14176 20276 14216
rect 1852 14092 1892 14132
rect 2236 14092 2276 14132
rect 4732 14092 4772 14132
rect 1228 14008 1268 14048
rect 1612 14008 1652 14048
rect 1996 14008 2036 14048
rect 3052 14008 3092 14048
rect 4492 14008 4532 14048
rect 5068 14008 5108 14048
rect 6028 14008 6068 14048
rect 8044 14008 8084 14048
rect 9331 14008 9371 14048
rect 9676 14008 9716 14048
rect 10252 14008 10292 14048
rect 10540 14008 10580 14048
rect 13612 14008 13652 14048
rect 15628 14008 15668 14048
rect 2563 13924 2603 13964
rect 2668 13924 2708 13964
rect 3148 13924 3188 13964
rect 3628 13924 3668 13964
rect 4116 13924 4156 13964
rect 5539 13924 5579 13964
rect 5644 13924 5684 13964
rect 6124 13924 6164 13964
rect 6604 13924 6644 13964
rect 7092 13924 7132 13964
rect 7555 13924 7595 13964
rect 7660 13924 7700 13964
rect 8140 13924 8180 13964
rect 8620 13924 8660 13964
rect 9108 13924 9148 13964
rect 10924 13924 10964 13964
rect 12172 13924 12212 13964
rect 13123 13924 13163 13964
rect 13228 13924 13268 13964
rect 13708 13924 13748 13964
rect 14188 13924 14228 13964
rect 14676 13924 14716 13964
rect 15139 13924 15179 13964
rect 15244 13924 15284 13964
rect 15724 13924 15764 13964
rect 16204 13924 16244 13964
rect 16723 13924 16763 13964
rect 17068 13924 17108 13964
rect 18316 13924 18356 13964
rect 18796 13924 18836 13964
rect 20044 13924 20084 13964
rect 1468 13840 1508 13880
rect 4828 13840 4868 13880
rect 4300 13756 4340 13796
rect 7276 13756 7316 13796
rect 10780 13756 10820 13796
rect 14860 13756 14900 13796
rect 16876 13756 16916 13796
rect 4928 13588 4968 13628
rect 5010 13588 5050 13628
rect 5092 13588 5132 13628
rect 5174 13588 5214 13628
rect 5256 13588 5296 13628
rect 20048 13588 20088 13628
rect 20130 13588 20170 13628
rect 20212 13588 20252 13628
rect 20294 13588 20334 13628
rect 20376 13588 20416 13628
rect 1468 13420 1508 13460
rect 3052 13420 3092 13460
rect 3580 13420 3620 13460
rect 14380 13420 14420 13460
rect 15484 13420 15524 13460
rect 17356 13420 17396 13460
rect 19852 13420 19892 13460
rect 20092 13420 20132 13460
rect 1612 13252 1652 13292
rect 2860 13243 2900 13283
rect 4108 13252 4148 13292
rect 5356 13243 5396 13283
rect 5836 13252 5876 13292
rect 7084 13243 7124 13283
rect 9580 13252 9620 13292
rect 10828 13243 10868 13283
rect 11212 13252 11252 13292
rect 12460 13243 12500 13283
rect 12940 13252 12980 13292
rect 14188 13243 14228 13283
rect 15916 13252 15956 13292
rect 17164 13243 17204 13283
rect 18115 13252 18155 13292
rect 18220 13252 18260 13292
rect 18604 13252 18644 13292
rect 19180 13243 19220 13283
rect 19660 13243 19700 13283
rect 1228 13168 1268 13208
rect 3244 13168 3284 13208
rect 3820 13168 3860 13208
rect 7948 13168 7988 13208
rect 8332 13168 8372 13208
rect 8716 13168 8756 13208
rect 15724 13168 15764 13208
rect 17740 13168 17780 13208
rect 18700 13168 18740 13208
rect 20332 13168 20372 13208
rect 7276 13084 7316 13124
rect 8092 13084 8132 13124
rect 17500 13084 17540 13124
rect 3484 13000 3524 13040
rect 5548 13000 5588 13040
rect 7708 13000 7748 13040
rect 8476 13000 8516 13040
rect 11020 13000 11060 13040
rect 12652 13000 12692 13040
rect 3688 12832 3728 12872
rect 3770 12832 3810 12872
rect 3852 12832 3892 12872
rect 3934 12832 3974 12872
rect 4016 12832 4056 12872
rect 18808 12832 18848 12872
rect 18890 12832 18930 12872
rect 18972 12832 19012 12872
rect 19054 12832 19094 12872
rect 19136 12832 19176 12872
rect 2236 12664 2276 12704
rect 7228 12664 7268 12704
rect 15244 12664 15284 12704
rect 16876 12664 16916 12704
rect 17404 12664 17444 12704
rect 7612 12580 7652 12620
rect 17020 12580 17060 12620
rect 1228 12496 1268 12536
rect 1612 12496 1652 12536
rect 1996 12496 2036 12536
rect 2956 12496 2996 12536
rect 4396 12496 4436 12536
rect 4636 12496 4676 12536
rect 4876 12496 4916 12536
rect 5116 12496 5156 12536
rect 5836 12496 5876 12536
rect 7123 12496 7163 12536
rect 7468 12496 7508 12536
rect 7852 12496 7892 12536
rect 8428 12496 8468 12536
rect 12364 12496 12404 12536
rect 17260 12496 17300 12536
rect 17644 12496 17684 12536
rect 18412 12496 18452 12536
rect 20332 12496 20372 12536
rect 2467 12412 2507 12452
rect 2572 12412 2612 12452
rect 3052 12412 3092 12452
rect 3532 12412 3572 12452
rect 4020 12412 4060 12452
rect 5347 12412 5387 12452
rect 5452 12412 5492 12452
rect 5932 12412 5972 12452
rect 6412 12412 6452 12452
rect 6904 12412 6944 12452
rect 8620 12412 8660 12452
rect 9868 12412 9908 12452
rect 11854 12412 11894 12452
rect 11977 12412 12017 12452
rect 12460 12412 12500 12452
rect 12940 12412 12980 12452
rect 13428 12412 13468 12452
rect 13804 12412 13844 12452
rect 15052 12412 15092 12452
rect 15436 12412 15476 12452
rect 16684 12412 16724 12452
rect 17902 12412 17942 12452
rect 18028 12412 18068 12452
rect 18508 12412 18548 12452
rect 18988 12412 19028 12452
rect 19476 12412 19516 12452
rect 20092 12328 20132 12368
rect 1468 12244 1508 12284
rect 1852 12244 1892 12284
rect 4204 12244 4244 12284
rect 8188 12244 8228 12284
rect 10060 12244 10100 12284
rect 13612 12244 13652 12284
rect 19660 12244 19700 12284
rect 4928 12076 4968 12116
rect 5010 12076 5050 12116
rect 5092 12076 5132 12116
rect 5174 12076 5214 12116
rect 5256 12076 5296 12116
rect 20048 12076 20088 12116
rect 20130 12076 20170 12116
rect 20212 12076 20252 12116
rect 20294 12076 20334 12116
rect 20376 12076 20416 12116
rect 1180 11908 1220 11948
rect 1564 11908 1604 11948
rect 3628 11908 3668 11948
rect 6508 11908 6548 11948
rect 8428 11908 8468 11948
rect 16444 11908 16484 11948
rect 18316 11908 18356 11948
rect 3772 11824 3812 11864
rect 13132 11824 13172 11864
rect 16348 11824 16388 11864
rect 20092 11824 20132 11864
rect 2188 11740 2228 11780
rect 3440 11731 3480 11771
rect 5068 11740 5108 11780
rect 6316 11731 6356 11771
rect 6988 11740 7028 11780
rect 8236 11731 8276 11771
rect 8707 11740 8747 11780
rect 8812 11740 8852 11780
rect 9196 11740 9236 11780
rect 9772 11731 9812 11771
rect 10252 11731 10292 11771
rect 11692 11740 11732 11780
rect 12940 11731 12980 11771
rect 13411 11740 13451 11780
rect 13516 11740 13556 11780
rect 13900 11740 13940 11780
rect 14476 11731 14516 11771
rect 14956 11731 14996 11771
rect 16876 11740 16916 11780
rect 18124 11731 18164 11771
rect 18508 11740 18548 11780
rect 19756 11731 19796 11771
rect 1420 11656 1460 11696
rect 1804 11656 1844 11696
rect 4012 11656 4052 11696
rect 4492 11656 4532 11696
rect 4876 11656 4916 11696
rect 9292 11656 9332 11696
rect 10483 11656 10523 11696
rect 10828 11656 10868 11696
rect 13996 11656 14036 11696
rect 15187 11656 15227 11696
rect 15532 11656 15572 11696
rect 16108 11656 16148 11696
rect 16684 11656 16724 11696
rect 20332 11656 20372 11696
rect 4252 11572 4292 11612
rect 4636 11572 4676 11612
rect 15292 11572 15332 11612
rect 19948 11572 19988 11612
rect 10588 11488 10628 11528
rect 3688 11320 3728 11360
rect 3770 11320 3810 11360
rect 3852 11320 3892 11360
rect 3934 11320 3974 11360
rect 4016 11320 4056 11360
rect 18808 11320 18848 11360
rect 18890 11320 18930 11360
rect 18972 11320 19012 11360
rect 19054 11320 19094 11360
rect 19136 11320 19176 11360
rect 2668 11152 2708 11192
rect 3484 11152 3524 11192
rect 8044 11152 8084 11192
rect 15052 11152 15092 11192
rect 19372 11152 19412 11192
rect 19708 11152 19748 11192
rect 20092 11152 20132 11192
rect 2812 11068 2852 11108
rect 3052 10984 3092 11024
rect 3244 10984 3284 11024
rect 3820 10984 3860 11024
rect 4012 10984 4052 11024
rect 6604 10984 6644 11024
rect 11980 10984 12020 11024
rect 15916 10984 15956 11024
rect 17203 10984 17243 11024
rect 17548 10984 17588 11024
rect 19948 10984 19988 11024
rect 20332 10984 20372 11024
rect 1228 10900 1268 10940
rect 2476 10900 2516 10940
rect 4396 10900 4436 10940
rect 5644 10900 5684 10940
rect 6115 10900 6155 10940
rect 6220 10900 6260 10940
rect 6700 10900 6740 10940
rect 7180 10900 7220 10940
rect 7699 10900 7739 10940
rect 8236 10900 8276 10940
rect 9484 10900 9524 10940
rect 9772 10900 9812 10940
rect 11020 10900 11060 10940
rect 11491 10900 11531 10940
rect 11596 10900 11636 10940
rect 12076 10900 12116 10940
rect 12556 10900 12596 10940
rect 13044 10900 13084 10940
rect 13612 10900 13652 10940
rect 14860 10900 14900 10940
rect 15427 10900 15467 10940
rect 15532 10900 15572 10940
rect 16012 10900 16052 10940
rect 16492 10900 16532 10940
rect 16980 10900 17020 10940
rect 17932 10900 17972 10940
rect 19180 10900 19220 10940
rect 5836 10816 5876 10856
rect 11212 10816 11252 10856
rect 3580 10732 3620 10772
rect 4252 10732 4292 10772
rect 7852 10732 7892 10772
rect 13228 10732 13268 10772
rect 17308 10732 17348 10772
rect 4928 10564 4968 10604
rect 5010 10564 5050 10604
rect 5092 10564 5132 10604
rect 5174 10564 5214 10604
rect 5256 10564 5296 10604
rect 20048 10564 20088 10604
rect 20130 10564 20170 10604
rect 20212 10564 20252 10604
rect 20294 10564 20334 10604
rect 20376 10564 20416 10604
rect 1180 10396 1220 10436
rect 2236 10396 2276 10436
rect 4588 10396 4628 10436
rect 7948 10396 7988 10436
rect 12172 10396 12212 10436
rect 14188 10396 14228 10436
rect 15820 10396 15860 10436
rect 17644 10396 17684 10436
rect 20092 10396 20132 10436
rect 17923 10312 17963 10352
rect 2830 10228 2870 10268
rect 2947 10261 2987 10301
rect 3340 10228 3380 10268
rect 3916 10219 3956 10259
rect 4396 10219 4436 10259
rect 4780 10228 4820 10268
rect 6028 10219 6068 10259
rect 6508 10228 6548 10268
rect 7756 10219 7796 10259
rect 10732 10228 10772 10268
rect 11980 10219 12020 10259
rect 12451 10228 12491 10268
rect 12556 10228 12596 10268
rect 12940 10228 12980 10268
rect 13516 10219 13556 10259
rect 13996 10219 14036 10259
rect 14380 10228 14420 10268
rect 15628 10219 15668 10259
rect 16204 10228 16244 10268
rect 17452 10219 17492 10259
rect 18115 10228 18155 10268
rect 18604 10219 18644 10259
rect 19084 10228 19124 10268
rect 19564 10228 19604 10268
rect 19677 10209 19717 10249
rect 1420 10144 1460 10184
rect 1900 10144 1940 10184
rect 2140 10144 2180 10184
rect 2476 10144 2516 10184
rect 3436 10144 3476 10184
rect 8332 10144 8372 10184
rect 13036 10144 13076 10184
rect 19180 10144 19220 10184
rect 20332 10144 20372 10184
rect 8092 10060 8132 10100
rect 6220 9976 6260 10016
rect 3688 9808 3728 9848
rect 3770 9808 3810 9848
rect 3852 9808 3892 9848
rect 3934 9808 3974 9848
rect 4016 9808 4056 9848
rect 18808 9808 18848 9848
rect 18890 9808 18930 9848
rect 18972 9808 19012 9848
rect 19054 9808 19094 9848
rect 19136 9808 19176 9848
rect 1180 9640 1220 9680
rect 3484 9640 3524 9680
rect 6076 9640 6116 9680
rect 14227 9640 14267 9680
rect 15292 9640 15332 9680
rect 16876 9640 16916 9680
rect 20092 9640 20132 9680
rect 3340 9556 3380 9596
rect 11164 9556 11204 9596
rect 1420 9472 1460 9512
rect 3724 9472 3764 9512
rect 4684 9472 4724 9512
rect 5971 9472 6011 9512
rect 6316 9472 6356 9512
rect 6892 9472 6932 9512
rect 9772 9472 9812 9512
rect 11059 9472 11099 9512
rect 11404 9472 11444 9512
rect 12940 9472 12980 9512
rect 14572 9472 14612 9512
rect 15052 9472 15092 9512
rect 17260 9472 17300 9512
rect 17644 9472 17684 9512
rect 18412 9472 18452 9512
rect 20332 9472 20372 9512
rect 1900 9388 1940 9428
rect 3148 9388 3188 9428
rect 4195 9388 4235 9428
rect 4300 9388 4340 9428
rect 4780 9388 4820 9428
rect 5260 9388 5300 9428
rect 5779 9388 5819 9428
rect 7564 9388 7604 9428
rect 8812 9388 8852 9428
rect 9283 9388 9323 9428
rect 9388 9388 9428 9428
rect 9868 9388 9908 9428
rect 10348 9388 10388 9428
rect 10836 9388 10876 9428
rect 12451 9388 12491 9428
rect 12556 9388 12596 9428
rect 13036 9388 13076 9428
rect 13516 9388 13556 9428
rect 14035 9388 14075 9428
rect 15436 9388 15476 9428
rect 16684 9388 16724 9428
rect 17923 9388 17963 9428
rect 18028 9388 18068 9428
rect 18508 9388 18548 9428
rect 18988 9388 19028 9428
rect 19507 9388 19547 9428
rect 9004 9304 9044 9344
rect 6652 9220 6692 9260
rect 14332 9220 14372 9260
rect 17020 9220 17060 9260
rect 17404 9220 17444 9260
rect 19660 9220 19700 9260
rect 4928 9052 4968 9092
rect 5010 9052 5050 9092
rect 5092 9052 5132 9092
rect 5174 9052 5214 9092
rect 5256 9052 5296 9092
rect 20048 9052 20088 9092
rect 20130 9052 20170 9092
rect 20212 9052 20252 9092
rect 20294 9052 20334 9092
rect 20376 9052 20416 9092
rect 2668 8884 2708 8924
rect 11884 8884 11924 8924
rect 13996 8884 14036 8924
rect 15292 8884 15332 8924
rect 17548 8884 17588 8924
rect 19180 8884 19220 8924
rect 20092 8884 20132 8924
rect 2812 8800 2852 8840
rect 3772 8800 3812 8840
rect 8188 8800 8228 8840
rect 15100 8800 15140 8840
rect 19708 8800 19748 8840
rect 1228 8716 1268 8756
rect 2476 8707 2516 8747
rect 4291 8716 4331 8756
rect 4396 8716 4436 8756
rect 4780 8716 4820 8756
rect 5356 8707 5396 8747
rect 5836 8707 5876 8747
rect 6307 8716 6347 8756
rect 6412 8716 6452 8756
rect 6796 8716 6836 8756
rect 7372 8707 7412 8747
rect 7852 8707 7892 8747
rect 8620 8716 8660 8756
rect 9868 8707 9908 8747
rect 10444 8716 10484 8756
rect 11692 8707 11732 8747
rect 12259 8716 12299 8756
rect 12364 8716 12404 8756
rect 12748 8716 12788 8756
rect 13324 8707 13364 8747
rect 13804 8707 13844 8747
rect 15811 8716 15851 8756
rect 15916 8716 15956 8756
rect 16300 8716 16340 8756
rect 16876 8707 16916 8747
rect 17356 8707 17396 8747
rect 17740 8716 17780 8756
rect 18988 8707 19028 8747
rect 3052 8632 3092 8672
rect 3244 8632 3284 8672
rect 3484 8632 3524 8672
rect 4012 8632 4052 8672
rect 4876 8632 4916 8672
rect 6067 8632 6107 8672
rect 6892 8632 6932 8672
rect 8083 8632 8123 8672
rect 8428 8632 8468 8672
rect 12844 8632 12884 8672
rect 14860 8632 14900 8672
rect 15532 8632 15572 8672
rect 16396 8632 16436 8672
rect 19324 8632 19364 8672
rect 19564 8632 19604 8672
rect 19948 8632 19988 8672
rect 20332 8632 20372 8672
rect 10060 8464 10100 8504
rect 3688 8296 3728 8336
rect 3770 8296 3810 8336
rect 3852 8296 3892 8336
rect 3934 8296 3974 8336
rect 4016 8296 4056 8336
rect 18808 8296 18848 8336
rect 18890 8296 18930 8336
rect 18972 8296 19012 8336
rect 19054 8296 19094 8336
rect 19136 8296 19176 8336
rect 2860 8128 2900 8168
rect 4492 8128 4532 8168
rect 6220 8128 6260 8168
rect 7948 8128 7988 8168
rect 11788 8128 11828 8168
rect 13804 8128 13844 8168
rect 13996 8128 14036 8168
rect 16156 8128 16196 8168
rect 17740 8128 17780 8168
rect 19948 8128 19988 8168
rect 20092 8044 20132 8084
rect 15916 7960 15956 8000
rect 18124 7960 18164 8000
rect 20332 7960 20372 8000
rect 1420 7876 1460 7916
rect 2668 7876 2708 7916
rect 3052 7876 3092 7916
rect 4300 7876 4340 7916
rect 4780 7876 4820 7916
rect 6028 7876 6068 7916
rect 6508 7876 6548 7916
rect 7756 7876 7796 7916
rect 8620 7876 8660 7916
rect 9868 7876 9908 7916
rect 10348 7876 10388 7916
rect 11596 7876 11636 7916
rect 12364 7876 12404 7916
rect 13612 7876 13652 7916
rect 14188 7876 14228 7916
rect 15436 7876 15476 7916
rect 16300 7876 16340 7916
rect 17548 7876 17588 7916
rect 18508 7876 18548 7916
rect 19756 7876 19796 7916
rect 10060 7708 10100 7748
rect 17884 7708 17924 7748
rect 4928 7540 4968 7580
rect 5010 7540 5050 7580
rect 5092 7540 5132 7580
rect 5174 7540 5214 7580
rect 5256 7540 5296 7580
rect 20048 7540 20088 7580
rect 20130 7540 20170 7580
rect 20212 7540 20252 7580
rect 20294 7540 20334 7580
rect 20376 7540 20416 7580
rect 3820 7372 3860 7412
rect 6700 7372 6740 7412
rect 2380 7204 2420 7244
rect 3628 7195 3668 7235
rect 5260 7204 5300 7244
rect 6508 7195 6548 7235
rect 6988 7204 7028 7244
rect 8236 7195 8276 7235
rect 8707 7204 8747 7244
rect 8812 7204 8852 7244
rect 9196 7204 9236 7244
rect 9772 7195 9812 7235
rect 10252 7195 10292 7235
rect 10636 7204 10676 7244
rect 11884 7195 11924 7235
rect 12844 7204 12884 7244
rect 14092 7195 14132 7235
rect 14668 7195 14708 7235
rect 15916 7204 15956 7244
rect 16300 7195 16340 7235
rect 17548 7204 17588 7244
rect 17932 7195 17972 7235
rect 19180 7204 19220 7244
rect 1180 7120 1220 7160
rect 1420 7120 1460 7160
rect 1804 7120 1844 7160
rect 1948 7120 1988 7160
rect 2188 7120 2228 7160
rect 4204 7120 4244 7160
rect 4588 7120 4628 7160
rect 4972 7120 5012 7160
rect 9292 7120 9332 7160
rect 16099 7120 16139 7160
rect 17731 7120 17771 7160
rect 19660 7120 19700 7160
rect 20332 7120 20372 7160
rect 4348 7036 4388 7076
rect 8428 7036 8468 7076
rect 10492 7036 10532 7076
rect 12076 7036 12116 7076
rect 14284 7036 14324 7076
rect 20092 7036 20132 7076
rect 1564 6952 1604 6992
rect 3964 6952 4004 6992
rect 4732 6952 4772 6992
rect 14476 6952 14516 6992
rect 19420 6952 19460 6992
rect 3688 6784 3728 6824
rect 3770 6784 3810 6824
rect 3852 6784 3892 6824
rect 3934 6784 3974 6824
rect 4016 6784 4056 6824
rect 18808 6784 18848 6824
rect 18890 6784 18930 6824
rect 18972 6784 19012 6824
rect 19054 6784 19094 6824
rect 19136 6784 19176 6824
rect 1180 6616 1220 6656
rect 1564 6616 1604 6656
rect 2812 6616 2852 6656
rect 3196 6616 3236 6656
rect 3916 6616 3956 6656
rect 19756 6616 19796 6656
rect 2332 6532 2372 6572
rect 10300 6532 10340 6572
rect 20092 6532 20132 6572
rect 1420 6448 1460 6488
rect 1804 6448 1844 6488
rect 1996 6448 2036 6488
rect 2572 6448 2612 6488
rect 3052 6448 3092 6488
rect 3436 6448 3476 6488
rect 8908 6448 8948 6488
rect 10540 6448 10580 6488
rect 15052 6448 15092 6488
rect 15916 6448 15956 6488
rect 17203 6448 17243 6488
rect 17548 6448 17588 6488
rect 20332 6448 20372 6488
rect 4108 6364 4148 6404
rect 5356 6364 5396 6404
rect 6508 6364 6548 6404
rect 7756 6364 7796 6404
rect 8419 6364 8459 6404
rect 8524 6364 8564 6404
rect 9004 6364 9044 6404
rect 9487 6364 9527 6404
rect 9972 6364 10012 6404
rect 11116 6364 11156 6404
rect 12364 6364 12404 6404
rect 13228 6364 13268 6404
rect 14476 6364 14516 6404
rect 15406 6364 15446 6404
rect 15532 6364 15572 6404
rect 16012 6364 16052 6404
rect 16492 6364 16532 6404
rect 16980 6364 17020 6404
rect 18316 6364 18356 6404
rect 19564 6364 19604 6404
rect 2236 6280 2276 6320
rect 7948 6196 7988 6236
rect 10156 6196 10196 6236
rect 12556 6196 12596 6236
rect 14668 6196 14708 6236
rect 14812 6196 14852 6236
rect 17308 6196 17348 6236
rect 4928 6028 4968 6068
rect 5010 6028 5050 6068
rect 5092 6028 5132 6068
rect 5174 6028 5214 6068
rect 5256 6028 5296 6068
rect 20048 6028 20088 6068
rect 20130 6028 20170 6068
rect 20212 6028 20252 6068
rect 20294 6028 20334 6068
rect 20376 6028 20416 6068
rect 14668 5860 14708 5900
rect 16300 5860 16340 5900
rect 16492 5860 16532 5900
rect 2332 5776 2372 5816
rect 5260 5692 5300 5732
rect 6508 5683 6548 5723
rect 6892 5692 6932 5732
rect 8140 5683 8180 5723
rect 8524 5692 8564 5732
rect 9772 5683 9812 5723
rect 10915 5692 10955 5732
rect 11020 5692 11060 5732
rect 11404 5692 11444 5732
rect 11980 5683 12020 5723
rect 12460 5683 12500 5723
rect 12931 5692 12971 5732
rect 13036 5692 13076 5732
rect 13420 5692 13460 5732
rect 13996 5683 14036 5723
rect 14476 5683 14516 5723
rect 14860 5692 14900 5732
rect 16108 5683 16148 5723
rect 16684 5683 16724 5723
rect 17932 5692 17972 5732
rect 1180 5608 1220 5648
rect 1420 5608 1460 5648
rect 1804 5608 1844 5648
rect 2188 5608 2228 5648
rect 2572 5608 2612 5648
rect 2764 5608 2804 5648
rect 3340 5608 3380 5648
rect 4300 5608 4340 5648
rect 4684 5608 4724 5648
rect 4924 5608 4964 5648
rect 10348 5608 10388 5648
rect 11500 5608 11540 5648
rect 13516 5608 13556 5648
rect 18940 5608 18980 5648
rect 19180 5608 19220 5648
rect 19564 5608 19604 5648
rect 19948 5608 19988 5648
rect 20332 5608 20372 5648
rect 3004 5524 3044 5564
rect 8332 5524 8372 5564
rect 19708 5524 19748 5564
rect 1564 5440 1604 5480
rect 1948 5440 1988 5480
rect 3100 5440 3140 5480
rect 4540 5440 4580 5480
rect 6700 5440 6740 5480
rect 9964 5440 10004 5480
rect 10108 5440 10148 5480
rect 12691 5440 12731 5480
rect 19324 5440 19364 5480
rect 20092 5440 20132 5480
rect 3688 5272 3728 5312
rect 3770 5272 3810 5312
rect 3852 5272 3892 5312
rect 3934 5272 3974 5312
rect 4016 5272 4056 5312
rect 18808 5272 18848 5312
rect 18890 5272 18930 5312
rect 18972 5272 19012 5312
rect 19054 5272 19094 5312
rect 19136 5272 19176 5312
rect 1180 5104 1220 5144
rect 1564 5104 1604 5144
rect 8044 5104 8084 5144
rect 10540 5104 10580 5144
rect 13084 5104 13124 5144
rect 15868 5104 15908 5144
rect 19324 5104 19364 5144
rect 20092 5104 20132 5144
rect 2332 5020 2372 5060
rect 19708 5020 19748 5060
rect 1420 4936 1460 4976
rect 1804 4936 1844 4976
rect 2188 4936 2228 4976
rect 2572 4936 2612 4976
rect 2956 4936 2996 4976
rect 11308 4936 11348 4976
rect 12595 4936 12635 4976
rect 12940 4936 12980 4976
rect 13324 4936 13364 4976
rect 14476 4936 14516 4976
rect 15763 4936 15803 4976
rect 16108 4936 16148 4976
rect 19564 4936 19604 4976
rect 19948 4936 19988 4976
rect 20332 4936 20372 4976
rect 6604 4852 6644 4892
rect 7852 4852 7892 4892
rect 9100 4852 9140 4892
rect 10348 4852 10388 4892
rect 10819 4852 10859 4892
rect 10924 4852 10964 4892
rect 11404 4852 11444 4892
rect 11884 4852 11924 4892
rect 12372 4852 12412 4892
rect 13987 4852 14027 4892
rect 14092 4852 14132 4892
rect 14572 4852 14612 4892
rect 15052 4852 15092 4892
rect 15571 4852 15611 4892
rect 2716 4768 2756 4808
rect 1948 4684 1988 4724
rect 12700 4684 12740 4724
rect 4928 4516 4968 4556
rect 5010 4516 5050 4556
rect 5092 4516 5132 4556
rect 5174 4516 5214 4556
rect 5256 4516 5296 4556
rect 20048 4516 20088 4556
rect 20130 4516 20170 4556
rect 20212 4516 20252 4556
rect 20294 4516 20334 4556
rect 20376 4516 20416 4556
rect 1180 4264 1220 4304
rect 1564 4264 1604 4304
rect 19708 4264 19748 4304
rect 10924 4180 10964 4220
rect 12172 4171 12212 4211
rect 1420 4096 1460 4136
rect 1804 4096 1844 4136
rect 2188 4096 2228 4136
rect 2572 4096 2612 4136
rect 2764 4096 2804 4136
rect 19948 4096 19988 4136
rect 20332 4096 20372 4136
rect 3004 4012 3044 4052
rect 20092 4012 20132 4052
rect 1948 3928 1988 3968
rect 2332 3928 2372 3968
rect 12364 3928 12404 3968
rect 3688 3760 3728 3800
rect 3770 3760 3810 3800
rect 3852 3760 3892 3800
rect 3934 3760 3974 3800
rect 4016 3760 4056 3800
rect 18808 3760 18848 3800
rect 18890 3760 18930 3800
rect 18972 3760 19012 3800
rect 19054 3760 19094 3800
rect 19136 3760 19176 3800
rect 1180 3592 1220 3632
rect 1564 3592 1604 3632
rect 3772 3592 3812 3632
rect 3388 3508 3428 3548
rect 1420 3424 1460 3464
rect 1804 3424 1844 3464
rect 2188 3424 2228 3464
rect 2380 3424 2420 3464
rect 2956 3424 2996 3464
rect 3148 3424 3188 3464
rect 3532 3424 3572 3464
rect 20332 3424 20372 3464
rect 1948 3256 1988 3296
rect 2620 3256 2660 3296
rect 2716 3172 2756 3212
rect 20092 3172 20132 3212
rect 4928 3004 4968 3044
rect 5010 3004 5050 3044
rect 5092 3004 5132 3044
rect 5174 3004 5214 3044
rect 5256 3004 5296 3044
rect 20048 3004 20088 3044
rect 20130 3004 20170 3044
rect 20212 3004 20252 3044
rect 20294 3004 20334 3044
rect 20376 3004 20416 3044
rect 1180 2836 1220 2876
rect 3868 2836 3908 2876
rect 4252 2836 4292 2876
rect 4636 2836 4676 2876
rect 5788 2836 5828 2876
rect 6172 2836 6212 2876
rect 8476 2836 8516 2876
rect 3484 2752 3524 2792
rect 5020 2752 5060 2792
rect 1420 2584 1460 2624
rect 1708 2584 1748 2624
rect 2092 2584 2132 2624
rect 2572 2584 2612 2624
rect 2812 2584 2852 2624
rect 3244 2584 3284 2624
rect 3628 2584 3668 2624
rect 4012 2584 4052 2624
rect 4396 2584 4436 2624
rect 4780 2584 4820 2624
rect 5164 2584 5204 2624
rect 5548 2584 5588 2624
rect 5932 2584 5972 2624
rect 8236 2584 8276 2624
rect 9196 2584 9236 2624
rect 9580 2584 9620 2624
rect 9964 2584 10004 2624
rect 10348 2584 10388 2624
rect 10732 2584 10772 2624
rect 11116 2584 11156 2624
rect 12844 2584 12884 2624
rect 13228 2584 13268 2624
rect 13612 2584 13652 2624
rect 13996 2584 14036 2624
rect 14380 2584 14420 2624
rect 14764 2584 14804 2624
rect 15148 2584 15188 2624
rect 15532 2584 15572 2624
rect 1948 2500 1988 2540
rect 2332 2416 2372 2456
rect 5404 2416 5444 2456
rect 8956 2416 8996 2456
rect 9340 2416 9380 2456
rect 9724 2416 9764 2456
rect 10108 2416 10148 2456
rect 10492 2416 10532 2456
rect 10876 2416 10916 2456
rect 12604 2416 12644 2456
rect 12988 2416 13028 2456
rect 13372 2416 13412 2456
rect 13756 2416 13796 2456
rect 14140 2416 14180 2456
rect 14524 2416 14564 2456
rect 14908 2416 14948 2456
rect 15292 2416 15332 2456
rect 3688 2248 3728 2288
rect 3770 2248 3810 2288
rect 3852 2248 3892 2288
rect 3934 2248 3974 2288
rect 4016 2248 4056 2288
rect 18808 2248 18848 2288
rect 18890 2248 18930 2288
rect 18972 2248 19012 2288
rect 19054 2248 19094 2288
rect 19136 2248 19176 2288
rect 1948 2080 1988 2120
rect 2812 2080 2852 2120
rect 3868 2080 3908 2120
rect 4252 2080 4292 2120
rect 5020 2080 5060 2120
rect 6172 2080 6212 2120
rect 6556 2080 6596 2120
rect 7036 2080 7076 2120
rect 7708 2080 7748 2120
rect 17404 2080 17444 2120
rect 4348 1996 4388 2036
rect 6940 1996 6980 2036
rect 14716 1996 14756 2036
rect 1324 1912 1364 1952
rect 1708 1912 1748 1952
rect 2092 1912 2132 1952
rect 2476 1912 2516 1952
rect 3052 1912 3092 1952
rect 3244 1912 3284 1952
rect 3628 1912 3668 1952
rect 4012 1912 4052 1952
rect 4588 1912 4628 1952
rect 4780 1912 4820 1952
rect 5164 1912 5204 1952
rect 5548 1912 5588 1952
rect 5932 1912 5972 1952
rect 6316 1912 6356 1952
rect 6700 1912 6740 1952
rect 7276 1912 7316 1952
rect 7468 1912 7508 1952
rect 8236 1912 8276 1952
rect 8620 1912 8660 1952
rect 9004 1912 9044 1952
rect 9388 1912 9428 1952
rect 9772 1912 9812 1952
rect 10156 1912 10196 1952
rect 10540 1912 10580 1952
rect 10924 1912 10964 1952
rect 11500 1912 11540 1952
rect 11884 1912 11924 1952
rect 12268 1912 12308 1952
rect 12652 1912 12692 1952
rect 13036 1912 13076 1952
rect 13420 1912 13460 1952
rect 13804 1912 13844 1952
rect 14188 1912 14228 1952
rect 14572 1912 14612 1952
rect 14956 1912 14996 1952
rect 15340 1912 15380 1952
rect 15724 1912 15764 1952
rect 16108 1912 16148 1952
rect 16492 1912 16532 1952
rect 17644 1912 17684 1952
rect 2716 1744 2756 1784
rect 5404 1744 5444 1784
rect 11164 1744 11204 1784
rect 12412 1744 12452 1784
rect 13564 1744 13604 1784
rect 15484 1744 15524 1784
rect 1564 1660 1604 1700
rect 2332 1660 2372 1700
rect 3484 1660 3524 1700
rect 5788 1660 5828 1700
rect 8476 1660 8516 1700
rect 8860 1660 8900 1700
rect 9244 1660 9284 1700
rect 9628 1660 9668 1700
rect 10012 1660 10052 1700
rect 10396 1660 10436 1700
rect 10780 1660 10820 1700
rect 11260 1660 11300 1700
rect 11644 1660 11684 1700
rect 12028 1660 12068 1700
rect 12796 1660 12836 1700
rect 13180 1660 13220 1700
rect 13948 1660 13988 1700
rect 14332 1660 14372 1700
rect 15100 1660 15140 1700
rect 15868 1660 15908 1700
rect 16252 1660 16292 1700
rect 4928 1492 4968 1532
rect 5010 1492 5050 1532
rect 5092 1492 5132 1532
rect 5174 1492 5214 1532
rect 5256 1492 5296 1532
rect 20048 1492 20088 1532
rect 20130 1492 20170 1532
rect 20212 1492 20252 1532
rect 20294 1492 20334 1532
rect 20376 1492 20416 1532
<< metal2 >>
rect 4919 95236 4928 95276
rect 4968 95236 5010 95276
rect 5050 95236 5092 95276
rect 5132 95236 5174 95276
rect 5214 95236 5256 95276
rect 5296 95236 5305 95276
rect 20039 95236 20048 95276
rect 20088 95236 20130 95276
rect 20170 95236 20212 95276
rect 20252 95236 20294 95276
rect 20334 95236 20376 95276
rect 20416 95236 20425 95276
rect 7315 95068 7324 95108
rect 7364 95068 7700 95108
rect 7660 95024 7700 95068
rect 7948 95068 8468 95108
rect 13507 95068 13516 95108
rect 13556 95068 13748 95108
rect 1555 94984 1564 95024
rect 1604 94984 2572 95024
rect 2612 94984 2621 95024
rect 2707 94984 2716 95024
rect 2756 94984 3340 95024
rect 3380 94984 3389 95024
rect 3475 94984 3484 95024
rect 3524 94984 4204 95024
rect 4244 94984 4253 95024
rect 4579 94984 4588 95024
rect 4628 94984 4636 95024
rect 4676 94984 4759 95024
rect 5011 94984 5020 95024
rect 5060 94984 5644 95024
rect 5684 94984 5693 95024
rect 5779 94984 5788 95024
rect 5828 94984 6412 95024
rect 6452 94984 6461 95024
rect 6931 94984 6940 95024
rect 6980 94984 7564 95024
rect 7604 94984 7613 95024
rect 7660 94984 7852 95024
rect 7892 94984 7901 95024
rect 7948 94940 7988 95068
rect 8428 95024 8468 95068
rect 13708 95024 13748 95068
rect 17740 95068 18548 95108
rect 17740 95024 17780 95068
rect 18508 95024 18548 95068
rect 8083 94984 8092 95024
rect 8132 94984 8332 95024
rect 8372 94984 8381 95024
rect 8428 94984 11308 95024
rect 11348 94984 11357 95024
rect 12739 94984 12748 95024
rect 12788 94984 13652 95024
rect 13708 94984 14420 95024
rect 15619 94984 15628 95024
rect 15668 94984 15676 95024
rect 15716 94984 15799 95024
rect 15907 94984 15916 95024
rect 15956 94984 16060 95024
rect 16100 94984 16109 95024
rect 16195 94984 16204 95024
rect 16244 94984 16828 95024
rect 16868 94984 16877 95024
rect 16972 94984 17212 95024
rect 17252 94984 17261 95024
rect 17347 94984 17356 95024
rect 17396 94984 17780 95024
rect 17836 94984 18364 95024
rect 18404 94984 18413 95024
rect 18508 94984 18748 95024
rect 18788 94984 18797 95024
rect 18988 94984 19900 95024
rect 19940 94984 19949 95024
rect 2860 94900 7988 94940
rect 8236 94900 8716 94940
rect 8756 94900 8765 94940
rect 9091 94900 9100 94940
rect 9140 94900 9149 94940
rect 9475 94900 9484 94940
rect 9524 94900 9533 94940
rect 9859 94900 9868 94940
rect 9908 94900 9917 94940
rect 9964 94900 10252 94940
rect 10292 94900 10301 94940
rect 10627 94900 10636 94940
rect 10676 94900 10685 94940
rect 10732 94900 11020 94940
rect 11060 94900 11069 94940
rect 11203 94900 11212 94940
rect 11252 94900 11261 94940
rect 11971 94900 11980 94940
rect 12020 94900 12029 94940
rect 12163 94900 12172 94940
rect 12212 94900 12884 94940
rect 13123 94900 13132 94940
rect 13172 94900 13556 94940
rect 2860 94856 2900 94900
rect 8236 94856 8276 94900
rect 9100 94856 9140 94900
rect 9484 94856 9524 94900
rect 9868 94856 9908 94900
rect 9964 94856 10004 94900
rect 10636 94856 10676 94900
rect 10732 94856 10772 94900
rect 11212 94856 11252 94900
rect 11980 94856 12020 94900
rect 12844 94856 12884 94900
rect 1193 94816 1324 94856
rect 1364 94816 1373 94856
rect 1577 94816 1708 94856
rect 1748 94816 1757 94856
rect 1961 94816 2092 94856
rect 2132 94816 2141 94856
rect 2345 94816 2476 94856
rect 2516 94816 2525 94856
rect 2851 94816 2860 94856
rect 2900 94816 2909 94856
rect 3113 94816 3244 94856
rect 3284 94816 3293 94856
rect 3497 94816 3628 94856
rect 3668 94816 3677 94856
rect 3881 94816 4012 94856
rect 4052 94816 4061 94856
rect 4265 94816 4396 94856
rect 4436 94816 4445 94856
rect 4771 94816 4780 94856
rect 4820 94816 4829 94856
rect 5155 94816 5164 94856
rect 5204 94816 5213 94856
rect 5417 94816 5548 94856
rect 5588 94816 5597 94856
rect 5801 94816 5932 94856
rect 5972 94816 5981 94856
rect 6185 94816 6316 94856
rect 6356 94816 6365 94856
rect 6569 94816 6700 94856
rect 6740 94816 6749 94856
rect 6953 94816 7084 94856
rect 7124 94816 7133 94856
rect 7459 94816 7468 94856
rect 7508 94816 7517 94856
rect 7564 94816 7852 94856
rect 7892 94816 7901 94856
rect 8227 94816 8236 94856
rect 8276 94816 8285 94856
rect 8611 94816 8620 94856
rect 8660 94816 9140 94856
rect 9187 94816 9196 94856
rect 9236 94816 9524 94856
rect 9571 94816 9580 94856
rect 9620 94816 9908 94856
rect 9955 94816 9964 94856
rect 10004 94816 10013 94856
rect 10147 94816 10156 94856
rect 10196 94816 10676 94856
rect 10723 94816 10732 94856
rect 10772 94816 10781 94856
rect 10915 94816 10924 94856
rect 10964 94816 11252 94856
rect 11299 94816 11308 94856
rect 11348 94816 11404 94856
rect 11444 94816 11479 94856
rect 11587 94816 11596 94856
rect 11636 94816 11884 94856
rect 11924 94816 11933 94856
rect 11980 94816 12076 94856
rect 12116 94816 12125 94856
rect 12172 94816 12652 94856
rect 12692 94816 12701 94856
rect 12835 94816 12844 94856
rect 12884 94816 12893 94856
rect 13411 94816 13420 94856
rect 13460 94816 13469 94856
rect 1939 94732 1948 94772
rect 1988 94732 2956 94772
rect 2996 94732 3005 94772
rect 3091 94732 3100 94772
rect 3140 94732 3724 94772
rect 3764 94732 3773 94772
rect 3859 94732 3868 94772
rect 3908 94732 4492 94772
rect 4532 94732 4541 94772
rect 4780 94688 4820 94816
rect 2323 94648 2332 94688
rect 2372 94648 2900 94688
rect 4243 94648 4252 94688
rect 4292 94648 4532 94688
rect 4780 94648 4916 94688
rect 2860 94604 2900 94648
rect 4492 94604 4532 94648
rect 2860 94564 3148 94604
rect 3188 94564 3197 94604
rect 4492 94564 4780 94604
rect 4820 94564 4829 94604
rect 3679 94480 3688 94520
rect 3728 94480 3770 94520
rect 3810 94480 3852 94520
rect 3892 94480 3934 94520
rect 3974 94480 4016 94520
rect 4056 94480 4065 94520
rect 4876 94436 4916 94648
rect 5164 94436 5204 94816
rect 5395 94732 5404 94772
rect 5444 94732 6028 94772
rect 6068 94732 6077 94772
rect 6163 94732 6172 94772
rect 6212 94732 6796 94772
rect 6836 94732 6845 94772
rect 6547 94648 6556 94688
rect 6596 94648 7180 94688
rect 7220 94648 7229 94688
rect 7468 94520 7508 94816
rect 7564 94772 7604 94816
rect 12172 94772 12212 94816
rect 7555 94732 7564 94772
rect 7604 94732 7613 94772
rect 7699 94732 7708 94772
rect 7748 94732 8140 94772
rect 8180 94732 8189 94772
rect 8851 94732 8860 94772
rect 8900 94732 10292 94772
rect 10387 94732 10396 94772
rect 10436 94732 10732 94772
rect 10772 94732 10781 94772
rect 11417 94732 11500 94772
rect 11540 94732 11548 94772
rect 11588 94732 11597 94772
rect 11779 94732 11788 94772
rect 11828 94732 12212 94772
rect 12307 94732 12316 94772
rect 12356 94732 12364 94772
rect 12404 94732 12487 94772
rect 13075 94732 13084 94772
rect 13124 94732 13228 94772
rect 13268 94732 13277 94772
rect 8345 94648 8428 94688
rect 8468 94648 8476 94688
rect 8516 94648 8525 94688
rect 8803 94648 8812 94688
rect 8852 94648 8956 94688
rect 8996 94648 9005 94688
rect 9331 94648 9340 94688
rect 9380 94648 9388 94688
rect 9428 94648 9511 94688
rect 9715 94648 9724 94688
rect 9764 94648 9772 94688
rect 9812 94648 9895 94688
rect 10252 94604 10292 94732
rect 10483 94648 10492 94688
rect 10532 94648 10540 94688
rect 10580 94648 10663 94688
rect 11155 94648 11164 94688
rect 11204 94648 11212 94688
rect 11252 94648 11335 94688
rect 11513 94648 11596 94688
rect 11636 94648 11644 94688
rect 11684 94648 11693 94688
rect 12163 94648 12172 94688
rect 12212 94648 12412 94688
rect 12452 94648 12461 94688
rect 13027 94648 13036 94688
rect 13076 94648 13180 94688
rect 13220 94648 13229 94688
rect 13420 94604 13460 94816
rect 13516 94772 13556 94900
rect 13612 94856 13652 94984
rect 14380 94856 14420 94984
rect 16972 94940 17012 94984
rect 17836 94940 17876 94984
rect 18988 94940 19028 94984
rect 16387 94900 16396 94940
rect 16436 94900 17012 94940
rect 17155 94900 17164 94940
rect 17204 94900 17876 94940
rect 18115 94900 18124 94940
rect 18164 94900 19028 94940
rect 19372 94900 19948 94940
rect 19988 94900 19997 94940
rect 19372 94856 19412 94900
rect 13603 94816 13612 94856
rect 13652 94816 13661 94856
rect 13708 94816 14188 94856
rect 14228 94816 14237 94856
rect 14371 94816 14380 94856
rect 14420 94816 14429 94856
rect 14947 94816 14956 94856
rect 14996 94816 15005 94856
rect 15907 94816 15916 94856
rect 15956 94816 15965 94856
rect 16217 94816 16300 94856
rect 16340 94816 16348 94856
rect 16388 94816 16397 94856
rect 16483 94816 16492 94856
rect 16532 94816 16684 94856
rect 16724 94816 16733 94856
rect 16937 94816 17068 94856
rect 17108 94816 17117 94856
rect 17321 94816 17452 94856
rect 17492 94816 17501 94856
rect 17635 94816 17644 94856
rect 17684 94816 17836 94856
rect 17876 94816 17885 94856
rect 18089 94816 18220 94856
rect 18260 94816 18269 94856
rect 18473 94816 18604 94856
rect 18644 94816 18653 94856
rect 18787 94816 18796 94856
rect 18836 94816 18988 94856
rect 19028 94816 19037 94856
rect 19363 94816 19372 94856
rect 19412 94816 19421 94856
rect 19625 94816 19756 94856
rect 19796 94816 19805 94856
rect 20131 94816 20140 94856
rect 20180 94816 20189 94856
rect 13708 94772 13748 94816
rect 13516 94732 13748 94772
rect 13843 94732 13852 94772
rect 13892 94732 14324 94772
rect 14371 94732 14380 94772
rect 14420 94732 14620 94772
rect 14660 94732 14669 94772
rect 14284 94688 14324 94732
rect 10252 94564 11788 94604
rect 11828 94564 11837 94604
rect 12451 94564 12460 94604
rect 12500 94564 13460 94604
rect 13516 94648 13948 94688
rect 13988 94648 13997 94688
rect 14284 94648 14572 94688
rect 14612 94648 14621 94688
rect 14707 94648 14716 94688
rect 14756 94648 14764 94688
rect 14804 94648 14887 94688
rect 7468 94480 13420 94520
rect 13460 94480 13469 94520
rect 1612 94396 2668 94436
rect 2708 94396 2717 94436
rect 3436 94396 4916 94436
rect 4972 94396 5204 94436
rect 6124 94396 12980 94436
rect 1612 94184 1652 94396
rect 3436 94352 3476 94396
rect 2227 94312 2236 94352
rect 2276 94312 2380 94352
rect 2420 94312 2429 94352
rect 2611 94312 2620 94352
rect 2660 94312 2764 94352
rect 2804 94312 2813 94352
rect 2995 94312 3004 94352
rect 3044 94312 3476 94352
rect 3523 94312 3532 94352
rect 3572 94312 3580 94352
rect 3620 94312 3703 94352
rect 3955 94312 3964 94352
rect 4004 94312 4108 94352
rect 4148 94312 4157 94352
rect 4291 94312 4300 94352
rect 4340 94312 4348 94352
rect 4388 94312 4471 94352
rect 4675 94312 4684 94352
rect 4724 94312 4732 94352
rect 4772 94312 4855 94352
rect 4972 94268 5012 94396
rect 5107 94312 5116 94352
rect 5156 94312 5356 94352
rect 5396 94312 5405 94352
rect 5827 94312 5836 94352
rect 5876 94312 5884 94352
rect 5924 94312 6007 94352
rect 6124 94268 6164 94396
rect 12940 94352 12980 94396
rect 13516 94352 13556 94648
rect 14956 94604 14996 94816
rect 15916 94772 15956 94816
rect 15916 94732 19660 94772
rect 19700 94732 19709 94772
rect 16003 94648 16012 94688
rect 16052 94648 16444 94688
rect 16484 94648 16493 94688
rect 16579 94648 16588 94688
rect 16628 94648 17596 94688
rect 17636 94648 17645 94688
rect 17740 94648 17980 94688
rect 18020 94648 18029 94688
rect 18115 94648 18124 94688
rect 18164 94648 19132 94688
rect 19172 94648 19181 94688
rect 19276 94648 19516 94688
rect 19556 94648 19565 94688
rect 17740 94604 17780 94648
rect 19276 94604 19316 94648
rect 13891 94564 13900 94604
rect 13940 94564 14996 94604
rect 15331 94564 15340 94604
rect 15380 94564 16492 94604
rect 16532 94564 16541 94604
rect 16771 94564 16780 94604
rect 16820 94564 17780 94604
rect 17827 94564 17836 94604
rect 17876 94564 19316 94604
rect 17260 94480 17452 94520
rect 17492 94480 17501 94520
rect 18211 94480 18220 94520
rect 18260 94480 18604 94520
rect 18644 94480 18653 94520
rect 18799 94480 18808 94520
rect 18848 94480 18890 94520
rect 18930 94480 18972 94520
rect 19012 94480 19054 94520
rect 19094 94480 19136 94520
rect 19176 94480 19185 94520
rect 17260 94436 17300 94480
rect 20140 94436 20180 94816
rect 6211 94312 6220 94352
rect 6260 94312 6268 94352
rect 6308 94312 6391 94352
rect 6595 94312 6604 94352
rect 6644 94312 6652 94352
rect 6692 94312 6775 94352
rect 6979 94312 6988 94352
rect 7028 94312 7036 94352
rect 7076 94312 7159 94352
rect 7363 94312 7372 94352
rect 7412 94312 7420 94352
rect 7460 94312 7543 94352
rect 7747 94312 7756 94352
rect 7796 94312 7804 94352
rect 7844 94312 7927 94352
rect 8515 94312 8524 94352
rect 8564 94312 8572 94352
rect 8612 94312 8695 94352
rect 12940 94312 13556 94352
rect 13900 94396 17300 94436
rect 17731 94396 17740 94436
rect 17780 94396 20180 94436
rect 1843 94228 1852 94268
rect 1892 94228 2188 94268
rect 2228 94228 2237 94268
rect 3379 94228 3388 94268
rect 3428 94228 5012 94268
rect 5443 94228 5452 94268
rect 5492 94228 5500 94268
rect 5540 94228 5623 94268
rect 5836 94228 6164 94268
rect 6508 94228 8188 94268
rect 8228 94228 8237 94268
rect 8899 94228 8908 94268
rect 8948 94228 8957 94268
rect 9667 94228 9676 94268
rect 9716 94228 9725 94268
rect 10435 94228 10444 94268
rect 10484 94228 10493 94268
rect 12931 94228 12940 94268
rect 12980 94228 12989 94268
rect 13699 94228 13708 94268
rect 13748 94228 13757 94268
rect 1097 94144 1228 94184
rect 1268 94144 1277 94184
rect 1603 94144 1612 94184
rect 1652 94144 1661 94184
rect 1987 94144 1996 94184
rect 2036 94144 2045 94184
rect 2371 94144 2380 94184
rect 2420 94144 2429 94184
rect 2633 94144 2764 94184
rect 2804 94144 2813 94184
rect 3017 94144 3148 94184
rect 3188 94144 3197 94184
rect 3811 94144 3820 94184
rect 3860 94144 3869 94184
rect 4195 94144 4204 94184
rect 4244 94144 4253 94184
rect 4457 94144 4588 94184
rect 4628 94144 4637 94184
rect 4841 94144 4972 94184
rect 5012 94144 5021 94184
rect 5225 94144 5356 94184
rect 5396 94144 5405 94184
rect 5609 94144 5740 94184
rect 5780 94144 5789 94184
rect 1459 93892 1468 93932
rect 1508 93892 1940 93932
rect 0 93848 90 93868
rect 0 93808 76 93848
rect 116 93808 125 93848
rect 0 93788 90 93808
rect 1900 93680 1940 93892
rect 1996 93764 2036 94144
rect 2380 94100 2420 94144
rect 2380 94060 2860 94100
rect 2900 94060 2909 94100
rect 3820 93932 3860 94144
rect 4204 94016 4244 94144
rect 5836 94100 5876 94228
rect 6508 94184 6548 94228
rect 8908 94184 8948 94228
rect 9676 94184 9716 94228
rect 10444 94184 10484 94228
rect 12940 94184 12980 94228
rect 13708 94184 13748 94228
rect 5993 94144 6124 94184
rect 6164 94144 6173 94184
rect 6499 94144 6508 94184
rect 6548 94144 6557 94184
rect 6761 94144 6892 94184
rect 6932 94144 6941 94184
rect 7145 94144 7276 94184
rect 7316 94144 7325 94184
rect 7651 94144 7660 94184
rect 7700 94144 7709 94184
rect 7913 94144 8044 94184
rect 8084 94144 8093 94184
rect 8227 94144 8236 94184
rect 8276 94144 8428 94184
rect 8468 94144 8477 94184
rect 8803 94144 8812 94184
rect 8852 94144 8861 94184
rect 8908 94144 9004 94184
rect 9044 94144 9053 94184
rect 9283 94144 9292 94184
rect 9332 94144 9580 94184
rect 9620 94144 9629 94184
rect 9676 94144 9772 94184
rect 9812 94144 9821 94184
rect 10051 94144 10060 94184
rect 10100 94144 10348 94184
rect 10388 94144 10397 94184
rect 10444 94144 10540 94184
rect 10580 94144 10589 94184
rect 10819 94144 10828 94184
rect 10868 94144 11116 94184
rect 11156 94144 11165 94184
rect 12547 94144 12556 94184
rect 12596 94144 12844 94184
rect 12884 94144 12893 94184
rect 12940 94144 13036 94184
rect 13076 94144 13085 94184
rect 13315 94144 13324 94184
rect 13364 94144 13612 94184
rect 13652 94144 13661 94184
rect 13708 94144 13804 94184
rect 13844 94144 13853 94184
rect 7660 94100 7700 94144
rect 4675 94060 4684 94100
rect 4724 94060 5876 94100
rect 7171 94060 7180 94100
rect 7220 94060 7700 94100
rect 8812 94100 8852 94144
rect 13900 94100 13940 94396
rect 16435 94312 16444 94352
rect 16484 94312 19508 94352
rect 14467 94228 14476 94268
rect 14516 94228 14996 94268
rect 15043 94228 15052 94268
rect 15092 94228 16820 94268
rect 17203 94228 17212 94268
rect 17252 94228 19124 94268
rect 14956 94184 14996 94228
rect 16780 94184 16820 94228
rect 19084 94184 19124 94228
rect 19468 94184 19508 94312
rect 14083 94144 14092 94184
rect 14132 94144 14572 94184
rect 14612 94144 14621 94184
rect 14947 94144 14956 94184
rect 14996 94144 15005 94184
rect 15209 94144 15244 94184
rect 15284 94144 15340 94184
rect 15380 94144 15389 94184
rect 16073 94144 16204 94184
rect 16244 94144 16253 94184
rect 16771 94144 16780 94184
rect 16820 94144 16829 94184
rect 16963 94144 16972 94184
rect 17012 94144 17143 94184
rect 17347 94144 17356 94184
rect 17396 94144 17527 94184
rect 17587 94144 17596 94184
rect 17636 94144 17740 94184
rect 17780 94144 17789 94184
rect 17923 94144 17932 94184
rect 17972 94144 17981 94184
rect 18115 94144 18124 94184
rect 18164 94144 18295 94184
rect 18569 94144 18604 94184
rect 18644 94144 18700 94184
rect 18740 94144 18749 94184
rect 18835 94144 18844 94184
rect 18884 94144 18932 94184
rect 19075 94144 19084 94184
rect 19124 94144 19133 94184
rect 19459 94144 19468 94184
rect 19508 94144 19517 94184
rect 19721 94144 19852 94184
rect 19892 94144 19901 94184
rect 20105 94144 20236 94184
rect 20276 94144 20285 94184
rect 17932 94100 17972 94144
rect 18892 94100 18932 94144
rect 8812 94060 9484 94100
rect 9524 94060 9533 94100
rect 11683 94060 11692 94100
rect 11732 94060 13940 94100
rect 14851 94060 14860 94100
rect 14900 94060 17972 94100
rect 18019 94060 18028 94100
rect 18068 94060 18932 94100
rect 4204 93976 8140 94016
rect 8180 93976 8189 94016
rect 9235 93976 9244 94016
rect 9284 93976 9580 94016
rect 9620 93976 9629 94016
rect 9881 93976 9964 94016
rect 10004 93976 10012 94016
rect 10052 93976 10061 94016
rect 10771 93976 10780 94016
rect 10820 93976 11020 94016
rect 11060 93976 11069 94016
rect 12067 93976 12076 94016
rect 12116 93976 13276 94016
rect 13316 93976 13325 94016
rect 13411 93976 13420 94016
rect 13460 93976 17300 94016
rect 18355 93976 18364 94016
rect 18404 93976 18836 94016
rect 17260 93932 17300 93976
rect 3820 93892 7468 93932
rect 7508 93892 7517 93932
rect 7651 93892 7660 93932
rect 7700 93892 9340 93932
rect 9380 93892 9389 93932
rect 10099 93892 10108 93932
rect 10148 93892 10156 93932
rect 10196 93892 10279 93932
rect 10745 93892 10828 93932
rect 10868 93892 10876 93932
rect 10916 93892 10925 93932
rect 12595 93892 12604 93932
rect 12644 93892 12652 93932
rect 12692 93892 12775 93932
rect 12931 93892 12940 93932
rect 12980 93892 13372 93932
rect 13412 93892 13421 93932
rect 13891 93892 13900 93932
rect 13940 93892 14044 93932
rect 14084 93892 14093 93932
rect 14201 93892 14284 93932
rect 14324 93892 14332 93932
rect 14372 93892 14381 93932
rect 14585 93892 14668 93932
rect 14708 93892 14716 93932
rect 14756 93892 14765 93932
rect 15091 93892 15100 93932
rect 15140 93892 15148 93932
rect 15188 93892 15271 93932
rect 16531 93892 16540 93932
rect 16580 93892 16588 93932
rect 16628 93892 16711 93932
rect 17260 93892 17452 93932
rect 17492 93892 17501 93932
rect 17683 93892 17692 93932
rect 17732 93892 17740 93932
rect 17780 93892 17863 93932
rect 18028 93892 18460 93932
rect 18500 93892 18509 93932
rect 18028 93848 18068 93892
rect 18796 93848 18836 93976
rect 18892 93892 19228 93932
rect 19268 93892 19277 93932
rect 19481 93892 19564 93932
rect 19604 93892 19612 93932
rect 19652 93892 19661 93932
rect 19747 93892 19756 93932
rect 19796 93892 19996 93932
rect 20036 93892 20045 93932
rect 2860 93808 8620 93848
rect 8660 93808 8669 93848
rect 14467 93808 14476 93848
rect 14516 93808 17492 93848
rect 17539 93808 17548 93848
rect 17588 93808 18068 93848
rect 18307 93808 18316 93848
rect 18356 93808 18644 93848
rect 18787 93808 18796 93848
rect 18836 93808 18845 93848
rect 2860 93764 2900 93808
rect 17452 93764 17492 93808
rect 18604 93764 18644 93808
rect 18892 93764 18932 93892
rect 1996 93724 2900 93764
rect 4919 93724 4928 93764
rect 4968 93724 5010 93764
rect 5050 93724 5092 93764
rect 5132 93724 5174 93764
rect 5214 93724 5256 93764
rect 5296 93724 5305 93764
rect 7459 93724 7468 93764
rect 7508 93724 12268 93764
rect 12308 93724 12317 93764
rect 14947 93724 14956 93764
rect 14996 93724 15572 93764
rect 16387 93724 16396 93764
rect 16436 93724 17396 93764
rect 17452 93724 18220 93764
rect 18260 93724 18269 93764
rect 18604 93724 18932 93764
rect 18979 93724 18988 93764
rect 19028 93724 19852 93764
rect 19892 93724 19901 93764
rect 20039 93724 20048 93764
rect 20088 93724 20130 93764
rect 20170 93724 20212 93764
rect 20252 93724 20294 93764
rect 20334 93724 20376 93764
rect 20416 93724 20425 93764
rect 15532 93680 15572 93724
rect 17356 93680 17396 93724
rect 67 93640 76 93680
rect 116 93640 212 93680
rect 1900 93640 6028 93680
rect 6068 93640 6077 93680
rect 14563 93640 14572 93680
rect 14612 93640 15436 93680
rect 15476 93640 15485 93680
rect 15532 93640 17300 93680
rect 17356 93640 18316 93680
rect 18356 93640 18365 93680
rect 18412 93640 19948 93680
rect 19988 93640 19997 93680
rect 172 93620 212 93640
rect 172 93596 288 93620
rect 17260 93596 17300 93640
rect 18412 93596 18452 93640
rect 163 93556 172 93596
rect 212 93580 288 93596
rect 212 93556 221 93580
rect 1987 93556 1996 93596
rect 2036 93556 2716 93596
rect 2756 93556 2765 93596
rect 17260 93556 18452 93596
rect 18499 93556 18508 93596
rect 18548 93556 18556 93596
rect 18596 93556 18679 93596
rect 19651 93556 19660 93596
rect 19700 93556 19708 93596
rect 19748 93556 19831 93596
rect 0 93512 90 93532
rect 0 93472 2420 93512
rect 2467 93472 2476 93512
rect 2516 93472 2620 93512
rect 2660 93472 2669 93512
rect 18451 93472 18460 93512
rect 18500 93472 18700 93512
rect 18740 93472 18749 93512
rect 0 93452 90 93472
rect 163 93388 172 93428
rect 212 93388 2132 93428
rect 451 93304 460 93344
rect 500 93304 1228 93344
rect 1268 93304 1277 93344
rect 1481 93304 1612 93344
rect 1652 93304 1661 93344
rect 1987 93304 1996 93344
rect 2036 93304 2045 93344
rect 1996 93260 2036 93304
rect 1324 93220 2036 93260
rect 2092 93260 2132 93388
rect 2380 93344 2420 93472
rect 2860 93388 3188 93428
rect 2860 93344 2900 93388
rect 3148 93344 3188 93388
rect 18220 93388 19756 93428
rect 19796 93388 19805 93428
rect 18220 93344 18260 93388
rect 2371 93304 2380 93344
rect 2420 93304 2429 93344
rect 2476 93304 2900 93344
rect 2947 93304 2956 93344
rect 2996 93304 3005 93344
rect 3139 93304 3148 93344
rect 3188 93304 3197 93344
rect 17827 93304 17836 93344
rect 17876 93304 17885 93344
rect 18211 93304 18220 93344
rect 18260 93304 18269 93344
rect 18665 93304 18796 93344
rect 18836 93304 18845 93344
rect 18979 93304 18988 93344
rect 19028 93304 19159 93344
rect 19555 93304 19564 93344
rect 19604 93304 19948 93344
rect 19988 93304 19997 93344
rect 20131 93304 20140 93344
rect 20180 93304 20311 93344
rect 2476 93260 2516 93304
rect 2092 93220 2516 93260
rect 2956 93260 2996 93304
rect 2956 93220 4780 93260
rect 4820 93220 4829 93260
rect 0 93176 90 93196
rect 0 93136 1228 93176
rect 1268 93136 1277 93176
rect 0 93116 90 93136
rect 0 92840 90 92860
rect 1324 92840 1364 93220
rect 1459 93136 1468 93176
rect 1508 93136 1708 93176
rect 1748 93136 1757 93176
rect 1843 93136 1852 93176
rect 1892 93136 2132 93176
rect 2227 93136 2236 93176
rect 2276 93136 2612 93176
rect 3379 93136 3388 93176
rect 3428 93136 4108 93176
rect 4148 93136 4157 93176
rect 0 92800 1364 92840
rect 0 92780 90 92800
rect 2092 92756 2132 93136
rect 2572 92924 2612 93136
rect 3679 92968 3688 93008
rect 3728 92968 3770 93008
rect 3810 92968 3852 93008
rect 3892 92968 3934 93008
rect 3974 92968 4016 93008
rect 4056 92968 4065 93008
rect 2572 92884 8716 92924
rect 8756 92884 8765 92924
rect 2179 92800 2188 92840
rect 2228 92800 2716 92840
rect 2756 92800 2765 92840
rect 2092 92716 13612 92756
rect 13652 92716 13661 92756
rect 1097 92632 1228 92672
rect 1268 92632 1277 92672
rect 1411 92632 1420 92672
rect 1460 92632 1612 92672
rect 1652 92632 1661 92672
rect 1865 92632 1996 92672
rect 2036 92632 2045 92672
rect 2092 92632 2236 92672
rect 2276 92632 2285 92672
rect 2371 92632 2380 92672
rect 2420 92632 2429 92672
rect 2947 92632 2956 92672
rect 2996 92632 3127 92672
rect 2092 92588 2132 92632
rect 1891 92548 1900 92588
rect 1940 92548 2132 92588
rect 0 92504 90 92524
rect 2380 92504 2420 92632
rect 17836 92504 17876 93304
rect 18067 93220 18076 93260
rect 18116 93220 19084 93260
rect 19124 93220 19133 93260
rect 19219 93220 19228 93260
rect 19268 93220 19564 93260
rect 19604 93220 19613 93260
rect 18691 93136 18700 93176
rect 18740 93136 19324 93176
rect 19364 93136 19373 93176
rect 20371 93136 20380 93176
rect 20420 93136 21004 93176
rect 21044 93136 21053 93176
rect 18799 92968 18808 93008
rect 18848 92968 18890 93008
rect 18930 92968 18972 93008
rect 19012 92968 19054 93008
rect 19094 92968 19136 93008
rect 19176 92968 19185 93008
rect 18931 92800 18940 92840
rect 18980 92800 19276 92840
rect 19316 92800 19325 92840
rect 19459 92800 19468 92840
rect 19508 92800 19517 92840
rect 19468 92756 19508 92800
rect 18835 92716 18844 92756
rect 18884 92716 19508 92756
rect 21510 92672 21600 92692
rect 18595 92632 18604 92672
rect 18644 92632 18653 92672
rect 19049 92632 19180 92672
rect 19220 92632 19229 92672
rect 19433 92632 19468 92672
rect 19508 92632 19564 92672
rect 19604 92632 19613 92672
rect 19747 92632 19756 92672
rect 19796 92632 19927 92672
rect 20131 92632 20140 92672
rect 20180 92632 20524 92672
rect 20564 92632 20573 92672
rect 20995 92632 21004 92672
rect 21044 92632 21600 92672
rect 18604 92588 18644 92632
rect 21510 92612 21600 92632
rect 18604 92548 19660 92588
rect 19700 92548 19709 92588
rect 0 92464 2420 92504
rect 2611 92464 2620 92504
rect 2660 92464 15532 92504
rect 15572 92464 15581 92504
rect 17836 92464 19324 92504
rect 19364 92464 19373 92504
rect 0 92444 90 92464
rect 1459 92380 1468 92420
rect 1508 92380 1517 92420
rect 1843 92380 1852 92420
rect 1892 92380 2132 92420
rect 2659 92380 2668 92420
rect 2708 92380 6796 92420
rect 6836 92380 6845 92420
rect 16003 92380 16012 92420
rect 16052 92380 19180 92420
rect 19220 92380 19229 92420
rect 19987 92380 19996 92420
rect 20036 92380 20045 92420
rect 20371 92380 20380 92420
rect 20420 92380 21004 92420
rect 21044 92380 21053 92420
rect 1468 92252 1508 92380
rect 2092 92336 2132 92380
rect 19996 92336 20036 92380
rect 2092 92296 3148 92336
rect 3188 92296 3197 92336
rect 19996 92296 20852 92336
rect 1468 92212 2956 92252
rect 2996 92212 3005 92252
rect 4919 92212 4928 92252
rect 4968 92212 5010 92252
rect 5050 92212 5092 92252
rect 5132 92212 5174 92252
rect 5214 92212 5256 92252
rect 5296 92212 5305 92252
rect 20039 92212 20048 92252
rect 20088 92212 20130 92252
rect 20170 92212 20212 92252
rect 20252 92212 20294 92252
rect 20334 92212 20376 92252
rect 20416 92212 20425 92252
rect 0 92168 90 92188
rect 20812 92168 20852 92296
rect 21510 92168 21600 92188
rect 0 92128 1612 92168
rect 1652 92128 1661 92168
rect 20812 92128 21600 92168
rect 0 92108 90 92128
rect 21510 92108 21600 92128
rect 5923 92044 5932 92084
rect 5972 92044 7804 92084
rect 7844 92044 7853 92084
rect 19241 92044 19324 92084
rect 19364 92044 19372 92084
rect 19412 92044 19421 92084
rect 1315 91960 1324 92000
rect 1364 91960 2420 92000
rect 1123 91876 1132 91916
rect 1172 91876 2036 91916
rect 0 91832 90 91852
rect 1996 91832 2036 91876
rect 2380 91832 2420 91960
rect 0 91792 460 91832
rect 500 91792 509 91832
rect 739 91792 748 91832
rect 788 91792 1228 91832
rect 1268 91792 1277 91832
rect 1481 91792 1516 91832
rect 1556 91792 1612 91832
rect 1652 91792 1661 91832
rect 1987 91792 1996 91832
rect 2036 91792 2045 91832
rect 2371 91792 2380 91832
rect 2420 91792 2429 91832
rect 2755 91792 2764 91832
rect 2804 91792 2813 91832
rect 7913 91792 8044 91832
rect 8084 91792 8093 91832
rect 19433 91792 19564 91832
rect 19604 91792 19613 91832
rect 19747 91792 19756 91832
rect 19796 91792 19927 91832
rect 20131 91792 20140 91832
rect 20180 91792 20908 91832
rect 20948 91792 20957 91832
rect 0 91772 90 91792
rect 2764 91748 2804 91792
rect 172 91708 2804 91748
rect 0 91496 90 91516
rect 172 91496 212 91708
rect 21510 91664 21600 91684
rect 1459 91624 1468 91664
rect 1508 91624 1517 91664
rect 1603 91624 1612 91664
rect 1652 91624 1852 91664
rect 1892 91624 1901 91664
rect 2105 91624 2188 91664
rect 2228 91624 2236 91664
rect 2276 91624 2285 91664
rect 2467 91624 2476 91664
rect 2516 91624 2620 91664
rect 2660 91624 2669 91664
rect 2995 91624 3004 91664
rect 3044 91624 9676 91664
rect 9716 91624 9725 91664
rect 19987 91624 19996 91664
rect 20036 91624 20045 91664
rect 20371 91624 20380 91664
rect 20420 91624 20812 91664
rect 20852 91624 20861 91664
rect 20995 91624 21004 91664
rect 21044 91624 21600 91664
rect 1468 91580 1508 91624
rect 1468 91540 18508 91580
rect 18548 91540 18557 91580
rect 19996 91496 20036 91624
rect 21510 91604 21600 91624
rect 0 91456 212 91496
rect 3679 91456 3688 91496
rect 3728 91456 3770 91496
rect 3810 91456 3852 91496
rect 3892 91456 3934 91496
rect 3974 91456 4016 91496
rect 4056 91456 4065 91496
rect 18799 91456 18808 91496
rect 18848 91456 18890 91496
rect 18930 91456 18972 91496
rect 19012 91456 19054 91496
rect 19094 91456 19136 91496
rect 19176 91456 19185 91496
rect 19996 91456 21575 91496
rect 0 91436 90 91456
rect 2563 91372 2572 91412
rect 2612 91372 10828 91412
rect 10868 91372 10877 91412
rect 21535 91328 21575 91456
rect 67 91288 76 91328
rect 116 91288 2804 91328
rect 6883 91288 6892 91328
rect 6932 91288 7708 91328
rect 7748 91288 7757 91328
rect 21388 91288 21575 91328
rect 748 91204 1996 91244
rect 2036 91204 2045 91244
rect 0 91160 90 91180
rect 748 91160 788 91204
rect 2764 91160 2804 91288
rect 7267 91204 7276 91244
rect 7316 91204 8092 91244
rect 8132 91204 8141 91244
rect 21388 91160 21428 91288
rect 21510 91160 21600 91180
rect 0 91120 788 91160
rect 835 91120 844 91160
rect 884 91120 1228 91160
rect 1268 91120 1277 91160
rect 1603 91120 1612 91160
rect 1652 91120 1661 91160
rect 1987 91120 1996 91160
rect 2036 91120 2324 91160
rect 2371 91120 2380 91160
rect 2420 91120 2572 91160
rect 2612 91120 2621 91160
rect 2755 91120 2764 91160
rect 2804 91120 2813 91160
rect 7817 91120 7948 91160
rect 7988 91120 7997 91160
rect 8201 91120 8332 91160
rect 8372 91120 8381 91160
rect 19625 91120 19660 91160
rect 19700 91120 19756 91160
rect 19796 91120 19805 91160
rect 20009 91120 20140 91160
rect 20180 91120 20189 91160
rect 21388 91120 21600 91160
rect 0 91100 90 91120
rect 1612 90992 1652 91120
rect 2284 91076 2324 91120
rect 21510 91100 21600 91120
rect 2284 91036 2380 91076
rect 2420 91036 2429 91076
rect 259 90952 268 90992
rect 308 90952 1652 90992
rect 2227 90952 2236 90992
rect 2276 90952 9964 90992
rect 10004 90952 10013 90992
rect 19987 90952 19996 90992
rect 20036 90952 20716 90992
rect 20756 90952 20765 90992
rect 1459 90868 1468 90908
rect 1508 90868 1517 90908
rect 1721 90868 1804 90908
rect 1844 90868 1852 90908
rect 1892 90868 1901 90908
rect 2611 90868 2620 90908
rect 2660 90868 2900 90908
rect 2995 90868 3004 90908
rect 3044 90868 3052 90908
rect 3092 90868 3175 90908
rect 20371 90868 20380 90908
rect 20420 90868 21004 90908
rect 21044 90868 21053 90908
rect 0 90824 90 90844
rect 0 90784 1324 90824
rect 1364 90784 1373 90824
rect 0 90764 90 90784
rect 1468 90740 1508 90868
rect 2860 90824 2900 90868
rect 2860 90784 4684 90824
rect 4724 90784 4733 90824
rect 4780 90784 6028 90824
rect 6068 90784 6077 90824
rect 4780 90740 4820 90784
rect 1468 90700 4820 90740
rect 4919 90700 4928 90740
rect 4968 90700 5010 90740
rect 5050 90700 5092 90740
rect 5132 90700 5174 90740
rect 5214 90700 5256 90740
rect 5296 90700 5305 90740
rect 20039 90700 20048 90740
rect 20088 90700 20130 90740
rect 20170 90700 20212 90740
rect 20252 90700 20294 90740
rect 20334 90700 20376 90740
rect 20416 90700 20425 90740
rect 21510 90656 21600 90676
rect 20803 90616 20812 90656
rect 20852 90616 21600 90656
rect 21510 90596 21600 90616
rect 2380 90532 4492 90572
rect 4532 90532 4541 90572
rect 16937 90532 17020 90572
rect 17060 90532 17068 90572
rect 17108 90532 17117 90572
rect 0 90488 90 90508
rect 0 90448 1420 90488
rect 1460 90448 1469 90488
rect 0 90428 90 90448
rect 2380 90320 2420 90532
rect 2476 90448 14188 90488
rect 14228 90448 14237 90488
rect 643 90280 652 90320
rect 692 90280 1228 90320
rect 1268 90280 1277 90320
rect 1337 90280 1420 90320
rect 1460 90280 1468 90320
rect 1508 90280 1517 90320
rect 1603 90280 1612 90320
rect 1652 90280 1661 90320
rect 1987 90280 1996 90320
rect 2036 90280 2092 90320
rect 2132 90280 2167 90320
rect 2371 90280 2380 90320
rect 2420 90280 2429 90320
rect 1612 90236 1652 90280
rect 2476 90236 2516 90448
rect 2860 90364 3956 90404
rect 11273 90364 11404 90404
rect 11444 90364 11453 90404
rect 12652 90395 13132 90404
rect 2633 90280 2668 90320
rect 2708 90280 2764 90320
rect 2804 90280 2813 90320
rect 2860 90236 2900 90364
rect 3916 90320 3956 90364
rect 12692 90364 13132 90395
rect 13172 90364 13181 90404
rect 14371 90364 14380 90404
rect 14420 90364 15340 90404
rect 15380 90364 15389 90404
rect 15497 90364 15628 90404
rect 15668 90364 15677 90404
rect 12652 90346 12692 90355
rect 15628 90346 15668 90355
rect 3209 90280 3340 90320
rect 3380 90280 3389 90320
rect 3523 90280 3532 90320
rect 3572 90280 3703 90320
rect 3907 90280 3916 90320
rect 3956 90280 3965 90320
rect 17129 90280 17260 90320
rect 17300 90280 17309 90320
rect 19241 90280 19276 90320
rect 19316 90280 19372 90320
rect 19412 90280 19421 90320
rect 19747 90280 19756 90320
rect 19796 90280 19805 90320
rect 20009 90280 20140 90320
rect 20180 90280 20189 90320
rect 19756 90236 19796 90280
rect 1027 90196 1036 90236
rect 1076 90196 1652 90236
rect 1843 90196 1852 90236
rect 1892 90196 2516 90236
rect 2764 90196 2900 90236
rect 2995 90196 3004 90236
rect 3044 90196 11020 90236
rect 11060 90196 11069 90236
rect 11116 90196 19796 90236
rect 20371 90196 20380 90236
rect 20420 90196 21292 90236
rect 21332 90196 21341 90236
rect 0 90152 90 90172
rect 0 90112 1228 90152
rect 1268 90112 1277 90152
rect 2227 90112 2236 90152
rect 2276 90112 2284 90152
rect 2324 90112 2407 90152
rect 2476 90112 2620 90152
rect 2660 90112 2669 90152
rect 0 90092 90 90112
rect 2476 90068 2516 90112
rect 1411 90028 1420 90068
rect 1460 90028 2516 90068
rect 2764 89984 2804 90196
rect 11116 90152 11156 90196
rect 21510 90152 21600 90172
rect 3091 90112 3100 90152
rect 3140 90112 3148 90152
rect 3188 90112 3271 90152
rect 3763 90112 3772 90152
rect 3812 90112 4012 90152
rect 4052 90112 4061 90152
rect 4147 90112 4156 90152
rect 4196 90112 4204 90152
rect 4244 90112 4327 90152
rect 5731 90112 5740 90152
rect 5780 90112 11156 90152
rect 12835 90112 12844 90152
rect 12884 90112 13036 90152
rect 13076 90112 13085 90152
rect 15811 90112 15820 90152
rect 15860 90112 16108 90152
rect 16148 90112 16157 90152
rect 19603 90112 19612 90152
rect 19652 90112 19661 90152
rect 19987 90112 19996 90152
rect 20036 90112 20045 90152
rect 20707 90112 20716 90152
rect 20756 90112 21600 90152
rect 19612 89984 19652 90112
rect 19996 90068 20036 90112
rect 21510 90092 21600 90112
rect 19996 90028 20812 90068
rect 20852 90028 20861 90068
rect 172 89944 2804 89984
rect 3679 89944 3688 89984
rect 3728 89944 3770 89984
rect 3810 89944 3852 89984
rect 3892 89944 3934 89984
rect 3974 89944 4016 89984
rect 4056 89944 4065 89984
rect 18799 89944 18808 89984
rect 18848 89944 18890 89984
rect 18930 89944 18972 89984
rect 19012 89944 19054 89984
rect 19094 89944 19136 89984
rect 19176 89944 19185 89984
rect 19612 89944 21575 89984
rect 0 89816 90 89836
rect 172 89816 212 89944
rect 1315 89860 1324 89900
rect 1364 89860 2668 89900
rect 2708 89860 2717 89900
rect 4012 89860 11596 89900
rect 11636 89860 11645 89900
rect 4012 89816 4052 89860
rect 21535 89816 21575 89944
rect 0 89776 212 89816
rect 2611 89776 2620 89816
rect 2660 89776 3628 89816
rect 3668 89776 3677 89816
rect 3763 89776 3772 89816
rect 3812 89776 4052 89816
rect 4147 89776 4156 89816
rect 4196 89776 11500 89816
rect 11540 89776 11549 89816
rect 21388 89776 21575 89816
rect 0 89756 90 89776
rect 2083 89692 2092 89732
rect 2132 89692 2668 89732
rect 2708 89692 2717 89732
rect 2851 89692 2860 89732
rect 2900 89692 2909 89732
rect 2995 89692 3004 89732
rect 3044 89692 10636 89732
rect 10676 89692 10685 89732
rect 13219 89692 13228 89732
rect 13268 89692 17164 89732
rect 17204 89692 17213 89732
rect 19987 89692 19996 89732
rect 20036 89692 21196 89732
rect 21236 89692 21245 89732
rect 2860 89648 2900 89692
rect 21388 89648 21428 89776
rect 21510 89648 21600 89668
rect 931 89608 940 89648
rect 980 89608 1228 89648
rect 1268 89608 1277 89648
rect 1603 89608 1612 89648
rect 1652 89608 1661 89648
rect 1865 89608 1996 89648
rect 2036 89608 2045 89648
rect 2371 89608 2380 89648
rect 2420 89608 2476 89648
rect 2516 89608 2580 89648
rect 2755 89608 2764 89648
rect 2804 89608 2813 89648
rect 2860 89608 3148 89648
rect 3188 89608 3197 89648
rect 3401 89608 3436 89648
rect 3476 89608 3532 89648
rect 3572 89608 3581 89648
rect 3785 89608 3820 89648
rect 3860 89608 3916 89648
rect 3956 89608 3965 89648
rect 4291 89608 4300 89648
rect 4340 89608 4349 89648
rect 13027 89608 13036 89648
rect 13076 89608 13172 89648
rect 13507 89608 13516 89648
rect 13556 89608 13612 89648
rect 13652 89608 13687 89648
rect 14716 89608 15043 89648
rect 15083 89608 15092 89648
rect 15331 89608 15340 89648
rect 15380 89608 18028 89648
rect 18068 89608 18077 89648
rect 18979 89608 18988 89648
rect 19028 89608 19316 89648
rect 19363 89608 19372 89648
rect 19412 89608 19468 89648
rect 19508 89608 19543 89648
rect 19747 89608 19756 89648
rect 19796 89608 19927 89648
rect 20009 89608 20140 89648
rect 20180 89608 20189 89648
rect 21388 89608 21600 89648
rect 1612 89564 1652 89608
rect 2380 89564 2420 89608
rect 163 89524 172 89564
rect 212 89524 1652 89564
rect 2083 89524 2092 89564
rect 2132 89524 2420 89564
rect 2476 89524 2708 89564
rect 0 89480 90 89500
rect 2476 89480 2516 89524
rect 0 89440 1420 89480
rect 1460 89440 1469 89480
rect 2227 89440 2236 89480
rect 2276 89440 2516 89480
rect 0 89420 90 89440
rect 2668 89396 2708 89524
rect 2764 89480 2804 89608
rect 4300 89564 4340 89608
rect 5932 89564 5972 89573
rect 12652 89564 12692 89573
rect 13132 89564 13172 89608
rect 14188 89564 14228 89573
rect 14716 89564 14756 89608
rect 2851 89524 2860 89564
rect 2900 89524 4340 89564
rect 4553 89524 4684 89564
rect 4724 89524 4733 89564
rect 5972 89524 9292 89564
rect 9332 89524 9341 89564
rect 11273 89524 11404 89564
rect 11444 89524 11453 89564
rect 12692 89524 12748 89564
rect 12788 89524 12823 89564
rect 13114 89524 13123 89564
rect 13163 89524 13172 89564
rect 13219 89524 13228 89564
rect 13268 89524 13277 89564
rect 13577 89524 13708 89564
rect 13748 89524 13757 89564
rect 13804 89524 14188 89564
rect 14698 89524 14707 89564
rect 14747 89524 14756 89564
rect 15244 89564 15284 89573
rect 16492 89564 16532 89608
rect 18124 89564 18164 89573
rect 19276 89564 19316 89608
rect 21510 89588 21600 89608
rect 16483 89524 16492 89564
rect 16532 89524 16541 89564
rect 16771 89524 16780 89564
rect 16820 89524 16876 89564
rect 16916 89524 16951 89564
rect 17993 89524 18124 89564
rect 18164 89524 18173 89564
rect 19276 89524 19564 89564
rect 19604 89524 19613 89564
rect 5932 89480 5972 89524
rect 2764 89440 3244 89480
rect 3284 89440 3293 89480
rect 4003 89440 4012 89480
rect 4052 89440 5972 89480
rect 6211 89440 6220 89480
rect 6260 89440 10060 89480
rect 10100 89440 10109 89480
rect 11404 89396 11444 89524
rect 12652 89515 12692 89524
rect 13228 89480 13268 89524
rect 13804 89480 13844 89524
rect 14188 89515 14228 89524
rect 15244 89480 15284 89524
rect 18124 89515 18164 89524
rect 12835 89440 12844 89480
rect 12884 89440 13268 89480
rect 13795 89440 13804 89480
rect 13844 89440 13853 89480
rect 15244 89440 17260 89480
rect 17300 89440 17309 89480
rect 19219 89440 19228 89480
rect 19268 89440 20620 89480
rect 20660 89440 20669 89480
rect 1459 89356 1468 89396
rect 1508 89356 1612 89396
rect 1652 89356 1661 89396
rect 1843 89356 1852 89396
rect 1892 89356 2420 89396
rect 2668 89356 3052 89396
rect 3092 89356 3101 89396
rect 3379 89356 3388 89396
rect 3428 89356 3628 89396
rect 3668 89356 3677 89396
rect 4531 89356 4540 89396
rect 4580 89356 6068 89396
rect 6115 89356 6124 89396
rect 6164 89356 6412 89396
rect 6452 89356 6461 89396
rect 11404 89356 12788 89396
rect 12835 89356 12844 89396
rect 12884 89356 14380 89396
rect 14420 89356 14429 89396
rect 14729 89356 14860 89396
rect 14900 89356 14909 89396
rect 2380 89312 2420 89356
rect 6028 89312 6068 89356
rect 1411 89272 1420 89312
rect 1460 89272 2036 89312
rect 2380 89272 5972 89312
rect 6028 89272 12556 89312
rect 12596 89272 12605 89312
rect 1996 89228 2036 89272
rect 5932 89228 5972 89272
rect 12748 89228 12788 89356
rect 15244 89312 15284 89440
rect 17635 89356 17644 89396
rect 17684 89356 18316 89396
rect 18356 89356 18365 89396
rect 19603 89356 19612 89396
rect 19652 89356 19661 89396
rect 20371 89356 20380 89396
rect 20420 89356 21100 89396
rect 21140 89356 21149 89396
rect 12940 89272 13076 89312
rect 13123 89272 13132 89312
rect 13172 89272 15284 89312
rect 19612 89312 19652 89356
rect 19612 89272 20716 89312
rect 20756 89272 20765 89312
rect 12940 89228 12980 89272
rect 1996 89188 3820 89228
rect 3860 89188 3869 89228
rect 4919 89188 4928 89228
rect 4968 89188 5010 89228
rect 5050 89188 5092 89228
rect 5132 89188 5174 89228
rect 5214 89188 5256 89228
rect 5296 89188 5305 89228
rect 5932 89188 6220 89228
rect 6260 89188 6269 89228
rect 12748 89188 12980 89228
rect 13036 89228 13076 89272
rect 13036 89188 13900 89228
rect 13940 89188 13949 89228
rect 20039 89188 20048 89228
rect 20088 89188 20130 89228
rect 20170 89188 20212 89228
rect 20252 89188 20294 89228
rect 20334 89188 20376 89228
rect 20416 89188 20425 89228
rect 0 89144 90 89164
rect 21510 89144 21600 89164
rect 0 89104 3532 89144
rect 3572 89104 3581 89144
rect 12835 89104 12844 89144
rect 12884 89104 14708 89144
rect 20995 89104 21004 89144
rect 21044 89104 21600 89144
rect 0 89084 90 89104
rect 2611 89020 2620 89060
rect 2660 89020 5356 89060
rect 5396 89020 5405 89060
rect 9427 89020 9436 89060
rect 9476 89020 11692 89060
rect 11732 89020 11741 89060
rect 12076 89020 13132 89060
rect 13172 89020 13181 89060
rect 14153 89020 14284 89060
rect 14324 89020 14333 89060
rect 172 88936 2420 88976
rect 3523 88936 3532 88976
rect 3572 88936 5780 88976
rect 0 88808 90 88828
rect 0 88768 76 88808
rect 116 88768 125 88808
rect 0 88748 90 88768
rect 172 88640 212 88936
rect 1219 88852 1228 88892
rect 1268 88852 2036 88892
rect 1996 88808 2036 88852
rect 2380 88808 2420 88936
rect 2633 88852 2764 88892
rect 2804 88852 2813 88892
rect 3043 88852 3052 88892
rect 3092 88852 4012 88892
rect 4052 88852 4061 88892
rect 4387 88852 4396 88892
rect 4436 88852 4492 88892
rect 4532 88852 4567 88892
rect 5740 88883 5780 88936
rect 12076 88892 12116 89020
rect 12259 88936 12268 88976
rect 12308 88936 14132 88976
rect 4012 88834 4052 88843
rect 355 88768 364 88808
rect 404 88768 1228 88808
rect 1268 88768 1277 88808
rect 1603 88768 1612 88808
rect 1652 88768 1661 88808
rect 1987 88768 1996 88808
rect 2036 88768 2045 88808
rect 2371 88768 2380 88808
rect 2420 88768 2429 88808
rect 1612 88724 1652 88768
rect 4492 88724 4532 88852
rect 5740 88834 5780 88843
rect 7276 88883 8468 88892
rect 7316 88852 8468 88883
rect 8515 88852 8524 88892
rect 8564 88852 8716 88892
rect 8756 88852 8765 88892
rect 10723 88852 10732 88892
rect 10772 88852 10828 88892
rect 10868 88852 10903 88892
rect 11945 88852 11980 88892
rect 12020 88883 12116 88892
rect 12020 88852 12076 88883
rect 7276 88834 7316 88843
rect 6115 88768 6124 88808
rect 6164 88768 6173 88808
rect 6124 88724 6164 88768
rect 451 88684 460 88724
rect 500 88684 1652 88724
rect 2227 88684 2236 88724
rect 2276 88684 2956 88724
rect 2996 88684 3005 88724
rect 4492 88684 6164 88724
rect 8428 88724 8468 88852
rect 12163 88852 12172 88892
rect 12212 88852 12547 88892
rect 12587 88852 12596 88892
rect 12643 88852 12652 88892
rect 12692 88852 12844 88892
rect 12884 88852 12893 88892
rect 13027 88852 13036 88892
rect 13076 88852 13516 88892
rect 13556 88852 13565 88892
rect 13612 88883 13996 88892
rect 12076 88834 12116 88843
rect 13652 88852 13996 88883
rect 14036 88852 14045 88892
rect 14092 88883 14132 88936
rect 14668 88892 14708 89104
rect 21510 89084 21600 89104
rect 16169 89020 16300 89060
rect 16340 89020 16349 89060
rect 19987 88936 19996 88976
rect 20036 88936 21484 88976
rect 21524 88936 21533 88976
rect 13612 88834 13652 88843
rect 14371 88852 14380 88892
rect 14420 88852 14563 88892
rect 14603 88852 14612 88892
rect 14659 88852 14668 88892
rect 14708 88852 14717 88892
rect 15043 88852 15052 88892
rect 15092 88852 15101 88892
rect 15628 88883 15668 88892
rect 14092 88834 14132 88843
rect 15052 88808 15092 88852
rect 15977 88852 16108 88892
rect 16148 88852 16157 88892
rect 16771 88852 16780 88892
rect 16820 88852 16876 88892
rect 16916 88852 16951 88892
rect 17251 88852 17260 88892
rect 17300 88883 18164 88892
rect 17300 88852 18124 88883
rect 9161 88768 9196 88808
rect 9236 88768 9292 88808
rect 9332 88768 9532 88808
rect 9572 88768 9581 88808
rect 9763 88768 9772 88808
rect 9812 88768 10156 88808
rect 10196 88768 10205 88808
rect 10505 88768 10636 88808
rect 10676 88768 10685 88808
rect 13123 88768 13132 88808
rect 13172 88768 13303 88808
rect 14275 88768 14284 88808
rect 14324 88768 15092 88808
rect 15139 88768 15148 88808
rect 15188 88768 15197 88808
rect 10156 88724 10196 88768
rect 15148 88724 15188 88768
rect 8428 88684 9908 88724
rect 10156 88684 10924 88724
rect 10964 88684 10973 88724
rect 13699 88684 13708 88724
rect 13748 88684 15188 88724
rect 9868 88640 9908 88684
rect 15628 88640 15668 88843
rect 16108 88834 16148 88843
rect 18124 88834 18164 88843
rect 18473 88768 18604 88808
rect 18644 88768 18653 88808
rect 18857 88768 18988 88808
rect 19028 88768 19037 88808
rect 19241 88768 19372 88808
rect 19412 88768 19421 88808
rect 19625 88768 19756 88808
rect 19796 88768 19805 88808
rect 20131 88768 20140 88808
rect 20180 88768 20311 88808
rect 20371 88768 20380 88808
rect 20420 88768 21388 88808
rect 21428 88768 21437 88808
rect 18835 88684 18844 88724
rect 18884 88684 20236 88724
rect 20276 88684 20285 88724
rect 21510 88640 21600 88660
rect 67 88600 76 88640
rect 116 88600 212 88640
rect 1459 88600 1468 88640
rect 1508 88600 1517 88640
rect 1843 88600 1852 88640
rect 1892 88600 2420 88640
rect 4195 88600 4204 88640
rect 4244 88600 4780 88640
rect 4820 88600 4829 88640
rect 5923 88600 5932 88640
rect 5972 88600 6220 88640
rect 6260 88600 6269 88640
rect 6355 88600 6364 88640
rect 6404 88600 6452 88640
rect 6953 88600 7084 88640
rect 7124 88600 7133 88640
rect 9859 88600 9868 88640
rect 9908 88600 9916 88640
rect 9956 88600 10039 88640
rect 10387 88600 10396 88640
rect 10436 88600 10540 88640
rect 10580 88600 10589 88640
rect 13795 88600 13804 88640
rect 13844 88600 15668 88640
rect 18307 88600 18316 88640
rect 18356 88600 18700 88640
rect 18740 88600 18749 88640
rect 19219 88600 19228 88640
rect 19268 88600 19277 88640
rect 19603 88600 19612 88640
rect 19652 88600 20332 88640
rect 20372 88600 20381 88640
rect 20611 88600 20620 88640
rect 20660 88600 21600 88640
rect 0 88472 90 88492
rect 0 88432 1132 88472
rect 1172 88432 1181 88472
rect 0 88412 90 88432
rect 1468 88388 1508 88600
rect 2380 88556 2420 88600
rect 6412 88556 6452 88600
rect 19228 88556 19268 88600
rect 21510 88580 21600 88600
rect 2380 88516 4340 88556
rect 4387 88516 4396 88556
rect 4436 88516 8524 88556
rect 8564 88516 8573 88556
rect 12940 88516 13132 88556
rect 13172 88516 13181 88556
rect 13507 88516 13516 88556
rect 13556 88516 14284 88556
rect 14324 88516 14333 88556
rect 19228 88516 21004 88556
rect 21044 88516 21053 88556
rect 4300 88472 4340 88516
rect 12940 88472 12980 88516
rect 3679 88432 3688 88472
rect 3728 88432 3770 88472
rect 3810 88432 3852 88472
rect 3892 88432 3934 88472
rect 3974 88432 4016 88472
rect 4056 88432 4065 88472
rect 4300 88432 10348 88472
rect 10388 88432 12980 88472
rect 18799 88432 18808 88472
rect 18848 88432 18890 88472
rect 18930 88432 18972 88472
rect 19012 88432 19054 88472
rect 19094 88432 19136 88472
rect 19176 88432 19185 88472
rect 1468 88348 12980 88388
rect 12940 88304 12980 88348
rect 1996 88264 2476 88304
rect 2516 88264 2525 88304
rect 8611 88264 8620 88304
rect 8660 88264 8668 88304
rect 8708 88264 8791 88304
rect 12041 88264 12172 88304
rect 12212 88264 12221 88304
rect 12665 88264 12748 88304
rect 12788 88264 12796 88304
rect 12836 88264 12845 88304
rect 12940 88264 18796 88304
rect 18836 88264 18845 88304
rect 547 88180 556 88220
rect 596 88180 1268 88220
rect 0 88136 90 88156
rect 1228 88136 1268 88180
rect 1996 88136 2036 88264
rect 0 88096 1172 88136
rect 1219 88096 1228 88136
rect 1268 88096 1277 88136
rect 1891 88096 1900 88136
rect 1940 88096 2036 88136
rect 2092 88180 3340 88220
rect 3380 88180 3389 88220
rect 9091 88180 9100 88220
rect 9140 88180 12980 88220
rect 13123 88180 13132 88220
rect 13172 88180 13652 88220
rect 0 88076 90 88096
rect 1132 88052 1172 88096
rect 2092 88052 2132 88180
rect 2275 88096 2284 88136
rect 2324 88096 2900 88136
rect 4265 88096 4396 88136
rect 4436 88096 4445 88136
rect 5321 88096 5356 88136
rect 5396 88096 5452 88136
rect 5492 88096 5501 88136
rect 8777 88096 8908 88136
rect 8948 88096 8957 88136
rect 10627 88096 10636 88136
rect 10676 88096 10685 88136
rect 10915 88096 10924 88136
rect 10964 88096 12556 88136
rect 12596 88096 12605 88136
rect 1132 88012 2132 88052
rect 2633 88012 2764 88052
rect 2804 88012 2813 88052
rect 2131 87928 2140 87968
rect 2180 87928 2476 87968
rect 2516 87928 2525 87968
rect 1459 87844 1468 87884
rect 1508 87844 2092 87884
rect 2132 87844 2141 87884
rect 2515 87844 2524 87884
rect 2564 87844 2764 87884
rect 2804 87844 2813 87884
rect 0 87800 90 87820
rect 0 87760 2572 87800
rect 2612 87760 2621 87800
rect 0 87740 90 87760
rect 2860 87632 2900 88096
rect 4012 88052 4052 88061
rect 5932 88052 5972 88061
rect 6988 88052 7028 88061
rect 9292 88052 9332 88061
rect 10636 88052 10676 88096
rect 12940 88052 12980 88180
rect 13385 88096 13516 88136
rect 13556 88096 13565 88136
rect 13612 88052 13652 88180
rect 13996 88180 16436 88220
rect 17923 88180 17932 88220
rect 17972 88180 19892 88220
rect 3523 88012 3532 88052
rect 3572 88012 4012 88052
rect 4052 88012 4061 88052
rect 4204 88012 4867 88052
rect 4907 88012 4916 88052
rect 4963 88012 4972 88052
rect 5012 88012 5021 88052
rect 5347 88012 5356 88052
rect 5396 88012 5452 88052
rect 5492 88012 5644 88052
rect 5684 88012 5693 88052
rect 5801 88012 5836 88052
rect 5876 88012 5932 88052
rect 6211 88012 6220 88052
rect 6260 88012 6420 88052
rect 6460 88012 6469 88052
rect 8227 88012 8236 88052
rect 8276 88012 8716 88052
rect 8756 88012 8765 88052
rect 9161 88012 9292 88052
rect 9332 88012 9341 88052
rect 10409 88012 10540 88052
rect 10580 88012 10589 88052
rect 10636 88012 10732 88052
rect 10772 88012 10781 88052
rect 11837 88012 11980 88052
rect 12028 88012 12556 88052
rect 12596 88012 12605 88052
rect 12940 88012 13027 88052
rect 13067 88012 13076 88052
rect 13123 88012 13132 88052
rect 13172 88012 13303 88052
rect 13603 88012 13612 88052
rect 13652 88012 13661 88052
rect 4012 88003 4052 88012
rect 4204 87968 4244 88012
rect 4978 87968 5018 88012
rect 5932 88003 5972 88012
rect 6988 87968 7028 88012
rect 4195 87928 4204 87968
rect 4244 87928 4253 87968
rect 4978 87928 5548 87968
rect 5588 87928 5597 87968
rect 6988 87928 8620 87968
rect 8660 87928 8669 87968
rect 8716 87884 8756 88012
rect 9292 88003 9332 88012
rect 10540 87968 10580 88012
rect 13996 87968 14036 88180
rect 14476 88096 15188 88136
rect 14092 88052 14132 88061
rect 14083 88012 14092 88052
rect 14132 88012 14263 88052
rect 14092 88003 14132 88012
rect 10540 87928 11116 87968
rect 11156 87928 11165 87968
rect 12076 87928 14036 87968
rect 12076 87884 12116 87928
rect 14476 87884 14516 88096
rect 15148 88052 15188 88096
rect 16396 88052 16436 88180
rect 18089 88096 18220 88136
rect 18260 88096 18269 88136
rect 17836 88052 17876 88061
rect 19852 88052 19892 88180
rect 21510 88136 21600 88156
rect 20803 88096 20812 88136
rect 20852 88096 21600 88136
rect 21510 88076 21600 88096
rect 14602 88012 14611 88052
rect 14651 88012 14996 88052
rect 14956 87968 14996 88012
rect 16387 88012 16396 88052
rect 16436 88012 16445 88052
rect 16579 88012 16588 88052
rect 16628 88012 16759 88052
rect 17876 88012 18124 88052
rect 18164 88012 18173 88052
rect 18499 88012 18508 88052
rect 18548 88012 18604 88052
rect 18644 88012 18679 88052
rect 15148 87968 15188 88012
rect 17836 87968 17876 88012
rect 19852 88003 19892 88012
rect 14947 87928 14956 87968
rect 14996 87928 15005 87968
rect 15148 87928 15628 87968
rect 15668 87928 17876 87968
rect 18019 87928 18028 87968
rect 18068 87928 19276 87968
rect 19316 87928 19325 87968
rect 20227 87928 20236 87968
rect 20276 87928 21575 87968
rect 4627 87844 4636 87884
rect 4676 87844 5356 87884
rect 5396 87844 5405 87884
rect 5923 87844 5932 87884
rect 5972 87844 6604 87884
rect 6644 87844 6653 87884
rect 6787 87844 6796 87884
rect 6836 87844 7372 87884
rect 7412 87844 7421 87884
rect 8716 87844 9292 87884
rect 9332 87844 9341 87884
rect 11299 87844 11308 87884
rect 11348 87844 12116 87884
rect 12739 87844 12748 87884
rect 12788 87844 14516 87884
rect 14755 87844 14764 87884
rect 14804 87844 15340 87884
rect 15380 87844 15389 87884
rect 18451 87844 18460 87884
rect 18500 87844 19796 87884
rect 19843 87844 19852 87884
rect 19892 87844 20044 87884
rect 20084 87844 20093 87884
rect 4483 87760 4492 87800
rect 4532 87760 9140 87800
rect 9187 87760 9196 87800
rect 9236 87760 12844 87800
rect 12884 87760 12893 87800
rect 9100 87716 9140 87760
rect 4919 87676 4928 87716
rect 4968 87676 5010 87716
rect 5050 87676 5092 87716
rect 5132 87676 5174 87716
rect 5214 87676 5256 87716
rect 5296 87676 5305 87716
rect 9100 87676 10060 87716
rect 10100 87676 10109 87716
rect 10435 87676 10444 87716
rect 10484 87676 17836 87716
rect 17876 87676 17885 87716
rect 2860 87592 4052 87632
rect 0 87464 90 87484
rect 2860 87464 2900 87592
rect 4012 87464 4052 87592
rect 9100 87592 9868 87632
rect 9908 87592 12884 87632
rect 12931 87592 12940 87632
rect 12980 87592 15140 87632
rect 6473 87508 6604 87548
rect 6644 87508 6653 87548
rect 8585 87508 8716 87548
rect 8756 87508 8765 87548
rect 0 87424 1516 87464
rect 1556 87424 1565 87464
rect 2467 87424 2476 87464
rect 2516 87424 2900 87464
rect 3859 87424 3868 87464
rect 3908 87424 4052 87464
rect 5164 87424 5548 87464
rect 5588 87424 5597 87464
rect 6988 87424 7084 87464
rect 7124 87424 7133 87464
rect 8899 87424 8908 87464
rect 8948 87424 8957 87464
rect 0 87404 90 87424
rect 2476 87380 2516 87424
rect 5164 87380 5204 87424
rect 6988 87380 7028 87424
rect 8908 87380 8948 87424
rect 1603 87340 1612 87380
rect 1652 87340 2516 87380
rect 2729 87340 2860 87380
rect 2900 87340 3052 87380
rect 3092 87340 3101 87380
rect 4715 87340 4780 87380
rect 4820 87340 4846 87380
rect 4886 87340 4895 87380
rect 4963 87340 4972 87380
rect 5012 87340 5164 87380
rect 5204 87340 5213 87380
rect 5347 87340 5356 87380
rect 5396 87340 5452 87380
rect 5492 87340 5556 87380
rect 5827 87340 5836 87380
rect 5876 87371 6007 87380
rect 5876 87340 5932 87371
rect 2860 87322 2900 87331
rect 1219 87256 1228 87296
rect 1268 87256 1324 87296
rect 1364 87256 1399 87296
rect 3331 87256 3340 87296
rect 3380 87256 3436 87296
rect 3476 87256 3511 87296
rect 3619 87256 3628 87296
rect 3668 87256 3799 87296
rect 4003 87256 4012 87296
rect 4052 87256 4061 87296
rect 4579 87256 4588 87296
rect 4628 87256 4637 87296
rect 4012 87212 4052 87256
rect 1603 87172 1612 87212
rect 1652 87172 4052 87212
rect 4108 87172 4252 87212
rect 4292 87172 4301 87212
rect 0 87128 90 87148
rect 4108 87128 4148 87172
rect 4588 87128 4628 87256
rect 5356 87212 5396 87340
rect 5972 87340 6007 87371
rect 6281 87340 6412 87380
rect 6452 87340 6461 87380
rect 6970 87340 6979 87380
rect 7019 87340 7028 87380
rect 7075 87340 7084 87380
rect 7124 87340 7171 87380
rect 7459 87340 7468 87380
rect 7508 87340 7700 87380
rect 7913 87340 7948 87380
rect 7988 87371 8084 87380
rect 7988 87340 8044 87371
rect 5932 87322 5972 87331
rect 6412 87322 6452 87331
rect 7084 87296 7124 87340
rect 5443 87256 5452 87296
rect 5492 87256 5644 87296
rect 5684 87256 5693 87296
rect 7075 87256 7084 87296
rect 7124 87256 7133 87296
rect 7555 87256 7564 87296
rect 7604 87256 7613 87296
rect 7564 87212 7604 87256
rect 5196 87172 5260 87212
rect 5300 87172 7604 87212
rect 7660 87128 7700 87340
rect 8044 87322 8084 87331
rect 8524 87371 8948 87380
rect 8564 87340 8948 87371
rect 9100 87371 9140 87592
rect 12844 87548 12884 87592
rect 12355 87508 12364 87548
rect 12404 87508 12692 87548
rect 12844 87508 13036 87548
rect 13076 87508 13085 87548
rect 13315 87508 13324 87548
rect 13364 87508 13516 87548
rect 13556 87508 13565 87548
rect 12652 87464 12692 87508
rect 12652 87424 12884 87464
rect 12844 87380 12884 87424
rect 12988 87424 13132 87464
rect 13172 87424 13181 87464
rect 12988 87380 13028 87424
rect 15100 87380 15140 87592
rect 19756 87548 19796 87844
rect 21535 87800 21575 87928
rect 21388 87760 21575 87800
rect 20039 87676 20048 87716
rect 20088 87676 20130 87716
rect 20170 87676 20212 87716
rect 20252 87676 20294 87716
rect 20334 87676 20376 87716
rect 20416 87676 20425 87716
rect 21388 87632 21428 87760
rect 21510 87632 21600 87652
rect 21388 87592 21600 87632
rect 21510 87572 21600 87592
rect 19756 87508 20236 87548
rect 20276 87508 20285 87548
rect 17321 87424 17443 87464
rect 17492 87424 17501 87464
rect 8524 87322 8564 87331
rect 9100 87322 9140 87331
rect 10060 87340 10348 87380
rect 10388 87340 10397 87380
rect 10732 87340 11116 87380
rect 11156 87340 11165 87380
rect 12163 87340 12172 87380
rect 12212 87371 12404 87380
rect 12212 87340 12364 87371
rect 10060 87212 10100 87340
rect 10732 87296 10772 87340
rect 12739 87340 12748 87380
rect 12788 87340 12797 87380
rect 12844 87340 12863 87380
rect 12903 87340 12912 87380
rect 12988 87340 13036 87380
rect 13076 87340 13085 87380
rect 13228 87359 13267 87380
rect 13132 87340 13267 87359
rect 13307 87340 13316 87380
rect 12364 87322 12404 87331
rect 10601 87256 10732 87296
rect 10772 87256 10781 87296
rect 12748 87212 12788 87340
rect 13132 87319 13268 87340
rect 13132 87212 13172 87319
rect 13360 87308 13369 87348
rect 13409 87308 13418 87348
rect 15100 87340 15724 87380
rect 15764 87340 16588 87380
rect 16628 87340 16637 87380
rect 16972 87371 17260 87380
rect 17012 87340 17260 87371
rect 17300 87340 17309 87380
rect 17513 87340 17635 87380
rect 17684 87340 17693 87380
rect 18124 87371 18316 87380
rect 16972 87322 17012 87331
rect 18164 87340 18316 87371
rect 18356 87340 18365 87380
rect 18473 87340 18604 87380
rect 18644 87340 18653 87380
rect 19075 87340 19084 87380
rect 19124 87340 19133 87380
rect 19193 87340 19202 87380
rect 19242 87340 19276 87380
rect 19316 87340 19382 87380
rect 18124 87322 18164 87331
rect 13378 87212 13418 87308
rect 18403 87256 18412 87296
rect 18452 87256 18700 87296
rect 18740 87256 18749 87296
rect 19084 87212 19124 87340
rect 19625 87256 19756 87296
rect 19796 87256 19805 87296
rect 20009 87256 20140 87296
rect 20180 87256 20189 87296
rect 20371 87256 20380 87296
rect 20420 87256 21484 87296
rect 21524 87256 21533 87296
rect 8803 87172 8812 87212
rect 8852 87172 10100 87212
rect 12547 87172 12556 87212
rect 12596 87172 13268 87212
rect 13315 87172 13324 87212
rect 13364 87172 13418 87212
rect 17731 87172 17740 87212
rect 17780 87172 19124 87212
rect 13228 87128 13268 87172
rect 21510 87128 21600 87148
rect 0 87088 748 87128
rect 788 87088 797 87128
rect 1459 87088 1468 87128
rect 1508 87088 1516 87128
rect 1556 87088 1639 87128
rect 2921 87088 3052 87128
rect 3092 87088 3101 87128
rect 3187 87088 3196 87128
rect 3236 87088 3340 87128
rect 3380 87088 3389 87128
rect 3523 87088 3532 87128
rect 3572 87088 4148 87128
rect 4339 87088 4348 87128
rect 4388 87088 4532 87128
rect 4588 87088 5452 87128
rect 5492 87088 5501 87128
rect 6403 87088 6412 87128
rect 6452 87088 9388 87128
rect 9428 87088 9437 87128
rect 10963 87088 10972 87128
rect 11012 87088 11308 87128
rect 11348 87088 11357 87128
rect 12739 87088 12748 87128
rect 12788 87088 12797 87128
rect 13219 87088 13228 87128
rect 13268 87088 13277 87128
rect 17155 87088 17164 87128
rect 17204 87088 17213 87128
rect 17635 87088 17644 87128
rect 17684 87088 17836 87128
rect 17876 87088 17885 87128
rect 18115 87088 18124 87128
rect 18164 87088 18604 87128
rect 18644 87088 18653 87128
rect 19987 87088 19996 87128
rect 20036 87088 20045 87128
rect 20707 87088 20716 87128
rect 20756 87088 21600 87128
rect 0 87068 90 87088
rect 4492 87044 4532 87088
rect 4492 87004 9100 87044
rect 9140 87004 9149 87044
rect 3679 86920 3688 86960
rect 3728 86920 3770 86960
rect 3810 86920 3852 86960
rect 3892 86920 3934 86960
rect 3974 86920 4016 86960
rect 4056 86920 4065 86960
rect 6844 86836 10732 86876
rect 10772 86836 10781 86876
rect 0 86792 90 86812
rect 6844 86792 6884 86836
rect 0 86752 1420 86792
rect 1460 86752 1469 86792
rect 1516 86752 1844 86792
rect 2633 86752 2764 86792
rect 2804 86752 2813 86792
rect 5635 86752 5644 86792
rect 5684 86752 5693 86792
rect 6835 86752 6844 86792
rect 6884 86752 6893 86792
rect 8899 86752 8908 86792
rect 8948 86752 9235 86792
rect 9275 86752 9284 86792
rect 9619 86752 9628 86792
rect 9668 86752 10060 86792
rect 10100 86752 10109 86792
rect 10291 86752 10300 86792
rect 10340 86752 10444 86792
rect 10484 86752 10493 86792
rect 10675 86752 10684 86792
rect 10724 86752 11212 86792
rect 11252 86752 11261 86792
rect 12233 86752 12268 86792
rect 12308 86752 12364 86792
rect 12404 86752 12413 86792
rect 0 86732 90 86752
rect 1516 86708 1556 86752
rect 1804 86708 1844 86752
rect 172 86668 1556 86708
rect 1603 86668 1612 86708
rect 1652 86668 1661 86708
rect 1804 86668 3436 86708
rect 3476 86668 3485 86708
rect 3532 86668 4492 86708
rect 4532 86668 5548 86708
rect 5588 86668 5597 86708
rect 0 86456 90 86476
rect 172 86456 212 86668
rect 1612 86624 1652 86668
rect 3532 86624 3572 86668
rect 5644 86624 5684 86752
rect 6115 86668 6124 86708
rect 6164 86668 6788 86708
rect 6748 86624 6788 86668
rect 8140 86668 10100 86708
rect 11683 86668 11692 86708
rect 11732 86668 12500 86708
rect 0 86416 212 86456
rect 1228 86584 1652 86624
rect 2572 86584 2860 86624
rect 2900 86584 2909 86624
rect 2956 86584 3572 86624
rect 5033 86584 5164 86624
rect 5204 86584 5213 86624
rect 5644 86584 5780 86624
rect 6019 86584 6028 86624
rect 6068 86584 6604 86624
rect 6644 86584 6653 86624
rect 6748 86584 6988 86624
rect 7028 86584 7180 86624
rect 7220 86584 7229 86624
rect 7843 86584 7852 86624
rect 7892 86584 7948 86624
rect 7988 86584 8023 86624
rect 0 86396 90 86416
rect 0 86120 90 86140
rect 0 86080 1132 86120
rect 1172 86080 1181 86120
rect 0 86060 90 86080
rect 1228 86036 1268 86584
rect 2572 86540 2612 86584
rect 2956 86540 2996 86584
rect 4204 86540 4244 86549
rect 5740 86540 5780 86584
rect 1315 86500 1324 86540
rect 1364 86500 1612 86540
rect 1652 86500 1940 86540
rect 1900 86372 1940 86500
rect 2947 86500 2956 86540
rect 2996 86500 3005 86540
rect 4003 86500 4012 86540
rect 4052 86500 4204 86540
rect 2572 86491 2612 86500
rect 4204 86491 4244 86500
rect 4396 86500 4675 86540
rect 4715 86500 4724 86540
rect 4771 86500 4780 86540
rect 4820 86500 4829 86540
rect 5129 86500 5260 86540
rect 5300 86500 5644 86540
rect 5684 86500 5693 86540
rect 5827 86500 5836 86540
rect 5876 86500 6228 86540
rect 6268 86500 6277 86540
rect 7307 86500 7372 86540
rect 7412 86500 7438 86540
rect 7478 86500 7487 86540
rect 7555 86500 7564 86540
rect 7604 86500 7613 86540
rect 7913 86500 7948 86540
rect 7988 86500 8044 86540
rect 8084 86500 8093 86540
rect 4396 86456 4436 86500
rect 4780 86456 4820 86500
rect 5740 86491 5780 86500
rect 7564 86456 7604 86500
rect 8140 86456 8180 86668
rect 10060 86624 10100 86668
rect 12460 86624 12500 86668
rect 9283 86584 9292 86624
rect 9332 86584 9388 86624
rect 9428 86584 9463 86624
rect 10051 86584 10060 86624
rect 10100 86584 10109 86624
rect 10435 86584 10444 86624
rect 10484 86584 10493 86624
rect 12451 86584 12460 86624
rect 12500 86584 12509 86624
rect 8523 86540 8563 86549
rect 8227 86500 8236 86540
rect 8276 86500 8523 86540
rect 8611 86500 8620 86540
rect 8660 86500 9012 86540
rect 9052 86500 9061 86540
rect 8523 86491 8563 86500
rect 10444 86456 10484 86584
rect 12076 86540 12116 86549
rect 12748 86540 12788 87088
rect 13027 86668 13036 86708
rect 13076 86668 15188 86708
rect 15148 86624 15188 86668
rect 12931 86584 12940 86624
rect 12980 86584 13130 86624
rect 13219 86584 13228 86624
rect 13268 86584 13315 86624
rect 15148 86584 16820 86624
rect 13090 86540 13130 86584
rect 13228 86540 13268 86584
rect 15148 86540 15188 86584
rect 16780 86540 16820 86584
rect 17164 86540 17204 87088
rect 18799 86920 18808 86960
rect 18848 86920 18890 86960
rect 18930 86920 18972 86960
rect 19012 86920 19054 86960
rect 19094 86920 19136 86960
rect 19176 86920 19185 86960
rect 19996 86792 20036 87088
rect 21510 87068 21600 87088
rect 19996 86752 20908 86792
rect 20948 86752 20957 86792
rect 21510 86624 21600 86644
rect 17251 86584 17260 86624
rect 17300 86584 18028 86624
rect 18068 86584 18412 86624
rect 18452 86584 18461 86624
rect 19625 86584 19756 86624
rect 19796 86584 19805 86624
rect 20009 86584 20140 86624
rect 20180 86584 20189 86624
rect 21283 86584 21292 86624
rect 21332 86584 21600 86624
rect 21510 86564 21600 86584
rect 18604 86540 18644 86549
rect 10627 86500 10636 86540
rect 10676 86500 10828 86540
rect 10868 86500 10877 86540
rect 12041 86500 12076 86540
rect 12116 86500 12172 86540
rect 12212 86500 12221 86540
rect 12748 86500 12835 86540
rect 12875 86500 12884 86540
rect 12940 86500 12953 86540
rect 12993 86500 13002 86540
rect 13076 86500 13085 86540
rect 13125 86500 13134 86540
rect 13210 86500 13219 86540
rect 13259 86500 13268 86540
rect 13354 86500 13363 86540
rect 13403 86500 13412 86540
rect 13603 86500 13612 86540
rect 13652 86500 13900 86540
rect 13940 86500 13949 86540
rect 15401 86500 15532 86540
rect 15572 86500 15581 86540
rect 16820 86500 16916 86540
rect 17164 86500 17539 86540
rect 17579 86500 17588 86540
rect 17635 86500 17644 86540
rect 17684 86500 17740 86540
rect 17780 86500 17815 86540
rect 17993 86500 18124 86540
rect 18164 86500 18173 86540
rect 18307 86500 18316 86540
rect 18356 86500 18604 86540
rect 18691 86500 18700 86540
rect 18740 86500 19092 86540
rect 19132 86500 19141 86540
rect 12076 86491 12116 86500
rect 12940 86456 12980 86500
rect 13372 86456 13412 86500
rect 15148 86491 15188 86500
rect 16780 86491 16820 86500
rect 4387 86416 4396 86456
rect 4436 86416 4445 86456
rect 4780 86416 5588 86456
rect 6115 86416 6124 86456
rect 6164 86416 7084 86456
rect 7124 86416 7604 86456
rect 7660 86416 8180 86456
rect 8707 86416 8716 86456
rect 8756 86416 10484 86456
rect 12259 86416 12268 86456
rect 12308 86416 12980 86456
rect 13027 86416 13036 86456
rect 13076 86416 13123 86456
rect 13219 86416 13228 86456
rect 13268 86416 13412 86456
rect 15331 86416 15340 86456
rect 15380 86416 15511 86456
rect 5548 86372 5588 86416
rect 6124 86372 6164 86416
rect 7660 86372 7700 86416
rect 13036 86372 13076 86416
rect 16876 86372 16916 86500
rect 18604 86491 18644 86500
rect 16963 86416 16972 86456
rect 17012 86416 17143 86456
rect 17260 86416 17452 86456
rect 17492 86416 17932 86456
rect 17972 86416 17981 86456
rect 18787 86416 18796 86456
rect 18836 86416 19316 86456
rect 20371 86416 20380 86456
rect 20420 86416 20716 86456
rect 20756 86416 20765 86456
rect 17260 86372 17300 86416
rect 19276 86372 19316 86416
rect 1900 86332 5452 86372
rect 5492 86332 5501 86372
rect 5548 86332 6164 86372
rect 6281 86332 6412 86372
rect 6452 86332 6461 86372
rect 6691 86332 6700 86372
rect 6740 86332 7228 86372
rect 7268 86332 7700 86372
rect 12547 86332 12556 86372
rect 12596 86332 12700 86372
rect 12740 86332 12749 86372
rect 13027 86332 13036 86372
rect 13076 86332 13085 86372
rect 16876 86332 17300 86372
rect 19267 86332 19276 86372
rect 19316 86332 19325 86372
rect 19865 86332 19948 86372
rect 19988 86332 19996 86372
rect 20036 86332 20045 86372
rect 20227 86332 20236 86372
rect 20276 86332 21292 86372
rect 21332 86332 21341 86372
rect 3235 86248 3244 86288
rect 3284 86248 4012 86288
rect 4052 86248 4780 86288
rect 4820 86248 4829 86288
rect 5356 86248 15724 86288
rect 15764 86248 15773 86288
rect 4919 86164 4928 86204
rect 4968 86164 5010 86204
rect 5050 86164 5092 86204
rect 5132 86164 5174 86204
rect 5214 86164 5256 86204
rect 5296 86164 5305 86204
rect 1411 86080 1420 86120
rect 1460 86080 2476 86120
rect 2516 86080 4396 86120
rect 4436 86080 4445 86120
rect 5356 86036 5396 86248
rect 8332 86164 12460 86204
rect 12500 86164 12509 86204
rect 12556 86164 15244 86204
rect 15284 86164 15293 86204
rect 20039 86164 20048 86204
rect 20088 86164 20130 86204
rect 20170 86164 20212 86204
rect 20252 86164 20294 86204
rect 20334 86164 20376 86204
rect 20416 86164 20425 86204
rect 8332 86036 8372 86164
rect 12556 86120 12596 86164
rect 21510 86120 21600 86140
rect 8812 86080 12596 86120
rect 12835 86080 12844 86120
rect 12884 86080 17932 86120
rect 17972 86080 18124 86120
rect 18164 86080 18173 86120
rect 20995 86080 21004 86120
rect 21044 86080 21600 86120
rect 1219 85996 1228 86036
rect 1268 85996 1277 86036
rect 2371 85996 2380 86036
rect 2420 85996 2429 86036
rect 3955 85996 3964 86036
rect 4004 85996 5396 86036
rect 5705 85996 5836 86036
rect 5876 85996 5885 86036
rect 6739 85996 6748 86036
rect 6788 85996 8372 86036
rect 8489 85996 8620 86036
rect 8660 85996 8669 86036
rect 2380 85952 2420 85996
rect 8812 85952 8852 86080
rect 21510 86060 21600 86080
rect 12425 85996 12508 86036
rect 12548 85996 12556 86036
rect 12596 85996 12605 86036
rect 12652 85996 14284 86036
rect 14324 85996 14333 86036
rect 940 85912 2420 85952
rect 3571 85912 3580 85952
rect 3620 85912 8852 85952
rect 0 85784 90 85804
rect 940 85784 980 85912
rect 12652 85868 12692 85996
rect 12739 85912 12748 85952
rect 12788 85912 12980 85952
rect 12940 85868 12980 85912
rect 13132 85912 13556 85952
rect 13603 85912 13612 85952
rect 13652 85912 13661 85952
rect 16483 85912 16492 85952
rect 16532 85912 18172 85952
rect 18212 85912 18221 85952
rect 13132 85868 13172 85912
rect 13516 85868 13556 85912
rect 13612 85868 13652 85912
rect 1699 85828 1708 85868
rect 1748 85828 2380 85868
rect 2420 85828 2429 85868
rect 2851 85828 2860 85868
rect 2900 85859 3031 85868
rect 2900 85828 2956 85859
rect 2996 85828 3031 85859
rect 3244 85828 3476 85868
rect 4387 85828 4396 85868
rect 4436 85828 4724 85868
rect 4771 85828 4780 85868
rect 4820 85859 5684 85868
rect 4820 85828 5644 85859
rect 2956 85810 2996 85819
rect 0 85744 980 85784
rect 1097 85744 1228 85784
rect 1268 85744 1277 85784
rect 0 85724 90 85744
rect 3244 85700 3284 85828
rect 3436 85784 3476 85828
rect 3331 85744 3340 85784
rect 3380 85744 3389 85784
rect 3436 85744 3724 85784
rect 3764 85744 3773 85784
rect 2467 85660 2476 85700
rect 2516 85660 3284 85700
rect 3340 85700 3380 85744
rect 4684 85700 4724 85828
rect 5644 85784 5684 85819
rect 6316 85828 6932 85868
rect 7049 85828 7180 85868
rect 7220 85828 7229 85868
rect 8428 85859 8563 85868
rect 6316 85784 6356 85828
rect 5644 85744 6076 85784
rect 6116 85744 6125 85784
rect 6307 85744 6316 85784
rect 6356 85744 6365 85784
rect 6499 85744 6508 85784
rect 6548 85744 6679 85784
rect 3340 85660 4492 85700
rect 4532 85660 4541 85700
rect 4684 85660 6700 85700
rect 6740 85660 6749 85700
rect 6892 85616 6932 85828
rect 8468 85828 8563 85859
rect 8681 85828 8812 85868
rect 8852 85828 8861 85868
rect 10060 85859 10252 85868
rect 8428 85810 8468 85819
rect 8523 85784 8563 85828
rect 10100 85828 10252 85859
rect 10292 85828 10301 85868
rect 10435 85828 10444 85868
rect 10484 85828 10493 85868
rect 11692 85859 11884 85868
rect 10060 85810 10100 85819
rect 8523 85744 9004 85784
rect 9044 85744 9053 85784
rect 10444 85700 10484 85828
rect 11732 85828 11884 85859
rect 11924 85828 11933 85868
rect 12233 85828 12364 85868
rect 12404 85828 12413 85868
rect 12643 85828 12652 85868
rect 12692 85828 12701 85868
rect 12826 85828 12835 85868
rect 12875 85828 12884 85868
rect 12940 85828 13132 85868
rect 13172 85828 13181 85868
rect 13360 85828 13369 85868
rect 13409 85828 13460 85868
rect 13507 85828 13516 85868
rect 13556 85828 13565 85868
rect 13612 85828 13804 85868
rect 13844 85828 14092 85868
rect 14132 85828 14141 85868
rect 14921 85828 15052 85868
rect 15092 85828 15101 85868
rect 15401 85828 15436 85868
rect 15476 85828 15532 85868
rect 15572 85828 15581 85868
rect 16684 85859 16724 85868
rect 11692 85810 11732 85819
rect 8803 85660 8812 85700
rect 8852 85660 10484 85700
rect 12844 85700 12884 85828
rect 13420 85784 13460 85828
rect 15052 85784 15092 85819
rect 16684 85784 16724 85819
rect 17260 85828 18508 85868
rect 18548 85828 18604 85868
rect 18644 85828 18679 85868
rect 18892 85859 20044 85868
rect 18892 85828 19852 85859
rect 17260 85784 17300 85828
rect 13027 85744 13036 85784
rect 13076 85744 13207 85784
rect 13258 85775 13316 85784
rect 13258 85735 13267 85775
rect 13307 85735 13316 85775
rect 13420 85744 13612 85784
rect 13652 85744 13661 85784
rect 15052 85744 17204 85784
rect 17251 85744 17260 85784
rect 17300 85744 17309 85784
rect 17443 85744 17452 85784
rect 17492 85744 17623 85784
rect 17827 85744 17836 85784
rect 17876 85744 18007 85784
rect 18281 85744 18412 85784
rect 18452 85744 18461 85784
rect 13258 85734 13316 85735
rect 13276 85700 13316 85734
rect 17164 85700 17204 85744
rect 12844 85660 13172 85700
rect 13276 85660 15820 85700
rect 15860 85660 15869 85700
rect 16675 85660 16684 85700
rect 16724 85660 17020 85700
rect 17060 85660 17069 85700
rect 17164 85660 17972 85700
rect 18067 85660 18076 85700
rect 18116 85660 18220 85700
rect 18260 85660 18269 85700
rect 1459 85576 1468 85616
rect 1508 85576 2572 85616
rect 2612 85576 2621 85616
rect 3139 85576 3148 85616
rect 3188 85576 3197 85616
rect 6892 85576 8908 85616
rect 8948 85576 8957 85616
rect 10243 85576 10252 85616
rect 10292 85576 10444 85616
rect 10484 85576 10493 85616
rect 11875 85576 11884 85616
rect 11924 85576 12556 85616
rect 12596 85576 12605 85616
rect 12713 85576 12835 85616
rect 12884 85576 12893 85616
rect 3148 85532 3188 85576
rect 13132 85532 13172 85660
rect 17932 85616 17972 85660
rect 18892 85616 18932 85828
rect 19892 85828 20044 85859
rect 20084 85828 20093 85868
rect 19852 85810 19892 85819
rect 21510 85616 21600 85636
rect 13651 85576 13660 85616
rect 13700 85576 14380 85616
rect 14420 85576 14429 85616
rect 15235 85576 15244 85616
rect 15284 85576 15293 85616
rect 16867 85576 16876 85616
rect 16916 85576 16925 85616
rect 17683 85576 17692 85616
rect 17732 85576 17741 85616
rect 17932 85576 18124 85616
rect 18164 85576 18932 85616
rect 19363 85576 19372 85616
rect 19412 85576 20044 85616
rect 20084 85576 20093 85616
rect 21187 85576 21196 85616
rect 21236 85576 21600 85616
rect 3148 85492 4300 85532
rect 4340 85492 4349 85532
rect 13132 85492 14860 85532
rect 14900 85492 14909 85532
rect 0 85448 90 85468
rect 0 85408 268 85448
rect 308 85408 317 85448
rect 3679 85408 3688 85448
rect 3728 85408 3770 85448
rect 3810 85408 3852 85448
rect 3892 85408 3934 85448
rect 3974 85408 4016 85448
rect 4056 85408 4065 85448
rect 4387 85408 4396 85448
rect 4436 85408 10636 85448
rect 10676 85408 10685 85448
rect 12355 85408 12364 85448
rect 12404 85408 12748 85448
rect 12788 85408 12797 85448
rect 0 85388 90 85408
rect 1411 85324 1420 85364
rect 1460 85324 8468 85364
rect 2851 85240 2860 85280
rect 2900 85240 4676 85280
rect 5443 85240 5452 85280
rect 5492 85240 8188 85280
rect 8228 85240 8237 85280
rect 2860 85156 3244 85196
rect 3284 85156 3293 85196
rect 0 85112 90 85132
rect 0 85072 844 85112
rect 884 85072 893 85112
rect 0 85052 90 85072
rect 2668 85028 2708 85037
rect 2860 85028 2900 85156
rect 4636 85112 4676 85240
rect 4745 85156 4780 85196
rect 4820 85156 4876 85196
rect 4916 85156 4925 85196
rect 8428 85112 8468 85324
rect 8707 85240 8716 85280
rect 8756 85240 8860 85280
rect 8900 85240 9868 85280
rect 9908 85240 9917 85280
rect 10060 85240 10540 85280
rect 10580 85240 10589 85280
rect 10060 85196 10100 85240
rect 8515 85156 8524 85196
rect 8564 85156 10100 85196
rect 13123 85156 13132 85196
rect 13172 85156 14284 85196
rect 14324 85156 14333 85196
rect 15244 85112 15284 85576
rect 3043 85072 3052 85112
rect 3092 85072 4396 85112
rect 4436 85072 4445 85112
rect 4636 85072 4724 85112
rect 4684 85028 4724 85072
rect 6508 85072 7180 85112
rect 7220 85072 7229 85112
rect 7337 85072 7468 85112
rect 7508 85072 7517 85112
rect 7699 85072 7708 85112
rect 7748 85072 7756 85112
rect 7796 85072 7879 85112
rect 8419 85072 8428 85112
rect 8468 85072 8477 85112
rect 8611 85072 8620 85112
rect 8660 85072 9004 85112
rect 9044 85072 9053 85112
rect 12317 85072 12364 85112
rect 12404 85072 12413 85112
rect 12739 85072 12748 85112
rect 12788 85072 12844 85112
rect 12884 85072 12919 85112
rect 13420 85072 13996 85112
rect 14036 85072 14045 85112
rect 14188 85072 14612 85112
rect 6508 85028 6548 85072
rect 10252 85028 10292 85037
rect 11884 85028 11924 85037
rect 12364 85028 12404 85072
rect 13420 85028 13460 85072
rect 14188 85028 14228 85072
rect 14572 85028 14612 85072
rect 15148 85072 15284 85112
rect 15497 85072 15628 85112
rect 15668 85072 15677 85112
rect 15811 85072 15820 85112
rect 15860 85072 15869 85112
rect 15148 85028 15188 85072
rect 15820 85028 15860 85072
rect 16204 85028 16244 85037
rect 16876 85028 16916 85576
rect 17692 85532 17732 85576
rect 21510 85556 21600 85576
rect 17692 85492 18604 85532
rect 18644 85492 18653 85532
rect 18799 85408 18808 85448
rect 18848 85408 18890 85448
rect 18930 85408 18972 85448
rect 19012 85408 19054 85448
rect 19094 85408 19136 85448
rect 19176 85408 19185 85448
rect 17059 85156 17068 85196
rect 17108 85156 18740 85196
rect 18316 85028 18356 85037
rect 18700 85028 18740 85156
rect 21510 85112 21600 85132
rect 21283 85072 21292 85112
rect 21332 85072 21600 85112
rect 21510 85052 21600 85072
rect 19948 85028 19988 85037
rect 1411 84988 1420 85028
rect 1460 84988 1612 85028
rect 1652 84988 1661 85028
rect 2708 84988 2860 85028
rect 2900 84988 2909 85028
rect 3331 84988 3340 85028
rect 3380 84988 3436 85028
rect 3476 84988 4108 85028
rect 4148 84988 4157 85028
rect 5251 84988 5260 85028
rect 5300 84988 5548 85028
rect 5588 84988 5597 85028
rect 6874 84988 6883 85028
rect 6923 84988 7564 85028
rect 7604 84988 7613 85028
rect 7721 84988 7852 85028
rect 7892 84988 7901 85028
rect 8035 84988 8044 85028
rect 8084 84988 8215 85028
rect 8995 84988 9004 85028
rect 9044 84988 9292 85028
rect 9332 84988 9341 85028
rect 10121 84988 10252 85028
rect 10292 84988 10301 85028
rect 10505 84988 10636 85028
rect 10676 84988 10685 85028
rect 11753 84988 11884 85028
rect 11924 84988 11933 85028
rect 12346 84988 12355 85028
rect 12395 84988 12404 85028
rect 12451 84988 12460 85028
rect 12500 84988 12631 85028
rect 12809 84988 12940 85028
rect 12980 84988 12989 85028
rect 13899 84988 13908 85028
rect 13948 84988 14228 85028
rect 14275 84988 14284 85028
rect 14324 84988 14333 85028
rect 14563 84988 14572 85028
rect 14612 84988 14621 85028
rect 15130 84988 15139 85028
rect 15179 84988 15188 85028
rect 15235 84988 15244 85028
rect 15284 84988 15415 85028
rect 15593 84988 15724 85028
rect 15764 84988 15773 85028
rect 15820 84988 16204 85028
rect 16714 84988 16723 85028
rect 16763 84988 16916 85028
rect 17059 84988 17068 85028
rect 17108 84988 17117 85028
rect 18115 84988 18124 85028
rect 18164 84988 18316 85028
rect 18691 84988 18700 85028
rect 18740 84988 18749 85028
rect 19913 84988 19948 85028
rect 19988 84988 20044 85028
rect 20084 84988 20093 85028
rect 2668 84979 2708 84988
rect 4684 84979 4724 84988
rect 6508 84979 6548 84988
rect 10252 84979 10292 84988
rect 11884 84979 11924 84988
rect 13420 84979 13460 84988
rect 3283 84904 3292 84944
rect 3332 84904 3628 84944
rect 3668 84904 3677 84944
rect 7075 84904 7084 84944
rect 7124 84904 7133 84944
rect 7185 84904 7194 84944
rect 7234 84904 7660 84944
rect 7700 84904 7709 84944
rect 7939 84904 7948 84944
rect 7988 84904 8332 84944
rect 8372 84904 8381 84944
rect 2851 84820 2860 84860
rect 2900 84820 2956 84860
rect 2996 84820 3031 84860
rect 4780 84820 5684 84860
rect 6569 84820 6700 84860
rect 6740 84820 6749 84860
rect 6857 84820 6892 84860
rect 6932 84820 6979 84860
rect 7019 84820 7037 84860
rect 0 84776 90 84796
rect 0 84736 1420 84776
rect 1460 84736 1469 84776
rect 0 84716 90 84736
rect 4780 84692 4820 84820
rect 5644 84776 5684 84820
rect 7084 84776 7124 84904
rect 13917 84860 13957 84988
rect 14284 84944 14324 84988
rect 16204 84979 16244 84988
rect 17068 84944 17108 84988
rect 18316 84979 18356 84988
rect 19948 84979 19988 84988
rect 14179 84904 14188 84944
rect 14228 84904 14324 84944
rect 16588 84904 17108 84944
rect 16588 84860 16628 84904
rect 8131 84820 8140 84860
rect 8180 84820 9292 84860
rect 9332 84820 9341 84860
rect 10313 84820 10444 84860
rect 10484 84820 10493 84860
rect 12067 84820 12076 84860
rect 12116 84820 12940 84860
rect 12980 84820 13612 84860
rect 13652 84820 13957 84860
rect 14083 84820 14092 84860
rect 14132 84820 14668 84860
rect 14708 84820 14717 84860
rect 16099 84820 16108 84860
rect 16148 84820 16628 84860
rect 16745 84820 16876 84860
rect 16916 84820 16925 84860
rect 18377 84820 18508 84860
rect 18548 84820 18557 84860
rect 20131 84820 20140 84860
rect 20180 84820 20716 84860
rect 20756 84820 20765 84860
rect 5644 84736 6836 84776
rect 7084 84736 8524 84776
rect 8564 84736 8573 84776
rect 8899 84736 8908 84776
rect 8948 84736 11692 84776
rect 11732 84736 12460 84776
rect 12500 84736 12509 84776
rect 12940 84736 14036 84776
rect 6796 84692 6836 84736
rect 12940 84692 12980 84736
rect 3619 84652 3628 84692
rect 3668 84652 4820 84692
rect 4919 84652 4928 84692
rect 4968 84652 5010 84692
rect 5050 84652 5092 84692
rect 5132 84652 5174 84692
rect 5214 84652 5256 84692
rect 5296 84652 5305 84692
rect 6796 84652 12980 84692
rect 13996 84692 14036 84736
rect 13996 84652 15628 84692
rect 15668 84652 17932 84692
rect 17972 84652 17981 84692
rect 20039 84652 20048 84692
rect 20088 84652 20130 84692
rect 20170 84652 20212 84692
rect 20252 84652 20294 84692
rect 20334 84652 20376 84692
rect 20416 84652 20425 84692
rect 21510 84608 21600 84628
rect 172 84568 6028 84608
rect 6068 84568 6077 84608
rect 7459 84568 7468 84608
rect 7508 84568 8468 84608
rect 20899 84568 20908 84608
rect 20948 84568 21600 84608
rect 0 84440 90 84460
rect 172 84440 212 84568
rect 8428 84524 8468 84568
rect 21510 84548 21600 84568
rect 3628 84484 4436 84524
rect 4483 84484 4492 84524
rect 4532 84484 5548 84524
rect 5588 84484 5597 84524
rect 5731 84484 5740 84524
rect 5780 84484 6836 84524
rect 7651 84484 7660 84524
rect 7700 84484 7852 84524
rect 7892 84484 7901 84524
rect 8419 84484 8428 84524
rect 8468 84484 8477 84524
rect 9139 84484 9148 84524
rect 9188 84484 11980 84524
rect 12020 84484 12029 84524
rect 12233 84484 12364 84524
rect 12404 84484 12413 84524
rect 12739 84484 12748 84524
rect 12788 84484 13844 84524
rect 14249 84484 14380 84524
rect 14420 84484 14429 84524
rect 14755 84484 14764 84524
rect 14804 84484 14860 84524
rect 14900 84484 14935 84524
rect 16745 84484 16876 84524
rect 16916 84484 16925 84524
rect 16972 84484 19564 84524
rect 19604 84484 19613 84524
rect 0 84400 212 84440
rect 2179 84400 2188 84440
rect 2228 84400 2237 84440
rect 2717 84400 2764 84440
rect 2804 84400 2813 84440
rect 2860 84400 3340 84440
rect 3380 84400 3389 84440
rect 0 84380 90 84400
rect 2188 84356 2228 84400
rect 2764 84356 2804 84400
rect 2860 84356 2900 84400
rect 2188 84316 2612 84356
rect 2746 84316 2755 84356
rect 2795 84316 2804 84356
rect 2851 84316 2860 84356
rect 2900 84316 2909 84356
rect 3235 84316 3244 84356
rect 3284 84316 3436 84356
rect 3476 84316 3485 84356
rect 2572 84272 2612 84316
rect 259 84232 268 84272
rect 308 84232 1228 84272
rect 1268 84232 1277 84272
rect 1411 84232 1420 84272
rect 1460 84232 1612 84272
rect 1652 84232 1661 84272
rect 1987 84232 1996 84272
rect 2036 84232 2188 84272
rect 2228 84232 2237 84272
rect 2572 84232 2764 84272
rect 2804 84232 2813 84272
rect 3235 84232 3244 84272
rect 3284 84232 3340 84272
rect 3380 84232 3415 84272
rect 3628 84188 3668 84484
rect 3715 84316 3724 84356
rect 3764 84347 3895 84356
rect 3764 84316 3820 84347
rect 3860 84316 3895 84347
rect 4169 84316 4300 84356
rect 4340 84316 4349 84356
rect 3820 84298 3860 84307
rect 4300 84298 4340 84307
rect 835 84148 844 84188
rect 884 84148 3668 84188
rect 4396 84188 4436 84484
rect 5635 84400 5644 84440
rect 5684 84400 5692 84440
rect 5732 84400 5815 84440
rect 5932 84400 6700 84440
rect 6740 84400 6749 84440
rect 4675 84316 4684 84356
rect 4724 84316 5492 84356
rect 5452 84272 5492 84316
rect 5644 84272 5684 84400
rect 5932 84356 5972 84400
rect 6796 84356 6836 84484
rect 13804 84440 13844 84484
rect 16972 84440 17012 84484
rect 8323 84400 8332 84440
rect 8372 84400 8468 84440
rect 12931 84400 12940 84440
rect 12980 84400 13364 84440
rect 13577 84400 13708 84440
rect 13748 84400 13757 84440
rect 13804 84400 14174 84440
rect 14214 84400 14223 84440
rect 14266 84400 14275 84440
rect 14324 84400 14455 84440
rect 14659 84400 14668 84440
rect 14708 84400 14717 84440
rect 15148 84400 15340 84440
rect 15380 84400 15389 84440
rect 16579 84400 16588 84440
rect 16628 84400 17012 84440
rect 17836 84400 18508 84440
rect 18548 84400 18557 84440
rect 8428 84356 8468 84400
rect 13324 84356 13364 84400
rect 14668 84356 14708 84400
rect 15148 84356 15188 84400
rect 17836 84356 17876 84400
rect 5772 84316 5836 84356
rect 5876 84316 5923 84356
rect 5963 84316 5972 84356
rect 6019 84316 6028 84356
rect 6068 84316 6199 84356
rect 6403 84316 6412 84356
rect 6452 84316 6836 84356
rect 6979 84316 6988 84356
rect 7028 84316 7159 84356
rect 7337 84316 7468 84356
rect 7508 84316 7517 84356
rect 7817 84316 7852 84356
rect 7892 84316 7948 84356
rect 7988 84316 7997 84356
rect 8165 84316 8179 84356
rect 8219 84316 8228 84356
rect 8324 84316 8333 84356
rect 8373 84316 8468 84356
rect 8515 84316 8524 84356
rect 8564 84316 8695 84356
rect 8899 84316 8908 84356
rect 8948 84316 8957 84356
rect 9283 84316 9292 84356
rect 9332 84316 9772 84356
rect 9812 84316 9821 84356
rect 10243 84316 10252 84356
rect 10292 84347 10580 84356
rect 10292 84316 10540 84347
rect 6988 84298 7028 84307
rect 7468 84298 7508 84307
rect 4483 84232 4492 84272
rect 4532 84232 4684 84272
rect 4724 84232 4733 84272
rect 5059 84232 5068 84272
rect 5108 84232 5117 84272
rect 5443 84232 5452 84272
rect 5492 84232 5501 84272
rect 5644 84232 6508 84272
rect 6548 84232 6557 84272
rect 7651 84232 7660 84272
rect 7700 84232 7852 84272
rect 7892 84232 7901 84272
rect 8058 84232 8067 84272
rect 8107 84232 8116 84272
rect 5068 84188 5108 84232
rect 4396 84148 5108 84188
rect 5299 84148 5308 84188
rect 5348 84148 5644 84188
rect 5684 84148 5693 84188
rect 0 84104 90 84124
rect 8067 84104 8107 84232
rect 8165 84188 8205 84316
rect 8908 84272 8948 84316
rect 10627 84316 10636 84356
rect 10676 84316 10924 84356
rect 10964 84316 10973 84356
rect 11491 84316 11500 84356
rect 11540 84316 11884 84356
rect 11924 84347 12212 84356
rect 11924 84316 12172 84347
rect 10540 84272 10580 84307
rect 12547 84316 12556 84356
rect 12596 84316 12844 84356
rect 12884 84316 12893 84356
rect 13001 84316 13081 84356
rect 13121 84316 13132 84356
rect 13172 84316 13181 84356
rect 13315 84316 13324 84356
rect 13364 84316 13373 84356
rect 13594 84316 13603 84356
rect 13643 84316 14380 84356
rect 14420 84316 14429 84356
rect 12172 84298 12212 84307
rect 14473 84291 14482 84331
rect 14522 84291 14612 84331
rect 14659 84316 14668 84356
rect 14708 84316 14755 84356
rect 14851 84316 14860 84356
rect 14900 84316 15031 84356
rect 15130 84316 15139 84356
rect 15179 84316 15188 84356
rect 15235 84316 15244 84356
rect 15284 84316 15415 84356
rect 15497 84316 15628 84356
rect 15668 84316 15677 84356
rect 15811 84316 15820 84356
rect 15860 84347 16244 84356
rect 15860 84316 16204 84347
rect 8899 84232 8908 84272
rect 8948 84232 8995 84272
rect 10540 84232 10828 84272
rect 10868 84232 10877 84272
rect 12970 84263 13036 84272
rect 12970 84223 12979 84263
rect 13019 84232 13036 84263
rect 13076 84232 13159 84272
rect 13019 84223 13028 84232
rect 12970 84222 13028 84223
rect 14572 84188 14612 84291
rect 15593 84232 15724 84272
rect 15764 84232 15773 84272
rect 15820 84188 15860 84316
rect 16204 84298 16244 84307
rect 16684 84347 16972 84356
rect 16724 84316 16972 84347
rect 17012 84316 17021 84356
rect 17818 84316 17827 84356
rect 17867 84316 17876 84356
rect 17923 84316 17932 84356
rect 17972 84316 18103 84356
rect 18172 84316 18316 84356
rect 18356 84316 18365 84356
rect 18691 84316 18700 84356
rect 18740 84347 18932 84356
rect 18740 84316 18892 84347
rect 16684 84298 16724 84307
rect 18172 84272 18212 84316
rect 19241 84316 19372 84356
rect 19412 84316 19421 84356
rect 18892 84298 18932 84307
rect 19372 84298 19412 84307
rect 17059 84232 17068 84272
rect 17108 84232 17117 84272
rect 18115 84232 18124 84272
rect 18164 84232 18212 84272
rect 18316 84232 18412 84272
rect 18452 84232 18461 84272
rect 19747 84232 19756 84272
rect 19796 84232 19805 84272
rect 20009 84232 20140 84272
rect 20180 84232 20189 84272
rect 17068 84188 17108 84232
rect 18316 84188 18356 84232
rect 19756 84188 19796 84232
rect 8165 84148 8332 84188
rect 8372 84148 8381 84188
rect 8812 84148 11348 84188
rect 13987 84148 13996 84188
rect 14036 84148 14612 84188
rect 14659 84148 14668 84188
rect 14708 84148 15860 84188
rect 16291 84148 16300 84188
rect 16340 84148 17108 84188
rect 17731 84148 17740 84188
rect 17780 84148 18356 84188
rect 19363 84148 19372 84188
rect 19412 84148 19796 84188
rect 0 84064 1364 84104
rect 1459 84064 1468 84104
rect 1508 84064 1612 84104
rect 1652 84064 1661 84104
rect 1843 84064 1852 84104
rect 1892 84064 1900 84104
rect 1940 84064 2023 84104
rect 2227 84064 2236 84104
rect 2276 84064 3628 84104
rect 3668 84064 3677 84104
rect 4915 84064 4924 84104
rect 4964 84064 4973 84104
rect 8067 84064 8524 84104
rect 8564 84064 8573 84104
rect 0 84044 90 84064
rect 1324 84020 1364 84064
rect 4924 84020 4964 84064
rect 8812 84020 8852 84148
rect 11308 84104 11348 84148
rect 21510 84104 21600 84124
rect 1324 83980 2668 84020
rect 2708 83980 2717 84020
rect 2851 83980 2860 84020
rect 2900 83980 2909 84020
rect 4924 83980 8852 84020
rect 9004 84064 9148 84104
rect 9188 84064 9197 84104
rect 10723 84064 10732 84104
rect 10772 84064 11212 84104
rect 11252 84064 11261 84104
rect 11308 84064 13652 84104
rect 13699 84064 13708 84104
rect 13748 84064 14188 84104
rect 14228 84064 14237 84104
rect 17299 84064 17308 84104
rect 17348 84064 18356 84104
rect 19987 84064 19996 84104
rect 20036 84064 20044 84104
rect 20084 84064 20167 84104
rect 20371 84064 20380 84104
rect 20420 84064 20908 84104
rect 20948 84064 20957 84104
rect 21091 84064 21100 84104
rect 21140 84064 21600 84104
rect 0 83768 90 83788
rect 2860 83768 2900 83980
rect 3679 83896 3688 83936
rect 3728 83896 3770 83936
rect 3810 83896 3852 83936
rect 3892 83896 3934 83936
rect 3974 83896 4016 83936
rect 4056 83896 4065 83936
rect 9004 83852 9044 84064
rect 13612 84020 13652 84064
rect 18316 84020 18356 84064
rect 21510 84044 21600 84064
rect 13612 83980 16972 84020
rect 17012 83980 17260 84020
rect 17300 83980 17309 84020
rect 18316 83980 21292 84020
rect 21332 83980 21341 84020
rect 9283 83896 9292 83936
rect 9332 83896 12556 83936
rect 12596 83896 12605 83936
rect 18799 83896 18808 83936
rect 18848 83896 18890 83936
rect 18930 83896 18972 83936
rect 19012 83896 19054 83936
rect 19094 83896 19136 83936
rect 19176 83896 19185 83936
rect 7747 83812 7756 83852
rect 7796 83812 9044 83852
rect 11395 83812 11404 83852
rect 11444 83812 13420 83852
rect 13460 83812 13469 83852
rect 15715 83812 15724 83852
rect 15764 83812 18124 83852
rect 18164 83812 18356 83852
rect 0 83728 2764 83768
rect 2804 83728 2813 83768
rect 2860 83728 2996 83768
rect 3235 83728 3244 83768
rect 3284 83728 3820 83768
rect 3860 83728 3869 83768
rect 4387 83728 4396 83768
rect 4436 83728 5260 83768
rect 5300 83728 5308 83768
rect 5348 83728 5357 83768
rect 5875 83728 5884 83768
rect 5924 83728 6892 83768
rect 6932 83728 6941 83768
rect 7555 83728 7564 83768
rect 7604 83728 7660 83768
rect 7700 83728 7735 83768
rect 9331 83728 9340 83768
rect 9380 83728 12748 83768
rect 12788 83728 12797 83768
rect 13066 83728 13075 83768
rect 13115 83728 13996 83768
rect 14036 83728 14045 83768
rect 14803 83728 14812 83768
rect 14852 83728 16300 83768
rect 16340 83728 16349 83768
rect 17827 83728 17836 83768
rect 17876 83728 18260 83768
rect 0 83708 90 83728
rect 2764 83516 2804 83525
rect 2956 83516 2996 83728
rect 3043 83644 3052 83684
rect 3092 83644 3284 83684
rect 7459 83644 7468 83684
rect 7508 83644 8044 83684
rect 8084 83644 8093 83684
rect 9964 83644 10636 83684
rect 10676 83644 10685 83684
rect 11011 83644 11020 83684
rect 11060 83644 12500 83684
rect 12835 83644 12844 83684
rect 12884 83644 14228 83684
rect 14275 83644 14284 83684
rect 14324 83644 14333 83684
rect 14956 83644 16684 83684
rect 16724 83644 16733 83684
rect 16963 83644 16972 83684
rect 17012 83644 18124 83684
rect 18164 83644 18173 83684
rect 1507 83476 1516 83516
rect 1556 83476 1900 83516
rect 1940 83476 1949 83516
rect 2633 83476 2764 83516
rect 2804 83476 2996 83516
rect 3244 83516 3284 83644
rect 3427 83560 3436 83600
rect 3476 83560 3916 83600
rect 3956 83560 3965 83600
rect 5539 83560 5548 83600
rect 5588 83560 6988 83600
rect 7028 83560 7037 83600
rect 8515 83560 8524 83600
rect 8564 83560 8908 83600
rect 8948 83560 8957 83600
rect 9004 83560 9100 83600
rect 9140 83560 9149 83600
rect 4492 83516 4532 83525
rect 7276 83516 7316 83525
rect 3244 83476 3427 83516
rect 3467 83476 3476 83516
rect 3523 83476 3532 83516
rect 3572 83476 3581 83516
rect 3715 83476 3724 83516
rect 3764 83476 4012 83516
rect 4052 83476 4061 83516
rect 4387 83476 4396 83516
rect 4436 83476 4492 83516
rect 4532 83476 4567 83516
rect 4771 83476 4780 83516
rect 4820 83476 4980 83516
rect 5020 83476 5029 83516
rect 5705 83476 5740 83516
rect 5780 83476 5836 83516
rect 5876 83476 5972 83516
rect 6019 83476 6028 83516
rect 6068 83476 6796 83516
rect 6836 83476 6845 83516
rect 7459 83476 7468 83516
rect 7508 83507 8084 83516
rect 7508 83476 8044 83507
rect 2764 83467 2804 83476
rect 0 83432 90 83452
rect 3532 83432 3572 83476
rect 4492 83467 4532 83476
rect 0 83392 1036 83432
rect 1076 83392 1085 83432
rect 3331 83392 3340 83432
rect 3380 83392 3572 83432
rect 0 83372 90 83392
rect 5932 83348 5972 83476
rect 7276 83432 7316 83476
rect 8201 83476 8332 83516
rect 8372 83476 8567 83516
rect 8607 83476 8616 83516
rect 8698 83476 8707 83516
rect 8747 83476 8756 83516
rect 8803 83476 8812 83516
rect 8852 83476 8861 83516
rect 8044 83458 8084 83467
rect 8716 83432 8756 83476
rect 7276 83392 7372 83432
rect 7412 83392 7421 83432
rect 7651 83392 7660 83432
rect 7700 83392 7948 83432
rect 7988 83392 7997 83432
rect 8515 83392 8524 83432
rect 8564 83392 8756 83432
rect 8812 83348 8852 83476
rect 2947 83308 2956 83348
rect 2996 83308 3127 83348
rect 5155 83308 5164 83348
rect 5204 83308 5684 83348
rect 5932 83308 8852 83348
rect 5644 83180 5684 83308
rect 9004 83264 9044 83560
rect 9964 83516 10004 83644
rect 11203 83560 11212 83600
rect 11252 83560 11261 83600
rect 11779 83560 11788 83600
rect 11828 83560 11980 83600
rect 12020 83560 12029 83600
rect 10828 83516 10868 83525
rect 11212 83516 11252 83560
rect 12364 83516 12404 83525
rect 9571 83476 9580 83516
rect 9620 83476 9629 83516
rect 9955 83476 9964 83516
rect 10004 83476 10013 83516
rect 10697 83476 10828 83516
rect 10868 83476 10877 83516
rect 11212 83476 11278 83516
rect 11318 83476 11327 83516
rect 11395 83476 11404 83516
rect 11444 83476 11575 83516
rect 11683 83476 11692 83516
rect 11732 83476 11884 83516
rect 11924 83476 11933 83516
rect 12067 83476 12076 83516
rect 12116 83476 12364 83516
rect 12460 83516 12500 83644
rect 14188 83600 14228 83644
rect 14284 83600 14324 83644
rect 14956 83600 14996 83644
rect 12547 83560 12556 83600
rect 12596 83560 13556 83600
rect 13603 83560 13612 83600
rect 13652 83560 13661 83600
rect 13843 83560 13852 83600
rect 13892 83560 13900 83600
rect 13940 83560 14023 83600
rect 14179 83560 14188 83600
rect 14228 83560 14237 83600
rect 14284 83560 14524 83600
rect 14564 83560 14573 83600
rect 14620 83560 14996 83600
rect 15043 83560 15052 83600
rect 15092 83560 15676 83600
rect 15716 83560 15725 83600
rect 15907 83560 15916 83600
rect 15956 83560 16087 83600
rect 17452 83560 17836 83600
rect 17876 83560 17885 83600
rect 12460 83476 12852 83516
rect 12892 83476 12901 83516
rect 7372 83224 9044 83264
rect 76 83140 652 83180
rect 692 83140 701 83180
rect 4919 83140 4928 83180
rect 4968 83140 5010 83180
rect 5050 83140 5092 83180
rect 5132 83140 5174 83180
rect 5214 83140 5256 83180
rect 5296 83140 5305 83180
rect 5635 83140 5644 83180
rect 5684 83140 5693 83180
rect 76 83116 116 83140
rect 0 83056 116 83116
rect 7372 83096 7412 83224
rect 9580 83180 9620 83476
rect 10828 83467 10868 83476
rect 12268 83432 12308 83476
rect 12364 83467 12404 83476
rect 13516 83432 13556 83560
rect 13612 83516 13652 83560
rect 14620 83516 14660 83560
rect 17356 83516 17396 83525
rect 17452 83516 17492 83560
rect 18220 83516 18260 83728
rect 18316 83600 18356 83812
rect 18979 83728 18988 83768
rect 19028 83728 19603 83768
rect 19643 83728 19652 83768
rect 21187 83728 21196 83768
rect 21236 83728 21428 83768
rect 18691 83644 18700 83684
rect 18740 83644 18749 83684
rect 19555 83644 19564 83684
rect 19604 83644 19756 83684
rect 19796 83644 19805 83684
rect 18307 83560 18316 83600
rect 18356 83560 18365 83600
rect 18700 83516 18740 83644
rect 21388 83600 21428 83728
rect 21510 83600 21600 83620
rect 19660 83560 19852 83600
rect 19892 83560 19901 83600
rect 20009 83560 20140 83600
rect 20180 83560 20189 83600
rect 20371 83560 20380 83600
rect 20420 83560 21196 83600
rect 21236 83560 21245 83600
rect 21388 83560 21600 83600
rect 18892 83516 18932 83525
rect 19660 83516 19700 83560
rect 21510 83540 21600 83560
rect 13612 83476 14660 83516
rect 14860 83476 14947 83516
rect 14987 83476 14996 83516
rect 15249 83476 15258 83516
rect 15298 83476 15820 83516
rect 15860 83476 15869 83516
rect 16003 83476 16012 83516
rect 16052 83476 16108 83516
rect 16148 83476 16183 83516
rect 17225 83476 17260 83516
rect 17300 83476 17356 83516
rect 17396 83476 17492 83516
rect 17548 83476 17827 83516
rect 17867 83476 17876 83516
rect 17923 83476 17932 83516
rect 17972 83476 18103 83516
rect 18220 83476 18412 83516
rect 18452 83476 18461 83516
rect 18604 83476 18892 83516
rect 19402 83476 19411 83516
rect 19451 83476 19700 83516
rect 19747 83476 19756 83516
rect 19796 83476 19805 83516
rect 19939 83476 19948 83516
rect 19988 83476 19997 83516
rect 12259 83392 12268 83432
rect 12308 83392 12317 83432
rect 13516 83392 13948 83432
rect 13988 83392 13997 83432
rect 8035 83140 8044 83180
rect 8084 83140 8428 83180
rect 8468 83140 9620 83180
rect 4387 83056 4396 83096
rect 4436 83056 4684 83096
rect 4724 83056 4733 83096
rect 4876 83056 7412 83096
rect 13795 83056 13804 83096
rect 13844 83056 14420 83096
rect 0 83036 90 83056
rect 4876 83012 4916 83056
rect 172 82972 4916 83012
rect 4963 82972 4972 83012
rect 5012 82972 5143 83012
rect 7555 82972 7564 83012
rect 7604 82972 8332 83012
rect 8372 82972 8428 83012
rect 8468 82972 8503 83012
rect 13123 82972 13132 83012
rect 13172 82972 14284 83012
rect 14324 82972 14333 83012
rect 172 82928 212 82972
rect 14380 82928 14420 83056
rect 14476 83056 14764 83096
rect 14804 83056 14813 83096
rect 14476 83012 14516 83056
rect 14860 83012 14900 83476
rect 17356 83467 17396 83476
rect 17548 83432 17588 83476
rect 15043 83392 15052 83432
rect 15092 83392 15223 83432
rect 17539 83392 17548 83432
rect 17588 83392 17597 83432
rect 18604 83348 18644 83476
rect 18892 83467 18932 83476
rect 19756 83432 19796 83476
rect 19948 83432 19988 83476
rect 19075 83392 19084 83432
rect 19124 83392 19796 83432
rect 19843 83392 19852 83432
rect 19892 83392 19988 83432
rect 15139 83308 15148 83348
rect 15188 83308 15197 83348
rect 15331 83308 15340 83348
rect 15380 83308 18644 83348
rect 15148 83012 15188 83308
rect 20039 83140 20048 83180
rect 20088 83140 20130 83180
rect 20170 83140 20212 83180
rect 20252 83140 20294 83180
rect 20334 83140 20376 83180
rect 20416 83140 20425 83180
rect 21510 83096 21600 83116
rect 21379 83056 21388 83096
rect 21428 83056 21600 83096
rect 21510 83036 21600 83056
rect 14467 82972 14476 83012
rect 14516 82972 14525 83012
rect 14860 82972 14908 83012
rect 14948 82972 14957 83012
rect 15148 82972 16532 83012
rect 17731 82972 17740 83012
rect 17780 82972 20180 83012
rect 76 82888 212 82928
rect 2633 82888 2764 82928
rect 2804 82888 4436 82928
rect 76 82780 116 82888
rect 1507 82804 1516 82844
rect 1556 82804 1565 82844
rect 2764 82835 2804 82888
rect 0 82720 116 82780
rect 0 82700 90 82720
rect 1516 82676 1556 82804
rect 2851 82804 2860 82844
rect 2900 82804 3235 82844
rect 3275 82804 3284 82844
rect 3331 82804 3340 82844
rect 3380 82804 3511 82844
rect 3715 82804 3724 82844
rect 3764 82804 3773 82844
rect 4169 82804 4300 82844
rect 4340 82804 4349 82844
rect 2764 82786 2804 82795
rect 3724 82760 3764 82804
rect 4300 82786 4340 82795
rect 3523 82720 3532 82760
rect 3572 82720 3764 82760
rect 3820 82720 3859 82760
rect 3899 82720 4204 82760
rect 4244 82720 4253 82760
rect 3820 82676 3860 82720
rect 4396 82676 4436 82888
rect 4780 82888 5164 82928
rect 5204 82888 5213 82928
rect 6988 82888 13076 82928
rect 4780 82835 4820 82888
rect 6988 82844 7028 82888
rect 4780 82786 4820 82795
rect 5356 82835 5396 82844
rect 6211 82804 6220 82844
rect 6260 82804 6604 82844
rect 6644 82804 6653 82844
rect 6979 82804 6988 82844
rect 7028 82804 7037 82844
rect 7363 82804 7372 82844
rect 7412 82835 8564 82844
rect 7412 82804 8236 82835
rect 5356 82676 5396 82795
rect 1516 82636 2764 82676
rect 2804 82636 3244 82676
rect 3284 82636 3293 82676
rect 3792 82636 3820 82676
rect 3860 82636 3869 82676
rect 4396 82636 5396 82676
rect 6604 82676 6644 82804
rect 8276 82804 8564 82835
rect 8611 82804 8620 82844
rect 8660 82804 8669 82844
rect 9868 82835 10252 82844
rect 8236 82786 8276 82795
rect 8524 82760 8564 82804
rect 8515 82720 8524 82760
rect 8564 82720 8573 82760
rect 8620 82676 8660 82804
rect 9908 82804 10252 82835
rect 10292 82804 10301 82844
rect 10435 82804 10444 82844
rect 10484 82804 11395 82844
rect 11435 82804 11444 82844
rect 11491 82804 11500 82844
rect 11540 82804 11549 82844
rect 11779 82804 11788 82844
rect 11828 82804 11884 82844
rect 11924 82804 11980 82844
rect 12020 82804 12084 82844
rect 12259 82804 12268 82844
rect 12308 82835 12500 82844
rect 12308 82804 12460 82835
rect 9868 82786 9908 82795
rect 11500 82760 11540 82804
rect 12739 82804 12748 82844
rect 12788 82835 12980 82844
rect 12788 82804 12940 82835
rect 12460 82786 12500 82795
rect 12940 82786 12980 82795
rect 11395 82720 11404 82760
rect 11444 82720 11540 82760
rect 11683 82720 11692 82760
rect 11732 82720 11980 82760
rect 12020 82720 12029 82760
rect 13036 82676 13076 82888
rect 13708 82888 14764 82928
rect 14804 82888 14813 82928
rect 15148 82888 15668 82928
rect 16003 82888 16012 82928
rect 16052 82888 16340 82928
rect 13708 82760 13748 82888
rect 15148 82844 15188 82888
rect 15628 82844 15668 82888
rect 16300 82844 16340 82888
rect 16492 82844 16532 82972
rect 16876 82888 19988 82928
rect 16876 82844 16916 82888
rect 19948 82844 19988 82888
rect 13795 82804 13804 82844
rect 13844 82804 14572 82844
rect 14612 82804 14621 82844
rect 14800 82804 14809 82844
rect 14849 82804 15188 82844
rect 15235 82804 15244 82844
rect 15284 82804 15293 82844
rect 15340 82804 15353 82844
rect 15393 82804 15427 82844
rect 15497 82804 15628 82844
rect 15668 82804 15677 82844
rect 15785 82804 15916 82844
rect 15956 82804 15965 82844
rect 16099 82804 16108 82844
rect 16148 82804 16244 82844
rect 16291 82804 16300 82844
rect 16340 82804 16349 82844
rect 16483 82804 16492 82844
rect 16532 82804 16541 82844
rect 16867 82804 16876 82844
rect 16916 82804 16972 82844
rect 17012 82804 17076 82844
rect 17731 82804 17740 82844
rect 17780 82835 18164 82844
rect 17780 82804 18124 82835
rect 15244 82760 15284 82804
rect 15340 82760 15380 82804
rect 16204 82760 16244 82804
rect 18499 82804 18508 82844
rect 18548 82835 18740 82844
rect 18548 82804 18700 82835
rect 18124 82786 18164 82795
rect 19939 82804 19948 82844
rect 19988 82804 19997 82844
rect 18700 82786 18740 82795
rect 20140 82760 20180 82972
rect 13411 82720 13420 82760
rect 13460 82720 13748 82760
rect 13961 82720 14092 82760
rect 14132 82720 14141 82760
rect 14659 82720 14668 82760
rect 14731 82720 14839 82760
rect 15139 82720 15148 82760
rect 15188 82720 15284 82760
rect 15331 82720 15340 82760
rect 15380 82720 15389 82760
rect 16195 82720 16204 82760
rect 16244 82720 16253 82760
rect 20131 82720 20140 82760
rect 20180 82720 20189 82760
rect 6604 82636 8428 82676
rect 8468 82636 8660 82676
rect 13027 82636 13036 82676
rect 13076 82636 13085 82676
rect 13651 82636 13660 82676
rect 13700 82636 14284 82676
rect 14324 82636 14333 82676
rect 16003 82636 16012 82676
rect 16052 82636 16300 82676
rect 16340 82636 16349 82676
rect 20371 82636 20380 82676
rect 20420 82636 21100 82676
rect 21140 82636 21149 82676
rect 21510 82592 21600 82612
rect 2947 82552 2956 82592
rect 2996 82552 4300 82592
rect 4340 82552 4349 82592
rect 6115 82552 6124 82592
rect 6164 82552 6796 82592
rect 6836 82552 6845 82592
rect 10051 82552 10060 82592
rect 10100 82552 12556 82592
rect 12596 82552 12605 82592
rect 14323 82552 14332 82592
rect 14372 82552 14381 82592
rect 18185 82552 18316 82592
rect 18356 82552 18365 82592
rect 18499 82552 18508 82592
rect 18548 82552 18679 82592
rect 20140 82552 21600 82592
rect 14332 82508 14372 82552
rect 20140 82508 20180 82552
rect 21510 82532 21600 82552
rect 2860 82468 6508 82508
rect 6548 82468 6557 82508
rect 14332 82468 20180 82508
rect 0 82424 90 82444
rect 2860 82424 2900 82468
rect 0 82384 2900 82424
rect 3679 82384 3688 82424
rect 3728 82384 3770 82424
rect 3810 82384 3852 82424
rect 3892 82384 3934 82424
rect 3974 82384 4016 82424
rect 4056 82384 4065 82424
rect 6883 82384 6892 82424
rect 6932 82384 14956 82424
rect 14996 82384 15005 82424
rect 18799 82384 18808 82424
rect 18848 82384 18890 82424
rect 18930 82384 18972 82424
rect 19012 82384 19054 82424
rect 19094 82384 19136 82424
rect 19176 82384 19185 82424
rect 0 82364 90 82384
rect 643 82300 652 82340
rect 692 82300 1420 82340
rect 1460 82300 1469 82340
rect 1891 82300 1900 82340
rect 1940 82300 16492 82340
rect 16532 82300 16541 82340
rect 1027 82216 1036 82256
rect 1076 82216 4396 82256
rect 4436 82216 4445 82256
rect 7267 82216 7276 82256
rect 7316 82216 8140 82256
rect 8180 82216 8189 82256
rect 13027 82216 13036 82256
rect 13076 82216 13660 82256
rect 13700 82216 13709 82256
rect 14371 82216 14380 82256
rect 14420 82216 15148 82256
rect 15188 82216 15197 82256
rect 2755 82132 2764 82172
rect 2804 82132 4436 82172
rect 6595 82132 6604 82172
rect 6644 82132 7468 82172
rect 7508 82132 7517 82172
rect 7564 82132 8084 82172
rect 13795 82132 13804 82172
rect 13844 82132 16436 82172
rect 0 82088 90 82108
rect 4396 82088 4436 82132
rect 7564 82088 7604 82132
rect 0 82048 1420 82088
rect 1460 82048 1469 82088
rect 2851 82048 2860 82088
rect 2900 82048 3628 82088
rect 3668 82048 3724 82088
rect 3764 82048 3773 82088
rect 4003 82048 4012 82088
rect 4052 82048 4340 82088
rect 4396 82048 5204 82088
rect 6499 82048 6508 82088
rect 6548 82048 7604 82088
rect 7660 82048 7988 82088
rect 0 82028 90 82048
rect 2764 82004 2804 82013
rect 4300 82004 4340 82048
rect 5164 82004 5204 82048
rect 6412 82004 6452 82013
rect 6988 82004 7028 82048
rect 1507 81964 1516 82004
rect 1556 81964 1996 82004
rect 2036 81964 2476 82004
rect 2516 81964 2525 82004
rect 2947 81964 2956 82004
rect 2996 81964 3235 82004
rect 3275 81964 3284 82004
rect 3331 81964 3340 82004
rect 3380 81964 3511 82004
rect 3811 81964 3820 82004
rect 3860 81964 3991 82004
rect 4387 81964 4396 82004
rect 4436 81964 4788 82004
rect 4828 81964 4837 82004
rect 5155 81964 5164 82004
rect 5204 81964 5213 82004
rect 5347 81964 5356 82004
rect 5396 81964 6412 82004
rect 6612 81964 6700 82004
rect 6740 81964 6743 82004
rect 6783 81964 6792 82004
rect 6874 81964 6883 82004
rect 6923 81964 6932 82004
rect 6979 81964 6988 82004
rect 7028 81964 7037 82004
rect 7145 81964 7276 82004
rect 7316 81964 7325 82004
rect 7433 81964 7564 82004
rect 7604 81964 7613 82004
rect 2764 81920 2804 81964
rect 3340 81920 3380 81964
rect 4300 81955 4340 81964
rect 6412 81955 6452 81964
rect 6892 81920 6932 81964
rect 7660 81920 7700 82048
rect 7948 82004 7988 82048
rect 7747 81964 7756 82004
rect 7796 81964 7805 82004
rect 7930 81964 7939 82004
rect 7979 81964 7988 82004
rect 8044 82004 8084 82132
rect 8297 82048 8428 82088
rect 8468 82048 8477 82088
rect 8611 82048 8620 82088
rect 8660 82048 8908 82088
rect 8948 82048 8957 82088
rect 9091 82048 9100 82088
rect 9140 82048 9332 82088
rect 11657 82048 11692 82088
rect 11732 82048 11788 82088
rect 11828 82048 11837 82088
rect 13385 82048 13420 82088
rect 13460 82048 13516 82088
rect 13556 82048 13565 82088
rect 14249 82048 14380 82088
rect 14420 82048 14429 82088
rect 15043 82048 15052 82088
rect 15092 82048 16252 82088
rect 16292 82048 16301 82088
rect 9292 82004 9332 82048
rect 10540 82004 10580 82013
rect 12268 82004 12308 82013
rect 14956 82004 14996 82013
rect 16396 82004 16436 82132
rect 21510 82088 21600 82108
rect 18115 82048 18124 82088
rect 18164 82048 18892 82088
rect 18932 82048 18941 82088
rect 21388 82048 21600 82088
rect 17836 82004 17876 82013
rect 19468 82004 19508 82013
rect 8044 81964 9100 82004
rect 9140 81964 9149 82004
rect 9283 81964 9292 82004
rect 9332 81964 9964 82004
rect 10004 81964 10013 82004
rect 10243 81964 10252 82004
rect 10292 81964 10540 82004
rect 2764 81880 3148 81920
rect 3188 81880 3197 81920
rect 3340 81880 3724 81920
rect 3764 81880 3773 81920
rect 6892 81880 6988 81920
rect 7028 81880 7037 81920
rect 7171 81880 7180 81920
rect 7220 81880 7700 81920
rect 2947 81796 2956 81836
rect 2996 81796 3436 81836
rect 3476 81796 3485 81836
rect 4841 81796 4972 81836
rect 5012 81796 5021 81836
rect 6953 81796 7075 81836
rect 7124 81796 7133 81836
rect 0 81752 90 81772
rect 0 81712 76 81752
rect 116 81712 125 81752
rect 0 81692 90 81712
rect 7756 81668 7796 81964
rect 7843 81880 7852 81920
rect 7892 81880 8428 81920
rect 8468 81880 8477 81920
rect 8851 81880 8860 81920
rect 8900 81880 10484 81920
rect 8179 81796 8188 81836
rect 8228 81796 8332 81836
rect 8372 81796 8381 81836
rect 8947 81796 8956 81836
rect 8996 81796 9005 81836
rect 8956 81752 8996 81796
rect 7843 81712 7852 81752
rect 7892 81712 8996 81752
rect 10444 81752 10484 81880
rect 10540 81836 10580 81964
rect 10732 81964 11203 82004
rect 11243 81964 11252 82004
rect 11299 81964 11308 82004
rect 11348 81964 11404 82004
rect 11444 81964 11479 82004
rect 11683 81964 11692 82004
rect 11732 81964 11788 82004
rect 11828 81964 11863 82004
rect 12233 81964 12268 82004
rect 12308 81964 12364 82004
rect 12404 81964 12413 82004
rect 12547 81964 12556 82004
rect 12596 81964 12756 82004
rect 12796 81964 12805 82004
rect 13027 81964 13036 82004
rect 13076 81964 13804 82004
rect 13844 81964 13891 82004
rect 13931 81964 13940 82004
rect 13987 81964 13996 82004
rect 14036 81964 14092 82004
rect 14132 81964 14167 82004
rect 14345 81964 14476 82004
rect 14516 81964 14525 82004
rect 14825 81964 14956 82004
rect 14996 81964 15005 82004
rect 15331 81964 15340 82004
rect 15380 81964 15444 82004
rect 15484 81964 15628 82004
rect 15668 81964 15811 82004
rect 15851 81964 15860 82004
rect 15977 81964 16012 82004
rect 16052 81964 16108 82004
rect 16148 81964 16157 82004
rect 16387 81964 16396 82004
rect 16436 81964 16445 82004
rect 16553 81964 16588 82004
rect 16628 81964 16684 82004
rect 16724 81964 16916 82004
rect 16963 81964 16972 82004
rect 17012 81964 17836 82004
rect 18251 81964 18316 82004
rect 18356 81964 18382 82004
rect 18422 81964 18431 82004
rect 18504 81964 18513 82004
rect 18553 81964 18562 82004
rect 18857 81964 18988 82004
rect 19028 81964 19037 82004
rect 19171 81964 19180 82004
rect 19220 81964 19468 82004
rect 19651 81964 19660 82004
rect 19700 81964 19956 82004
rect 19996 81964 20005 82004
rect 10732 81920 10772 81964
rect 12268 81955 12308 81964
rect 14956 81920 14996 81964
rect 16876 81920 16916 81964
rect 17836 81955 17876 81964
rect 18508 81920 18548 81964
rect 19468 81955 19508 81964
rect 10723 81880 10732 81920
rect 10772 81880 10781 81920
rect 13987 81880 13996 81920
rect 14036 81880 14996 81920
rect 16003 81880 16012 81920
rect 16052 81880 16780 81920
rect 16820 81880 16829 81920
rect 16876 81880 17068 81920
rect 17108 81880 17117 81920
rect 18316 81880 18548 81920
rect 21388 81920 21428 82048
rect 21510 82028 21600 82048
rect 21388 81880 21524 81920
rect 18316 81836 18356 81880
rect 21484 81836 21524 81880
rect 10540 81796 11884 81836
rect 11924 81796 11933 81836
rect 12931 81796 12940 81836
rect 12980 81796 12989 81836
rect 13420 81796 13660 81836
rect 13700 81796 13709 81836
rect 15619 81796 15628 81836
rect 15668 81796 15916 81836
rect 15956 81796 15965 81836
rect 18019 81796 18028 81836
rect 18068 81796 18077 81836
rect 18307 81796 18316 81836
rect 18356 81796 18365 81836
rect 20131 81796 20140 81836
rect 20180 81796 21388 81836
rect 21428 81796 21437 81836
rect 21484 81796 21575 81836
rect 10444 81712 10732 81752
rect 10772 81712 10781 81752
rect 4919 81628 4928 81668
rect 4968 81628 5010 81668
rect 5050 81628 5092 81668
rect 5132 81628 5174 81668
rect 5214 81628 5256 81668
rect 5296 81628 5305 81668
rect 7459 81628 7468 81668
rect 7508 81628 7796 81668
rect 4553 81460 4636 81500
rect 4676 81460 4684 81500
rect 4724 81460 4733 81500
rect 6595 81460 6604 81500
rect 6644 81460 7180 81500
rect 7220 81460 7229 81500
rect 7721 81460 7843 81500
rect 7892 81460 7901 81500
rect 8851 81460 8860 81500
rect 8900 81460 9484 81500
rect 9524 81460 9533 81500
rect 10348 81460 10828 81500
rect 10868 81460 10972 81500
rect 11012 81460 11021 81500
rect 0 81416 90 81436
rect 0 81376 172 81416
rect 212 81376 221 81416
rect 2467 81376 2476 81416
rect 2516 81376 4108 81416
rect 4148 81376 4157 81416
rect 4876 81376 5836 81416
rect 5876 81376 6412 81416
rect 6452 81376 6461 81416
rect 7267 81376 7276 81416
rect 7316 81376 7660 81416
rect 7700 81376 7709 81416
rect 7939 81376 7948 81416
rect 7988 81376 8276 81416
rect 0 81356 90 81376
rect 2476 81332 2516 81376
rect 4876 81332 4916 81376
rect 8236 81332 8276 81376
rect 1603 81292 1612 81332
rect 1652 81292 2516 81332
rect 2729 81292 2860 81332
rect 2900 81292 2909 81332
rect 3523 81292 3532 81332
rect 3572 81292 3764 81332
rect 3811 81292 3820 81332
rect 3860 81292 4676 81332
rect 4858 81292 4867 81332
rect 4907 81292 4916 81332
rect 4963 81292 4972 81332
rect 5012 81292 5143 81332
rect 5225 81292 5356 81332
rect 5396 81292 5405 81332
rect 5801 81292 5932 81332
rect 5972 81292 6124 81332
rect 6164 81292 6173 81332
rect 6412 81323 6700 81332
rect 2860 81274 2900 81283
rect 3724 81248 3764 81292
rect 4636 81248 4676 81292
rect 5356 81248 5396 81292
rect 5932 81274 5972 81283
rect 6452 81292 6700 81323
rect 6740 81292 6892 81332
rect 6932 81292 6941 81332
rect 7049 81292 7171 81332
rect 7220 81292 7372 81332
rect 7412 81292 7421 81332
rect 7564 81292 7747 81332
rect 7787 81292 7796 81332
rect 7843 81292 7852 81332
rect 7892 81292 8055 81332
rect 8095 81292 8104 81332
rect 8227 81292 8236 81332
rect 8276 81292 8285 81332
rect 8410 81292 8419 81332
rect 8468 81292 8599 81332
rect 8803 81292 8812 81332
rect 8852 81292 9100 81332
rect 9140 81292 9149 81332
rect 10348 81323 10388 81460
rect 12940 81416 12980 81796
rect 13420 81584 13460 81796
rect 18028 81752 18068 81796
rect 21535 81752 21575 81796
rect 13507 81712 13516 81752
rect 13556 81712 15724 81752
rect 15764 81712 15773 81752
rect 18019 81712 18028 81752
rect 18068 81712 18115 81752
rect 18595 81712 18604 81752
rect 18644 81712 21575 81752
rect 20039 81628 20048 81668
rect 20088 81628 20130 81668
rect 20170 81628 20212 81668
rect 20252 81628 20294 81668
rect 20334 81628 20376 81668
rect 20416 81628 20425 81668
rect 21510 81584 21600 81604
rect 13420 81544 18164 81584
rect 18211 81544 18220 81584
rect 18260 81544 21600 81584
rect 13027 81460 13036 81500
rect 13076 81460 14860 81500
rect 14900 81460 14909 81500
rect 15811 81460 15820 81500
rect 15860 81460 17059 81500
rect 17099 81460 17108 81500
rect 17417 81460 17500 81500
rect 17540 81460 17548 81500
rect 17588 81460 17597 81500
rect 18124 81416 18164 81544
rect 21510 81524 21600 81544
rect 19075 81460 19084 81500
rect 19124 81460 20140 81500
rect 20180 81460 20189 81500
rect 10531 81376 10540 81416
rect 10580 81376 11348 81416
rect 12940 81376 14668 81416
rect 14708 81376 14717 81416
rect 14947 81376 14956 81416
rect 14996 81376 16204 81416
rect 16244 81376 17012 81416
rect 18124 81376 18220 81416
rect 18260 81376 18269 81416
rect 18412 81376 18508 81416
rect 18548 81376 18557 81416
rect 11308 81332 11348 81376
rect 16972 81332 17012 81376
rect 18412 81332 18452 81376
rect 6412 81274 6452 81283
rect 67 81208 76 81248
rect 116 81208 1228 81248
rect 1268 81208 1277 81248
rect 3113 81208 3244 81248
rect 3284 81208 3293 81248
rect 3497 81208 3628 81248
rect 3668 81208 3677 81248
rect 3724 81208 3964 81248
rect 4004 81208 4013 81248
rect 4099 81208 4108 81248
rect 4148 81208 4204 81248
rect 4244 81208 4279 81248
rect 4387 81208 4396 81248
rect 4436 81208 4567 81248
rect 4636 81208 5396 81248
rect 5443 81208 5452 81248
rect 5492 81208 5501 81248
rect 5452 81164 5492 81208
rect 7564 81164 7604 81292
rect 11290 81292 11299 81332
rect 11339 81292 11348 81332
rect 11395 81292 11404 81332
rect 11444 81292 11575 81332
rect 11657 81292 11788 81332
rect 11828 81292 11837 81332
rect 12233 81292 12364 81332
rect 12404 81292 12413 81332
rect 12460 81323 12884 81332
rect 12460 81292 12844 81323
rect 10348 81274 10388 81283
rect 12364 81274 12404 81283
rect 8428 81208 8620 81248
rect 8660 81208 8669 81248
rect 10435 81208 10444 81248
rect 10484 81208 10732 81248
rect 10772 81208 10781 81248
rect 11683 81208 11692 81248
rect 11732 81208 11884 81248
rect 11924 81208 11933 81248
rect 8428 81164 8468 81208
rect 3708 81124 3724 81164
rect 3764 81124 3868 81164
rect 3908 81124 5492 81164
rect 7555 81124 7564 81164
rect 7604 81124 7613 81164
rect 8410 81124 8419 81164
rect 8459 81124 8468 81164
rect 0 81080 90 81100
rect 12460 81080 12500 81292
rect 13507 81292 13516 81332
rect 13556 81292 13708 81332
rect 13748 81292 13757 81332
rect 14633 81292 14764 81332
rect 14804 81292 14813 81332
rect 15340 81323 15380 81332
rect 12844 81274 12884 81283
rect 14764 81274 14804 81283
rect 15715 81292 15724 81332
rect 15764 81292 16588 81332
rect 16628 81292 16637 81332
rect 16963 81292 16972 81332
rect 17012 81292 17021 81332
rect 18394 81292 18403 81332
rect 18443 81292 18452 81332
rect 18499 81292 18508 81332
rect 18548 81292 18604 81332
rect 18644 81292 18679 81332
rect 18761 81292 18892 81332
rect 18932 81292 18941 81332
rect 19171 81292 19180 81332
rect 19220 81323 19508 81332
rect 19220 81292 19468 81323
rect 15340 81164 15380 81283
rect 14371 81124 14380 81164
rect 14420 81124 15380 81164
rect 16684 81250 16732 81290
rect 16772 81250 16781 81290
rect 16684 81164 16724 81250
rect 16858 81208 16867 81248
rect 16907 81208 17260 81248
rect 17300 81208 17309 81248
rect 17731 81208 17740 81248
rect 17780 81208 17789 81248
rect 17923 81208 17932 81248
rect 17972 81208 18103 81248
rect 18499 81208 18508 81248
rect 18548 81208 18988 81248
rect 19028 81208 19037 81248
rect 17740 81164 17780 81208
rect 16684 81124 16780 81164
rect 16820 81124 16829 81164
rect 17740 81124 19372 81164
rect 19412 81124 19421 81164
rect 19468 81080 19508 81283
rect 19948 81323 20716 81332
rect 19988 81292 20716 81323
rect 20756 81292 20765 81332
rect 19948 81274 19988 81283
rect 21510 81080 21600 81100
rect 0 81040 940 81080
rect 980 81040 989 81080
rect 1459 81040 1468 81080
rect 1508 81040 1996 81080
rect 2036 81040 2045 81080
rect 2921 81040 3052 81080
rect 3092 81040 3101 81080
rect 3475 81040 3484 81080
rect 3524 81040 3533 81080
rect 7555 81040 7564 81080
rect 7604 81040 12500 81080
rect 15139 81040 15148 81080
rect 15188 81040 15319 81080
rect 18163 81040 18172 81080
rect 18212 81040 18604 81080
rect 18644 81040 18653 81080
rect 19372 81040 19508 81080
rect 20995 81040 21004 81080
rect 21044 81040 21600 81080
rect 0 81020 90 81040
rect 3484 80996 3524 81040
rect 3484 80956 17932 80996
rect 17972 80956 18316 80996
rect 18356 80956 18365 80996
rect 3679 80872 3688 80912
rect 3728 80872 3770 80912
rect 3810 80872 3852 80912
rect 3892 80872 3934 80912
rect 3974 80872 4016 80912
rect 4056 80872 4065 80912
rect 7267 80872 7276 80912
rect 7316 80872 8908 80912
rect 8948 80872 8957 80912
rect 18799 80872 18808 80912
rect 18848 80872 18890 80912
rect 18930 80872 18972 80912
rect 19012 80872 19054 80912
rect 19094 80872 19136 80912
rect 19176 80872 19185 80912
rect 19372 80828 19412 81040
rect 21510 81020 21600 81040
rect 1411 80788 1420 80828
rect 1460 80788 2188 80828
rect 2228 80788 2237 80828
rect 14275 80788 14284 80828
rect 14324 80788 14708 80828
rect 0 80744 90 80764
rect 0 80704 1132 80744
rect 1172 80704 1181 80744
rect 2764 80704 3476 80744
rect 5923 80704 5932 80744
rect 5972 80704 6700 80744
rect 6740 80704 6749 80744
rect 11884 80704 13460 80744
rect 0 80684 90 80704
rect 2764 80660 2804 80704
rect 3436 80660 3476 80704
rect 652 80620 2804 80660
rect 2860 80620 3380 80660
rect 3436 80620 4148 80660
rect 4339 80620 4348 80660
rect 4388 80620 6028 80660
rect 6068 80620 6077 80660
rect 652 80492 692 80620
rect 2860 80576 2900 80620
rect 3340 80576 3380 80620
rect 4108 80576 4148 80620
rect 739 80536 748 80576
rect 788 80536 1228 80576
rect 1268 80536 1277 80576
rect 1420 80536 2900 80576
rect 3331 80536 3340 80576
rect 3380 80536 3389 80576
rect 3593 80536 3628 80576
rect 3668 80536 3724 80576
rect 3764 80536 3773 80576
rect 4099 80536 4108 80576
rect 4148 80536 4157 80576
rect 1420 80492 1460 80536
rect 2956 80492 2996 80501
rect 5740 80492 5780 80501
rect 6124 80492 6164 80704
rect 8236 80620 11212 80660
rect 11252 80620 11261 80660
rect 6682 80536 6691 80576
rect 6731 80536 7084 80576
rect 7124 80536 7133 80576
rect 8236 80492 8276 80620
rect 11884 80576 11924 80704
rect 13420 80660 13460 80704
rect 14188 80704 14612 80744
rect 14188 80660 14228 80704
rect 13420 80620 14228 80660
rect 14572 80576 14612 80704
rect 14668 80660 14708 80788
rect 18988 80788 19412 80828
rect 18988 80744 19028 80788
rect 18979 80704 18988 80744
rect 19028 80704 19037 80744
rect 14668 80620 18316 80660
rect 18356 80620 18365 80660
rect 20707 80620 20716 80660
rect 20756 80620 21388 80660
rect 21428 80620 21437 80660
rect 21510 80576 21600 80596
rect 10313 80536 10348 80576
rect 10388 80536 10444 80576
rect 10484 80536 10493 80576
rect 10636 80536 11924 80576
rect 12451 80536 12460 80576
rect 12500 80536 12692 80576
rect 12739 80536 12748 80576
rect 12788 80536 12844 80576
rect 12884 80536 12919 80576
rect 13132 80536 13708 80576
rect 13748 80536 13757 80576
rect 14572 80536 15532 80576
rect 15572 80536 15581 80576
rect 16204 80536 16972 80576
rect 17012 80536 17021 80576
rect 17155 80536 17164 80576
rect 17204 80536 17213 80576
rect 17539 80536 17548 80576
rect 17588 80536 17780 80576
rect 18115 80536 18124 80576
rect 18164 80536 18644 80576
rect 21475 80536 21484 80576
rect 21524 80536 21600 80576
rect 652 80452 788 80492
rect 1123 80452 1132 80492
rect 1172 80452 1460 80492
rect 1699 80452 1708 80492
rect 1748 80452 2476 80492
rect 2516 80452 2525 80492
rect 2851 80452 2860 80492
rect 2900 80452 2956 80492
rect 2996 80452 3148 80492
rect 3188 80452 3197 80492
rect 4291 80452 4300 80492
rect 4340 80452 4492 80492
rect 4532 80452 4541 80492
rect 6106 80452 6115 80492
rect 6155 80452 6164 80492
rect 6220 80452 6412 80492
rect 6452 80452 6461 80492
rect 6508 80452 6551 80492
rect 6591 80452 6600 80492
rect 6700 80452 6796 80492
rect 6836 80452 6845 80492
rect 7075 80452 7084 80492
rect 7124 80452 8276 80492
rect 8332 80492 8372 80501
rect 8908 80492 8948 80501
rect 10636 80492 10676 80536
rect 11980 80492 12020 80501
rect 12652 80492 12692 80536
rect 13132 80492 13172 80536
rect 14476 80492 14516 80501
rect 16204 80492 16244 80536
rect 8372 80452 8908 80492
rect 8948 80452 10100 80492
rect 10147 80452 10156 80492
rect 10196 80452 10676 80492
rect 10723 80452 10732 80492
rect 10772 80452 10903 80492
rect 11849 80452 11980 80492
rect 12020 80452 12500 80492
rect 12652 80452 13172 80492
rect 13219 80452 13228 80492
rect 13268 80452 13324 80492
rect 13364 80452 13399 80492
rect 14516 80452 14764 80492
rect 14804 80452 14813 80492
rect 14947 80452 14956 80492
rect 14996 80452 15860 80492
rect 15907 80452 15916 80492
rect 15956 80452 16204 80492
rect 0 80408 90 80428
rect 0 80368 652 80408
rect 692 80368 701 80408
rect 0 80348 90 80368
rect 748 80240 788 80452
rect 2956 80443 2996 80452
rect 3571 80368 3580 80408
rect 3620 80368 5684 80408
rect 1459 80284 1468 80324
rect 1508 80284 1517 80324
rect 3139 80284 3148 80324
rect 3188 80284 3197 80324
rect 3955 80284 3964 80324
rect 4004 80284 4204 80324
rect 4244 80284 4253 80324
rect 643 80200 652 80240
rect 692 80200 788 80240
rect 1468 80240 1508 80284
rect 3148 80240 3188 80284
rect 5644 80240 5684 80368
rect 5740 80324 5780 80452
rect 6220 80408 6260 80452
rect 6508 80408 6548 80452
rect 6019 80368 6028 80408
rect 6068 80368 6260 80408
rect 6307 80368 6316 80408
rect 6356 80368 6548 80408
rect 6700 80324 6740 80452
rect 8332 80443 8372 80452
rect 8908 80443 8948 80452
rect 10060 80408 10100 80452
rect 11980 80443 12020 80452
rect 12460 80408 12500 80452
rect 14476 80408 14516 80452
rect 6874 80368 6883 80408
rect 6923 80368 7852 80408
rect 7892 80368 7901 80408
rect 10051 80368 10060 80408
rect 10100 80368 10109 80408
rect 10627 80368 10636 80408
rect 10676 80368 11788 80408
rect 11828 80368 11837 80408
rect 12163 80368 12172 80408
rect 12212 80368 12268 80408
rect 12308 80368 12343 80408
rect 12460 80368 14516 80408
rect 14659 80368 14668 80408
rect 14708 80368 15340 80408
rect 15380 80368 15389 80408
rect 15820 80324 15860 80452
rect 16204 80443 16244 80452
rect 16396 80452 16675 80492
rect 16715 80452 16724 80492
rect 16771 80452 16780 80492
rect 16820 80452 16951 80492
rect 16396 80408 16436 80452
rect 16387 80368 16396 80408
rect 16436 80368 16445 80408
rect 5740 80284 6508 80324
rect 6548 80284 6557 80324
rect 6700 80284 7468 80324
rect 7508 80284 7517 80324
rect 8515 80284 8524 80324
rect 8564 80284 8573 80324
rect 8707 80284 8716 80324
rect 8756 80284 8765 80324
rect 10579 80284 10588 80324
rect 10628 80284 12172 80324
rect 12212 80284 12221 80324
rect 12355 80284 12364 80324
rect 12404 80284 12596 80324
rect 12691 80284 12700 80324
rect 12740 80284 12748 80324
rect 12788 80284 12871 80324
rect 13075 80284 13084 80324
rect 13124 80284 14284 80324
rect 14324 80284 14333 80324
rect 15820 80284 16300 80324
rect 16340 80284 16780 80324
rect 16820 80284 16829 80324
rect 1468 80200 1612 80240
rect 1652 80200 1661 80240
rect 3148 80200 4684 80240
rect 4724 80200 4733 80240
rect 5644 80200 7564 80240
rect 7604 80200 7613 80240
rect 4919 80116 4928 80156
rect 4968 80116 5010 80156
rect 5050 80116 5092 80156
rect 5132 80116 5174 80156
rect 5214 80116 5256 80156
rect 5296 80116 5305 80156
rect 0 80072 90 80092
rect 0 80032 460 80072
rect 500 80032 509 80072
rect 0 80012 90 80032
rect 3610 79948 3619 79988
rect 3659 79948 5260 79988
rect 5300 79948 5309 79988
rect 7337 79948 7468 79988
rect 7508 79948 7517 79988
rect 8524 79904 8564 80284
rect 3043 79864 3052 79904
rect 3092 79864 3340 79904
rect 3380 79895 3476 79904
rect 3380 79864 3427 79895
rect 3418 79855 3427 79864
rect 3467 79855 3476 79895
rect 3418 79854 3476 79855
rect 3532 79864 5452 79904
rect 5492 79864 5501 79904
rect 5827 79864 5836 79904
rect 5876 79864 6007 79904
rect 7756 79864 8564 79904
rect 8716 79904 8756 80284
rect 12556 80240 12596 80284
rect 17164 80240 17204 80536
rect 17740 80492 17780 80536
rect 18604 80492 18644 80536
rect 21510 80516 21600 80536
rect 19852 80492 19892 80501
rect 17251 80452 17260 80492
rect 17300 80452 17684 80492
rect 17644 80324 17684 80452
rect 18019 80452 18028 80492
rect 18068 80452 18228 80492
rect 18268 80452 18277 80492
rect 18595 80452 18604 80492
rect 18644 80452 18653 80492
rect 18787 80452 18796 80492
rect 18836 80452 19852 80492
rect 17740 80443 17780 80452
rect 19852 80443 19892 80452
rect 20035 80368 20044 80408
rect 20084 80368 20948 80408
rect 17644 80284 17836 80324
rect 17876 80284 17885 80324
rect 18281 80284 18412 80324
rect 18452 80284 18461 80324
rect 19948 80284 20044 80324
rect 20084 80284 20093 80324
rect 12556 80200 17204 80240
rect 9283 80116 9292 80156
rect 9332 80116 10636 80156
rect 10676 80116 10685 80156
rect 11596 80116 13228 80156
rect 13268 80116 13277 80156
rect 11596 79988 11636 80116
rect 9449 79948 9484 79988
rect 9524 79948 9580 79988
rect 9620 79948 9629 79988
rect 10291 79948 10300 79988
rect 10340 79948 11636 79988
rect 11692 80032 19796 80072
rect 11692 79904 11732 80032
rect 11779 79948 11788 79988
rect 11828 79948 17020 79988
rect 17060 79948 17069 79988
rect 8716 79864 9332 79904
rect 3532 79820 3572 79864
rect 7756 79820 7796 79864
rect 1507 79780 1516 79820
rect 1556 79780 1804 79820
rect 1844 79780 1853 79820
rect 2633 79780 2764 79820
rect 2804 79780 2813 79820
rect 3017 79780 3139 79820
rect 3188 79780 3197 79820
rect 3244 79811 3284 79820
rect 2764 79762 2804 79771
rect 3514 79780 3523 79820
rect 3563 79780 3572 79820
rect 3628 79780 3657 79820
rect 3697 79780 3706 79820
rect 4387 79780 4396 79820
rect 4436 79780 4445 79820
rect 5644 79811 5684 79820
rect 0 79736 90 79756
rect 3244 79736 3284 79771
rect 3628 79736 3668 79780
rect 0 79696 364 79736
rect 404 79696 413 79736
rect 3043 79696 3052 79736
rect 3092 79696 3284 79736
rect 3523 79696 3532 79736
rect 3572 79696 3668 79736
rect 3907 79696 3916 79736
rect 3956 79696 3965 79736
rect 0 79676 90 79696
rect 3916 79652 3956 79696
rect 1228 79612 3956 79652
rect 4396 79652 4436 79780
rect 5897 79780 6028 79820
rect 6068 79780 6077 79820
rect 7241 79811 7372 79820
rect 7241 79780 7276 79811
rect 5644 79736 5684 79771
rect 7316 79780 7372 79811
rect 7412 79780 7421 79820
rect 7738 79780 7747 79820
rect 7787 79780 7796 79820
rect 7843 79780 7852 79820
rect 7892 79780 8023 79820
rect 8105 79780 8236 79820
rect 8276 79780 8285 79820
rect 8681 79780 8812 79820
rect 8852 79780 8861 79820
rect 9292 79811 9332 79864
rect 7276 79736 7316 79771
rect 8812 79762 8852 79771
rect 9292 79762 9332 79771
rect 9388 79864 9676 79904
rect 9716 79864 9725 79904
rect 9907 79864 9916 79904
rect 9956 79864 11732 79904
rect 12499 79864 12508 79904
rect 12548 79864 12844 79904
rect 12884 79864 12893 79904
rect 14179 79864 14188 79904
rect 14228 79864 14804 79904
rect 5644 79696 7316 79736
rect 7459 79696 7468 79736
rect 7508 79696 8332 79736
rect 8372 79696 8381 79736
rect 9388 79652 9428 79864
rect 14764 79820 14804 79864
rect 15436 79864 19412 79904
rect 9868 79780 10732 79820
rect 10772 79780 10781 79820
rect 11683 79780 11692 79820
rect 11732 79780 11924 79820
rect 11971 79780 11980 79820
rect 12020 79780 12172 79820
rect 12212 79780 12221 79820
rect 9868 79736 9908 79780
rect 11884 79736 11924 79780
rect 12268 79756 12300 79796
rect 12340 79756 12349 79796
rect 12460 79780 12638 79820
rect 12678 79780 12687 79820
rect 12739 79780 12748 79820
rect 12788 79780 12797 79820
rect 12931 79780 12940 79820
rect 12980 79780 12989 79820
rect 13123 79780 13132 79820
rect 13172 79780 13324 79820
rect 13364 79780 14092 79820
rect 14132 79780 14141 79820
rect 14249 79780 14380 79820
rect 14420 79780 14429 79820
rect 14755 79780 14764 79820
rect 14804 79780 15340 79820
rect 15380 79780 15389 79820
rect 12268 79736 12308 79756
rect 9545 79696 9676 79736
rect 9716 79696 9908 79736
rect 10051 79696 10060 79736
rect 10100 79696 10109 79736
rect 10627 79696 10636 79736
rect 10676 79696 10685 79736
rect 11081 79696 11116 79736
rect 11156 79696 11212 79736
rect 11252 79696 11261 79736
rect 11657 79696 11788 79736
rect 11828 79696 11837 79736
rect 11884 79696 12308 79736
rect 10060 79652 10100 79696
rect 4396 79612 9292 79652
rect 9332 79612 9341 79652
rect 9388 79612 10100 79652
rect 0 79400 90 79420
rect 0 79360 556 79400
rect 596 79360 605 79400
rect 0 79340 90 79360
rect 1228 79232 1268 79612
rect 2947 79528 2956 79568
rect 2996 79528 3127 79568
rect 4147 79528 4156 79568
rect 4196 79528 6356 79568
rect 7267 79528 7276 79568
rect 7316 79528 10396 79568
rect 10436 79528 10445 79568
rect 6316 79484 6356 79528
rect 10636 79484 10676 79696
rect 12460 79652 12500 79780
rect 12748 79736 12788 79780
rect 12940 79736 12980 79780
rect 14380 79762 14420 79771
rect 12547 79696 12556 79736
rect 12596 79696 12788 79736
rect 12931 79696 12940 79736
rect 12980 79696 13228 79736
rect 13268 79696 13277 79736
rect 15436 79652 15476 79864
rect 15811 79780 15820 79820
rect 15860 79811 16052 79820
rect 15860 79780 16012 79811
rect 16483 79780 16492 79820
rect 16532 79780 17452 79820
rect 17492 79780 17501 79820
rect 18665 79811 18796 79820
rect 18665 79780 18700 79811
rect 16012 79762 16052 79771
rect 18740 79780 18796 79811
rect 18836 79780 18845 79820
rect 18700 79762 18740 79771
rect 19372 79736 19412 79864
rect 19756 79736 19796 80032
rect 19948 79820 19988 80284
rect 20039 80116 20048 80156
rect 20088 80116 20130 80156
rect 20170 80116 20212 80156
rect 20252 80116 20294 80156
rect 20334 80116 20376 80156
rect 20416 80116 20425 80156
rect 20908 80072 20948 80368
rect 21510 80072 21600 80092
rect 20908 80032 21600 80072
rect 21510 80012 21600 80032
rect 19939 79780 19948 79820
rect 19988 79780 19997 79820
rect 16291 79696 16300 79736
rect 16340 79696 16684 79736
rect 16724 79696 16733 79736
rect 17129 79696 17260 79736
rect 17300 79696 17309 79736
rect 19363 79696 19372 79736
rect 19412 79696 19421 79736
rect 19747 79696 19756 79736
rect 19796 79696 19805 79736
rect 20009 79696 20140 79736
rect 20180 79696 20189 79736
rect 20236 79696 21388 79736
rect 21428 79696 21437 79736
rect 20236 79652 20276 79696
rect 11395 79612 11404 79652
rect 11444 79612 12500 79652
rect 12617 79612 12748 79652
rect 12788 79612 12797 79652
rect 14179 79612 14188 79652
rect 14228 79612 15476 79652
rect 19603 79612 19612 79652
rect 19652 79612 20276 79652
rect 20371 79612 20380 79652
rect 20420 79612 21004 79652
rect 21044 79612 21053 79652
rect 21510 79568 21600 79588
rect 11203 79528 11212 79568
rect 11252 79528 11356 79568
rect 11396 79528 11405 79568
rect 12019 79528 12028 79568
rect 12068 79528 12077 79568
rect 14441 79528 14572 79568
rect 14612 79528 14621 79568
rect 15811 79528 15820 79568
rect 15860 79528 16204 79568
rect 16244 79528 16253 79568
rect 16915 79528 16924 79568
rect 16964 79528 18508 79568
rect 18548 79528 18557 79568
rect 18883 79528 18892 79568
rect 18932 79528 19372 79568
rect 19412 79528 19421 79568
rect 19987 79528 19996 79568
rect 20036 79528 20428 79568
rect 20468 79528 20477 79568
rect 20524 79528 21600 79568
rect 6316 79444 8524 79484
rect 8564 79444 8573 79484
rect 8620 79444 10676 79484
rect 12028 79484 12068 79528
rect 20524 79484 20564 79528
rect 21510 79508 21600 79528
rect 12028 79444 20564 79484
rect 8620 79400 8660 79444
rect 3679 79360 3688 79400
rect 3728 79360 3770 79400
rect 3810 79360 3852 79400
rect 3892 79360 3934 79400
rect 3974 79360 4016 79400
rect 4056 79360 4065 79400
rect 6403 79360 6412 79400
rect 6452 79360 8660 79400
rect 9283 79360 9292 79400
rect 9332 79360 13324 79400
rect 13364 79360 13373 79400
rect 18799 79360 18808 79400
rect 18848 79360 18890 79400
rect 18930 79360 18972 79400
rect 19012 79360 19054 79400
rect 19094 79360 19136 79400
rect 19176 79360 19185 79400
rect 10627 79276 10636 79316
rect 10676 79276 11212 79316
rect 11252 79276 11261 79316
rect 13027 79276 13036 79316
rect 13076 79276 20140 79316
rect 20180 79276 20189 79316
rect 547 79192 556 79232
rect 596 79192 1268 79232
rect 2755 79192 2764 79232
rect 2804 79192 2900 79232
rect 3139 79192 3148 79232
rect 3188 79192 3244 79232
rect 3284 79192 3319 79232
rect 12835 79192 12844 79232
rect 12884 79192 12893 79232
rect 15619 79192 15628 79232
rect 15668 79192 15860 79232
rect 19171 79192 19180 79232
rect 19220 79192 19948 79232
rect 19988 79192 19997 79232
rect 76 79108 1036 79148
rect 1076 79108 1085 79148
rect 76 79084 116 79108
rect 0 79024 116 79084
rect 163 79024 172 79064
rect 212 79024 1228 79064
rect 1268 79024 1277 79064
rect 0 79004 90 79024
rect 2860 78980 2900 79192
rect 4291 79108 4300 79148
rect 4340 79108 5396 79148
rect 5443 79108 5452 79148
rect 5492 79108 5500 79148
rect 5540 79108 5623 79148
rect 8236 79108 8812 79148
rect 8852 79108 8861 79148
rect 9667 79108 9676 79148
rect 9716 79108 11212 79148
rect 11252 79108 11261 79148
rect 4300 79064 4340 79108
rect 3331 79024 3340 79064
rect 3380 79024 3389 79064
rect 3916 79024 4340 79064
rect 5356 79064 5396 79108
rect 5356 79024 7028 79064
rect 3340 78980 3380 79024
rect 3916 78980 3956 79024
rect 5164 78980 5204 78989
rect 1481 78940 1612 78980
rect 1652 78940 2188 78980
rect 2228 78940 2237 78980
rect 3113 78940 3244 78980
rect 3284 78940 3293 78980
rect 3340 78940 3359 78980
rect 3399 78940 3427 78980
rect 3523 78940 3532 78980
rect 3572 78940 3703 78980
rect 3907 78940 3916 78980
rect 3956 78940 3965 78980
rect 4291 78940 4300 78980
rect 4340 78940 5164 78980
rect 2860 78896 2900 78940
rect 4300 78896 4340 78940
rect 5164 78931 5204 78940
rect 5260 78940 5644 78980
rect 5684 78940 5693 78980
rect 5827 78940 5836 78980
rect 5876 78940 6007 78980
rect 2860 78856 4340 78896
rect 1459 78772 1468 78812
rect 1508 78772 2188 78812
rect 2228 78772 2237 78812
rect 3043 78772 3052 78812
rect 3092 78772 3340 78812
rect 3380 78772 3389 78812
rect 0 78728 90 78748
rect 5260 78728 5300 78940
rect 6988 78812 7028 79024
rect 7084 79024 7468 79064
rect 7508 79024 7517 79064
rect 8009 79024 8140 79064
rect 8180 79024 8189 79064
rect 7084 78980 7124 79024
rect 8236 78980 8276 79108
rect 9004 79024 9772 79064
rect 9812 79024 9964 79064
rect 10004 79024 10013 79064
rect 10601 79024 10732 79064
rect 10772 79024 10781 79064
rect 12508 79024 12556 79064
rect 12596 79024 12605 79064
rect 12701 79024 12748 79064
rect 12788 79024 12797 79064
rect 7084 78931 7124 78940
rect 7276 78940 7651 78980
rect 7691 78940 7700 78980
rect 7747 78940 7756 78980
rect 7796 78940 7852 78980
rect 7892 78940 7956 78980
rect 8227 78940 8236 78980
rect 8276 78940 8285 78980
rect 8710 78940 8719 78980
rect 8759 78940 8908 78980
rect 8948 78940 8957 78980
rect 7276 78896 7316 78940
rect 7756 78896 7796 78940
rect 9004 78896 9044 79024
rect 12364 78980 12404 78989
rect 9195 78940 9204 78980
rect 9244 78940 9253 78980
rect 11107 78940 11116 78980
rect 11156 78940 11788 78980
rect 11828 78940 11837 78980
rect 7267 78856 7276 78896
rect 7316 78856 7325 78896
rect 7651 78856 7660 78896
rect 7700 78856 7796 78896
rect 8620 78856 9044 78896
rect 8620 78812 8660 78856
rect 5347 78772 5356 78812
rect 5396 78772 5405 78812
rect 6988 78772 8660 78812
rect 0 78688 1900 78728
rect 1940 78688 1949 78728
rect 3139 78688 3148 78728
rect 3188 78688 4108 78728
rect 4148 78688 5300 78728
rect 0 78668 90 78688
rect 4919 78604 4928 78644
rect 4968 78604 5010 78644
rect 5050 78604 5092 78644
rect 5132 78604 5174 78644
rect 5214 78604 5256 78644
rect 5296 78604 5305 78644
rect 5356 78560 5396 78772
rect 9196 78728 9236 78940
rect 9283 78856 9292 78896
rect 9332 78856 9532 78896
rect 9572 78856 9581 78896
rect 10060 78856 10540 78896
rect 10580 78856 10589 78896
rect 9379 78772 9388 78812
rect 9428 78772 9437 78812
rect 9100 78688 9236 78728
rect 9100 78644 9140 78688
rect 3148 78520 3532 78560
rect 3572 78520 4340 78560
rect 2921 78436 3043 78476
rect 3092 78436 3101 78476
rect 0 78392 90 78412
rect 3148 78392 3188 78520
rect 0 78352 844 78392
rect 884 78352 893 78392
rect 3148 78352 3380 78392
rect 0 78332 90 78352
rect 3340 78308 3380 78352
rect 1219 78268 1228 78308
rect 1268 78268 2092 78308
rect 2132 78268 2141 78308
rect 2345 78268 2380 78308
rect 2420 78299 2516 78308
rect 2420 78268 2476 78299
rect 2476 78250 2516 78259
rect 3195 78254 3204 78294
rect 3244 78254 3253 78294
rect 3331 78268 3340 78308
rect 3380 78268 3389 78308
rect 3580 78284 3598 78308
rect 3532 78268 3598 78284
rect 3638 78268 3647 78308
rect 3715 78268 3724 78308
rect 3764 78268 3773 78308
rect 4003 78268 4012 78308
rect 4052 78268 4108 78308
rect 4148 78268 4183 78308
rect 3213 78140 3253 78254
rect 3532 78244 3620 78268
rect 3532 78224 3572 78244
rect 3724 78224 3764 78268
rect 3427 78184 3436 78224
rect 3476 78184 3572 78224
rect 3677 78184 3724 78224
rect 3764 78184 3773 78224
rect 4073 78184 4108 78224
rect 4148 78184 4204 78224
rect 4244 78184 4253 78224
rect 4108 78140 4148 78184
rect 3213 78100 4148 78140
rect 4300 78140 4340 78520
rect 4876 78520 5396 78560
rect 8716 78604 9140 78644
rect 9388 78644 9428 78772
rect 10060 78728 10100 78856
rect 12364 78812 12404 78940
rect 12508 78896 12548 79024
rect 12748 78980 12788 79024
rect 12844 78991 12884 79192
rect 15820 79148 15860 79192
rect 15820 79108 16532 79148
rect 17155 79108 17164 79148
rect 17204 79108 17876 79148
rect 17923 79108 17932 79148
rect 17972 79108 19660 79148
rect 19700 79108 19709 79148
rect 12931 79024 12940 79064
rect 12980 79024 13172 79064
rect 12730 78940 12739 78980
rect 12779 78940 12788 78980
rect 12835 78951 12844 78991
rect 12884 78951 12893 78991
rect 13132 78980 13172 79024
rect 13516 79024 14036 79064
rect 14275 79024 14284 79064
rect 14324 79024 14476 79064
rect 14516 79024 14525 79064
rect 15562 79024 15571 79064
rect 15611 79024 15916 79064
rect 15956 79024 15965 79064
rect 16099 79024 16108 79064
rect 16148 79024 16157 79064
rect 12940 78940 12989 78980
rect 13029 78940 13038 78980
rect 13114 78940 13123 78980
rect 13163 78940 13172 78980
rect 13219 78940 13228 78980
rect 13297 78940 13399 78980
rect 12940 78896 12980 78940
rect 13516 78896 13556 79024
rect 12508 78856 12556 78896
rect 12596 78856 12980 78896
rect 13228 78856 13556 78896
rect 13708 78940 13795 78980
rect 13835 78940 13844 78980
rect 13891 78940 13900 78980
rect 13940 78940 13949 78980
rect 13228 78812 13268 78856
rect 10195 78772 10204 78812
rect 10244 78772 10388 78812
rect 10483 78772 10492 78812
rect 10532 78772 12172 78812
rect 12212 78772 12221 78812
rect 12364 78772 12748 78812
rect 12788 78772 12797 78812
rect 13097 78772 13219 78812
rect 13268 78772 13277 78812
rect 9475 78688 9484 78728
rect 9524 78688 10100 78728
rect 10348 78728 10388 78772
rect 10348 78688 13036 78728
rect 13076 78688 13085 78728
rect 9388 78604 10636 78644
rect 10676 78604 10685 78644
rect 4876 78308 4916 78520
rect 8716 78476 8756 78604
rect 10060 78520 10540 78560
rect 10580 78520 10589 78560
rect 5347 78436 5356 78476
rect 5396 78436 7180 78476
rect 7220 78436 7229 78476
rect 8707 78436 8716 78476
rect 8756 78436 8765 78476
rect 10060 78392 10100 78520
rect 13708 78476 13748 78940
rect 13900 78896 13940 78940
rect 13795 78856 13804 78896
rect 13844 78856 13940 78896
rect 13996 78896 14036 79024
rect 14860 78980 14900 78989
rect 16108 78980 16148 79024
rect 16492 78980 16532 79108
rect 17740 78980 17780 78989
rect 17836 78980 17876 79108
rect 19372 78980 19412 78989
rect 19948 78980 19988 79192
rect 21510 79064 21600 79084
rect 20803 79024 20812 79064
rect 20852 79024 21600 79064
rect 21510 79004 21600 79024
rect 14371 78940 14380 78980
rect 14420 78940 14764 78980
rect 14804 78940 14813 78980
rect 15139 78940 15148 78980
rect 15188 78940 15348 78980
rect 15388 78940 15397 78980
rect 15619 78940 15628 78980
rect 15668 78940 16148 78980
rect 16483 78940 16492 78980
rect 16532 78940 16541 78980
rect 17609 78940 17740 78980
rect 17780 78940 17789 78980
rect 17836 78940 18124 78980
rect 18164 78940 18220 78980
rect 18260 78940 18324 78980
rect 19075 78940 19084 78980
rect 19124 78940 19372 78980
rect 14860 78896 14900 78940
rect 17740 78931 17780 78940
rect 19372 78931 19412 78940
rect 19660 78940 19703 78980
rect 19743 78940 19752 78980
rect 19834 78940 19843 78980
rect 19883 78940 19892 78980
rect 19939 78940 19948 78980
rect 19988 78940 19997 78980
rect 13996 78856 14900 78896
rect 13891 78772 13900 78812
rect 13940 78772 15676 78812
rect 15716 78772 15725 78812
rect 16339 78772 16348 78812
rect 16388 78772 18988 78812
rect 19028 78772 19037 78812
rect 19433 78772 19564 78812
rect 19604 78772 19613 78812
rect 14764 78520 19180 78560
rect 19220 78520 19229 78560
rect 10339 78436 10348 78476
rect 10388 78436 10924 78476
rect 10964 78436 11732 78476
rect 11849 78436 11980 78476
rect 12020 78436 12029 78476
rect 12307 78436 12316 78476
rect 12356 78436 12940 78476
rect 12980 78436 12989 78476
rect 13708 78436 13900 78476
rect 13940 78436 13949 78476
rect 11692 78392 11732 78436
rect 7276 78352 10100 78392
rect 10243 78352 10252 78392
rect 10292 78352 10580 78392
rect 11692 78352 12212 78392
rect 7276 78308 7316 78352
rect 10540 78308 10580 78352
rect 12172 78308 12212 78352
rect 14764 78308 14804 78520
rect 14851 78436 14860 78476
rect 14900 78436 16492 78476
rect 16532 78436 16541 78476
rect 16841 78436 16972 78476
rect 17012 78436 17021 78476
rect 17923 78436 17932 78476
rect 17972 78436 19508 78476
rect 14956 78352 17539 78392
rect 17579 78352 17588 78392
rect 17740 78352 18028 78392
rect 18068 78352 18077 78392
rect 18364 78352 18796 78392
rect 18836 78352 18845 78392
rect 14956 78308 14996 78352
rect 17740 78308 17780 78352
rect 4387 78268 4396 78308
rect 4436 78268 4588 78308
rect 4628 78299 4759 78308
rect 4628 78268 4684 78299
rect 4724 78268 4759 78299
rect 4876 78299 5204 78308
rect 4876 78268 5164 78299
rect 4684 78250 4724 78259
rect 5164 78250 5204 78259
rect 5740 78299 5780 78308
rect 6691 78268 6700 78308
rect 6740 78268 6892 78308
rect 6932 78268 6988 78308
rect 7028 78268 7063 78308
rect 7267 78268 7276 78308
rect 7316 78268 7325 78308
rect 7459 78268 7468 78308
rect 7508 78268 8428 78308
rect 8468 78287 8564 78308
rect 8468 78268 8524 78287
rect 5740 78224 5780 78259
rect 8515 78247 8524 78268
rect 8564 78247 8573 78287
rect 8899 78268 8908 78308
rect 8948 78268 8957 78308
rect 9996 78268 10060 78308
rect 10100 78299 10348 78308
rect 10100 78268 10156 78299
rect 8908 78224 8948 78268
rect 10196 78268 10348 78299
rect 10388 78268 10397 78308
rect 10531 78268 10540 78308
rect 10580 78268 10589 78308
rect 11753 78299 11884 78308
rect 11753 78268 11788 78299
rect 10156 78250 10196 78259
rect 11828 78268 11884 78299
rect 11924 78268 11933 78308
rect 12163 78268 12172 78308
rect 12212 78268 12221 78308
rect 12355 78268 12364 78308
rect 12404 78268 12460 78308
rect 12500 78268 12556 78308
rect 12596 78268 12660 78308
rect 13708 78299 14380 78308
rect 11788 78250 11828 78259
rect 13748 78268 14380 78299
rect 14420 78268 14429 78308
rect 14755 78268 14764 78308
rect 14804 78268 14813 78308
rect 14938 78268 14947 78308
rect 14987 78268 14996 78308
rect 15226 78268 15235 78308
rect 15275 78268 15284 78308
rect 15331 78268 15340 78308
rect 15380 78268 15389 78308
rect 15715 78268 15724 78308
rect 15764 78268 15773 78308
rect 16300 78299 16340 78308
rect 13708 78224 13748 78259
rect 5251 78184 5260 78224
rect 5300 78184 8468 78224
rect 8908 78184 9964 78224
rect 10004 78184 10013 78224
rect 13228 78184 13748 78224
rect 13961 78184 14092 78224
rect 14132 78184 14141 78224
rect 4300 78100 5548 78140
rect 5588 78100 5597 78140
rect 0 78056 90 78076
rect 0 78016 1324 78056
rect 1364 78016 1373 78056
rect 2659 78016 2668 78056
rect 2708 78016 3148 78056
rect 3188 78016 3197 78056
rect 0 77996 90 78016
rect 172 77932 6412 77972
rect 6452 77932 6461 77972
rect 0 77720 90 77740
rect 172 77720 212 77932
rect 8428 77888 8468 78184
rect 9100 78140 9140 78184
rect 9091 78100 9100 78140
rect 9140 78100 9149 78140
rect 10339 78100 10348 78140
rect 10388 78100 12364 78140
rect 12404 78100 12413 78140
rect 13228 78056 13268 78184
rect 15244 78140 15284 78268
rect 15340 78224 15380 78268
rect 15340 78184 15628 78224
rect 15668 78184 15677 78224
rect 13603 78100 13612 78140
rect 13652 78100 15284 78140
rect 9859 78016 9868 78056
rect 9908 78016 13268 78056
rect 13315 78016 13324 78056
rect 13364 78016 13900 78056
rect 13940 78016 14332 78056
rect 14372 78016 14381 78056
rect 15724 77972 15764 78268
rect 16483 78268 16492 78308
rect 16532 78299 16820 78308
rect 16532 78268 16780 78299
rect 15811 78184 15820 78224
rect 15860 78184 16108 78224
rect 16148 78184 16157 78224
rect 16300 78140 16340 78259
rect 17722 78268 17731 78308
rect 17771 78268 17780 78308
rect 18364 78307 18404 78352
rect 19468 78308 19508 78436
rect 18316 78288 18404 78307
rect 16780 78250 16820 78259
rect 18211 78248 18220 78288
rect 18260 78267 18404 78288
rect 18691 78268 18700 78308
rect 18740 78268 18892 78308
rect 18932 78268 18941 78308
rect 19049 78268 19180 78308
rect 19220 78268 19229 78308
rect 19289 78268 19298 78308
rect 19338 78268 19412 78308
rect 19468 78268 19564 78308
rect 19604 78268 19613 78308
rect 18260 78248 18356 78267
rect 17033 78184 17164 78224
rect 17204 78184 17213 78224
rect 18316 78140 18356 78248
rect 19372 78224 19412 78268
rect 18665 78184 18796 78224
rect 18836 78184 18845 78224
rect 19372 78184 19564 78224
rect 19604 78184 19613 78224
rect 16300 78100 17932 78140
rect 17972 78100 17981 78140
rect 18316 78100 19412 78140
rect 17155 78016 17164 78056
rect 17204 78016 17404 78056
rect 17444 78016 17453 78056
rect 18979 78016 18988 78056
rect 19028 78016 19037 78056
rect 18988 77972 19028 78016
rect 8515 77932 8524 77972
rect 8564 77932 15724 77972
rect 15764 77932 15773 77972
rect 18988 77932 19316 77972
rect 19276 77888 19316 77932
rect 19372 77888 19412 78100
rect 19468 78056 19508 78184
rect 19660 78140 19700 78940
rect 19852 78896 19892 78940
rect 19756 78856 19892 78896
rect 20035 78856 20044 78896
rect 20084 78856 20948 78896
rect 19756 78476 19796 78856
rect 19913 78772 19948 78812
rect 19988 78772 20035 78812
rect 20075 78772 20093 78812
rect 20039 78604 20048 78644
rect 20088 78604 20130 78644
rect 20170 78604 20212 78644
rect 20252 78604 20294 78644
rect 20334 78604 20376 78644
rect 20416 78604 20425 78644
rect 20908 78560 20948 78856
rect 21510 78560 21600 78580
rect 20908 78520 21600 78560
rect 21510 78500 21600 78520
rect 19756 78436 20323 78476
rect 20363 78436 20372 78476
rect 19852 78352 20044 78392
rect 20084 78352 20093 78392
rect 19852 78308 19892 78352
rect 19843 78268 19852 78308
rect 19892 78268 19991 78308
rect 20031 78268 20052 78308
rect 20131 78268 20140 78308
rect 20180 78268 20236 78308
rect 20276 78268 20311 78308
rect 20122 78184 20131 78224
rect 20171 78184 20180 78224
rect 20140 78140 20180 78184
rect 19555 78100 19564 78140
rect 19604 78100 19700 78140
rect 20035 78100 20044 78140
rect 20084 78100 20180 78140
rect 21510 78056 21600 78076
rect 19468 78016 20140 78056
rect 20180 78016 20189 78056
rect 20899 78016 20908 78056
rect 20948 78016 21600 78056
rect 21510 77996 21600 78016
rect 3679 77848 3688 77888
rect 3728 77848 3770 77888
rect 3810 77848 3852 77888
rect 3892 77848 3934 77888
rect 3974 77848 4016 77888
rect 4056 77848 4065 77888
rect 8428 77848 12844 77888
rect 12884 77848 12893 77888
rect 13612 77848 16492 77888
rect 16532 77848 16541 77888
rect 18799 77848 18808 77888
rect 18848 77848 18890 77888
rect 18930 77848 18972 77888
rect 19012 77848 19054 77888
rect 19094 77848 19136 77888
rect 19176 77848 19185 77888
rect 19267 77848 19276 77888
rect 19316 77848 19325 77888
rect 19372 77848 20908 77888
rect 20948 77848 20957 77888
rect 3148 77764 6548 77804
rect 3148 77720 3188 77764
rect 0 77680 212 77720
rect 2275 77680 2284 77720
rect 2324 77680 3188 77720
rect 6508 77720 6548 77764
rect 13612 77720 13652 77848
rect 14467 77764 14476 77804
rect 14516 77764 16108 77804
rect 16148 77764 16157 77804
rect 16675 77764 16684 77804
rect 16724 77764 17164 77804
rect 17204 77764 17213 77804
rect 17692 77764 20180 77804
rect 17692 77720 17732 77764
rect 20140 77720 20180 77764
rect 6508 77680 9100 77720
rect 9140 77680 9149 77720
rect 10531 77680 10540 77720
rect 10580 77680 13652 77720
rect 15283 77680 15292 77720
rect 15332 77680 17732 77720
rect 19843 77680 19852 77720
rect 19892 77680 20035 77720
rect 20075 77680 20084 77720
rect 20140 77680 21292 77720
rect 21332 77680 21341 77720
rect 0 77660 90 77680
rect 1459 77596 1468 77636
rect 1508 77596 13516 77636
rect 13556 77596 13565 77636
rect 14441 77596 14476 77636
rect 14516 77596 14572 77636
rect 14612 77596 14621 77636
rect 15715 77596 15724 77636
rect 15764 77596 16052 77636
rect 19363 77596 19372 77636
rect 19412 77596 19421 77636
rect 19843 77596 19852 77636
rect 19892 77596 19901 77636
rect 16012 77552 16052 77596
rect 19372 77552 19412 77596
rect 451 77512 460 77552
rect 500 77512 1228 77552
rect 1268 77512 1277 77552
rect 1324 77512 1612 77552
rect 1652 77512 1661 77552
rect 6988 77512 7852 77552
rect 7892 77512 9868 77552
rect 9908 77512 9917 77552
rect 12547 77512 12556 77552
rect 12596 77512 12748 77552
rect 12788 77512 12797 77552
rect 14921 77512 15052 77552
rect 15092 77512 15101 77552
rect 15532 77512 15820 77552
rect 15860 77512 15869 77552
rect 16003 77512 16012 77552
rect 16052 77512 16061 77552
rect 17827 77512 17836 77552
rect 17876 77512 19028 77552
rect 1324 77468 1364 77512
rect 3436 77468 3476 77477
rect 5068 77468 5108 77477
rect 6988 77468 7028 77512
rect 10348 77468 10388 77477
rect 11980 77468 12020 77477
rect 14380 77468 14420 77477
rect 15532 77468 15572 77512
rect 16588 77468 16628 77477
rect 17644 77468 17684 77477
rect 1315 77428 1324 77468
rect 1364 77428 1373 77468
rect 2153 77428 2188 77468
rect 2228 77428 2284 77468
rect 2324 77428 2333 77468
rect 3305 77428 3436 77468
rect 3476 77428 3485 77468
rect 3689 77428 3820 77468
rect 3860 77428 3869 77468
rect 4291 77428 4300 77468
rect 4340 77428 5068 77468
rect 5731 77428 5740 77468
rect 5780 77428 5789 77468
rect 7555 77428 7564 77468
rect 7604 77428 7756 77468
rect 7796 77428 7805 77468
rect 8515 77428 8524 77468
rect 8564 77428 8812 77468
rect 8852 77428 8861 77468
rect 9091 77428 9100 77468
rect 9140 77428 9908 77468
rect 10217 77428 10348 77468
rect 10388 77428 10397 77468
rect 10531 77428 10540 77468
rect 10580 77428 10732 77468
rect 10772 77428 10781 77468
rect 12163 77428 12172 77468
rect 12212 77428 13132 77468
rect 13172 77428 13181 77468
rect 15514 77428 15523 77468
rect 15563 77428 15572 77468
rect 15619 77428 15628 77468
rect 15668 77428 15799 77468
rect 15977 77428 16108 77468
rect 16148 77428 16157 77468
rect 16628 77428 16684 77468
rect 16724 77428 16759 77468
rect 17098 77428 17107 77468
rect 17147 77428 17156 77468
rect 17513 77428 17644 77468
rect 17684 77428 17693 77468
rect 18761 77428 18892 77468
rect 18932 77428 18941 77468
rect 3436 77419 3476 77428
rect 5068 77419 5108 77428
rect 0 77384 90 77404
rect 0 77344 3148 77384
rect 3188 77344 3197 77384
rect 0 77324 90 77344
rect 1843 77260 1852 77300
rect 1892 77260 1900 77300
rect 1940 77260 2023 77300
rect 3619 77260 3628 77300
rect 3668 77260 4588 77300
rect 4628 77260 4637 77300
rect 5251 77260 5260 77300
rect 5300 77260 5356 77300
rect 5396 77260 5431 77300
rect 5740 77216 5780 77428
rect 6988 77419 7028 77428
rect 8812 77300 8852 77428
rect 9868 77384 9908 77428
rect 10348 77419 10388 77428
rect 11980 77384 12020 77428
rect 14380 77384 14420 77428
rect 16588 77419 16628 77428
rect 17116 77384 17156 77428
rect 17644 77419 17684 77428
rect 18988 77384 19028 77512
rect 19180 77512 19412 77552
rect 19852 77552 19892 77596
rect 21510 77552 21600 77572
rect 19852 77512 20372 77552
rect 21187 77512 21196 77552
rect 21236 77512 21600 77552
rect 19180 77468 19220 77512
rect 20332 77468 20372 77512
rect 21510 77492 21600 77512
rect 19171 77428 19180 77468
rect 19220 77428 19229 77468
rect 19337 77428 19372 77468
rect 19412 77428 19459 77468
rect 19499 77428 19517 77468
rect 19939 77428 19948 77468
rect 19988 77428 20030 77468
rect 20070 77428 20119 77468
rect 20332 77419 20372 77428
rect 9859 77344 9868 77384
rect 9908 77344 9917 77384
rect 11491 77344 11500 77384
rect 11540 77344 12316 77384
rect 12356 77344 12365 77384
rect 12828 77344 12940 77384
rect 12980 77344 12988 77384
rect 13028 77344 16300 77384
rect 16340 77344 16349 77384
rect 17116 77344 17452 77384
rect 17492 77344 17501 77384
rect 18988 77344 19564 77384
rect 19604 77344 19852 77384
rect 19892 77344 19901 77384
rect 7049 77260 7180 77300
rect 7220 77260 7229 77300
rect 7363 77260 7372 77300
rect 7412 77260 8044 77300
rect 8084 77260 8093 77300
rect 8812 77260 10444 77300
rect 10484 77260 10493 77300
rect 12041 77260 12172 77300
rect 12212 77260 12221 77300
rect 17129 77260 17260 77300
rect 17300 77260 17309 77300
rect 20227 77260 20236 77300
rect 20276 77260 20285 77300
rect 20236 77216 20276 77260
rect 2467 77176 2476 77216
rect 2516 77176 5780 77216
rect 6307 77176 6316 77216
rect 6356 77176 12364 77216
rect 12404 77176 12413 77216
rect 15523 77176 15532 77216
rect 15572 77176 15668 77216
rect 2659 77092 2668 77132
rect 2708 77092 4868 77132
rect 4919 77092 4928 77132
rect 4968 77092 5010 77132
rect 5050 77092 5092 77132
rect 5132 77092 5174 77132
rect 5214 77092 5256 77132
rect 5296 77092 5305 77132
rect 10243 77092 10252 77132
rect 10292 77092 10732 77132
rect 10772 77092 11444 77132
rect 14851 77092 14860 77132
rect 14900 77092 15572 77132
rect 0 77048 90 77068
rect 4828 77048 4868 77092
rect 0 77008 4492 77048
rect 4532 77008 4541 77048
rect 4828 77008 11348 77048
rect 0 76988 90 77008
rect 4716 76924 4780 76964
rect 4820 76924 4876 76964
rect 4916 76924 5836 76964
rect 5876 76924 5885 76964
rect 6307 76924 6316 76964
rect 6356 76924 8140 76964
rect 8180 76924 8468 76964
rect 10121 76924 10204 76964
rect 10244 76924 10252 76964
rect 10292 76924 10301 76964
rect 1027 76840 1036 76880
rect 1076 76840 5684 76880
rect 1411 76756 1420 76796
rect 1460 76756 1612 76796
rect 1652 76756 1661 76796
rect 2668 76787 2860 76796
rect 2708 76756 2860 76787
rect 2900 76756 2909 76796
rect 3130 76756 3139 76796
rect 3179 76756 3188 76796
rect 3235 76756 3244 76796
rect 3284 76756 3293 76796
rect 3523 76756 3532 76796
rect 3572 76756 3628 76796
rect 3668 76756 3703 76796
rect 4204 76787 4396 76796
rect 2668 76738 2708 76747
rect 0 76712 90 76732
rect 3148 76712 3188 76756
rect 0 76672 1228 76712
rect 1268 76672 1277 76712
rect 2947 76672 2956 76712
rect 2996 76672 3188 76712
rect 3244 76712 3284 76756
rect 4244 76756 4396 76787
rect 4436 76756 4445 76796
rect 4553 76756 4684 76796
rect 4724 76756 4733 76796
rect 5059 76756 5068 76796
rect 5108 76756 5356 76796
rect 5396 76756 5405 76796
rect 4204 76738 4244 76747
rect 4684 76738 4724 76747
rect 5644 76712 5684 76840
rect 6316 76840 8044 76880
rect 8084 76840 8093 76880
rect 6316 76796 6356 76840
rect 8428 76796 8468 76924
rect 8899 76840 8908 76880
rect 8948 76840 8957 76880
rect 9379 76840 9388 76880
rect 9428 76840 10972 76880
rect 11012 76840 11021 76880
rect 8908 76796 8948 76840
rect 6115 76756 6124 76796
rect 6164 76756 6173 76796
rect 6298 76756 6307 76796
rect 6347 76756 6356 76796
rect 6403 76756 6412 76796
rect 6452 76756 6461 76796
rect 6595 76756 6604 76796
rect 6644 76756 6775 76796
rect 7747 76756 7756 76796
rect 7796 76787 7927 76796
rect 7796 76756 7852 76787
rect 6124 76712 6164 76756
rect 3244 76672 3668 76712
rect 3715 76672 3724 76712
rect 3764 76672 4012 76712
rect 4052 76672 4061 76712
rect 5059 76672 5068 76712
rect 5108 76672 5117 76712
rect 5635 76672 5644 76712
rect 5684 76672 5693 76712
rect 6124 76672 6316 76712
rect 6356 76672 6365 76712
rect 0 76652 90 76672
rect 3628 76628 3668 76672
rect 4012 76628 4052 76672
rect 5068 76628 5108 76672
rect 6412 76628 6452 76756
rect 7892 76756 7927 76787
rect 8314 76756 8323 76796
rect 8363 76756 8372 76796
rect 8419 76756 8428 76796
rect 8468 76756 8477 76796
rect 8681 76756 8812 76796
rect 8852 76756 8861 76796
rect 8908 76787 9428 76796
rect 8908 76756 9388 76787
rect 7852 76738 7892 76747
rect 8332 76712 8372 76756
rect 9737 76756 9868 76796
rect 9908 76756 9917 76796
rect 10588 76756 10636 76796
rect 10676 76756 10704 76796
rect 9388 76712 9428 76747
rect 9868 76738 9908 76747
rect 10588 76712 10628 76756
rect 8323 76672 8332 76712
rect 8372 76672 8419 76712
rect 8899 76672 8908 76712
rect 8948 76672 9100 76712
rect 9140 76672 9149 76712
rect 9379 76672 9388 76712
rect 9428 76672 9504 76712
rect 10090 76672 10099 76712
rect 10139 76672 10444 76712
rect 10484 76672 10493 76712
rect 10540 76672 10588 76712
rect 10628 76672 10637 76712
rect 11203 76672 11212 76712
rect 11252 76672 11261 76712
rect 9100 76628 9140 76672
rect 3619 76588 3628 76628
rect 3668 76588 3677 76628
rect 4012 76588 4300 76628
rect 4340 76588 4349 76628
rect 4675 76588 4684 76628
rect 4724 76588 5108 76628
rect 5164 76588 5404 76628
rect 5444 76588 5453 76628
rect 6412 76588 8044 76628
rect 8084 76588 8236 76628
rect 8276 76588 8285 76628
rect 9100 76588 9964 76628
rect 10004 76588 10013 76628
rect 10060 76588 10444 76628
rect 10484 76588 10493 76628
rect 5164 76544 5204 76588
rect 10060 76544 10100 76588
rect 10540 76544 10580 76672
rect 10867 76588 10876 76628
rect 10916 76588 10924 76628
rect 10964 76588 11047 76628
rect 11212 76544 11252 76672
rect 11308 76628 11348 77008
rect 11404 76796 11444 77092
rect 14467 77008 14476 77048
rect 14516 77008 14525 77048
rect 14476 76964 14516 77008
rect 13996 76924 14092 76964
rect 14132 76924 14141 76964
rect 14476 76924 14852 76964
rect 15113 76924 15148 76964
rect 15188 76924 15244 76964
rect 15284 76924 15293 76964
rect 13027 76840 13036 76880
rect 13076 76840 13085 76880
rect 13036 76796 13076 76840
rect 13996 76796 14036 76924
rect 14812 76796 14852 76924
rect 15532 76880 15572 77092
rect 15628 76964 15668 77176
rect 19948 77176 20276 77216
rect 19948 76964 19988 77176
rect 20039 77092 20048 77132
rect 20088 77092 20130 77132
rect 20170 77092 20212 77132
rect 20252 77092 20294 77132
rect 20334 77092 20376 77132
rect 20416 77092 20425 77132
rect 21510 77048 21600 77068
rect 20140 77008 21600 77048
rect 15628 76924 15772 76964
rect 15812 76924 15820 76964
rect 15860 76924 15972 76964
rect 16204 76924 18892 76964
rect 18932 76924 18941 76964
rect 19948 76924 19996 76964
rect 20036 76924 20045 76964
rect 15532 76840 15676 76880
rect 15716 76840 15725 76880
rect 16204 76796 16244 76924
rect 20140 76880 20180 77008
rect 21510 76988 21600 77008
rect 17452 76840 18356 76880
rect 18595 76840 18604 76880
rect 18644 76840 20180 76880
rect 17452 76796 17492 76840
rect 18316 76796 18356 76840
rect 11404 76756 11596 76796
rect 11636 76756 11645 76796
rect 12809 76787 12940 76796
rect 12809 76756 12844 76787
rect 12884 76756 12940 76787
rect 12980 76756 12989 76796
rect 13036 76756 13507 76796
rect 13547 76756 13556 76796
rect 13603 76756 13612 76796
rect 13652 76756 13804 76796
rect 13844 76756 13853 76796
rect 13987 76756 13996 76796
rect 14036 76756 14045 76796
rect 14537 76787 14668 76796
rect 14537 76756 14572 76787
rect 12844 76738 12884 76747
rect 14612 76756 14668 76787
rect 14708 76756 14717 76796
rect 14812 76787 15092 76796
rect 14812 76756 15052 76787
rect 14572 76738 14612 76747
rect 15052 76738 15092 76747
rect 16012 76756 16204 76796
rect 16244 76756 16253 76796
rect 16963 76756 16972 76796
rect 17012 76787 17492 76796
rect 17012 76756 17452 76787
rect 16012 76712 16052 76756
rect 18089 76756 18220 76796
rect 18260 76756 18269 76796
rect 18316 76787 19508 76796
rect 18316 76756 19468 76787
rect 17452 76738 17492 76747
rect 19843 76756 19852 76796
rect 19892 76756 19948 76796
rect 19988 76756 20023 76796
rect 20093 76756 20140 76796
rect 20180 76756 20189 76796
rect 19468 76738 19508 76747
rect 20140 76712 20180 76756
rect 13961 76672 14092 76712
rect 14132 76672 14141 76712
rect 15305 76672 15340 76712
rect 15380 76672 15436 76712
rect 15476 76672 15485 76712
rect 16003 76672 16012 76712
rect 16052 76672 16061 76712
rect 17827 76672 17836 76712
rect 17876 76672 17885 76712
rect 20131 76672 20140 76712
rect 20180 76672 20189 76712
rect 20371 76672 20380 76712
rect 20420 76672 21428 76712
rect 16012 76628 16052 76672
rect 11308 76588 16052 76628
rect 2659 76504 2668 76544
rect 2708 76504 2860 76544
rect 2900 76504 2909 76544
rect 4483 76504 4492 76544
rect 4532 76504 5204 76544
rect 5299 76504 5308 76544
rect 5348 76504 5357 76544
rect 6281 76504 6412 76544
rect 6452 76504 6461 76544
rect 6595 76504 6604 76544
rect 6644 76504 10100 76544
rect 10444 76504 10580 76544
rect 10828 76504 11252 76544
rect 17513 76504 17644 76544
rect 17684 76504 17693 76544
rect 5308 76460 5348 76504
rect 10444 76460 10484 76504
rect 10828 76460 10868 76504
rect 2860 76420 4148 76460
rect 5308 76420 10060 76460
rect 10100 76420 10109 76460
rect 10435 76420 10444 76460
rect 10484 76420 10493 76460
rect 10732 76420 10868 76460
rect 11212 76420 15628 76460
rect 15668 76420 15677 76460
rect 0 76376 90 76396
rect 2860 76376 2900 76420
rect 4108 76376 4148 76420
rect 10732 76376 10772 76420
rect 11212 76376 11252 76420
rect 17836 76376 17876 76672
rect 21388 76628 21428 76672
rect 18067 76588 18076 76628
rect 18116 76588 20428 76628
rect 20468 76588 20477 76628
rect 21379 76588 21388 76628
rect 21428 76588 21437 76628
rect 21510 76544 21600 76564
rect 19651 76504 19660 76544
rect 19700 76504 19892 76544
rect 19852 76460 19892 76504
rect 21388 76504 21600 76544
rect 18499 76420 18508 76460
rect 18548 76420 19796 76460
rect 19843 76420 19852 76460
rect 19892 76420 19901 76460
rect 0 76336 2900 76376
rect 3679 76336 3688 76376
rect 3728 76336 3770 76376
rect 3810 76336 3852 76376
rect 3892 76336 3934 76376
rect 3974 76336 4016 76376
rect 4056 76336 4065 76376
rect 4108 76336 10772 76376
rect 10828 76336 11252 76376
rect 12355 76336 12364 76376
rect 12404 76336 17876 76376
rect 18799 76336 18808 76376
rect 18848 76336 18890 76376
rect 18930 76336 18972 76376
rect 19012 76336 19054 76376
rect 19094 76336 19136 76376
rect 19176 76336 19185 76376
rect 0 76316 90 76336
rect 10828 76292 10868 76336
rect 19756 76292 19796 76420
rect 21388 76376 21428 76504
rect 21510 76484 21600 76504
rect 19948 76336 21428 76376
rect 19948 76292 19988 76336
rect 8044 76252 10868 76292
rect 13324 76252 14092 76292
rect 14132 76252 14764 76292
rect 14804 76252 14813 76292
rect 17059 76252 17068 76292
rect 17108 76252 18220 76292
rect 18260 76252 18269 76292
rect 19756 76252 19988 76292
rect 8044 76208 8084 76252
rect 5971 76168 5980 76208
rect 6020 76168 8084 76208
rect 8201 76168 8332 76208
rect 8372 76168 8381 76208
rect 9833 76168 9868 76208
rect 9908 76168 9964 76208
rect 10004 76168 10013 76208
rect 11923 76168 11932 76208
rect 11972 76168 12364 76208
rect 12404 76168 12413 76208
rect 7939 76084 7948 76124
rect 7988 76084 8549 76124
rect 8899 76084 8908 76124
rect 8948 76084 10732 76124
rect 10772 76084 10781 76124
rect 11683 76084 11692 76124
rect 11732 76084 12844 76124
rect 12884 76084 12893 76124
rect 0 76040 90 76060
rect 0 76000 1420 76040
rect 1460 76000 1469 76040
rect 2851 76000 2860 76040
rect 2900 76000 3031 76040
rect 3523 76000 3532 76040
rect 3572 76000 3916 76040
rect 3956 76000 3965 76040
rect 4291 76000 4300 76040
rect 4340 76000 4349 76040
rect 5417 76000 5548 76040
rect 5588 76000 5597 76040
rect 5731 76000 5740 76040
rect 5780 76000 5789 76040
rect 5923 76000 5932 76040
rect 5972 76000 6124 76040
rect 6164 76000 6173 76040
rect 6499 76000 6508 76040
rect 6548 76000 7468 76040
rect 7508 76000 7517 76040
rect 0 75980 90 76000
rect 2476 75956 2516 75965
rect 4300 75956 4340 76000
rect 4492 75956 4532 75965
rect 5740 75956 5780 76000
rect 8140 75956 8180 75965
rect 1097 75916 1228 75956
rect 1268 75916 1277 75956
rect 2371 75916 2380 75956
rect 2420 75916 2476 75956
rect 2516 75916 2551 75956
rect 3275 75916 3340 75956
rect 3380 75916 3406 75956
rect 3446 75916 3455 75956
rect 3523 75916 3532 75956
rect 3572 75916 3628 75956
rect 3668 75916 3703 75956
rect 4003 75916 4012 75956
rect 4052 75916 4340 75956
rect 4387 75916 4396 75956
rect 4436 75916 4492 75956
rect 4532 75916 4567 75956
rect 4937 75916 5011 75956
rect 5051 75916 5068 75956
rect 5108 75916 5117 75956
rect 5251 75916 5260 75956
rect 5300 75916 5780 75956
rect 6857 75916 6892 75956
rect 6932 75916 6988 75956
rect 7028 75916 7037 75956
rect 7843 75916 7852 75956
rect 7892 75916 8140 75956
rect 8509 75956 8549 76084
rect 13324 76040 13364 76252
rect 15043 76168 15052 76208
rect 15092 76168 17876 76208
rect 18115 76168 18124 76208
rect 18164 76168 18364 76208
rect 18404 76168 18413 76208
rect 15331 76084 15340 76124
rect 15380 76084 15476 76124
rect 9772 76000 10924 76040
rect 10964 76000 10973 76040
rect 13123 76000 13132 76040
rect 13172 76000 13364 76040
rect 13678 76000 13708 76040
rect 13748 76000 13765 76040
rect 9772 75956 9812 76000
rect 11500 75956 11540 75965
rect 13725 75956 13765 76000
rect 15340 75956 15380 75965
rect 8509 75916 8524 75956
rect 8564 75916 9484 75956
rect 9524 75916 9533 75956
rect 2476 75907 2516 75916
rect 4492 75907 4532 75916
rect 8140 75872 8180 75916
rect 9772 75872 9812 75916
rect 5164 75832 6124 75872
rect 6164 75832 6892 75872
rect 6932 75832 6941 75872
rect 8140 75832 9812 75872
rect 9868 75916 10252 75956
rect 10292 75916 10301 75956
rect 11369 75916 11500 75956
rect 11540 75916 11549 75956
rect 12041 75916 12163 75956
rect 12212 75916 12221 75956
rect 12648 75916 12657 75956
rect 12697 75916 13036 75956
rect 13076 75916 13085 75956
rect 13193 75916 13228 75956
rect 13268 75916 13324 75956
rect 13364 75916 13373 75956
rect 13481 75916 13612 75956
rect 13652 75916 13661 75956
rect 13716 75916 13725 75956
rect 13765 75916 13774 75956
rect 14083 75916 14092 75956
rect 14132 75916 14141 75956
rect 14371 75916 14380 75956
rect 14420 75916 15340 75956
rect 15436 75956 15476 76084
rect 17836 76040 17876 76168
rect 19267 76084 19276 76124
rect 19316 76084 20276 76124
rect 20236 76040 20276 76084
rect 21510 76040 21600 76060
rect 17635 76000 17644 76040
rect 17684 76000 17780 76040
rect 17836 76000 18124 76040
rect 18164 76000 18892 76040
rect 18932 76000 18941 76040
rect 20009 76000 20140 76040
rect 20180 76000 20189 76040
rect 20236 76000 21600 76040
rect 16972 75956 17012 75965
rect 17740 75956 17780 76000
rect 21510 75980 21600 76000
rect 19756 75956 19796 75965
rect 15436 75916 15724 75956
rect 15764 75916 15773 75956
rect 17059 75916 17068 75956
rect 17108 75916 17347 75956
rect 17387 75916 17396 75956
rect 17482 75916 17491 75956
rect 17531 75916 17540 75956
rect 17622 75916 17631 75956
rect 17671 75916 17680 75956
rect 17722 75916 17731 75956
rect 17771 75916 17780 75956
rect 17827 75916 17836 75956
rect 17905 75916 18007 75956
rect 18211 75916 18220 75956
rect 18260 75916 18508 75956
rect 18548 75916 18557 75956
rect 5164 75788 5204 75832
rect 9868 75788 9908 75916
rect 11500 75907 11540 75916
rect 14092 75872 14132 75916
rect 15340 75907 15380 75916
rect 16972 75872 17012 75916
rect 17500 75872 17540 75916
rect 12451 75832 12460 75872
rect 12500 75832 12844 75872
rect 12884 75832 14132 75872
rect 16841 75832 16972 75872
rect 17012 75832 17060 75872
rect 2659 75748 2668 75788
rect 2708 75748 2764 75788
rect 2804 75748 2839 75788
rect 3091 75748 3100 75788
rect 3140 75748 5108 75788
rect 5155 75748 5164 75788
rect 5204 75748 5213 75788
rect 5299 75748 5308 75788
rect 5348 75748 5452 75788
rect 5492 75748 5501 75788
rect 6355 75748 6364 75788
rect 6404 75748 6452 75788
rect 6499 75748 6508 75788
rect 6548 75748 6748 75788
rect 6788 75748 6797 75788
rect 6979 75748 6988 75788
rect 7028 75748 7372 75788
rect 7412 75748 9908 75788
rect 9964 75748 13708 75788
rect 13748 75748 13996 75788
rect 14036 75748 14045 75788
rect 15401 75748 15532 75788
rect 15572 75748 15581 75788
rect 0 75704 90 75724
rect 5068 75704 5108 75748
rect 6412 75704 6452 75748
rect 9964 75704 10004 75748
rect 17020 75704 17060 75832
rect 17260 75832 17540 75872
rect 17640 75872 17680 75916
rect 19756 75872 19796 75916
rect 17640 75832 17740 75872
rect 17780 75832 17789 75872
rect 18499 75832 18508 75872
rect 18548 75832 19796 75872
rect 17260 75788 17300 75832
rect 17129 75748 17164 75788
rect 17204 75748 17260 75788
rect 17300 75748 17309 75788
rect 17417 75748 17548 75788
rect 17588 75748 17597 75788
rect 19817 75748 19948 75788
rect 19988 75748 19997 75788
rect 20371 75748 20380 75788
rect 20420 75748 20908 75788
rect 20948 75748 20957 75788
rect 0 75664 940 75704
rect 980 75664 989 75704
rect 5068 75664 6356 75704
rect 6412 75664 10004 75704
rect 10060 75664 15340 75704
rect 15380 75664 15389 75704
rect 17020 75664 17588 75704
rect 0 75644 90 75664
rect 6316 75620 6356 75664
rect 10060 75620 10100 75664
rect 1603 75580 1612 75620
rect 1652 75580 4684 75620
rect 4724 75580 4733 75620
rect 4919 75580 4928 75620
rect 4968 75580 5010 75620
rect 5050 75580 5092 75620
rect 5132 75580 5174 75620
rect 5214 75580 5256 75620
rect 5296 75580 5305 75620
rect 6316 75580 10100 75620
rect 12940 75580 15052 75620
rect 15092 75580 15101 75620
rect 12940 75536 12980 75580
rect 17548 75536 17588 75664
rect 20039 75580 20048 75620
rect 20088 75580 20130 75620
rect 20170 75580 20212 75620
rect 20252 75580 20294 75620
rect 20334 75580 20376 75620
rect 20416 75580 20425 75620
rect 21510 75536 21600 75556
rect 2860 75496 8908 75536
rect 8948 75496 8957 75536
rect 10252 75496 12980 75536
rect 13603 75496 13612 75536
rect 13652 75496 15092 75536
rect 17539 75496 17548 75536
rect 17588 75496 17597 75536
rect 21091 75496 21100 75536
rect 21140 75496 21600 75536
rect 2860 75452 2900 75496
rect 10252 75452 10292 75496
rect 2227 75412 2236 75452
rect 2276 75412 2900 75452
rect 7939 75412 7948 75452
rect 7988 75412 8180 75452
rect 8419 75412 8428 75452
rect 8468 75412 9004 75452
rect 9044 75412 9053 75452
rect 10051 75412 10060 75452
rect 10100 75412 10292 75452
rect 11155 75412 11164 75452
rect 11204 75412 13036 75452
rect 13076 75412 13085 75452
rect 13411 75412 13420 75452
rect 13460 75412 14044 75452
rect 14084 75412 14093 75452
rect 0 75368 90 75388
rect 0 75328 268 75368
rect 308 75328 317 75368
rect 556 75328 2476 75368
rect 2516 75328 2525 75368
rect 6403 75328 6412 75368
rect 6452 75328 7988 75368
rect 0 75308 90 75328
rect 0 75032 90 75052
rect 556 75032 596 75328
rect 7948 75284 7988 75328
rect 8140 75284 8180 75412
rect 8340 75328 8660 75368
rect 10723 75328 10732 75368
rect 10772 75328 14996 75368
rect 8340 75284 8380 75328
rect 8620 75284 8660 75328
rect 14956 75284 14996 75328
rect 15052 75284 15092 75496
rect 21510 75476 21600 75496
rect 16553 75412 16588 75452
rect 16628 75412 16684 75452
rect 16724 75412 16733 75452
rect 16195 75328 16204 75368
rect 16244 75328 18796 75368
rect 18836 75328 20180 75368
rect 2275 75244 2284 75284
rect 2324 75244 2668 75284
rect 2708 75244 2717 75284
rect 2860 75275 3956 75284
rect 2860 75244 3916 75275
rect 2860 75200 2900 75244
rect 4675 75244 4684 75284
rect 4724 75244 4876 75284
rect 4916 75244 4925 75284
rect 5932 75275 6124 75284
rect 3916 75226 3956 75235
rect 5972 75244 6124 75275
rect 6164 75244 6173 75284
rect 6307 75244 6316 75284
rect 6356 75244 6988 75284
rect 7028 75244 7037 75284
rect 7564 75275 7756 75284
rect 5932 75226 5972 75235
rect 7604 75244 7756 75275
rect 7796 75244 7805 75284
rect 7930 75244 7939 75284
rect 7979 75244 7988 75284
rect 8044 75275 8084 75284
rect 7564 75226 7604 75235
rect 8140 75275 8228 75284
rect 8140 75244 8188 75275
rect 8044 75200 8084 75235
rect 8340 75244 8362 75284
rect 8402 75244 8411 75284
rect 8491 75244 8500 75284
rect 8540 75281 8549 75284
rect 8540 75244 8569 75281
rect 8611 75244 8620 75284
rect 8660 75244 8716 75284
rect 8756 75244 8791 75284
rect 8849 75244 8858 75284
rect 8898 75244 8908 75284
rect 8948 75244 9236 75284
rect 9283 75244 9292 75284
rect 9332 75244 9341 75284
rect 10243 75244 10252 75284
rect 10292 75275 11500 75284
rect 10292 75244 10540 75275
rect 8509 75241 8569 75244
rect 8188 75226 8228 75235
rect 643 75160 652 75200
rect 692 75160 1228 75200
rect 1268 75160 1277 75200
rect 1411 75160 1420 75200
rect 1460 75160 1612 75200
rect 1652 75160 1661 75200
rect 1987 75160 1996 75200
rect 2036 75160 2045 75200
rect 2371 75160 2380 75200
rect 2420 75160 2900 75200
rect 4483 75160 4492 75200
rect 4532 75160 4684 75200
rect 4724 75160 4733 75200
rect 8035 75160 8044 75200
rect 8084 75160 8131 75200
rect 1996 75116 2036 75160
rect 8529 75116 8569 75241
rect 9196 75200 9236 75244
rect 9187 75160 9196 75200
rect 9236 75160 9245 75200
rect 835 75076 844 75116
rect 884 75076 2036 75116
rect 3331 75076 3340 75116
rect 3380 75076 4252 75116
rect 4292 75076 4301 75116
rect 4867 75076 4876 75116
rect 4916 75076 8276 75116
rect 8419 75076 8428 75116
rect 8468 75076 8569 75116
rect 8236 75032 8276 75076
rect 9292 75032 9332 75244
rect 10580 75244 11500 75275
rect 11540 75244 11549 75284
rect 12748 75244 13364 75284
rect 13411 75244 13420 75284
rect 13460 75244 13708 75284
rect 13748 75244 13757 75284
rect 14275 75244 14284 75284
rect 14324 75244 14516 75284
rect 14938 75244 14947 75284
rect 14987 75244 14996 75284
rect 15043 75244 15052 75284
rect 15092 75244 15101 75284
rect 15331 75244 15340 75284
rect 15380 75244 15436 75284
rect 15476 75244 15511 75284
rect 16003 75244 16012 75284
rect 16052 75244 16396 75284
rect 16436 75244 16445 75284
rect 16492 75275 16532 75284
rect 10540 75226 10580 75235
rect 12748 75200 12788 75244
rect 13324 75200 13364 75244
rect 14476 75200 14516 75244
rect 16012 75226 16052 75235
rect 16716 75244 16780 75284
rect 16820 75244 16876 75284
rect 16916 75244 17012 75284
rect 17059 75244 17068 75284
rect 17108 75275 18508 75284
rect 17108 75244 18124 75275
rect 16492 75200 16532 75235
rect 16972 75200 17012 75244
rect 18164 75244 18508 75275
rect 18548 75244 18557 75284
rect 18761 75244 18892 75284
rect 18932 75244 18941 75284
rect 20140 75275 20180 75328
rect 18124 75226 18164 75235
rect 20140 75226 20180 75235
rect 10636 75160 10924 75200
rect 10964 75160 11884 75200
rect 11924 75160 11933 75200
rect 12617 75160 12748 75200
rect 12788 75160 12797 75200
rect 12931 75160 12940 75200
rect 12980 75160 12989 75200
rect 13164 75160 13180 75200
rect 13220 75160 13324 75200
rect 13364 75160 13373 75200
rect 13699 75160 13708 75200
rect 13748 75160 13996 75200
rect 14036 75160 14045 75200
rect 14153 75160 14188 75200
rect 14228 75160 14284 75200
rect 14324 75160 14333 75200
rect 14467 75160 14476 75200
rect 14516 75160 14525 75200
rect 14851 75160 14860 75200
rect 14900 75160 15532 75200
rect 15572 75160 15628 75200
rect 15668 75160 15732 75200
rect 16099 75160 16108 75200
rect 16148 75160 16532 75200
rect 16963 75160 16972 75200
rect 17012 75160 17021 75200
rect 18307 75160 18316 75200
rect 18356 75160 18508 75200
rect 18548 75160 18557 75200
rect 10636 75116 10676 75160
rect 12940 75116 12980 75160
rect 10243 75076 10252 75116
rect 10292 75076 10676 75116
rect 10915 75076 10924 75116
rect 10964 75076 12980 75116
rect 13315 75076 13324 75116
rect 13364 75076 13564 75116
rect 13604 75076 13613 75116
rect 13939 75076 13948 75116
rect 13988 75076 20332 75116
rect 20372 75076 20381 75116
rect 21510 75032 21600 75052
rect 0 74992 596 75032
rect 1459 74992 1468 75032
rect 1508 74992 1612 75032
rect 1652 74992 1661 75032
rect 1843 74992 1852 75032
rect 1892 74992 2132 75032
rect 3977 74992 4108 75032
rect 4148 74992 4157 75032
rect 5731 74992 5740 75032
rect 5780 74992 6124 75032
rect 6164 74992 6173 75032
rect 7625 74992 7756 75032
rect 7796 74992 7805 75032
rect 7930 74992 7939 75032
rect 7988 74992 8119 75032
rect 8236 74992 9332 75032
rect 12163 74992 12172 75032
rect 12212 74992 12508 75032
rect 12548 74992 14036 75032
rect 14707 74992 14716 75032
rect 14756 74992 17492 75032
rect 18019 74992 18028 75032
rect 18068 74992 18316 75032
rect 18356 74992 18365 75032
rect 18739 74992 18748 75032
rect 18788 74992 19276 75032
rect 19316 74992 19325 75032
rect 20035 74992 20044 75032
rect 20084 74992 20332 75032
rect 20372 74992 20381 75032
rect 21283 74992 21292 75032
rect 21332 74992 21600 75032
rect 0 74972 90 74992
rect 2092 74948 2132 74992
rect 13996 74948 14036 74992
rect 17452 74948 17492 74992
rect 21510 74972 21600 74992
rect 931 74908 940 74948
rect 980 74908 989 74948
rect 2092 74908 13804 74948
rect 13844 74908 13853 74948
rect 13996 74908 17068 74948
rect 17108 74908 17117 74948
rect 17452 74908 21100 74948
rect 21140 74908 21149 74948
rect 940 74864 980 74908
rect 259 74824 268 74864
rect 308 74824 980 74864
rect 3679 74824 3688 74864
rect 3728 74824 3770 74864
rect 3810 74824 3852 74864
rect 3892 74824 3934 74864
rect 3974 74824 4016 74864
rect 4056 74824 4065 74864
rect 12451 74824 12460 74864
rect 12500 74824 18316 74864
rect 18356 74824 18365 74864
rect 18799 74824 18808 74864
rect 18848 74824 18890 74864
rect 18930 74824 18972 74864
rect 19012 74824 19054 74864
rect 19094 74824 19136 74864
rect 19176 74824 19185 74864
rect 4012 74740 4300 74780
rect 4340 74740 4349 74780
rect 8899 74740 8908 74780
rect 8948 74740 20180 74780
rect 0 74696 90 74716
rect 0 74656 556 74696
rect 596 74656 605 74696
rect 0 74636 90 74656
rect 2729 74488 2860 74528
rect 2900 74488 2909 74528
rect 3523 74488 3532 74528
rect 3572 74488 3916 74528
rect 3956 74488 3965 74528
rect 2476 74444 2516 74453
rect 4012 74444 4052 74740
rect 4204 74656 5260 74696
rect 5300 74656 5309 74696
rect 5491 74656 5500 74696
rect 5540 74656 8428 74696
rect 8468 74656 8477 74696
rect 9475 74656 9484 74696
rect 9524 74656 11636 74696
rect 11683 74656 11692 74696
rect 11732 74656 12748 74696
rect 12788 74656 12797 74696
rect 15331 74656 15340 74696
rect 15380 74656 17068 74696
rect 17108 74656 17156 74696
rect 17225 74656 17356 74696
rect 17396 74656 17405 74696
rect 17683 74656 17692 74696
rect 17732 74656 17836 74696
rect 17876 74656 17885 74696
rect 1097 74404 1228 74444
rect 1268 74404 1277 74444
rect 2345 74404 2476 74444
rect 2516 74404 2525 74444
rect 2659 74404 2668 74444
rect 2708 74404 3427 74444
rect 3467 74404 3476 74444
rect 3523 74404 3532 74444
rect 3572 74404 3619 74444
rect 3881 74404 4012 74444
rect 4052 74404 4061 74444
rect 2476 74395 2516 74404
rect 0 74360 90 74380
rect 3532 74360 3572 74404
rect 0 74320 1804 74360
rect 1844 74320 1853 74360
rect 3523 74320 3532 74360
rect 3572 74320 3581 74360
rect 0 74300 90 74320
rect 4204 74276 4244 74656
rect 5059 74572 5068 74612
rect 5108 74572 10060 74612
rect 10100 74572 10109 74612
rect 5693 74488 5740 74528
rect 5780 74488 5789 74528
rect 6089 74488 6220 74528
rect 6260 74488 6269 74528
rect 6316 74488 6700 74528
rect 6740 74488 6749 74528
rect 7817 74488 7852 74528
rect 7892 74488 7948 74528
rect 7988 74488 7997 74528
rect 8419 74488 8428 74528
rect 8468 74488 8477 74528
rect 9868 74488 10252 74528
rect 10292 74488 10301 74528
rect 4492 74444 4532 74453
rect 5740 74444 5780 74488
rect 6316 74444 6356 74488
rect 6796 74444 6836 74453
rect 8428 74444 8468 74488
rect 9868 74444 9908 74488
rect 11500 74444 11540 74453
rect 11596 74444 11636 74656
rect 13315 74488 13324 74528
rect 13364 74488 13612 74528
rect 13652 74488 13661 74528
rect 14380 74488 14572 74528
rect 14612 74488 14621 74528
rect 14851 74488 14860 74528
rect 14900 74488 14909 74528
rect 15619 74488 15628 74528
rect 15668 74488 16100 74528
rect 13228 74444 13268 74453
rect 14380 74444 14420 74488
rect 4387 74404 4396 74444
rect 4436 74404 4492 74444
rect 4532 74404 4780 74444
rect 4820 74404 4829 74444
rect 4937 74404 5011 74444
rect 5051 74404 5068 74444
rect 5108 74404 5117 74444
rect 5347 74404 5356 74444
rect 5396 74404 5405 74444
rect 5722 74404 5731 74444
rect 5771 74404 5780 74444
rect 5827 74404 5836 74444
rect 5876 74404 5885 74444
rect 6307 74404 6316 74444
rect 6356 74404 6365 74444
rect 6700 74404 6796 74444
rect 6836 74404 7084 74444
rect 7124 74404 7133 74444
rect 7180 74404 7284 74444
rect 7324 74404 7333 74444
rect 7852 74404 8468 74444
rect 8585 74404 8620 74444
rect 8660 74404 8716 74444
rect 8756 74404 9100 74444
rect 9140 74404 9149 74444
rect 10243 74404 10252 74444
rect 10292 74404 10301 74444
rect 11369 74404 11500 74444
rect 11540 74404 11549 74444
rect 11596 74404 11980 74444
rect 12020 74404 12029 74444
rect 12739 74404 12748 74444
rect 12788 74404 13228 74444
rect 13795 74404 13804 74444
rect 13844 74404 14228 74444
rect 14362 74404 14371 74444
rect 14411 74404 14420 74444
rect 14467 74404 14476 74444
rect 14516 74404 14647 74444
rect 4492 74395 4532 74404
rect 5356 74360 5396 74404
rect 5836 74360 5876 74404
rect 5356 74320 5444 74360
rect 5827 74320 5836 74360
rect 5876 74320 5923 74360
rect 5404 74276 5444 74320
rect 6700 74276 6740 74404
rect 6796 74395 6836 74404
rect 7180 74276 7220 74404
rect 7852 74360 7892 74404
rect 9868 74395 9908 74404
rect 7363 74320 7372 74360
rect 7412 74320 7892 74360
rect 8035 74320 8044 74360
rect 8084 74320 8092 74360
rect 8132 74320 8215 74360
rect 2537 74236 2668 74276
rect 2708 74236 2717 74276
rect 3091 74236 3100 74276
rect 3140 74236 4244 74276
rect 4684 74236 4876 74276
rect 4916 74236 4925 74276
rect 5033 74236 5164 74276
rect 5204 74236 5213 74276
rect 5404 74236 6740 74276
rect 6796 74236 7220 74276
rect 7337 74236 7468 74276
rect 7508 74236 7517 74276
rect 7651 74236 7660 74276
rect 7700 74236 8188 74276
rect 8228 74236 8237 74276
rect 0 74024 90 74044
rect 0 73984 364 74024
rect 404 73984 413 74024
rect 0 73964 90 73984
rect 1987 73900 1996 73940
rect 2036 73900 4396 73940
rect 4436 73900 4445 73940
rect 3052 73816 3244 73856
rect 3284 73816 3293 73856
rect 3436 73816 3532 73856
rect 3572 73816 3581 73856
rect 3052 73772 3092 73816
rect 3436 73772 3476 73816
rect 4684 73772 4724 74236
rect 6796 74108 6836 74236
rect 10252 74108 10292 74404
rect 11500 74395 11540 74404
rect 13228 74395 13268 74404
rect 14188 74360 14228 74404
rect 14476 74360 14516 74404
rect 14860 74360 14900 74488
rect 15436 74444 15476 74453
rect 16060 74444 16100 74488
rect 17116 74479 17156 74656
rect 17836 74572 18452 74612
rect 17836 74528 17876 74572
rect 18412 74528 18452 74572
rect 20140 74528 20180 74740
rect 21510 74528 21600 74548
rect 17251 74488 17260 74528
rect 17300 74488 17347 74528
rect 17404 74488 17644 74528
rect 17684 74488 17693 74528
rect 17827 74488 17836 74528
rect 17876 74488 17885 74528
rect 17932 74488 18028 74528
rect 18068 74488 18077 74528
rect 18403 74488 18412 74528
rect 18452 74488 18461 74528
rect 20131 74488 20140 74528
rect 20180 74488 20189 74528
rect 20323 74488 20332 74528
rect 20372 74488 21600 74528
rect 17050 74470 17156 74479
rect 14947 74404 14956 74444
rect 14996 74404 15340 74444
rect 15380 74404 15389 74444
rect 15523 74404 15532 74444
rect 15572 74404 15924 74444
rect 15964 74404 15973 74444
rect 16060 74404 16396 74444
rect 16436 74404 16732 74444
rect 16772 74404 16781 74444
rect 16867 74404 16876 74444
rect 16916 74404 16925 74444
rect 17050 74430 17059 74470
rect 17099 74439 17156 74470
rect 17260 74444 17300 74488
rect 17404 74444 17444 74488
rect 17932 74444 17972 74488
rect 21510 74468 21600 74488
rect 18988 74444 19028 74453
rect 17099 74430 17108 74439
rect 17050 74429 17108 74430
rect 17242 74404 17251 74444
rect 17291 74404 17300 74444
rect 17347 74404 17356 74444
rect 17396 74404 17444 74444
rect 17539 74404 17548 74444
rect 17588 74404 17597 74444
rect 17914 74404 17923 74444
rect 17963 74404 17972 74444
rect 18019 74404 18028 74444
rect 18068 74404 18077 74444
rect 18348 74404 18412 74444
rect 18452 74404 18508 74444
rect 18548 74404 18892 74444
rect 18932 74404 18941 74444
rect 19498 74404 19507 74444
rect 19547 74404 19948 74444
rect 19988 74404 19997 74444
rect 13324 74320 13852 74360
rect 13892 74320 13901 74360
rect 14188 74320 14516 74360
rect 14563 74320 14572 74360
rect 14612 74320 14900 74360
rect 15436 74360 15476 74404
rect 16876 74360 16916 74404
rect 17356 74360 17396 74404
rect 15436 74320 15628 74360
rect 15668 74320 15677 74360
rect 16876 74320 17396 74360
rect 17548 74360 17588 74404
rect 17548 74320 17932 74360
rect 17972 74320 17981 74360
rect 13324 74276 13364 74320
rect 18028 74276 18068 74404
rect 13027 74236 13036 74276
rect 13076 74236 13364 74276
rect 13411 74236 13420 74276
rect 13460 74236 13804 74276
rect 13844 74236 13853 74276
rect 16099 74236 16108 74276
rect 16148 74236 16340 74276
rect 16570 74236 16579 74276
rect 16619 74236 17740 74276
rect 17780 74236 17789 74276
rect 17932 74236 18068 74276
rect 16300 74108 16340 74236
rect 17932 74192 17972 74236
rect 17059 74152 17068 74192
rect 17108 74152 17972 74192
rect 4919 74068 4928 74108
rect 4968 74068 5010 74108
rect 5050 74068 5092 74108
rect 5132 74068 5174 74108
rect 5214 74068 5256 74108
rect 5296 74068 5305 74108
rect 6604 74068 6836 74108
rect 8227 74068 8236 74108
rect 8276 74068 10292 74108
rect 15811 74068 15820 74108
rect 15860 74068 16340 74108
rect 6604 73940 6644 74068
rect 18988 74024 19028 74404
rect 19075 74236 19084 74276
rect 19124 74236 19660 74276
rect 19700 74236 19709 74276
rect 20371 74236 20380 74276
rect 20420 74236 21292 74276
rect 21332 74236 21341 74276
rect 20039 74068 20048 74108
rect 20088 74068 20130 74108
rect 20170 74068 20212 74108
rect 20252 74068 20294 74108
rect 20334 74068 20376 74108
rect 20416 74068 20425 74108
rect 21510 74024 21600 74044
rect 6979 73984 6988 74024
rect 7028 73984 8084 74024
rect 8131 73984 8140 74024
rect 8180 73984 14420 74024
rect 14659 73984 14668 74024
rect 14708 73984 15628 74024
rect 15668 73984 17780 74024
rect 17827 73984 17836 74024
rect 17876 73984 19028 74024
rect 21187 73984 21196 74024
rect 21236 73984 21600 74024
rect 8044 73940 8084 73984
rect 4771 73900 4780 73940
rect 4820 73900 5548 73940
rect 5588 73900 5597 73940
rect 6595 73900 6604 73940
rect 6644 73900 6653 73940
rect 6988 73900 7604 73940
rect 8044 73900 8660 73940
rect 6988 73856 7028 73900
rect 5347 73816 5356 73856
rect 5396 73816 7028 73856
rect 7075 73816 7084 73856
rect 7124 73816 7508 73856
rect 1315 73732 1324 73772
rect 1364 73732 2284 73772
rect 2324 73732 2333 73772
rect 2467 73732 2476 73772
rect 2516 73763 2647 73772
rect 2516 73732 2572 73763
rect 2612 73732 2647 73763
rect 3034 73732 3043 73772
rect 3083 73732 3092 73772
rect 3139 73732 3148 73772
rect 3188 73732 3476 73772
rect 3523 73732 3532 73772
rect 3572 73732 3581 73772
rect 4108 73763 4300 73772
rect 2572 73714 2612 73723
rect 0 73688 90 73708
rect 0 73648 268 73688
rect 308 73648 317 73688
rect 0 73628 90 73648
rect 3532 73604 3572 73732
rect 4148 73732 4300 73763
rect 4340 73732 4349 73772
rect 4457 73732 4588 73772
rect 4628 73732 4637 73772
rect 4684 73732 5164 73772
rect 5204 73732 5213 73772
rect 6211 73732 6220 73772
rect 6260 73763 6452 73772
rect 6260 73732 6412 73763
rect 4108 73714 4148 73723
rect 4588 73714 4628 73723
rect 6970 73732 6979 73772
rect 7019 73732 7180 73772
rect 7220 73732 7229 73772
rect 7363 73732 7372 73772
rect 7412 73732 7421 73772
rect 7468 73763 7508 73816
rect 6412 73714 6452 73723
rect 7372 73688 7412 73732
rect 7564 73772 7604 73900
rect 7747 73816 7756 73856
rect 7796 73816 8564 73856
rect 8524 73772 8564 73816
rect 7564 73732 7948 73772
rect 7988 73732 7997 73772
rect 8419 73732 8428 73772
rect 8468 73732 8477 73772
rect 8520 73732 8529 73772
rect 8569 73732 8578 73772
rect 7468 73714 7508 73723
rect 3619 73648 3628 73688
rect 3668 73648 4012 73688
rect 4052 73648 4061 73688
rect 6739 73648 6748 73688
rect 6788 73648 7412 73688
rect 7555 73648 7564 73688
rect 7604 73648 8044 73688
rect 8084 73648 8140 73688
rect 8180 73648 8244 73688
rect 3532 73564 8276 73604
rect 2755 73480 2764 73520
rect 2804 73480 4300 73520
rect 4340 73480 4349 73520
rect 8236 73436 8276 73564
rect 8428 73520 8468 73732
rect 8620 73688 8660 73900
rect 9100 73900 11500 73940
rect 11540 73900 11549 73940
rect 11875 73900 11884 73940
rect 11924 73900 12220 73940
rect 12260 73900 12269 73940
rect 9100 73772 9140 73900
rect 14380 73856 14420 73984
rect 14467 73900 14476 73940
rect 14516 73900 15436 73940
rect 15476 73900 15485 73940
rect 16483 73900 16492 73940
rect 16532 73900 17644 73940
rect 17684 73900 17693 73940
rect 17740 73856 17780 73984
rect 21510 73964 21600 73984
rect 18316 73900 19276 73940
rect 19316 73900 19325 73940
rect 18316 73856 18356 73900
rect 10252 73816 11116 73856
rect 11156 73816 11165 73856
rect 12067 73816 12076 73856
rect 12116 73816 12788 73856
rect 10252 73772 10292 73816
rect 12748 73772 12788 73816
rect 12844 73816 13708 73856
rect 13748 73816 13757 73856
rect 14380 73816 17548 73856
rect 17588 73816 17684 73856
rect 17740 73816 18356 73856
rect 18499 73816 18508 73856
rect 18548 73816 18740 73856
rect 18883 73816 18892 73856
rect 18932 73816 20372 73856
rect 12844 73772 12884 73816
rect 17644 73772 17684 73816
rect 18700 73772 18740 73816
rect 20332 73772 20372 73816
rect 8995 73732 9004 73772
rect 9044 73732 9140 73772
rect 10121 73732 10252 73772
rect 10292 73732 10301 73772
rect 10627 73732 10636 73772
rect 10676 73732 10685 73772
rect 11491 73732 11500 73772
rect 11540 73763 12596 73772
rect 11540 73732 11884 73763
rect 10636 73688 10676 73732
rect 11924 73732 12596 73763
rect 12730 73732 12739 73772
rect 12779 73732 12788 73772
rect 12835 73732 12844 73772
rect 12884 73732 12893 73772
rect 13132 73732 13228 73772
rect 13268 73732 13516 73772
rect 13556 73732 13565 73772
rect 13673 73732 13804 73772
rect 13844 73732 13853 73772
rect 14153 73732 14188 73772
rect 14228 73763 14324 73772
rect 14228 73732 14284 73763
rect 11884 73714 11924 73723
rect 12556 73688 12596 73732
rect 13132 73688 13172 73732
rect 13804 73714 13844 73723
rect 14371 73732 14380 73772
rect 14420 73732 15668 73772
rect 15811 73732 15820 73772
rect 15860 73732 15869 73772
rect 16265 73732 16396 73772
rect 16436 73732 16445 73772
rect 17644 73763 18124 73772
rect 14284 73714 14324 73723
rect 8620 73648 10676 73688
rect 11980 73648 12212 73688
rect 12329 73648 12460 73688
rect 12500 73648 12509 73688
rect 12556 73648 12748 73688
rect 12788 73648 12797 73688
rect 13123 73648 13132 73688
rect 13172 73648 13181 73688
rect 13289 73648 13324 73688
rect 13364 73648 13420 73688
rect 13460 73648 13469 73688
rect 14659 73648 14668 73688
rect 14708 73648 14860 73688
rect 14900 73648 14909 73688
rect 14969 73648 15052 73688
rect 15092 73648 15100 73688
rect 15140 73648 15149 73688
rect 15244 73648 15484 73688
rect 15524 73648 15533 73688
rect 8524 73564 10924 73604
rect 10964 73564 10973 73604
rect 8419 73480 8428 73520
rect 8468 73480 8477 73520
rect 8524 73436 8564 73564
rect 11980 73520 12020 73648
rect 12172 73604 12212 73648
rect 15244 73604 15284 73648
rect 15628 73604 15668 73732
rect 15820 73688 15860 73732
rect 17684 73732 18124 73763
rect 18164 73732 18173 73772
rect 18473 73732 18604 73772
rect 18644 73732 18653 73772
rect 18700 73763 19892 73772
rect 18700 73732 19852 73763
rect 17644 73714 17684 73723
rect 20323 73732 20332 73772
rect 20372 73732 20381 73772
rect 19852 73714 19892 73723
rect 15715 73648 15724 73688
rect 15764 73648 15860 73688
rect 15907 73648 15916 73688
rect 15956 73648 16087 73688
rect 18211 73648 18220 73688
rect 18260 73648 18269 73688
rect 18220 73604 18260 73648
rect 12067 73564 12076 73604
rect 12116 73564 12125 73604
rect 12172 73564 15284 73604
rect 15379 73564 15388 73604
rect 15428 73564 15572 73604
rect 15628 73564 18260 73604
rect 19651 73564 19660 73604
rect 19700 73564 20188 73604
rect 20228 73564 20237 73604
rect 20803 73564 20812 73604
rect 20852 73564 21236 73604
rect 8803 73480 8812 73520
rect 8852 73480 8908 73520
rect 8948 73480 8983 73520
rect 9091 73480 9100 73520
rect 9140 73480 12020 73520
rect 12076 73520 12116 73564
rect 15532 73520 15572 73564
rect 21196 73520 21236 73564
rect 21510 73520 21600 73540
rect 12076 73480 14620 73520
rect 14660 73480 14669 73520
rect 15532 73480 15628 73520
rect 15668 73480 15677 73520
rect 16147 73480 16156 73520
rect 16196 73480 16396 73520
rect 16436 73480 16445 73520
rect 17705 73480 17836 73520
rect 17876 73480 17885 73520
rect 18451 73480 18460 73520
rect 18500 73480 19700 73520
rect 19747 73480 19756 73520
rect 19796 73480 20044 73520
rect 20084 73480 20093 73520
rect 20140 73480 21140 73520
rect 21196 73480 21600 73520
rect 3331 73396 3340 73436
rect 3380 73396 5300 73436
rect 8236 73396 8564 73436
rect 19660 73436 19700 73480
rect 20140 73436 20180 73480
rect 19660 73396 20180 73436
rect 0 73352 90 73372
rect 5260 73352 5300 73396
rect 21100 73352 21140 73480
rect 21510 73460 21600 73480
rect 0 73312 364 73352
rect 404 73312 413 73352
rect 3679 73312 3688 73352
rect 3728 73312 3770 73352
rect 3810 73312 3852 73352
rect 3892 73312 3934 73352
rect 3974 73312 4016 73352
rect 4056 73312 4065 73352
rect 5251 73312 5260 73352
rect 5300 73312 5309 73352
rect 6700 73312 10060 73352
rect 10100 73312 10109 73352
rect 13795 73312 13804 73352
rect 13844 73312 17068 73352
rect 17108 73312 17117 73352
rect 18799 73312 18808 73352
rect 18848 73312 18890 73352
rect 18930 73312 18972 73352
rect 19012 73312 19054 73352
rect 19094 73312 19136 73352
rect 19176 73312 19185 73352
rect 20899 73312 20908 73352
rect 20948 73312 21140 73352
rect 0 73292 90 73312
rect 1324 73144 3340 73184
rect 3380 73144 3389 73184
rect 4819 73144 4828 73184
rect 4868 73144 5932 73184
rect 5972 73144 5981 73184
rect 0 73016 90 73036
rect 0 72976 76 73016
rect 116 72976 125 73016
rect 0 72956 90 72976
rect 1324 72932 1364 73144
rect 3820 73060 4628 73100
rect 2572 72932 2612 72941
rect 1315 72892 1324 72932
rect 1364 72892 1373 72932
rect 2441 72892 2572 72932
rect 2612 72892 2621 72932
rect 2825 72892 2956 72932
rect 2996 72892 3005 72932
rect 2572 72883 2612 72892
rect 3820 72848 3860 73060
rect 4588 73016 4628 73060
rect 6700 73016 6740 73312
rect 6787 73228 6796 73268
rect 6836 73228 14188 73268
rect 14228 73228 14237 73268
rect 17452 73228 19796 73268
rect 17452 73184 17492 73228
rect 6931 73144 6940 73184
rect 6980 73144 7084 73184
rect 7124 73144 7133 73184
rect 8131 73144 8140 73184
rect 8180 73144 8380 73184
rect 10819 73144 10828 73184
rect 10868 73144 14900 73184
rect 17443 73144 17452 73184
rect 17492 73144 17501 73184
rect 19145 73144 19267 73184
rect 19316 73144 19325 73184
rect 8340 73016 8380 73144
rect 11011 73060 11020 73100
rect 11060 73060 13556 73100
rect 4579 72976 4588 73016
rect 4628 72976 4637 73016
rect 6691 72976 6700 73016
rect 6740 72976 6749 73016
rect 8057 72976 8140 73016
rect 8180 72976 8188 73016
rect 8228 72976 8237 73016
rect 8322 72976 8331 73016
rect 8371 72976 8380 73016
rect 8428 72976 9100 73016
rect 9140 72976 9149 73016
rect 9580 72976 11500 73016
rect 11540 72976 11549 73016
rect 13289 72976 13324 73016
rect 13364 72976 13420 73016
rect 13460 72976 13469 73016
rect 4204 72932 4244 72941
rect 6220 72932 6260 72941
rect 7756 72932 7796 72941
rect 8428 72932 8468 72976
rect 9580 72932 9620 72976
rect 12268 72932 12308 72941
rect 13516 72932 13556 73060
rect 14860 73016 14900 73144
rect 15475 73060 15484 73100
rect 15524 73060 19028 73100
rect 19075 73060 19084 73100
rect 19124 73060 19508 73100
rect 14851 72976 14860 73016
rect 14900 72976 14909 73016
rect 15113 72976 15244 73016
rect 15284 72976 15293 73016
rect 15497 72976 15628 73016
rect 15668 72976 15677 73016
rect 13996 72932 14036 72941
rect 17260 72932 17300 72941
rect 18892 72932 18932 72941
rect 67 72808 76 72848
rect 116 72808 212 72848
rect 172 72764 212 72808
rect 2668 72808 3860 72848
rect 4012 72892 4204 72932
rect 4841 72892 4972 72932
rect 5012 72892 5548 72932
rect 5588 72892 5597 72932
rect 6089 72892 6220 72932
rect 6260 72892 6269 72932
rect 7258 72892 7267 72932
rect 7307 72892 7316 72932
rect 2668 72764 2708 72808
rect 4012 72764 4052 72892
rect 4204 72883 4244 72892
rect 6220 72883 6260 72892
rect 6499 72808 6508 72848
rect 6548 72808 7075 72848
rect 7115 72808 7124 72848
rect 7276 72764 7316 72892
rect 7796 72892 8468 72932
rect 8585 72892 8620 72932
rect 8660 72892 8716 72932
rect 8756 72892 8765 72932
rect 8825 72892 8834 72932
rect 8874 72892 8908 72932
rect 8948 72892 9014 72932
rect 10697 72892 10828 72932
rect 10868 72892 10877 72932
rect 11011 72892 11020 72932
rect 11060 72892 11191 72932
rect 11971 72892 11980 72932
rect 12020 72892 12172 72932
rect 12212 72892 12268 72932
rect 7756 72883 7796 72892
rect 9580 72883 9620 72892
rect 10828 72848 10868 72892
rect 12268 72883 12308 72892
rect 12460 72892 12931 72932
rect 12971 72892 12980 72932
rect 13027 72892 13036 72932
rect 13076 72892 13132 72932
rect 13172 72892 13207 72932
rect 13507 72892 13516 72932
rect 13556 72892 13565 72932
rect 13795 72892 13804 72932
rect 13844 72892 13996 72932
rect 14506 72892 14515 72932
rect 14555 72892 14804 72932
rect 15907 72892 15916 72932
rect 15956 72892 16012 72932
rect 16052 72892 16087 72932
rect 17635 72892 17644 72932
rect 17684 72892 18412 72932
rect 18452 72892 18461 72932
rect 12460 72848 12500 72892
rect 13996 72883 14036 72892
rect 10828 72808 11308 72848
rect 11348 72808 11357 72848
rect 12451 72808 12460 72848
rect 12500 72808 12509 72848
rect 172 72724 2708 72764
rect 2755 72724 2764 72764
rect 2804 72724 3052 72764
rect 3092 72724 3101 72764
rect 3427 72724 3436 72764
rect 3476 72724 4052 72764
rect 4265 72724 4396 72764
rect 4436 72724 4445 72764
rect 6115 72724 6124 72764
rect 6164 72724 6412 72764
rect 6452 72724 6461 72764
rect 7276 72724 9388 72764
rect 9428 72724 9437 72764
rect 9763 72724 9772 72764
rect 9812 72724 14420 72764
rect 14537 72724 14668 72764
rect 14708 72724 14717 72764
rect 0 72680 90 72700
rect 0 72640 748 72680
rect 788 72640 797 72680
rect 9379 72640 9388 72680
rect 9428 72640 11020 72680
rect 11060 72640 11069 72680
rect 0 72620 90 72640
rect 4919 72556 4928 72596
rect 4968 72556 5010 72596
rect 5050 72556 5092 72596
rect 5132 72556 5174 72596
rect 5214 72556 5256 72596
rect 5296 72556 5305 72596
rect 7267 72556 7276 72596
rect 7316 72556 10636 72596
rect 10676 72556 10685 72596
rect 14380 72512 14420 72724
rect 14764 72596 14804 72892
rect 17260 72848 17300 72892
rect 18892 72848 18932 72892
rect 15091 72808 15100 72848
rect 15140 72808 17164 72848
rect 17204 72808 17213 72848
rect 17260 72808 17932 72848
rect 17972 72808 17981 72848
rect 18307 72808 18316 72848
rect 18356 72808 18508 72848
rect 18548 72808 18932 72848
rect 18988 72848 19028 73060
rect 19075 72892 19084 72932
rect 19124 72892 19267 72932
rect 19307 72892 19316 72932
rect 19363 72903 19372 72943
rect 19412 72903 19421 72943
rect 19468 72932 19508 73060
rect 19651 72976 19660 73016
rect 19700 72976 19709 73016
rect 19660 72932 19700 72976
rect 18988 72808 19180 72848
rect 19220 72808 19229 72848
rect 15859 72724 15868 72764
rect 15908 72724 17260 72764
rect 17300 72724 17309 72764
rect 17443 72724 17452 72764
rect 17492 72724 17644 72764
rect 17684 72724 17693 72764
rect 18028 72724 18836 72764
rect 18953 72724 19084 72764
rect 19124 72724 19133 72764
rect 18028 72596 18068 72724
rect 18796 72680 18836 72724
rect 19372 72680 19412 72903
rect 19468 72892 19517 72932
rect 19557 72892 19566 72932
rect 19613 72892 19647 72932
rect 19687 72892 19700 72932
rect 19756 72943 19796 73228
rect 20140 73144 21484 73184
rect 21524 73144 21533 73184
rect 20140 73016 20180 73144
rect 21510 73016 21600 73036
rect 20131 72976 20140 73016
rect 20180 72976 20189 73016
rect 21091 72976 21100 73016
rect 21140 72976 21600 73016
rect 21510 72956 21600 72976
rect 19756 72903 19777 72943
rect 19817 72903 19826 72943
rect 20371 72724 20380 72764
rect 20420 72724 21484 72764
rect 21524 72724 21533 72764
rect 18796 72640 19412 72680
rect 14659 72556 14668 72596
rect 14708 72556 14804 72596
rect 17164 72556 18068 72596
rect 20039 72556 20048 72596
rect 20088 72556 20130 72596
rect 20170 72556 20212 72596
rect 20252 72556 20294 72596
rect 20334 72556 20376 72596
rect 20416 72556 20425 72596
rect 172 72472 940 72512
rect 980 72472 989 72512
rect 1699 72472 1708 72512
rect 1748 72472 13132 72512
rect 13172 72472 13181 72512
rect 14380 72472 16724 72512
rect 0 72344 90 72364
rect 0 72302 116 72344
rect 172 72302 212 72472
rect 3436 72388 6796 72428
rect 6836 72388 6845 72428
rect 6979 72388 6988 72428
rect 7028 72388 8564 72428
rect 9187 72388 9196 72428
rect 9236 72388 10492 72428
rect 10532 72388 10541 72428
rect 11251 72388 11260 72428
rect 11300 72388 11500 72428
rect 11540 72388 11549 72428
rect 14659 72388 14668 72428
rect 14708 72388 15052 72428
rect 15092 72388 15101 72428
rect 3436 72344 3476 72388
rect 931 72304 940 72344
rect 980 72304 2332 72344
rect 2372 72304 2381 72344
rect 2572 72304 3476 72344
rect 3523 72304 3532 72344
rect 3572 72304 5116 72344
rect 5156 72304 5165 72344
rect 5491 72304 5500 72344
rect 5540 72304 5644 72344
rect 5684 72304 5693 72344
rect 0 72284 212 72302
rect 76 72262 212 72284
rect 1420 72220 1708 72260
rect 1748 72220 1757 72260
rect 1420 72176 1460 72220
rect 2572 72176 2612 72304
rect 2659 72220 2668 72260
rect 2708 72220 2851 72260
rect 2891 72220 2900 72260
rect 2947 72220 2956 72260
rect 2996 72220 3127 72260
rect 3209 72220 3340 72260
rect 3380 72220 3389 72260
rect 3916 72251 3956 72260
rect 4265 72220 4300 72260
rect 4340 72251 4436 72260
rect 4340 72220 4396 72251
rect 3916 72176 3956 72211
rect 4618 72220 4627 72260
rect 4667 72220 5396 72260
rect 6115 72220 6124 72260
rect 6164 72220 6286 72260
rect 6326 72220 6335 72260
rect 6403 72220 6412 72260
rect 6452 72220 6461 72260
rect 6691 72220 6700 72260
rect 6740 72220 6796 72260
rect 6836 72220 6871 72260
rect 7241 72220 7372 72260
rect 7412 72220 7421 72260
rect 7721 72220 7852 72260
rect 7892 72220 7901 72260
rect 4396 72202 4436 72211
rect 5356 72176 5396 72220
rect 6412 72176 6452 72220
rect 7372 72202 7412 72211
rect 7852 72202 7892 72211
rect 8524 72176 8564 72388
rect 8611 72304 8620 72344
rect 8660 72304 10108 72344
rect 10148 72304 10157 72344
rect 11971 72304 11980 72344
rect 12020 72304 14900 72344
rect 9763 72220 9772 72260
rect 9812 72220 10388 72260
rect 10819 72220 10828 72260
rect 10868 72220 11980 72260
rect 12020 72220 12029 72260
rect 12835 72220 12844 72260
rect 12884 72251 13268 72260
rect 12884 72220 13228 72251
rect 10348 72176 10388 72220
rect 13603 72220 13612 72260
rect 13652 72220 14668 72260
rect 14708 72220 14717 72260
rect 14860 72251 14900 72304
rect 16684 72260 16724 72472
rect 17164 72428 17204 72556
rect 21510 72512 21600 72532
rect 18595 72472 18604 72512
rect 18644 72472 20180 72512
rect 20995 72472 21004 72512
rect 21044 72472 21600 72512
rect 20140 72428 20180 72472
rect 21510 72452 21600 72472
rect 17146 72388 17155 72428
rect 17195 72388 17204 72428
rect 17251 72388 17260 72428
rect 17300 72388 17972 72428
rect 20131 72388 20140 72428
rect 20180 72388 20189 72428
rect 17932 72344 17972 72388
rect 17539 72304 17548 72344
rect 17588 72304 17876 72344
rect 17932 72304 20332 72344
rect 20372 72304 20381 72344
rect 17836 72260 17876 72304
rect 13228 72202 13268 72211
rect 14947 72220 14956 72260
rect 14996 72220 15244 72260
rect 15284 72220 15293 72260
rect 15811 72220 15820 72260
rect 15860 72220 16396 72260
rect 16436 72251 16567 72260
rect 16436 72220 16492 72251
rect 14860 72202 14900 72211
rect 16532 72220 16567 72251
rect 16684 72220 17308 72260
rect 17348 72220 17357 72260
rect 17443 72220 17452 72260
rect 17492 72220 17644 72260
rect 17684 72220 17693 72260
rect 17818 72220 17827 72260
rect 17867 72220 17876 72260
rect 17923 72220 17932 72260
rect 17972 72220 18164 72260
rect 18251 72220 18316 72260
rect 18356 72220 18382 72260
rect 18422 72220 18431 72260
rect 18504 72220 18513 72260
rect 18553 72220 18562 72260
rect 18787 72220 18796 72260
rect 18836 72220 18892 72260
rect 18932 72220 18967 72260
rect 19075 72220 19084 72260
rect 19124 72251 19508 72260
rect 19124 72220 19468 72251
rect 16492 72202 16532 72211
rect 259 72136 268 72176
rect 308 72136 1364 72176
rect 1411 72136 1420 72176
rect 1460 72136 1469 72176
rect 1795 72136 1804 72176
rect 1844 72136 2132 72176
rect 2179 72136 2188 72176
rect 2228 72136 2237 72176
rect 2563 72136 2572 72176
rect 2612 72136 2621 72176
rect 3427 72136 3436 72176
rect 3476 72136 3628 72176
rect 3668 72136 3677 72176
rect 3916 72136 4204 72176
rect 4244 72136 4253 72176
rect 4579 72136 4588 72176
rect 4628 72136 4732 72176
rect 4772 72136 4781 72176
rect 4963 72136 4972 72176
rect 5012 72136 5164 72176
rect 5204 72136 5213 72176
rect 5347 72136 5356 72176
rect 5396 72136 5405 72176
rect 5609 72136 5740 72176
rect 5780 72136 5789 72176
rect 5923 72136 5932 72176
rect 5972 72136 6452 72176
rect 6761 72136 6892 72176
rect 6932 72136 6941 72176
rect 8074 72136 8083 72176
rect 8123 72136 8428 72176
rect 8468 72136 8477 72176
rect 8524 72136 8620 72176
rect 8660 72136 8669 72176
rect 8716 72136 8956 72176
rect 8996 72136 9005 72176
rect 9065 72136 9196 72176
rect 9236 72136 9245 72176
rect 9379 72136 9388 72176
rect 9428 72136 9559 72176
rect 9833 72136 9964 72176
rect 10004 72136 10013 72176
rect 10339 72136 10348 72176
rect 10388 72136 10397 72176
rect 10601 72136 10636 72176
rect 10676 72136 10732 72176
rect 10772 72136 10781 72176
rect 11203 72136 11212 72176
rect 11252 72136 11500 72176
rect 11540 72136 11549 72176
rect 1324 72092 1364 72136
rect 355 72052 364 72092
rect 404 72052 1180 72092
rect 1220 72052 1229 72092
rect 1324 72052 1564 72092
rect 1604 72052 1613 72092
rect 1699 72052 1708 72092
rect 1748 72052 1948 72092
rect 1988 72052 1997 72092
rect 0 72008 90 72028
rect 2092 72008 2132 72136
rect 2188 72092 2228 72136
rect 8716 72092 8756 72136
rect 2188 72052 8188 72092
rect 8228 72052 8237 72092
rect 8611 72052 8620 72092
rect 8660 72052 8756 72092
rect 8851 72052 8860 72092
rect 8900 72052 8908 72092
rect 8948 72052 9100 72092
rect 9140 72052 9149 72092
rect 9619 72052 9628 72092
rect 9668 72052 17164 72092
rect 17204 72052 17213 72092
rect 17308 72008 17348 72220
rect 18124 72176 18164 72220
rect 18508 72176 18548 72220
rect 19817 72220 19948 72260
rect 19988 72220 19997 72260
rect 19468 72202 19508 72211
rect 19948 72202 19988 72211
rect 18115 72136 18124 72176
rect 18164 72136 18548 72176
rect 18979 72136 18988 72176
rect 19028 72136 19037 72176
rect 17923 72052 17932 72092
rect 17972 72052 18892 72092
rect 18932 72052 18941 72092
rect 18988 72008 19028 72136
rect 21510 72008 21600 72028
rect 0 71968 556 72008
rect 596 71968 605 72008
rect 2092 71968 2380 72008
rect 2420 71968 2429 72008
rect 6595 71968 6604 72008
rect 6644 71968 9724 72008
rect 9764 71968 9773 72008
rect 13289 71968 13420 72008
rect 13460 71968 13469 72008
rect 14659 71968 14668 72008
rect 14708 71968 14956 72008
rect 14996 71968 15005 72008
rect 16553 71968 16684 72008
rect 16724 71968 16733 72008
rect 17308 71968 19028 72008
rect 19075 71968 19084 72008
rect 19124 71968 19316 72008
rect 21091 71968 21100 72008
rect 21140 71968 21600 72008
rect 0 71948 90 71968
rect 14668 71924 14708 71968
rect 18412 71924 18452 71968
rect 2179 71884 2188 71924
rect 2228 71884 5780 71924
rect 9283 71884 9292 71924
rect 9332 71884 14708 71924
rect 18403 71884 18412 71924
rect 18452 71884 18528 71924
rect 5740 71840 5780 71884
rect 3679 71800 3688 71840
rect 3728 71800 3770 71840
rect 3810 71800 3852 71840
rect 3892 71800 3934 71840
rect 3974 71800 4016 71840
rect 4056 71800 4065 71840
rect 5740 71800 12076 71840
rect 12116 71800 12125 71840
rect 12940 71800 15628 71840
rect 15668 71800 15677 71840
rect 18799 71800 18808 71840
rect 18848 71800 18890 71840
rect 18930 71800 18972 71840
rect 19012 71800 19054 71840
rect 19094 71800 19136 71840
rect 19176 71800 19185 71840
rect 12940 71756 12980 71800
rect 19276 71756 19316 71968
rect 21510 71948 21600 71968
rect 7756 71716 12980 71756
rect 19180 71716 19316 71756
rect 0 71672 90 71692
rect 0 71632 1228 71672
rect 1268 71632 1277 71672
rect 2131 71632 2140 71672
rect 2180 71632 7660 71672
rect 7700 71632 7709 71672
rect 0 71612 90 71632
rect 7756 71588 7796 71716
rect 19180 71672 19220 71716
rect 7843 71632 7852 71672
rect 7892 71632 8140 71672
rect 8180 71632 8189 71672
rect 15523 71632 15532 71672
rect 15572 71632 19220 71672
rect 1420 71548 7796 71588
rect 7852 71548 12172 71588
rect 12212 71548 12500 71588
rect 1420 71504 1460 71548
rect 7852 71504 7892 71548
rect 12460 71504 12500 71548
rect 12940 71548 14572 71588
rect 14612 71548 14621 71588
rect 14764 71548 15436 71588
rect 15476 71548 15485 71588
rect 16387 71548 16396 71588
rect 16436 71548 17684 71588
rect 1411 71464 1420 71504
rect 1460 71464 1469 71504
rect 1699 71464 1708 71504
rect 1748 71464 1900 71504
rect 1940 71464 1949 71504
rect 2275 71464 2284 71504
rect 2324 71464 2476 71504
rect 2516 71464 2525 71504
rect 2572 71464 2860 71504
rect 2900 71464 2909 71504
rect 3331 71464 3340 71504
rect 3380 71464 3511 71504
rect 3916 71464 4588 71504
rect 4628 71464 5260 71504
rect 5300 71464 5309 71504
rect 6124 71464 7892 71504
rect 9868 71464 10348 71504
rect 10388 71464 10397 71504
rect 12451 71464 12460 71504
rect 12500 71464 12509 71504
rect 1900 71420 1940 71464
rect 2572 71420 2612 71464
rect 3916 71420 3956 71464
rect 6028 71420 6068 71429
rect 1900 71380 2612 71420
rect 2699 71380 2764 71420
rect 2804 71380 2830 71420
rect 2870 71380 2879 71420
rect 2947 71380 2956 71420
rect 2996 71380 3005 71420
rect 3427 71380 3436 71420
rect 3476 71380 3820 71420
rect 3860 71380 3869 71420
rect 4099 71380 4108 71420
rect 4148 71380 4404 71420
rect 4444 71380 4453 71420
rect 4771 71380 4780 71420
rect 4820 71380 5548 71420
rect 5588 71380 5597 71420
rect 0 71336 90 71356
rect 2380 71336 2420 71380
rect 2956 71336 2996 71380
rect 3916 71371 3956 71380
rect 6028 71336 6068 71380
rect 0 71296 2284 71336
rect 2324 71296 2333 71336
rect 2380 71296 2524 71336
rect 2564 71296 2573 71336
rect 2956 71296 3724 71336
rect 3764 71296 3773 71336
rect 4492 71296 5932 71336
rect 5972 71296 6068 71336
rect 0 71276 90 71296
rect 4492 71252 4532 71296
rect 547 71212 556 71252
rect 596 71212 1180 71252
rect 1220 71212 1229 71252
rect 2860 71212 4532 71252
rect 4579 71212 4588 71252
rect 4628 71212 5740 71252
rect 5780 71212 5789 71252
rect 2860 71084 2900 71212
rect 6124 71168 6164 71464
rect 7948 71420 7988 71429
rect 9868 71420 9908 71464
rect 11500 71420 11540 71429
rect 12940 71420 12980 71548
rect 14764 71504 14804 71548
rect 17644 71504 17684 71548
rect 13738 71464 13747 71504
rect 13787 71464 14092 71504
rect 14132 71464 14141 71504
rect 14755 71464 14764 71504
rect 14804 71464 14813 71504
rect 15401 71464 15532 71504
rect 15572 71464 15581 71504
rect 17129 71464 17260 71504
rect 17300 71464 17309 71504
rect 17635 71464 17644 71504
rect 17684 71464 17693 71504
rect 18499 71464 18508 71504
rect 18548 71464 18604 71504
rect 18644 71464 18679 71504
rect 13036 71420 13076 71429
rect 16108 71420 16148 71429
rect 19180 71420 19220 71632
rect 21510 71504 21600 71524
rect 19939 71464 19948 71504
rect 19988 71464 20140 71504
rect 20180 71464 20189 71504
rect 20323 71464 20332 71504
rect 20372 71464 21600 71504
rect 21510 71444 21600 71464
rect 6595 71380 6604 71420
rect 6644 71380 6700 71420
rect 6740 71380 6775 71420
rect 7913 71380 7948 71420
rect 7988 71380 8044 71420
rect 8084 71380 8093 71420
rect 8585 71380 8620 71420
rect 8660 71380 8716 71420
rect 8756 71380 8765 71420
rect 10121 71380 10252 71420
rect 10292 71380 10636 71420
rect 10676 71380 10685 71420
rect 11369 71380 11500 71420
rect 11540 71380 11549 71420
rect 11692 71380 11971 71420
rect 12011 71380 12020 71420
rect 12067 71380 12076 71420
rect 12116 71380 12247 71420
rect 12547 71380 12556 71420
rect 12596 71380 12844 71420
rect 12884 71380 12980 71420
rect 13027 71380 13036 71420
rect 13076 71380 13207 71420
rect 13411 71380 13420 71420
rect 13460 71380 13524 71420
rect 13564 71380 13591 71420
rect 15034 71380 15043 71420
rect 15083 71380 15092 71420
rect 15139 71380 15148 71420
rect 15188 71380 15197 71420
rect 15331 71380 15340 71420
rect 15380 71380 15628 71420
rect 15668 71380 15677 71420
rect 15811 71380 15820 71420
rect 15860 71380 16108 71420
rect 16148 71380 16157 71420
rect 16553 71380 16627 71420
rect 16667 71380 16684 71420
rect 16724 71380 16733 71420
rect 17827 71380 17836 71420
rect 17876 71380 18115 71420
rect 18155 71380 18164 71420
rect 18211 71380 18220 71420
rect 18260 71380 18269 71420
rect 18403 71380 18412 71420
rect 18452 71380 18700 71420
rect 18740 71380 18749 71420
rect 19690 71380 19699 71420
rect 19739 71380 19756 71420
rect 19796 71380 19879 71420
rect 7948 71336 7988 71380
rect 9868 71371 9908 71380
rect 11500 71371 11540 71380
rect 11692 71336 11732 71380
rect 13036 71336 13076 71380
rect 6211 71296 6220 71336
rect 6260 71296 7988 71336
rect 11683 71296 11692 71336
rect 11732 71296 11741 71336
rect 13036 71296 13324 71336
rect 13364 71296 13373 71336
rect 6211 71212 6220 71252
rect 6260 71212 6269 71252
rect 10051 71212 10060 71252
rect 10100 71212 12844 71252
rect 12884 71212 12893 71252
rect 13411 71212 13420 71252
rect 13460 71212 13852 71252
rect 13892 71212 13901 71252
rect 14515 71212 14524 71252
rect 14564 71212 14572 71252
rect 14612 71212 14695 71252
rect 2563 71044 2572 71084
rect 2612 71044 2900 71084
rect 4012 71128 6164 71168
rect 0 71000 90 71020
rect 4012 71000 4052 71128
rect 6220 71084 6260 71212
rect 7651 71128 7660 71168
rect 7700 71128 13804 71168
rect 13844 71128 13853 71168
rect 15052 71084 15092 71380
rect 15148 71336 15188 71380
rect 16108 71371 16148 71380
rect 18220 71336 18260 71380
rect 15148 71296 15532 71336
rect 15572 71296 15581 71336
rect 18115 71296 18124 71336
rect 18164 71296 18260 71336
rect 16771 71212 16780 71252
rect 16820 71212 16829 71252
rect 17491 71212 17500 71252
rect 17540 71212 17549 71252
rect 17875 71212 17884 71252
rect 17924 71212 18988 71252
rect 19028 71212 19037 71252
rect 4919 71044 4928 71084
rect 4968 71044 5010 71084
rect 5050 71044 5092 71084
rect 5132 71044 5174 71084
rect 5214 71044 5256 71084
rect 5296 71044 5305 71084
rect 6019 71044 6028 71084
rect 6068 71044 6260 71084
rect 6940 71044 10100 71084
rect 15052 71044 15332 71084
rect 0 70960 1228 71000
rect 1268 70960 1277 71000
rect 2083 70960 2092 71000
rect 2132 70960 4052 71000
rect 0 70940 90 70960
rect 6940 70916 6980 71044
rect 10060 71000 10100 71044
rect 10060 70960 13036 71000
rect 13076 70960 13085 71000
rect 15292 70916 15332 71044
rect 1123 70876 1132 70916
rect 1172 70876 1564 70916
rect 1604 70876 1613 70916
rect 3820 70876 6980 70916
rect 7337 70876 7468 70916
rect 7508 70876 7517 70916
rect 11971 70876 11980 70916
rect 12020 70876 13420 70916
rect 13460 70876 13469 70916
rect 15235 70876 15244 70916
rect 15284 70876 15332 70916
rect 739 70708 748 70748
rect 788 70708 797 70748
rect 1987 70708 1996 70748
rect 2036 70708 2764 70748
rect 2804 70708 2813 70748
rect 3244 70739 3436 70748
rect 0 70664 90 70684
rect 748 70664 788 70708
rect 3284 70708 3436 70739
rect 3476 70708 3764 70748
rect 3244 70690 3284 70699
rect 0 70624 788 70664
rect 1289 70624 1420 70664
rect 1460 70624 1469 70664
rect 1795 70624 1804 70664
rect 1844 70624 2668 70664
rect 2708 70624 2717 70664
rect 0 70604 90 70624
rect 3724 70580 3764 70708
rect 3820 70664 3860 70876
rect 16780 70832 16820 71212
rect 17500 71000 17540 71212
rect 19180 71168 19220 71380
rect 19843 71212 19852 71252
rect 19892 71212 20044 71252
rect 20084 71212 20093 71252
rect 20371 71212 20380 71252
rect 20420 71212 21100 71252
rect 21140 71212 21149 71252
rect 19180 71128 19756 71168
rect 19796 71128 19805 71168
rect 20039 71044 20048 71084
rect 20088 71044 20130 71084
rect 20170 71044 20212 71084
rect 20252 71044 20294 71084
rect 20334 71044 20376 71084
rect 20416 71044 20425 71084
rect 21510 71000 21600 71020
rect 17500 70960 18836 71000
rect 19267 70960 19276 71000
rect 19316 70960 21600 71000
rect 18796 70916 18836 70960
rect 21510 70940 21600 70960
rect 17539 70876 17548 70916
rect 17588 70876 18364 70916
rect 18404 70876 18413 70916
rect 18796 70876 20332 70916
rect 20372 70876 20381 70916
rect 4349 70792 4396 70832
rect 4436 70792 4445 70832
rect 4972 70792 6796 70832
rect 6836 70792 6845 70832
rect 7171 70792 7180 70832
rect 7220 70792 9524 70832
rect 10915 70792 10924 70832
rect 10964 70792 11732 70832
rect 4396 70748 4436 70792
rect 4378 70708 4387 70748
rect 4427 70708 4436 70748
rect 4483 70708 4492 70748
rect 4532 70708 4541 70748
rect 4745 70708 4876 70748
rect 4916 70708 4925 70748
rect 4492 70664 4532 70708
rect 4972 70664 5012 70792
rect 9484 70748 9524 70792
rect 11692 70748 11732 70792
rect 11788 70792 12076 70832
rect 12116 70792 12125 70832
rect 12451 70792 12460 70832
rect 12500 70792 16148 70832
rect 16780 70792 17204 70832
rect 18979 70792 18988 70832
rect 19028 70792 20428 70832
rect 20468 70792 20477 70832
rect 11788 70748 11828 70792
rect 16108 70748 16148 70792
rect 5452 70739 5492 70748
rect 5897 70739 6028 70748
rect 5897 70708 5932 70739
rect 3811 70624 3820 70664
rect 3860 70624 3869 70664
rect 4291 70624 4300 70664
rect 4340 70624 4532 70664
rect 4963 70624 4972 70664
rect 5012 70624 5021 70664
rect 739 70540 748 70580
rect 788 70540 1180 70580
rect 1220 70540 1229 70580
rect 1420 70540 3580 70580
rect 3620 70540 3629 70580
rect 3724 70540 4108 70580
rect 4148 70540 4157 70580
rect 1420 70496 1460 70540
rect 1411 70456 1420 70496
rect 1460 70456 1469 70496
rect 3427 70456 3436 70496
rect 3476 70456 4300 70496
rect 4340 70456 4349 70496
rect 5452 70412 5492 70699
rect 5972 70708 6028 70739
rect 6068 70708 6077 70748
rect 7171 70708 7180 70748
rect 7220 70708 7229 70748
rect 7313 70708 7322 70748
rect 7362 70708 7372 70748
rect 7412 70708 7502 70748
rect 7852 70739 7892 70748
rect 5932 70690 5972 70699
rect 7180 70664 7220 70708
rect 9091 70708 9100 70748
rect 9140 70708 9292 70748
rect 9332 70708 9341 70748
rect 9475 70708 9484 70748
rect 9524 70708 9533 70748
rect 9763 70708 9772 70748
rect 9812 70708 10348 70748
rect 10388 70739 10772 70748
rect 10388 70708 10732 70739
rect 7852 70664 7892 70699
rect 9772 70664 9812 70708
rect 6028 70624 6316 70664
rect 6356 70624 6365 70664
rect 6508 70624 6892 70664
rect 6932 70624 6941 70664
rect 7180 70624 7276 70664
rect 7316 70624 7325 70664
rect 7852 70624 9812 70664
rect 11674 70708 11683 70748
rect 11723 70708 11732 70748
rect 11779 70708 11788 70748
rect 11828 70708 11837 70748
rect 12041 70708 12172 70748
rect 12212 70708 12221 70748
rect 12748 70739 13132 70748
rect 10732 70664 10772 70699
rect 12788 70708 13132 70739
rect 13172 70708 13181 70748
rect 13228 70739 13268 70748
rect 12748 70690 12788 70699
rect 13603 70708 13612 70748
rect 13652 70708 13804 70748
rect 13844 70708 13853 70748
rect 14563 70708 14572 70748
rect 14612 70739 15724 70748
rect 14612 70708 15052 70739
rect 13228 70664 13268 70699
rect 15092 70708 15724 70739
rect 15764 70708 15773 70748
rect 16099 70708 16108 70748
rect 16148 70708 17068 70748
rect 17108 70708 17117 70748
rect 15052 70690 15092 70699
rect 17164 70664 17204 70792
rect 17251 70708 17260 70748
rect 17300 70739 17932 70748
rect 17300 70708 17356 70739
rect 17396 70708 17932 70739
rect 17972 70708 17981 70748
rect 18211 70708 18220 70748
rect 18260 70708 18796 70748
rect 18836 70708 19276 70748
rect 19316 70708 19325 70748
rect 20044 70739 20084 70748
rect 17356 70690 17396 70699
rect 20044 70664 20084 70699
rect 10732 70624 11068 70664
rect 11108 70624 11117 70664
rect 11203 70624 11212 70664
rect 11252 70624 11308 70664
rect 11348 70624 11383 70664
rect 12259 70624 12268 70664
rect 12308 70624 12706 70664
rect 12835 70624 12844 70664
rect 12884 70624 13268 70664
rect 15907 70624 15916 70664
rect 15956 70624 17204 70664
rect 17897 70624 18028 70664
rect 18068 70624 18077 70664
rect 18473 70624 18604 70664
rect 18644 70624 18653 70664
rect 18700 70624 20084 70664
rect 6028 70580 6068 70624
rect 6508 70580 6548 70624
rect 12666 70580 12706 70624
rect 18700 70580 18740 70624
rect 5932 70540 6068 70580
rect 6163 70540 6172 70580
rect 6212 70540 6548 70580
rect 6595 70540 6604 70580
rect 6644 70540 6652 70580
rect 6692 70540 6775 70580
rect 12666 70540 12980 70580
rect 13027 70540 13036 70580
rect 13076 70540 15676 70580
rect 15716 70540 15725 70580
rect 18259 70540 18268 70580
rect 18308 70540 18508 70580
rect 18548 70540 18557 70580
rect 18604 70540 18740 70580
rect 19843 70540 19852 70580
rect 19892 70540 20236 70580
rect 20276 70540 20285 70580
rect 5932 70496 5972 70540
rect 12940 70496 12980 70540
rect 18604 70496 18644 70540
rect 21510 70496 21600 70516
rect 5731 70456 5740 70496
rect 5780 70456 5972 70496
rect 6019 70456 6028 70496
rect 6068 70456 6556 70496
rect 6596 70456 6605 70496
rect 7171 70456 7180 70496
rect 7220 70456 7660 70496
rect 7700 70456 7709 70496
rect 12940 70456 13228 70496
rect 13268 70456 13277 70496
rect 17417 70456 17548 70496
rect 17588 70456 17597 70496
rect 17827 70456 17836 70496
rect 17876 70456 18644 70496
rect 18700 70456 21600 70496
rect 18700 70412 18740 70456
rect 21510 70436 21600 70456
rect 4867 70372 4876 70412
rect 4916 70372 9004 70412
rect 9044 70372 9053 70412
rect 11491 70372 11500 70412
rect 11540 70372 14764 70412
rect 14804 70372 15436 70412
rect 15476 70372 15485 70412
rect 17347 70372 17356 70412
rect 17396 70372 18740 70412
rect 0 70328 90 70348
rect 0 70288 172 70328
rect 212 70288 221 70328
rect 3679 70288 3688 70328
rect 3728 70288 3770 70328
rect 3810 70288 3852 70328
rect 3892 70288 3934 70328
rect 3974 70288 4016 70328
rect 4056 70288 4065 70328
rect 12940 70288 16396 70328
rect 16436 70288 16445 70328
rect 18799 70288 18808 70328
rect 18848 70288 18890 70328
rect 18930 70288 18972 70328
rect 19012 70288 19054 70328
rect 19094 70288 19136 70328
rect 19176 70288 19185 70328
rect 19651 70288 19660 70328
rect 19700 70288 21575 70328
rect 0 70268 90 70288
rect 2860 70204 9196 70244
rect 9236 70204 9245 70244
rect 2860 70160 2900 70204
rect 12940 70160 12980 70288
rect 16099 70204 16108 70244
rect 16148 70204 17164 70244
rect 17204 70204 17213 70244
rect 21535 70160 21575 70288
rect 76 70120 2900 70160
rect 6892 70120 8140 70160
rect 8180 70120 8189 70160
rect 12595 70120 12604 70160
rect 12644 70120 12980 70160
rect 16003 70120 16012 70160
rect 16052 70120 16060 70160
rect 16100 70120 16183 70160
rect 17321 70120 17404 70160
rect 17444 70120 17452 70160
rect 17492 70120 17501 70160
rect 18787 70120 18796 70160
rect 18836 70120 19756 70160
rect 19796 70120 19805 70160
rect 21388 70120 21575 70160
rect 76 70012 116 70120
rect 0 69952 116 70012
rect 3532 70036 4492 70076
rect 4532 70036 4541 70076
rect 4675 70036 4684 70076
rect 4724 70036 5396 70076
rect 3532 69992 3572 70036
rect 3523 69952 3532 69992
rect 3572 69952 3581 69992
rect 0 69932 90 69952
rect 2764 69908 2804 69917
rect 3916 69908 3956 69917
rect 5356 69908 5396 70036
rect 6604 69908 6644 69917
rect 6892 69908 6932 70120
rect 7555 70036 7564 70076
rect 7604 70036 7796 70076
rect 13699 70036 13708 70076
rect 13748 70036 16732 70076
rect 16772 70036 16781 70076
rect 16972 70036 19660 70076
rect 19700 70036 19709 70076
rect 7660 69908 7700 69917
rect 1507 69868 1516 69908
rect 1556 69868 1708 69908
rect 1748 69868 1757 69908
rect 2563 69868 2572 69908
rect 2612 69868 2764 69908
rect 2851 69868 2860 69908
rect 2900 69868 3916 69908
rect 4963 69868 4972 69908
rect 5012 69868 5164 69908
rect 5204 69868 5213 69908
rect 5347 69868 5356 69908
rect 5396 69868 5405 69908
rect 6644 69868 6892 69908
rect 6932 69868 6941 69908
rect 7049 69868 7171 69908
rect 7220 69868 7229 69908
rect 7363 69868 7372 69908
rect 7412 69868 7660 69908
rect 7756 69908 7796 70036
rect 16972 69992 17012 70036
rect 21388 69992 21428 70120
rect 21510 69992 21600 70012
rect 8105 69952 8140 69992
rect 8180 69952 8236 69992
rect 8276 69952 8285 69992
rect 8707 69952 8716 69992
rect 8756 69952 9196 69992
rect 9236 69952 9245 69992
rect 9562 69952 9571 69992
rect 9611 69952 9620 69992
rect 10339 69952 10348 69992
rect 10388 69952 10828 69992
rect 10868 69952 11212 69992
rect 11252 69952 11261 69992
rect 12067 69952 12076 69992
rect 12116 69952 12364 69992
rect 12404 69952 12652 69992
rect 12692 69952 12701 69992
rect 13996 69952 14572 69992
rect 14612 69952 14621 69992
rect 16156 69952 16300 69992
rect 16340 69952 16349 69992
rect 16963 69952 16972 69992
rect 17012 69952 17021 69992
rect 17155 69952 17164 69992
rect 17204 69952 17335 69992
rect 17923 69952 17932 69992
rect 17972 69952 18124 69992
rect 18164 69952 18316 69992
rect 18356 69952 18365 69992
rect 19625 69952 19756 69992
rect 19796 69952 19805 69992
rect 20009 69952 20140 69992
rect 20180 69952 20189 69992
rect 21388 69952 21600 69992
rect 9580 69908 9620 69952
rect 9772 69908 9812 69917
rect 13996 69908 14036 69952
rect 15724 69908 15764 69917
rect 7756 69868 8236 69908
rect 8276 69868 8285 69908
rect 8489 69868 8620 69908
rect 8660 69868 8669 69908
rect 8729 69868 8738 69908
rect 8778 69868 9620 69908
rect 9763 69868 9772 69908
rect 9812 69868 9943 69908
rect 10531 69868 10540 69908
rect 10580 69868 11020 69908
rect 11060 69868 11308 69908
rect 11348 69868 11357 69908
rect 12617 69868 12748 69908
rect 12788 69868 12797 69908
rect 14083 69868 14092 69908
rect 14132 69868 14476 69908
rect 14516 69868 14525 69908
rect 15764 69868 16012 69908
rect 16052 69868 16061 69908
rect 0 69656 90 69676
rect 0 69616 1324 69656
rect 1364 69616 1373 69656
rect 0 69596 90 69616
rect 0 69320 90 69340
rect 0 69280 460 69320
rect 500 69280 509 69320
rect 0 69260 90 69280
rect 1516 69236 1556 69868
rect 2764 69859 2804 69868
rect 3916 69859 3956 69868
rect 5164 69824 5204 69868
rect 6604 69859 6644 69868
rect 7660 69824 7700 69868
rect 9772 69859 9812 69868
rect 12748 69824 12788 69868
rect 13996 69824 14036 69868
rect 4003 69784 4012 69824
rect 4052 69784 4876 69824
rect 4916 69784 4925 69824
rect 5164 69784 6124 69824
rect 6164 69784 6173 69824
rect 7660 69784 8140 69824
rect 8180 69784 8189 69824
rect 12547 69784 12556 69824
rect 12596 69784 12788 69824
rect 12940 69784 14036 69824
rect 2947 69700 2956 69740
rect 2996 69700 3127 69740
rect 3283 69700 3292 69740
rect 3332 69700 3341 69740
rect 3715 69700 3724 69740
rect 3764 69700 4588 69740
rect 4628 69700 4637 69740
rect 5842 69700 6796 69740
rect 6836 69700 6845 69740
rect 6979 69700 6988 69740
rect 7028 69700 7180 69740
rect 7220 69700 7229 69740
rect 8227 69700 8236 69740
rect 8276 69700 8956 69740
rect 8996 69700 9005 69740
rect 11299 69700 11308 69740
rect 11348 69700 11452 69740
rect 11492 69700 11501 69740
rect 3292 69656 3332 69700
rect 2083 69616 2092 69656
rect 2132 69616 3332 69656
rect 4919 69532 4928 69572
rect 4968 69532 5010 69572
rect 5050 69532 5092 69572
rect 5132 69532 5174 69572
rect 5214 69532 5256 69572
rect 5296 69532 5305 69572
rect 5356 69532 5740 69572
rect 5780 69532 5789 69572
rect 5356 69488 5396 69532
rect 2860 69448 3956 69488
rect 2860 69404 2900 69448
rect 1699 69364 1708 69404
rect 1748 69364 2900 69404
rect 3916 69320 3956 69448
rect 4876 69448 5396 69488
rect 4876 69404 4916 69448
rect 5842 69404 5882 69700
rect 7363 69448 7372 69488
rect 7412 69448 7892 69488
rect 4867 69364 4876 69404
rect 4916 69364 4925 69404
rect 5842 69364 7371 69404
rect 7433 69364 7555 69404
rect 7604 69364 7613 69404
rect 5842 69320 5882 69364
rect 7331 69320 7371 69364
rect 7852 69320 7892 69448
rect 12940 69404 12980 69784
rect 14092 69740 14132 69868
rect 15724 69859 15764 69868
rect 13507 69700 13516 69740
rect 13556 69700 14132 69740
rect 14179 69700 14188 69740
rect 14228 69700 14237 69740
rect 15523 69700 15532 69740
rect 15572 69700 15916 69740
rect 15956 69700 15965 69740
rect 8035 69364 8044 69404
rect 8084 69364 12980 69404
rect 3916 69280 5020 69320
rect 5060 69280 5069 69320
rect 5644 69280 5882 69320
rect 5932 69280 6988 69320
rect 7028 69280 7037 69320
rect 7331 69280 7700 69320
rect 5644 69236 5684 69280
rect 5932 69236 5972 69280
rect 1411 69196 1420 69236
rect 1460 69196 1652 69236
rect 2633 69227 2764 69236
rect 2633 69196 2668 69227
rect 0 68984 90 69004
rect 0 68944 1228 68984
rect 1268 68944 1277 68984
rect 0 68924 90 68944
rect 0 68648 90 68668
rect 0 68608 76 68648
rect 116 68608 125 68648
rect 0 68588 90 68608
rect 1193 68356 1228 68396
rect 1268 68356 1324 68396
rect 1364 68356 1373 68396
rect 0 68312 90 68332
rect 0 68272 1036 68312
rect 1076 68272 1085 68312
rect 0 68252 90 68272
rect 1612 68228 1652 69196
rect 2708 69196 2764 69227
rect 2804 69196 2813 69236
rect 2987 69196 3052 69236
rect 3092 69196 3118 69236
rect 3158 69196 3167 69236
rect 3235 69196 3244 69236
rect 3284 69196 3380 69236
rect 3497 69196 3628 69236
rect 3668 69196 3677 69236
rect 4003 69196 4012 69236
rect 4052 69227 4244 69236
rect 4052 69196 4204 69227
rect 2668 69178 2708 69187
rect 2851 69112 2860 69152
rect 2900 69112 2909 69152
rect 2860 69068 2900 69112
rect 3340 69068 3380 69196
rect 4291 69196 4300 69236
rect 4340 69227 4724 69236
rect 4340 69196 4684 69227
rect 4204 69178 4244 69187
rect 5251 69196 5260 69236
rect 5300 69196 5452 69236
rect 5492 69196 5501 69236
rect 5626 69196 5635 69236
rect 5675 69196 5684 69236
rect 5731 69196 5740 69236
rect 5780 69196 5876 69236
rect 5923 69196 5932 69236
rect 5972 69196 5981 69236
rect 6883 69196 6892 69236
rect 6932 69227 7220 69236
rect 6932 69196 7180 69227
rect 4684 69178 4724 69187
rect 5836 69152 5876 69196
rect 7363 69196 7372 69236
rect 7412 69196 7555 69236
rect 7595 69196 7604 69236
rect 7660 69227 7700 69280
rect 7834 69311 7892 69320
rect 7834 69271 7843 69311
rect 7883 69271 7892 69311
rect 8227 69280 8236 69320
rect 8276 69280 8468 69320
rect 7834 69270 7892 69271
rect 8428 69236 8468 69280
rect 7180 69178 7220 69187
rect 7930 69196 7939 69236
rect 7979 69196 7988 69236
rect 8035 69196 8044 69236
rect 8113 69196 8215 69236
rect 8419 69196 8428 69236
rect 8468 69196 8477 69236
rect 9676 69227 9716 69364
rect 10675 69280 10684 69320
rect 10724 69280 11020 69320
rect 11060 69280 11069 69320
rect 14188 69236 14228 69700
rect 16156 69656 16196 69952
rect 21510 69932 21600 69952
rect 18700 69908 18740 69917
rect 17483 69868 17548 69908
rect 17588 69868 17614 69908
rect 17654 69868 17663 69908
rect 17731 69868 17740 69908
rect 17780 69868 17789 69908
rect 18211 69868 18220 69908
rect 18260 69868 18412 69908
rect 18452 69868 18548 69908
rect 18665 69868 18700 69908
rect 18740 69868 18796 69908
rect 18836 69868 18845 69908
rect 19145 69868 19219 69908
rect 19259 69868 19276 69908
rect 19316 69868 19325 69908
rect 21187 69868 21196 69908
rect 21236 69868 21332 69908
rect 17740 69824 17780 69868
rect 17740 69784 18124 69824
rect 18164 69784 18173 69824
rect 18508 69740 18548 69868
rect 18700 69859 18740 69868
rect 19987 69784 19996 69824
rect 20036 69784 21004 69824
rect 21044 69784 21053 69824
rect 18508 69700 18892 69740
rect 18932 69700 18941 69740
rect 19363 69700 19372 69740
rect 19412 69700 19421 69740
rect 19747 69700 19756 69740
rect 19796 69700 20044 69740
rect 20084 69700 20093 69740
rect 20371 69700 20380 69740
rect 20420 69700 21196 69740
rect 21236 69700 21245 69740
rect 19372 69656 19412 69700
rect 21292 69656 21332 69868
rect 16012 69616 16196 69656
rect 19075 69616 19084 69656
rect 19124 69616 19412 69656
rect 21100 69616 21332 69656
rect 14755 69448 14764 69488
rect 14804 69448 15052 69488
rect 15092 69448 15101 69488
rect 16012 69404 16052 69616
rect 20039 69532 20048 69572
rect 20088 69532 20130 69572
rect 20170 69532 20212 69572
rect 20252 69532 20294 69572
rect 20334 69532 20376 69572
rect 20416 69532 20425 69572
rect 21100 69488 21140 69616
rect 21510 69488 21600 69508
rect 17923 69448 17932 69488
rect 17972 69448 21140 69488
rect 21379 69448 21388 69488
rect 21428 69448 21600 69488
rect 20044 69404 20084 69448
rect 21510 69428 21600 69448
rect 16003 69364 16012 69404
rect 16052 69364 16061 69404
rect 17932 69364 19508 69404
rect 20035 69364 20044 69404
rect 20084 69364 20093 69404
rect 17932 69320 17972 69364
rect 19468 69320 19508 69364
rect 14673 69280 17972 69320
rect 18019 69280 18028 69320
rect 18068 69280 18356 69320
rect 18403 69280 18412 69320
rect 18452 69280 18548 69320
rect 18787 69280 18796 69320
rect 18836 69280 19412 69320
rect 19468 69280 20236 69320
rect 20276 69280 20285 69320
rect 7660 69178 7700 69187
rect 3715 69112 3724 69152
rect 3764 69112 4148 69152
rect 5251 69112 5260 69152
rect 5300 69112 5548 69152
rect 5588 69112 5597 69152
rect 5836 69112 7124 69152
rect 4108 69068 4148 69112
rect 7084 69068 7124 69112
rect 7948 69068 7988 69196
rect 11369 69196 11500 69236
rect 11540 69196 11549 69236
rect 11779 69196 11788 69236
rect 11828 69227 12788 69236
rect 11828 69196 12748 69227
rect 9676 69178 9716 69187
rect 12748 69178 12788 69187
rect 13036 69196 13940 69236
rect 14188 69196 14275 69236
rect 14315 69196 14324 69236
rect 14371 69196 14380 69236
rect 14420 69196 14572 69236
rect 14612 69196 14621 69236
rect 10121 69112 10252 69152
rect 10292 69112 10301 69152
rect 10409 69112 10444 69152
rect 10484 69112 10540 69152
rect 10580 69112 10589 69152
rect 13036 69068 13076 69196
rect 13193 69112 13324 69152
rect 13364 69112 13373 69152
rect 13673 69112 13804 69152
rect 13844 69112 13853 69152
rect 13900 69068 13940 69196
rect 14673 69152 14713 69280
rect 18316 69236 18356 69280
rect 18508 69236 18548 69280
rect 14851 69196 14860 69236
rect 14900 69196 15244 69236
rect 15284 69196 15293 69236
rect 15340 69227 15380 69236
rect 15523 69196 15532 69236
rect 15572 69227 15860 69236
rect 15572 69196 15820 69227
rect 14035 69112 14044 69152
rect 14084 69112 14713 69152
rect 14755 69112 14764 69152
rect 14804 69112 14935 69152
rect 2860 69028 3052 69068
rect 3092 69028 3101 69068
rect 3331 69028 3340 69068
rect 3380 69028 3389 69068
rect 4108 69028 6740 69068
rect 7084 69028 7276 69068
rect 7316 69028 7372 69068
rect 7412 69028 7988 69068
rect 8227 69028 8236 69068
rect 8276 69028 9772 69068
rect 9812 69028 10196 69068
rect 10339 69028 10348 69068
rect 10388 69028 13076 69068
rect 13219 69028 13228 69068
rect 13268 69028 13564 69068
rect 13604 69028 13613 69068
rect 13900 69028 14900 69068
rect 6700 68984 6740 69028
rect 10156 68984 10196 69028
rect 2851 68944 2860 68984
rect 2900 68944 3031 68984
rect 5731 68944 5740 68984
rect 5780 68944 5789 68984
rect 6691 68944 6700 68984
rect 6740 68944 7564 68984
rect 7604 68944 7613 68984
rect 9737 68944 9868 68984
rect 9908 68944 9917 68984
rect 10003 68944 10012 68984
rect 10052 68944 10100 68984
rect 10156 68944 12460 68984
rect 12500 68944 12509 68984
rect 12931 68944 12940 68984
rect 12980 68944 13460 68984
rect 5740 68816 5780 68944
rect 3679 68776 3688 68816
rect 3728 68776 3770 68816
rect 3810 68776 3852 68816
rect 3892 68776 3934 68816
rect 3974 68776 4016 68816
rect 4056 68776 4065 68816
rect 5740 68776 7372 68816
rect 7412 68776 7421 68816
rect 10060 68732 10100 68944
rect 13420 68900 13460 68944
rect 14860 68900 14900 69028
rect 15340 68984 15380 69187
rect 16579 69196 16588 69236
rect 16628 69196 16972 69236
rect 17012 69196 17021 69236
rect 17705 69196 17836 69236
rect 17876 69196 17885 69236
rect 18298 69196 18307 69236
rect 18347 69196 18356 69236
rect 18403 69196 18412 69236
rect 18452 69196 18461 69236
rect 18508 69196 18796 69236
rect 18836 69196 18845 69236
rect 19372 69227 19412 69280
rect 15820 69178 15860 69187
rect 17836 69178 17876 69187
rect 18412 69152 18452 69196
rect 19721 69196 19852 69236
rect 19892 69196 19901 69236
rect 19372 69178 19412 69187
rect 19852 69178 19892 69187
rect 16003 69112 16012 69152
rect 16052 69112 16156 69152
rect 16196 69112 16205 69152
rect 16387 69112 16396 69152
rect 16436 69112 16588 69152
rect 16628 69112 16637 69152
rect 18115 69112 18124 69152
rect 18164 69112 18452 69152
rect 18761 69112 18892 69152
rect 18932 69112 18941 69152
rect 18892 69068 18932 69112
rect 18403 69028 18412 69068
rect 18452 69028 18932 69068
rect 21510 68984 21600 69004
rect 14947 68944 14956 68984
rect 14996 68944 15380 68984
rect 20803 68944 20812 68984
rect 20852 68944 21600 68984
rect 21510 68924 21600 68944
rect 13420 68860 13804 68900
rect 13844 68860 13853 68900
rect 14860 68860 17548 68900
rect 17588 68860 17597 68900
rect 13132 68776 14572 68816
rect 14612 68776 14621 68816
rect 18799 68776 18808 68816
rect 18848 68776 18890 68816
rect 18930 68776 18972 68816
rect 19012 68776 19054 68816
rect 19094 68776 19136 68816
rect 19176 68776 19185 68816
rect 13132 68732 13172 68776
rect 1804 68692 2900 68732
rect 1804 68312 1844 68692
rect 2860 68648 2900 68692
rect 3340 68692 10100 68732
rect 10915 68692 10924 68732
rect 10964 68692 12460 68732
rect 12500 68692 13172 68732
rect 2179 68608 2188 68648
rect 2228 68608 2476 68648
rect 2516 68608 2525 68648
rect 2860 68608 3196 68648
rect 3236 68608 3245 68648
rect 1900 68524 2812 68564
rect 2852 68524 2861 68564
rect 1795 68272 1804 68312
rect 1844 68272 1853 68312
rect 1603 68188 1612 68228
rect 1652 68188 1661 68228
rect 1900 68060 1940 68524
rect 3340 68480 3380 68692
rect 4963 68608 4972 68648
rect 5012 68608 6220 68648
rect 6260 68608 8516 68648
rect 10003 68608 10012 68648
rect 10052 68608 10060 68648
rect 10100 68608 10212 68648
rect 13228 68608 15244 68648
rect 15284 68608 15293 68648
rect 16483 68608 16492 68648
rect 16532 68608 16828 68648
rect 16868 68608 16877 68648
rect 18979 68608 18988 68648
rect 19028 68608 19276 68648
rect 19316 68608 19325 68648
rect 3436 68524 7468 68564
rect 7508 68524 7517 68564
rect 3436 68480 3476 68524
rect 8476 68480 8516 68608
rect 8707 68524 8716 68564
rect 8756 68524 12652 68564
rect 12692 68524 12701 68564
rect 12748 68524 12940 68564
rect 12980 68524 12989 68564
rect 12748 68480 12788 68524
rect 13228 68480 13268 68608
rect 3043 68440 3052 68480
rect 3092 68440 3380 68480
rect 3427 68440 3436 68480
rect 3476 68440 3485 68480
rect 4003 68440 4012 68480
rect 4052 68440 4300 68480
rect 4340 68440 4349 68480
rect 6115 68440 6124 68480
rect 6164 68440 7124 68480
rect 7171 68440 7180 68480
rect 7220 68440 7372 68480
rect 7412 68440 7421 68480
rect 7555 68440 7564 68480
rect 7604 68440 8084 68480
rect 8201 68440 8236 68480
rect 8276 68440 8332 68480
rect 8372 68440 8381 68480
rect 8458 68440 8467 68480
rect 8507 68440 8516 68480
rect 9475 68440 9484 68480
rect 9524 68440 9772 68480
rect 9812 68440 9821 68480
rect 12739 68440 12748 68480
rect 12788 68440 12797 68480
rect 12844 68440 13268 68480
rect 13420 68524 19420 68564
rect 19460 68524 19469 68564
rect 20899 68524 20908 68564
rect 20948 68524 20957 68564
rect 2476 68396 2516 68405
rect 4876 68396 4916 68405
rect 5932 68396 5972 68405
rect 7084 68396 7124 68440
rect 8044 68396 8084 68440
rect 8908 68396 8948 68405
rect 11692 68396 11732 68405
rect 12844 68396 12884 68440
rect 13324 68396 13364 68405
rect 1987 68356 1996 68396
rect 2036 68356 2476 68396
rect 2516 68356 2804 68396
rect 2947 68356 2956 68396
rect 2996 68356 3811 68396
rect 3851 68356 3860 68396
rect 3907 68356 3916 68396
rect 3956 68356 4087 68396
rect 4204 68356 4396 68396
rect 4436 68356 4445 68396
rect 5386 68356 5395 68396
rect 5435 68356 5780 68396
rect 5923 68356 5932 68396
rect 5972 68356 6103 68396
rect 7084 68356 7180 68396
rect 7220 68356 7229 68396
rect 7363 68356 7372 68396
rect 7412 68356 7843 68396
rect 7883 68356 7892 68396
rect 7939 68356 7948 68396
rect 7988 68356 7997 68396
rect 8044 68356 8908 68396
rect 9418 68356 9427 68396
rect 9467 68356 9868 68396
rect 9908 68356 9917 68396
rect 10435 68356 10444 68396
rect 10484 68356 10493 68396
rect 11657 68356 11692 68396
rect 11732 68356 11788 68396
rect 11828 68356 11837 68396
rect 12250 68356 12259 68396
rect 12299 68356 12308 68396
rect 12355 68356 12364 68396
rect 12404 68356 12460 68396
rect 12500 68356 12535 68396
rect 12835 68356 12844 68396
rect 12884 68356 12893 68396
rect 13193 68356 13228 68396
rect 13268 68356 13324 68396
rect 2476 68347 2516 68356
rect 2537 68188 2572 68228
rect 2612 68188 2668 68228
rect 2708 68188 2717 68228
rect 2764 68144 2804 68356
rect 4204 68228 4244 68356
rect 4876 68312 4916 68356
rect 5740 68312 5780 68356
rect 5932 68347 5972 68356
rect 4291 68272 4300 68312
rect 4340 68272 4916 68312
rect 5731 68272 5740 68312
rect 5780 68272 5789 68312
rect 7180 68228 7220 68356
rect 7948 68312 7988 68356
rect 8908 68347 8948 68356
rect 7459 68272 7468 68312
rect 7508 68272 7988 68312
rect 9580 68272 10252 68312
rect 10292 68272 10301 68312
rect 9580 68228 9620 68272
rect 10444 68228 10484 68356
rect 11692 68347 11732 68356
rect 12268 68312 12308 68356
rect 13324 68347 13364 68356
rect 11875 68272 11884 68312
rect 11924 68272 12308 68312
rect 12931 68272 12940 68312
rect 12980 68272 12989 68312
rect 12940 68228 12980 68272
rect 4204 68188 4972 68228
rect 5012 68188 5021 68228
rect 5417 68188 5548 68228
rect 5588 68188 5597 68228
rect 7171 68188 7180 68228
rect 7220 68188 7229 68228
rect 7603 68188 7612 68228
rect 7652 68188 8236 68228
rect 8276 68188 8285 68228
rect 9571 68188 9580 68228
rect 9620 68188 9629 68228
rect 10444 68188 12980 68228
rect 13420 68144 13460 68524
rect 20908 68480 20948 68524
rect 21510 68480 21600 68500
rect 14026 68440 14035 68480
rect 14075 68440 14380 68480
rect 14420 68440 14429 68480
rect 15331 68440 15340 68480
rect 15380 68440 15532 68480
rect 15572 68440 15581 68480
rect 16108 68440 17068 68480
rect 17108 68440 17117 68480
rect 19651 68440 19660 68480
rect 19700 68440 19852 68480
rect 19892 68440 19901 68480
rect 20131 68440 20140 68480
rect 20180 68440 20189 68480
rect 20908 68440 21600 68480
rect 15916 68396 15956 68405
rect 16108 68396 16148 68440
rect 18796 68396 18836 68405
rect 13795 68356 13804 68396
rect 13852 68356 13975 68396
rect 14371 68356 14380 68396
rect 14420 68356 14851 68396
rect 14891 68356 14900 68396
rect 14947 68356 14956 68396
rect 14996 68356 15005 68396
rect 15427 68356 15436 68396
rect 15476 68356 15820 68396
rect 15860 68356 15869 68396
rect 15956 68356 16148 68396
rect 16195 68356 16204 68396
rect 16244 68356 16404 68396
rect 16444 68356 16453 68396
rect 17417 68356 17548 68396
rect 17588 68356 17597 68396
rect 18665 68356 18796 68396
rect 18836 68356 18845 68396
rect 14956 68312 14996 68356
rect 15916 68347 15956 68356
rect 16108 68312 16148 68356
rect 18796 68347 18836 68356
rect 13987 68272 13996 68312
rect 14036 68272 14516 68312
rect 14563 68272 14572 68312
rect 14612 68272 14996 68312
rect 16099 68272 16108 68312
rect 16148 68272 16157 68312
rect 2764 68104 4204 68144
rect 4244 68104 10060 68144
rect 10100 68104 10109 68144
rect 10243 68104 10252 68144
rect 10292 68104 13460 68144
rect 13516 68188 14140 68228
rect 14180 68188 14189 68228
rect 13516 68060 13556 68188
rect 14476 68144 14516 68272
rect 20140 68228 20180 68440
rect 21510 68420 21600 68440
rect 16457 68188 16588 68228
rect 16628 68188 16637 68228
rect 17251 68188 17260 68228
rect 17300 68188 20180 68228
rect 20227 68188 20236 68228
rect 20276 68188 20285 68228
rect 20371 68188 20380 68228
rect 20420 68188 21388 68228
rect 21428 68188 21437 68228
rect 20236 68144 20276 68188
rect 14476 68104 14860 68144
rect 14900 68104 16492 68144
rect 16532 68104 17972 68144
rect 20236 68104 20948 68144
rect 1315 68020 1324 68060
rect 1364 68020 1940 68060
rect 4919 68020 4928 68060
rect 4968 68020 5010 68060
rect 5050 68020 5092 68060
rect 5132 68020 5174 68060
rect 5214 68020 5256 68060
rect 5296 68020 5305 68060
rect 7555 68020 7564 68060
rect 7604 68020 13556 68060
rect 13987 68020 13996 68060
rect 14036 68020 17780 68060
rect 0 67976 90 67996
rect 0 67936 844 67976
rect 884 67936 893 67976
rect 7075 67936 7084 67976
rect 7124 67936 9620 67976
rect 10627 67936 10636 67976
rect 10676 67936 11116 67976
rect 11156 67936 11165 67976
rect 11875 67936 11884 67976
rect 11924 67936 12980 67976
rect 0 67916 90 67936
rect 9580 67808 9620 67936
rect 10531 67852 10540 67892
rect 10580 67852 12748 67892
rect 12788 67852 12797 67892
rect 12940 67808 12980 67936
rect 13027 67852 13036 67892
rect 13076 67852 15532 67892
rect 15572 67852 15581 67892
rect 16073 67852 16204 67892
rect 16244 67852 16253 67892
rect 3148 67768 3916 67808
rect 3956 67768 3965 67808
rect 4108 67768 5396 67808
rect 7171 67768 7180 67808
rect 7220 67768 9484 67808
rect 9524 67768 9533 67808
rect 9580 67768 10676 67808
rect 3148 67724 3188 67768
rect 4108 67724 4148 67768
rect 5356 67724 5396 67768
rect 835 67684 844 67724
rect 884 67684 1324 67724
rect 1364 67684 2476 67724
rect 2516 67684 2525 67724
rect 2572 67715 2668 67724
rect 2612 67684 2668 67715
rect 2708 67684 2743 67724
rect 2851 67684 2860 67724
rect 2900 67684 3043 67724
rect 3083 67684 3092 67724
rect 3139 67684 3148 67724
rect 3188 67684 3197 67724
rect 3523 67684 3532 67724
rect 3572 67684 3581 67724
rect 3977 67684 4108 67724
rect 4148 67684 4157 67724
rect 4457 67684 4588 67724
rect 4628 67684 4637 67724
rect 5347 67684 5356 67724
rect 5396 67684 5405 67724
rect 5609 67684 5644 67724
rect 5684 67684 5740 67724
rect 5780 67684 5789 67724
rect 6761 67684 6892 67724
rect 6932 67684 7316 67724
rect 7363 67684 7372 67724
rect 7412 67684 8236 67724
rect 8276 67684 8428 67724
rect 8468 67684 8477 67724
rect 8524 67715 9292 67724
rect 8524 67684 8620 67715
rect 2572 67666 2612 67675
rect 0 67640 90 67660
rect 3532 67640 3572 67684
rect 4108 67666 4148 67675
rect 4588 67666 4628 67675
rect 6892 67666 6932 67675
rect 7276 67640 7316 67684
rect 8524 67640 8564 67684
rect 8660 67684 9292 67715
rect 9332 67684 9341 67724
rect 9475 67684 9484 67724
rect 9524 67684 10348 67724
rect 10388 67684 10397 67724
rect 8620 67666 8660 67675
rect 0 67600 1420 67640
rect 1460 67600 1469 67640
rect 3331 67600 3340 67640
rect 3380 67600 3572 67640
rect 3619 67600 3628 67640
rect 3668 67600 3677 67640
rect 4771 67600 4780 67640
rect 4820 67600 5164 67640
rect 5204 67600 5213 67640
rect 7276 67600 8564 67640
rect 8873 67600 9004 67640
rect 9044 67600 9053 67640
rect 9235 67600 9244 67640
rect 9284 67600 9676 67640
rect 9716 67600 9725 67640
rect 0 67580 90 67600
rect 3628 67556 3668 67600
rect 10636 67556 10676 67768
rect 10732 67768 12884 67808
rect 12940 67768 14420 67808
rect 15427 67768 15436 67808
rect 15476 67768 16628 67808
rect 10732 67715 10772 67768
rect 10985 67684 11116 67724
rect 11156 67684 11165 67724
rect 11212 67684 12172 67724
rect 12212 67684 12221 67724
rect 12364 67715 12404 67768
rect 12844 67724 12884 67768
rect 14380 67724 14420 67768
rect 16588 67724 16628 67768
rect 17740 67724 17780 68020
rect 17932 67808 17972 68104
rect 20039 68020 20048 68060
rect 20088 68020 20130 68060
rect 20170 68020 20212 68060
rect 20252 68020 20294 68060
rect 20334 68020 20376 68060
rect 20416 68020 20425 68060
rect 20908 67976 20948 68104
rect 21510 67976 21600 67996
rect 20908 67936 21600 67976
rect 21510 67916 21600 67936
rect 17932 67768 18644 67808
rect 18604 67724 18644 67768
rect 10732 67666 10772 67675
rect 11212 67556 11252 67684
rect 12617 67684 12748 67724
rect 12788 67684 12797 67724
rect 12844 67684 13940 67724
rect 12364 67666 12404 67675
rect 3628 67516 4300 67556
rect 4340 67516 4349 67556
rect 4819 67516 4828 67556
rect 4868 67516 4876 67556
rect 4916 67516 4999 67556
rect 5491 67516 5500 67556
rect 5540 67516 8044 67556
rect 8084 67516 8093 67556
rect 10636 67516 11252 67556
rect 13900 67556 13940 67684
rect 13996 67715 14092 67724
rect 14036 67684 14092 67715
rect 14132 67684 14167 67724
rect 14380 67684 14764 67724
rect 14804 67684 15244 67724
rect 15284 67684 15293 67724
rect 16012 67715 16052 67724
rect 13996 67666 14036 67675
rect 14380 67640 14420 67684
rect 16579 67684 16588 67724
rect 16628 67684 16972 67724
rect 17012 67684 17021 67724
rect 17740 67715 18548 67724
rect 17740 67684 18220 67715
rect 16012 67640 16052 67675
rect 18260 67684 18548 67715
rect 18595 67684 18604 67724
rect 18644 67684 18653 67724
rect 18700 67715 20140 67724
rect 18700 67684 19852 67715
rect 18220 67666 18260 67675
rect 18508 67640 18548 67684
rect 18700 67640 18740 67684
rect 19892 67684 20140 67715
rect 20180 67684 20189 67724
rect 19852 67666 19892 67675
rect 14371 67600 14380 67640
rect 14420 67600 14429 67640
rect 14851 67600 14860 67640
rect 14900 67600 16052 67640
rect 16483 67600 16492 67640
rect 16532 67600 16588 67640
rect 16628 67600 16663 67640
rect 16819 67600 16828 67640
rect 16868 67600 17260 67640
rect 17300 67600 17309 67640
rect 18508 67600 18740 67640
rect 13900 67516 13996 67556
rect 14036 67516 14045 67556
rect 14179 67516 14188 67556
rect 14228 67516 14380 67556
rect 14420 67516 14429 67556
rect 15811 67516 15820 67556
rect 15860 67516 18796 67556
rect 18836 67516 18845 67556
rect 21510 67472 21600 67492
rect 2467 67432 2476 67472
rect 2516 67432 2764 67472
rect 2804 67432 2813 67472
rect 2860 67432 4924 67472
rect 4964 67432 4973 67472
rect 7075 67432 7084 67472
rect 7124 67432 7133 67472
rect 8803 67432 8812 67472
rect 8852 67432 8861 67472
rect 10915 67432 10924 67472
rect 10964 67432 10973 67472
rect 12547 67432 12556 67472
rect 12596 67432 12605 67472
rect 14537 67432 14620 67472
rect 14660 67432 14668 67472
rect 14708 67432 15436 67472
rect 15476 67432 15485 67472
rect 18403 67432 18412 67472
rect 18452 67432 18461 67472
rect 20035 67432 20044 67472
rect 20084 67432 20093 67472
rect 21283 67432 21292 67472
rect 21332 67432 21600 67472
rect 0 67304 90 67324
rect 2860 67304 2900 67432
rect 0 67264 652 67304
rect 692 67264 701 67304
rect 2083 67264 2092 67304
rect 2132 67264 2900 67304
rect 3679 67264 3688 67304
rect 3728 67264 3770 67304
rect 3810 67264 3852 67304
rect 3892 67264 3934 67304
rect 3974 67264 4016 67304
rect 4056 67264 4065 67304
rect 0 67244 90 67264
rect 172 67096 5836 67136
rect 5876 67096 5885 67136
rect 0 66968 90 66988
rect 172 66968 212 67096
rect 4387 67012 4396 67052
rect 4436 67012 4972 67052
rect 5012 67012 5212 67052
rect 5252 67012 5261 67052
rect 0 66928 212 66968
rect 1289 66928 1420 66968
rect 1460 66928 1469 66968
rect 4099 66928 4108 66968
rect 4148 66928 4972 66968
rect 5012 66928 5021 66968
rect 0 66908 90 66928
rect 2956 66884 2996 66893
rect 3532 66884 3572 66893
rect 6604 66884 6644 66893
rect 7084 66884 7124 67432
rect 7372 67012 8620 67052
rect 8660 67012 8669 67052
rect 7372 66884 7412 67012
rect 7529 66928 7564 66968
rect 7604 66928 7660 66968
rect 7700 66928 7709 66968
rect 8140 66884 8180 66893
rect 8812 66884 8852 67432
rect 8899 67096 8908 67136
rect 8948 67096 8956 67136
rect 8996 67096 9079 67136
rect 9187 66928 9196 66968
rect 9236 66928 9245 66968
rect 1699 66844 1708 66884
rect 1748 66844 1996 66884
rect 2036 66844 2045 66884
rect 2825 66844 2956 66884
rect 2996 66844 3005 66884
rect 3572 66844 4204 66884
rect 4244 66844 4253 66884
rect 4745 66844 4780 66884
rect 4820 66844 4876 66884
rect 4916 66844 4925 66884
rect 5347 66844 5356 66884
rect 5396 66844 5836 66884
rect 5876 66844 5885 66884
rect 6211 66844 6220 66884
rect 6260 66844 6604 66884
rect 7066 66844 7075 66884
rect 7115 66844 7124 66884
rect 7171 66844 7180 66884
rect 7220 66844 7412 66884
rect 7564 66844 7660 66884
rect 7700 66844 7709 66884
rect 8009 66844 8140 66884
rect 8180 66844 8189 66884
rect 8650 66844 8659 66884
rect 8699 66844 8852 66884
rect 2956 66835 2996 66844
rect 3532 66835 3572 66844
rect 6604 66835 6644 66844
rect 6787 66760 6796 66800
rect 6836 66760 7372 66800
rect 7412 66760 7421 66800
rect 7564 66716 7604 66844
rect 8140 66800 8180 66844
rect 9196 66800 9236 66928
rect 10732 66884 10772 66893
rect 9353 66844 9484 66884
rect 9524 66844 9533 66884
rect 10147 66844 10156 66884
rect 10196 66844 10732 66884
rect 10924 66884 10964 67432
rect 11491 66928 11500 66968
rect 11540 66928 11692 66968
rect 11732 66928 11741 66968
rect 12268 66884 12308 66893
rect 10924 66844 11203 66884
rect 11243 66844 11252 66884
rect 11299 66844 11308 66884
rect 11348 66844 11404 66884
rect 11444 66844 11479 66884
rect 11683 66844 11692 66884
rect 11732 66844 11788 66884
rect 11828 66844 11863 66884
rect 12556 66884 12596 67432
rect 13123 67096 13132 67136
rect 13172 67096 13372 67136
rect 13412 67096 13421 67136
rect 15475 67096 15484 67136
rect 15524 67096 18028 67136
rect 18068 67096 18077 67136
rect 12835 67012 12844 67052
rect 12884 67012 15668 67052
rect 15859 67012 15868 67052
rect 15908 67012 17164 67052
rect 17204 67012 17213 67052
rect 15628 66968 15668 67012
rect 18412 66968 18452 67432
rect 18799 67264 18808 67304
rect 18848 67264 18890 67304
rect 18930 67264 18972 67304
rect 19012 67264 19054 67304
rect 19094 67264 19136 67304
rect 19176 67264 19185 67304
rect 13123 66928 13132 66968
rect 13172 66928 13996 66968
rect 14036 66928 14045 66968
rect 15113 66928 15244 66968
rect 15284 66928 15293 66968
rect 15619 66928 15628 66968
rect 15668 66928 15677 66968
rect 15811 66928 15820 66968
rect 15860 66928 16012 66968
rect 16052 66928 16061 66968
rect 18124 66928 18452 66968
rect 18595 66928 18604 66968
rect 18644 66928 18653 66968
rect 14860 66884 14900 66893
rect 17644 66884 17684 66893
rect 18124 66884 18164 66928
rect 18604 66884 18644 66928
rect 19180 66884 19220 66893
rect 20044 66884 20084 67432
rect 21510 67412 21600 67432
rect 20803 67012 20812 67052
rect 20852 67012 20861 67052
rect 20812 66968 20852 67012
rect 21510 66968 21600 66988
rect 20227 66928 20236 66968
rect 20276 66928 20716 66968
rect 20756 66928 20765 66968
rect 20812 66928 21600 66968
rect 21510 66908 21600 66928
rect 12556 66844 12756 66884
rect 12796 66844 12805 66884
rect 13507 66844 13516 66884
rect 13556 66844 13612 66884
rect 13652 66844 13687 66884
rect 14083 66844 14092 66884
rect 14132 66844 14860 66884
rect 14900 66844 14909 66884
rect 16291 66844 16300 66884
rect 16340 66844 16396 66884
rect 16436 66844 16588 66884
rect 16628 66844 16637 66884
rect 17609 66844 17644 66884
rect 17684 66844 17740 66884
rect 17780 66844 17789 66884
rect 18106 66844 18115 66884
rect 18155 66844 18164 66884
rect 18211 66844 18220 66884
rect 18260 66844 18269 66884
rect 18403 66844 18412 66884
rect 18452 66844 18644 66884
rect 18691 66844 18700 66884
rect 18740 66844 18796 66884
rect 18836 66844 18871 66884
rect 19690 66844 19699 66884
rect 19739 66844 20084 66884
rect 10732 66835 10772 66844
rect 7651 66760 7660 66800
rect 7700 66760 8180 66800
rect 8812 66760 9236 66800
rect 12268 66800 12308 66844
rect 14860 66835 14900 66844
rect 17644 66835 17684 66844
rect 18220 66800 18260 66844
rect 19180 66800 19220 66844
rect 12268 66760 12748 66800
rect 12788 66760 12797 66800
rect 18115 66760 18124 66800
rect 18164 66760 18260 66800
rect 18307 66760 18316 66800
rect 18356 66760 19220 66800
rect 8812 66716 8852 66760
rect 643 66676 652 66716
rect 692 66676 1180 66716
rect 1220 66676 1229 66716
rect 2659 66676 2668 66716
rect 2708 66676 3148 66716
rect 3188 66676 3197 66716
rect 3331 66676 3340 66716
rect 3380 66676 4204 66716
rect 4244 66676 4253 66716
rect 7564 66676 8332 66716
rect 8372 66676 8381 66716
rect 8803 66676 8812 66716
rect 8852 66676 8861 66716
rect 10915 66676 10924 66716
rect 10964 66676 11116 66716
rect 11156 66676 11165 66716
rect 12876 66676 12940 66716
rect 12980 66676 13036 66716
rect 13076 66676 13111 66716
rect 14921 66676 15052 66716
rect 15092 66676 15101 66716
rect 16099 66676 16108 66716
rect 16148 66676 16252 66716
rect 16292 66676 17356 66716
rect 17396 66676 17405 66716
rect 17705 66676 17836 66716
rect 17876 66676 17885 66716
rect 19721 66676 19756 66716
rect 19796 66676 19852 66716
rect 19892 66676 19901 66716
rect 19948 66676 19996 66716
rect 20036 66676 20045 66716
rect 20419 66676 20428 66716
rect 20468 66676 20660 66716
rect 0 66632 90 66652
rect 19948 66632 19988 66676
rect 0 66592 940 66632
rect 980 66592 989 66632
rect 11875 66592 11884 66632
rect 11924 66592 13516 66632
rect 13556 66592 13565 66632
rect 16483 66592 16492 66632
rect 16532 66592 19988 66632
rect 0 66572 90 66592
rect 4919 66508 4928 66548
rect 4968 66508 5010 66548
rect 5050 66508 5092 66548
rect 5132 66508 5174 66548
rect 5214 66508 5256 66548
rect 5296 66508 5305 66548
rect 6403 66508 6412 66548
rect 6452 66508 7604 66548
rect 20039 66508 20048 66548
rect 20088 66508 20130 66548
rect 20170 66508 20212 66548
rect 20252 66508 20294 66548
rect 20334 66508 20376 66548
rect 20416 66508 20425 66548
rect 4387 66340 4396 66380
rect 4436 66340 4780 66380
rect 4820 66340 4829 66380
rect 5932 66340 6988 66380
rect 7028 66340 7276 66380
rect 7316 66340 7325 66380
rect 0 66296 90 66316
rect 0 66256 1228 66296
rect 1268 66256 1277 66296
rect 2729 66256 2860 66296
rect 2900 66256 4492 66296
rect 4532 66256 5356 66296
rect 5396 66256 5405 66296
rect 0 66236 90 66256
rect 2764 66212 2804 66256
rect 5932 66212 5972 66340
rect 6220 66256 6844 66296
rect 6884 66256 6893 66296
rect 6220 66212 6260 66256
rect 1411 66172 1420 66212
rect 1460 66172 1612 66212
rect 1652 66172 1661 66212
rect 2507 66172 2572 66212
rect 2612 66172 2638 66212
rect 2678 66172 2687 66212
rect 2755 66172 2764 66212
rect 2804 66172 2813 66212
rect 3139 66172 3148 66212
rect 3188 66172 3628 66212
rect 3668 66172 3677 66212
rect 3724 66203 3820 66212
rect 3764 66172 3820 66203
rect 3860 66172 3895 66212
rect 4073 66172 4204 66212
rect 4244 66172 4253 66212
rect 4771 66172 4780 66212
rect 4820 66172 5972 66212
rect 6028 66203 6220 66212
rect 3724 66154 3764 66163
rect 4204 66154 4244 66163
rect 6068 66172 6220 66203
rect 6260 66172 6269 66212
rect 6028 66154 6068 66163
rect 7564 66128 7604 66508
rect 20620 66464 20660 66676
rect 21510 66464 21600 66484
rect 20620 66424 21600 66464
rect 21510 66404 21600 66424
rect 13795 66340 13804 66380
rect 13844 66340 17116 66380
rect 17156 66340 17165 66380
rect 20323 66340 20332 66380
rect 20372 66340 21292 66380
rect 21332 66340 21341 66380
rect 12643 66256 12652 66296
rect 12692 66256 14324 66296
rect 14659 66256 14668 66296
rect 14708 66256 14996 66296
rect 14284 66212 14324 66256
rect 14956 66212 14996 66256
rect 15820 66256 16732 66296
rect 16772 66256 16781 66296
rect 18019 66256 18028 66296
rect 18068 66256 18740 66296
rect 15820 66212 15860 66256
rect 18700 66212 18740 66256
rect 7817 66172 7948 66212
rect 7988 66172 7997 66212
rect 9196 66203 9236 66212
rect 9475 66172 9484 66212
rect 9524 66172 9868 66212
rect 9908 66172 9917 66212
rect 11116 66203 11788 66212
rect 9196 66128 9236 66163
rect 11156 66172 11788 66203
rect 11828 66172 11837 66212
rect 12067 66172 12076 66212
rect 12116 66172 12460 66212
rect 12500 66172 13036 66212
rect 13076 66172 13085 66212
rect 14249 66203 14380 66212
rect 14249 66172 14284 66203
rect 11116 66128 11156 66163
rect 14324 66172 14380 66203
rect 14420 66172 14429 66212
rect 14476 66172 14851 66212
rect 14891 66172 14900 66212
rect 14947 66172 14956 66212
rect 14996 66172 15005 66212
rect 15209 66172 15340 66212
rect 15380 66172 15389 66212
rect 15619 66172 15628 66212
rect 15668 66172 15860 66212
rect 15916 66203 15956 66212
rect 14284 66154 14324 66163
rect 1411 66088 1420 66128
rect 1460 66088 1469 66128
rect 1673 66088 1804 66128
rect 1844 66088 1853 66128
rect 1987 66088 1996 66128
rect 2036 66088 2045 66128
rect 2179 66088 2188 66128
rect 2228 66088 2237 66128
rect 3235 66088 3244 66128
rect 3284 66088 3293 66128
rect 6595 66088 6604 66128
rect 6683 66088 6775 66128
rect 6883 66088 6892 66128
rect 6932 66088 6988 66128
rect 7028 66088 7063 66128
rect 7555 66088 7564 66128
rect 7604 66088 7613 66128
rect 9196 66088 11156 66128
rect 11203 66088 11212 66128
rect 11252 66088 11540 66128
rect 12835 66088 12844 66128
rect 12884 66088 13036 66128
rect 13076 66088 13085 66128
rect 13219 66088 13228 66128
rect 13268 66088 13516 66128
rect 13556 66088 13565 66128
rect 1420 66044 1460 66088
rect 1996 66044 2036 66088
rect 1420 66004 2036 66044
rect 0 65960 90 65980
rect 2188 65960 2228 66088
rect 3244 66044 3284 66088
rect 11500 66044 11540 66088
rect 14476 66044 14516 66172
rect 16265 66172 16396 66212
rect 16436 66172 16445 66212
rect 17827 66172 17836 66212
rect 17876 66172 18211 66212
rect 18251 66172 18260 66212
rect 18307 66172 18316 66212
rect 18356 66172 18487 66212
rect 18691 66172 18700 66212
rect 18740 66172 18749 66212
rect 19145 66172 19276 66212
rect 19316 66172 19325 66212
rect 19756 66203 20180 66212
rect 14755 66088 14764 66128
rect 14804 66088 15436 66128
rect 15476 66088 15724 66128
rect 15764 66088 15773 66128
rect 15916 66044 15956 66163
rect 16396 66154 16436 66163
rect 19276 66154 19316 66163
rect 19796 66172 20180 66203
rect 19756 66154 19796 66163
rect 16618 66088 16627 66128
rect 16667 66088 16972 66128
rect 17012 66088 17021 66128
rect 17347 66088 17356 66128
rect 17396 66088 17405 66128
rect 17609 66088 17740 66128
rect 17780 66088 17789 66128
rect 18787 66088 18796 66128
rect 18836 66088 19180 66128
rect 19220 66088 19229 66128
rect 2851 66004 2860 66044
rect 2900 66004 3284 66044
rect 7171 66004 7180 66044
rect 7220 66004 7228 66044
rect 7268 66004 7351 66044
rect 11500 66004 14420 66044
rect 14467 66004 14476 66044
rect 14516 66004 14525 66044
rect 15756 66004 15820 66044
rect 15860 66004 16780 66044
rect 16820 66004 16829 66044
rect 14380 65960 14420 66004
rect 0 65920 460 65960
rect 500 65920 509 65960
rect 931 65920 940 65960
rect 980 65920 1180 65960
rect 1220 65920 1229 65960
rect 1555 65920 1564 65960
rect 1604 65920 1612 65960
rect 1652 65920 1735 65960
rect 1939 65920 1948 65960
rect 1988 65920 1996 65960
rect 2036 65920 2119 65960
rect 2188 65920 5356 65960
rect 5396 65920 5405 65960
rect 5827 65920 5836 65960
rect 5876 65920 6220 65960
rect 6260 65920 6269 65960
rect 7315 65920 7324 65960
rect 7364 65920 7373 65960
rect 9379 65920 9388 65960
rect 9428 65920 9484 65960
rect 9524 65920 9559 65960
rect 9955 65920 9964 65960
rect 10004 65920 10636 65960
rect 10676 65920 10685 65960
rect 11011 65920 11020 65960
rect 11060 65920 11308 65960
rect 11348 65920 11357 65960
rect 11491 65920 11500 65960
rect 11540 65920 12604 65960
rect 12644 65920 12653 65960
rect 14380 65920 16492 65960
rect 16532 65920 16541 65960
rect 0 65900 90 65920
rect 7324 65876 7364 65920
rect 1219 65836 1228 65876
rect 1268 65836 7364 65876
rect 7468 65836 11212 65876
rect 11252 65836 11261 65876
rect 13132 65836 13804 65876
rect 13844 65836 13853 65876
rect 7468 65792 7508 65836
rect 13132 65792 13172 65836
rect 3244 65752 3476 65792
rect 3679 65752 3688 65792
rect 3728 65752 3770 65792
rect 3810 65752 3852 65792
rect 3892 65752 3934 65792
rect 3974 65752 4016 65792
rect 4056 65752 4065 65792
rect 5347 65752 5356 65792
rect 5396 65752 7508 65792
rect 7852 65752 13172 65792
rect 3244 65708 3284 65752
rect 1795 65668 1804 65708
rect 1844 65668 3284 65708
rect 3436 65708 3476 65752
rect 7852 65708 7892 65752
rect 3436 65668 7892 65708
rect 8803 65668 8812 65708
rect 8852 65668 9716 65708
rect 0 65624 90 65644
rect 0 65584 268 65624
rect 308 65584 317 65624
rect 1411 65584 1420 65624
rect 1460 65584 2900 65624
rect 2947 65584 2956 65624
rect 2996 65584 3100 65624
rect 3140 65584 3149 65624
rect 4003 65584 4012 65624
rect 4052 65584 5932 65624
rect 5972 65584 6220 65624
rect 6260 65584 6269 65624
rect 0 65564 90 65584
rect 2860 65540 2900 65584
rect 2860 65500 7948 65540
rect 7988 65500 7997 65540
rect 9283 65500 9292 65540
rect 9332 65500 9620 65540
rect 2851 65416 2860 65456
rect 2900 65416 3340 65456
rect 3380 65416 3389 65456
rect 3523 65416 3532 65456
rect 3572 65416 3724 65456
rect 3764 65416 3773 65456
rect 4169 65416 4300 65456
rect 4340 65416 4349 65456
rect 4396 65416 5684 65456
rect 3340 65372 3380 65416
rect 4396 65372 4436 65416
rect 1385 65332 1420 65372
rect 1460 65332 1516 65372
rect 1556 65332 1565 65372
rect 2763 65332 2772 65372
rect 2812 65332 2956 65372
rect 2996 65332 3005 65372
rect 3340 65332 4436 65372
rect 4483 65332 4492 65372
rect 4532 65332 5164 65372
rect 5204 65332 5213 65372
rect 0 65288 90 65308
rect 0 65248 364 65288
rect 404 65248 413 65288
rect 1027 65248 1036 65288
rect 1076 65248 3484 65288
rect 3524 65248 3533 65288
rect 0 65228 90 65248
rect 2947 65164 2956 65204
rect 2996 65164 3127 65204
rect 3523 65164 3532 65204
rect 3572 65164 4060 65204
rect 4100 65164 4109 65204
rect 4492 65120 4532 65332
rect 4003 65080 4012 65120
rect 4052 65080 4532 65120
rect 5644 65036 5684 65416
rect 5740 65372 5780 65381
rect 6124 65372 6164 65500
rect 7372 65372 7412 65381
rect 7756 65372 7796 65500
rect 9437 65416 9484 65456
rect 9524 65416 9533 65456
rect 9004 65372 9044 65381
rect 9484 65372 9524 65416
rect 9580 65372 9620 65500
rect 9676 65372 9716 65668
rect 17356 65624 17396 66088
rect 18595 66004 18604 66044
rect 18644 66004 19996 66044
rect 20036 66004 20045 66044
rect 17971 65920 17980 65960
rect 18020 65920 20044 65960
rect 20084 65920 20093 65960
rect 18799 65752 18808 65792
rect 18848 65752 18890 65792
rect 18930 65752 18972 65792
rect 19012 65752 19054 65792
rect 19094 65752 19136 65792
rect 19176 65752 19185 65792
rect 20140 65624 20180 66172
rect 21510 65960 21600 65980
rect 21475 65920 21484 65960
rect 21524 65920 21600 65960
rect 21510 65900 21600 65920
rect 12019 65584 12028 65624
rect 12068 65584 12652 65624
rect 12692 65584 12701 65624
rect 13228 65584 15340 65624
rect 15380 65584 15389 65624
rect 16906 65584 16915 65624
rect 16955 65584 17396 65624
rect 20131 65584 20140 65624
rect 20180 65584 20189 65624
rect 9955 65416 9964 65456
rect 10004 65416 10292 65456
rect 11683 65416 11692 65456
rect 11732 65416 11788 65456
rect 11828 65416 12124 65456
rect 12164 65416 12173 65456
rect 12355 65416 12364 65456
rect 12404 65416 12844 65456
rect 12884 65416 12893 65456
rect 13001 65416 13132 65456
rect 13172 65416 13181 65456
rect 10252 65372 10292 65416
rect 10540 65372 10580 65381
rect 13228 65372 13268 65584
rect 16387 65500 16396 65540
rect 16436 65500 17068 65540
rect 17108 65500 17117 65540
rect 18499 65500 18508 65540
rect 18548 65500 20084 65540
rect 20044 65456 20084 65500
rect 21510 65456 21600 65476
rect 13507 65416 13516 65456
rect 13556 65416 13632 65456
rect 14410 65416 14419 65456
rect 14459 65416 14764 65456
rect 14804 65416 14813 65456
rect 15497 65416 15628 65456
rect 15668 65416 15677 65456
rect 20044 65416 21600 65456
rect 13516 65372 13556 65416
rect 21510 65396 21600 65416
rect 13708 65372 13748 65381
rect 16204 65372 16244 65381
rect 17260 65372 17300 65381
rect 19948 65372 19988 65381
rect 6115 65332 6124 65372
rect 6164 65332 6173 65372
rect 7747 65332 7756 65372
rect 7796 65332 7805 65372
rect 9466 65332 9475 65372
rect 9515 65332 9524 65372
rect 9571 65332 9580 65372
rect 9620 65332 9629 65372
rect 9676 65332 10060 65372
rect 10100 65332 10109 65372
rect 10243 65332 10252 65372
rect 10292 65332 10301 65372
rect 10409 65332 10540 65372
rect 10580 65332 10589 65372
rect 11011 65332 11020 65372
rect 11068 65332 11191 65372
rect 11404 65332 12308 65372
rect 12634 65332 12643 65372
rect 12683 65332 12692 65372
rect 12739 65332 12748 65372
rect 12788 65332 12919 65372
rect 13219 65332 13228 65372
rect 13268 65332 13277 65372
rect 13411 65332 13420 65372
rect 13460 65332 13708 65372
rect 14083 65332 14092 65372
rect 14132 65332 14196 65372
rect 14236 65332 14263 65372
rect 14987 65332 15052 65372
rect 15092 65332 15118 65372
rect 15158 65332 15167 65372
rect 5740 65288 5780 65332
rect 7372 65288 7412 65332
rect 9004 65288 9044 65332
rect 10540 65323 10580 65332
rect 11404 65288 11444 65332
rect 5740 65248 6700 65288
rect 6740 65248 6749 65288
rect 7372 65248 7756 65288
rect 7796 65248 7805 65288
rect 9004 65248 10156 65288
rect 10196 65248 10205 65288
rect 10636 65248 11444 65288
rect 5801 65164 5932 65204
rect 5972 65164 5981 65204
rect 6700 65120 6740 65248
rect 10636 65204 10676 65248
rect 12268 65204 12308 65332
rect 12652 65288 12692 65332
rect 13708 65323 13748 65332
rect 15235 65331 15244 65371
rect 15284 65331 15293 65371
rect 15593 65332 15724 65372
rect 15764 65332 15773 65372
rect 16169 65332 16204 65372
rect 16244 65332 16300 65372
rect 16340 65332 16349 65372
rect 16675 65332 16684 65372
rect 16732 65332 16855 65372
rect 17225 65332 17260 65372
rect 17300 65332 17356 65372
rect 17396 65332 17405 65372
rect 18377 65332 18508 65372
rect 18548 65332 18557 65372
rect 18691 65332 18700 65372
rect 18740 65332 18749 65372
rect 19075 65332 19084 65372
rect 19124 65332 19948 65372
rect 15244 65288 15284 65331
rect 16204 65323 16244 65332
rect 12652 65248 13516 65288
rect 13556 65248 13565 65288
rect 13804 65248 14524 65288
rect 14564 65248 14573 65288
rect 14659 65248 14668 65288
rect 14708 65248 15284 65288
rect 16300 65288 16340 65332
rect 17260 65323 17300 65332
rect 18700 65288 18740 65332
rect 19948 65323 19988 65332
rect 16300 65248 16876 65288
rect 16916 65248 16925 65288
rect 17635 65248 17644 65288
rect 17684 65248 19180 65288
rect 19220 65248 19229 65288
rect 13804 65204 13844 65248
rect 7555 65164 7564 65204
rect 7604 65164 8524 65204
rect 8564 65164 8573 65204
rect 9187 65164 9196 65204
rect 9236 65164 9484 65204
rect 9524 65164 9533 65204
rect 9955 65164 9964 65204
rect 10004 65164 10676 65204
rect 11081 65164 11212 65204
rect 11252 65164 11261 65204
rect 11897 65164 11980 65204
rect 12020 65164 12028 65204
rect 12068 65164 12077 65204
rect 12268 65164 13844 65204
rect 14563 65164 14572 65204
rect 14612 65164 17740 65204
rect 17780 65164 17789 65204
rect 20131 65164 20140 65204
rect 20180 65164 21388 65204
rect 21428 65164 21437 65204
rect 6700 65080 11692 65120
rect 11732 65080 11741 65120
rect 4919 64996 4928 65036
rect 4968 64996 5010 65036
rect 5050 64996 5092 65036
rect 5132 64996 5174 65036
rect 5214 64996 5256 65036
rect 5296 64996 5305 65036
rect 5644 64996 8620 65036
rect 8660 64996 8669 65036
rect 8803 64996 8812 65036
rect 8852 64996 12940 65036
rect 12980 64996 12989 65036
rect 20039 64996 20048 65036
rect 20088 64996 20130 65036
rect 20170 64996 20212 65036
rect 20252 64996 20294 65036
rect 20334 64996 20376 65036
rect 20416 64996 20425 65036
rect 0 64952 90 64972
rect 21510 64952 21600 64972
rect 0 64912 556 64952
rect 596 64912 605 64952
rect 10147 64912 10156 64952
rect 10196 64912 11212 64952
rect 11252 64912 11261 64952
rect 21091 64912 21100 64952
rect 21140 64912 21600 64952
rect 0 64892 90 64912
rect 21510 64892 21600 64912
rect 3820 64828 4300 64868
rect 4340 64828 4349 64868
rect 9283 64828 9292 64868
rect 9332 64828 9341 64868
rect 9667 64828 9676 64868
rect 9716 64828 10252 64868
rect 10292 64828 10301 64868
rect 13961 64828 14092 64868
rect 14132 64828 14141 64868
rect 16099 64828 16108 64868
rect 16148 64828 16684 64868
rect 16724 64828 16733 64868
rect 19171 64828 19180 64868
rect 19220 64828 20428 64868
rect 20468 64828 20477 64868
rect 3820 64784 3860 64828
rect 9292 64784 9332 64828
rect 2170 64744 2179 64784
rect 2219 64744 3860 64784
rect 4108 64744 4492 64784
rect 4532 64744 4541 64784
rect 5356 64744 8276 64784
rect 8323 64744 8332 64784
rect 8372 64744 9140 64784
rect 9292 64744 9721 64784
rect 4108 64700 4148 64744
rect 2362 64660 2371 64700
rect 2411 64660 2668 64700
rect 2708 64660 2717 64700
rect 2860 64691 3052 64700
rect 2900 64660 3052 64691
rect 3092 64660 3101 64700
rect 3209 64660 3340 64700
rect 3380 64660 3389 64700
rect 3689 64660 3820 64700
rect 3860 64660 3869 64700
rect 3929 64660 3938 64700
rect 3978 64660 4148 64700
rect 4282 64660 4291 64700
rect 4331 64660 4340 64700
rect 4387 64660 4396 64700
rect 4436 64660 4532 64700
rect 4649 64660 4684 64700
rect 4724 64660 4780 64700
rect 4820 64660 4829 64700
rect 5356 64691 5396 64744
rect 2860 64642 2900 64651
rect 0 64616 90 64636
rect 4300 64616 4340 64660
rect 0 64576 1228 64616
rect 1268 64576 1277 64616
rect 1411 64576 1420 64616
rect 1460 64576 1469 64616
rect 1673 64576 1708 64616
rect 1748 64576 1804 64616
rect 1844 64576 1853 64616
rect 3427 64576 3436 64616
rect 3476 64576 3628 64616
rect 3668 64576 3677 64616
rect 4012 64576 4340 64616
rect 0 64556 90 64576
rect 1420 64532 1460 64576
rect 4012 64532 4052 64576
rect 4492 64532 4532 64660
rect 5705 64660 5836 64700
rect 5876 64660 5885 64700
rect 6883 64660 6892 64700
rect 6932 64660 7180 64700
rect 7220 64660 7229 64700
rect 7747 64660 7756 64700
rect 7796 64660 8140 64700
rect 8180 64660 8189 64700
rect 5356 64642 5396 64651
rect 5836 64642 5876 64651
rect 8140 64642 8180 64651
rect 8236 64616 8276 64744
rect 9100 64700 9140 64744
rect 9681 64700 9721 64744
rect 10060 64700 10100 64828
rect 10147 64744 10156 64784
rect 10196 64744 11252 64784
rect 12067 64744 12076 64784
rect 12116 64744 12652 64784
rect 12692 64744 12701 64784
rect 14515 64744 14524 64784
rect 14564 64744 21100 64784
rect 21140 64744 21149 64784
rect 8393 64660 8515 64700
rect 8564 64660 8573 64700
rect 8681 64660 8812 64700
rect 8852 64660 8861 64700
rect 9091 64660 9100 64700
rect 9140 64660 9292 64700
rect 9332 64660 9341 64700
rect 9449 64660 9484 64700
rect 9524 64660 9571 64700
rect 9611 64660 9629 64700
rect 9672 64660 9681 64700
rect 9721 64660 9730 64700
rect 10051 64660 10060 64700
rect 10100 64660 10109 64700
rect 10476 64660 10540 64700
rect 10580 64691 10676 64700
rect 10580 64660 10636 64691
rect 10985 64660 11116 64700
rect 11156 64660 11165 64700
rect 10636 64616 10676 64651
rect 11116 64642 11156 64651
rect 11212 64616 11252 64744
rect 12268 64660 12652 64700
rect 12692 64660 12701 64700
rect 13795 64660 13804 64700
rect 13844 64691 13975 64700
rect 13844 64660 13900 64691
rect 12268 64616 12308 64660
rect 13940 64660 13975 64691
rect 14380 64660 14668 64700
rect 14708 64660 14717 64700
rect 15715 64660 15724 64700
rect 15764 64691 15956 64700
rect 15764 64660 15916 64691
rect 13900 64642 13940 64651
rect 4745 64576 4876 64616
rect 4916 64576 4925 64616
rect 6058 64576 6067 64616
rect 6107 64576 6412 64616
rect 6452 64576 6461 64616
rect 8236 64576 9004 64616
rect 9044 64576 9053 64616
rect 10051 64576 10060 64616
rect 10100 64576 10156 64616
rect 10196 64576 10231 64616
rect 10636 64576 11020 64616
rect 11060 64576 11069 64616
rect 11212 64576 12076 64616
rect 12116 64576 12268 64616
rect 12308 64576 12317 64616
rect 12451 64576 12460 64616
rect 12500 64576 12508 64616
rect 12548 64576 12748 64616
rect 12788 64576 12797 64616
rect 14275 64576 14284 64616
rect 14324 64576 14333 64616
rect 14284 64532 14324 64576
rect 1420 64492 2228 64532
rect 2467 64492 2476 64532
rect 2516 64492 4052 64532
rect 4291 64492 4300 64532
rect 4340 64492 4532 64532
rect 6115 64492 6124 64532
rect 6164 64492 6172 64532
rect 6212 64492 6295 64532
rect 8611 64492 8620 64532
rect 8660 64492 8956 64532
rect 8996 64492 9005 64532
rect 10060 64492 14324 64532
rect 2188 64448 2228 64492
rect 547 64408 556 64448
rect 596 64408 1180 64448
rect 1220 64408 1229 64448
rect 1555 64408 1564 64448
rect 1604 64408 1804 64448
rect 1844 64408 1853 64448
rect 2188 64408 3052 64448
rect 3092 64408 3101 64448
rect 4003 64408 4012 64448
rect 4052 64408 4061 64448
rect 8681 64408 8812 64448
rect 8852 64408 8861 64448
rect 4012 64364 4052 64408
rect 10060 64364 10100 64492
rect 14380 64448 14420 64660
rect 16579 64660 16588 64700
rect 16628 64660 16780 64700
rect 16820 64660 16972 64700
rect 17012 64660 17021 64700
rect 17836 64691 17876 64700
rect 15916 64642 15956 64651
rect 18211 64660 18220 64700
rect 18260 64660 18316 64700
rect 18356 64660 18391 64700
rect 19564 64691 19604 64700
rect 17836 64616 17876 64651
rect 19564 64616 19604 64651
rect 16387 64576 16396 64616
rect 16436 64576 17260 64616
rect 17300 64576 19604 64616
rect 20009 64576 20140 64616
rect 20180 64576 20189 64616
rect 20899 64576 20908 64616
rect 20948 64576 21044 64616
rect 11107 64408 11116 64448
rect 11156 64408 11347 64448
rect 11387 64408 11396 64448
rect 12451 64408 12460 64448
rect 12500 64408 14420 64448
rect 17897 64408 18028 64448
rect 18068 64408 18077 64448
rect 1411 64324 1420 64364
rect 1460 64324 2900 64364
rect 4012 64324 4300 64364
rect 4340 64324 4349 64364
rect 7939 64324 7948 64364
rect 7988 64324 10100 64364
rect 0 64280 90 64300
rect 0 64240 1132 64280
rect 1172 64240 1181 64280
rect 0 64220 90 64240
rect 2860 64196 2900 64324
rect 3679 64240 3688 64280
rect 3728 64240 3770 64280
rect 3810 64240 3852 64280
rect 3892 64240 3934 64280
rect 3974 64240 4016 64280
rect 4056 64240 4065 64280
rect 5059 64240 5068 64280
rect 5108 64240 5836 64280
rect 5876 64240 5885 64280
rect 7747 64240 7756 64280
rect 7796 64240 9868 64280
rect 9908 64240 12556 64280
rect 12596 64240 12605 64280
rect 12931 64240 12940 64280
rect 12980 64240 15436 64280
rect 15476 64240 15485 64280
rect 18799 64240 18808 64280
rect 18848 64240 18890 64280
rect 18930 64240 18972 64280
rect 19012 64240 19054 64280
rect 19094 64240 19136 64280
rect 19176 64240 19185 64280
rect 2860 64156 6124 64196
rect 6164 64156 6173 64196
rect 11299 64156 11308 64196
rect 11348 64156 12980 64196
rect 12940 64112 12980 64156
rect 4771 64072 4780 64112
rect 4820 64072 5692 64112
rect 5732 64072 5741 64112
rect 6316 64072 8756 64112
rect 9187 64072 9196 64112
rect 9236 64072 9436 64112
rect 9476 64072 9485 64112
rect 12940 64072 14804 64112
rect 14995 64072 15004 64112
rect 15044 64072 16684 64112
rect 16724 64072 16733 64112
rect 2947 63988 2956 64028
rect 2996 63988 3340 64028
rect 3380 63988 3389 64028
rect 6067 63988 6076 64028
rect 6116 63988 6220 64028
rect 6260 63988 6269 64028
rect 0 63944 90 63964
rect 6316 63944 6356 64072
rect 8716 64028 8756 64072
rect 8332 63988 8620 64028
rect 8660 63988 8669 64028
rect 8716 63988 11692 64028
rect 11732 63988 11741 64028
rect 12067 63988 12076 64028
rect 12116 63988 12404 64028
rect 8332 63944 8372 63988
rect 0 63904 748 63944
rect 788 63904 797 63944
rect 3331 63904 3340 63944
rect 3380 63904 3389 63944
rect 3715 63904 3724 63944
rect 3764 63904 5068 63944
rect 5108 63904 5117 63944
rect 5923 63904 5932 63944
rect 5972 63904 6316 63944
rect 6356 63904 6365 63944
rect 6569 63904 6700 63944
rect 6740 63904 6749 63944
rect 6892 63904 7756 63944
rect 7796 63904 7805 63944
rect 8093 63904 8140 63944
rect 8180 63904 8189 63944
rect 8236 63904 8372 63944
rect 8419 63904 8428 63944
rect 8468 63904 8660 63944
rect 8995 63904 9004 63944
rect 9044 63904 9091 63944
rect 9131 63904 9175 63944
rect 9545 63904 9676 63944
rect 9716 63904 9725 63944
rect 11683 63904 11692 63944
rect 11732 63904 12268 63944
rect 12308 63904 12317 63944
rect 0 63884 90 63904
rect 2764 63860 2804 63869
rect 1411 63820 1420 63860
rect 1460 63820 1516 63860
rect 1556 63820 1591 63860
rect 2729 63820 2764 63860
rect 2804 63820 2860 63860
rect 2900 63820 2909 63860
rect 2764 63811 2804 63820
rect 3340 63776 3380 63904
rect 5164 63860 5204 63869
rect 6892 63860 6932 63904
rect 8140 63860 8180 63904
rect 3785 63820 3916 63860
rect 3956 63820 4300 63860
rect 4340 63820 4349 63860
rect 5204 63820 6220 63860
rect 6260 63820 6269 63860
rect 6883 63820 6892 63860
rect 6932 63820 6941 63860
rect 7267 63820 7276 63860
rect 7316 63820 8140 63860
rect 5164 63811 5204 63820
rect 8140 63811 8180 63820
rect 8236 63776 8276 63904
rect 8620 63860 8660 63904
rect 11308 63860 11348 63869
rect 12364 63860 12404 63988
rect 14764 63944 14804 64072
rect 15043 63988 15052 64028
rect 15092 63988 15484 64028
rect 15524 63988 15533 64028
rect 15907 63988 15916 64028
rect 15956 63988 16148 64028
rect 12547 63904 12556 63944
rect 12596 63904 12652 63944
rect 12692 63904 12727 63944
rect 14563 63904 14572 63944
rect 14612 63904 14621 63944
rect 14755 63904 14764 63944
rect 14804 63904 14813 63944
rect 15139 63904 15148 63944
rect 15188 63904 15436 63944
rect 15476 63904 15485 63944
rect 15593 63904 15724 63944
rect 15764 63904 15773 63944
rect 13996 63860 14036 63869
rect 8393 63820 8515 63860
rect 8564 63820 8573 63860
rect 8620 63820 8951 63860
rect 8991 63820 9000 63860
rect 9187 63820 9196 63860
rect 9236 63820 9292 63860
rect 9332 63820 9484 63860
rect 9524 63820 9533 63860
rect 10051 63820 10060 63860
rect 10100 63820 10732 63860
rect 10772 63820 10781 63860
rect 11348 63820 11500 63860
rect 11540 63820 11980 63860
rect 12020 63820 12029 63860
rect 12364 63820 12748 63860
rect 12788 63820 12797 63860
rect 13123 63820 13132 63860
rect 13172 63820 13996 63860
rect 14036 63820 14045 63860
rect 14572 63859 14612 63904
rect 16108 63860 16148 63988
rect 18892 63988 19276 64028
rect 19316 63988 19325 64028
rect 16195 63904 16204 63944
rect 16244 63904 17356 63944
rect 17396 63904 17405 63944
rect 18473 63904 18508 63944
rect 18548 63904 18604 63944
rect 18644 63904 18653 63944
rect 17644 63860 17684 63869
rect 18892 63860 18932 63988
rect 19564 63944 19604 64576
rect 21004 64448 21044 64576
rect 21510 64448 21600 64468
rect 19747 64408 19756 64448
rect 19796 64408 19805 64448
rect 20371 64408 20380 64448
rect 20420 64408 20908 64448
rect 20948 64408 20957 64448
rect 21004 64408 21600 64448
rect 19555 63904 19564 63944
rect 19604 63904 19613 63944
rect 19180 63860 19220 63869
rect 19756 63860 19796 64408
rect 21510 64388 21600 64408
rect 19913 64072 19996 64112
rect 20036 64072 20044 64112
rect 20084 64072 20093 64112
rect 14764 63859 15916 63860
rect 14572 63820 15916 63859
rect 15956 63820 15965 63860
rect 16108 63820 16396 63860
rect 16436 63820 16445 63860
rect 17251 63820 17260 63860
rect 17300 63820 17644 63860
rect 11308 63811 11348 63820
rect 13996 63811 14036 63820
rect 14572 63819 14804 63820
rect 17644 63811 17684 63820
rect 17836 63820 18115 63860
rect 18155 63820 18164 63860
rect 18211 63820 18220 63860
rect 18260 63820 18391 63860
rect 18665 63820 18700 63860
rect 18740 63820 18796 63860
rect 18836 63820 18932 63860
rect 18979 63820 18988 63860
rect 19028 63820 19180 63860
rect 19220 63820 19229 63860
rect 19663 63820 19672 63860
rect 19712 63820 19796 63860
rect 20140 63988 20812 64028
rect 20852 63988 20861 64028
rect 17836 63776 17876 63820
rect 19180 63811 19220 63820
rect 20140 63776 20180 63988
rect 21510 63944 21600 63964
rect 20227 63904 20236 63944
rect 20276 63904 20285 63944
rect 21091 63904 21100 63944
rect 21140 63904 21600 63944
rect 2860 63736 3100 63776
rect 3140 63736 3149 63776
rect 3340 63736 4204 63776
rect 4244 63736 4253 63776
rect 5731 63736 5740 63776
rect 5780 63736 6460 63776
rect 6500 63736 6509 63776
rect 8236 63736 8660 63776
rect 8817 63736 8826 63776
rect 8866 63736 9196 63776
rect 9236 63736 9245 63776
rect 11772 63736 11788 63776
rect 11828 63736 11932 63776
rect 11972 63736 13228 63776
rect 13268 63736 13277 63776
rect 13324 63736 13748 63776
rect 14083 63736 14092 63776
rect 14132 63736 14332 63776
rect 14372 63736 14381 63776
rect 15379 63736 15388 63776
rect 15428 63736 17588 63776
rect 17827 63736 17836 63776
rect 17876 63736 17885 63776
rect 19564 63736 20180 63776
rect 2860 63692 2900 63736
rect 8620 63692 8660 63736
rect 13324 63692 13364 63736
rect 1228 63652 1708 63692
rect 1748 63652 1757 63692
rect 2083 63652 2092 63692
rect 2132 63652 2900 63692
rect 3148 63652 3484 63692
rect 3524 63652 3533 63692
rect 5225 63652 5356 63692
rect 5396 63652 5405 63692
rect 6115 63652 6124 63692
rect 6164 63652 7756 63692
rect 7796 63652 7805 63692
rect 8323 63652 8332 63692
rect 8372 63652 8381 63692
rect 8602 63652 8611 63692
rect 8651 63652 8660 63692
rect 8707 63652 8716 63692
rect 8756 63652 8765 63692
rect 8995 63652 9004 63692
rect 9044 63652 9283 63692
rect 9323 63652 9332 63692
rect 10051 63652 10060 63692
rect 10100 63652 11500 63692
rect 11540 63652 11549 63692
rect 12067 63652 12076 63692
rect 12116 63652 12316 63692
rect 12356 63652 12365 63692
rect 12940 63652 13364 63692
rect 13708 63692 13748 63736
rect 17548 63692 17588 63736
rect 19564 63692 19604 63736
rect 13708 63652 14036 63692
rect 14179 63652 14188 63692
rect 14228 63652 14380 63692
rect 14420 63652 14429 63692
rect 15235 63652 15244 63692
rect 15284 63652 15964 63692
rect 16004 63652 16013 63692
rect 17548 63652 19604 63692
rect 19721 63652 19852 63692
rect 19892 63652 19901 63692
rect 0 63608 90 63628
rect 1228 63608 1268 63652
rect 3148 63608 3188 63652
rect 0 63568 1268 63608
rect 1315 63568 1324 63608
rect 1364 63568 3188 63608
rect 3244 63568 7948 63608
rect 7988 63568 7997 63608
rect 0 63548 90 63568
rect 3244 63524 3284 63568
rect 1699 63484 1708 63524
rect 1748 63484 3284 63524
rect 4919 63484 4928 63524
rect 4968 63484 5010 63524
rect 5050 63484 5092 63524
rect 5132 63484 5174 63524
rect 5214 63484 5256 63524
rect 5296 63484 5305 63524
rect 4483 63400 4492 63440
rect 4532 63400 5588 63440
rect 5548 63356 5588 63400
rect 8332 63356 8372 63652
rect 8716 63608 8756 63652
rect 8716 63568 9428 63608
rect 11299 63568 11308 63608
rect 11348 63568 12652 63608
rect 12692 63568 12701 63608
rect 9388 63524 9428 63568
rect 12940 63524 12980 63652
rect 13996 63608 14036 63652
rect 20236 63608 20276 63904
rect 21510 63884 21600 63904
rect 20419 63652 20428 63692
rect 20468 63652 20564 63692
rect 13996 63568 15188 63608
rect 16675 63568 16684 63608
rect 16724 63568 18604 63608
rect 18644 63568 18653 63608
rect 18700 63568 20276 63608
rect 15148 63524 15188 63568
rect 18700 63524 18740 63568
rect 8611 63484 8620 63524
rect 8660 63484 8908 63524
rect 8948 63484 8957 63524
rect 9379 63484 9388 63524
rect 9428 63484 9437 63524
rect 11107 63484 11116 63524
rect 11156 63484 12980 63524
rect 13603 63484 13612 63524
rect 13652 63484 15052 63524
rect 15092 63484 15101 63524
rect 15148 63484 16300 63524
rect 16340 63484 16349 63524
rect 17251 63484 17260 63524
rect 17300 63484 18740 63524
rect 20039 63484 20048 63524
rect 20088 63484 20130 63524
rect 20170 63484 20212 63524
rect 20252 63484 20294 63524
rect 20334 63484 20376 63524
rect 20416 63484 20425 63524
rect 9955 63400 9964 63440
rect 10004 63400 12940 63440
rect 12980 63400 12989 63440
rect 13564 63400 13900 63440
rect 13940 63400 13949 63440
rect 18412 63400 18836 63440
rect 13564 63356 13604 63400
rect 18412 63356 18452 63400
rect 5539 63316 5548 63356
rect 5588 63316 5597 63356
rect 6691 63316 6700 63356
rect 6740 63316 7220 63356
rect 8332 63316 8948 63356
rect 9065 63316 9187 63356
rect 9236 63316 9245 63356
rect 9475 63316 9484 63356
rect 9524 63316 9676 63356
rect 9716 63316 9725 63356
rect 12403 63316 12412 63356
rect 12452 63316 12556 63356
rect 12596 63316 12605 63356
rect 13555 63316 13564 63356
rect 13604 63316 13613 63356
rect 13900 63316 14668 63356
rect 14708 63316 14717 63356
rect 15523 63316 15532 63356
rect 15572 63316 15724 63356
rect 15764 63316 15773 63356
rect 15907 63316 15916 63356
rect 15956 63316 18452 63356
rect 18796 63356 18836 63400
rect 20524 63356 20564 63652
rect 21510 63440 21600 63460
rect 21187 63400 21196 63440
rect 21236 63400 21600 63440
rect 21510 63380 21600 63400
rect 18796 63316 19852 63356
rect 19892 63316 19901 63356
rect 20227 63316 20236 63356
rect 20276 63316 20564 63356
rect 0 63272 90 63292
rect 7180 63272 7220 63316
rect 8908 63272 8948 63316
rect 0 63232 1228 63272
rect 1268 63232 1277 63272
rect 5404 63232 7124 63272
rect 7180 63232 8428 63272
rect 8468 63232 8477 63272
rect 8803 63232 8812 63272
rect 8852 63232 8861 63272
rect 8908 63232 9140 63272
rect 0 63212 90 63232
rect 5404 63188 5444 63232
rect 7084 63188 7124 63232
rect 1411 63148 1420 63188
rect 1460 63148 1708 63188
rect 1748 63148 1757 63188
rect 2659 63148 2668 63188
rect 2708 63179 2996 63188
rect 2708 63148 2956 63179
rect 3785 63148 3916 63188
rect 3956 63148 3965 63188
rect 4771 63148 4780 63188
rect 4820 63179 5444 63188
rect 4820 63148 5164 63179
rect 2956 63130 2996 63139
rect 5204 63148 5444 63179
rect 5740 63179 5780 63188
rect 5164 63130 5204 63139
rect 6595 63148 6604 63188
rect 6644 63148 6988 63188
rect 7028 63148 7037 63188
rect 7084 63148 7756 63188
rect 7796 63148 7805 63188
rect 7913 63148 8044 63188
rect 8084 63148 8093 63188
rect 8236 63148 8299 63188
rect 8339 63148 8348 63188
rect 5740 63104 5780 63139
rect 1411 63064 1420 63104
rect 1460 63064 1516 63104
rect 1556 63064 1591 63104
rect 3523 63064 3532 63104
rect 3572 63064 3581 63104
rect 5260 63064 5780 63104
rect 7363 63064 7372 63104
rect 7412 63064 7564 63104
rect 7604 63064 7613 63104
rect 7747 63064 7756 63104
rect 7796 63064 8140 63104
rect 8180 63064 8189 63104
rect 3532 63020 3572 63064
rect 5260 63020 5300 63064
rect 8236 63020 8276 63148
rect 1891 62980 1900 63020
rect 1940 62980 3292 63020
rect 3332 62980 3341 63020
rect 3532 62980 4012 63020
rect 4052 62980 4061 63020
rect 4963 62980 4972 63020
rect 5012 62980 5300 63020
rect 5347 62980 5356 63020
rect 5396 62980 5452 63020
rect 5492 62980 5527 63020
rect 6691 62980 6700 63020
rect 6740 62980 8276 63020
rect 0 62936 90 62956
rect 8428 62936 8468 63232
rect 8812 63188 8852 63232
rect 9100 63188 9140 63232
rect 9580 63232 9868 63272
rect 9908 63232 9917 63272
rect 9580 63188 9620 63232
rect 13900 63188 13940 63316
rect 13996 63232 20948 63272
rect 8812 63148 8855 63188
rect 8895 63148 8904 63188
rect 9091 63148 9100 63188
rect 9140 63148 9149 63188
rect 9257 63148 9388 63188
rect 9428 63148 9437 63188
rect 9562 63148 9571 63188
rect 9611 63148 9620 63188
rect 9667 63148 9676 63188
rect 9716 63148 9772 63188
rect 9812 63148 9847 63188
rect 9955 63148 9964 63188
rect 10004 63148 10013 63188
rect 10217 63148 10348 63188
rect 10388 63148 10828 63188
rect 10868 63148 10877 63188
rect 11465 63148 11500 63188
rect 11540 63179 11636 63188
rect 11540 63148 11596 63179
rect 9100 63104 9140 63148
rect 9964 63104 10004 63148
rect 11683 63148 11692 63188
rect 11732 63148 12748 63188
rect 12788 63148 13364 63188
rect 13603 63148 13612 63188
rect 13652 63148 13795 63188
rect 13835 63148 13844 63188
rect 13891 63148 13900 63188
rect 13940 63148 13949 63188
rect 11596 63130 11636 63139
rect 13324 63104 13364 63148
rect 8873 63064 8995 63104
rect 9044 63064 9053 63104
rect 9100 63064 10004 63104
rect 12041 63064 12172 63104
rect 12212 63064 12221 63104
rect 12931 63064 12940 63104
rect 12980 63064 12989 63104
rect 13315 63064 13324 63104
rect 13364 63064 13373 63104
rect 12940 63020 12980 63064
rect 13996 63020 14036 63232
rect 14249 63148 14284 63188
rect 14324 63148 14380 63188
rect 14420 63148 14429 63188
rect 14825 63179 14956 63188
rect 14825 63148 14860 63179
rect 14900 63148 14956 63179
rect 14996 63148 15005 63188
rect 15340 63179 15380 63188
rect 14860 63130 14900 63139
rect 15340 63104 15380 63139
rect 15916 63179 15956 63188
rect 16963 63148 16972 63188
rect 17012 63148 17164 63188
rect 17204 63148 17213 63188
rect 17963 63148 18028 63188
rect 18068 63148 18094 63188
rect 18134 63148 18143 63188
rect 18209 63148 18218 63188
rect 18260 63148 18391 63188
rect 18499 63148 18508 63188
rect 18548 63148 18604 63188
rect 18644 63148 18679 63188
rect 19049 63148 19180 63188
rect 19220 63148 19229 63188
rect 19660 63179 20276 63188
rect 15916 63104 15956 63139
rect 18220 63104 18260 63148
rect 19180 63104 19220 63139
rect 19700 63148 20276 63179
rect 19660 63130 19700 63139
rect 14083 63064 14092 63104
rect 14132 63064 14380 63104
rect 14420 63064 14429 63104
rect 15043 63064 15052 63104
rect 15092 63064 15380 63104
rect 15436 63064 15956 63104
rect 17635 63064 17644 63104
rect 17684 63064 17693 63104
rect 17827 63064 17836 63104
rect 17876 63064 18260 63104
rect 18665 63064 18700 63104
rect 18740 63064 18796 63104
rect 18836 63064 18845 63104
rect 19180 63064 19468 63104
rect 19508 63064 19517 63104
rect 20131 63064 20140 63104
rect 20180 63064 20189 63104
rect 8515 62980 8524 63020
rect 8564 62980 8716 63020
rect 8756 62980 8765 63020
rect 9379 62980 9388 63020
rect 9428 62980 12980 63020
rect 13171 62980 13180 63020
rect 13220 62980 14036 63020
rect 14380 62936 14420 63064
rect 15436 62936 15476 63064
rect 17644 63020 17684 63064
rect 15532 62980 17684 63020
rect 0 62896 404 62936
rect 451 62896 460 62936
rect 500 62896 1180 62936
rect 1220 62896 1229 62936
rect 3017 62896 3148 62936
rect 3188 62896 3197 62936
rect 5731 62896 5740 62936
rect 5780 62896 7132 62936
rect 7172 62896 7181 62936
rect 7507 62896 7516 62936
rect 7556 62896 7565 62936
rect 8428 62896 11020 62936
rect 11060 62896 11069 62936
rect 11657 62896 11692 62936
rect 11732 62896 11788 62936
rect 11828 62896 11837 62936
rect 14371 62896 14380 62936
rect 14420 62896 14429 62936
rect 15427 62896 15436 62936
rect 15476 62896 15485 62936
rect 0 62876 90 62896
rect 364 62852 404 62896
rect 7516 62852 7556 62896
rect 364 62812 7556 62852
rect 10060 62812 15052 62852
rect 15092 62812 15101 62852
rect 10060 62768 10100 62812
rect 15532 62768 15572 62980
rect 15715 62896 15724 62936
rect 15764 62896 16012 62936
rect 16052 62896 16061 62936
rect 17875 62896 17884 62936
rect 17924 62896 18028 62936
rect 18068 62896 18077 62936
rect 18700 62852 18740 63064
rect 20140 63020 20180 63064
rect 18979 62980 18988 63020
rect 19028 62980 20180 63020
rect 20236 62936 20276 63148
rect 20908 62936 20948 63232
rect 21510 62936 21600 62956
rect 15811 62812 15820 62852
rect 15860 62812 18740 62852
rect 20140 62896 20276 62936
rect 20371 62896 20380 62936
rect 20420 62896 20812 62936
rect 20852 62896 20861 62936
rect 20908 62896 21600 62936
rect 1507 62728 1516 62768
rect 1556 62728 3620 62768
rect 3679 62728 3688 62768
rect 3728 62728 3770 62768
rect 3810 62728 3852 62768
rect 3892 62728 3934 62768
rect 3974 62728 4016 62768
rect 4056 62728 4065 62768
rect 4867 62728 4876 62768
rect 4916 62728 6604 62768
rect 6644 62728 6653 62768
rect 7084 62728 10100 62768
rect 10627 62728 10636 62768
rect 10676 62728 15572 62768
rect 18799 62728 18808 62768
rect 18848 62728 18890 62768
rect 18930 62728 18972 62768
rect 19012 62728 19054 62768
rect 19094 62728 19136 62768
rect 19176 62728 19185 62768
rect 3580 62684 3620 62728
rect 7084 62684 7124 62728
rect 1420 62644 2860 62684
rect 2900 62644 2909 62684
rect 3580 62644 7124 62684
rect 7747 62644 7756 62684
rect 7796 62644 13132 62684
rect 13172 62644 13420 62684
rect 13460 62644 13469 62684
rect 16012 62644 17260 62684
rect 17300 62644 17316 62684
rect 0 62600 90 62620
rect 1420 62600 1460 62644
rect 0 62560 1460 62600
rect 1612 62560 5740 62600
rect 5780 62560 5789 62600
rect 6220 62560 6700 62600
rect 6740 62560 7084 62600
rect 7124 62560 7133 62600
rect 8899 62560 8908 62600
rect 8948 62560 9388 62600
rect 9428 62560 9437 62600
rect 9514 62560 9523 62600
rect 9563 62560 9676 62600
rect 9716 62560 9725 62600
rect 10435 62560 10444 62600
rect 10484 62560 10580 62600
rect 13385 62560 13516 62600
rect 13556 62560 13565 62600
rect 13987 62560 13996 62600
rect 14036 62560 14332 62600
rect 14372 62560 14381 62600
rect 0 62540 90 62560
rect 1219 62308 1228 62348
rect 1268 62308 1420 62348
rect 1460 62308 1469 62348
rect 0 62264 90 62284
rect 1612 62264 1652 62560
rect 2851 62476 2860 62516
rect 2900 62476 5644 62516
rect 5684 62476 5693 62516
rect 6220 62432 6260 62560
rect 6307 62476 6316 62516
rect 6356 62476 6365 62516
rect 7555 62476 7564 62516
rect 7604 62476 8180 62516
rect 10147 62476 10156 62516
rect 10196 62476 10484 62516
rect 6316 62432 6356 62476
rect 3043 62392 3052 62432
rect 3092 62392 3860 62432
rect 3907 62392 3916 62432
rect 3956 62392 4204 62432
rect 4244 62392 4253 62432
rect 5740 62392 5932 62432
rect 5972 62392 5981 62432
rect 6211 62392 6220 62432
rect 6260 62392 6269 62432
rect 6316 62392 6836 62432
rect 2476 62348 2516 62357
rect 2516 62308 2764 62348
rect 2804 62308 2813 62348
rect 2947 62308 2956 62348
rect 2996 62308 3427 62348
rect 3467 62308 3476 62348
rect 3523 62308 3532 62348
rect 3572 62308 3628 62348
rect 3668 62308 3703 62348
rect 2476 62299 2516 62308
rect 0 62224 1652 62264
rect 0 62204 90 62224
rect 2275 62140 2284 62180
rect 2324 62140 2668 62180
rect 2708 62140 2717 62180
rect 2764 62140 2812 62180
rect 2852 62140 2861 62180
rect 2764 62096 2804 62140
rect 1507 62056 1516 62096
rect 1556 62056 2804 62096
rect 3820 62096 3860 62392
rect 4492 62348 4532 62357
rect 5740 62348 5780 62392
rect 6796 62348 6836 62392
rect 7756 62392 8044 62432
rect 8084 62392 8093 62432
rect 7756 62348 7796 62392
rect 8140 62348 8180 62476
rect 10444 62432 10484 62476
rect 8227 62392 8236 62432
rect 8276 62392 8524 62432
rect 8564 62392 8573 62432
rect 9964 62392 10060 62432
rect 10100 62392 10109 62432
rect 10435 62392 10444 62432
rect 10484 62392 10493 62432
rect 8812 62348 8852 62357
rect 9964 62348 10004 62392
rect 10540 62348 10580 62560
rect 16012 62516 16052 62644
rect 12259 62476 12268 62516
rect 12308 62476 12748 62516
rect 12788 62476 13748 62516
rect 13708 62432 13748 62476
rect 14284 62476 16052 62516
rect 13699 62392 13708 62432
rect 13748 62392 13757 62432
rect 13987 62392 13996 62432
rect 14036 62392 14092 62432
rect 14132 62392 14167 62432
rect 11020 62348 11060 62357
rect 13324 62348 13364 62357
rect 14284 62348 14324 62476
rect 14371 62392 14380 62432
rect 14420 62392 14996 62432
rect 15113 62392 15244 62432
rect 15284 62392 15293 62432
rect 14956 62348 14996 62392
rect 15820 62348 15860 62357
rect 17116 62348 17156 62644
rect 20140 62600 20180 62896
rect 21510 62876 21600 62896
rect 18019 62560 18028 62600
rect 18068 62560 18796 62600
rect 18836 62560 18845 62600
rect 19843 62560 19852 62600
rect 19892 62560 20180 62600
rect 17251 62476 17260 62516
rect 17300 62476 18452 62516
rect 18595 62476 18604 62516
rect 18644 62476 20276 62516
rect 17932 62348 17972 62357
rect 18412 62348 18452 62476
rect 20236 62432 20276 62476
rect 21510 62432 21600 62452
rect 20009 62392 20044 62432
rect 20084 62392 20140 62432
rect 20180 62392 20189 62432
rect 20236 62392 21600 62432
rect 21510 62372 21600 62392
rect 19660 62348 19700 62357
rect 4003 62308 4012 62348
rect 4052 62308 4183 62348
rect 4361 62308 4492 62348
rect 4532 62308 4541 62348
rect 5002 62308 5011 62348
rect 5051 62308 5356 62348
rect 5396 62308 5405 62348
rect 5718 62308 5727 62348
rect 5767 62308 5780 62348
rect 5827 62308 5836 62348
rect 5876 62308 6260 62348
rect 6307 62308 6316 62348
rect 6356 62308 6644 62348
rect 4492 62299 4532 62308
rect 6220 62264 6260 62308
rect 6220 62224 6316 62264
rect 6356 62224 6365 62264
rect 6604 62180 6644 62308
rect 7306 62308 7315 62348
rect 7355 62308 7372 62348
rect 7412 62308 7495 62348
rect 7738 62308 7747 62348
rect 7787 62308 7796 62348
rect 7843 62308 7852 62348
rect 7892 62308 8180 62348
rect 8323 62308 8332 62348
rect 8372 62308 8716 62348
rect 8756 62308 8765 62348
rect 9322 62308 9331 62348
rect 9371 62308 9484 62348
rect 9524 62308 9533 62348
rect 9946 62308 9955 62348
rect 9995 62308 10004 62348
rect 10051 62308 10060 62348
rect 10100 62308 10109 62348
rect 10531 62308 10540 62348
rect 10580 62308 10589 62348
rect 10819 62308 10828 62348
rect 10868 62308 11020 62348
rect 11530 62308 11539 62348
rect 11579 62308 11692 62348
rect 11732 62308 11741 62348
rect 12041 62308 12076 62348
rect 12116 62308 12172 62348
rect 12212 62308 12221 62348
rect 6796 62299 6836 62308
rect 8812 62264 8852 62308
rect 10060 62264 10100 62308
rect 6892 62224 8852 62264
rect 9955 62224 9964 62264
rect 10004 62224 10100 62264
rect 10540 62264 10580 62308
rect 11020 62299 11060 62308
rect 13324 62264 13364 62308
rect 13948 62308 14324 62348
rect 14746 62308 14755 62348
rect 14795 62308 14804 62348
rect 14851 62308 14860 62348
rect 14900 62308 14909 62348
rect 14956 62308 15340 62348
rect 15380 62308 15724 62348
rect 15764 62308 15773 62348
rect 15860 62308 15956 62348
rect 16003 62308 16012 62348
rect 16052 62308 16308 62348
rect 16348 62308 16357 62348
rect 16553 62308 16684 62348
rect 16724 62308 16733 62348
rect 17116 62308 17932 62348
rect 17972 62308 18220 62348
rect 18260 62308 18269 62348
rect 18403 62308 18412 62348
rect 18452 62308 18461 62348
rect 19555 62308 19564 62348
rect 19604 62308 19660 62348
rect 19700 62308 19735 62348
rect 13948 62264 13988 62308
rect 14764 62264 14804 62308
rect 10540 62224 10964 62264
rect 13324 62224 13948 62264
rect 13988 62224 13997 62264
rect 14476 62224 14804 62264
rect 14860 62264 14900 62308
rect 15820 62299 15860 62308
rect 15916 62264 15956 62308
rect 17932 62299 17972 62308
rect 14860 62224 15244 62264
rect 15284 62224 15293 62264
rect 15907 62224 15916 62264
rect 15956 62224 16492 62264
rect 16532 62224 16541 62264
rect 6892 62180 6932 62224
rect 8812 62180 8852 62224
rect 10924 62180 10964 62224
rect 5155 62140 5164 62180
rect 5204 62140 5548 62180
rect 5588 62140 5597 62180
rect 6595 62140 6604 62180
rect 6644 62140 6932 62180
rect 7459 62140 7468 62180
rect 7508 62140 7756 62180
rect 7796 62140 7805 62180
rect 8812 62140 10828 62180
rect 10868 62140 10877 62180
rect 10924 62140 11500 62180
rect 11540 62140 11549 62180
rect 11683 62140 11692 62180
rect 11732 62140 14380 62180
rect 14420 62140 14429 62180
rect 3820 62056 9964 62096
rect 10004 62056 10013 62096
rect 2179 61972 2188 62012
rect 2228 61972 4820 62012
rect 4919 61972 4928 62012
rect 4968 61972 5010 62012
rect 5050 61972 5092 62012
rect 5132 61972 5174 62012
rect 5214 61972 5256 62012
rect 5296 61972 5305 62012
rect 5356 61972 7412 62012
rect 7459 61972 7468 62012
rect 7508 61972 9484 62012
rect 9524 61972 9533 62012
rect 0 61928 90 61948
rect 4780 61928 4820 61972
rect 5356 61928 5396 61972
rect 0 61888 1036 61928
rect 1076 61888 1085 61928
rect 4780 61888 5396 61928
rect 7372 61928 7412 61972
rect 7372 61888 7564 61928
rect 7604 61888 7613 61928
rect 0 61868 90 61888
rect 14476 61844 14516 62224
rect 14860 62180 14900 62224
rect 18412 62180 18452 62308
rect 19660 62299 19700 62308
rect 14659 62140 14668 62180
rect 14708 62140 14900 62180
rect 15811 62140 15820 62180
rect 15860 62140 16492 62180
rect 16532 62140 16541 62180
rect 17993 62140 18124 62180
rect 18164 62140 18173 62180
rect 18412 62140 19564 62180
rect 19604 62140 19613 62180
rect 20371 62140 20380 62180
rect 20420 62140 20908 62180
rect 20948 62140 20957 62180
rect 19948 62056 21044 62096
rect 19948 62012 19988 62056
rect 18787 61972 18796 62012
rect 18836 61972 19988 62012
rect 20039 61972 20048 62012
rect 20088 61972 20130 62012
rect 20170 61972 20212 62012
rect 20252 61972 20294 62012
rect 20334 61972 20376 62012
rect 20416 61972 20425 62012
rect 16867 61888 16876 61928
rect 16916 61888 17932 61928
rect 17972 61888 17981 61928
rect 4771 61804 4780 61844
rect 4820 61804 5308 61844
rect 5348 61804 5357 61844
rect 5404 61804 6316 61844
rect 6356 61804 6365 61844
rect 7241 61804 7372 61844
rect 7412 61804 7421 61844
rect 7948 61804 10732 61844
rect 10772 61804 10781 61844
rect 11107 61804 11116 61844
rect 11156 61804 11404 61844
rect 11444 61804 11453 61844
rect 11731 61804 11740 61844
rect 11780 61804 12268 61844
rect 12308 61804 12317 61844
rect 13481 61804 13612 61844
rect 13652 61804 13661 61844
rect 14476 61804 15244 61844
rect 15284 61804 15293 61844
rect 17347 61804 17356 61844
rect 17396 61804 18124 61844
rect 18164 61804 18173 61844
rect 18499 61804 18508 61844
rect 18548 61804 19028 61844
rect 20131 61804 20140 61844
rect 20180 61804 20716 61844
rect 20756 61804 20765 61844
rect 5404 61760 5444 61804
rect 1708 61720 2956 61760
rect 2996 61720 3005 61760
rect 3532 61720 5444 61760
rect 5635 61720 5644 61760
rect 5684 61720 7516 61760
rect 7556 61720 7565 61760
rect 1708 61676 1748 61720
rect 3532 61676 3572 61720
rect 7948 61676 7988 61804
rect 9379 61720 9388 61760
rect 9428 61720 9437 61760
rect 12835 61720 12844 61760
rect 12884 61720 15092 61760
rect 16195 61720 16204 61760
rect 16244 61720 17492 61760
rect 9388 61676 9428 61720
rect 15052 61676 15092 61720
rect 1699 61636 1708 61676
rect 1748 61636 1757 61676
rect 2755 61636 2764 61676
rect 2804 61667 2996 61676
rect 2804 61636 2956 61667
rect 3275 61636 3340 61676
rect 3380 61636 3406 61676
rect 3446 61636 3455 61676
rect 3523 61636 3532 61676
rect 3572 61636 3581 61676
rect 3907 61636 3916 61676
rect 3956 61636 4204 61676
rect 4244 61636 4253 61676
rect 4361 61636 4492 61676
rect 4532 61636 4780 61676
rect 4820 61636 4829 61676
rect 4972 61667 5452 61676
rect 2956 61618 2996 61627
rect 4492 61618 4532 61627
rect 5012 61636 5452 61667
rect 5492 61636 5501 61676
rect 5923 61636 5932 61676
rect 5972 61636 6124 61676
rect 6164 61636 6173 61676
rect 6691 61636 6700 61676
rect 6740 61667 7220 61676
rect 6740 61636 7180 61667
rect 4972 61618 5012 61627
rect 7939 61636 7948 61676
rect 7988 61636 7997 61676
rect 9196 61667 9332 61676
rect 7180 61618 7220 61627
rect 9236 61636 9332 61667
rect 9388 61636 9667 61676
rect 9707 61636 9716 61676
rect 9763 61636 9772 61676
rect 9812 61636 9868 61676
rect 9908 61636 9943 61676
rect 10025 61636 10156 61676
rect 10196 61636 10205 61676
rect 10697 61667 10828 61676
rect 10697 61636 10732 61667
rect 9196 61618 9236 61627
rect 0 61592 90 61612
rect 0 61552 652 61592
rect 692 61552 701 61592
rect 1411 61552 1420 61592
rect 1460 61552 2900 61592
rect 3881 61552 4012 61592
rect 4052 61552 4061 61592
rect 5417 61552 5548 61592
rect 5588 61552 5597 61592
rect 7625 61552 7756 61592
rect 7796 61552 7805 61592
rect 0 61532 90 61552
rect 2860 61508 2900 61552
rect 2860 61468 6260 61508
rect 163 61384 172 61424
rect 212 61384 1180 61424
rect 1220 61384 1229 61424
rect 3139 61384 3148 61424
rect 3188 61384 3532 61424
rect 3572 61384 3581 61424
rect 5164 61384 5203 61424
rect 5243 61384 5252 61424
rect 5164 61340 5204 61384
rect 5164 61300 6164 61340
rect 0 61256 90 61276
rect 0 61216 1996 61256
rect 2036 61216 2045 61256
rect 3679 61216 3688 61256
rect 3728 61216 3770 61256
rect 3810 61216 3852 61256
rect 3892 61216 3934 61256
rect 3974 61216 4016 61256
rect 4056 61216 4065 61256
rect 0 61196 90 61216
rect 2563 60964 2572 61004
rect 2612 60964 5500 61004
rect 5540 60964 5549 61004
rect 0 60920 90 60940
rect 6124 60920 6164 61300
rect 6220 61172 6260 61468
rect 9292 61424 9332 61636
rect 10772 61636 10828 61667
rect 10868 61636 10877 61676
rect 11212 61667 11252 61676
rect 10732 61618 10772 61627
rect 12041 61636 12172 61676
rect 12212 61636 12221 61676
rect 13289 61636 13420 61676
rect 13460 61636 13469 61676
rect 13699 61636 13708 61676
rect 13748 61636 13804 61676
rect 13844 61636 13879 61676
rect 15052 61667 15436 61676
rect 11212 61592 11252 61627
rect 13420 61618 13460 61627
rect 15092 61636 15436 61667
rect 15476 61636 15485 61676
rect 16378 61636 16387 61676
rect 16427 61636 16436 61676
rect 16483 61636 16492 61676
rect 16532 61636 16541 61676
rect 16867 61636 16876 61676
rect 16916 61636 17068 61676
rect 17108 61636 17117 61676
rect 17452 61667 17492 61720
rect 18988 61676 19028 61804
rect 21004 61760 21044 62056
rect 21510 61928 21600 61948
rect 21091 61888 21100 61928
rect 21140 61888 21600 61928
rect 21510 61868 21600 61888
rect 21004 61720 21100 61760
rect 21140 61720 21149 61760
rect 15052 61618 15092 61627
rect 10243 61552 10252 61592
rect 10292 61552 10676 61592
rect 11107 61552 11116 61592
rect 11156 61552 11252 61592
rect 11971 61552 11980 61592
rect 12020 61552 12844 61592
rect 12884 61552 12893 61592
rect 15689 61552 15724 61592
rect 15764 61552 15820 61592
rect 15860 61552 15869 61592
rect 16099 61552 16108 61592
rect 16148 61552 16300 61592
rect 16340 61552 16349 61592
rect 10636 61508 10676 61552
rect 16396 61508 16436 61636
rect 16492 61508 16532 61636
rect 17452 61618 17492 61627
rect 17932 61667 17972 61676
rect 18115 61636 18124 61676
rect 18164 61636 18403 61676
rect 18443 61636 18452 61676
rect 18499 61636 18508 61676
rect 18548 61636 18604 61676
rect 18644 61636 18679 61676
rect 18796 61636 18892 61676
rect 18932 61636 19028 61676
rect 19337 61636 19468 61676
rect 19508 61636 19517 61676
rect 19948 61667 20084 61676
rect 16867 61552 16876 61592
rect 16916 61552 16972 61592
rect 17012 61552 17047 61592
rect 17932 61508 17972 61627
rect 18796 61592 18836 61636
rect 19468 61618 19508 61627
rect 19988 61636 20084 61667
rect 19948 61618 19988 61627
rect 18019 61552 18028 61592
rect 18068 61552 18836 61592
rect 18979 61552 18988 61592
rect 19028 61552 19159 61592
rect 10636 61468 11500 61508
rect 11540 61468 11549 61508
rect 12931 61468 12940 61508
rect 12980 61468 15868 61508
rect 15908 61468 15917 61508
rect 16387 61468 16396 61508
rect 16436 61468 16445 61508
rect 16492 61468 17356 61508
rect 17396 61468 17405 61508
rect 17932 61468 18164 61508
rect 9292 61384 12172 61424
rect 12212 61384 12221 61424
rect 14371 61384 14380 61424
rect 14420 61384 15484 61424
rect 15524 61384 15533 61424
rect 8803 61216 8812 61256
rect 8852 61216 14708 61256
rect 6220 61132 13612 61172
rect 13652 61132 13661 61172
rect 11107 61048 11116 61088
rect 11156 61048 11500 61088
rect 11540 61048 11549 61088
rect 14057 61048 14140 61088
rect 14180 61048 14188 61088
rect 14228 61048 14237 61088
rect 7555 60964 7564 61004
rect 7604 60964 7756 61004
rect 7796 60964 8180 61004
rect 0 60880 1612 60920
rect 1652 60880 1661 60920
rect 3043 60880 3052 60920
rect 3092 60880 3436 60920
rect 3476 60880 3485 60920
rect 4003 60880 4012 60920
rect 4052 60880 4108 60920
rect 4148 60880 4183 60920
rect 5386 60880 5395 60920
rect 5435 60880 5740 60920
rect 5780 60880 5789 60920
rect 6115 60880 6124 60920
rect 6164 60880 6173 60920
rect 0 60860 90 60880
rect 2476 60836 2516 60845
rect 4684 60836 4724 60845
rect 7564 60836 7604 60845
rect 8140 60836 8180 60964
rect 9964 60964 12556 61004
rect 12596 60964 12605 61004
rect 8323 60880 8332 60920
rect 8372 60880 8524 60920
rect 8564 60880 8573 60920
rect 9100 60836 9140 60845
rect 9964 60836 10004 60964
rect 14668 60920 14708 61216
rect 18124 61088 18164 61468
rect 18799 61216 18808 61256
rect 18848 61216 18890 61256
rect 18930 61216 18972 61256
rect 19012 61216 19054 61256
rect 19094 61216 19136 61256
rect 19176 61216 19185 61256
rect 20044 61088 20084 61636
rect 21510 61424 21600 61444
rect 21379 61384 21388 61424
rect 21428 61384 21600 61424
rect 21510 61364 21600 61384
rect 16361 61048 16396 61088
rect 16436 61048 16492 61088
rect 16532 61048 16541 61088
rect 18115 61048 18124 61088
rect 18164 61048 18173 61088
rect 20035 61048 20044 61088
rect 20084 61048 20093 61088
rect 15778 60964 17932 61004
rect 17972 60964 18068 61004
rect 11587 60880 11596 60920
rect 11636 60880 12172 60920
rect 12212 60880 12221 60920
rect 14371 60880 14380 60920
rect 14420 60880 14429 60920
rect 14659 60880 14668 60920
rect 14708 60880 14717 60920
rect 11308 60836 11348 60845
rect 12748 60836 12788 60845
rect 14380 60836 14420 60880
rect 15778 60836 15818 60964
rect 1219 60796 1228 60836
rect 1268 60796 1996 60836
rect 2036 60796 2045 60836
rect 2516 60796 2668 60836
rect 2708 60796 2717 60836
rect 3139 60796 3148 60836
rect 3188 60796 3619 60836
rect 3659 60796 3668 60836
rect 3715 60796 3724 60836
rect 3764 60796 3820 60836
rect 3860 60796 3895 60836
rect 4195 60796 4204 60836
rect 4244 60796 4253 60836
rect 4579 60796 4588 60836
rect 4628 60796 4684 60836
rect 4724 60796 4759 60836
rect 5194 60796 5203 60836
rect 5243 60796 5548 60836
rect 5588 60796 5597 60836
rect 6307 60796 6316 60836
rect 6356 60796 6365 60836
rect 7267 60796 7276 60836
rect 7316 60796 7564 60836
rect 8026 60796 8035 60836
rect 8075 60796 8084 60836
rect 8131 60796 8140 60836
rect 8180 60796 8189 60836
rect 8585 60796 8620 60836
rect 8660 60796 8716 60836
rect 8756 60796 8765 60836
rect 9140 60796 9484 60836
rect 9524 60796 9533 60836
rect 9610 60796 9619 60836
rect 9659 60796 10004 60836
rect 10051 60796 10060 60836
rect 10100 60796 10348 60836
rect 10388 60796 10397 60836
rect 11348 60796 12172 60836
rect 12212 60796 12221 60836
rect 13865 60796 13996 60836
rect 14036 60796 14045 60836
rect 14380 60796 15052 60836
rect 15092 60796 15818 60836
rect 16300 60880 17740 60920
rect 17780 60880 17972 60920
rect 16300 60836 16340 60880
rect 17932 60836 17972 60880
rect 16675 60796 16684 60836
rect 16724 60796 16855 60836
rect 18028 60836 18068 60964
rect 21510 60920 21600 60940
rect 18211 60880 18220 60920
rect 18260 60880 19180 60920
rect 19220 60880 19892 60920
rect 21475 60880 21484 60920
rect 21524 60880 21600 60920
rect 19852 60836 19892 60880
rect 21510 60860 21600 60880
rect 18028 60796 18604 60836
rect 18644 60796 18653 60836
rect 2476 60787 2516 60796
rect 4204 60752 4244 60796
rect 4684 60787 4724 60796
rect 3907 60712 3916 60752
rect 3956 60712 4244 60752
rect 2537 60628 2668 60668
rect 2708 60628 2717 60668
rect 2764 60628 2812 60668
rect 2852 60628 2861 60668
rect 2947 60628 2956 60668
rect 2996 60628 4012 60668
rect 4052 60628 4061 60668
rect 4579 60628 4588 60668
rect 4628 60628 5884 60668
rect 5924 60628 5933 60668
rect 0 60584 90 60604
rect 2764 60584 2804 60628
rect 0 60544 940 60584
rect 980 60544 989 60584
rect 1507 60544 1516 60584
rect 1556 60544 2804 60584
rect 6316 60584 6356 60796
rect 7564 60787 7604 60796
rect 8044 60752 8084 60796
rect 9100 60787 9140 60796
rect 11308 60787 11348 60796
rect 12748 60752 12788 60796
rect 7747 60712 7756 60752
rect 7796 60712 8084 60752
rect 12316 60712 12596 60752
rect 12643 60712 12652 60752
rect 12692 60712 12788 60752
rect 9641 60628 9772 60668
rect 9812 60628 9821 60668
rect 12316 60584 12356 60712
rect 12556 60668 12596 60712
rect 14380 60668 14420 60796
rect 16300 60787 16340 60796
rect 17932 60787 17972 60796
rect 19852 60787 19892 60796
rect 12403 60628 12412 60668
rect 12452 60628 12500 60668
rect 12556 60628 14420 60668
rect 14899 60628 14908 60668
rect 14948 60628 18220 60668
rect 18260 60628 18269 60668
rect 6316 60544 12356 60584
rect 12460 60584 12500 60628
rect 12460 60544 20852 60584
rect 0 60524 90 60544
rect 4919 60460 4928 60500
rect 4968 60460 5010 60500
rect 5050 60460 5092 60500
rect 5132 60460 5174 60500
rect 5214 60460 5256 60500
rect 5296 60460 5305 60500
rect 7267 60460 7276 60500
rect 7316 60460 12652 60500
rect 12692 60460 12980 60500
rect 16195 60460 16204 60500
rect 16244 60460 16684 60500
rect 16724 60460 16733 60500
rect 20039 60460 20048 60500
rect 20088 60460 20130 60500
rect 20170 60460 20212 60500
rect 20252 60460 20294 60500
rect 20334 60460 20376 60500
rect 20416 60460 20425 60500
rect 12940 60416 12980 60460
rect 20812 60416 20852 60544
rect 21510 60416 21600 60436
rect 1420 60376 5356 60416
rect 5396 60376 5405 60416
rect 12940 60376 13556 60416
rect 0 60248 90 60268
rect 0 60208 1324 60248
rect 1364 60208 1373 60248
rect 0 60188 90 60208
rect 1420 60080 1460 60376
rect 13516 60332 13556 60376
rect 15340 60376 20716 60416
rect 20756 60376 20765 60416
rect 20812 60376 21600 60416
rect 15340 60332 15380 60376
rect 21510 60356 21600 60376
rect 1987 60292 1996 60332
rect 2036 60292 4396 60332
rect 4436 60292 4445 60332
rect 5417 60292 5548 60332
rect 5588 60292 5597 60332
rect 7891 60292 7900 60332
rect 7940 60292 8236 60332
rect 8276 60292 8285 60332
rect 12521 60292 12604 60332
rect 12644 60292 12652 60332
rect 12692 60292 12701 60332
rect 13516 60292 14140 60332
rect 14180 60292 14189 60332
rect 14899 60292 14908 60332
rect 14948 60292 15380 60332
rect 15427 60292 15436 60332
rect 15476 60292 17260 60332
rect 17300 60292 17309 60332
rect 2188 60208 2284 60248
rect 2324 60208 2333 60248
rect 2572 60208 12268 60248
rect 12308 60208 12317 60248
rect 15820 60208 16012 60248
rect 16052 60208 16061 60248
rect 16108 60208 16204 60248
rect 16244 60208 16253 60248
rect 17155 60208 17164 60248
rect 17204 60208 19468 60248
rect 19508 60208 19517 60248
rect 2188 60164 2228 60208
rect 2170 60124 2179 60164
rect 2219 60124 2228 60164
rect 2275 60124 2284 60164
rect 2324 60124 2476 60164
rect 2516 60124 2525 60164
rect 2572 60080 2612 60208
rect 15820 60164 15860 60208
rect 16108 60164 16148 60208
rect 2659 60124 2668 60164
rect 2708 60124 2764 60164
rect 2804 60124 2839 60164
rect 3209 60155 3340 60164
rect 3209 60124 3244 60155
rect 3284 60124 3340 60155
rect 3380 60124 3389 60164
rect 3523 60124 3532 60164
rect 3572 60155 3764 60164
rect 3572 60124 3724 60155
rect 3244 60106 3284 60115
rect 4003 60124 4012 60164
rect 4052 60124 4108 60164
rect 4148 60124 4183 60164
rect 5356 60155 5644 60164
rect 3724 60106 3764 60115
rect 5396 60124 5644 60155
rect 5684 60124 5693 60164
rect 5801 60124 5836 60164
rect 5876 60124 5932 60164
rect 5972 60124 5981 60164
rect 6115 60124 6124 60164
rect 6164 60155 7124 60164
rect 6164 60124 7084 60155
rect 5356 60106 5396 60115
rect 7084 60106 7124 60115
rect 7660 60124 9100 60164
rect 9140 60124 10060 60164
rect 10100 60124 10109 60164
rect 10348 60155 10388 60164
rect 7660 60080 7700 60124
rect 10601 60124 10732 60164
rect 10772 60124 10781 60164
rect 11980 60155 12020 60164
rect 10348 60080 10388 60115
rect 15401 60124 15532 60164
rect 15572 60124 15581 60164
rect 15760 60124 15769 60164
rect 15809 60124 15860 60164
rect 15906 60124 15915 60164
rect 15955 60124 16148 60164
rect 16198 60124 16207 60164
rect 16247 60124 16291 60164
rect 16387 60124 16396 60164
rect 16436 60124 16567 60164
rect 16771 60124 16780 60164
rect 16820 60124 16829 60164
rect 16937 60124 17059 60164
rect 17108 60124 17117 60164
rect 17347 60124 17356 60164
rect 17396 60124 17644 60164
rect 17684 60124 17693 60164
rect 17818 60124 17827 60164
rect 17876 60124 18007 60164
rect 18499 60124 18508 60164
rect 18548 60124 18700 60164
rect 18740 60124 19660 60164
rect 19700 60124 19709 60164
rect 19913 60155 20044 60164
rect 19913 60124 19948 60155
rect 11980 60080 12020 60115
rect 67 60040 76 60080
rect 116 60040 1180 60080
rect 1220 60040 1229 60080
rect 1411 60040 1420 60080
rect 1460 60040 1469 60080
rect 1795 60040 1804 60080
rect 1844 60040 2612 60080
rect 2729 60040 2764 60080
rect 2804 60040 2860 60080
rect 2900 60040 2909 60080
rect 7651 60040 7660 60080
rect 7700 60040 7709 60080
rect 10348 60040 10924 60080
rect 10964 60040 12364 60080
rect 12404 60040 12460 60080
rect 12500 60040 12509 60080
rect 13001 60040 13036 60080
rect 13076 60040 13132 60080
rect 13172 60040 13181 60080
rect 13411 60040 13420 60080
rect 13460 60040 13469 60080
rect 14249 60040 14380 60080
rect 14420 60040 14429 60080
rect 14537 60040 14668 60080
rect 14708 60040 14717 60080
rect 14892 60040 14956 60080
rect 14996 60040 15052 60080
rect 15092 60040 15436 60080
rect 15476 60040 15485 60080
rect 15658 60071 15820 60080
rect 13420 59996 13460 60040
rect 15658 60031 15667 60071
rect 15707 60040 15820 60071
rect 15860 60040 15869 60080
rect 15707 60031 15716 60040
rect 15658 60030 15716 60031
rect 172 59956 2092 59996
rect 2132 59956 2141 59996
rect 3436 59956 3724 59996
rect 3764 59956 3773 59996
rect 4003 59956 4012 59996
rect 4052 59956 4148 59996
rect 0 59912 90 59932
rect 172 59912 212 59956
rect 0 59872 212 59912
rect 259 59872 268 59912
rect 308 59872 1564 59912
rect 1604 59872 1613 59912
rect 0 59852 90 59872
rect 0 59576 90 59596
rect 0 59536 1900 59576
rect 1940 59536 1949 59576
rect 0 59516 90 59536
rect 1289 59368 1420 59408
rect 1460 59368 1469 59408
rect 2860 59324 2900 59333
rect 3436 59324 3476 59956
rect 3532 59872 3955 59912
rect 3995 59872 4004 59912
rect 3532 59408 3572 59872
rect 3679 59704 3688 59744
rect 3728 59704 3770 59744
rect 3810 59704 3852 59744
rect 3892 59704 3934 59744
rect 3974 59704 4016 59744
rect 4056 59704 4065 59744
rect 4108 59660 4148 59956
rect 5932 59956 8812 59996
rect 8852 59956 8861 59996
rect 10444 59956 11156 59996
rect 11203 59956 11212 59996
rect 11252 59956 12796 59996
rect 12836 59956 13460 59996
rect 13987 59956 13996 59996
rect 14036 59956 14045 59996
rect 5932 59912 5972 59956
rect 10444 59912 10484 59956
rect 11116 59912 11156 59956
rect 5635 59872 5644 59912
rect 5684 59872 5972 59912
rect 7145 59872 7276 59912
rect 7316 59872 7325 59912
rect 8611 59872 8620 59912
rect 8660 59872 10484 59912
rect 10531 59872 10540 59912
rect 10580 59872 10589 59912
rect 11116 59872 11972 59912
rect 12041 59872 12172 59912
rect 12212 59872 12221 59912
rect 12643 59872 12652 59912
rect 12692 59872 13180 59912
rect 13220 59872 13229 59912
rect 10540 59828 10580 59872
rect 5731 59788 5740 59828
rect 5780 59788 6124 59828
rect 6164 59788 6173 59828
rect 10540 59788 10828 59828
rect 10868 59788 10877 59828
rect 11932 59744 11972 59872
rect 13996 59828 14036 59956
rect 15916 59912 15956 60124
rect 16204 60080 16244 60124
rect 16780 60080 16820 60124
rect 19988 60124 20044 60155
rect 20084 60124 20093 60164
rect 19948 60080 19988 60115
rect 16195 60040 16204 60080
rect 16244 60040 16820 60080
rect 18185 60040 18316 60080
rect 18356 60040 18365 60080
rect 19171 60040 19180 60080
rect 19220 60040 19988 60080
rect 16531 59956 16540 59996
rect 16580 59956 17548 59996
rect 17588 59956 17597 59996
rect 19948 59956 20428 59996
rect 20468 59956 20477 59996
rect 15283 59872 15292 59912
rect 15332 59872 16972 59912
rect 17012 59872 17021 59912
rect 17321 59872 17452 59912
rect 17492 59872 17501 59912
rect 17818 59872 17827 59912
rect 17867 59872 18412 59912
rect 18452 59872 18461 59912
rect 18547 59872 18556 59912
rect 18596 59872 19660 59912
rect 19700 59872 19709 59912
rect 19948 59828 19988 59956
rect 21510 59912 21600 59932
rect 20131 59872 20140 59912
rect 20180 59872 20189 59912
rect 21283 59872 21292 59912
rect 21332 59872 21600 59912
rect 13996 59788 19988 59828
rect 11932 59704 12980 59744
rect 18799 59704 18808 59744
rect 18848 59704 18890 59744
rect 18930 59704 18972 59744
rect 19012 59704 19054 59744
rect 19094 59704 19136 59744
rect 19176 59704 19185 59744
rect 4012 59620 4148 59660
rect 6691 59620 6700 59660
rect 6740 59620 11116 59660
rect 11156 59620 11165 59660
rect 3619 59536 3628 59576
rect 3668 59536 3676 59576
rect 3716 59536 3799 59576
rect 4012 59492 4052 59620
rect 12940 59576 12980 59704
rect 7721 59536 7804 59576
rect 7844 59536 7852 59576
rect 7892 59536 7901 59576
rect 8131 59536 8140 59576
rect 8180 59536 8188 59576
rect 8228 59536 8311 59576
rect 9283 59536 9292 59576
rect 9332 59536 11348 59576
rect 12931 59536 12940 59576
rect 12980 59536 12989 59576
rect 14659 59536 14668 59576
rect 14708 59536 15916 59576
rect 15956 59536 16396 59576
rect 16436 59536 16445 59576
rect 18796 59536 20044 59576
rect 20084 59536 20093 59576
rect 11308 59492 11348 59536
rect 18796 59492 18836 59536
rect 3715 59452 3724 59492
rect 3764 59452 4052 59492
rect 6115 59452 6124 59492
rect 6164 59452 6316 59492
rect 6356 59452 6365 59492
rect 10819 59452 10828 59492
rect 10868 59452 10877 59492
rect 11308 59452 11788 59492
rect 11828 59452 11837 59492
rect 15523 59452 15532 59492
rect 15572 59452 16300 59492
rect 16340 59452 16349 59492
rect 17932 59452 18796 59492
rect 18836 59452 18845 59492
rect 19084 59452 19468 59492
rect 19508 59452 19517 59492
rect 10828 59408 10868 59452
rect 3523 59368 3532 59408
rect 3572 59368 3581 59408
rect 3785 59368 3916 59408
rect 3956 59368 3965 59408
rect 5356 59368 5740 59408
rect 5780 59368 5789 59408
rect 5923 59368 5932 59408
rect 5972 59368 6316 59408
rect 6356 59368 6365 59408
rect 7913 59368 8044 59408
rect 8084 59368 8093 59408
rect 8419 59368 8428 59408
rect 8468 59368 8477 59408
rect 10732 59368 10868 59408
rect 11081 59368 11212 59408
rect 11252 59368 11261 59408
rect 5356 59324 5396 59368
rect 6892 59324 6932 59333
rect 8428 59324 8468 59368
rect 9004 59324 9044 59333
rect 10732 59324 10772 59368
rect 11308 59324 11348 59452
rect 12163 59368 12172 59408
rect 12212 59368 12356 59408
rect 12490 59368 12499 59408
rect 12539 59368 12844 59408
rect 12884 59368 12893 59408
rect 14476 59368 16148 59408
rect 12316 59324 12356 59368
rect 14476 59324 14516 59368
rect 16108 59324 16148 59368
rect 17932 59324 17972 59452
rect 18019 59368 18028 59408
rect 18068 59368 18892 59408
rect 18932 59368 18941 59408
rect 1603 59284 1612 59324
rect 1652 59284 2284 59324
rect 2324 59284 2333 59324
rect 2900 59284 3436 59324
rect 3476 59284 3485 59324
rect 4099 59284 4108 59324
rect 4148 59284 4396 59324
rect 4436 59284 4445 59324
rect 5818 59284 5827 59324
rect 5867 59284 5876 59324
rect 5923 59284 5932 59324
rect 5972 59284 6124 59324
rect 6164 59284 6173 59324
rect 6403 59284 6412 59324
rect 6452 59284 6604 59324
rect 6644 59284 6653 59324
rect 7267 59284 7276 59324
rect 7316 59284 7380 59324
rect 7420 59284 7447 59324
rect 7564 59284 8468 59324
rect 8611 59284 8620 59324
rect 8660 59284 8669 59324
rect 8873 59284 9004 59324
rect 9044 59284 9053 59324
rect 10217 59284 10252 59324
rect 10292 59284 10348 59324
rect 10388 59284 10397 59324
rect 10714 59284 10723 59324
rect 10763 59284 10772 59324
rect 10819 59284 10828 59324
rect 10868 59284 10999 59324
rect 11299 59284 11308 59324
rect 11348 59284 11357 59324
rect 11782 59284 11791 59324
rect 11831 59284 11924 59324
rect 12298 59284 12307 59324
rect 12347 59284 12356 59324
rect 12931 59284 12940 59324
rect 12980 59284 13228 59324
rect 13268 59284 13277 59324
rect 14345 59284 14380 59324
rect 14420 59284 14476 59324
rect 14851 59284 14860 59324
rect 14900 59284 14956 59324
rect 14996 59284 15031 59324
rect 16387 59284 16396 59324
rect 16436 59284 16588 59324
rect 16628 59284 16684 59324
rect 16724 59284 16733 59324
rect 18394 59284 18403 59324
rect 18443 59284 18452 59324
rect 18499 59284 18508 59324
rect 18548 59284 18604 59324
rect 18644 59284 18679 59324
rect 2860 59275 2900 59284
rect 5356 59275 5396 59284
rect 0 59240 90 59260
rect 5836 59240 5876 59284
rect 6892 59240 6932 59284
rect 0 59200 1804 59240
rect 1844 59200 1853 59240
rect 3043 59200 3052 59240
rect 3092 59200 3820 59240
rect 3860 59200 3869 59240
rect 5539 59200 5548 59240
rect 5588 59200 5876 59240
rect 6403 59200 6412 59240
rect 6452 59200 6932 59240
rect 0 59180 90 59200
rect 7564 59156 7604 59284
rect 8620 59240 8660 59284
rect 9004 59275 9044 59284
rect 7843 59200 7852 59240
rect 7892 59200 8660 59240
rect 11884 59240 11924 59284
rect 14476 59275 14516 59284
rect 16108 59275 16148 59284
rect 17932 59275 17972 59284
rect 18412 59240 18452 59284
rect 11884 59200 12268 59240
rect 12308 59200 12317 59240
rect 18115 59200 18124 59240
rect 18164 59200 18452 59240
rect 18892 59156 18932 59368
rect 19084 59324 19124 59452
rect 19468 59324 19508 59333
rect 20140 59324 20180 59872
rect 21510 59852 21600 59872
rect 21510 59408 21600 59428
rect 20419 59368 20428 59408
rect 20468 59368 21600 59408
rect 21510 59348 21600 59368
rect 18979 59284 18988 59324
rect 19028 59284 19124 59324
rect 19337 59284 19468 59324
rect 19508 59284 19517 59324
rect 19978 59284 19987 59324
rect 20027 59284 20180 59324
rect 19468 59275 19508 59284
rect 19564 59200 21292 59240
rect 21332 59200 21341 59240
rect 19564 59156 19604 59200
rect 739 59116 748 59156
rect 788 59116 1180 59156
rect 1220 59116 1229 59156
rect 3043 59116 3052 59156
rect 3092 59116 3292 59156
rect 3332 59116 3341 59156
rect 7555 59116 7564 59156
rect 7604 59116 7613 59156
rect 8611 59116 8620 59156
rect 8660 59116 8812 59156
rect 8852 59116 8861 59156
rect 10147 59116 10156 59156
rect 10196 59116 10828 59156
rect 10868 59116 10877 59156
rect 10924 59116 12604 59156
rect 12644 59116 12653 59156
rect 16291 59116 16300 59156
rect 16340 59116 18028 59156
rect 18068 59116 18077 59156
rect 18892 59116 19604 59156
rect 20131 59116 20140 59156
rect 20180 59116 20189 59156
rect 10924 59072 10964 59116
rect 20140 59072 20180 59116
rect 4780 59032 5396 59072
rect 7555 59032 7564 59072
rect 7604 59032 10964 59072
rect 16291 59032 16300 59072
rect 16340 59032 20180 59072
rect 4780 58988 4820 59032
rect 5356 58988 5396 59032
rect 2755 58948 2764 58988
rect 2804 58948 4820 58988
rect 4919 58948 4928 58988
rect 4968 58948 5010 58988
rect 5050 58948 5092 58988
rect 5132 58948 5174 58988
rect 5214 58948 5256 58988
rect 5296 58948 5305 58988
rect 5356 58948 5932 58988
rect 5972 58948 5981 58988
rect 6796 58948 13708 58988
rect 13748 58948 13757 58988
rect 20039 58948 20048 58988
rect 20088 58948 20130 58988
rect 20170 58948 20212 58988
rect 20252 58948 20294 58988
rect 20334 58948 20376 58988
rect 20416 58948 20425 58988
rect 0 58904 90 58924
rect 0 58864 556 58904
rect 596 58864 605 58904
rect 1804 58864 6740 58904
rect 0 58844 90 58864
rect 1324 58612 1612 58652
rect 1652 58612 1661 58652
rect 0 58568 90 58588
rect 1324 58568 1364 58612
rect 1804 58568 1844 58864
rect 3881 58780 3916 58820
rect 3956 58780 4012 58820
rect 4052 58780 4061 58820
rect 4867 58780 4876 58820
rect 4916 58780 5588 58820
rect 5705 58780 5788 58820
rect 5828 58780 5836 58820
rect 5876 58780 5885 58820
rect 5548 58736 5588 58780
rect 2284 58696 2668 58736
rect 2708 58696 2717 58736
rect 2851 58696 2860 58736
rect 2900 58696 2909 58736
rect 3427 58696 3436 58736
rect 3476 58696 5492 58736
rect 5548 58696 6548 58736
rect 2284 58652 2324 58696
rect 2266 58612 2275 58652
rect 2315 58612 2324 58652
rect 2371 58612 2380 58652
rect 2420 58612 2476 58652
rect 2516 58612 2551 58652
rect 2633 58612 2764 58652
rect 2804 58612 2813 58652
rect 2860 58568 2900 58696
rect 5452 58652 5492 58696
rect 3209 58612 3340 58652
rect 3380 58612 3389 58652
rect 3689 58612 3820 58652
rect 3860 58612 3869 58652
rect 4195 58612 4204 58652
rect 4244 58612 4876 58652
rect 4916 58612 4925 58652
rect 5452 58643 5644 58652
rect 3340 58594 3380 58603
rect 3820 58594 3860 58603
rect 4204 58568 4244 58612
rect 5492 58612 5644 58643
rect 5684 58612 5693 58652
rect 6019 58612 6028 58652
rect 6068 58612 6452 58652
rect 5452 58594 5492 58603
rect 6412 58568 6452 58612
rect 0 58528 1364 58568
rect 1411 58528 1420 58568
rect 1460 58528 1469 58568
rect 1795 58528 1804 58568
rect 1844 58528 1853 58568
rect 2659 58528 2668 58568
rect 2708 58528 2860 58568
rect 2900 58528 2909 58568
rect 3907 58528 3916 58568
rect 3956 58528 4244 58568
rect 5539 58528 5548 58568
rect 5588 58528 6028 58568
rect 6068 58528 6077 58568
rect 6403 58528 6412 58568
rect 6452 58528 6461 58568
rect 0 58508 90 58528
rect 1420 58484 1460 58528
rect 1420 58444 2380 58484
rect 2420 58444 2429 58484
rect 2860 58444 6172 58484
rect 6212 58444 6221 58484
rect 643 58360 652 58400
rect 692 58360 1180 58400
rect 1220 58360 1229 58400
rect 1411 58360 1420 58400
rect 1460 58360 1564 58400
rect 1604 58360 1613 58400
rect 0 58232 90 58252
rect 0 58192 460 58232
rect 500 58192 509 58232
rect 0 58172 90 58192
rect 2860 58148 2900 58444
rect 6508 58400 6548 58696
rect 6700 58484 6740 58864
rect 6796 58652 6836 58948
rect 21510 58904 21600 58924
rect 7171 58864 7180 58904
rect 7220 58864 8812 58904
rect 8852 58864 9292 58904
rect 9332 58864 9341 58904
rect 9475 58864 9484 58904
rect 9524 58864 10772 58904
rect 10732 58820 10772 58864
rect 8227 58780 8236 58820
rect 8276 58780 10196 58820
rect 10714 58780 10723 58820
rect 10763 58780 10772 58820
rect 10828 58864 11348 58904
rect 11683 58864 11692 58904
rect 11732 58864 12076 58904
rect 12116 58864 12125 58904
rect 14755 58864 14764 58904
rect 14804 58864 16012 58904
rect 16052 58864 16061 58904
rect 18211 58864 18220 58904
rect 18260 58864 21600 58904
rect 8393 58696 8419 58736
rect 8459 58696 8524 58736
rect 8564 58696 8573 58736
rect 9100 58696 9676 58736
rect 9716 58696 9725 58736
rect 6787 58612 6796 58652
rect 6836 58612 6845 58652
rect 8044 58643 8084 58652
rect 8489 58612 8611 58652
rect 8660 58612 8669 58652
rect 9100 58643 9140 58696
rect 10156 58672 10196 58780
rect 10828 58736 10868 58864
rect 11308 58736 11348 58864
rect 21510 58844 21600 58864
rect 12979 58780 12988 58820
rect 13028 58780 13036 58820
rect 13076 58780 13159 58820
rect 15043 58780 15052 58820
rect 15092 58780 16204 58820
rect 16244 58780 16253 58820
rect 17155 58780 17164 58820
rect 17204 58780 17780 58820
rect 17827 58780 17836 58820
rect 17876 58780 17932 58820
rect 17972 58780 18007 58820
rect 16204 58736 16244 58780
rect 10749 58696 10868 58736
rect 11251 58696 11260 58736
rect 11300 58696 11348 58736
rect 12163 58696 12172 58736
rect 12212 58696 14956 58736
rect 14996 58696 15005 58736
rect 15436 58696 15916 58736
rect 15956 58696 15965 58736
rect 16204 58696 17012 58736
rect 17211 58696 17260 58736
rect 17300 58696 17342 58736
rect 17382 58696 17391 58736
rect 17443 58696 17452 58736
rect 17492 58696 17684 58736
rect 8044 58568 8084 58603
rect 9283 58612 9292 58652
rect 9332 58612 9580 58652
rect 9620 58612 9629 58652
rect 10051 58612 10060 58652
rect 10100 58612 10109 58652
rect 10156 58632 10173 58672
rect 10213 58632 10222 58672
rect 10749 58652 10789 58696
rect 15436 58652 15476 58696
rect 10442 58612 10540 58652
rect 10604 58612 10622 58652
rect 10714 58612 10723 58652
rect 10763 58612 10789 58652
rect 10840 58612 10867 58652
rect 10907 58612 10916 58652
rect 9100 58594 9140 58603
rect 10060 58568 10100 58612
rect 10840 58568 10880 58612
rect 11002 58601 11011 58641
rect 11051 58601 11060 58641
rect 11104 58612 11113 58652
rect 11156 58612 11287 58652
rect 11395 58612 11404 58652
rect 11444 58612 11500 58652
rect 11540 58612 11575 58652
rect 12172 58612 13612 58652
rect 13652 58612 13996 58652
rect 14036 58612 14045 58652
rect 14371 58612 14380 58652
rect 14420 58643 14900 58652
rect 14420 58612 14860 58643
rect 8044 58528 9004 58568
rect 9044 58528 9053 58568
rect 9571 58528 9580 58568
rect 9620 58528 9676 58568
rect 9716 58528 9751 58568
rect 10060 58528 10156 58568
rect 10196 58528 10205 58568
rect 10819 58528 10828 58568
rect 10868 58528 10880 58568
rect 11020 58484 11060 58601
rect 11596 58528 11788 58568
rect 11828 58528 11837 58568
rect 6700 58444 10924 58484
rect 10964 58444 10973 58484
rect 11020 58444 11212 58484
rect 11252 58444 11261 58484
rect 5635 58360 5644 58400
rect 5684 58360 5693 58400
rect 6508 58360 10444 58400
rect 10484 58360 10493 58400
rect 3679 58192 3688 58232
rect 3728 58192 3770 58232
rect 3810 58192 3852 58232
rect 3892 58192 3934 58232
rect 3974 58192 4016 58232
rect 4056 58192 4065 58232
rect 1420 58108 2900 58148
rect 0 57896 90 57916
rect 1420 57896 1460 58108
rect 5290 58024 5299 58064
rect 5339 58024 5548 58064
rect 5588 58024 5597 58064
rect 5644 57980 5684 58360
rect 11107 58108 11116 58148
rect 11156 58108 11540 58148
rect 11500 58064 11540 58108
rect 10531 58024 10540 58064
rect 10580 58024 11308 58064
rect 11348 58024 11357 58064
rect 11491 58024 11500 58064
rect 11540 58024 11549 58064
rect 11596 57980 11636 58528
rect 12172 58484 12212 58612
rect 15418 58612 15427 58652
rect 15467 58612 15476 58652
rect 15523 58612 15532 58652
rect 15572 58612 15581 58652
rect 14860 58594 14900 58603
rect 12739 58528 12748 58568
rect 12788 58528 12797 58568
rect 13001 58528 13132 58568
rect 13172 58528 13181 58568
rect 12748 58484 12788 58528
rect 15532 58484 15572 58612
rect 12163 58444 12172 58484
rect 12212 58444 12221 58484
rect 12748 58444 13420 58484
rect 13460 58444 13469 58484
rect 14467 58444 14476 58484
rect 14516 58444 15572 58484
rect 12019 58360 12028 58400
rect 12068 58360 12980 58400
rect 13363 58360 13372 58400
rect 13412 58360 14188 58400
rect 14228 58360 14237 58400
rect 12940 58316 12980 58360
rect 12940 58276 15052 58316
rect 15092 58276 15101 58316
rect 12067 58192 12076 58232
rect 12116 58192 15428 58232
rect 15388 58064 15428 58192
rect 11779 58024 11788 58064
rect 11828 58024 11837 58064
rect 14275 58024 14284 58064
rect 14324 58024 14332 58064
rect 14372 58024 14455 58064
rect 14947 58024 14956 58064
rect 14996 58024 15004 58064
rect 15044 58024 15127 58064
rect 15379 58024 15388 58064
rect 15428 58024 15437 58064
rect 5068 57940 5684 57980
rect 6691 57940 6700 57980
rect 6740 57940 10924 57980
rect 10964 57940 10973 57980
rect 11116 57940 11636 57980
rect 11788 57980 11828 58024
rect 11788 57940 12116 57980
rect 14563 57940 14572 57980
rect 14612 57940 14908 57980
rect 14948 57940 14957 57980
rect 15043 57940 15052 57980
rect 15092 57940 15668 57980
rect 0 57856 1460 57896
rect 2860 57856 3436 57896
rect 3476 57856 3485 57896
rect 4003 57856 4012 57896
rect 4052 57856 4204 57896
rect 4244 57856 4253 57896
rect 0 57836 90 57856
rect 2764 57812 2804 57821
rect 2860 57812 2900 57856
rect 5068 57845 5108 57940
rect 6953 57856 7084 57896
rect 7124 57856 7133 57896
rect 8995 57856 9004 57896
rect 9044 57856 11020 57896
rect 11060 57856 11069 57896
rect 4588 57812 4628 57821
rect 1315 57772 1324 57812
rect 1364 57772 1516 57812
rect 1556 57772 2420 57812
rect 0 57560 90 57580
rect 2380 57560 2420 57772
rect 2804 57772 2900 57812
rect 3514 57772 3523 57812
rect 3563 57772 3572 57812
rect 3619 57772 3628 57812
rect 3668 57772 3677 57812
rect 4003 57772 4012 57812
rect 4052 57772 4108 57812
rect 4148 57772 4183 57812
rect 4628 57772 4876 57812
rect 4916 57772 4925 57812
rect 8716 57812 8756 57821
rect 11116 57812 11156 57940
rect 12076 57854 12116 57940
rect 15628 57896 15668 57940
rect 14083 57856 14092 57896
rect 14132 57856 14141 57896
rect 14537 57856 14668 57896
rect 14708 57856 14717 57896
rect 15235 57856 15244 57896
rect 15284 57856 15572 57896
rect 15619 57856 15628 57896
rect 15668 57856 15677 57896
rect 12076 57845 12159 57854
rect 12076 57814 12119 57845
rect 5068 57796 5108 57805
rect 5627 57772 5636 57812
rect 5684 57772 5815 57812
rect 6761 57772 6892 57812
rect 6932 57772 6941 57812
rect 7459 57772 7468 57812
rect 7508 57772 7852 57812
rect 7892 57772 8140 57812
rect 8180 57772 8189 57812
rect 8611 57772 8620 57812
rect 8660 57772 8716 57812
rect 8756 57772 9196 57812
rect 9236 57772 9245 57812
rect 9859 57772 9868 57812
rect 9908 57772 10540 57812
rect 10580 57772 10589 57812
rect 10985 57772 11116 57812
rect 11156 57772 11165 57812
rect 11299 57772 11308 57812
rect 11348 57772 11500 57812
rect 11540 57772 11549 57812
rect 11606 57772 11615 57812
rect 11655 57772 11664 57812
rect 11779 57772 11788 57812
rect 11828 57772 11980 57812
rect 12020 57772 12029 57812
rect 13708 57812 13748 57821
rect 12119 57796 12159 57805
rect 12425 57772 12460 57812
rect 12500 57772 12556 57812
rect 12596 57772 12605 57812
rect 13315 57772 13324 57812
rect 13364 57772 13708 57812
rect 13748 57772 13900 57812
rect 13940 57772 13949 57812
rect 2764 57763 2804 57772
rect 3532 57728 3572 57772
rect 2947 57688 2956 57728
rect 2996 57688 3572 57728
rect 3628 57644 3668 57772
rect 4588 57763 4628 57772
rect 8716 57763 8756 57772
rect 11116 57763 11156 57772
rect 11615 57728 11655 57772
rect 10060 57688 10924 57728
rect 10964 57688 10973 57728
rect 11212 57688 11655 57728
rect 2467 57604 2476 57644
rect 2516 57604 3668 57644
rect 5443 57604 5452 57644
rect 5492 57604 6412 57644
rect 6452 57604 6461 57644
rect 7315 57604 7324 57644
rect 7364 57604 8044 57644
rect 8084 57604 8093 57644
rect 8899 57604 8908 57644
rect 8948 57604 9292 57644
rect 9332 57604 9341 57644
rect 10060 57560 10100 57688
rect 11212 57644 11252 57688
rect 11788 57644 11828 57772
rect 13708 57763 13748 57772
rect 14092 57728 14132 57856
rect 12067 57688 12076 57728
rect 12116 57688 12980 57728
rect 12940 57644 12980 57688
rect 13804 57688 14132 57728
rect 13804 57644 13844 57688
rect 15532 57644 15572 57856
rect 15724 57812 15764 58696
rect 15881 58612 15916 58652
rect 15956 58612 16012 58652
rect 16052 58612 16061 58652
rect 16492 58643 16876 58652
rect 16532 58612 16876 58643
rect 16916 58612 16925 58652
rect 16972 58643 17012 58696
rect 16492 58594 16532 58603
rect 17417 58612 17548 58652
rect 17588 58612 17597 58652
rect 17644 58643 17684 58696
rect 16972 58594 17012 58603
rect 17740 58652 17780 58780
rect 18787 58696 18796 58736
rect 18836 58696 19988 58736
rect 17740 58612 17836 58652
rect 17876 58612 17885 58652
rect 18019 58612 18028 58652
rect 18068 58612 18199 58652
rect 18691 58612 18700 58652
rect 18740 58612 19564 58652
rect 19604 58612 19613 58652
rect 19948 58643 19988 58696
rect 17644 58594 17684 58603
rect 16003 58528 16012 58568
rect 16052 58528 16300 58568
rect 16340 58528 16349 58568
rect 18281 58528 18412 58568
rect 18452 58528 18461 58568
rect 17225 58360 17347 58400
rect 17396 58360 17405 58400
rect 18163 58360 18172 58400
rect 18212 58360 18220 58400
rect 18260 58360 18343 58400
rect 19372 58316 19412 58612
rect 19948 58594 19988 58603
rect 21510 58400 21600 58420
rect 20131 58360 20140 58400
rect 20180 58360 20189 58400
rect 21091 58360 21100 58400
rect 21140 58360 21600 58400
rect 19363 58276 19372 58316
rect 19412 58276 19421 58316
rect 18799 58192 18808 58232
rect 18848 58192 18890 58232
rect 18930 58192 18972 58232
rect 19012 58192 19054 58232
rect 19094 58192 19136 58232
rect 19176 58192 19185 58232
rect 15811 58024 15820 58064
rect 15860 58024 15869 58064
rect 15820 57896 15860 58024
rect 16963 57940 16972 57980
rect 17012 57940 19412 57980
rect 15811 57856 15820 57896
rect 15860 57856 15869 57896
rect 16042 57887 16684 57896
rect 16042 57847 16051 57887
rect 16091 57856 16684 57887
rect 16724 57856 16733 57896
rect 18665 57856 18796 57896
rect 18836 57856 18845 57896
rect 16091 57847 16100 57856
rect 16042 57846 16100 57847
rect 17836 57812 17876 57821
rect 19372 57812 19412 57940
rect 20140 57812 20180 58360
rect 21510 58340 21600 58360
rect 21510 57896 21600 57916
rect 20707 57856 20716 57896
rect 20756 57856 21600 57896
rect 21510 57836 21600 57856
rect 15724 57772 15916 57812
rect 15956 57772 15965 57812
rect 16144 57772 16153 57812
rect 16193 57772 16204 57812
rect 16244 57772 16333 57812
rect 16428 57772 16492 57812
rect 16532 57772 16588 57812
rect 16628 57772 16780 57812
rect 16820 57772 16829 57812
rect 17876 57772 18028 57812
rect 18068 57772 18077 57812
rect 18298 57772 18307 57812
rect 18347 57772 18356 57812
rect 18403 57772 18412 57812
rect 18452 57772 18583 57812
rect 18761 57772 18892 57812
rect 18932 57772 18941 57812
rect 19882 57772 19891 57812
rect 19931 57772 20180 57812
rect 17836 57763 17876 57772
rect 18316 57728 18356 57772
rect 19372 57763 19412 57772
rect 18019 57688 18028 57728
rect 18068 57688 18356 57728
rect 10147 57604 10156 57644
rect 10196 57604 10772 57644
rect 10819 57604 10828 57644
rect 10868 57604 11252 57644
rect 11299 57604 11308 57644
rect 11348 57604 11828 57644
rect 12076 57604 12268 57644
rect 12308 57604 12317 57644
rect 12940 57604 13844 57644
rect 13891 57604 13900 57644
rect 13940 57604 14860 57644
rect 14900 57604 14909 57644
rect 15532 57604 20044 57644
rect 20084 57604 20093 57644
rect 0 57520 1516 57560
rect 1556 57520 1565 57560
rect 2380 57520 10100 57560
rect 10732 57560 10772 57604
rect 12076 57560 12116 57604
rect 10732 57520 11308 57560
rect 11348 57520 11357 57560
rect 12067 57520 12076 57560
rect 12116 57520 12125 57560
rect 12739 57520 12748 57560
rect 12788 57520 19852 57560
rect 19892 57520 19901 57560
rect 0 57500 90 57520
rect 4919 57436 4928 57476
rect 4968 57436 5010 57476
rect 5050 57436 5092 57476
rect 5132 57436 5174 57476
rect 5214 57436 5256 57476
rect 5296 57436 5305 57476
rect 5347 57436 5356 57476
rect 5396 57436 10100 57476
rect 13027 57436 13036 57476
rect 13076 57436 16820 57476
rect 20039 57436 20048 57476
rect 20088 57436 20130 57476
rect 20170 57436 20212 57476
rect 20252 57436 20294 57476
rect 20334 57436 20376 57476
rect 20416 57436 20425 57476
rect 10060 57392 10100 57436
rect 10060 57352 12884 57392
rect 14179 57352 14188 57392
rect 14228 57352 16436 57392
rect 2227 57268 2236 57308
rect 2276 57268 2668 57308
rect 2708 57268 2717 57308
rect 3139 57268 3148 57308
rect 3188 57268 6748 57308
rect 6788 57268 6797 57308
rect 10819 57268 10828 57308
rect 10868 57268 11308 57308
rect 11348 57268 11357 57308
rect 0 57224 90 57244
rect 0 57184 172 57224
rect 212 57184 221 57224
rect 2572 57184 3052 57224
rect 3092 57184 3101 57224
rect 4195 57184 4204 57224
rect 4244 57184 4253 57224
rect 4972 57184 5932 57224
rect 5972 57184 5981 57224
rect 6172 57184 8276 57224
rect 0 57164 90 57184
rect 2572 57056 2612 57184
rect 4204 57140 4244 57184
rect 4972 57140 5012 57184
rect 2659 57100 2668 57140
rect 2708 57100 2764 57140
rect 2804 57100 2839 57140
rect 3427 57100 3436 57140
rect 3476 57131 4052 57140
rect 3476 57100 4012 57131
rect 4204 57100 4867 57140
rect 4907 57100 4916 57140
rect 4963 57100 4972 57140
rect 5012 57100 5021 57140
rect 5347 57100 5356 57140
rect 5396 57100 5405 57140
rect 5539 57100 5548 57140
rect 5588 57131 5972 57140
rect 5588 57100 5932 57131
rect 4012 57082 4052 57091
rect 1411 57016 1420 57056
rect 1460 57016 1469 57056
rect 1673 57016 1804 57056
rect 1844 57016 1853 57056
rect 1987 57016 1996 57056
rect 2036 57016 2167 57056
rect 2563 57016 2572 57056
rect 2612 57016 2621 57056
rect 4457 57016 4588 57056
rect 4628 57016 4637 57056
rect 1420 56972 1460 57016
rect 5356 56972 5396 57100
rect 5932 57082 5972 57091
rect 5443 57016 5452 57056
rect 5492 57016 5876 57056
rect 5836 56972 5876 57016
rect 6172 56972 6212 57184
rect 8236 57140 8276 57184
rect 8812 57184 9484 57224
rect 9524 57184 9533 57224
rect 9868 57184 12556 57224
rect 12596 57184 12605 57224
rect 6281 57100 6412 57140
rect 6452 57100 6461 57140
rect 7738 57100 7747 57140
rect 7787 57100 7796 57140
rect 7843 57100 7852 57140
rect 7892 57100 8023 57140
rect 8227 57100 8236 57140
rect 8276 57100 8524 57140
rect 8564 57100 8573 57140
rect 8812 57131 8852 57184
rect 9868 57140 9908 57184
rect 6412 57082 6452 57091
rect 6634 57016 6643 57056
rect 6683 57016 6988 57056
rect 7028 57016 7037 57056
rect 1420 56932 2572 56972
rect 2612 56932 2621 56972
rect 2860 56932 4532 56972
rect 5356 56932 5644 56972
rect 5684 56932 5693 56972
rect 5836 56932 6124 56972
rect 6164 56932 6212 56972
rect 7756 56972 7796 57100
rect 9161 57100 9292 57140
rect 9332 57100 9341 57140
rect 9859 57100 9868 57140
rect 9908 57100 9917 57140
rect 10985 57100 11116 57140
rect 11156 57100 11165 57140
rect 11491 57100 11500 57140
rect 11540 57100 11788 57140
rect 11828 57100 11837 57140
rect 12617 57100 12652 57140
rect 12692 57131 12788 57140
rect 12692 57100 12748 57131
rect 8812 57082 8852 57091
rect 9292 57082 9332 57091
rect 11116 57082 11156 57091
rect 12748 57082 12788 57091
rect 12844 57056 12884 57352
rect 13324 57268 14476 57308
rect 14516 57268 14525 57308
rect 14947 57268 14956 57308
rect 14996 57268 15724 57308
rect 15764 57268 15773 57308
rect 12931 57184 12940 57224
rect 12980 57184 13268 57224
rect 13228 57140 13268 57184
rect 13324 57140 13364 57268
rect 13804 57184 16300 57224
rect 16340 57184 16349 57224
rect 13210 57100 13219 57140
rect 13259 57100 13268 57140
rect 13315 57100 13324 57140
rect 13364 57100 13420 57140
rect 13460 57100 13524 57140
rect 13699 57100 13708 57140
rect 13748 57100 13757 57140
rect 13708 57056 13748 57100
rect 13804 57056 13844 57184
rect 16396 57140 16436 57352
rect 16780 57224 16820 57436
rect 21510 57392 21600 57412
rect 20611 57352 20620 57392
rect 20660 57352 21600 57392
rect 21510 57332 21600 57352
rect 16867 57268 16876 57308
rect 16916 57268 18508 57308
rect 18548 57268 18557 57308
rect 16780 57184 17300 57224
rect 18115 57184 18124 57224
rect 18164 57184 18644 57224
rect 17260 57140 17300 57184
rect 18604 57140 18644 57184
rect 14153 57100 14284 57140
rect 14324 57100 14333 57140
rect 14764 57131 14804 57140
rect 14284 57082 14324 57091
rect 15305 57100 15340 57140
rect 15380 57100 15436 57140
rect 15476 57100 15724 57140
rect 15764 57100 15773 57140
rect 16396 57131 16628 57140
rect 16396 57100 16588 57131
rect 8297 57016 8332 57056
rect 8372 57016 8428 57056
rect 8468 57016 8477 57056
rect 12844 57016 13748 57056
rect 13795 57016 13804 57056
rect 13844 57016 13900 57056
rect 13940 57016 14004 57056
rect 13708 56972 13748 57016
rect 7756 56932 7852 56972
rect 7892 56932 7901 56972
rect 13708 56932 13804 56972
rect 13844 56932 13853 56972
rect 0 56888 90 56908
rect 2860 56888 2900 56932
rect 4492 56888 4532 56932
rect 0 56848 268 56888
rect 308 56848 317 56888
rect 451 56848 460 56888
rect 500 56848 1180 56888
rect 1220 56848 1229 56888
rect 1315 56848 1324 56888
rect 1364 56848 1564 56888
rect 1604 56848 1613 56888
rect 1795 56848 1804 56888
rect 1844 56848 2332 56888
rect 2372 56848 2381 56888
rect 2604 56848 2668 56888
rect 2708 56848 2900 56888
rect 3532 56848 4348 56888
rect 4388 56848 4397 56888
rect 4492 56848 6836 56888
rect 9514 56848 9523 56888
rect 9563 56848 9964 56888
rect 10004 56848 10013 56888
rect 0 56828 90 56848
rect 2764 56804 2804 56848
rect 835 56764 844 56804
rect 884 56764 2804 56804
rect 3532 56720 3572 56848
rect 172 56680 3572 56720
rect 3679 56680 3688 56720
rect 3728 56680 3770 56720
rect 3810 56680 3852 56720
rect 3892 56680 3934 56720
rect 3974 56680 4016 56720
rect 4056 56680 4065 56720
rect 0 56552 90 56572
rect 0 56512 76 56552
rect 116 56512 125 56552
rect 0 56492 90 56512
rect 0 56216 90 56236
rect 172 56216 212 56680
rect 3619 56512 3628 56552
rect 3668 56512 5932 56552
rect 5972 56512 5981 56552
rect 6796 56468 6836 56848
rect 6979 56764 6988 56804
rect 7028 56764 8084 56804
rect 8323 56764 8332 56804
rect 8372 56764 13900 56804
rect 13940 56764 13949 56804
rect 8044 56720 8084 56764
rect 8044 56680 12980 56720
rect 8323 56596 8332 56636
rect 8372 56596 12172 56636
rect 12212 56596 12221 56636
rect 7843 56512 7852 56552
rect 7892 56512 8044 56552
rect 8084 56512 8093 56552
rect 10051 56512 10060 56552
rect 10100 56512 10108 56552
rect 10148 56512 10231 56552
rect 12940 56468 12980 56680
rect 14764 56552 14804 57091
rect 16963 57100 16972 57140
rect 17012 57100 17164 57140
rect 17204 57100 17213 57140
rect 17260 57131 18260 57140
rect 17260 57100 18220 57131
rect 16588 57082 16628 57091
rect 18595 57100 18604 57140
rect 18644 57100 18653 57140
rect 19852 57131 19892 57140
rect 18220 57056 18260 57091
rect 19852 57056 19892 57091
rect 18220 57016 19892 57056
rect 18316 56932 20716 56972
rect 20756 56932 20765 56972
rect 16771 56848 16780 56888
rect 16820 56848 16876 56888
rect 16916 56848 16951 56888
rect 18316 56552 18356 56932
rect 21510 56888 21600 56908
rect 18403 56848 18412 56888
rect 18452 56848 18461 56888
rect 18700 56848 18796 56888
rect 18836 56848 18845 56888
rect 20035 56848 20044 56888
rect 20084 56848 20093 56888
rect 20803 56848 20812 56888
rect 20852 56848 21600 56888
rect 13027 56512 13036 56552
rect 13076 56512 14804 56552
rect 17971 56512 17980 56552
rect 18020 56512 18356 56552
rect 2860 56428 5404 56468
rect 5444 56428 5453 56468
rect 6796 56428 9908 56468
rect 12940 56428 17308 56468
rect 17348 56428 17357 56468
rect 2860 56384 2900 56428
rect 1411 56344 1420 56384
rect 1460 56344 2900 56384
rect 3139 56344 3148 56384
rect 3188 56344 4012 56384
rect 4052 56344 4204 56384
rect 4244 56344 4253 56384
rect 5290 56344 5299 56384
rect 5339 56344 5644 56384
rect 5684 56344 5693 56384
rect 6281 56344 6412 56384
rect 6452 56344 6461 56384
rect 6595 56344 6604 56384
rect 6644 56344 6653 56384
rect 7363 56344 7372 56384
rect 7412 56344 7756 56384
rect 7796 56344 7805 56384
rect 2956 56300 2996 56309
rect 4588 56300 4628 56309
rect 6604 56300 6644 56344
rect 7852 56300 7892 56309
rect 9772 56300 9812 56309
rect 835 56260 844 56300
rect 884 56260 1708 56300
rect 1748 56260 1757 56300
rect 2947 56260 2956 56300
rect 2996 56260 3127 56300
rect 3514 56260 3523 56300
rect 3563 56260 3572 56300
rect 3619 56260 3628 56300
rect 3668 56260 3799 56300
rect 4099 56260 4108 56300
rect 4148 56260 4492 56300
rect 4532 56260 4541 56300
rect 4628 56260 4780 56300
rect 4820 56260 4829 56300
rect 5098 56260 5107 56300
rect 5147 56260 5356 56300
rect 5396 56260 5405 56300
rect 5827 56260 5836 56300
rect 5876 56260 6609 56300
rect 6649 56260 6658 56300
rect 8323 56260 8332 56300
rect 8372 56260 8524 56300
rect 8564 56260 8573 56300
rect 9283 56260 9292 56300
rect 9332 56260 9772 56300
rect 9868 56300 9908 56428
rect 18412 56384 18452 56848
rect 18700 56384 18740 56848
rect 18799 56680 18808 56720
rect 18848 56680 18890 56720
rect 18930 56680 18972 56720
rect 19012 56680 19054 56720
rect 19094 56680 19136 56720
rect 19176 56680 19185 56720
rect 20044 56468 20084 56848
rect 21510 56828 21600 56848
rect 19756 56428 20084 56468
rect 9955 56344 9964 56384
rect 10004 56344 10348 56384
rect 10388 56344 10397 56384
rect 13411 56344 13420 56384
rect 13460 56344 13469 56384
rect 13673 56344 13804 56384
rect 13844 56344 13853 56384
rect 15689 56344 15820 56384
rect 15860 56344 16300 56384
rect 16340 56344 16349 56384
rect 16396 56344 17068 56384
rect 17108 56344 17117 56384
rect 17539 56344 17548 56384
rect 17588 56344 17597 56384
rect 17731 56344 17740 56384
rect 17780 56344 17911 56384
rect 18172 56344 18452 56384
rect 18665 56344 18700 56384
rect 18740 56344 18796 56384
rect 18836 56344 18845 56384
rect 12844 56300 12884 56309
rect 13420 56300 13460 56344
rect 14380 56300 14420 56309
rect 16396 56300 16436 56344
rect 9868 56260 10828 56300
rect 10868 56260 10877 56300
rect 11587 56260 11596 56300
rect 11636 56260 12076 56300
rect 12116 56260 12556 56300
rect 12596 56260 12605 56300
rect 13306 56260 13315 56300
rect 13355 56260 13364 56300
rect 13411 56260 13420 56300
rect 13460 56260 13507 56300
rect 13769 56260 13900 56300
rect 13940 56260 13949 56300
rect 14275 56260 14284 56300
rect 14324 56260 14380 56300
rect 14420 56260 14455 56300
rect 14746 56260 14860 56300
rect 14908 56260 14926 56300
rect 15043 56260 15052 56300
rect 15092 56260 15331 56300
rect 15371 56260 15380 56300
rect 15427 56260 15436 56300
rect 15476 56260 15607 56300
rect 15881 56260 15916 56300
rect 15956 56260 16012 56300
rect 16052 56260 16061 56300
rect 16771 56260 16780 56300
rect 16820 56260 16884 56300
rect 16924 56260 16951 56300
rect 2956 56251 2996 56260
rect 3532 56216 3572 56260
rect 0 56176 212 56216
rect 547 56176 556 56216
rect 596 56176 1180 56216
rect 1220 56176 1229 56216
rect 3139 56176 3148 56216
rect 3188 56176 3572 56216
rect 4588 56216 4628 56260
rect 4588 56176 5452 56216
rect 5492 56176 5501 56216
rect 0 56156 90 56176
rect 7852 56132 7892 56260
rect 9772 56251 9812 56260
rect 12844 56216 12884 56260
rect 10060 56176 12268 56216
rect 12308 56176 12317 56216
rect 12643 56176 12652 56216
rect 12692 56176 12884 56216
rect 13324 56216 13364 56260
rect 14380 56251 14420 56260
rect 16396 56216 16436 56260
rect 13324 56176 13420 56216
rect 13460 56176 13469 56216
rect 14659 56176 14668 56216
rect 14708 56176 15092 56216
rect 16291 56176 16300 56216
rect 16340 56176 16436 56216
rect 17059 56176 17068 56216
rect 17108 56176 17155 56216
rect 3043 56092 3052 56132
rect 3092 56092 5260 56132
rect 5300 56092 5309 56132
rect 6163 56092 6172 56132
rect 6212 56092 6221 56132
rect 7852 56092 8620 56132
rect 8660 56092 8669 56132
rect 9833 56092 9964 56132
rect 10004 56092 10013 56132
rect 6172 56048 6212 56092
rect 10060 56048 10100 56176
rect 15052 56132 15092 56176
rect 17068 56132 17108 56176
rect 17548 56132 17588 56344
rect 18172 56300 18212 56344
rect 19756 56333 19796 56428
rect 21510 56384 21600 56404
rect 19843 56344 19852 56384
rect 19892 56344 20140 56384
rect 20180 56344 20189 56384
rect 20899 56344 20908 56384
rect 20948 56344 21600 56384
rect 19276 56300 19316 56309
rect 18172 56260 18211 56300
rect 18251 56260 18260 56300
rect 18307 56260 18316 56300
rect 18356 56260 18365 56300
rect 18499 56260 18508 56300
rect 18548 56260 18796 56300
rect 18836 56260 18845 56300
rect 19171 56260 19180 56300
rect 19220 56260 19276 56300
rect 19316 56260 19351 56300
rect 21510 56324 21600 56344
rect 19756 56284 19796 56293
rect 18316 56216 18356 56260
rect 19276 56251 19316 56260
rect 18211 56176 18220 56216
rect 18260 56176 18356 56216
rect 20371 56176 20380 56216
rect 20420 56176 21004 56216
rect 21044 56176 21053 56216
rect 15043 56092 15052 56132
rect 15092 56092 15101 56132
rect 17059 56092 17068 56132
rect 17108 56092 17117 56132
rect 17548 56092 19948 56132
rect 19988 56092 19997 56132
rect 6172 56008 10100 56048
rect 4919 55924 4928 55964
rect 4968 55924 5010 55964
rect 5050 55924 5092 55964
rect 5132 55924 5174 55964
rect 5214 55924 5256 55964
rect 5296 55924 5305 55964
rect 20039 55924 20048 55964
rect 20088 55924 20130 55964
rect 20170 55924 20212 55964
rect 20252 55924 20294 55964
rect 20334 55924 20376 55964
rect 20416 55924 20425 55964
rect 0 55880 90 55900
rect 21510 55880 21600 55900
rect 0 55840 748 55880
rect 788 55840 797 55880
rect 4195 55840 4204 55880
rect 4244 55840 4492 55880
rect 4532 55840 5492 55880
rect 9283 55840 9292 55880
rect 9332 55840 10868 55880
rect 15331 55840 15340 55880
rect 15380 55840 17204 55880
rect 19651 55840 19660 55880
rect 19700 55840 21600 55880
rect 0 55820 90 55840
rect 5452 55796 5492 55840
rect 2275 55756 2284 55796
rect 2324 55756 3092 55796
rect 3283 55756 3292 55796
rect 3332 55756 3436 55796
rect 3476 55756 3485 55796
rect 5225 55756 5356 55796
rect 5396 55756 5405 55796
rect 5452 55756 5500 55796
rect 5540 55756 5549 55796
rect 5644 55756 6316 55796
rect 6356 55756 6892 55796
rect 6932 55756 6941 55796
rect 8995 55756 9004 55796
rect 9044 55756 9580 55796
rect 9620 55756 9629 55796
rect 2659 55672 2668 55712
rect 2708 55672 2860 55712
rect 2900 55672 2909 55712
rect 1411 55588 1420 55628
rect 1460 55588 1996 55628
rect 2036 55588 2045 55628
rect 2537 55588 2572 55628
rect 2612 55619 2708 55628
rect 2612 55588 2668 55619
rect 2668 55570 2708 55579
rect 0 55544 90 55564
rect 3052 55544 3092 55756
rect 5644 55712 5684 55756
rect 3916 55672 5684 55712
rect 5836 55672 6412 55712
rect 6452 55672 7660 55712
rect 7700 55672 7709 55712
rect 8035 55672 8044 55712
rect 8084 55672 8093 55712
rect 8524 55672 8908 55712
rect 8948 55672 10156 55712
rect 10196 55672 10205 55712
rect 3916 55628 3956 55672
rect 3907 55588 3916 55628
rect 3956 55588 3965 55628
rect 5164 55619 5204 55628
rect 0 55504 1420 55544
rect 1460 55504 1469 55544
rect 3043 55504 3052 55544
rect 3092 55504 3101 55544
rect 3619 55504 3628 55544
rect 3668 55504 3677 55544
rect 0 55484 90 55504
rect 2764 55420 3388 55460
rect 3428 55420 3437 55460
rect 2764 55376 2804 55420
rect 2755 55336 2764 55376
rect 2804 55336 2813 55376
rect 3628 55292 3668 55504
rect 5164 55460 5204 55579
rect 5836 55544 5876 55672
rect 8044 55628 8084 55672
rect 8524 55628 8564 55672
rect 6569 55588 6604 55628
rect 6644 55588 6700 55628
rect 6740 55588 6749 55628
rect 7852 55619 7892 55628
rect 8044 55588 8419 55628
rect 8459 55588 8468 55628
rect 8515 55588 8524 55628
rect 8564 55588 8573 55628
rect 8873 55588 8908 55628
rect 8948 55588 9004 55628
rect 9044 55588 9053 55628
rect 9484 55619 9676 55628
rect 7852 55544 7892 55579
rect 9524 55588 9676 55619
rect 9716 55588 9725 55628
rect 9833 55588 9964 55628
rect 10004 55588 10013 55628
rect 10828 55619 10868 55840
rect 17164 55796 17204 55840
rect 21510 55820 21600 55840
rect 17059 55756 17068 55796
rect 17108 55756 17117 55796
rect 17164 55756 17212 55796
rect 17252 55756 17261 55796
rect 17068 55712 17108 55756
rect 15043 55672 15052 55712
rect 15092 55672 15380 55712
rect 17068 55672 19892 55712
rect 15340 55628 15380 55672
rect 9484 55570 9524 55579
rect 9964 55570 10004 55579
rect 11945 55588 12076 55628
rect 12116 55588 12748 55628
rect 12788 55588 12797 55628
rect 13577 55588 13612 55628
rect 13652 55588 13708 55628
rect 13748 55588 13757 55628
rect 14179 55588 14188 55628
rect 14228 55619 14900 55628
rect 14228 55588 14860 55619
rect 10828 55570 10868 55579
rect 15322 55588 15331 55628
rect 15371 55588 15380 55628
rect 15427 55588 15436 55628
rect 15476 55588 15607 55628
rect 15689 55588 15820 55628
rect 15860 55588 15869 55628
rect 16291 55588 16300 55628
rect 16340 55619 16471 55628
rect 16340 55588 16396 55619
rect 14860 55570 14900 55579
rect 16436 55588 16471 55619
rect 16745 55588 16876 55628
rect 16916 55588 16925 55628
rect 17993 55588 18028 55628
rect 18068 55588 18124 55628
rect 18164 55588 18173 55628
rect 18307 55588 18316 55628
rect 18356 55619 19316 55628
rect 18356 55588 19276 55619
rect 16396 55570 16436 55579
rect 16876 55570 16916 55579
rect 19276 55570 19316 55579
rect 19852 55544 19892 55672
rect 5731 55504 5740 55544
rect 5780 55504 5876 55544
rect 5923 55504 5932 55544
rect 5972 55504 6508 55544
rect 6548 55504 6557 55544
rect 7852 55504 8044 55544
rect 8084 55504 8093 55544
rect 8803 55504 8812 55544
rect 8852 55504 9004 55544
rect 9044 55504 9053 55544
rect 12137 55504 12268 55544
rect 12308 55504 12317 55544
rect 15881 55504 15916 55544
rect 15956 55504 16012 55544
rect 16052 55504 16061 55544
rect 17155 55504 17164 55544
rect 17204 55504 17452 55544
rect 17492 55504 17501 55544
rect 17635 55504 17644 55544
rect 17684 55504 17693 55544
rect 19625 55504 19660 55544
rect 19700 55504 19756 55544
rect 19796 55504 19805 55544
rect 19852 55504 20140 55544
rect 20180 55504 20189 55544
rect 17644 55460 17684 55504
rect 5164 55420 14092 55460
rect 14132 55420 14141 55460
rect 16579 55420 16588 55460
rect 16628 55420 17684 55460
rect 19987 55420 19996 55460
rect 20036 55420 20812 55460
rect 20852 55420 20861 55460
rect 21510 55376 21600 55396
rect 6163 55336 6172 55376
rect 6212 55336 6220 55376
rect 6260 55336 6343 55376
rect 7267 55336 7276 55376
rect 7316 55336 10195 55376
rect 10235 55336 10244 55376
rect 10627 55336 10636 55376
rect 10676 55336 10924 55376
rect 10964 55336 10973 55376
rect 12499 55336 12508 55376
rect 12548 55336 14860 55376
rect 14900 55336 14909 55376
rect 17875 55336 17884 55376
rect 17924 55336 19412 55376
rect 19459 55336 19468 55376
rect 19508 55336 19852 55376
rect 19892 55336 19901 55376
rect 20371 55336 20380 55376
rect 20420 55336 20908 55376
rect 20948 55336 20957 55376
rect 21004 55336 21600 55376
rect 19372 55292 19412 55336
rect 3628 55252 17068 55292
rect 17108 55252 17117 55292
rect 19372 55252 20620 55292
rect 20660 55252 20669 55292
rect 0 55208 90 55228
rect 0 55168 652 55208
rect 692 55168 701 55208
rect 3679 55168 3688 55208
rect 3728 55168 3770 55208
rect 3810 55168 3852 55208
rect 3892 55168 3934 55208
rect 3974 55168 4016 55208
rect 4056 55168 4065 55208
rect 18799 55168 18808 55208
rect 18848 55168 18890 55208
rect 18930 55168 18972 55208
rect 19012 55168 19054 55208
rect 19094 55168 19136 55208
rect 19176 55168 19185 55208
rect 0 55148 90 55168
rect 2659 55084 2668 55124
rect 2708 55084 2717 55124
rect 7756 55084 13324 55124
rect 13364 55084 13373 55124
rect 2668 54956 2708 55084
rect 2668 54916 3764 54956
rect 0 54872 90 54892
rect 3724 54872 3764 54916
rect 0 54832 1804 54872
rect 1844 54832 1853 54872
rect 2851 54832 2860 54872
rect 2900 54832 3332 54872
rect 3593 54832 3724 54872
rect 3764 54832 3773 54872
rect 4195 54832 4204 54872
rect 4244 54832 4253 54872
rect 5548 54832 7508 54872
rect 0 54812 90 54832
rect 2668 54788 2708 54797
rect 3292 54788 3332 54832
rect 3724 54788 3764 54832
rect 4204 54788 4244 54832
rect 5548 54788 5588 54832
rect 7468 54788 7508 54832
rect 7756 54788 7796 55084
rect 21004 55040 21044 55336
rect 21510 55316 21600 55336
rect 7852 55000 11788 55040
rect 11828 55000 11837 55040
rect 13289 55000 13420 55040
rect 13460 55000 13469 55040
rect 14921 55000 15052 55040
rect 15092 55000 15101 55040
rect 16649 55000 16780 55040
rect 16820 55000 16829 55040
rect 18883 55000 18892 55040
rect 18932 55000 21044 55040
rect 7852 54788 7892 55000
rect 9667 54916 9676 54956
rect 9716 54916 10292 54956
rect 12163 54916 12172 54956
rect 12212 54916 12844 54956
rect 12884 54916 17300 54956
rect 19939 54916 19948 54956
rect 19988 54916 20332 54956
rect 20372 54916 20381 54956
rect 9571 54832 9580 54872
rect 9620 54832 10060 54872
rect 10100 54832 10109 54872
rect 9100 54788 9140 54797
rect 10252 54788 10292 54916
rect 10723 54832 10732 54872
rect 10772 54832 11347 54872
rect 11387 54832 11396 54872
rect 14860 54832 16300 54872
rect 16340 54832 16628 54872
rect 10636 54788 10676 54797
rect 13228 54788 13268 54797
rect 14860 54788 14900 54832
rect 16588 54788 16628 54832
rect 17260 54788 17300 54916
rect 21510 54872 21600 54892
rect 18307 54832 18316 54872
rect 18356 54832 18432 54872
rect 20707 54832 20716 54872
rect 20756 54832 21600 54872
rect 18316 54788 18356 54832
rect 21510 54812 21600 54832
rect 20140 54788 20180 54797
rect 1411 54748 1420 54788
rect 1460 54748 2284 54788
rect 2324 54748 2333 54788
rect 2563 54748 2572 54788
rect 2612 54748 2668 54788
rect 2708 54748 2743 54788
rect 2860 54748 3052 54788
rect 3092 54748 3101 54788
rect 3148 54748 3191 54788
rect 3231 54748 3240 54788
rect 3292 54748 3532 54788
rect 3572 54748 3581 54788
rect 3706 54748 3715 54788
rect 3755 54748 3764 54788
rect 3811 54748 3820 54788
rect 3860 54748 3869 54788
rect 4003 54748 4012 54788
rect 4052 54748 4244 54788
rect 4291 54748 4300 54788
rect 4340 54748 4492 54788
rect 4532 54748 4541 54788
rect 5417 54748 5548 54788
rect 5588 54748 5597 54788
rect 6019 54748 6028 54788
rect 6068 54748 6220 54788
rect 6260 54748 6892 54788
rect 6932 54748 6941 54788
rect 7508 54748 7796 54788
rect 7843 54748 7852 54788
rect 7892 54748 7901 54788
rect 8969 54748 9004 54788
rect 9044 54748 9100 54788
rect 9187 54748 9196 54788
rect 9236 54748 9571 54788
rect 9611 54748 9620 54788
rect 9667 54748 9676 54788
rect 9716 54748 9847 54788
rect 9964 54748 10156 54788
rect 10196 54748 10205 54788
rect 10252 54748 10444 54788
rect 10484 54748 10636 54788
rect 11146 54748 11155 54788
rect 11195 54748 11308 54788
rect 11348 54748 11357 54788
rect 11779 54748 11788 54788
rect 11828 54748 11980 54788
rect 12020 54748 12029 54788
rect 13193 54748 13228 54788
rect 13268 54748 13324 54788
rect 13364 54748 13373 54788
rect 13577 54748 13612 54788
rect 13652 54748 13708 54788
rect 13748 54748 13757 54788
rect 14729 54748 14860 54788
rect 14900 54748 14909 54788
rect 15331 54748 15340 54788
rect 15380 54748 15724 54788
rect 15764 54748 15773 54788
rect 17033 54748 17068 54788
rect 17108 54748 17164 54788
rect 17204 54748 17213 54788
rect 17260 54748 18316 54788
rect 18403 54748 18412 54788
rect 18452 54748 18892 54788
rect 18932 54748 18941 54788
rect 19459 54748 19468 54788
rect 19508 54748 20140 54788
rect 2668 54739 2708 54748
rect 2860 54620 2900 54748
rect 3148 54620 3188 54748
rect 3820 54704 3860 54748
rect 5548 54739 5588 54748
rect 7468 54739 7508 54748
rect 9100 54739 9140 54748
rect 3497 54664 3619 54704
rect 3668 54664 3677 54704
rect 3820 54664 3916 54704
rect 3956 54664 3965 54704
rect 2851 54580 2860 54620
rect 2900 54580 2909 54620
rect 3043 54580 3052 54620
rect 3092 54580 3188 54620
rect 3331 54580 3340 54620
rect 3380 54580 3532 54620
rect 3572 54580 3581 54620
rect 4147 54580 4156 54620
rect 4196 54580 4204 54620
rect 4244 54580 4327 54620
rect 5731 54580 5740 54620
rect 5780 54580 5789 54620
rect 7651 54580 7660 54620
rect 7700 54580 7756 54620
rect 7796 54580 7831 54620
rect 9161 54580 9292 54620
rect 9332 54580 9341 54620
rect 0 54536 90 54556
rect 2860 54536 2900 54580
rect 0 54496 2764 54536
rect 2804 54496 2813 54536
rect 2860 54496 3916 54536
rect 3956 54496 3965 54536
rect 0 54476 90 54496
rect 4919 54412 4928 54452
rect 4968 54412 5010 54452
rect 5050 54412 5092 54452
rect 5132 54412 5174 54452
rect 5214 54412 5256 54452
rect 5296 54412 5305 54452
rect 3523 54328 3532 54368
rect 3572 54328 4052 54368
rect 1699 54244 1708 54284
rect 1748 54244 1948 54284
rect 1988 54244 1997 54284
rect 3484 54244 3820 54284
rect 3860 54244 3869 54284
rect 0 54200 90 54220
rect 0 54160 1324 54200
rect 1364 54160 1373 54200
rect 0 54140 90 54160
rect 3484 54116 3524 54244
rect 4012 54200 4052 54328
rect 3715 54160 3724 54200
rect 3764 54160 3860 54200
rect 1961 54076 2092 54116
rect 2132 54076 2141 54116
rect 2467 54076 2476 54116
rect 2516 54107 3524 54116
rect 2516 54076 3340 54107
rect 3380 54076 3524 54107
rect 3579 54076 3628 54116
rect 3668 54105 3677 54116
rect 3820 54107 3860 54160
rect 3994 54191 4052 54200
rect 3994 54151 4003 54191
rect 4043 54151 4052 54191
rect 5740 54200 5780 54580
rect 9964 54536 10004 54748
rect 10636 54739 10676 54748
rect 13228 54739 13268 54748
rect 14860 54739 14900 54748
rect 16588 54739 16628 54748
rect 18316 54739 18356 54748
rect 20140 54739 20180 54748
rect 16675 54664 16684 54704
rect 16724 54664 17260 54704
rect 17300 54664 17309 54704
rect 17260 54536 17300 54664
rect 18377 54580 18508 54620
rect 18548 54580 18557 54620
rect 8803 54496 8812 54536
rect 8852 54496 9964 54536
rect 10004 54496 10013 54536
rect 17260 54496 19084 54536
rect 19124 54496 19133 54536
rect 13603 54412 13612 54452
rect 13652 54412 17156 54452
rect 20039 54412 20048 54452
rect 20088 54412 20130 54452
rect 20170 54412 20212 54452
rect 20252 54412 20294 54452
rect 20334 54412 20376 54452
rect 20416 54412 20425 54452
rect 14755 54328 14764 54368
rect 14804 54328 17060 54368
rect 17020 54284 17060 54328
rect 6211 54244 6220 54284
rect 6260 54244 6356 54284
rect 7267 54244 7276 54284
rect 7316 54244 7325 54284
rect 7817 54244 7948 54284
rect 7988 54244 7997 54284
rect 8515 54244 8524 54284
rect 8564 54244 9004 54284
rect 9044 54244 11060 54284
rect 11299 54244 11308 54284
rect 11348 54244 11479 54284
rect 12809 54244 12892 54284
rect 12932 54244 12940 54284
rect 12980 54244 12989 54284
rect 14947 54244 14956 54284
rect 14996 54244 15284 54284
rect 17011 54244 17020 54284
rect 17060 54244 17069 54284
rect 5740 54160 6260 54200
rect 3994 54150 4052 54151
rect 6220 54116 6260 54160
rect 6316 54116 6356 54244
rect 7276 54200 7316 54244
rect 7276 54160 7852 54200
rect 7892 54160 7901 54200
rect 9571 54160 9580 54200
rect 9620 54160 9908 54200
rect 3668 54076 3699 54105
rect 3340 54058 3380 54067
rect 3628 54065 3699 54076
rect 3739 54065 3748 54105
rect 4090 54076 4099 54116
rect 4139 54076 4148 54116
rect 4195 54076 4204 54116
rect 4273 54076 4375 54116
rect 4483 54076 4492 54116
rect 4532 54076 4663 54116
rect 5609 54076 5740 54116
rect 5780 54076 5789 54116
rect 6202 54076 6211 54116
rect 6251 54076 6260 54116
rect 6307 54076 6316 54116
rect 6356 54076 6365 54116
rect 6691 54076 6700 54116
rect 6740 54076 6749 54116
rect 7171 54076 7180 54116
rect 7220 54076 7229 54116
rect 7276 54107 7316 54160
rect 9868 54116 9908 54160
rect 11020 54116 11060 54244
rect 11779 54160 11788 54200
rect 11828 54160 12980 54200
rect 14851 54160 14860 54200
rect 14900 54160 15188 54200
rect 12940 54116 12980 54160
rect 15148 54116 15188 54160
rect 15244 54116 15284 54244
rect 17116 54200 17156 54412
rect 21510 54368 21600 54388
rect 17932 54328 18892 54368
rect 18932 54328 18941 54368
rect 20611 54328 20620 54368
rect 20660 54328 21600 54368
rect 17932 54284 17972 54328
rect 21510 54308 21600 54328
rect 17683 54244 17692 54284
rect 17732 54244 17972 54284
rect 18028 54244 20044 54284
rect 20084 54244 20093 54284
rect 17116 54160 17788 54200
rect 17828 54160 17837 54200
rect 3820 54058 3860 54067
rect 4108 54032 4148 54076
rect 5740 54058 5780 54067
rect 1411 53992 1420 54032
rect 1460 53992 1469 54032
rect 1577 53992 1708 54032
rect 1748 53992 1757 54032
rect 3907 53992 3916 54032
rect 3956 53992 4148 54032
rect 0 53864 90 53884
rect 0 53824 460 53864
rect 500 53824 509 53864
rect 643 53824 652 53864
rect 692 53824 1180 53864
rect 1220 53824 1229 53864
rect 0 53804 90 53824
rect 1420 53780 1460 53992
rect 6700 53948 6740 54076
rect 7180 54032 7220 54076
rect 7625 54076 7756 54116
rect 7796 54076 7805 54116
rect 9257 54076 9292 54116
rect 9332 54076 9379 54116
rect 9419 54076 9437 54116
rect 9480 54076 9489 54116
rect 9529 54076 9676 54116
rect 9716 54076 9725 54116
rect 9859 54076 9868 54116
rect 9908 54076 9917 54116
rect 10313 54076 10444 54116
rect 10484 54076 10493 54116
rect 10793 54076 10924 54116
rect 10964 54076 10973 54116
rect 11020 54107 11540 54116
rect 11020 54076 11500 54107
rect 7276 54058 7316 54067
rect 7756 54058 7796 54067
rect 9484 54032 9524 54076
rect 10444 54058 10484 54067
rect 10924 54058 10964 54067
rect 12739 54076 12748 54116
rect 12788 54076 12797 54116
rect 12940 54076 13420 54116
rect 13460 54076 13469 54116
rect 14083 54076 14092 54116
rect 14132 54107 14708 54116
rect 14132 54076 14668 54107
rect 11500 54058 11540 54067
rect 6787 53992 6796 54032
rect 6836 53992 7220 54032
rect 8899 53992 8908 54032
rect 8948 53992 9524 54032
rect 9833 53992 9964 54032
rect 10004 53992 10013 54032
rect 12748 53948 12788 54076
rect 15130 54076 15139 54116
rect 15179 54076 15188 54116
rect 15235 54076 15244 54116
rect 15284 54076 15415 54116
rect 15497 54076 15628 54116
rect 15668 54076 16012 54116
rect 16052 54076 16061 54116
rect 16204 54107 16588 54116
rect 14668 54058 14708 54067
rect 16244 54076 16588 54107
rect 16628 54076 16637 54116
rect 16684 54107 16724 54116
rect 16204 54058 16244 54067
rect 17923 54076 17932 54116
rect 17972 54076 17981 54116
rect 13123 53992 13132 54032
rect 13172 53992 13324 54032
rect 13364 53992 13373 54032
rect 15689 53992 15724 54032
rect 15764 53992 15820 54032
rect 15860 53992 15869 54032
rect 3523 53908 3532 53948
rect 3572 53908 4204 53948
rect 4244 53908 4253 53948
rect 5923 53908 5932 53948
rect 5972 53908 7180 53948
rect 7220 53908 7229 53948
rect 8803 53908 8812 53948
rect 8852 53908 15724 53948
rect 15764 53908 15773 53948
rect 3593 53824 3715 53864
rect 3764 53824 3773 53864
rect 5923 53824 5932 53864
rect 5972 53824 6604 53864
rect 6644 53824 6653 53864
rect 10051 53824 10060 53864
rect 10100 53824 10348 53864
rect 10388 53824 10397 53864
rect 10627 53824 10636 53864
rect 10676 53824 11155 53864
rect 11195 53824 11500 53864
rect 11540 53824 11549 53864
rect 1420 53740 14708 53780
rect 1891 53656 1900 53696
rect 1940 53656 3572 53696
rect 3679 53656 3688 53696
rect 3728 53656 3770 53696
rect 3810 53656 3852 53696
rect 3892 53656 3934 53696
rect 3974 53656 4016 53696
rect 4056 53656 4065 53696
rect 5731 53656 5740 53696
rect 5780 53656 6988 53696
rect 7028 53656 12652 53696
rect 12692 53656 12701 53696
rect 3532 53612 3572 53656
rect 1420 53572 3476 53612
rect 3532 53572 5932 53612
rect 5972 53572 5981 53612
rect 6028 53572 9964 53612
rect 10004 53572 10013 53612
rect 10060 53572 14572 53612
rect 14612 53572 14621 53612
rect 0 53528 90 53548
rect 0 53488 556 53528
rect 596 53488 605 53528
rect 0 53468 90 53488
rect 1420 53360 1460 53572
rect 3436 53528 3476 53572
rect 6028 53528 6068 53572
rect 10060 53528 10100 53572
rect 2057 53488 2140 53528
rect 2180 53488 2188 53528
rect 2228 53488 2237 53528
rect 3436 53488 6068 53528
rect 8458 53488 8467 53528
rect 8507 53488 10100 53528
rect 10483 53488 10492 53528
rect 10532 53488 10676 53528
rect 12403 53488 12412 53528
rect 12452 53488 12748 53528
rect 12788 53488 14380 53528
rect 14420 53488 14429 53528
rect 10636 53444 10676 53488
rect 14668 53444 14708 53740
rect 16684 53528 16724 54067
rect 17932 54032 17972 54076
rect 18028 54032 18068 54244
rect 18316 54160 18508 54200
rect 18548 54160 18557 54200
rect 18316 54116 18356 54160
rect 18298 54076 18307 54116
rect 18347 54076 18356 54116
rect 18403 54076 18412 54116
rect 18452 54076 18604 54116
rect 18644 54076 18653 54116
rect 18787 54076 18796 54116
rect 18836 54076 18967 54116
rect 19075 54076 19084 54116
rect 19124 54107 19468 54116
rect 19124 54076 19372 54107
rect 19412 54076 19468 54107
rect 19508 54076 19572 54116
rect 19721 54076 19852 54116
rect 19892 54076 19901 54116
rect 19372 54058 19412 54067
rect 19852 54058 19892 54067
rect 16906 53992 16915 54032
rect 16955 53992 17260 54032
rect 17300 53992 17309 54032
rect 17443 53992 17452 54032
rect 17492 53992 17972 54032
rect 18019 53992 18028 54032
rect 18068 53992 18077 54032
rect 18761 53992 18892 54032
rect 18932 53992 18941 54032
rect 21510 53864 21600 53884
rect 18700 53824 18796 53864
rect 18836 53824 18845 53864
rect 20995 53824 21004 53864
rect 21044 53824 21600 53864
rect 18700 53612 18740 53824
rect 21510 53804 21600 53824
rect 18799 53656 18808 53696
rect 18848 53656 18890 53696
rect 18930 53656 18972 53696
rect 19012 53656 19054 53696
rect 19094 53656 19136 53696
rect 19176 53656 19185 53696
rect 17155 53572 17164 53612
rect 17204 53572 19028 53612
rect 15235 53488 15244 53528
rect 15284 53488 16724 53528
rect 16780 53488 17788 53528
rect 17828 53488 17837 53528
rect 16780 53444 16820 53488
rect 3043 53404 3052 53444
rect 3092 53404 3188 53444
rect 3235 53404 3244 53444
rect 3284 53404 3293 53444
rect 3340 53404 6892 53444
rect 6932 53404 6941 53444
rect 7267 53404 7276 53444
rect 7316 53404 8428 53444
rect 8468 53404 8477 53444
rect 9929 53404 10060 53444
rect 10100 53404 10109 53444
rect 10156 53404 10444 53444
rect 10484 53404 10493 53444
rect 10627 53404 10636 53444
rect 10676 53404 10685 53444
rect 10915 53404 10924 53444
rect 10964 53404 10973 53444
rect 11779 53404 11788 53444
rect 11828 53404 12508 53444
rect 12548 53404 12557 53444
rect 14668 53404 16820 53444
rect 17299 53404 17308 53444
rect 17348 53404 18068 53444
rect 3148 53360 3188 53404
rect 547 53320 556 53360
rect 596 53320 1180 53360
rect 1220 53320 1229 53360
rect 1411 53320 1420 53360
rect 1460 53320 1469 53360
rect 1891 53320 1900 53360
rect 1940 53320 2092 53360
rect 2132 53320 3092 53360
rect 3139 53320 3148 53360
rect 3188 53320 3197 53360
rect 2650 53236 2659 53276
rect 2699 53236 2708 53276
rect 2755 53236 2764 53276
rect 2804 53236 2900 53276
rect 0 53192 90 53212
rect 0 53152 1324 53192
rect 1364 53152 1373 53192
rect 0 53132 90 53152
rect 0 52856 90 52876
rect 0 52816 652 52856
rect 692 52816 701 52856
rect 0 52796 90 52816
rect 2668 52772 2708 53236
rect 2860 53192 2900 53236
rect 3052 53192 3092 53320
rect 3244 53276 3284 53404
rect 3235 53236 3244 53276
rect 3284 53236 3293 53276
rect 3340 53192 3380 53404
rect 7049 53320 7180 53360
rect 7220 53320 7229 53360
rect 8140 53320 9620 53360
rect 3724 53276 3764 53285
rect 6124 53276 6164 53285
rect 7756 53276 7796 53285
rect 8140 53276 8180 53320
rect 9580 53276 9620 53320
rect 10156 53276 10196 53404
rect 10924 53360 10964 53404
rect 18028 53360 18068 53404
rect 18988 53360 19028 53572
rect 21510 53360 21600 53380
rect 10243 53320 10252 53360
rect 10292 53320 10348 53360
rect 10388 53320 10423 53360
rect 10579 53320 10588 53360
rect 10628 53320 10964 53360
rect 12163 53320 12172 53360
rect 12212 53320 12460 53360
rect 12500 53320 12509 53360
rect 12739 53320 12748 53360
rect 12788 53320 13324 53360
rect 13364 53320 13373 53360
rect 15881 53320 16012 53360
rect 16052 53320 16061 53360
rect 16963 53320 16972 53360
rect 17012 53320 17300 53360
rect 17395 53320 17404 53360
rect 17444 53320 17452 53360
rect 17492 53320 17575 53360
rect 17635 53320 17644 53360
rect 17684 53320 17693 53360
rect 18019 53320 18028 53360
rect 18068 53320 18077 53360
rect 18499 53320 18508 53360
rect 18548 53320 18932 53360
rect 18979 53320 18988 53360
rect 19028 53320 19037 53360
rect 20803 53320 20812 53360
rect 20852 53320 21600 53360
rect 15052 53276 15092 53285
rect 16588 53276 16628 53285
rect 17260 53276 17300 53320
rect 17644 53276 17684 53320
rect 18892 53276 18932 53320
rect 21510 53300 21600 53320
rect 19564 53276 19604 53285
rect 3764 53236 4012 53276
rect 4052 53236 4061 53276
rect 4195 53236 4204 53276
rect 4252 53236 4375 53276
rect 4867 53236 4876 53276
rect 4916 53236 4925 53276
rect 5539 53236 5548 53276
rect 5588 53236 5740 53276
rect 5780 53236 6124 53276
rect 6539 53236 6604 53276
rect 6644 53236 6670 53276
rect 6710 53236 6719 53276
rect 6787 53236 6796 53276
rect 6836 53236 6845 53276
rect 7145 53236 7276 53276
rect 7316 53236 7325 53276
rect 7721 53236 7756 53276
rect 7796 53236 7852 53276
rect 7892 53236 8180 53276
rect 8227 53236 8236 53276
rect 8284 53236 8407 53276
rect 8707 53236 8716 53276
rect 8756 53236 8765 53276
rect 8995 53236 9004 53276
rect 9044 53236 9388 53276
rect 9428 53236 9484 53276
rect 9524 53236 9533 53276
rect 9580 53236 9643 53276
rect 9683 53236 9692 53276
rect 9754 53236 9763 53276
rect 9803 53236 10196 53276
rect 10723 53236 10732 53276
rect 10772 53236 12596 53276
rect 12835 53236 12844 53276
rect 12884 53236 13804 53276
rect 13844 53236 13853 53276
rect 14371 53236 14380 53276
rect 14420 53236 15052 53276
rect 15514 53236 15523 53276
rect 15563 53236 15572 53276
rect 15619 53236 15628 53276
rect 15668 53236 15799 53276
rect 16073 53236 16108 53276
rect 16148 53236 16204 53276
rect 16244 53236 16253 53276
rect 16628 53236 16684 53276
rect 16724 53236 16759 53276
rect 17098 53236 17107 53276
rect 17147 53236 17204 53276
rect 17260 53236 17684 53276
rect 18490 53236 18499 53276
rect 18539 53236 18548 53276
rect 18595 53236 18604 53276
rect 18644 53236 18775 53276
rect 18892 53236 19084 53276
rect 19124 53236 19133 53276
rect 19363 53236 19372 53276
rect 19412 53236 19564 53276
rect 19939 53236 19948 53276
rect 19988 53236 20052 53276
rect 20092 53236 20119 53276
rect 3724 53227 3764 53236
rect 2851 53152 2860 53192
rect 2900 53152 2909 53192
rect 3052 53152 3380 53192
rect 4876 53192 4916 53236
rect 6124 53227 6164 53236
rect 6796 53192 6836 53236
rect 7756 53227 7796 53236
rect 8716 53192 8756 53236
rect 10732 53192 10772 53236
rect 4876 53152 5836 53192
rect 5876 53152 5885 53192
rect 6220 53152 6836 53192
rect 7852 53152 8756 53192
rect 9667 53152 9676 53192
rect 9716 53152 10772 53192
rect 6220 53108 6260 53152
rect 4265 53068 4396 53108
rect 4436 53068 4445 53108
rect 6019 53068 6028 53108
rect 6068 53068 6260 53108
rect 6307 53068 6316 53108
rect 6356 53068 6604 53108
rect 6644 53068 6653 53108
rect 7852 53024 7892 53152
rect 8794 53068 8803 53108
rect 8843 53068 9964 53108
rect 10004 53068 10013 53108
rect 5347 52984 5356 53024
rect 5396 52984 7892 53024
rect 9283 52984 9292 53024
rect 9332 52984 10732 53024
rect 10772 52984 10781 53024
rect 4919 52900 4928 52940
rect 4968 52900 5010 52940
rect 5050 52900 5092 52940
rect 5132 52900 5174 52940
rect 5214 52900 5256 52940
rect 5296 52900 5305 52940
rect 9475 52816 9484 52856
rect 9524 52816 10964 52856
rect 10924 52772 10964 52816
rect 12556 52772 12596 53236
rect 15052 53227 15092 53236
rect 15532 52772 15572 53236
rect 16588 53227 16628 53236
rect 17164 52772 17204 53236
rect 18508 52772 18548 53236
rect 19564 53227 19604 53236
rect 19651 53068 19660 53108
rect 19700 53068 20236 53108
rect 20276 53068 20285 53108
rect 20039 52900 20048 52940
rect 20088 52900 20130 52940
rect 20170 52900 20212 52940
rect 20252 52900 20294 52940
rect 20334 52900 20376 52940
rect 20416 52900 20425 52940
rect 21510 52856 21600 52876
rect 20899 52816 20908 52856
rect 20948 52816 21600 52856
rect 21510 52796 21600 52816
rect 2659 52732 2668 52772
rect 2708 52732 2717 52772
rect 4876 52732 5740 52772
rect 5780 52732 5789 52772
rect 6595 52732 6604 52772
rect 6644 52732 6892 52772
rect 6932 52732 6941 52772
rect 9859 52732 9868 52772
rect 9908 52732 10100 52772
rect 10627 52732 10636 52772
rect 10676 52732 10732 52772
rect 10772 52732 10807 52772
rect 10915 52732 10924 52772
rect 10964 52732 10973 52772
rect 12547 52732 12556 52772
rect 12596 52732 12605 52772
rect 12835 52732 12844 52772
rect 12884 52732 15476 52772
rect 15532 52732 15628 52772
rect 15668 52732 15677 52772
rect 17164 52732 17260 52772
rect 17300 52732 17309 52772
rect 18508 52732 18892 52772
rect 18932 52732 18941 52772
rect 19027 52732 19036 52772
rect 19076 52732 19084 52772
rect 19124 52732 19207 52772
rect 1219 52564 1228 52604
rect 1268 52564 1708 52604
rect 1748 52564 1757 52604
rect 2345 52564 2476 52604
rect 2516 52564 2525 52604
rect 3619 52564 3628 52604
rect 3668 52564 4108 52604
rect 4148 52564 4157 52604
rect 4876 52595 4916 52732
rect 10060 52688 10100 52732
rect 5059 52648 5068 52688
rect 5108 52648 5117 52688
rect 5548 52648 7372 52688
rect 7412 52648 7421 52688
rect 8140 52648 9484 52688
rect 9524 52648 9533 52688
rect 10060 52648 10540 52688
rect 10580 52648 10589 52688
rect 11116 52648 12788 52688
rect 13699 52648 13708 52688
rect 13748 52648 14228 52688
rect 2476 52546 2516 52555
rect 5068 52604 5108 52648
rect 5548 52604 5588 52648
rect 5068 52564 5347 52604
rect 5387 52564 5396 52604
rect 5443 52564 5452 52604
rect 5492 52564 5548 52604
rect 5588 52564 5623 52604
rect 5827 52564 5836 52604
rect 5876 52564 6028 52604
rect 6068 52564 6077 52604
rect 6307 52564 6316 52604
rect 6356 52595 6487 52604
rect 6356 52564 6412 52595
rect 4876 52546 4916 52555
rect 6452 52564 6487 52595
rect 6761 52564 6892 52604
rect 6932 52564 6941 52604
rect 6412 52546 6452 52555
rect 6892 52546 6932 52555
rect 0 52520 90 52540
rect 7372 52520 7412 52648
rect 8140 52604 8180 52648
rect 8122 52564 8131 52604
rect 8171 52564 8180 52604
rect 8227 52564 8236 52604
rect 8276 52564 8285 52604
rect 8332 52564 8620 52604
rect 8660 52564 8669 52604
rect 9196 52595 9292 52604
rect 8236 52520 8276 52564
rect 0 52480 652 52520
rect 692 52480 701 52520
rect 3043 52480 3052 52520
rect 3092 52480 4684 52520
rect 4724 52480 4733 52520
rect 5801 52480 5932 52520
rect 5972 52480 5981 52520
rect 7372 52480 8276 52520
rect 0 52460 90 52480
rect 5932 52436 5972 52480
rect 8332 52436 8372 52564
rect 9236 52564 9292 52595
rect 9332 52564 9367 52604
rect 9545 52564 9676 52604
rect 9716 52564 9725 52604
rect 9955 52564 9964 52604
rect 10004 52564 10007 52604
rect 10047 52564 10135 52604
rect 10243 52564 10252 52604
rect 10292 52564 10301 52604
rect 10409 52564 10444 52604
rect 10484 52564 10540 52604
rect 10580 52564 10589 52604
rect 10714 52564 10723 52604
rect 10763 52564 10772 52604
rect 9196 52546 9236 52555
rect 9676 52546 9716 52555
rect 8419 52480 8428 52520
rect 8468 52480 8716 52520
rect 8756 52480 8765 52520
rect 10138 52480 10147 52520
rect 10187 52480 10196 52520
rect 10156 52436 10196 52480
rect 5932 52396 6508 52436
rect 6548 52396 8372 52436
rect 9955 52396 9964 52436
rect 10004 52396 10196 52436
rect 10252 52436 10292 52564
rect 10732 52520 10772 52564
rect 11116 52595 11156 52648
rect 12748 52604 12788 52648
rect 14188 52604 14228 52648
rect 12355 52564 12364 52604
rect 12404 52564 12413 52604
rect 12617 52564 12748 52604
rect 12788 52564 12797 52604
rect 13987 52564 13996 52604
rect 14036 52564 14045 52604
rect 14179 52564 14188 52604
rect 14228 52564 14359 52604
rect 15436 52595 15476 52732
rect 17059 52648 17068 52688
rect 17108 52648 19420 52688
rect 19460 52648 19469 52688
rect 11116 52546 11156 52555
rect 10339 52480 10348 52520
rect 10388 52480 10519 52520
rect 10627 52480 10636 52520
rect 10676 52480 10772 52520
rect 10252 52396 10924 52436
rect 10964 52396 10973 52436
rect 172 52312 2812 52352
rect 2852 52312 2861 52352
rect 7114 52312 7123 52352
rect 7163 52312 10004 52352
rect 0 52184 90 52204
rect 172 52184 212 52312
rect 9964 52268 10004 52312
rect 9964 52228 10580 52268
rect 0 52144 212 52184
rect 3679 52144 3688 52184
rect 3728 52144 3770 52184
rect 3810 52144 3852 52184
rect 3892 52144 3934 52184
rect 3974 52144 4016 52184
rect 4056 52144 4065 52184
rect 0 52124 90 52144
rect 10540 52100 10580 52228
rect 12364 52184 12404 52564
rect 12748 52546 12788 52555
rect 13996 52352 14036 52564
rect 15689 52564 15724 52604
rect 15764 52564 15820 52604
rect 15860 52564 15869 52604
rect 17068 52595 17108 52604
rect 15436 52520 15476 52555
rect 17251 52564 17260 52604
rect 17300 52564 17452 52604
rect 17492 52564 17501 52604
rect 18700 52595 19948 52604
rect 17068 52520 17108 52555
rect 18740 52564 19948 52595
rect 19988 52564 19997 52604
rect 18700 52520 18740 52555
rect 15436 52480 18740 52520
rect 19267 52480 19276 52520
rect 19316 52480 19325 52520
rect 19529 52480 19660 52520
rect 19700 52480 19709 52520
rect 20009 52480 20140 52520
rect 20180 52480 20189 52520
rect 19276 52436 19316 52480
rect 17443 52396 17452 52436
rect 17492 52396 17836 52436
rect 17876 52396 19316 52436
rect 19747 52396 19756 52436
rect 19796 52396 20564 52436
rect 20524 52352 20564 52396
rect 21510 52352 21600 52372
rect 13996 52312 17644 52352
rect 17684 52312 18412 52352
rect 18452 52312 18461 52352
rect 20297 52312 20380 52352
rect 20420 52312 20428 52352
rect 20468 52312 20477 52352
rect 20524 52312 21600 52352
rect 21510 52292 21600 52312
rect 12364 52144 16396 52184
rect 16436 52144 17260 52184
rect 17300 52144 17309 52184
rect 18799 52144 18808 52184
rect 18848 52144 18890 52184
rect 18930 52144 18972 52184
rect 19012 52144 19054 52184
rect 19094 52144 19136 52184
rect 19176 52144 19185 52184
rect 10348 52060 10444 52100
rect 10484 52060 10493 52100
rect 10540 52060 14092 52100
rect 14132 52060 14141 52100
rect 10348 52016 10388 52060
rect 6019 51976 6028 52016
rect 6068 51976 6164 52016
rect 7843 51976 7852 52016
rect 7892 51976 8236 52016
rect 8276 51976 8285 52016
rect 8707 51976 8716 52016
rect 8756 51976 10292 52016
rect 10339 51976 10348 52016
rect 10388 51976 10397 52016
rect 10505 51976 10540 52016
rect 10580 51976 10636 52016
rect 10676 51976 10685 52016
rect 10793 51976 10924 52016
rect 10964 51976 10973 52016
rect 2851 51892 2860 51932
rect 2900 51892 4052 51932
rect 0 51848 90 51868
rect 4012 51848 4052 51892
rect 4300 51892 5548 51932
rect 5588 51892 6068 51932
rect 0 51808 556 51848
rect 596 51808 605 51848
rect 1411 51808 1420 51848
rect 1460 51808 1469 51848
rect 1673 51808 1804 51848
rect 1844 51808 1853 51848
rect 2083 51808 2092 51848
rect 2132 51808 2476 51848
rect 2516 51808 2572 51848
rect 2612 51808 2621 51848
rect 2668 51808 2716 51848
rect 2756 51808 2765 51848
rect 4003 51808 4012 51848
rect 4052 51808 4061 51848
rect 0 51788 90 51808
rect 1420 51680 1460 51808
rect 2668 51680 2708 51808
rect 3532 51764 3572 51773
rect 4300 51764 4340 51892
rect 4387 51808 4396 51848
rect 4436 51808 5068 51848
rect 5108 51808 5117 51848
rect 6028 51764 6068 51892
rect 6124 51848 6164 51976
rect 10252 51932 10292 51976
rect 7948 51892 8180 51932
rect 7948 51848 7988 51892
rect 6124 51808 6412 51848
rect 6452 51808 6461 51848
rect 7075 51808 7084 51848
rect 7124 51808 7988 51848
rect 8140 51848 8180 51892
rect 9868 51892 9964 51932
rect 10004 51892 10013 51932
rect 10252 51892 12844 51932
rect 12884 51892 12893 51932
rect 16012 51892 16820 51932
rect 17251 51892 17260 51932
rect 17300 51892 18452 51932
rect 9868 51848 9908 51892
rect 16012 51848 16052 51892
rect 8140 51808 9332 51848
rect 9667 51808 9676 51848
rect 9716 51808 9812 51848
rect 9859 51808 9868 51848
rect 9908 51808 9917 51848
rect 10492 51808 10540 51848
rect 10580 51808 10589 51848
rect 11299 51808 11308 51848
rect 11348 51808 12556 51848
rect 12596 51808 12605 51848
rect 14860 51808 16052 51848
rect 16780 51848 16820 51892
rect 16780 51808 18316 51848
rect 18356 51808 18365 51848
rect 6988 51764 7028 51773
rect 8044 51764 8084 51773
rect 9292 51764 9332 51808
rect 9772 51764 9812 51808
rect 10492 51764 10532 51808
rect 11116 51764 11156 51773
rect 13420 51764 13460 51773
rect 14860 51764 14900 51808
rect 16108 51764 16148 51773
rect 16684 51764 16724 51773
rect 18412 51764 18452 51892
rect 21510 51848 21600 51868
rect 20009 51808 20140 51848
rect 20180 51808 20189 51848
rect 20419 51808 20428 51848
rect 20468 51808 21600 51848
rect 21510 51788 21600 51808
rect 19468 51764 19508 51773
rect 3034 51724 3043 51764
rect 3083 51724 3092 51764
rect 1420 51640 2180 51680
rect 2249 51640 2332 51680
rect 2372 51640 2380 51680
rect 2420 51640 2429 51680
rect 2572 51640 2708 51680
rect 3052 51680 3092 51724
rect 3619 51724 3628 51764
rect 3668 51724 4108 51764
rect 4148 51724 4157 51764
rect 4300 51724 4492 51764
rect 4532 51724 4541 51764
rect 4601 51724 4610 51764
rect 4650 51724 5780 51764
rect 5914 51724 5923 51764
rect 5963 51724 5972 51764
rect 6019 51724 6028 51764
rect 6068 51724 6077 51764
rect 6377 51724 6508 51764
rect 6548 51724 6557 51764
rect 7471 51724 7480 51764
rect 7520 51724 7529 51764
rect 7939 51724 7948 51764
rect 7988 51724 8044 51764
rect 8084 51724 8119 51764
rect 9283 51724 9292 51764
rect 9332 51724 9341 51764
rect 9396 51724 9484 51764
rect 9524 51724 9527 51764
rect 9567 51724 9576 51764
rect 9658 51724 9667 51764
rect 9707 51724 9716 51764
rect 9763 51724 9772 51764
rect 9812 51724 9821 51764
rect 9929 51724 10051 51764
rect 10100 51724 10109 51764
rect 10228 51724 10348 51764
rect 10399 51724 10408 51764
rect 10492 51724 10540 51764
rect 10580 51724 10589 51764
rect 10720 51724 10729 51764
rect 10769 51724 10964 51764
rect 3052 51640 3476 51680
rect 547 51556 556 51596
rect 596 51556 1180 51596
rect 1220 51556 1229 51596
rect 1324 51556 1564 51596
rect 1604 51556 1613 51596
rect 0 51512 90 51532
rect 1324 51512 1364 51556
rect 0 51472 1364 51512
rect 0 51452 90 51472
rect 643 51220 652 51260
rect 692 51220 1180 51260
rect 1220 51220 1229 51260
rect 1315 51220 1324 51260
rect 1364 51220 1564 51260
rect 1604 51220 1613 51260
rect 0 51176 90 51196
rect 0 51136 556 51176
rect 596 51136 605 51176
rect 0 51116 90 51136
rect 1411 50968 1420 51008
rect 1460 50968 1469 51008
rect 1795 50968 1804 51008
rect 1844 50968 1996 51008
rect 2036 50968 2045 51008
rect 1420 50672 1460 50968
rect 2140 50756 2180 51640
rect 2572 51176 2612 51640
rect 2851 51556 2860 51596
rect 2900 51556 3031 51596
rect 2572 51136 2900 51176
rect 2563 50968 2572 51008
rect 2612 50968 2764 51008
rect 2804 50968 2813 51008
rect 2860 50840 2900 51136
rect 3436 50924 3476 51640
rect 3532 51596 3572 51724
rect 4483 51640 4492 51680
rect 4532 51640 4828 51680
rect 4868 51640 4877 51680
rect 3532 51556 5356 51596
rect 5396 51556 5405 51596
rect 4919 51388 4928 51428
rect 4968 51388 5010 51428
rect 5050 51388 5092 51428
rect 5132 51388 5174 51428
rect 5214 51388 5256 51428
rect 5296 51388 5305 51428
rect 5740 51176 5780 51724
rect 5932 51260 5972 51724
rect 6988 51680 7028 51724
rect 6307 51640 6316 51680
rect 6356 51640 6988 51680
rect 7028 51640 7037 51680
rect 7485 51260 7525 51724
rect 8044 51715 8084 51724
rect 9676 51680 9716 51724
rect 10924 51680 10964 51724
rect 11875 51724 11884 51764
rect 11924 51724 12364 51764
rect 12404 51724 12556 51764
rect 12596 51724 12605 51764
rect 12739 51724 12748 51764
rect 12788 51724 13420 51764
rect 14659 51724 14668 51764
rect 14708 51724 14860 51764
rect 14900 51724 14909 51764
rect 14956 51724 16108 51764
rect 16148 51724 16684 51764
rect 17923 51724 17932 51764
rect 17972 51724 17981 51764
rect 18211 51724 18220 51764
rect 18260 51724 18452 51764
rect 18892 51724 19468 51764
rect 8419 51640 8428 51680
rect 8468 51640 9716 51680
rect 10025 51640 10156 51680
rect 10196 51640 10205 51680
rect 10915 51640 10924 51680
rect 10964 51640 10973 51680
rect 11116 51596 11156 51724
rect 13420 51715 13460 51724
rect 12163 51640 12172 51680
rect 12212 51640 12796 51680
rect 12836 51640 12845 51680
rect 13219 51640 13228 51680
rect 13268 51640 13364 51680
rect 13324 51596 13364 51640
rect 14956 51596 14996 51724
rect 16108 51715 16148 51724
rect 16684 51715 16724 51724
rect 16204 51640 16492 51680
rect 16532 51640 16628 51680
rect 16204 51596 16244 51640
rect 16588 51596 16628 51640
rect 17932 51596 17972 51724
rect 7651 51556 7660 51596
rect 7700 51556 7709 51596
rect 11116 51556 12748 51596
rect 12788 51556 12797 51596
rect 13219 51556 13228 51596
rect 13268 51556 13277 51596
rect 13324 51556 14996 51596
rect 15331 51556 15340 51596
rect 15380 51556 16244 51596
rect 16291 51556 16300 51596
rect 16340 51556 16349 51596
rect 16483 51556 16492 51596
rect 16532 51556 16541 51596
rect 16588 51556 17972 51596
rect 7660 51512 7700 51556
rect 7660 51472 13132 51512
rect 13172 51472 13181 51512
rect 13228 51344 13268 51556
rect 8812 51304 13268 51344
rect 5923 51220 5932 51260
rect 5972 51220 5981 51260
rect 7485 51220 7564 51260
rect 7604 51220 7613 51260
rect 8812 51176 8852 51304
rect 12115 51220 12124 51260
rect 12164 51220 12460 51260
rect 12500 51220 12509 51260
rect 14371 51220 14380 51260
rect 14420 51220 16204 51260
rect 16244 51220 16253 51260
rect 16300 51176 16340 51556
rect 5740 51136 8852 51176
rect 9004 51136 13324 51176
rect 13364 51136 13373 51176
rect 15724 51136 16340 51176
rect 16492 51176 16532 51556
rect 17321 51220 17452 51260
rect 17492 51220 17501 51260
rect 16492 51136 17300 51176
rect 4099 51052 4108 51092
rect 4148 51052 4492 51092
rect 4532 51052 4541 51092
rect 5740 51083 5780 51092
rect 5827 51052 5836 51092
rect 5876 51052 6124 51092
rect 6164 51052 6508 51092
rect 6548 51052 6557 51092
rect 7372 51083 7948 51092
rect 5740 51008 5780 51043
rect 7412 51052 7948 51083
rect 7988 51052 7997 51092
rect 8899 51052 8908 51092
rect 8948 51052 8957 51092
rect 7372 51008 7412 51043
rect 8908 51008 8948 51052
rect 5740 50968 7180 51008
rect 7220 50968 7412 51008
rect 7747 50968 7756 51008
rect 7796 50968 8948 51008
rect 9004 50924 9044 51136
rect 15724 51092 15764 51136
rect 10156 51083 10196 51092
rect 10531 51052 10540 51092
rect 10580 51052 10828 51092
rect 10868 51052 10877 51092
rect 11683 51052 11692 51092
rect 11732 51083 12500 51092
rect 11732 51052 11788 51083
rect 10156 51008 10196 51043
rect 11828 51052 12500 51083
rect 12739 51052 12748 51092
rect 12788 51083 13556 51092
rect 12788 51052 13516 51083
rect 11788 51034 11828 51043
rect 12460 51008 12500 51052
rect 14755 51052 14764 51092
rect 14804 51052 15340 51092
rect 15380 51052 15389 51092
rect 15706 51052 15715 51092
rect 15755 51052 15764 51092
rect 15811 51052 15820 51092
rect 15860 51052 15869 51092
rect 16073 51052 16204 51092
rect 16244 51052 16253 51092
rect 16649 51052 16780 51092
rect 16820 51052 16829 51092
rect 17260 51083 17300 51136
rect 18892 51092 18932 51724
rect 19468 51715 19508 51724
rect 19529 51556 19660 51596
rect 19700 51556 19709 51596
rect 20371 51556 20380 51596
rect 20420 51556 20429 51596
rect 20380 51512 20420 51556
rect 20380 51472 21044 51512
rect 20039 51388 20048 51428
rect 20088 51388 20130 51428
rect 20170 51388 20212 51428
rect 20252 51388 20294 51428
rect 20334 51388 20376 51428
rect 20416 51388 20425 51428
rect 21004 51344 21044 51472
rect 21510 51344 21600 51364
rect 21004 51304 21600 51344
rect 21510 51284 21600 51304
rect 19603 51220 19612 51260
rect 19652 51220 19756 51260
rect 19796 51220 19805 51260
rect 13516 51034 13556 51043
rect 15820 51008 15860 51052
rect 16780 51034 16820 51043
rect 17513 51052 17644 51092
rect 17684 51052 17693 51092
rect 17740 51083 18932 51092
rect 17740 51052 18892 51083
rect 17260 51034 17300 51043
rect 10156 50968 10444 51008
rect 10484 50968 11020 51008
rect 11060 50968 11069 51008
rect 11875 50968 11884 51008
rect 11924 50968 12364 51008
rect 12404 50968 12413 51008
rect 12460 50968 13228 51008
rect 13268 50968 13277 51008
rect 15523 50968 15532 51008
rect 15572 50968 15860 51008
rect 16169 50968 16300 51008
rect 16340 50968 16349 51008
rect 3436 50884 9044 50924
rect 11020 50924 11060 50968
rect 17740 50924 17780 51052
rect 18892 51034 18932 51043
rect 19756 51052 21196 51092
rect 21236 51052 21245 51092
rect 19756 51008 19796 51052
rect 19241 50968 19372 51008
rect 19412 50968 19421 51008
rect 19747 50968 19756 51008
rect 19796 50968 19805 51008
rect 20131 50968 20140 51008
rect 20180 50968 21100 51008
rect 21140 50968 21149 51008
rect 11020 50884 17780 50924
rect 19987 50884 19996 50924
rect 20036 50884 20852 50924
rect 20812 50840 20852 50884
rect 21510 50840 21600 50860
rect 2371 50800 2380 50840
rect 2420 50800 2524 50840
rect 2564 50800 2573 50840
rect 2860 50800 8716 50840
rect 8756 50800 8765 50840
rect 10217 50800 10348 50840
rect 10388 50800 10397 50840
rect 11849 50800 11980 50840
rect 12020 50800 12029 50840
rect 19075 50800 19084 50840
rect 19124 50800 19133 50840
rect 20371 50800 20380 50840
rect 20420 50800 20716 50840
rect 20756 50800 20765 50840
rect 20812 50800 21600 50840
rect 19084 50756 19124 50800
rect 21510 50780 21600 50800
rect 2140 50716 7564 50756
rect 7604 50716 7613 50756
rect 19084 50716 20236 50756
rect 20276 50716 20285 50756
rect 1420 50632 2956 50672
rect 2996 50632 3005 50672
rect 3679 50632 3688 50672
rect 3728 50632 3770 50672
rect 3810 50632 3852 50672
rect 3892 50632 3934 50672
rect 3974 50632 4016 50672
rect 4056 50632 4065 50672
rect 4483 50632 4492 50672
rect 4532 50632 7756 50672
rect 7796 50632 7805 50672
rect 18799 50632 18808 50672
rect 18848 50632 18890 50672
rect 18930 50632 18972 50672
rect 19012 50632 19054 50672
rect 19094 50632 19136 50672
rect 19176 50632 19185 50672
rect 2860 50464 8332 50504
rect 8372 50464 8381 50504
rect 8812 50464 9332 50504
rect 11011 50464 11020 50504
rect 11060 50464 11828 50504
rect 2860 50252 2900 50464
rect 8812 50420 8852 50464
rect 9292 50420 9332 50464
rect 11788 50420 11828 50464
rect 5260 50380 8852 50420
rect 8899 50380 8908 50420
rect 8948 50380 9196 50420
rect 9236 50380 9245 50420
rect 9292 50380 10964 50420
rect 11616 50380 11692 50420
rect 11732 50380 11741 50420
rect 11788 50380 11932 50420
rect 11972 50380 11981 50420
rect 15619 50380 15628 50420
rect 15668 50380 18460 50420
rect 18500 50380 18509 50420
rect 19084 50380 19660 50420
rect 19700 50380 19709 50420
rect 2083 50212 2092 50252
rect 2132 50212 2900 50252
rect 3340 50252 3380 50261
rect 5260 50252 5300 50380
rect 8995 50296 9004 50336
rect 9044 50296 9332 50336
rect 9667 50296 9676 50336
rect 9716 50296 10060 50336
rect 10100 50296 10109 50336
rect 8716 50252 8756 50261
rect 9292 50252 9332 50296
rect 10252 50252 10292 50261
rect 10924 50252 10964 50380
rect 11692 50336 11732 50380
rect 11273 50296 11404 50336
rect 11444 50296 11453 50336
rect 11683 50296 11692 50336
rect 11732 50296 11741 50336
rect 12137 50296 12268 50336
rect 12308 50296 12317 50336
rect 13804 50296 15916 50336
rect 15956 50296 15965 50336
rect 16265 50296 16396 50336
rect 16436 50296 16445 50336
rect 13804 50252 13844 50296
rect 15436 50252 15476 50296
rect 16972 50252 17012 50261
rect 19084 50252 19124 50380
rect 21510 50336 21600 50356
rect 19459 50296 19468 50336
rect 19508 50296 19660 50336
rect 19700 50296 19709 50336
rect 20227 50296 20236 50336
rect 20276 50296 20285 50336
rect 20707 50296 20716 50336
rect 20756 50296 21600 50336
rect 19180 50252 19220 50261
rect 20236 50252 20276 50296
rect 21510 50276 21600 50296
rect 4003 50212 4012 50252
rect 4052 50212 4300 50252
rect 4340 50212 4349 50252
rect 7459 50212 7468 50252
rect 7508 50212 7604 50252
rect 8131 50212 8140 50252
rect 8180 50212 8524 50252
rect 8564 50212 8716 50252
rect 9178 50212 9187 50252
rect 9227 50212 9236 50252
rect 9283 50212 9292 50252
rect 9332 50212 9341 50252
rect 9641 50212 9772 50252
rect 9812 50212 9821 50252
rect 10121 50212 10156 50252
rect 10196 50212 10252 50252
rect 10339 50212 10348 50252
rect 10388 50212 10740 50252
rect 10780 50212 10789 50252
rect 10924 50212 12116 50252
rect 12425 50212 12556 50252
rect 12596 50212 12605 50252
rect 12940 50212 13804 50252
rect 13987 50212 13996 50252
rect 14036 50212 14188 50252
rect 14228 50212 14237 50252
rect 15898 50212 15907 50252
rect 15947 50212 15956 50252
rect 16003 50212 16012 50252
rect 16052 50212 16061 50252
rect 16483 50212 16492 50252
rect 16532 50212 16876 50252
rect 16916 50212 16925 50252
rect 17451 50212 17460 50252
rect 17500 50212 17509 50252
rect 18682 50212 18691 50252
rect 18731 50212 19124 50252
rect 19171 50212 19180 50252
rect 19220 50212 19351 50252
rect 19625 50212 19756 50252
rect 19796 50212 19805 50252
rect 20131 50212 20140 50252
rect 20180 50212 20189 50252
rect 20232 50212 20241 50252
rect 20281 50212 20323 50252
rect 3340 50168 3380 50212
rect 5260 50168 5300 50212
rect 3340 50128 5300 50168
rect 3401 50044 3532 50084
rect 3572 50044 3581 50084
rect 5260 50000 5300 50128
rect 5443 50044 5452 50084
rect 5492 50044 5740 50084
rect 5780 50044 5789 50084
rect 4780 49960 5300 50000
rect 2860 49624 3340 49664
rect 3380 49624 3389 49664
rect 2860 49580 2900 49624
rect 4780 49580 4820 49960
rect 4919 49876 4928 49916
rect 4968 49876 5010 49916
rect 5050 49876 5092 49916
rect 5132 49876 5174 49916
rect 5214 49876 5256 49916
rect 5296 49876 5305 49916
rect 7564 49664 7604 50212
rect 8716 50203 8756 50212
rect 9196 49748 9236 50212
rect 10252 50203 10292 50212
rect 12076 50168 12116 50212
rect 12940 50168 12980 50212
rect 13804 50203 13844 50212
rect 15436 50203 15476 50212
rect 12076 50128 12980 50168
rect 9283 50044 9292 50084
rect 9332 50044 10924 50084
rect 10964 50044 10973 50084
rect 11155 50044 11164 50084
rect 11204 50044 11308 50084
rect 11348 50044 11357 50084
rect 11875 50044 11884 50084
rect 11924 50044 12028 50084
rect 12068 50044 12077 50084
rect 13987 50044 13996 50084
rect 14036 50044 15340 50084
rect 15380 50044 15389 50084
rect 15619 50044 15628 50084
rect 15668 50044 15820 50084
rect 15860 50044 15869 50084
rect 9292 49792 14188 49832
rect 14228 49792 14237 49832
rect 9187 49708 9196 49748
rect 9236 49708 9245 49748
rect 9292 49664 9332 49792
rect 15916 49748 15956 50212
rect 16012 50084 16052 50212
rect 16972 50168 17012 50212
rect 16195 50128 16204 50168
rect 16244 50128 17012 50168
rect 16012 50044 16300 50084
rect 16340 50044 17068 50084
rect 17108 50044 17117 50084
rect 17452 49748 17492 50212
rect 19180 50203 19220 50212
rect 20140 50168 20180 50212
rect 20140 50128 20524 50168
rect 20564 50128 20573 50168
rect 17635 50044 17644 50084
rect 17684 50044 17693 50084
rect 10915 49708 10924 49748
rect 10964 49708 11404 49748
rect 11444 49708 11453 49748
rect 15811 49708 15820 49748
rect 15860 49708 15956 49748
rect 17443 49708 17452 49748
rect 17492 49708 17501 49748
rect 17644 49664 17684 50044
rect 20039 49876 20048 49916
rect 20088 49876 20130 49916
rect 20170 49876 20212 49916
rect 20252 49876 20294 49916
rect 20334 49876 20376 49916
rect 20416 49876 20425 49916
rect 21510 49832 21600 49852
rect 20380 49792 21600 49832
rect 20380 49748 20420 49792
rect 21510 49772 21600 49792
rect 20371 49708 20380 49748
rect 20420 49708 20429 49748
rect 7564 49624 9332 49664
rect 9388 49624 10444 49664
rect 10484 49624 10493 49664
rect 11107 49624 11116 49664
rect 11156 49624 11836 49664
rect 11876 49624 11885 49664
rect 16195 49624 16204 49664
rect 16244 49624 17684 49664
rect 7564 49580 7604 49624
rect 9388 49580 9428 49624
rect 1987 49540 1996 49580
rect 2036 49540 2900 49580
rect 3244 49571 4820 49580
rect 3284 49540 4204 49571
rect 3244 49522 3284 49531
rect 4244 49540 4820 49571
rect 5443 49540 5452 49580
rect 5492 49540 6124 49580
rect 6164 49540 6173 49580
rect 6316 49571 7180 49580
rect 4204 49522 4244 49531
rect 6356 49540 7180 49571
rect 7220 49540 7229 49580
rect 7555 49540 7564 49580
rect 7604 49540 7613 49580
rect 7747 49540 7756 49580
rect 7796 49540 7805 49580
rect 7939 49540 7948 49580
rect 7988 49571 9428 49580
rect 7988 49540 9004 49571
rect 6316 49522 6356 49531
rect 7756 49496 7796 49540
rect 9044 49540 9428 49571
rect 9475 49540 9484 49580
rect 9524 49540 9667 49580
rect 9707 49540 9716 49580
rect 9763 49540 9772 49580
rect 9812 49540 9943 49580
rect 10025 49540 10156 49580
rect 10196 49540 10205 49580
rect 10601 49540 10732 49580
rect 10772 49540 10781 49580
rect 11081 49540 11212 49580
rect 11252 49540 11261 49580
rect 11971 49540 11980 49580
rect 12020 49540 12029 49580
rect 13097 49540 13228 49580
rect 13268 49540 13277 49580
rect 14371 49540 14380 49580
rect 14420 49540 14429 49580
rect 15497 49540 15628 49580
rect 15668 49540 15677 49580
rect 16003 49540 16012 49580
rect 16052 49540 16876 49580
rect 16916 49540 16925 49580
rect 17260 49571 17300 49580
rect 9004 49522 9044 49531
rect 10732 49522 10772 49531
rect 11212 49522 11252 49531
rect 6499 49456 6508 49496
rect 6548 49456 7796 49496
rect 10121 49456 10252 49496
rect 10292 49456 10301 49496
rect 11299 49456 11308 49496
rect 11348 49456 11596 49496
rect 11636 49456 11645 49496
rect 11980 49412 12020 49540
rect 13228 49522 13268 49531
rect 14380 49412 14420 49540
rect 15628 49496 15668 49531
rect 17260 49496 17300 49531
rect 15628 49456 17300 49496
rect 17827 49456 17836 49496
rect 17876 49456 17885 49496
rect 19241 49456 19372 49496
rect 19412 49456 19421 49496
rect 19747 49456 19756 49496
rect 19796 49456 19805 49496
rect 19939 49456 19948 49496
rect 19988 49456 20140 49496
rect 20180 49456 20189 49496
rect 17836 49412 17876 49456
rect 19756 49412 19796 49456
rect 3427 49372 3436 49412
rect 3476 49372 4108 49412
rect 4148 49372 4157 49412
rect 6211 49372 6220 49412
rect 6260 49372 12020 49412
rect 12835 49372 12844 49412
rect 12884 49372 14420 49412
rect 16291 49372 16300 49412
rect 16340 49372 17876 49412
rect 17932 49372 19796 49412
rect 19987 49372 19996 49412
rect 20036 49372 20852 49412
rect 4003 49288 4012 49328
rect 4052 49288 4684 49328
rect 4724 49288 4733 49328
rect 6115 49288 6124 49328
rect 6164 49288 6604 49328
rect 6644 49288 6653 49328
rect 13289 49288 13420 49328
rect 13460 49288 13469 49328
rect 17587 49288 17596 49328
rect 17636 49288 17644 49328
rect 17684 49288 17767 49328
rect 17932 49244 17972 49372
rect 20812 49328 20852 49372
rect 21510 49328 21600 49348
rect 19603 49288 19612 49328
rect 19652 49288 20428 49328
rect 20468 49288 20477 49328
rect 20812 49288 21600 49328
rect 21510 49268 21600 49288
rect 15715 49204 15724 49244
rect 15764 49204 17972 49244
rect 3679 49120 3688 49160
rect 3728 49120 3770 49160
rect 3810 49120 3852 49160
rect 3892 49120 3934 49160
rect 3974 49120 4016 49160
rect 4056 49120 4065 49160
rect 18799 49120 18808 49160
rect 18848 49120 18890 49160
rect 18930 49120 18972 49160
rect 19012 49120 19054 49160
rect 19094 49120 19136 49160
rect 19176 49120 19185 49160
rect 11203 48952 11212 48992
rect 11252 48952 11404 48992
rect 11444 48952 11453 48992
rect 15811 48952 15820 48992
rect 15860 48952 15869 48992
rect 19084 48952 19468 48992
rect 19508 48952 19517 48992
rect 15820 48908 15860 48952
rect 19084 48908 19124 48952
rect 4195 48868 4204 48908
rect 4244 48868 4540 48908
rect 4580 48868 4589 48908
rect 5164 48868 6988 48908
rect 7028 48868 7037 48908
rect 8489 48868 8572 48908
rect 8612 48868 8620 48908
rect 8660 48868 8669 48908
rect 14467 48868 14476 48908
rect 14516 48868 14716 48908
rect 14756 48868 14765 48908
rect 15820 48868 16916 48908
rect 18211 48868 18220 48908
rect 18260 48868 19124 48908
rect 19180 48868 19756 48908
rect 19796 48868 19805 48908
rect 20419 48868 20428 48908
rect 20468 48868 21236 48908
rect 5164 48824 5204 48868
rect 2755 48784 2764 48824
rect 2804 48784 3820 48824
rect 3860 48784 3869 48824
rect 4649 48784 4780 48824
rect 4820 48784 4829 48824
rect 5068 48784 5204 48824
rect 5539 48784 5548 48824
rect 5588 48784 5876 48824
rect 8777 48784 8812 48824
rect 8852 48784 8908 48824
rect 8948 48784 8956 48824
rect 8996 48784 9005 48824
rect 9065 48784 9196 48824
rect 9236 48784 9245 48824
rect 9545 48784 9676 48824
rect 9716 48784 9725 48824
rect 11692 48784 11980 48824
rect 12020 48784 12029 48824
rect 12163 48784 12172 48824
rect 12212 48784 12343 48824
rect 14947 48784 14956 48824
rect 14996 48784 15532 48824
rect 15572 48784 15581 48824
rect 15916 48784 16300 48824
rect 16340 48784 16349 48824
rect 5068 48740 5108 48784
rect 5050 48700 5059 48740
rect 5099 48700 5108 48740
rect 5155 48700 5164 48740
rect 5204 48700 5213 48740
rect 5513 48700 5644 48740
rect 5684 48700 5693 48740
rect 5164 48656 5204 48700
rect 4387 48616 4396 48656
rect 4436 48616 5204 48656
rect 4051 48532 4060 48572
rect 4100 48532 4204 48572
rect 4244 48532 4253 48572
rect 5836 48488 5876 48784
rect 6124 48740 6164 48749
rect 7180 48740 7220 48749
rect 11212 48740 11252 48749
rect 11692 48740 11732 48784
rect 12748 48740 12788 48749
rect 15820 48740 15860 48749
rect 5993 48700 6124 48740
rect 6164 48700 6173 48740
rect 6595 48700 6604 48740
rect 6652 48700 6775 48740
rect 7049 48700 7180 48740
rect 7220 48700 7948 48740
rect 7988 48700 7997 48740
rect 8419 48700 8428 48740
rect 8468 48700 8812 48740
rect 8852 48700 8861 48740
rect 9833 48700 9964 48740
rect 10004 48700 10013 48740
rect 10627 48700 10636 48740
rect 10676 48700 11212 48740
rect 11674 48700 11683 48740
rect 11723 48700 11732 48740
rect 11779 48700 11788 48740
rect 11828 48700 11837 48740
rect 12137 48700 12268 48740
rect 12308 48700 12317 48740
rect 12617 48700 12748 48740
rect 12788 48700 12797 48740
rect 13258 48700 13267 48740
rect 13307 48700 13420 48740
rect 13460 48700 13469 48740
rect 15209 48700 15331 48740
rect 15380 48700 15389 48740
rect 15689 48700 15820 48740
rect 15860 48700 15869 48740
rect 6124 48691 6164 48700
rect 7180 48691 7220 48700
rect 11212 48691 11252 48700
rect 11788 48656 11828 48700
rect 12748 48691 12788 48700
rect 15820 48691 15860 48700
rect 11788 48616 12652 48656
rect 12692 48616 12701 48656
rect 6665 48532 6796 48572
rect 6836 48532 6845 48572
rect 9388 48532 9436 48572
rect 9476 48532 9485 48572
rect 13385 48532 13420 48572
rect 13460 48532 13516 48572
rect 13556 48532 13565 48572
rect 15139 48532 15148 48572
rect 15188 48532 15820 48572
rect 15860 48532 15869 48572
rect 5705 48448 5836 48488
rect 5876 48448 8236 48488
rect 8276 48448 8285 48488
rect 4919 48364 4928 48404
rect 4968 48364 5010 48404
rect 5050 48364 5092 48404
rect 5132 48364 5174 48404
rect 5214 48364 5256 48404
rect 5296 48364 5305 48404
rect 3907 48196 3916 48236
rect 3956 48196 4492 48236
rect 4532 48196 4541 48236
rect 5923 48196 5932 48236
rect 5972 48196 6412 48236
rect 6452 48196 6461 48236
rect 1987 48112 1996 48152
rect 2036 48112 2324 48152
rect 3197 48112 3244 48152
rect 3284 48112 3293 48152
rect 5260 48112 7468 48152
rect 7508 48112 7517 48152
rect 2284 48068 2324 48112
rect 2170 48028 2179 48068
rect 2219 48028 2228 48068
rect 2275 48028 2284 48068
rect 2324 48028 2333 48068
rect 2537 48028 2668 48068
rect 2708 48028 2717 48068
rect 3244 48059 3284 48112
rect 2188 47984 2228 48028
rect 3331 48028 3340 48068
rect 3380 48059 3764 48068
rect 3380 48028 3724 48059
rect 3244 48010 3284 48019
rect 4043 48028 4108 48068
rect 4148 48028 4174 48068
rect 4214 48028 4223 48068
rect 4289 48028 4298 48068
rect 4338 48028 4347 48068
rect 4553 48028 4588 48068
rect 4628 48028 4684 48068
rect 4724 48028 4733 48068
rect 5260 48059 5300 48112
rect 9388 48068 9428 48532
rect 15916 48068 15956 48784
rect 16876 48759 16916 48868
rect 17539 48784 17548 48824
rect 17588 48784 18316 48824
rect 18356 48784 18365 48824
rect 18473 48784 18604 48824
rect 18644 48784 18653 48824
rect 16265 48700 16396 48740
rect 16436 48700 16445 48740
rect 16771 48700 16780 48740
rect 16820 48700 16829 48740
rect 16876 48719 16893 48759
rect 16933 48719 16942 48759
rect 19180 48740 19220 48868
rect 21196 48824 21236 48868
rect 21510 48824 21600 48844
rect 19363 48784 19372 48824
rect 19412 48784 19996 48824
rect 20036 48784 20045 48824
rect 20227 48784 20236 48824
rect 20276 48784 20524 48824
rect 20564 48784 21100 48824
rect 21140 48784 21149 48824
rect 21196 48784 21600 48824
rect 21510 48764 21600 48784
rect 18106 48700 18115 48740
rect 18155 48700 18164 48740
rect 18211 48700 18220 48740
rect 18260 48700 18391 48740
rect 18691 48700 18700 48740
rect 18740 48700 18749 48740
rect 19459 48700 19468 48740
rect 19508 48700 19668 48740
rect 19708 48700 19717 48740
rect 16780 48656 16820 48700
rect 16780 48616 16972 48656
rect 17012 48616 17021 48656
rect 18124 48236 18164 48700
rect 18700 48656 18740 48700
rect 19180 48691 19220 48700
rect 18307 48616 18316 48656
rect 18356 48616 18740 48656
rect 19843 48532 19852 48572
rect 19892 48532 20812 48572
rect 20852 48532 20861 48572
rect 20039 48364 20048 48404
rect 20088 48364 20130 48404
rect 20170 48364 20212 48404
rect 20252 48364 20294 48404
rect 20334 48364 20376 48404
rect 20416 48364 20425 48404
rect 21510 48320 21600 48340
rect 20380 48280 21600 48320
rect 20380 48236 20420 48280
rect 21510 48260 21600 48280
rect 17321 48196 17452 48236
rect 17492 48196 17501 48236
rect 18124 48196 19084 48236
rect 19124 48196 19133 48236
rect 20371 48196 20380 48236
rect 20420 48196 20429 48236
rect 3724 48010 3764 48019
rect 4300 47984 4340 48028
rect 5609 48028 5740 48068
rect 5780 48028 5789 48068
rect 9292 48028 10388 48068
rect 12809 48028 12940 48068
rect 12980 48028 12989 48068
rect 13219 48028 13228 48068
rect 13268 48059 14284 48068
rect 13268 48028 14188 48059
rect 5260 48010 5300 48019
rect 5740 48010 5780 48019
rect 9292 47984 9332 48028
rect 10348 47984 10388 48028
rect 14228 48028 14284 48059
rect 14324 48028 14333 48068
rect 15706 48028 15715 48068
rect 15755 48028 15764 48068
rect 15811 48028 15820 48068
rect 15860 48028 15956 48068
rect 16073 48028 16204 48068
rect 16244 48028 16253 48068
rect 16387 48028 16396 48068
rect 16436 48059 16820 48068
rect 16436 48028 16780 48059
rect 14188 48010 14228 48019
rect 15724 47984 15764 48028
rect 2179 47944 2188 47984
rect 2228 47944 2275 47984
rect 2633 47944 2764 47984
rect 2804 47944 2813 47984
rect 4195 47944 4204 47984
rect 4244 47944 4340 47984
rect 4745 47944 4780 47984
rect 4820 47944 4876 47984
rect 4916 47944 4925 47984
rect 7913 47944 7948 47984
rect 7988 47944 8044 47984
rect 8084 47944 8093 47984
rect 9283 47944 9292 47984
rect 9332 47944 9341 47984
rect 9667 47944 9676 47984
rect 9716 47944 9725 47984
rect 10339 47944 10348 47984
rect 10388 47944 10924 47984
rect 10964 47944 11308 47984
rect 11348 47944 11357 47984
rect 15724 47944 15820 47984
rect 15860 47944 15869 47984
rect 9676 47900 9716 47944
rect 15916 47900 15956 48028
rect 17129 48028 17260 48068
rect 17300 48028 17309 48068
rect 17635 48028 17644 48068
rect 17684 48028 17693 48068
rect 17788 48059 19276 48068
rect 17788 48028 18892 48059
rect 16780 48010 16820 48019
rect 17260 48010 17300 48019
rect 16169 47944 16300 47984
rect 16340 47944 16349 47984
rect 17644 47900 17684 48028
rect 8899 47860 8908 47900
rect 8948 47860 9716 47900
rect 10505 47860 10588 47900
rect 10628 47860 10636 47900
rect 10676 47860 10685 47900
rect 12940 47860 15956 47900
rect 16771 47860 16780 47900
rect 16820 47860 17684 47900
rect 8131 47776 8140 47816
rect 8180 47776 8188 47816
rect 8228 47776 8311 47816
rect 8803 47776 8812 47816
rect 8852 47776 9052 47816
rect 9092 47776 9101 47816
rect 9907 47776 9916 47816
rect 9956 47776 10540 47816
rect 10580 47776 10589 47816
rect 10675 47776 10684 47816
rect 10724 47776 10732 47816
rect 10772 47776 10855 47816
rect 12940 47732 12980 47860
rect 14371 47776 14380 47816
rect 14420 47776 14956 47816
rect 14996 47776 15005 47816
rect 6307 47692 6316 47732
rect 6356 47692 12980 47732
rect 17788 47648 17828 48028
rect 18932 48028 19276 48059
rect 19316 48028 19325 48068
rect 18892 48010 18932 48019
rect 19625 47944 19756 47984
rect 19796 47944 19805 47984
rect 20009 47944 20140 47984
rect 20180 47944 20189 47984
rect 19987 47860 19996 47900
rect 20036 47860 20852 47900
rect 20812 47816 20852 47860
rect 21510 47816 21600 47836
rect 20812 47776 21600 47816
rect 21510 47756 21600 47776
rect 3679 47608 3688 47648
rect 3728 47608 3770 47648
rect 3810 47608 3852 47648
rect 3892 47608 3934 47648
rect 3974 47608 4016 47648
rect 4056 47608 4065 47648
rect 10723 47608 10732 47648
rect 10772 47608 17828 47648
rect 18799 47608 18808 47648
rect 18848 47608 18890 47648
rect 18930 47608 18972 47648
rect 19012 47608 19054 47648
rect 19094 47608 19136 47648
rect 19176 47608 19185 47648
rect 3043 47440 3052 47480
rect 3092 47440 3340 47480
rect 3380 47440 3389 47480
rect 9379 47440 9388 47480
rect 9428 47440 9811 47480
rect 9851 47440 9860 47480
rect 15689 47440 15820 47480
rect 15860 47440 15869 47480
rect 17251 47440 17260 47480
rect 17300 47440 17452 47480
rect 17492 47440 17501 47480
rect 19337 47440 19468 47480
rect 19508 47440 19517 47480
rect 3235 47356 3244 47396
rect 3284 47356 3860 47396
rect 3820 47312 3860 47356
rect 4396 47356 7660 47396
rect 7700 47356 7709 47396
rect 8524 47356 10828 47396
rect 10868 47356 10877 47396
rect 3340 47272 3532 47312
rect 3572 47272 3581 47312
rect 3811 47272 3820 47312
rect 3860 47272 3869 47312
rect 2860 47228 2900 47237
rect 3340 47228 3380 47272
rect 4396 47228 4436 47356
rect 8524 47312 8564 47356
rect 21510 47312 21600 47332
rect 1603 47188 1612 47228
rect 1652 47188 1661 47228
rect 2729 47188 2860 47228
rect 2900 47188 2909 47228
rect 3322 47188 3331 47228
rect 3371 47188 3380 47228
rect 3427 47188 3436 47228
rect 3476 47188 3607 47228
rect 3785 47188 3916 47228
rect 3956 47188 3965 47228
rect 1612 47060 1652 47188
rect 2860 47179 2900 47188
rect 4396 47179 4436 47188
rect 4588 47272 6356 47312
rect 8515 47272 8524 47312
rect 8564 47272 8573 47312
rect 9100 47272 11500 47312
rect 11540 47272 11549 47312
rect 15628 47272 17300 47312
rect 19625 47272 19660 47312
rect 19700 47272 19756 47312
rect 19796 47272 19805 47312
rect 20131 47272 20140 47312
rect 20180 47272 20189 47312
rect 20371 47272 20380 47312
rect 20420 47272 21600 47312
rect 4588 47060 4628 47272
rect 6316 47228 6356 47272
rect 7564 47228 7604 47237
rect 9100 47228 9140 47272
rect 12076 47228 12116 47237
rect 13996 47228 14036 47237
rect 15628 47228 15668 47272
rect 17260 47228 17300 47272
rect 19276 47228 19316 47237
rect 20140 47228 20180 47272
rect 21510 47252 21600 47272
rect 4675 47188 4684 47228
rect 4724 47188 4884 47228
rect 4924 47188 4933 47228
rect 6115 47188 6124 47228
rect 6164 47188 6173 47228
rect 6307 47188 6316 47228
rect 6356 47188 6365 47228
rect 1612 47020 4628 47060
rect 4771 47020 4780 47060
rect 4820 47020 5068 47060
rect 5108 47020 5117 47060
rect 5635 47020 5644 47060
rect 5684 47020 5980 47060
rect 6020 47020 6029 47060
rect 4919 46852 4928 46892
rect 4968 46852 5010 46892
rect 5050 46852 5092 46892
rect 5132 46852 5174 46892
rect 5214 46852 5256 46892
rect 5296 46852 5305 46892
rect 6124 46724 6164 47188
rect 6316 46976 6356 47188
rect 7564 47060 7604 47188
rect 7756 47188 8035 47228
rect 8075 47188 8084 47228
rect 8131 47188 8140 47228
rect 8180 47188 8189 47228
rect 8611 47188 8620 47228
rect 8660 47188 8791 47228
rect 9379 47188 9388 47228
rect 9428 47188 9588 47228
rect 9628 47188 9637 47228
rect 10435 47188 10444 47228
rect 10484 47188 10615 47228
rect 10819 47188 10828 47228
rect 10868 47188 10877 47228
rect 11587 47188 11596 47228
rect 11636 47188 12076 47228
rect 12259 47188 12268 47228
rect 12308 47188 12748 47228
rect 12788 47188 12844 47228
rect 12884 47188 12948 47228
rect 13865 47188 13996 47228
rect 14036 47188 14045 47228
rect 14371 47188 14380 47228
rect 14420 47188 14572 47228
rect 14612 47188 14621 47228
rect 15497 47188 15628 47228
rect 15668 47188 15677 47228
rect 15811 47188 15820 47228
rect 15860 47188 16012 47228
rect 16052 47188 16061 47228
rect 17897 47188 18028 47228
rect 18068 47188 18077 47228
rect 19145 47188 19276 47228
rect 19316 47188 19325 47228
rect 20140 47188 20524 47228
rect 20564 47188 20573 47228
rect 7756 47144 7796 47188
rect 8140 47144 8180 47188
rect 9100 47179 9140 47188
rect 7747 47104 7756 47144
rect 7796 47104 7805 47144
rect 8140 47104 9044 47144
rect 7564 47020 8908 47060
rect 8948 47020 8957 47060
rect 6316 46936 8524 46976
rect 8564 46936 8573 46976
rect 9004 46892 9044 47104
rect 10828 47060 10868 47188
rect 12076 47179 12116 47188
rect 13996 47179 14036 47188
rect 15628 47179 15668 47188
rect 17260 47179 17300 47188
rect 19276 47179 19316 47188
rect 12172 47104 12980 47144
rect 12172 47060 12212 47104
rect 10579 47020 10588 47060
rect 10628 47020 10637 47060
rect 10828 47020 12212 47060
rect 12259 47020 12268 47060
rect 12308 47020 12556 47060
rect 12596 47020 12605 47060
rect 10588 46976 10628 47020
rect 10588 46936 11212 46976
rect 11252 46936 11261 46976
rect 12940 46892 12980 47104
rect 14057 47020 14188 47060
rect 14228 47020 14237 47060
rect 19987 47020 19996 47060
rect 20036 47020 20756 47060
rect 9004 46852 10772 46892
rect 12940 46852 15820 46892
rect 15860 46852 15869 46892
rect 20039 46852 20048 46892
rect 20088 46852 20130 46892
rect 20170 46852 20212 46892
rect 20252 46852 20294 46892
rect 20334 46852 20376 46892
rect 20416 46852 20425 46892
rect 2179 46684 2188 46724
rect 2228 46684 2764 46724
rect 2804 46684 2813 46724
rect 3331 46684 3340 46724
rect 3380 46684 3868 46724
rect 3908 46684 3917 46724
rect 4339 46684 4348 46724
rect 4388 46684 4684 46724
rect 4724 46684 4733 46724
rect 5347 46684 5356 46724
rect 5396 46684 6164 46724
rect 9257 46684 9388 46724
rect 9428 46684 9437 46724
rect 10217 46684 10348 46724
rect 10388 46684 10397 46724
rect 10732 46640 10772 46852
rect 20716 46808 20756 47020
rect 21510 46808 21600 46828
rect 11683 46768 11692 46808
rect 11732 46768 12076 46808
rect 12116 46768 12125 46808
rect 20716 46768 21600 46808
rect 21510 46748 21600 46768
rect 14755 46684 14764 46724
rect 14804 46684 15148 46724
rect 15188 46684 15197 46724
rect 1324 46600 5492 46640
rect 1324 46556 1364 46600
rect 1315 46516 1324 46556
rect 1364 46516 1373 46556
rect 2572 46547 2860 46556
rect 2612 46516 2860 46547
rect 2900 46516 2909 46556
rect 4954 46516 4963 46556
rect 5003 46516 5356 46556
rect 5396 46516 5405 46556
rect 2572 46498 2612 46507
rect 3427 46432 3436 46472
rect 3476 46432 3628 46472
rect 3668 46432 3677 46472
rect 4099 46432 4108 46472
rect 4148 46432 4157 46472
rect 4361 46432 4492 46472
rect 4532 46432 4541 46472
rect 4108 46388 4148 46432
rect 5452 46388 5492 46600
rect 5548 46600 8140 46640
rect 8180 46600 8189 46640
rect 9772 46600 10100 46640
rect 5548 46547 5588 46600
rect 9772 46556 9812 46600
rect 10060 46556 10100 46600
rect 10732 46600 13556 46640
rect 13987 46600 13996 46640
rect 14036 46600 15572 46640
rect 10732 46556 10772 46600
rect 13516 46556 13556 46600
rect 6625 46516 6700 46556
rect 6740 46516 6756 46556
rect 6796 46516 6805 46556
rect 6857 46516 6988 46556
rect 7028 46516 7037 46556
rect 7171 46516 7180 46556
rect 7220 46516 7324 46556
rect 7364 46516 7380 46556
rect 7459 46516 7468 46556
rect 7508 46516 7639 46556
rect 7939 46516 7948 46556
rect 7988 46516 8852 46556
rect 8899 46516 8908 46556
rect 8948 46547 9236 46556
rect 8948 46516 9196 46547
rect 5548 46498 5588 46507
rect 8812 46388 8852 46516
rect 9449 46516 9580 46556
rect 9620 46516 9629 46556
rect 9754 46516 9763 46556
rect 9803 46516 9812 46556
rect 9859 46516 9868 46556
rect 9908 46516 9917 46556
rect 10051 46516 10060 46556
rect 10100 46516 10109 46556
rect 10193 46516 10202 46556
rect 10242 46516 10252 46556
rect 10292 46516 10382 46556
rect 10618 46516 10627 46556
rect 10667 46516 10676 46556
rect 10723 46516 10732 46556
rect 10772 46516 10781 46556
rect 10985 46516 11116 46556
rect 11156 46516 11165 46556
rect 11299 46516 11308 46556
rect 11348 46516 11500 46556
rect 11540 46547 11732 46556
rect 11540 46516 11692 46547
rect 9196 46498 9236 46507
rect 9772 46472 9812 46516
rect 9868 46472 9908 46516
rect 10636 46472 10676 46516
rect 11692 46498 11732 46507
rect 12172 46547 12556 46556
rect 12212 46516 12556 46547
rect 12596 46516 12605 46556
rect 13402 46516 13411 46556
rect 13451 46516 13460 46556
rect 13507 46516 13516 46556
rect 13556 46516 13612 46556
rect 13652 46516 13687 46556
rect 13769 46516 13900 46556
rect 13940 46516 13949 46556
rect 14345 46516 14476 46556
rect 14516 46516 14525 46556
rect 14825 46516 14956 46556
rect 14996 46516 15005 46556
rect 15532 46547 15572 46600
rect 12172 46498 12212 46507
rect 13420 46472 13460 46516
rect 14476 46498 14516 46507
rect 14956 46498 14996 46507
rect 16745 46516 16780 46556
rect 16820 46516 16876 46556
rect 16916 46516 16925 46556
rect 17539 46516 17548 46556
rect 17588 46516 17836 46556
rect 17876 46516 17885 46556
rect 19084 46547 19124 46556
rect 15532 46472 15572 46507
rect 19084 46472 19124 46507
rect 9725 46432 9772 46472
rect 9812 46432 9821 46472
rect 9868 46432 10444 46472
rect 10484 46432 10493 46472
rect 10627 46432 10636 46472
rect 10676 46432 10723 46472
rect 10819 46432 10828 46472
rect 10868 46432 11212 46472
rect 11252 46432 11636 46472
rect 12394 46432 12403 46472
rect 12443 46432 12748 46472
rect 12788 46432 12797 46472
rect 13411 46432 13420 46472
rect 13460 46432 13507 46472
rect 13987 46432 13996 46472
rect 14036 46432 14380 46472
rect 14420 46432 14429 46472
rect 15532 46432 17356 46472
rect 17396 46432 19124 46472
rect 19747 46432 19756 46472
rect 19796 46432 19805 46472
rect 20009 46432 20140 46472
rect 20180 46432 20189 46472
rect 11596 46388 11636 46432
rect 19756 46388 19796 46432
rect 4108 46348 4300 46388
rect 4340 46348 4349 46388
rect 4841 46348 4935 46388
rect 5012 46348 5021 46388
rect 5146 46348 5155 46388
rect 5195 46348 5356 46388
rect 5396 46348 5405 46388
rect 5452 46348 11500 46388
rect 11540 46348 11549 46388
rect 11596 46348 14476 46388
rect 14516 46348 14525 46388
rect 17251 46348 17260 46388
rect 17300 46348 19796 46388
rect 19987 46348 19996 46388
rect 20036 46348 20620 46388
rect 20660 46348 20669 46388
rect 21510 46304 21600 46324
rect 4195 46264 4204 46304
rect 4244 46264 4732 46304
rect 4772 46264 4781 46304
rect 6595 46264 6604 46304
rect 6644 46264 7084 46304
rect 7124 46264 7133 46304
rect 9859 46264 9868 46304
rect 9908 46264 10828 46304
rect 10868 46264 10877 46304
rect 11683 46264 11692 46304
rect 11732 46264 12268 46304
rect 12308 46264 12317 46304
rect 12499 46264 12508 46304
rect 12548 46264 12556 46304
rect 12596 46264 12679 46304
rect 15209 46264 15340 46304
rect 15380 46264 15389 46304
rect 19145 46264 19276 46304
rect 19316 46264 19325 46304
rect 20371 46264 20380 46304
rect 20420 46264 21600 46304
rect 21510 46244 21600 46264
rect 2860 46180 6740 46220
rect 2860 46136 2900 46180
rect 6700 46136 6740 46180
rect 12940 46180 17548 46220
rect 17588 46180 17597 46220
rect 12940 46136 12980 46180
rect 2275 46096 2284 46136
rect 2324 46096 2900 46136
rect 3679 46096 3688 46136
rect 3728 46096 3770 46136
rect 3810 46096 3852 46136
rect 3892 46096 3934 46136
rect 3974 46096 4016 46136
rect 4056 46096 4065 46136
rect 5443 46096 5452 46136
rect 5492 46096 5876 46136
rect 6691 46096 6700 46136
rect 6740 46096 12980 46136
rect 18799 46096 18808 46136
rect 18848 46096 18890 46136
rect 18930 46096 18972 46136
rect 19012 46096 19054 46136
rect 19094 46096 19136 46136
rect 19176 46096 19185 46136
rect 5836 46052 5876 46096
rect 5251 46012 5260 46052
rect 5300 46012 5740 46052
rect 5780 46012 5789 46052
rect 5836 46012 6220 46052
rect 6260 46012 6269 46052
rect 6316 46012 8236 46052
rect 8276 46012 8285 46052
rect 12940 46012 18412 46052
rect 18452 46012 18461 46052
rect 6316 45968 6356 46012
rect 12940 45968 12980 46012
rect 1843 45928 1852 45968
rect 1892 45928 3916 45968
rect 3956 45928 3965 45968
rect 4675 45928 4684 45968
rect 4724 45928 5401 45968
rect 5443 45928 5452 45968
rect 5492 45928 6356 45968
rect 6403 45928 6412 45968
rect 6452 45928 7852 45968
rect 7892 45928 7901 45968
rect 9641 45928 9772 45968
rect 9812 45928 9821 45968
rect 10147 45928 10156 45968
rect 10196 45928 10205 45968
rect 10627 45928 10636 45968
rect 10676 45928 11404 45968
rect 11444 45928 11453 45968
rect 11692 45928 12980 45968
rect 13289 45928 13420 45968
rect 13460 45928 13469 45968
rect 15043 45928 15052 45968
rect 15092 45928 19564 45968
rect 19604 45928 19613 45968
rect 5361 45884 5401 45928
rect 10156 45884 10196 45928
rect 11692 45884 11732 45928
rect 1459 45844 1468 45884
rect 1508 45844 2900 45884
rect 4771 45844 4780 45884
rect 4820 45844 4868 45884
rect 5059 45844 5068 45884
rect 5108 45844 5164 45884
rect 5204 45844 5239 45884
rect 5361 45844 5492 45884
rect 2860 45800 2900 45844
rect 67 45760 76 45800
rect 116 45760 1228 45800
rect 1268 45760 1277 45800
rect 1603 45760 1612 45800
rect 1652 45760 1661 45800
rect 2860 45760 4012 45800
rect 4052 45760 4061 45800
rect 4396 45760 4492 45800
rect 4532 45760 4541 45800
rect 4674 45760 4684 45800
rect 4724 45760 4761 45800
rect 0 45464 90 45484
rect 0 45424 76 45464
rect 116 45424 125 45464
rect 0 45404 90 45424
rect 0 45128 90 45148
rect 1612 45128 1652 45760
rect 4396 45716 4436 45760
rect 4674 45716 4714 45760
rect 4828 45716 4868 45844
rect 5155 45760 5164 45800
rect 5204 45760 5260 45800
rect 5300 45760 5335 45800
rect 4979 45718 5000 45758
rect 5040 45751 5049 45758
rect 5040 45737 5060 45751
rect 5040 45718 5108 45737
rect 5000 45716 5108 45718
rect 5452 45716 5492 45844
rect 5836 45844 7180 45884
rect 7220 45844 7229 45884
rect 7459 45844 7468 45884
rect 7508 45844 8140 45884
rect 8180 45844 8189 45884
rect 10156 45844 11732 45884
rect 11827 45844 11836 45884
rect 11876 45844 20524 45884
rect 20564 45844 20573 45884
rect 5836 45716 5876 45844
rect 21510 45800 21600 45820
rect 6787 45760 6796 45800
rect 6836 45760 6915 45800
rect 6955 45760 6967 45800
rect 7564 45760 8428 45800
rect 8468 45760 8477 45800
rect 9580 45760 10156 45800
rect 10196 45760 10205 45800
rect 11587 45760 11596 45800
rect 11636 45760 11788 45800
rect 11828 45760 12940 45800
rect 12980 45760 12989 45800
rect 14141 45760 14188 45800
rect 14228 45760 14237 45800
rect 14371 45760 14380 45800
rect 14420 45760 14668 45800
rect 14708 45760 14717 45800
rect 17417 45760 17548 45800
rect 17588 45760 17597 45800
rect 18185 45760 18316 45800
rect 18356 45760 18365 45800
rect 19555 45760 19564 45800
rect 19604 45760 19756 45800
rect 19796 45760 19805 45800
rect 20131 45760 20140 45800
rect 20180 45760 20189 45800
rect 20611 45760 20620 45800
rect 20660 45760 21600 45800
rect 7564 45716 7604 45760
rect 9580 45716 9620 45760
rect 11212 45716 11252 45725
rect 13228 45716 13268 45725
rect 14188 45716 14228 45760
rect 15244 45716 15284 45725
rect 18892 45716 18932 45725
rect 20140 45716 20180 45760
rect 21510 45740 21600 45760
rect 3785 45676 3916 45716
rect 3956 45676 3965 45716
rect 4049 45676 4058 45716
rect 4098 45676 4108 45716
rect 4148 45676 4238 45716
rect 4387 45676 4396 45716
rect 4436 45676 4445 45716
rect 4542 45676 4551 45716
rect 4591 45676 4600 45716
rect 4665 45676 4674 45716
rect 4714 45676 4723 45716
rect 4828 45676 4852 45716
rect 4892 45676 4901 45716
rect 5000 45711 5068 45716
rect 5020 45697 5068 45711
rect 5059 45676 5068 45697
rect 5108 45676 5117 45716
rect 5276 45676 5285 45716
rect 5325 45676 5334 45716
rect 5434 45676 5443 45716
rect 5483 45676 5492 45716
rect 5578 45676 5587 45716
rect 5627 45676 5636 45716
rect 5692 45676 5701 45716
rect 5741 45676 5750 45716
rect 5818 45676 5827 45716
rect 5867 45676 5876 45716
rect 5923 45676 5932 45716
rect 5972 45676 6004 45716
rect 6044 45676 6220 45716
rect 6260 45676 6269 45716
rect 6353 45676 6362 45716
rect 6402 45676 6412 45716
rect 6452 45676 6542 45716
rect 6595 45676 6604 45716
rect 6644 45676 6796 45716
rect 6836 45676 6845 45716
rect 7024 45676 7033 45716
rect 7073 45676 7089 45716
rect 7168 45676 7177 45716
rect 7217 45676 7226 45716
rect 7306 45676 7315 45716
rect 7355 45676 7364 45716
rect 7420 45676 7429 45716
rect 7469 45676 7604 45716
rect 7747 45676 7756 45716
rect 7796 45676 7805 45716
rect 7852 45676 7875 45716
rect 7915 45676 7924 45716
rect 7984 45676 7993 45716
rect 8033 45676 8042 45716
rect 8227 45676 8236 45716
rect 8276 45676 8332 45716
rect 8372 45676 8407 45716
rect 9379 45676 9388 45716
rect 9428 45676 9580 45716
rect 9955 45676 9964 45716
rect 10004 45676 10013 45716
rect 11252 45676 11596 45716
rect 11636 45676 11645 45716
rect 11971 45676 11980 45716
rect 12020 45676 12029 45716
rect 13097 45676 13228 45716
rect 13268 45676 13516 45716
rect 13556 45676 13565 45716
rect 14170 45676 14179 45716
rect 14219 45676 14228 45716
rect 14275 45676 14284 45716
rect 14324 45676 14333 45716
rect 14729 45676 14764 45716
rect 14804 45676 14860 45716
rect 14900 45676 14909 45716
rect 15331 45676 15340 45716
rect 15380 45676 15732 45716
rect 15772 45676 15781 45716
rect 17818 45676 17827 45716
rect 17867 45676 17876 45716
rect 17923 45676 17932 45716
rect 17972 45676 18124 45716
rect 18164 45676 18173 45716
rect 18281 45676 18412 45716
rect 18452 45676 18461 45716
rect 18761 45676 18892 45716
rect 18932 45676 18941 45716
rect 19267 45676 19276 45716
rect 19316 45676 19380 45716
rect 19420 45676 19447 45716
rect 20140 45676 21428 45716
rect 3916 45632 3956 45676
rect 4551 45632 4591 45676
rect 5285 45632 5325 45676
rect 5596 45632 5636 45676
rect 3916 45592 4591 45632
rect 5260 45592 5325 45632
rect 5500 45592 5636 45632
rect 5698 45632 5738 45676
rect 7049 45632 7089 45676
rect 7180 45632 7220 45676
rect 7324 45632 7364 45676
rect 5698 45592 6068 45632
rect 6569 45592 6700 45632
rect 6740 45592 6749 45632
rect 6979 45592 6988 45632
rect 7028 45592 7089 45632
rect 7171 45592 7180 45632
rect 7220 45592 7264 45632
rect 7324 45592 7660 45632
rect 7700 45592 7709 45632
rect 5260 45590 5300 45592
rect 5199 45550 5300 45590
rect 4195 45508 4204 45548
rect 4244 45508 4972 45548
rect 5012 45508 5021 45548
rect 4492 45464 4532 45508
rect 5199 45464 5239 45550
rect 4483 45424 4492 45464
rect 4532 45424 4541 45464
rect 4771 45424 4780 45464
rect 4820 45424 5239 45464
rect 4919 45340 4928 45380
rect 4968 45340 5010 45380
rect 5050 45340 5092 45380
rect 5132 45340 5174 45380
rect 5214 45340 5256 45380
rect 5296 45340 5305 45380
rect 5500 45296 5540 45592
rect 6028 45548 6068 45592
rect 5914 45508 5923 45548
rect 5963 45508 5972 45548
rect 6028 45508 6508 45548
rect 6548 45508 6557 45548
rect 4565 45256 5540 45296
rect 4099 45172 4108 45212
rect 4148 45172 4204 45212
rect 4244 45172 4279 45212
rect 4565 45128 4605 45256
rect 5321 45172 5452 45212
rect 5492 45172 5501 45212
rect 5609 45172 5731 45212
rect 5780 45172 5789 45212
rect 0 45088 1652 45128
rect 3907 45088 3916 45128
rect 3956 45088 4605 45128
rect 0 45068 90 45088
rect 4565 45044 4605 45088
rect 5068 45088 5356 45128
rect 5396 45088 5405 45128
rect 5513 45088 5633 45128
rect 5684 45088 5693 45128
rect 5068 45044 5108 45088
rect 2755 45004 2764 45044
rect 2804 45004 2813 45044
rect 4012 45035 4108 45044
rect 67 44920 76 44960
rect 116 44920 1228 44960
rect 1268 44920 1277 44960
rect 1481 44920 1612 44960
rect 1652 44920 1661 44960
rect 2764 44876 2804 45004
rect 4052 45004 4108 45035
rect 4148 45004 4183 45044
rect 4387 45004 4396 45044
rect 4436 45004 4445 45044
rect 4556 45004 4565 45044
rect 4605 45004 4628 45044
rect 4675 45004 4684 45044
rect 4724 45004 4820 45044
rect 5059 45004 5068 45044
rect 5108 45004 5117 45044
rect 5164 45004 5190 45044
rect 5230 45004 5239 45044
rect 5407 45035 5452 45044
rect 4012 44986 4052 44995
rect 4396 44960 4436 45004
rect 4588 44960 4628 45004
rect 4204 44920 4492 44960
rect 4532 44920 4541 44960
rect 4588 44920 4684 44960
rect 4724 44920 4733 44960
rect 4204 44876 4244 44920
rect 2563 44836 2572 44876
rect 2612 44836 2900 44876
rect 4195 44836 4204 44876
rect 4244 44836 4253 44876
rect 0 44792 90 44812
rect 0 44752 76 44792
rect 116 44752 125 44792
rect 1337 44752 1420 44792
rect 1460 44752 1468 44792
rect 1508 44752 1517 44792
rect 1843 44752 1852 44792
rect 1892 44752 2380 44792
rect 2420 44752 2429 44792
rect 0 44732 90 44752
rect 2860 44708 2900 44836
rect 4780 44792 4820 45004
rect 5164 44960 5204 45004
rect 4876 44920 5204 44960
rect 5305 45002 5345 45011
rect 5447 45004 5452 45035
rect 5492 45004 5578 45044
rect 5827 45004 5836 45044
rect 5876 45004 5885 45044
rect 5932 45035 5972 45508
rect 7756 45464 7796 45676
rect 7651 45424 7660 45464
rect 7700 45424 7796 45464
rect 7852 45380 7892 45676
rect 8002 45632 8042 45676
rect 9580 45667 9620 45676
rect 8002 45592 8332 45632
rect 8372 45592 8381 45632
rect 9763 45508 9772 45548
rect 9812 45508 9821 45548
rect 6403 45340 6412 45380
rect 6452 45340 6892 45380
rect 6932 45340 6941 45380
rect 7555 45340 7564 45380
rect 7604 45340 7892 45380
rect 9772 45380 9812 45508
rect 9964 45464 10004 45676
rect 11212 45667 11252 45676
rect 11980 45632 12020 45676
rect 13228 45667 13268 45676
rect 14284 45632 14324 45676
rect 11491 45592 11500 45632
rect 11540 45592 12020 45632
rect 13891 45592 13900 45632
rect 13940 45592 14324 45632
rect 15244 45548 15284 45676
rect 15916 45592 17260 45632
rect 17300 45592 17309 45632
rect 15916 45548 15956 45592
rect 15244 45508 15340 45548
rect 15380 45508 15389 45548
rect 15907 45508 15916 45548
rect 15956 45508 15965 45548
rect 17299 45508 17308 45548
rect 17348 45508 17740 45548
rect 17780 45508 17789 45548
rect 9964 45424 14572 45464
rect 14612 45424 15244 45464
rect 15284 45424 15293 45464
rect 9772 45340 11636 45380
rect 6211 45256 6220 45296
rect 6260 45256 6700 45296
rect 6740 45256 7084 45296
rect 7124 45256 7133 45296
rect 7939 45256 7948 45296
rect 7988 45256 9332 45296
rect 6019 45172 6028 45212
rect 6068 45172 6892 45212
rect 6932 45172 6941 45212
rect 8131 45172 8140 45212
rect 8180 45172 9196 45212
rect 9236 45172 9245 45212
rect 9292 45128 9332 45256
rect 10435 45172 10444 45212
rect 10484 45172 10636 45212
rect 10676 45172 11156 45212
rect 11203 45172 11212 45212
rect 11252 45172 11261 45212
rect 11116 45128 11156 45172
rect 6185 45088 6316 45128
rect 6356 45088 6796 45128
rect 6836 45088 6845 45128
rect 6979 45088 6988 45128
rect 7028 45088 7268 45128
rect 7529 45088 7660 45128
rect 7700 45088 7948 45128
rect 7988 45088 7997 45128
rect 8611 45088 8620 45128
rect 8660 45088 8875 45128
rect 7228 45044 7268 45088
rect 7660 45044 7700 45088
rect 8835 45044 8875 45088
rect 9004 45088 9332 45128
rect 10339 45088 10348 45128
rect 10388 45088 10964 45128
rect 9004 45044 9044 45088
rect 5407 44986 5447 44995
rect 4876 44876 4916 44920
rect 5305 44876 5345 44962
rect 4867 44836 4876 44876
rect 4916 44836 4925 44876
rect 5155 44836 5164 44876
rect 5204 44836 5345 44876
rect 5836 44876 5876 45004
rect 6019 45004 6028 45044
rect 6068 45004 6110 45044
rect 6150 45004 6199 45044
rect 6412 45035 6452 45044
rect 5932 44986 5972 44995
rect 6691 45004 6700 45044
rect 6740 45004 6748 45044
rect 6788 45004 6871 45044
rect 6988 45004 7049 45044
rect 7089 45004 7098 45044
rect 7210 45004 7219 45044
rect 7259 45004 7468 45044
rect 7508 45035 7604 45044
rect 7508 45004 7564 45035
rect 6412 44876 6452 44995
rect 6988 44960 7028 45004
rect 7660 45035 7715 45044
rect 7660 45004 7675 45035
rect 7564 44986 7604 44995
rect 7675 44986 7715 44995
rect 7786 45035 7852 45044
rect 7786 44995 7795 45035
rect 7835 45004 7852 45035
rect 7892 45004 7975 45044
rect 8131 45004 8140 45044
rect 8180 45004 8236 45044
rect 8276 45004 8311 45044
rect 8419 45004 8428 45044
rect 8493 45004 8599 45044
rect 8707 45004 8716 45044
rect 8756 45004 8765 45044
rect 8826 45004 8835 45044
rect 8875 45004 8884 45044
rect 8944 45004 8953 45044
rect 8993 45004 9044 45044
rect 9187 45004 9196 45044
rect 9236 45004 9245 45044
rect 10147 45004 10156 45044
rect 10196 45035 10484 45044
rect 10196 45004 10444 45035
rect 7835 44995 7844 45004
rect 7786 44994 7844 44995
rect 6761 44920 6892 44960
rect 6932 44920 6941 44960
rect 6988 44920 7276 44960
rect 7316 44920 7325 44960
rect 8362 44951 8620 44960
rect 8362 44911 8371 44951
rect 8411 44920 8620 44951
rect 8660 44920 8669 44960
rect 8411 44911 8420 44920
rect 8362 44910 8420 44911
rect 5836 44836 6700 44876
rect 6740 44836 6749 44876
rect 6979 44836 6988 44876
rect 7028 44836 7180 44876
rect 7220 44836 7229 44876
rect 8716 44792 8756 45004
rect 9196 44960 9236 45004
rect 10697 45004 10819 45044
rect 10868 45004 10877 45044
rect 10924 45035 10964 45088
rect 11098 45119 11156 45128
rect 11098 45079 11107 45119
rect 11147 45079 11156 45119
rect 11098 45078 11156 45079
rect 11212 45044 11252 45172
rect 11596 45128 11636 45340
rect 15148 45256 16492 45296
rect 16532 45256 16541 45296
rect 11923 45172 11932 45212
rect 11972 45172 15052 45212
rect 15092 45172 15101 45212
rect 15148 45128 15188 45256
rect 17836 45212 17876 45676
rect 18892 45667 18932 45676
rect 21388 45632 21428 45676
rect 19987 45592 19996 45632
rect 20036 45592 21004 45632
rect 21044 45592 21053 45632
rect 21388 45592 21484 45632
rect 21524 45592 21533 45632
rect 19555 45508 19564 45548
rect 19604 45508 19613 45548
rect 20371 45508 20380 45548
rect 20420 45508 20948 45548
rect 19564 45464 19604 45508
rect 19564 45424 20524 45464
rect 20564 45424 20573 45464
rect 20039 45340 20048 45380
rect 20088 45340 20130 45380
rect 20170 45340 20212 45380
rect 20252 45340 20294 45380
rect 20334 45340 20376 45380
rect 20416 45340 20425 45380
rect 20908 45296 20948 45508
rect 21510 45296 21600 45316
rect 20908 45256 21600 45296
rect 21510 45236 21600 45256
rect 15235 45172 15244 45212
rect 15284 45172 15293 45212
rect 17443 45172 17452 45212
rect 17492 45172 17876 45212
rect 18403 45172 18412 45212
rect 18452 45172 18461 45212
rect 18883 45172 18892 45212
rect 18932 45172 19756 45212
rect 19796 45172 19805 45212
rect 11500 45088 11636 45128
rect 12940 45088 15188 45128
rect 15244 45128 15284 45172
rect 18412 45128 18452 45172
rect 15244 45088 17588 45128
rect 18412 45088 18644 45128
rect 11500 45044 11540 45088
rect 10444 44960 10484 44995
rect 11190 45004 11199 45044
rect 11239 45004 11252 45044
rect 11371 45004 11380 45044
rect 11420 45004 11540 45044
rect 10924 44986 10964 44995
rect 12940 44960 12980 45088
rect 13355 45004 13420 45044
rect 13460 45004 13486 45044
rect 13526 45004 13535 45044
rect 13608 45004 13617 45044
rect 13657 45004 13699 45044
rect 13891 45004 13900 45044
rect 13940 45004 13996 45044
rect 14036 45004 14071 45044
rect 14412 45004 14476 45044
rect 14516 45035 14612 45044
rect 14516 45004 14572 45035
rect 13612 44960 13652 45004
rect 14921 45004 15052 45044
rect 15092 45004 15101 45044
rect 16003 45004 16012 45044
rect 16052 45004 16061 45044
rect 17129 45004 17260 45044
rect 17300 45004 17309 45044
rect 14572 44960 14612 44995
rect 15052 44986 15092 44995
rect 16012 44960 16052 45004
rect 17260 44986 17300 44995
rect 8899 44920 8908 44960
rect 8948 44920 9292 44960
rect 9332 44920 9396 44960
rect 10444 44920 10636 44960
rect 10676 44920 10685 44960
rect 11491 44920 11500 44960
rect 11540 44920 11692 44960
rect 11732 44920 11741 44960
rect 12643 44920 12652 44960
rect 12692 44920 12980 44960
rect 13603 44920 13612 44960
rect 13652 44920 13661 44960
rect 14057 44920 14092 44960
rect 14132 44920 14188 44960
rect 14228 44920 14237 44960
rect 14572 44920 14860 44960
rect 14900 44920 14909 44960
rect 15715 44920 15724 44960
rect 15764 44920 16052 44960
rect 15724 44876 15764 44920
rect 4780 44752 5932 44792
rect 5972 44752 5981 44792
rect 6106 44752 6115 44792
rect 6155 44752 6316 44792
rect 6356 44752 6365 44792
rect 7939 44752 7948 44792
rect 7988 44752 8756 44792
rect 9004 44836 15764 44876
rect 17548 44876 17588 45088
rect 17635 45004 17644 45044
rect 17684 45004 18019 45044
rect 18059 45004 18068 45044
rect 18115 45004 18124 45044
rect 18164 45004 18295 45044
rect 18377 45004 18412 45044
rect 18452 45004 18508 45044
rect 18548 45004 18557 45044
rect 18604 44960 18644 45088
rect 18924 45004 18988 45044
rect 19028 45035 19276 45044
rect 19028 45004 19084 45035
rect 19124 45004 19276 45035
rect 19316 45004 19325 45044
rect 19564 45035 20140 45044
rect 19084 44986 19124 44995
rect 19604 45004 20140 45035
rect 20180 45004 20189 45044
rect 19564 44986 19604 44995
rect 18595 44920 18604 44960
rect 18644 44920 18653 44960
rect 20131 44920 20140 44960
rect 20180 44920 21292 44960
rect 21332 44920 21341 44960
rect 17548 44836 19948 44876
rect 19988 44836 19997 44876
rect 9004 44708 9044 44836
rect 21510 44792 21600 44812
rect 10810 44752 10819 44792
rect 10859 44752 11212 44792
rect 11252 44752 11261 44792
rect 12403 44752 12412 44792
rect 12452 44752 12844 44792
rect 12884 44752 12893 44792
rect 15475 44752 15484 44792
rect 15524 44752 16204 44792
rect 16244 44752 16253 44792
rect 20371 44752 20380 44792
rect 20420 44752 21600 44792
rect 21510 44732 21600 44752
rect 2860 44668 9044 44708
rect 10819 44668 10828 44708
rect 10868 44668 19564 44708
rect 19604 44668 19613 44708
rect 3679 44584 3688 44624
rect 3728 44584 3770 44624
rect 3810 44584 3852 44624
rect 3892 44584 3934 44624
rect 3974 44584 4016 44624
rect 4056 44584 4065 44624
rect 4300 44584 8660 44624
rect 8707 44584 8716 44624
rect 8756 44584 11308 44624
rect 11348 44584 11500 44624
rect 11540 44584 11549 44624
rect 18799 44584 18808 44624
rect 18848 44584 18890 44624
rect 18930 44584 18972 44624
rect 19012 44584 19054 44624
rect 19094 44584 19136 44624
rect 19176 44584 19185 44624
rect 1708 44500 4148 44540
rect 0 44456 90 44476
rect 0 44416 1612 44456
rect 1652 44416 1661 44456
rect 0 44396 90 44416
rect 1708 44372 1748 44500
rect 1843 44416 1852 44456
rect 1892 44416 4012 44456
rect 4052 44416 4061 44456
rect 4108 44372 4148 44500
rect 1459 44332 1468 44372
rect 1508 44332 1748 44372
rect 3907 44332 3916 44372
rect 3956 44332 4148 44372
rect 67 44248 76 44288
rect 116 44248 1228 44288
rect 1268 44248 1277 44288
rect 1603 44248 1612 44288
rect 1652 44248 1661 44288
rect 2851 44248 2860 44288
rect 2900 44248 3052 44288
rect 3092 44248 3101 44288
rect 3436 44248 4204 44288
rect 4244 44248 4253 44288
rect 0 44120 90 44140
rect 0 44080 76 44120
rect 116 44080 125 44120
rect 0 44060 90 44080
rect 1612 43868 1652 44248
rect 3436 44204 3476 44248
rect 2362 44164 2371 44204
rect 2411 44164 2420 44204
rect 2467 44164 2476 44204
rect 2516 44164 2647 44204
rect 2947 44164 2956 44204
rect 2996 44164 3005 44204
rect 3276 44164 3340 44204
rect 3380 44164 3436 44204
rect 3523 44164 3532 44204
rect 3572 44164 3924 44204
rect 3964 44164 3973 44204
rect 2380 44120 2420 44164
rect 2956 44120 2996 44164
rect 3436 44155 3476 44164
rect 2380 44080 2668 44120
rect 2708 44080 2717 44120
rect 2956 44080 3244 44120
rect 3284 44080 3293 44120
rect 3427 43996 3436 44036
rect 3476 43996 4108 44036
rect 4148 43996 4157 44036
rect 4300 43952 4340 44584
rect 4684 44500 6028 44540
rect 6068 44500 6077 44540
rect 6691 44500 6700 44540
rect 6740 44500 6884 44540
rect 4684 44456 4724 44500
rect 6844 44456 6884 44500
rect 8620 44456 8660 44584
rect 9379 44500 9388 44540
rect 9428 44500 9868 44540
rect 9908 44500 9917 44540
rect 14179 44500 14188 44540
rect 14228 44500 19276 44540
rect 19316 44500 19325 44540
rect 4666 44416 4675 44456
rect 4715 44416 4724 44456
rect 4972 44416 5260 44456
rect 5300 44416 5309 44456
rect 5356 44416 5452 44456
rect 5492 44416 5501 44456
rect 5548 44416 6604 44456
rect 6644 44416 6653 44456
rect 6835 44416 6844 44456
rect 6884 44416 6893 44456
rect 7145 44416 7180 44456
rect 7220 44416 7276 44456
rect 7316 44416 7325 44456
rect 8620 44416 11164 44456
rect 11204 44416 11213 44456
rect 13289 44416 13420 44456
rect 13460 44416 13469 44456
rect 14921 44416 15052 44456
rect 15092 44416 15101 44456
rect 17513 44416 17644 44456
rect 17684 44416 17693 44456
rect 18019 44416 18028 44456
rect 18068 44416 18172 44456
rect 18212 44416 18221 44456
rect 20009 44416 20140 44456
rect 20180 44416 20189 44456
rect 4972 44372 5012 44416
rect 5356 44372 5396 44416
rect 5548 44372 5588 44416
rect 4460 44363 4492 44372
rect 4532 44332 4631 44372
rect 4876 44332 5012 44372
rect 5059 44332 5068 44372
rect 5108 44332 5396 44372
rect 5500 44332 5588 44372
rect 5731 44332 5740 44372
rect 5780 44332 6124 44372
rect 6164 44332 6173 44372
rect 6499 44332 6508 44372
rect 6548 44332 11548 44372
rect 11588 44332 13652 44372
rect 15881 44332 15916 44372
rect 15956 44332 16012 44372
rect 16052 44332 16061 44372
rect 16483 44332 16492 44372
rect 16532 44332 17876 44372
rect 4460 44314 4500 44323
rect 4876 44288 4916 44332
rect 4745 44248 4876 44288
rect 4916 44248 4925 44288
rect 5020 44248 5260 44288
rect 5300 44248 5309 44288
rect 4876 44204 4916 44248
rect 5020 44246 5060 44248
rect 5500 44246 5540 44332
rect 5923 44248 5932 44288
rect 5972 44248 6220 44288
rect 6260 44248 6269 44288
rect 6403 44248 6412 44288
rect 6452 44248 6980 44288
rect 9641 44248 9763 44288
rect 9812 44248 9821 44288
rect 10339 44248 10348 44288
rect 10388 44248 10540 44288
rect 10580 44248 10589 44288
rect 11299 44248 11308 44288
rect 11348 44248 11404 44288
rect 11444 44248 11479 44288
rect 11657 44248 11788 44288
rect 11828 44248 11837 44288
rect 5015 44237 5060 44246
rect 172 43828 1652 43868
rect 2860 43912 4340 43952
rect 4396 44164 4483 44204
rect 4523 44164 4684 44204
rect 4724 44164 4733 44204
rect 4876 44164 4915 44204
rect 4955 44164 4964 44204
rect 5055 44206 5060 44237
rect 5470 44206 5479 44246
rect 5519 44206 5540 44246
rect 5689 44237 5735 44246
rect 5689 44204 5695 44237
rect 5015 44188 5055 44197
rect 5347 44164 5356 44204
rect 5396 44164 5405 44204
rect 5584 44164 5593 44204
rect 5633 44164 5642 44204
rect 5687 44197 5695 44204
rect 6940 44204 6980 44248
rect 8812 44204 8852 44213
rect 13228 44204 13268 44213
rect 13612 44204 13652 44332
rect 17836 44288 17876 44332
rect 21510 44288 21600 44308
rect 17827 44248 17836 44288
rect 17876 44248 17885 44288
rect 18281 44248 18412 44288
rect 18452 44248 18461 44288
rect 20995 44248 21004 44288
rect 21044 44248 21600 44288
rect 21510 44228 21600 44248
rect 14860 44204 14900 44213
rect 17452 44204 17492 44213
rect 19948 44204 19988 44213
rect 5687 44188 5735 44197
rect 5687 44164 5729 44188
rect 5836 44164 5884 44204
rect 5924 44164 5933 44204
rect 6210 44164 6316 44204
rect 6381 44164 6390 44204
rect 4396 43952 4436 44164
rect 5356 44120 5396 44164
rect 5596 44120 5636 44164
rect 4684 44080 5396 44120
rect 5443 44080 5452 44120
rect 5492 44080 5636 44120
rect 4684 44036 4724 44080
rect 4675 43996 4684 44036
rect 4724 43996 4733 44036
rect 5033 43996 5164 44036
rect 5204 43996 5213 44036
rect 5687 43952 5727 44164
rect 5836 44120 5876 44164
rect 6047 44122 6056 44162
rect 6096 44122 6164 44162
rect 6496 44137 6505 44177
rect 6545 44137 6554 44177
rect 6700 44164 6709 44204
rect 6749 44164 6788 44204
rect 6931 44164 6940 44204
rect 6980 44164 6989 44204
rect 7171 44164 7180 44204
rect 7220 44164 7321 44204
rect 7363 44164 7372 44204
rect 7412 44164 7421 44204
rect 7555 44164 7564 44204
rect 7604 44164 8236 44204
rect 8276 44164 8285 44204
rect 8777 44164 8812 44204
rect 8852 44164 8908 44204
rect 8948 44164 8957 44204
rect 9065 44164 9187 44204
rect 9236 44164 9245 44204
rect 9634 44164 9643 44204
rect 9683 44164 9716 44204
rect 9859 44164 9868 44204
rect 9908 44164 10039 44204
rect 11971 44164 11980 44204
rect 12020 44164 12029 44204
rect 13603 44164 13612 44204
rect 13652 44164 13661 44204
rect 15043 44164 15052 44204
rect 15092 44164 15340 44204
rect 15380 44164 15389 44204
rect 15497 44164 15619 44204
rect 15668 44164 15677 44204
rect 16073 44164 16204 44204
rect 16244 44164 16253 44204
rect 17731 44164 17740 44204
rect 17780 44164 17932 44204
rect 17972 44164 18700 44204
rect 18740 44164 18749 44204
rect 5836 44080 5932 44120
rect 5972 44080 5981 44120
rect 4396 43912 5727 43952
rect 0 43784 90 43804
rect 172 43784 212 43828
rect 2860 43784 2900 43912
rect 0 43744 212 43784
rect 1219 43744 1228 43784
rect 1268 43744 2900 43784
rect 0 43724 90 43744
rect 4396 43700 4436 43912
rect 4919 43828 4928 43868
rect 4968 43828 5010 43868
rect 5050 43828 5092 43868
rect 5132 43828 5174 43868
rect 5214 43828 5256 43868
rect 5296 43828 5305 43868
rect 5347 43828 5356 43868
rect 5396 43828 5405 43868
rect 5356 43784 5396 43828
rect 4483 43744 4492 43784
rect 4532 43744 5012 43784
rect 1459 43660 1468 43700
rect 1508 43660 2764 43700
rect 2804 43660 2813 43700
rect 3907 43660 3916 43700
rect 3956 43660 4916 43700
rect 2092 43576 4204 43616
rect 4244 43576 4253 43616
rect 0 43448 90 43468
rect 2092 43448 2132 43576
rect 4876 43532 4916 43660
rect 2467 43492 2476 43532
rect 2516 43492 3628 43532
rect 3668 43492 3677 43532
rect 3724 43523 4108 43532
rect 3764 43492 4108 43523
rect 4148 43492 4157 43532
rect 4577 43492 4586 43532
rect 4626 43492 4635 43532
rect 4858 43492 4867 43532
rect 4907 43492 4916 43532
rect 4972 43532 5012 43744
rect 5068 43744 5396 43784
rect 5068 43700 5108 43744
rect 6124 43700 6164 44122
rect 6508 44036 6548 44137
rect 6748 44120 6788 44164
rect 6691 44080 6700 44120
rect 6740 44080 6788 44120
rect 7281 44036 7321 44164
rect 7372 44120 7412 44164
rect 8812 44155 8852 44164
rect 9676 44120 9716 44164
rect 11980 44120 12020 44164
rect 7372 44080 7948 44120
rect 7988 44080 7997 44120
rect 9257 44080 9388 44120
rect 9428 44080 9437 44120
rect 9489 44080 9498 44120
rect 9538 44080 9547 44120
rect 9676 44080 10100 44120
rect 11155 44080 11164 44120
rect 11204 44080 12020 44120
rect 13228 44120 13268 44164
rect 14860 44120 14900 44164
rect 17452 44120 17492 44164
rect 19948 44120 19988 44164
rect 13228 44080 14900 44120
rect 15715 44080 15724 44120
rect 15764 44080 15773 44120
rect 17452 44080 17644 44120
rect 17684 44080 19988 44120
rect 9498 44036 9538 44080
rect 6508 43996 7180 44036
rect 7220 43996 7229 44036
rect 7281 43996 7468 44036
rect 7508 43996 8332 44036
rect 8372 43996 9004 44036
rect 9044 43996 9053 44036
rect 9274 43996 9283 44036
rect 9323 43996 9332 44036
rect 9498 43996 9955 44036
rect 9995 43996 10004 44036
rect 9292 43952 9332 43996
rect 10060 43952 10100 44080
rect 10243 43996 10252 44036
rect 10292 43996 10300 44036
rect 10340 43996 10423 44036
rect 9292 43912 10388 43952
rect 6787 43828 6796 43868
rect 6836 43828 9868 43868
rect 9908 43828 9917 43868
rect 10348 43700 10388 43912
rect 13228 43868 13268 44080
rect 14860 44036 14900 44080
rect 14860 43996 14956 44036
rect 14996 43996 15005 44036
rect 15724 43868 15764 44080
rect 18067 43996 18076 44036
rect 18116 43996 18316 44036
rect 18356 43996 18365 44036
rect 13084 43828 13268 43868
rect 14275 43828 14284 43868
rect 14324 43828 18124 43868
rect 18164 43828 18173 43868
rect 20039 43828 20048 43868
rect 20088 43828 20130 43868
rect 20170 43828 20212 43868
rect 20252 43828 20294 43868
rect 20334 43828 20376 43868
rect 20416 43828 20425 43868
rect 10588 43744 12844 43784
rect 12884 43744 12893 43784
rect 5059 43660 5068 43700
rect 5108 43660 5117 43700
rect 5914 43660 5923 43700
rect 5963 43660 6164 43700
rect 8105 43660 8236 43700
rect 8276 43660 8285 43700
rect 10339 43660 10348 43700
rect 10388 43660 10397 43700
rect 5251 43576 5260 43616
rect 5300 43576 5439 43616
rect 5816 43576 5825 43616
rect 5876 43576 5996 43616
rect 6124 43576 6700 43616
rect 6740 43576 6749 43616
rect 8707 43576 8716 43616
rect 8756 43576 8908 43616
rect 8948 43576 10196 43616
rect 5399 43532 5439 43576
rect 4972 43492 5164 43532
rect 5204 43492 5213 43532
rect 5390 43492 5399 43532
rect 5439 43492 5448 43532
rect 5491 43492 5500 43532
rect 5540 43492 5549 43532
rect 5635 43492 5644 43532
rect 5684 43492 5740 43532
rect 5780 43492 5815 43532
rect 5897 43492 6028 43532
rect 6068 43492 6077 43532
rect 6124 43523 6164 43576
rect 10156 43532 10196 43576
rect 10588 43532 10628 43744
rect 13084 43700 13124 43828
rect 21510 43784 21600 43804
rect 13219 43744 13228 43784
rect 13268 43744 19124 43784
rect 12451 43660 12460 43700
rect 12500 43660 12652 43700
rect 12692 43660 12701 43700
rect 13075 43660 13084 43700
rect 13124 43660 13133 43700
rect 14188 43660 15052 43700
rect 15092 43660 15101 43700
rect 11020 43576 12172 43616
rect 12212 43576 12221 43616
rect 11020 43532 11060 43576
rect 14188 43532 14228 43660
rect 15436 43616 15476 43744
rect 16147 43660 16156 43700
rect 16196 43660 16780 43700
rect 16820 43660 16829 43700
rect 14323 43576 14332 43616
rect 14372 43576 14804 43616
rect 15427 43576 15436 43616
rect 15476 43576 15485 43616
rect 17731 43576 17740 43616
rect 17780 43576 18068 43616
rect 14764 43532 14804 43576
rect 18028 43532 18068 43576
rect 19084 43532 19124 43744
rect 20380 43744 21600 43784
rect 20380 43700 20420 43744
rect 21510 43724 21600 43744
rect 19625 43660 19756 43700
rect 19796 43660 19805 43700
rect 20371 43660 20380 43700
rect 20420 43660 20429 43700
rect 3724 43474 3764 43483
rect 4300 43450 4348 43490
rect 4388 43450 4397 43490
rect 4300 43448 4340 43450
rect 0 43408 1228 43448
rect 1268 43408 1277 43448
rect 1603 43408 1612 43448
rect 1652 43408 1661 43448
rect 2083 43408 2092 43448
rect 2132 43408 2141 43448
rect 4003 43408 4012 43448
rect 4052 43408 4340 43448
rect 4474 43408 4483 43448
rect 4523 43408 4532 43448
rect 0 43388 90 43408
rect 0 43112 90 43132
rect 1612 43112 1652 43408
rect 2179 43324 2188 43364
rect 2228 43324 2332 43364
rect 2372 43324 2381 43364
rect 1843 43240 1852 43280
rect 1892 43240 2092 43280
rect 2132 43240 2141 43280
rect 0 43072 1652 43112
rect 3679 43072 3688 43112
rect 3728 43072 3770 43112
rect 3810 43072 3852 43112
rect 3892 43072 3934 43112
rect 3974 43072 4016 43112
rect 4056 43072 4065 43112
rect 0 43052 90 43072
rect 4492 42860 4532 43408
rect 4588 43364 4628 43492
rect 5500 43448 5540 43492
rect 6490 43492 6499 43532
rect 6539 43492 6548 43532
rect 6595 43492 6604 43532
rect 6644 43492 6653 43532
rect 6857 43492 6988 43532
rect 7028 43492 7037 43532
rect 7564 43523 7756 43532
rect 6124 43474 6164 43483
rect 6508 43448 6548 43492
rect 4675 43408 4684 43448
rect 4724 43408 5540 43448
rect 6461 43408 6508 43448
rect 6548 43408 6557 43448
rect 6604 43364 6644 43492
rect 7604 43492 7756 43523
rect 7796 43492 7805 43532
rect 7939 43492 7948 43532
rect 7988 43523 8119 43532
rect 7988 43492 8044 43523
rect 7564 43474 7604 43483
rect 8084 43492 8119 43523
rect 8899 43492 8908 43532
rect 8948 43492 9292 43532
rect 9332 43492 9341 43532
rect 10156 43523 10628 43532
rect 8044 43474 8084 43483
rect 10196 43492 10628 43523
rect 10723 43492 10732 43532
rect 10772 43492 10915 43532
rect 10955 43492 10964 43532
rect 11011 43492 11020 43532
rect 11060 43492 11191 43532
rect 11273 43492 11404 43532
rect 11444 43492 11453 43532
rect 11980 43523 12364 43532
rect 10156 43474 10196 43483
rect 12020 43492 12364 43523
rect 12404 43492 12413 43532
rect 12460 43523 12500 43532
rect 11980 43474 12020 43483
rect 14179 43492 14188 43532
rect 14228 43492 14237 43532
rect 14441 43492 14572 43532
rect 14612 43492 14621 43532
rect 14764 43492 14809 43532
rect 14849 43492 14996 43532
rect 15043 43492 15052 43532
rect 15092 43492 15223 43532
rect 15322 43492 15331 43532
rect 15380 43492 15511 43532
rect 16291 43492 16300 43532
rect 16340 43492 16416 43532
rect 17251 43492 17260 43532
rect 17300 43523 17588 43532
rect 17300 43492 17548 43523
rect 6953 43408 7084 43448
rect 7124 43408 7133 43448
rect 11369 43408 11500 43448
rect 11540 43408 11549 43448
rect 12460 43364 12500 43483
rect 14956 43448 14996 43492
rect 16300 43448 16340 43492
rect 18010 43492 18019 43532
rect 18059 43492 18068 43532
rect 18115 43492 18124 43532
rect 18164 43492 18295 43532
rect 18499 43492 18508 43532
rect 18548 43492 18679 43532
rect 19084 43523 19276 43532
rect 12713 43408 12844 43448
rect 12884 43408 12893 43448
rect 13289 43408 13420 43448
rect 13460 43408 13469 43448
rect 14345 43408 14476 43448
rect 14516 43408 14525 43448
rect 14668 43408 14691 43448
rect 14731 43408 14740 43448
rect 14956 43408 15628 43448
rect 15668 43408 15677 43448
rect 15907 43408 15916 43448
rect 15956 43408 16300 43448
rect 16340 43408 16349 43448
rect 14668 43364 14708 43408
rect 17548 43364 17588 43483
rect 19124 43492 19276 43523
rect 19316 43492 19325 43532
rect 19433 43492 19564 43532
rect 19604 43492 19613 43532
rect 19084 43474 19124 43483
rect 19564 43474 19604 43483
rect 18473 43408 18604 43448
rect 18644 43408 18653 43448
rect 20131 43408 20140 43448
rect 20180 43408 20524 43448
rect 20564 43408 20573 43448
rect 4588 43324 4972 43364
rect 5012 43324 5021 43364
rect 5251 43324 5260 43364
rect 5300 43324 6644 43364
rect 11395 43324 11404 43364
rect 11444 43324 12500 43364
rect 13027 43324 13036 43364
rect 13076 43324 13180 43364
rect 13220 43324 13229 43364
rect 13699 43324 13708 43364
rect 13748 43324 14188 43364
rect 14228 43324 14708 43364
rect 15331 43324 15340 43364
rect 15380 43324 15389 43364
rect 15715 43324 15724 43364
rect 15764 43324 16108 43364
rect 16148 43324 16157 43364
rect 17548 43324 18700 43364
rect 18740 43324 18749 43364
rect 15340 43280 15380 43324
rect 21510 43280 21600 43300
rect 4771 43240 4780 43280
rect 4820 43240 5356 43280
rect 5396 43240 5405 43280
rect 9859 43240 9868 43280
rect 9908 43240 11788 43280
rect 11828 43240 11837 43280
rect 14371 43240 14380 43280
rect 14420 43240 15380 43280
rect 21388 43240 21600 43280
rect 6700 43156 11116 43196
rect 11156 43156 11165 43196
rect 12835 43156 12844 43196
rect 12884 43156 15052 43196
rect 15092 43156 15101 43196
rect 6700 43028 6740 43156
rect 15052 43112 15092 43156
rect 6307 42988 6316 43028
rect 6356 42988 6740 43028
rect 6796 43072 11500 43112
rect 11540 43072 11549 43112
rect 13315 43072 13324 43112
rect 13364 43072 14996 43112
rect 15052 43072 15436 43112
rect 15476 43072 15485 43112
rect 18799 43072 18808 43112
rect 18848 43072 18890 43112
rect 18930 43072 18972 43112
rect 19012 43072 19054 43112
rect 19094 43072 19136 43112
rect 19176 43072 19185 43112
rect 6796 42944 6836 43072
rect 14956 43028 14996 43072
rect 14956 42988 17684 43028
rect 4579 42904 4588 42944
rect 4628 42904 4684 42944
rect 4724 42904 4759 42944
rect 4963 42904 4972 42944
rect 5012 42904 5347 42944
rect 5387 42904 5396 42944
rect 5801 42904 5932 42944
rect 5972 42904 5981 42944
rect 6115 42904 6124 42944
rect 6164 42904 6836 42944
rect 8995 42904 9004 42944
rect 9044 42904 9772 42944
rect 9812 42904 9821 42944
rect 11971 42904 11980 42944
rect 12020 42904 12892 42944
rect 12932 42904 12941 42944
rect 15619 42904 15628 42944
rect 15668 42904 16148 42944
rect 1027 42820 1036 42860
rect 1076 42820 2236 42860
rect 2276 42820 2285 42860
rect 4003 42820 4012 42860
rect 4052 42820 4532 42860
rect 5155 42820 5164 42860
rect 5204 42820 5335 42860
rect 6019 42820 6028 42860
rect 6068 42820 6740 42860
rect 0 42776 90 42796
rect 4492 42776 4532 42820
rect 0 42736 1228 42776
rect 1268 42736 1277 42776
rect 1603 42736 1612 42776
rect 1652 42736 1661 42776
rect 1987 42736 1996 42776
rect 2036 42736 2045 42776
rect 4099 42736 4108 42776
rect 4148 42736 4157 42776
rect 4492 42736 5684 42776
rect 0 42716 90 42736
rect 1612 42608 1652 42736
rect 1996 42692 2036 42736
rect 3820 42692 3860 42701
rect 4108 42692 4148 42736
rect 4492 42692 4532 42736
rect 4972 42692 5012 42736
rect 5644 42692 5684 42736
rect 6316 42736 6508 42776
rect 6548 42736 6557 42776
rect 6316 42692 6356 42736
rect 6700 42692 6740 42820
rect 6796 42776 6836 42904
rect 7468 42820 15956 42860
rect 6787 42736 6796 42776
rect 6836 42736 6845 42776
rect 7372 42692 7412 42701
rect 1996 42652 2132 42692
rect 2563 42652 2572 42692
rect 2612 42652 3148 42692
rect 3188 42652 3197 42692
rect 3860 42652 4148 42692
rect 4195 42652 4204 42692
rect 4244 42652 4253 42692
rect 4483 42652 4492 42692
rect 4532 42652 4541 42692
rect 4675 42652 4684 42692
rect 4724 42652 4855 42692
rect 4963 42652 4972 42692
rect 5012 42652 5021 42692
rect 5336 42652 5345 42692
rect 5396 42652 5516 42692
rect 5635 42652 5644 42692
rect 5684 42652 5836 42692
rect 5876 42652 5885 42692
rect 5993 42652 6028 42692
rect 6068 42652 6124 42692
rect 6164 42652 6173 42692
rect 6298 42652 6307 42692
rect 6347 42652 6356 42692
rect 6403 42652 6412 42692
rect 6452 42652 6583 42692
rect 6700 42652 6892 42692
rect 6932 42652 6941 42692
rect 172 42568 1652 42608
rect 1795 42568 1804 42608
rect 1844 42568 1852 42608
rect 1892 42568 1975 42608
rect 0 42440 90 42460
rect 172 42440 212 42568
rect 1459 42484 1468 42524
rect 1508 42484 1708 42524
rect 1748 42484 1757 42524
rect 0 42400 212 42440
rect 0 42380 90 42400
rect 2092 42356 2132 42652
rect 3820 42643 3860 42652
rect 4204 42608 4244 42652
rect 5644 42643 5684 42652
rect 6412 42608 6452 42652
rect 7372 42608 7412 42652
rect 4204 42568 5260 42608
rect 5300 42568 5309 42608
rect 6019 42568 6028 42608
rect 6068 42568 6452 42608
rect 6883 42568 6892 42608
rect 6932 42568 7412 42608
rect 4204 42524 4244 42568
rect 2467 42484 2476 42524
rect 2516 42484 4244 42524
rect 4339 42484 4348 42524
rect 4388 42484 4684 42524
rect 4724 42484 4733 42524
rect 4858 42484 4867 42524
rect 4907 42484 4916 42524
rect 5539 42484 5548 42524
rect 5588 42484 6988 42524
rect 7028 42484 7037 42524
rect 4876 42440 4916 42484
rect 4876 42400 6892 42440
rect 6932 42400 6941 42440
rect 7468 42356 7508 42820
rect 8227 42736 8236 42776
rect 8276 42736 8756 42776
rect 12643 42736 12652 42776
rect 12692 42736 13132 42776
rect 13172 42736 13181 42776
rect 13795 42736 13804 42776
rect 13844 42736 13891 42776
rect 15427 42736 15436 42776
rect 15476 42736 15523 42776
rect 15563 42736 15607 42776
rect 8716 42692 8756 42736
rect 10924 42692 10964 42701
rect 12556 42692 12596 42701
rect 13804 42692 13844 42736
rect 15052 42692 15092 42701
rect 15916 42692 15956 42820
rect 16108 42692 16148 42904
rect 17644 42776 17684 42988
rect 21388 42944 21428 43240
rect 21510 43220 21600 43240
rect 20371 42904 20380 42944
rect 20420 42904 21428 42944
rect 21510 42776 21600 42796
rect 17644 42736 18508 42776
rect 18548 42736 18557 42776
rect 20131 42736 20140 42776
rect 20180 42736 20189 42776
rect 20515 42736 20524 42776
rect 20564 42736 21600 42776
rect 17548 42692 17588 42701
rect 19084 42692 19124 42701
rect 20140 42692 20180 42736
rect 21510 42716 21600 42736
rect 7817 42652 7891 42692
rect 7931 42652 7948 42692
rect 7988 42652 7997 42692
rect 8201 42652 8332 42692
rect 8372 42652 8381 42692
rect 8428 42652 8587 42692
rect 8627 42652 8636 42692
rect 8698 42652 8707 42692
rect 8747 42652 8756 42692
rect 9667 42652 9676 42692
rect 9716 42652 9868 42692
rect 9908 42652 9917 42692
rect 11177 42652 11212 42692
rect 11252 42652 11308 42692
rect 11348 42652 11357 42692
rect 13193 42652 13315 42692
rect 13364 42652 13373 42692
rect 13795 42652 13804 42692
rect 13844 42652 13853 42692
rect 14179 42652 14188 42692
rect 14228 42652 15052 42692
rect 15235 42652 15244 42692
rect 15284 42652 15383 42692
rect 15423 42652 15432 42692
rect 15619 42652 15628 42692
rect 15668 42652 15799 42692
rect 15907 42652 15916 42692
rect 15956 42652 15965 42692
rect 16099 42652 16108 42692
rect 16148 42652 16157 42692
rect 16291 42652 16300 42692
rect 16340 42652 16471 42692
rect 17588 42652 17684 42692
rect 8428 42608 8468 42652
rect 8044 42568 8468 42608
rect 10924 42608 10964 42652
rect 12556 42608 12596 42652
rect 15052 42643 15092 42652
rect 17548 42643 17588 42652
rect 10924 42568 12596 42608
rect 12739 42568 12748 42608
rect 12788 42568 12980 42608
rect 13617 42568 13626 42608
rect 13666 42568 13804 42608
rect 13844 42568 13853 42608
rect 15614 42568 16148 42608
rect 8044 42524 8084 42568
rect 8035 42484 8044 42524
rect 8084 42484 8093 42524
rect 172 42316 2132 42356
rect 4684 42316 4780 42356
rect 4820 42316 4829 42356
rect 4919 42316 4928 42356
rect 4968 42316 5010 42356
rect 5050 42316 5092 42356
rect 5132 42316 5174 42356
rect 5214 42316 5256 42356
rect 5296 42316 5305 42356
rect 7180 42316 7508 42356
rect 0 42104 90 42124
rect 172 42104 212 42316
rect 4684 42272 4724 42316
rect 7180 42272 7220 42316
rect 10924 42272 10964 42568
rect 12940 42524 12980 42568
rect 11107 42484 11116 42524
rect 11156 42484 11165 42524
rect 12940 42484 13076 42524
rect 13402 42484 13411 42524
rect 13451 42484 13460 42524
rect 13507 42484 13516 42524
rect 13556 42484 14284 42524
rect 14324 42484 14333 42524
rect 15043 42484 15052 42524
rect 15092 42484 15244 42524
rect 15284 42484 15293 42524
rect 0 42064 212 42104
rect 1420 42232 4724 42272
rect 4780 42232 7220 42272
rect 7363 42232 7372 42272
rect 7412 42232 10964 42272
rect 0 42044 90 42064
rect 1420 42020 1460 42232
rect 4780 42188 4820 42232
rect 7180 42188 7220 42232
rect 2947 42148 2956 42188
rect 2996 42148 3292 42188
rect 3332 42148 3341 42188
rect 3619 42148 3628 42188
rect 3668 42148 4820 42188
rect 6979 42148 6988 42188
rect 7028 42148 7220 42188
rect 7939 42148 7948 42188
rect 7988 42148 9100 42188
rect 9140 42148 9149 42188
rect 9868 42148 10444 42188
rect 10484 42148 10493 42188
rect 10601 42148 10732 42188
rect 10772 42148 10781 42188
rect 2851 42064 2860 42104
rect 2900 42064 3532 42104
rect 3572 42064 3581 42104
rect 4963 42064 4972 42104
rect 5012 42064 5300 42104
rect 5260 42020 5300 42064
rect 9868 42020 9908 42148
rect 11116 42020 11156 42484
rect 11203 42400 11212 42440
rect 11252 42400 12940 42440
rect 12980 42400 12989 42440
rect 13036 42272 13076 42484
rect 13420 42440 13460 42484
rect 15614 42440 15654 42568
rect 15706 42484 15715 42524
rect 15755 42484 15820 42524
rect 15860 42484 15895 42524
rect 16003 42484 16012 42524
rect 16052 42484 16061 42524
rect 13420 42400 14476 42440
rect 14516 42400 14525 42440
rect 15052 42400 15654 42440
rect 13027 42232 13036 42272
rect 13076 42232 13085 42272
rect 15052 42188 15092 42400
rect 16012 42356 16052 42484
rect 15772 42316 16052 42356
rect 15772 42272 15812 42316
rect 15532 42232 15812 42272
rect 13219 42148 13228 42188
rect 13268 42148 13420 42188
rect 13460 42148 13469 42188
rect 15043 42148 15052 42188
rect 15092 42148 15101 42188
rect 11779 42064 11788 42104
rect 11828 42064 12020 42104
rect 11980 42020 12020 42064
rect 12940 42064 13036 42104
rect 13076 42064 13085 42104
rect 15292 42064 15436 42104
rect 15476 42064 15485 42104
rect 12940 42020 12980 42064
rect 15292 42020 15332 42064
rect 15532 42020 15572 42232
rect 16108 42188 16148 42568
rect 17644 42524 17684 42652
rect 17740 42652 18019 42692
rect 18059 42652 18068 42692
rect 18115 42652 18124 42692
rect 18164 42652 18295 42692
rect 18473 42652 18604 42692
rect 18644 42652 18653 42692
rect 19124 42652 19276 42692
rect 19316 42652 19325 42692
rect 19372 42652 19572 42692
rect 19612 42652 19621 42692
rect 20140 42652 20812 42692
rect 20852 42652 20861 42692
rect 17740 42608 17780 42652
rect 19084 42643 19124 42652
rect 17731 42568 17740 42608
rect 17780 42568 17789 42608
rect 19372 42524 19412 42652
rect 17644 42484 17836 42524
rect 17876 42484 17885 42524
rect 18028 42484 19412 42524
rect 19747 42484 19756 42524
rect 19796 42484 19805 42524
rect 16195 42232 16204 42272
rect 16244 42232 16291 42272
rect 16204 42188 16244 42232
rect 18028 42188 18068 42484
rect 19756 42272 19796 42484
rect 20039 42316 20048 42356
rect 20088 42316 20130 42356
rect 20170 42316 20212 42356
rect 20252 42316 20294 42356
rect 20334 42316 20376 42356
rect 20416 42316 20425 42356
rect 21510 42272 21600 42292
rect 18124 42232 19796 42272
rect 20611 42232 20620 42272
rect 20660 42232 21600 42272
rect 15619 42148 15628 42188
rect 15668 42148 15677 42188
rect 16012 42148 16148 42188
rect 16195 42148 16204 42188
rect 16244 42148 16253 42188
rect 18019 42148 18028 42188
rect 18068 42148 18077 42188
rect 15628 42104 15668 42148
rect 16012 42104 16052 42148
rect 18124 42104 18164 42232
rect 21510 42212 21600 42232
rect 19555 42148 19564 42188
rect 19604 42148 19660 42188
rect 19700 42148 19735 42188
rect 20371 42148 20380 42188
rect 20420 42148 20524 42188
rect 20564 42148 20573 42188
rect 1411 41980 1420 42020
rect 1460 41980 1469 42020
rect 2467 41980 2476 42020
rect 2516 42011 2708 42020
rect 2516 41980 2668 42011
rect 2851 41980 2860 42020
rect 2900 41980 3476 42020
rect 3523 41980 3532 42020
rect 3572 41980 4588 42020
rect 4628 41980 4637 42020
rect 4780 42011 4820 42020
rect 2668 41962 2708 41971
rect 3436 41936 3476 41980
rect 5242 41980 5251 42020
rect 5291 41980 5300 42020
rect 5347 41980 5356 42020
rect 5396 41980 5443 42020
rect 5731 41980 5740 42020
rect 5780 41980 6220 42020
rect 6260 41980 6269 42020
rect 6316 42011 6356 42020
rect 4780 41936 4820 41971
rect 5356 41936 5396 41980
rect 3017 41896 3052 41936
rect 3092 41896 3148 41936
rect 3188 41896 3197 41936
rect 3436 41896 4820 41936
rect 5347 41896 5356 41936
rect 5396 41896 5405 41936
rect 5635 41896 5644 41936
rect 5684 41896 5836 41936
rect 5876 41896 5932 41936
rect 5972 41896 6036 41936
rect 6316 41852 6356 41971
rect 6796 42011 6836 42020
rect 7651 41980 7660 42020
rect 7700 41980 8428 42020
rect 8468 41980 8477 42020
rect 8707 41980 8716 42020
rect 8756 42011 8948 42020
rect 8756 41980 8908 42011
rect 6796 41936 6836 41971
rect 9283 41980 9292 42020
rect 9332 41980 9868 42020
rect 9908 41980 9917 42020
rect 10060 42011 10636 42020
rect 10060 41980 10540 42011
rect 8908 41962 8948 41971
rect 10060 41936 10100 41980
rect 10580 41980 10636 42011
rect 10676 41980 10685 42020
rect 11116 41980 11491 42020
rect 11531 41980 11540 42020
rect 11587 41980 11596 42020
rect 11636 41980 11683 42020
rect 11971 41980 11980 42020
rect 12020 41980 12029 42020
rect 12451 41980 12460 42020
rect 12500 42011 12631 42020
rect 12500 41980 12556 42011
rect 10540 41962 10580 41971
rect 11596 41936 11636 41980
rect 12596 41980 12631 42011
rect 12940 42011 13076 42020
rect 12940 41980 13036 42011
rect 12556 41962 12596 41971
rect 13411 41980 13420 42020
rect 13460 41980 13469 42020
rect 13699 41980 13708 42020
rect 13748 41980 14188 42020
rect 14228 42011 14708 42020
rect 14228 41980 14668 42011
rect 13036 41962 13076 41971
rect 6796 41896 7948 41936
rect 7988 41896 7997 41936
rect 9763 41896 9772 41936
rect 9812 41896 10100 41936
rect 11587 41896 11596 41936
rect 11636 41896 11645 41936
rect 12067 41896 12076 41936
rect 12116 41896 12125 41936
rect 12076 41852 12116 41896
rect 13420 41852 13460 41980
rect 15017 41980 15052 42020
rect 15092 41980 15148 42020
rect 15188 41980 15197 42020
rect 15274 42011 15332 42020
rect 14668 41962 14708 41971
rect 15274 41971 15283 42011
rect 15323 41971 15332 42011
rect 15376 41980 15385 42020
rect 15425 41980 15572 42020
rect 15614 42064 15668 42104
rect 15992 42064 16001 42104
rect 16041 42064 16052 42104
rect 16099 42064 16108 42104
rect 16148 42064 16340 42104
rect 15614 42020 15654 42064
rect 16300 42020 16340 42064
rect 16396 42064 18164 42104
rect 15614 41980 15627 42020
rect 15667 41980 15676 42020
rect 15811 41980 15820 42020
rect 15885 41980 15991 42020
rect 16300 42011 16342 42020
rect 16300 41980 16302 42011
rect 15274 41970 15332 41971
rect 16302 41962 16342 41971
rect 15401 41896 15436 41936
rect 15476 41896 15532 41936
rect 15572 41896 15581 41936
rect 15754 41927 15812 41936
rect 15754 41887 15763 41927
rect 15803 41887 15812 41927
rect 15754 41886 15812 41887
rect 15772 41852 15812 41886
rect 16396 41852 16436 42064
rect 16553 41980 16588 42020
rect 16628 41980 16684 42020
rect 16724 41980 16733 42020
rect 17705 41980 17836 42020
rect 17876 41980 17885 42020
rect 18211 41980 18220 42020
rect 18260 41980 18412 42020
rect 18452 41980 18461 42020
rect 18691 41980 18700 42020
rect 18740 42011 19508 42020
rect 18740 41980 19468 42011
rect 17836 41962 17876 41971
rect 18220 41852 18260 41980
rect 19468 41962 19508 41971
rect 20131 41896 20140 41936
rect 20180 41896 21388 41936
rect 21428 41896 21437 41936
rect 4099 41812 4108 41852
rect 4148 41812 4780 41852
rect 4820 41812 4829 41852
rect 5827 41812 5836 41852
rect 5876 41812 6796 41852
rect 6836 41812 6845 41852
rect 7171 41812 7180 41852
rect 7220 41812 7852 41852
rect 7892 41812 7901 41852
rect 11491 41812 11500 41852
rect 11540 41812 12116 41852
rect 12259 41812 12268 41852
rect 12308 41812 13460 41852
rect 13795 41812 13804 41852
rect 13844 41812 14996 41852
rect 15772 41812 15820 41852
rect 15860 41812 15869 41852
rect 16291 41812 16300 41852
rect 16340 41812 16436 41852
rect 16675 41812 16684 41852
rect 16724 41812 18260 41852
rect 0 41768 90 41788
rect 14956 41768 14996 41812
rect 21510 41768 21600 41788
rect 0 41728 172 41768
rect 212 41728 221 41768
rect 1891 41728 1900 41768
rect 1940 41728 14188 41768
rect 14228 41728 14237 41768
rect 14851 41728 14860 41768
rect 14900 41728 14909 41768
rect 14956 41728 16003 41768
rect 16043 41728 16052 41768
rect 18403 41728 18412 41768
rect 18452 41728 21600 41768
rect 0 41708 90 41728
rect 14860 41684 14900 41728
rect 21510 41708 21600 41728
rect 7843 41644 7852 41684
rect 7892 41644 13804 41684
rect 13844 41644 13853 41684
rect 14860 41644 16108 41684
rect 16148 41644 16157 41684
rect 16483 41644 16492 41684
rect 16532 41644 18508 41684
rect 18548 41644 18557 41684
rect 3679 41560 3688 41600
rect 3728 41560 3770 41600
rect 3810 41560 3852 41600
rect 3892 41560 3934 41600
rect 3974 41560 4016 41600
rect 4056 41560 4065 41600
rect 4108 41560 7180 41600
rect 7220 41560 7229 41600
rect 8035 41560 8044 41600
rect 8084 41560 13996 41600
rect 14036 41560 14045 41600
rect 15619 41560 15628 41600
rect 15668 41560 17836 41600
rect 17876 41560 17885 41600
rect 18799 41560 18808 41600
rect 18848 41560 18890 41600
rect 18930 41560 18972 41600
rect 19012 41560 19054 41600
rect 19094 41560 19136 41600
rect 19176 41560 19185 41600
rect 19756 41560 21004 41600
rect 21044 41560 21053 41600
rect 4108 41516 4148 41560
rect 2860 41476 4148 41516
rect 4204 41476 12980 41516
rect 0 41432 90 41452
rect 2860 41432 2900 41476
rect 4204 41432 4244 41476
rect 12940 41432 12980 41476
rect 19756 41432 19796 41560
rect 0 41392 1612 41432
rect 1652 41392 1661 41432
rect 2537 41392 2668 41432
rect 2708 41392 2717 41432
rect 2764 41392 2900 41432
rect 4099 41392 4108 41432
rect 4148 41392 4244 41432
rect 4457 41392 4540 41432
rect 4580 41392 4588 41432
rect 4628 41392 4637 41432
rect 6499 41392 6508 41432
rect 6548 41392 8908 41432
rect 8948 41392 8957 41432
rect 9475 41392 9484 41432
rect 9524 41392 10540 41432
rect 10580 41392 10589 41432
rect 12451 41392 12460 41432
rect 12500 41392 12692 41432
rect 12940 41392 14188 41432
rect 14228 41392 14237 41432
rect 14818 41392 15619 41432
rect 15659 41392 15668 41432
rect 16195 41392 16204 41432
rect 16244 41392 16252 41432
rect 16292 41392 16375 41432
rect 16483 41392 16492 41432
rect 16532 41392 18028 41432
rect 18068 41392 18077 41432
rect 19180 41392 19796 41432
rect 19852 41476 21100 41516
rect 21140 41476 21149 41516
rect 0 41372 90 41392
rect 2764 41348 2804 41392
rect 1507 41308 1516 41348
rect 1556 41308 2804 41348
rect 2860 41308 12596 41348
rect 2476 41180 2516 41189
rect 2860 41180 2900 41308
rect 4483 41224 4492 41264
rect 4532 41224 4780 41264
rect 4820 41224 4829 41264
rect 5309 41224 5356 41264
rect 5396 41224 5405 41264
rect 5548 41224 6164 41264
rect 6499 41224 6508 41264
rect 6548 41224 6584 41264
rect 11177 41224 11308 41264
rect 11348 41224 11357 41264
rect 11884 41224 12460 41264
rect 12500 41224 12509 41264
rect 4108 41180 4148 41189
rect 5356 41180 5396 41224
rect 5548 41180 5588 41224
rect 6124 41180 6164 41224
rect 6508 41180 6548 41224
rect 6796 41180 6836 41189
rect 8716 41180 8756 41189
rect 10348 41180 10388 41189
rect 11884 41180 11924 41224
rect 12556 41180 12596 41308
rect 12652 41264 12692 41392
rect 14818 41348 14858 41392
rect 13315 41308 13324 41348
rect 13364 41308 14858 41348
rect 15139 41308 15148 41348
rect 15188 41308 15244 41348
rect 15284 41308 15319 41348
rect 16003 41308 16012 41348
rect 16052 41308 18700 41348
rect 18740 41308 18749 41348
rect 12652 41224 14572 41264
rect 14612 41224 14621 41264
rect 15283 41224 15292 41264
rect 15332 41224 15820 41264
rect 15860 41224 15869 41264
rect 18595 41224 18604 41264
rect 18644 41224 18988 41264
rect 19028 41224 19037 41264
rect 14956 41180 14996 41189
rect 15916 41180 15956 41189
rect 17644 41180 17684 41189
rect 19180 41180 19220 41392
rect 451 41140 460 41180
rect 500 41140 1228 41180
rect 1268 41140 1277 41180
rect 2345 41140 2476 41180
rect 2516 41140 2668 41180
rect 2708 41140 2717 41180
rect 2851 41140 2860 41180
rect 2900 41140 2909 41180
rect 3043 41140 3052 41180
rect 3092 41140 4108 41180
rect 4148 41140 4157 41180
rect 5033 41140 5164 41180
rect 5204 41140 5213 41180
rect 5347 41140 5356 41180
rect 5396 41140 5405 41180
rect 5539 41140 5548 41180
rect 5588 41140 5597 41180
rect 5644 41140 5687 41180
rect 5727 41140 5736 41180
rect 5897 41140 6019 41180
rect 6068 41140 6077 41180
rect 6124 41140 6316 41180
rect 6356 41140 6365 41180
rect 6488 41140 6497 41180
rect 6537 41140 6548 41180
rect 6665 41140 6796 41180
rect 6836 41140 6845 41180
rect 7049 41140 7084 41180
rect 7124 41140 7180 41180
rect 7220 41140 7229 41180
rect 7337 41140 7468 41180
rect 7508 41140 7517 41180
rect 8585 41140 8716 41180
rect 8756 41140 8765 41180
rect 9091 41140 9100 41180
rect 9140 41140 10156 41180
rect 10196 41140 10205 41180
rect 10627 41140 10636 41180
rect 10676 41140 10798 41180
rect 10838 41140 10847 41180
rect 10896 41140 10905 41180
rect 10945 41140 10964 41180
rect 2476 41131 2516 41140
rect 4108 41131 4148 41140
rect 0 41096 90 41116
rect 0 41056 76 41096
rect 116 41056 125 41096
rect 5068 41056 5260 41096
rect 5300 41056 5309 41096
rect 0 41036 90 41056
rect 4003 40972 4012 41012
rect 4052 40972 4300 41012
rect 4340 40972 4349 41012
rect 5068 40928 5108 41056
rect 5225 40972 5347 41012
rect 5396 40972 5405 41012
rect 5644 40928 5684 41140
rect 6124 41096 6164 41140
rect 6796 41131 6836 41140
rect 8716 41131 8756 41140
rect 10348 41096 10388 41140
rect 10924 41096 10964 41140
rect 11116 41140 11404 41180
rect 11444 41140 11500 41180
rect 11540 41140 11604 41180
rect 12250 41140 12364 41180
rect 12412 41140 12430 41180
rect 12556 41140 12980 41180
rect 13577 41140 13708 41180
rect 13748 41140 13757 41180
rect 14284 41140 14956 41180
rect 15305 41140 15436 41180
rect 15476 41140 15485 41180
rect 15785 41140 15916 41180
rect 15956 41140 15965 41180
rect 16099 41140 16108 41180
rect 16148 41140 16279 41180
rect 16387 41140 16396 41180
rect 16436 41140 16532 41180
rect 6115 41056 6124 41096
rect 6164 41056 6173 41096
rect 6569 41056 6604 41096
rect 6644 41056 6700 41096
rect 6740 41056 6749 41096
rect 10348 41056 10732 41096
rect 10772 41056 10781 41096
rect 10915 41056 10924 41096
rect 10964 41056 10992 41096
rect 11116 41012 11156 41140
rect 11884 41131 11924 41140
rect 12940 41096 12980 41140
rect 12940 41056 14188 41096
rect 14228 41056 14237 41096
rect 14284 41012 14324 41140
rect 14956 41096 14996 41140
rect 15916 41131 15956 41140
rect 14956 41056 15244 41096
rect 15284 41056 15293 41096
rect 15436 41056 15614 41096
rect 15654 41056 15663 41096
rect 15436 41012 15476 41056
rect 5866 40972 5875 41012
rect 5915 40972 5932 41012
rect 5972 40972 6055 41012
rect 6211 40972 6220 41012
rect 6260 40972 6391 41012
rect 6473 40972 6508 41012
rect 6548 40972 6595 41012
rect 6635 40972 6653 41012
rect 6700 40972 6940 41012
rect 6980 40972 6989 41012
rect 7171 40972 7180 41012
rect 7220 40972 11156 41012
rect 12547 40972 12556 41012
rect 12596 40972 12652 41012
rect 12692 40972 12727 41012
rect 13795 40972 13804 41012
rect 13844 40972 14324 41012
rect 15427 40972 15436 41012
rect 15476 40972 15485 41012
rect 15811 40972 15820 41012
rect 15860 40972 16204 41012
rect 16244 40972 16253 41012
rect 6700 40928 6740 40972
rect 16492 40928 16532 41140
rect 17731 41140 17740 41180
rect 17780 41140 18115 41180
rect 18155 41140 18164 41180
rect 18211 41140 18220 41180
rect 18260 41140 18391 41180
rect 18499 41140 18508 41180
rect 18548 41140 18700 41180
rect 18740 41140 18749 41180
rect 18883 41140 18892 41180
rect 18932 41140 19180 41180
rect 17644 41096 17684 41140
rect 19180 41131 19220 41140
rect 19276 41140 19668 41180
rect 19708 41140 19717 41180
rect 17597 41056 17644 41096
rect 17684 41056 17693 41096
rect 17740 41056 19124 41096
rect 1411 40888 1420 40928
rect 1460 40888 4108 40928
rect 4148 40888 4157 40928
rect 5068 40888 5684 40928
rect 6595 40888 6604 40928
rect 6644 40888 6740 40928
rect 7459 40888 7468 40928
rect 7508 40888 16244 40928
rect 16483 40888 16492 40928
rect 16532 40888 16541 40928
rect 0 40760 90 40780
rect 0 40720 1228 40760
rect 1268 40720 1277 40760
rect 0 40700 90 40720
rect 1769 40636 1852 40676
rect 1892 40636 1900 40676
rect 1940 40636 1949 40676
rect 2153 40636 2236 40676
rect 2276 40636 2284 40676
rect 2324 40636 2333 40676
rect 67 40552 76 40592
rect 116 40552 212 40592
rect 1459 40552 1468 40592
rect 1508 40552 1516 40592
rect 1556 40552 1639 40592
rect 2284 40552 2668 40592
rect 2708 40552 2717 40592
rect 172 40508 212 40552
rect 2284 40508 2324 40552
rect 172 40468 2036 40508
rect 2275 40468 2284 40508
rect 2324 40468 2333 40508
rect 2537 40468 2572 40508
rect 2612 40468 2659 40508
rect 2699 40468 2717 40508
rect 2760 40468 2769 40508
rect 2809 40468 2818 40508
rect 0 40424 90 40444
rect 1996 40424 2036 40468
rect 2764 40424 2804 40468
rect 0 40364 116 40424
rect 163 40384 172 40424
rect 212 40384 1228 40424
rect 1268 40384 1277 40424
rect 1481 40384 1612 40424
rect 1652 40384 1661 40424
rect 1987 40384 1996 40424
rect 2036 40384 2045 40424
rect 2659 40384 2668 40424
rect 2708 40384 2804 40424
rect 2860 40424 2900 40888
rect 4919 40804 4928 40844
rect 4968 40804 5010 40844
rect 5050 40804 5092 40844
rect 5132 40804 5174 40844
rect 5214 40804 5256 40844
rect 5296 40804 5305 40844
rect 5356 40676 5396 40888
rect 6019 40804 6028 40844
rect 6068 40804 12940 40844
rect 12980 40804 12989 40844
rect 13324 40804 16012 40844
rect 16052 40804 16061 40844
rect 13324 40760 13364 40804
rect 6787 40720 6796 40760
rect 6836 40720 7412 40760
rect 8707 40720 8716 40760
rect 8756 40720 9964 40760
rect 10004 40720 10013 40760
rect 10732 40720 13364 40760
rect 13411 40720 13420 40760
rect 13460 40720 15436 40760
rect 15476 40720 15485 40760
rect 4387 40636 4396 40676
rect 4436 40636 4492 40676
rect 4532 40636 4567 40676
rect 4963 40636 4972 40676
rect 5012 40636 5396 40676
rect 6211 40636 6220 40676
rect 6260 40636 6269 40676
rect 6787 40636 6796 40676
rect 6836 40636 7180 40676
rect 7220 40636 7229 40676
rect 6220 40592 6260 40636
rect 5068 40552 6124 40592
rect 6164 40552 6173 40592
rect 6220 40552 7014 40592
rect 7075 40552 7084 40592
rect 7124 40552 7217 40592
rect 5068 40508 5108 40552
rect 6974 40508 7014 40552
rect 7177 40508 7217 40552
rect 7372 40508 7412 40720
rect 9580 40676 9620 40720
rect 8236 40636 9484 40676
rect 9524 40636 9533 40676
rect 9580 40636 9628 40676
rect 9668 40636 9677 40676
rect 7738 40552 7747 40592
rect 7796 40552 7927 40592
rect 3017 40468 3148 40508
rect 3188 40468 3197 40508
rect 3331 40468 3340 40508
rect 3380 40499 3764 40508
rect 3380 40468 3724 40499
rect 4003 40468 4012 40508
rect 4052 40468 4216 40508
rect 4256 40468 4265 40508
rect 5050 40468 5059 40508
rect 5099 40468 5108 40508
rect 5155 40468 5164 40508
rect 5204 40468 5335 40508
rect 5539 40468 5548 40508
rect 5588 40468 5780 40508
rect 6019 40468 6028 40508
rect 6068 40468 6077 40508
rect 6124 40499 6164 40508
rect 3724 40450 3764 40459
rect 2860 40384 3244 40424
rect 3284 40384 3293 40424
rect 5251 40384 5260 40424
rect 5300 40384 5644 40424
rect 5684 40384 5693 40424
rect 76 40340 116 40364
rect 5740 40340 5780 40468
rect 76 40300 1420 40340
rect 1460 40300 1469 40340
rect 1699 40300 1708 40340
rect 1748 40300 2476 40340
rect 2516 40300 4876 40340
rect 4916 40300 4925 40340
rect 5635 40300 5644 40340
rect 5684 40300 5780 40340
rect 6028 40256 6068 40468
rect 6211 40468 6220 40508
rect 6260 40499 6644 40508
rect 6260 40468 6604 40499
rect 6124 40424 6164 40459
rect 6965 40468 6974 40508
rect 7014 40468 7023 40508
rect 7075 40468 7084 40508
rect 7124 40468 7133 40508
rect 7177 40468 7276 40508
rect 7316 40468 7325 40508
rect 7372 40468 7415 40508
rect 7455 40468 7464 40508
rect 7649 40468 7658 40508
rect 7698 40484 7707 40508
rect 6604 40424 6644 40459
rect 7084 40424 7124 40468
rect 7651 40444 7660 40468
rect 7700 40444 7805 40484
rect 8236 40424 8276 40636
rect 10732 40592 10772 40720
rect 11203 40636 11212 40676
rect 11252 40636 12364 40676
rect 12404 40636 12413 40676
rect 12844 40636 13507 40676
rect 13547 40636 13556 40676
rect 13603 40636 13612 40676
rect 13652 40636 14092 40676
rect 14132 40636 14141 40676
rect 15619 40636 15628 40676
rect 15668 40636 15744 40676
rect 8467 40552 8476 40592
rect 8516 40552 10772 40592
rect 12844 40592 12884 40636
rect 15628 40592 15668 40636
rect 12844 40552 12926 40592
rect 12966 40552 12975 40592
rect 13018 40552 13027 40592
rect 13067 40552 13076 40592
rect 13123 40552 13132 40592
rect 13172 40552 13181 40592
rect 13228 40552 13987 40592
rect 14027 40552 14036 40592
rect 14563 40552 14572 40592
rect 14612 40552 15676 40592
rect 15716 40552 15725 40592
rect 9641 40468 9772 40508
rect 9812 40468 9821 40508
rect 10243 40468 10252 40508
rect 10292 40468 10828 40508
rect 10868 40499 11060 40508
rect 10868 40468 11020 40499
rect 11020 40450 11060 40459
rect 13036 40424 13076 40552
rect 13132 40424 13172 40552
rect 13228 40499 13268 40552
rect 16204 40508 16244 40888
rect 17740 40676 17780 41056
rect 19084 41012 19124 41056
rect 19276 41012 19316 41140
rect 19852 41012 19892 41476
rect 20140 41392 20524 41432
rect 20564 41392 20573 41432
rect 20140 41264 20180 41392
rect 20371 41308 20380 41348
rect 20420 41308 20620 41348
rect 20660 41308 20669 41348
rect 21510 41264 21600 41284
rect 20131 41224 20140 41264
rect 20180 41224 20189 41264
rect 20236 41224 21600 41264
rect 20236 41180 20276 41224
rect 21510 41204 21600 41224
rect 20035 41140 20044 41180
rect 20084 41140 20276 41180
rect 17827 40972 17836 41012
rect 17876 40972 18007 41012
rect 19084 40972 19316 41012
rect 19843 40972 19852 41012
rect 19892 40972 19901 41012
rect 20039 40804 20048 40844
rect 20088 40804 20130 40844
rect 20170 40804 20212 40844
rect 20252 40804 20294 40844
rect 20334 40804 20376 40844
rect 20416 40804 20425 40844
rect 21510 40760 21600 40780
rect 20044 40720 21600 40760
rect 20044 40676 20084 40720
rect 21510 40700 21600 40720
rect 17635 40636 17644 40676
rect 17684 40636 17780 40676
rect 18281 40636 18364 40676
rect 18404 40636 18412 40676
rect 18452 40636 18461 40676
rect 20035 40636 20044 40676
rect 20084 40636 20093 40676
rect 20323 40636 20332 40676
rect 20372 40636 21100 40676
rect 21140 40636 21149 40676
rect 17356 40552 21292 40592
rect 21332 40552 21341 40592
rect 13315 40468 13324 40508
rect 13364 40468 13406 40508
rect 13446 40468 13495 40508
rect 13708 40499 13748 40508
rect 13228 40450 13268 40459
rect 13795 40468 13804 40508
rect 13844 40468 13886 40508
rect 13926 40468 13975 40508
rect 14188 40499 14228 40508
rect 6124 40384 6316 40424
rect 6356 40384 6365 40424
rect 6604 40384 7124 40424
rect 7363 40384 7372 40424
rect 7412 40384 7421 40424
rect 7546 40384 7555 40424
rect 7595 40384 7604 40424
rect 8035 40384 8044 40424
rect 8084 40384 8236 40424
rect 8276 40384 8285 40424
rect 8489 40384 8620 40424
rect 8660 40384 8669 40424
rect 8995 40384 9004 40424
rect 9044 40384 9196 40424
rect 9236 40384 9245 40424
rect 9353 40384 9388 40424
rect 9428 40384 9484 40424
rect 9524 40384 9533 40424
rect 12547 40384 12556 40424
rect 12596 40384 13076 40424
rect 13123 40384 13132 40424
rect 13172 40384 13181 40424
rect 7372 40340 7412 40384
rect 7564 40340 7604 40384
rect 7372 40300 7604 40340
rect 8851 40300 8860 40340
rect 8900 40300 10196 40340
rect 12713 40300 12796 40340
rect 12836 40300 12844 40340
rect 12884 40300 12893 40340
rect 10156 40256 10196 40300
rect 2947 40216 2956 40256
rect 2996 40216 6068 40256
rect 6307 40216 6316 40256
rect 6356 40216 6988 40256
rect 7028 40216 7037 40256
rect 8899 40216 8908 40256
rect 8948 40216 8956 40256
rect 8996 40216 9079 40256
rect 10156 40216 10580 40256
rect 1891 40132 1900 40172
rect 1940 40132 9964 40172
rect 10004 40132 10013 40172
rect 0 40088 90 40108
rect 10540 40088 10580 40216
rect 13708 40172 13748 40459
rect 14659 40468 14668 40508
rect 14708 40468 15092 40508
rect 14188 40424 14228 40459
rect 15052 40424 15092 40468
rect 15436 40468 15628 40508
rect 15668 40468 15677 40508
rect 16195 40468 16204 40508
rect 16244 40468 16253 40508
rect 16483 40468 16492 40508
rect 16532 40468 16876 40508
rect 16916 40468 16925 40508
rect 15436 40424 15476 40468
rect 17356 40424 17396 40552
rect 17452 40499 17548 40508
rect 17492 40468 17548 40499
rect 17588 40468 17623 40508
rect 17827 40468 17836 40508
rect 17876 40468 18595 40508
rect 18635 40468 18644 40508
rect 18691 40468 18700 40508
rect 18740 40468 18749 40508
rect 19075 40468 19084 40508
rect 19124 40468 19276 40508
rect 19316 40468 19325 40508
rect 19555 40468 19564 40508
rect 19604 40499 19735 40508
rect 19604 40468 19660 40499
rect 17452 40450 17492 40459
rect 18700 40424 18740 40468
rect 19700 40468 19735 40499
rect 20009 40468 20140 40508
rect 20180 40468 20189 40508
rect 19660 40450 19700 40459
rect 20140 40450 20180 40459
rect 14179 40384 14188 40424
rect 14228 40384 14275 40424
rect 14659 40384 14668 40424
rect 14708 40384 14717 40424
rect 15043 40384 15052 40424
rect 15092 40384 15101 40424
rect 15305 40384 15436 40424
rect 15476 40384 15485 40424
rect 15689 40384 15820 40424
rect 15860 40384 15869 40424
rect 16051 40384 16060 40424
rect 16100 40384 17396 40424
rect 17993 40384 18124 40424
rect 18164 40384 18173 40424
rect 18595 40384 18604 40424
rect 18644 40384 18740 40424
rect 18979 40384 18988 40424
rect 19028 40384 19180 40424
rect 19220 40384 19604 40424
rect 14668 40340 14708 40384
rect 19564 40340 19604 40384
rect 14083 40300 14092 40340
rect 14132 40300 14708 40340
rect 15283 40300 15292 40340
rect 15332 40300 19508 40340
rect 19564 40300 19852 40340
rect 19892 40300 19901 40340
rect 19468 40256 19508 40300
rect 21510 40256 21600 40276
rect 14899 40216 14908 40256
rect 14948 40216 19412 40256
rect 19468 40216 21600 40256
rect 13708 40132 14092 40172
rect 14132 40132 14141 40172
rect 19372 40088 19412 40216
rect 21510 40196 21600 40216
rect 0 40048 364 40088
rect 404 40048 413 40088
rect 3679 40048 3688 40088
rect 3728 40048 3770 40088
rect 3810 40048 3852 40088
rect 3892 40048 3934 40088
rect 3974 40048 4016 40088
rect 4056 40048 4065 40088
rect 8611 40048 8620 40088
rect 8660 40048 8812 40088
rect 8852 40048 8861 40088
rect 10252 40048 10419 40088
rect 10540 40048 16492 40088
rect 16532 40048 16541 40088
rect 18799 40048 18808 40088
rect 18848 40048 18890 40088
rect 18930 40048 18972 40088
rect 19012 40048 19054 40088
rect 19094 40048 19136 40088
rect 19176 40048 19185 40088
rect 19372 40048 20948 40088
rect 0 40028 90 40048
rect 10252 40004 10292 40048
rect 1468 39964 10292 40004
rect 10379 40004 10419 40048
rect 10379 39964 11980 40004
rect 12020 39964 12029 40004
rect 12547 39964 12556 40004
rect 12596 39964 14372 40004
rect 1468 39920 1508 39964
rect 1459 39880 1468 39920
rect 1508 39880 1517 39920
rect 1843 39880 1852 39920
rect 1892 39880 1900 39920
rect 1940 39880 2023 39920
rect 6028 39880 6124 39920
rect 6164 39880 6173 39920
rect 6281 39880 6403 39920
rect 6452 39880 6461 39920
rect 6874 39880 6883 39920
rect 6923 39880 6932 39920
rect 8419 39880 8428 39920
rect 8468 39880 12364 39920
rect 12404 39880 12413 39920
rect 13891 39880 13900 39920
rect 13940 39880 14228 39920
rect 6028 39836 6068 39880
rect 6892 39836 6932 39880
rect 1996 39796 2860 39836
rect 2900 39796 2909 39836
rect 4723 39796 4732 39836
rect 4772 39796 5164 39836
rect 5204 39796 5213 39836
rect 5260 39796 5836 39836
rect 5876 39796 5885 39836
rect 6019 39796 6028 39836
rect 6068 39796 6077 39836
rect 6139 39796 6932 39836
rect 9763 39796 9772 39836
rect 9812 39796 10060 39836
rect 10100 39796 10109 39836
rect 11011 39796 11020 39836
rect 11060 39796 11068 39836
rect 11108 39796 11191 39836
rect 12019 39796 12028 39836
rect 12068 39796 13844 39836
rect 0 39752 90 39772
rect 1996 39752 2036 39796
rect 0 39712 884 39752
rect 1097 39712 1228 39752
rect 1268 39712 1277 39752
rect 1411 39712 1420 39752
rect 1460 39712 1612 39752
rect 1652 39712 1661 39752
rect 1708 39712 1996 39752
rect 2036 39712 2045 39752
rect 2476 39712 2668 39752
rect 2708 39712 2804 39752
rect 3017 39712 3148 39752
rect 3188 39712 3197 39752
rect 4387 39712 4396 39752
rect 4436 39712 4780 39752
rect 4820 39712 5204 39752
rect 0 39692 90 39712
rect 844 39668 884 39712
rect 844 39628 1612 39668
rect 1652 39628 1661 39668
rect 1708 39584 1748 39712
rect 2476 39668 2516 39712
rect 2764 39668 2804 39712
rect 3724 39668 3764 39677
rect 5164 39668 5204 39712
rect 5260 39668 5300 39796
rect 6139 39752 6179 39796
rect 5347 39712 5356 39752
rect 5396 39712 5780 39752
rect 6118 39712 6127 39752
rect 6167 39712 6179 39752
rect 6508 39712 6604 39752
rect 6644 39712 6653 39752
rect 9100 39712 10348 39752
rect 10388 39712 10397 39752
rect 10819 39712 10828 39752
rect 10868 39712 10924 39752
rect 10964 39712 10999 39752
rect 12378 39712 12387 39752
rect 12427 39712 12940 39752
rect 12980 39712 12989 39752
rect 13507 39712 13516 39752
rect 13556 39712 13699 39752
rect 13739 39712 13748 39752
rect 5740 39668 5780 39712
rect 1795 39628 1804 39668
rect 1844 39628 2516 39668
rect 2650 39628 2659 39668
rect 2699 39628 2708 39668
rect 2755 39628 2764 39668
rect 2804 39628 2813 39668
rect 2947 39628 2956 39668
rect 2996 39628 3244 39668
rect 3284 39628 3293 39668
rect 3764 39628 3860 39668
rect 2668 39584 2708 39628
rect 3724 39619 3764 39628
rect 1699 39544 1708 39584
rect 1748 39544 1757 39584
rect 1891 39544 1900 39584
rect 1940 39544 2236 39584
rect 2276 39544 2285 39584
rect 2659 39544 2668 39584
rect 2708 39544 2755 39584
rect 931 39460 940 39500
rect 980 39460 3148 39500
rect 3188 39460 3197 39500
rect 0 39416 90 39436
rect 0 39376 1364 39416
rect 0 39356 90 39376
rect 0 39080 90 39100
rect 0 39040 1228 39080
rect 1268 39040 1277 39080
rect 0 39020 90 39040
rect 1324 38996 1364 39376
rect 1459 39124 1468 39164
rect 1508 39124 3724 39164
rect 3764 39124 3773 39164
rect 3820 39080 3860 39628
rect 3916 39628 4212 39668
rect 4252 39628 4261 39668
rect 4457 39628 4492 39668
rect 4532 39628 4588 39668
rect 4628 39628 4637 39668
rect 4723 39628 4732 39668
rect 4772 39628 4876 39668
rect 4916 39628 4925 39668
rect 5050 39628 5059 39668
rect 5099 39628 5108 39668
rect 5155 39628 5164 39668
rect 5204 39628 5213 39668
rect 5260 39628 5303 39668
rect 5343 39628 5352 39668
rect 5434 39628 5443 39668
rect 5483 39628 5492 39668
rect 5539 39628 5548 39668
rect 5588 39628 5597 39668
rect 5740 39628 5788 39668
rect 5828 39628 5837 39668
rect 5923 39628 5932 39668
rect 5993 39628 6103 39668
rect 6185 39628 6259 39668
rect 6299 39628 6316 39668
rect 6356 39628 6365 39668
rect 3916 39164 3956 39628
rect 4954 39544 4963 39584
rect 5003 39544 5012 39584
rect 4195 39460 4204 39500
rect 4244 39460 4396 39500
rect 4436 39460 4445 39500
rect 4828 39460 4876 39500
rect 4916 39460 4925 39500
rect 4828 39248 4868 39460
rect 4972 39416 5012 39544
rect 5068 39500 5108 39628
rect 5068 39460 5164 39500
rect 5204 39460 5213 39500
rect 4972 39376 5401 39416
rect 4919 39292 4928 39332
rect 4968 39292 5010 39332
rect 5050 39292 5092 39332
rect 5132 39292 5174 39332
rect 5214 39292 5256 39332
rect 5296 39292 5305 39332
rect 4828 39208 4916 39248
rect 4876 39164 4916 39208
rect 5361 39164 5401 39376
rect 5452 39248 5492 39628
rect 5548 39584 5588 39628
rect 6508 39584 6548 39712
rect 6700 39668 6740 39677
rect 7180 39668 7220 39677
rect 9100 39668 9140 39712
rect 12748 39668 12788 39712
rect 13804 39668 13844 39796
rect 14044 39796 14092 39836
rect 14132 39796 14141 39836
rect 6740 39628 7084 39668
rect 7124 39628 7133 39668
rect 7555 39628 7564 39668
rect 7604 39628 7852 39668
rect 7892 39628 8180 39668
rect 8227 39628 8236 39668
rect 8276 39628 8820 39668
rect 8860 39628 9140 39668
rect 9187 39628 9196 39668
rect 9236 39628 9484 39668
rect 9524 39628 9533 39668
rect 10443 39628 10452 39668
rect 10492 39628 10828 39668
rect 10868 39628 10877 39668
rect 11875 39628 11884 39668
rect 11924 39628 12212 39668
rect 6700 39619 6740 39628
rect 5548 39544 6028 39584
rect 6068 39544 6077 39584
rect 6211 39544 6220 39584
rect 6260 39544 6401 39584
rect 6452 39544 6461 39584
rect 6508 39544 6604 39584
rect 6644 39544 6653 39584
rect 6796 39544 6878 39584
rect 6918 39544 6927 39584
rect 6796 39500 6836 39544
rect 5626 39460 5635 39500
rect 5675 39460 5836 39500
rect 5876 39460 5885 39500
rect 6604 39460 6836 39500
rect 6953 39460 6988 39500
rect 7028 39460 7084 39500
rect 7124 39460 7133 39500
rect 6604 39248 6644 39460
rect 7180 39416 7220 39628
rect 8140 39500 8180 39628
rect 12172 39584 12212 39628
rect 12259 39610 12268 39668
rect 12308 39650 12317 39668
rect 12308 39610 12421 39650
rect 12496 39628 12505 39668
rect 12545 39628 12556 39668
rect 12596 39628 12685 39668
rect 12739 39628 12748 39668
rect 12788 39628 12797 39668
rect 12940 39628 13027 39668
rect 13067 39628 13076 39668
rect 13411 39628 13420 39668
rect 13460 39628 13559 39668
rect 13599 39628 13608 39668
rect 13795 39628 13804 39668
rect 13844 39628 13853 39668
rect 12940 39584 12980 39628
rect 14044 39584 14084 39796
rect 14188 39752 14228 39880
rect 14332 39836 14372 39964
rect 17609 39880 17740 39920
rect 17780 39880 17789 39920
rect 18739 39880 18748 39920
rect 18788 39880 19948 39920
rect 19988 39880 19997 39920
rect 20131 39880 20140 39920
rect 20180 39880 20332 39920
rect 20372 39880 20381 39920
rect 14332 39796 14420 39836
rect 14467 39796 14476 39836
rect 14516 39796 15284 39836
rect 18355 39796 18364 39836
rect 18404 39796 20044 39836
rect 20084 39796 20093 39836
rect 14188 39712 14324 39752
rect 14284 39668 14324 39712
rect 14380 39668 14420 39796
rect 14659 39712 14668 39752
rect 14708 39712 14900 39752
rect 14170 39628 14179 39668
rect 14219 39628 14228 39668
rect 14275 39628 14284 39668
rect 14324 39628 14333 39668
rect 14380 39628 14764 39668
rect 14804 39628 14813 39668
rect 8908 39544 10100 39584
rect 12163 39544 12172 39584
rect 12212 39544 12221 39584
rect 12643 39544 12652 39584
rect 12692 39544 12980 39584
rect 13027 39544 13036 39584
rect 13076 39544 13132 39584
rect 13172 39544 13207 39584
rect 13459 39544 13468 39584
rect 13508 39544 14084 39584
rect 14188 39584 14228 39628
rect 14188 39544 14668 39584
rect 14708 39544 14717 39584
rect 8908 39500 8948 39544
rect 10060 39500 10100 39544
rect 8140 39460 8948 39500
rect 8995 39460 9004 39500
rect 9044 39460 9292 39500
rect 9332 39460 9341 39500
rect 10060 39460 10292 39500
rect 10505 39460 10636 39500
rect 10676 39460 10685 39500
rect 13123 39460 13132 39500
rect 13172 39460 13891 39500
rect 13931 39460 13940 39500
rect 10252 39416 10292 39460
rect 14860 39416 14900 39712
rect 15244 39668 15284 39796
rect 20908 39752 20948 40048
rect 21510 39752 21600 39772
rect 15811 39712 15820 39752
rect 15860 39712 16340 39752
rect 17993 39712 18124 39752
rect 18164 39712 18173 39752
rect 18377 39712 18508 39752
rect 18548 39712 18557 39752
rect 20908 39712 21600 39752
rect 16300 39668 16340 39712
rect 21510 39692 21600 39712
rect 17548 39668 17588 39677
rect 20140 39668 20180 39677
rect 15754 39628 15763 39668
rect 15803 39628 15860 39668
rect 16291 39628 16300 39668
rect 16340 39628 16349 39668
rect 17417 39628 17548 39668
rect 17588 39628 17597 39668
rect 18761 39628 18892 39668
rect 18932 39628 18941 39668
rect 15244 39619 15284 39628
rect 6691 39376 6700 39416
rect 6740 39376 7220 39416
rect 9475 39376 9484 39416
rect 9524 39376 10060 39416
rect 10100 39376 10109 39416
rect 10252 39376 11500 39416
rect 11540 39376 11549 39416
rect 13612 39376 14900 39416
rect 13612 39332 13652 39376
rect 8515 39292 8524 39332
rect 8564 39292 10924 39332
rect 10964 39292 10973 39332
rect 13219 39292 13228 39332
rect 13268 39292 13652 39332
rect 5452 39208 6644 39248
rect 6979 39208 6988 39248
rect 7028 39208 8620 39248
rect 8660 39208 8669 39248
rect 8803 39208 8812 39248
rect 8852 39208 13036 39248
rect 13076 39208 13085 39248
rect 13411 39208 13420 39248
rect 13460 39208 13469 39248
rect 6604 39164 6644 39208
rect 13420 39164 13460 39208
rect 3907 39124 3916 39164
rect 3956 39124 3965 39164
rect 4867 39124 4876 39164
rect 4916 39124 4925 39164
rect 5361 39124 5548 39164
rect 5588 39124 5597 39164
rect 5897 39124 5932 39164
rect 5972 39124 6028 39164
rect 6068 39124 6077 39164
rect 6595 39124 6604 39164
rect 6644 39124 6653 39164
rect 8777 39124 8812 39164
rect 8852 39124 8908 39164
rect 8948 39124 8957 39164
rect 9004 39124 9292 39164
rect 9332 39124 9341 39164
rect 12521 39124 12556 39164
rect 12596 39124 12652 39164
rect 12692 39124 12701 39164
rect 12940 39124 13460 39164
rect 5932 39080 5972 39124
rect 9004 39080 9044 39124
rect 3820 39040 5972 39080
rect 6211 39040 6220 39080
rect 6260 39040 6269 39080
rect 6604 39040 6796 39080
rect 6836 39040 6845 39080
rect 7564 39040 8332 39080
rect 8372 39040 8381 39080
rect 8620 39040 9044 39080
rect 9100 39040 11116 39080
rect 11156 39040 12788 39080
rect 6220 38996 6260 39040
rect 6604 38996 6644 39040
rect 7170 39029 7220 39038
rect 1324 38956 2036 38996
rect 2345 38956 2476 38996
rect 2516 38956 2525 38996
rect 3724 38987 4012 38996
rect 1996 38912 2036 38956
rect 3764 38956 4012 38987
rect 4052 38956 4061 38996
rect 4186 38956 4195 38996
rect 4235 38956 4244 38996
rect 4291 38956 4300 38996
rect 4340 38956 4471 38996
rect 4553 38956 4684 38996
rect 4724 38956 4733 38996
rect 5260 38987 5452 38996
rect 3724 38938 3764 38947
rect 4204 38912 4244 38956
rect 5300 38956 5452 38987
rect 5492 38956 5501 38996
rect 5609 38956 5740 38996
rect 5780 38956 5789 38996
rect 5993 38956 6124 38996
rect 6164 38956 6173 38996
rect 6220 38956 6239 38996
rect 6279 38956 6307 38996
rect 6403 38956 6412 38996
rect 6452 38956 6461 38996
rect 6595 38956 6604 38996
rect 6644 38956 6653 38996
rect 6787 38956 6796 38996
rect 6836 38956 6845 38996
rect 6923 38956 6988 38996
rect 7028 38956 7054 38996
rect 7094 38956 7103 38996
rect 7170 38989 7171 39029
rect 7211 38996 7220 39029
rect 7564 38996 7604 39040
rect 7211 38989 7276 38996
rect 7170 38980 7276 38989
rect 7180 38956 7276 38980
rect 7316 38956 7325 38996
rect 7555 38956 7564 38996
rect 7604 38956 7613 38996
rect 8140 38987 8180 38996
rect 5260 38938 5300 38947
rect 5740 38938 5780 38947
rect 6412 38912 6452 38956
rect 6796 38912 6836 38956
rect 355 38872 364 38912
rect 404 38872 1228 38912
rect 1268 38872 1277 38912
rect 1481 38872 1612 38912
rect 1652 38872 1661 38912
rect 1987 38872 1996 38912
rect 2036 38872 2045 38912
rect 2227 38872 2236 38912
rect 2276 38872 3668 38912
rect 4195 38872 4204 38912
rect 4244 38872 4291 38912
rect 4649 38872 4780 38912
rect 4820 38872 4829 38912
rect 6412 38872 6700 38912
rect 6740 38872 6749 38912
rect 6796 38872 6892 38912
rect 6932 38872 6941 38912
rect 7171 38872 7180 38912
rect 7220 38872 7660 38912
rect 7700 38872 7709 38912
rect 3628 38828 3668 38872
rect 8140 38828 8180 38947
rect 8620 38987 8660 39040
rect 8803 38956 8812 38996
rect 8852 38956 9004 38996
rect 9044 38956 9053 38996
rect 8620 38938 8660 38947
rect 9100 38912 9140 39040
rect 12748 38996 12788 39040
rect 12940 38996 12980 39124
rect 13612 39080 13652 39292
rect 15820 39164 15860 39628
rect 17548 39619 17588 39628
rect 20140 39584 20180 39628
rect 17635 39544 17644 39584
rect 17684 39544 20180 39584
rect 15907 39460 15916 39500
rect 15956 39460 21292 39500
rect 21332 39460 21341 39500
rect 20039 39292 20048 39332
rect 20088 39292 20130 39332
rect 20170 39292 20212 39332
rect 20252 39292 20294 39332
rect 20334 39292 20376 39332
rect 20416 39292 20425 39332
rect 21510 39248 21600 39268
rect 20611 39208 20620 39248
rect 20660 39208 21600 39248
rect 21510 39188 21600 39208
rect 13939 39124 13948 39164
rect 13988 39124 14188 39164
rect 14228 39124 14237 39164
rect 15820 39124 15916 39164
rect 15956 39124 15965 39164
rect 16723 39124 16732 39164
rect 16772 39124 18508 39164
rect 18548 39124 18557 39164
rect 13603 39040 13612 39080
rect 13652 39040 13661 39080
rect 14323 39040 14332 39080
rect 14372 39040 21004 39080
rect 21044 39040 21053 39080
rect 10252 38987 10772 38996
rect 10292 38956 10772 38987
rect 10915 38956 10924 38996
rect 10964 38956 11116 38996
rect 11156 38956 11203 38996
rect 11875 38956 11884 38996
rect 11924 38987 12404 38996
rect 11924 38956 12364 38987
rect 10252 38938 10292 38947
rect 10732 38912 10772 38956
rect 11116 38912 11156 38956
rect 12739 38956 12748 38996
rect 12788 38956 12797 38996
rect 12931 38956 12940 38996
rect 12980 38956 12989 38996
rect 13097 38956 13228 38996
rect 13268 38956 13277 38996
rect 13385 38956 13507 38996
rect 13556 38956 13565 38996
rect 13612 38956 13708 38996
rect 13748 38956 14476 38996
rect 14516 38956 14525 38996
rect 15689 38987 15820 38996
rect 15689 38956 15724 38987
rect 12364 38938 12404 38947
rect 12940 38912 12980 38956
rect 13612 38912 13652 38956
rect 15764 38956 15820 38987
rect 15860 38956 15869 38996
rect 16867 38956 16876 38996
rect 16916 38956 16972 38996
rect 17012 38956 17047 38996
rect 18019 38956 18028 38996
rect 18068 38987 18260 38996
rect 18068 38956 18220 38987
rect 15724 38938 15764 38947
rect 18220 38938 18260 38947
rect 18316 38956 18700 38996
rect 18740 38956 18749 38996
rect 19948 38987 19988 38996
rect 8716 38872 9140 38912
rect 9196 38872 10196 38912
rect 8716 38828 8756 38872
rect 3628 38788 6356 38828
rect 8140 38788 8428 38828
rect 8468 38788 8756 38828
rect 0 38744 90 38764
rect 6316 38744 6356 38788
rect 9196 38744 9236 38872
rect 10156 38828 10196 38872
rect 10348 38872 10636 38912
rect 10676 38872 10685 38912
rect 10732 38872 10828 38912
rect 10868 38872 10877 38912
rect 11107 38872 11116 38912
rect 11156 38872 11165 38912
rect 12451 38872 12460 38912
rect 12500 38872 12980 38912
rect 13027 38872 13036 38912
rect 13076 38872 13652 38912
rect 13961 38872 13996 38912
rect 14036 38872 14092 38912
rect 14132 38872 14141 38912
rect 16291 38872 16300 38912
rect 16340 38872 16492 38912
rect 16532 38872 16541 38912
rect 10348 38828 10388 38872
rect 10156 38788 10388 38828
rect 10732 38828 10772 38872
rect 18316 38828 18356 38956
rect 19948 38912 19988 38947
rect 18499 38872 18508 38912
rect 18548 38872 19988 38912
rect 10732 38788 11020 38828
rect 11060 38788 11069 38828
rect 15427 38788 15436 38828
rect 15476 38788 18124 38828
rect 18164 38788 18356 38828
rect 21510 38744 21600 38764
rect 0 38704 1612 38744
rect 1652 38704 1661 38744
rect 1843 38704 1852 38744
rect 1892 38704 1900 38744
rect 1940 38704 2023 38744
rect 5164 38704 6124 38744
rect 6164 38704 6173 38744
rect 6316 38704 9236 38744
rect 10313 38704 10444 38744
rect 10484 38704 10493 38744
rect 12739 38704 12748 38744
rect 12788 38704 12797 38744
rect 16003 38704 16012 38744
rect 16052 38704 16060 38744
rect 16100 38704 16183 38744
rect 18281 38704 18412 38744
rect 18452 38704 18461 38744
rect 19939 38704 19948 38744
rect 19988 38704 20140 38744
rect 20180 38704 20189 38744
rect 20236 38704 21600 38744
rect 0 38684 90 38704
rect 3679 38536 3688 38576
rect 3728 38536 3770 38576
rect 3810 38536 3852 38576
rect 3892 38536 3934 38576
rect 3974 38536 4016 38576
rect 4056 38536 4065 38576
rect 3523 38452 3532 38492
rect 3572 38452 3581 38492
rect 0 38408 90 38428
rect 0 38368 1460 38408
rect 2563 38368 2572 38408
rect 2612 38368 2668 38408
rect 2708 38368 2743 38408
rect 0 38348 90 38368
rect 1420 38324 1460 38368
rect 1420 38284 2764 38324
rect 2804 38284 2813 38324
rect 2476 38200 3052 38240
rect 3092 38200 3101 38240
rect 2476 38156 2516 38200
rect 3532 38156 3572 38452
rect 4291 38368 4300 38408
rect 4340 38368 4471 38408
rect 5164 38240 5204 38704
rect 12748 38660 12788 38704
rect 20236 38660 20276 38704
rect 21510 38684 21600 38704
rect 12643 38620 12652 38660
rect 12692 38620 12788 38660
rect 19843 38620 19852 38660
rect 19892 38620 20276 38660
rect 5443 38536 5452 38576
rect 5492 38536 16780 38576
rect 16820 38536 16829 38576
rect 18799 38536 18808 38576
rect 18848 38536 18890 38576
rect 18930 38536 18972 38576
rect 19012 38536 19054 38576
rect 19094 38536 19136 38576
rect 19176 38536 19185 38576
rect 6691 38452 6700 38492
rect 6740 38452 11596 38492
rect 11636 38452 11645 38492
rect 12076 38452 12268 38492
rect 12308 38452 12748 38492
rect 12788 38452 12797 38492
rect 12076 38408 12116 38452
rect 12067 38368 12076 38408
rect 12116 38368 12125 38408
rect 12403 38368 12412 38408
rect 12452 38368 12460 38408
rect 12500 38368 12583 38408
rect 14537 38368 14668 38408
rect 14708 38368 14717 38408
rect 15593 38368 15676 38408
rect 15716 38368 15724 38408
rect 15764 38368 15773 38408
rect 18028 38368 18508 38408
rect 18548 38368 18557 38408
rect 5827 38284 5836 38324
rect 5876 38284 5885 38324
rect 5993 38284 6124 38324
rect 6164 38284 6173 38324
rect 6499 38284 6508 38324
rect 6548 38284 6988 38324
rect 7028 38284 7037 38324
rect 8611 38284 8620 38324
rect 8660 38284 9964 38324
rect 10004 38284 10013 38324
rect 10636 38284 12172 38324
rect 12212 38284 12221 38324
rect 12503 38284 13228 38324
rect 13268 38284 13277 38324
rect 4291 38200 4300 38240
rect 4340 38200 4492 38240
rect 4532 38200 4541 38240
rect 5164 38200 5283 38240
rect 5323 38200 5332 38240
rect 5539 38200 5548 38240
rect 5588 38200 5597 38240
rect 4108 38156 4148 38165
rect 5548 38156 5588 38200
rect 5836 38156 5876 38284
rect 5923 38200 5932 38240
rect 5972 38200 6356 38240
rect 6586 38200 6595 38240
rect 6635 38200 7756 38240
rect 7796 38200 7805 38240
rect 8297 38200 8428 38240
rect 8468 38200 8477 38240
rect 8803 38200 8812 38240
rect 8852 38200 9196 38240
rect 9236 38200 9245 38240
rect 9475 38200 9484 38240
rect 9524 38200 9676 38240
rect 9716 38200 9725 38240
rect 6316 38156 6356 38200
rect 10636 38156 10676 38284
rect 11884 38156 11924 38165
rect 12503 38156 12543 38284
rect 12634 38200 12643 38240
rect 12683 38200 12844 38240
rect 12884 38200 12893 38240
rect 14921 38200 15052 38240
rect 15092 38200 15101 38240
rect 15305 38200 15436 38240
rect 15476 38200 15485 38240
rect 15811 38200 15820 38240
rect 15860 38200 16012 38240
rect 16052 38200 16061 38240
rect 16483 38200 16492 38240
rect 16532 38200 16876 38240
rect 16916 38200 16925 38240
rect 14476 38156 14516 38165
rect 15820 38156 15860 38200
rect 16780 38156 16820 38200
rect 18028 38156 18068 38368
rect 18364 38284 18412 38324
rect 18452 38284 18461 38324
rect 18364 38198 18404 38284
rect 21510 38240 21600 38260
rect 18979 38200 18988 38240
rect 19028 38200 19276 38240
rect 19316 38200 19325 38240
rect 19651 38200 19660 38240
rect 19700 38200 21600 38240
rect 18364 38174 18548 38198
rect 21510 38180 21600 38200
rect 18364 38158 18499 38174
rect 1193 38116 1228 38156
rect 1268 38116 1324 38156
rect 1364 38116 1373 38156
rect 2851 38116 2860 38156
rect 2900 38116 3572 38156
rect 3977 38116 4108 38156
rect 4148 38116 4157 38156
rect 5155 38116 5164 38156
rect 5204 38116 5213 38156
rect 5392 38116 5401 38156
rect 5441 38116 5492 38156
rect 5539 38116 5548 38156
rect 5588 38116 5635 38156
rect 5722 38116 5731 38156
rect 5771 38116 5780 38156
rect 5827 38116 5836 38156
rect 5876 38116 5885 38156
rect 6019 38116 6028 38156
rect 6068 38116 6077 38156
rect 6144 38116 6153 38156
rect 6193 38116 6260 38156
rect 6307 38116 6316 38156
rect 6356 38116 6365 38156
rect 6466 38116 6475 38156
rect 6515 38116 6548 38156
rect 2476 38107 2516 38116
rect 0 38072 90 38092
rect 4108 38072 4148 38116
rect 0 38032 748 38072
rect 788 38032 797 38072
rect 2860 38032 4148 38072
rect 0 38012 90 38032
rect 2860 37904 2900 38032
rect 5164 37988 5204 38116
rect 5452 38072 5492 38116
rect 5740 38072 5780 38116
rect 6028 38072 6068 38116
rect 6220 38072 6260 38116
rect 5452 38032 5635 38072
rect 5675 38032 5684 38072
rect 5740 38032 5836 38072
rect 5876 38032 5885 38072
rect 6028 38032 6124 38072
rect 6164 38032 6173 38072
rect 6220 38032 6316 38072
rect 6356 38032 6365 38072
rect 6508 37988 6548 38116
rect 4723 37948 4732 37988
rect 4772 37948 4820 37988
rect 5059 37948 5068 37988
rect 5108 37948 5117 37988
rect 5164 37948 5452 37988
rect 5492 37948 6548 37988
rect 6604 38116 6700 38156
rect 6740 38116 6749 38156
rect 6979 38116 6988 38156
rect 7028 38116 7037 38156
rect 7084 38116 7103 38156
rect 7143 38116 7171 38156
rect 7241 38116 7276 38156
rect 7316 38116 7372 38156
rect 7412 38116 7421 38156
rect 10627 38116 10636 38156
rect 10676 38116 10685 38156
rect 11753 38116 11884 38156
rect 11924 38116 11933 38156
rect 12163 38116 12172 38156
rect 12212 38116 12268 38156
rect 12308 38116 12503 38156
rect 12543 38116 12552 38156
rect 12617 38116 12748 38156
rect 12788 38116 13172 38156
rect 13219 38116 13228 38156
rect 13268 38116 13804 38156
rect 13844 38116 13853 38156
rect 2851 37864 2860 37904
rect 2900 37864 2909 37904
rect 0 37736 90 37756
rect 4780 37736 4820 37948
rect 5068 37904 5108 37948
rect 5068 37864 5401 37904
rect 5361 37820 5401 37864
rect 6604 37820 6644 38116
rect 6988 38072 7028 38116
rect 7084 38072 7124 38116
rect 11884 38107 11924 38116
rect 13132 38072 13172 38116
rect 6883 38032 6892 38072
rect 6932 38032 7028 38072
rect 7075 38032 7084 38072
rect 7124 38032 7133 38072
rect 10819 38032 10828 38072
rect 10868 38032 11596 38072
rect 11636 38032 11645 38072
rect 12556 38032 12980 38072
rect 13132 38032 13516 38072
rect 13556 38032 13565 38072
rect 12556 37988 12596 38032
rect 12940 37988 12980 38032
rect 13612 37988 13652 38116
rect 14476 38072 14516 38116
rect 15436 38116 15860 38156
rect 16771 38116 16780 38156
rect 16820 38116 16896 38156
rect 18490 38134 18499 38158
rect 18539 38134 18548 38174
rect 19564 38156 19604 38165
rect 18490 38133 18548 38134
rect 18592 38116 18601 38156
rect 18641 38116 18740 38156
rect 18953 38116 19084 38156
rect 19124 38116 19133 38156
rect 20074 38116 20083 38156
rect 20123 38116 20524 38156
rect 20564 38116 20573 38156
rect 15436 38072 15476 38116
rect 18028 38107 18068 38116
rect 18700 38072 18740 38116
rect 14476 38032 15436 38072
rect 15476 38032 15485 38072
rect 15811 38032 15820 38072
rect 15860 38032 16060 38072
rect 16100 38032 16492 38072
rect 16532 38032 16541 38072
rect 18403 38032 18412 38072
rect 18452 38032 18604 38072
rect 18644 38032 18740 38072
rect 6778 37948 6787 37988
rect 6836 37948 6967 37988
rect 7363 37948 7372 37988
rect 7412 37948 8188 37988
rect 8228 37948 8237 37988
rect 8489 37948 8572 37988
rect 8612 37948 8620 37988
rect 8660 37948 8669 37988
rect 9427 37948 9436 37988
rect 9476 37948 10484 37988
rect 10531 37948 10540 37988
rect 10580 37948 12596 37988
rect 12713 37948 12748 37988
rect 12788 37948 12835 37988
rect 12875 37948 12893 37988
rect 12940 37948 13652 37988
rect 14729 37948 14812 37988
rect 14852 37948 14860 37988
rect 14900 37948 15244 37988
rect 15284 37948 15293 37988
rect 15340 37948 16252 37988
rect 16292 37948 16301 37988
rect 18211 37948 18220 37988
rect 18260 37948 18269 37988
rect 10444 37904 10484 37948
rect 15340 37904 15380 37948
rect 10444 37864 11500 37904
rect 11540 37864 11549 37904
rect 12259 37864 12268 37904
rect 12308 37864 15380 37904
rect 4919 37780 4928 37820
rect 4968 37780 5010 37820
rect 5050 37780 5092 37820
rect 5132 37780 5174 37820
rect 5214 37780 5256 37820
rect 5296 37780 5305 37820
rect 5361 37780 6644 37820
rect 9475 37780 9484 37820
rect 9524 37780 10540 37820
rect 10580 37780 10589 37820
rect 11587 37780 11596 37820
rect 11636 37780 12844 37820
rect 12884 37780 12893 37820
rect 0 37696 844 37736
rect 884 37696 893 37736
rect 4780 37696 12556 37736
rect 12596 37696 12605 37736
rect 0 37676 90 37696
rect 2083 37612 2092 37652
rect 2132 37612 5204 37652
rect 5321 37612 5452 37652
rect 5492 37612 5501 37652
rect 5827 37612 5836 37652
rect 5876 37612 8035 37652
rect 8075 37612 8084 37652
rect 12041 37612 12172 37652
rect 12212 37612 12221 37652
rect 12940 37612 13132 37652
rect 13172 37612 13181 37652
rect 13289 37612 13372 37652
rect 13412 37612 13420 37652
rect 13460 37612 13469 37652
rect 5164 37568 5204 37612
rect 3427 37528 3436 37568
rect 3476 37528 4052 37568
rect 5164 37528 5684 37568
rect 7075 37528 7084 37568
rect 7124 37528 7988 37568
rect 8035 37528 8044 37568
rect 8084 37528 8247 37568
rect 8287 37528 8296 37568
rect 9292 37528 10060 37568
rect 10100 37528 10109 37568
rect 11820 37528 11884 37568
rect 11924 37528 12844 37568
rect 12884 37528 12893 37568
rect 4012 37484 4052 37528
rect 5644 37484 5684 37528
rect 1219 37444 1228 37484
rect 1268 37444 1708 37484
rect 1748 37444 1757 37484
rect 2476 37475 2860 37484
rect 2516 37444 2860 37475
rect 2900 37444 2909 37484
rect 3100 37444 3820 37484
rect 3860 37444 3869 37484
rect 4003 37444 4012 37484
rect 4052 37444 4061 37484
rect 4771 37444 4780 37484
rect 4820 37475 5300 37484
rect 4820 37444 5260 37475
rect 2476 37426 2516 37435
rect 0 37400 90 37420
rect 3100 37400 3140 37444
rect 5635 37444 5644 37484
rect 5684 37444 5932 37484
rect 5972 37444 5981 37484
rect 6115 37444 6124 37484
rect 6164 37444 6700 37484
rect 6740 37475 6932 37484
rect 6740 37444 6892 37475
rect 5260 37426 5300 37435
rect 6892 37426 6932 37435
rect 7372 37475 7412 37528
rect 7948 37484 7988 37528
rect 7594 37475 7660 37484
rect 7372 37426 7412 37435
rect 7462 37424 7471 37464
rect 7511 37424 7520 37464
rect 7594 37435 7603 37475
rect 7643 37444 7660 37475
rect 7700 37444 7783 37484
rect 7930 37444 7939 37484
rect 7979 37444 7988 37484
rect 9292 37475 9332 37528
rect 7643 37435 7652 37444
rect 7594 37434 7652 37435
rect 9955 37444 9964 37484
rect 10004 37444 10292 37484
rect 10409 37444 10540 37484
rect 10580 37444 10589 37484
rect 10636 37444 10732 37484
rect 10772 37444 11500 37484
rect 11540 37444 11549 37484
rect 11980 37475 12020 37528
rect 12940 37484 12980 37612
rect 13180 37528 13324 37568
rect 13364 37528 13373 37568
rect 17827 37528 17836 37568
rect 17876 37528 17884 37568
rect 17924 37528 18007 37568
rect 13180 37484 13220 37528
rect 18220 37484 18260 37948
rect 19564 37568 19604 38116
rect 20227 37948 20236 37988
rect 20276 37948 20908 37988
rect 20948 37948 20957 37988
rect 20039 37780 20048 37820
rect 20088 37780 20130 37820
rect 20170 37780 20212 37820
rect 20252 37780 20294 37820
rect 20334 37780 20376 37820
rect 20416 37780 20425 37820
rect 21510 37736 21600 37756
rect 20995 37696 21004 37736
rect 21044 37696 21600 37736
rect 21510 37676 21600 37696
rect 18403 37528 18412 37568
rect 18452 37528 18644 37568
rect 18883 37528 18892 37568
rect 18932 37528 19604 37568
rect 18604 37484 18644 37528
rect 9292 37426 9332 37435
rect 0 37360 212 37400
rect 2729 37360 2764 37400
rect 2804 37360 2860 37400
rect 2900 37360 2964 37400
rect 3091 37360 3100 37400
rect 3140 37360 3149 37400
rect 3235 37360 3244 37400
rect 3284 37360 3293 37400
rect 3619 37360 3628 37400
rect 3668 37360 3677 37400
rect 0 37340 90 37360
rect 172 37232 212 37360
rect 3244 37316 3284 37360
rect 2537 37276 2668 37316
rect 2708 37276 2717 37316
rect 2860 37276 3284 37316
rect 2860 37232 2900 37276
rect 172 37192 2900 37232
rect 3331 37192 3340 37232
rect 3380 37192 3484 37232
rect 3524 37192 3533 37232
rect 3628 37148 3668 37360
rect 7471 37316 7511 37424
rect 10252 37400 10292 37444
rect 10636 37400 10676 37444
rect 12521 37444 12619 37484
rect 12692 37444 12701 37484
rect 12835 37444 12844 37484
rect 12884 37444 12980 37484
rect 13036 37444 13220 37484
rect 13385 37444 13516 37484
rect 13556 37444 13565 37484
rect 13673 37444 13804 37484
rect 13844 37444 13853 37484
rect 14921 37444 15052 37484
rect 15092 37444 15101 37484
rect 15235 37444 15244 37484
rect 15284 37475 15668 37484
rect 15284 37444 15628 37475
rect 11980 37426 12020 37435
rect 13036 37400 13076 37444
rect 15052 37426 15092 37435
rect 16579 37444 16588 37484
rect 16628 37444 16876 37484
rect 16916 37444 16925 37484
rect 18220 37444 18499 37484
rect 18539 37444 18548 37484
rect 18595 37444 18604 37484
rect 18644 37444 18653 37484
rect 18979 37444 18988 37484
rect 19028 37444 19276 37484
rect 19316 37444 19325 37484
rect 19564 37475 19604 37528
rect 15628 37426 15668 37435
rect 19939 37444 19948 37484
rect 19988 37475 20119 37484
rect 19988 37444 20044 37475
rect 19564 37426 19604 37435
rect 20084 37444 20119 37475
rect 20044 37426 20084 37435
rect 7747 37360 7756 37400
rect 7796 37360 8620 37400
rect 8660 37360 8716 37400
rect 8756 37360 8765 37400
rect 10252 37360 10676 37400
rect 12617 37360 12739 37400
rect 12788 37360 12797 37400
rect 12876 37360 12940 37400
rect 12980 37360 13076 37400
rect 13123 37360 13132 37400
rect 13172 37360 13181 37400
rect 13603 37360 13612 37400
rect 13652 37360 13660 37400
rect 13700 37360 13783 37400
rect 16867 37360 16876 37400
rect 16916 37360 17068 37400
rect 17108 37360 17117 37400
rect 17225 37360 17308 37400
rect 17348 37360 17356 37400
rect 17396 37360 17405 37400
rect 17513 37360 17644 37400
rect 17684 37360 17693 37400
rect 17993 37360 18124 37400
rect 18164 37360 18604 37400
rect 18644 37360 18653 37400
rect 18953 37360 19084 37400
rect 19124 37360 19133 37400
rect 7267 37276 7276 37316
rect 7316 37276 7511 37316
rect 7660 37276 8812 37316
rect 8852 37276 8861 37316
rect 8947 37276 8956 37316
rect 8996 37276 10348 37316
rect 10388 37276 10397 37316
rect 3859 37192 3868 37232
rect 3908 37192 4108 37232
rect 4148 37192 4157 37232
rect 6307 37192 6316 37232
rect 6356 37192 7084 37232
rect 7124 37192 7133 37232
rect 7660 37148 7700 37276
rect 13132 37232 13172 37360
rect 19084 37316 19124 37360
rect 15235 37276 15244 37316
rect 15284 37276 17164 37316
rect 17204 37276 17213 37316
rect 17539 37276 17548 37316
rect 17588 37276 19124 37316
rect 21510 37232 21600 37252
rect 7747 37192 7756 37232
rect 7796 37192 7805 37232
rect 8105 37192 8236 37232
rect 8276 37192 8285 37232
rect 9091 37192 9100 37232
rect 9140 37192 9149 37232
rect 13132 37192 14860 37232
rect 14900 37192 14909 37232
rect 15427 37192 15436 37232
rect 15476 37192 15485 37232
rect 17251 37192 17260 37232
rect 17300 37192 17404 37232
rect 17444 37192 17453 37232
rect 18115 37192 18124 37232
rect 18164 37192 20275 37232
rect 20315 37192 20324 37232
rect 21283 37192 21292 37232
rect 21332 37192 21600 37232
rect 2860 37108 3668 37148
rect 4108 37108 7700 37148
rect 0 37064 90 37084
rect 2860 37064 2900 37108
rect 0 37024 2900 37064
rect 3679 37024 3688 37064
rect 3728 37024 3770 37064
rect 3810 37024 3852 37064
rect 3892 37024 3934 37064
rect 3974 37024 4016 37064
rect 4056 37024 4065 37064
rect 0 37004 90 37024
rect 4108 36980 4148 37108
rect 2860 36940 4148 36980
rect 4204 36940 5452 36980
rect 5492 36940 5501 36980
rect 2860 36896 2900 36940
rect 4204 36896 4244 36940
rect 1843 36856 1852 36896
rect 1892 36856 2900 36896
rect 2956 36856 4244 36896
rect 0 36728 90 36748
rect 2956 36728 2996 36856
rect 7756 36812 7796 37192
rect 7939 36856 7948 36896
rect 7988 36856 8119 36896
rect 3043 36772 3052 36812
rect 3092 36772 6796 36812
rect 6836 36772 6845 36812
rect 7756 36772 8372 36812
rect 0 36688 652 36728
rect 692 36688 701 36728
rect 1097 36688 1228 36728
rect 1268 36688 1277 36728
rect 1481 36688 1612 36728
rect 1652 36688 1661 36728
rect 2284 36688 2572 36728
rect 2612 36688 2621 36728
rect 2755 36688 2764 36728
rect 2804 36688 2996 36728
rect 3340 36688 3628 36728
rect 3668 36688 4204 36728
rect 4244 36688 4253 36728
rect 0 36668 90 36688
rect 2284 36644 2324 36688
rect 3340 36644 3380 36688
rect 4876 36644 4916 36772
rect 8105 36688 8227 36728
rect 8276 36688 8285 36728
rect 6124 36644 6164 36653
rect 7756 36644 7796 36653
rect 8332 36644 8372 36772
rect 9100 36644 9140 37192
rect 15436 37064 15476 37192
rect 21510 37172 21600 37192
rect 18211 37108 18220 37148
rect 18260 37108 19948 37148
rect 19988 37108 19997 37148
rect 15340 37024 15476 37064
rect 18799 37024 18808 37064
rect 18848 37024 18890 37064
rect 18930 37024 18972 37064
rect 19012 37024 19054 37064
rect 19094 37024 19136 37064
rect 19176 37024 19185 37064
rect 12355 36772 12364 36812
rect 12404 36772 14328 36812
rect 14851 36772 14860 36812
rect 14900 36772 14909 36812
rect 9475 36688 9484 36728
rect 9524 36688 9772 36728
rect 9812 36688 9821 36728
rect 10156 36688 11788 36728
rect 11828 36688 11837 36728
rect 13577 36688 13708 36728
rect 13748 36688 13757 36728
rect 9292 36644 9332 36653
rect 2266 36604 2275 36644
rect 2315 36604 2324 36644
rect 2371 36604 2380 36644
rect 2420 36604 2551 36644
rect 2851 36604 2860 36644
rect 2900 36604 3284 36644
rect 1459 36520 1468 36560
rect 1508 36520 2900 36560
rect 0 36392 90 36412
rect 0 36352 1420 36392
rect 1460 36352 1469 36392
rect 0 36332 90 36352
rect 2860 36224 2900 36520
rect 3244 36476 3284 36604
rect 3523 36604 3532 36644
rect 3572 36604 3828 36644
rect 3868 36604 3877 36644
rect 4867 36604 4876 36644
rect 4916 36604 4925 36644
rect 5993 36604 6124 36644
rect 6164 36604 6173 36644
rect 6499 36604 6508 36644
rect 6548 36604 6700 36644
rect 6740 36604 6749 36644
rect 7625 36604 7756 36644
rect 7796 36604 7805 36644
rect 7852 36604 8087 36644
rect 8127 36604 8136 36644
rect 8323 36604 8332 36644
rect 8372 36604 8381 36644
rect 8794 36604 8803 36644
rect 8843 36604 9140 36644
rect 9283 36604 9292 36644
rect 9332 36604 9463 36644
rect 9859 36604 9868 36644
rect 9908 36604 9964 36644
rect 10004 36604 10039 36644
rect 3340 36595 3380 36604
rect 6124 36595 6164 36604
rect 7756 36595 7796 36604
rect 3436 36520 3820 36560
rect 3860 36520 4148 36560
rect 4435 36520 4444 36560
rect 4484 36520 4684 36560
rect 4724 36520 4733 36560
rect 3436 36476 3476 36520
rect 4108 36476 4148 36520
rect 7852 36476 7892 36604
rect 9292 36595 9332 36604
rect 8602 36520 8611 36560
rect 8651 36520 9100 36560
rect 9140 36520 9149 36560
rect 3244 36436 3476 36476
rect 4003 36436 4012 36476
rect 4052 36436 4061 36476
rect 4108 36436 6124 36476
rect 6164 36436 6173 36476
rect 6307 36436 6316 36476
rect 6356 36436 7660 36476
rect 7700 36436 7892 36476
rect 8297 36436 8419 36476
rect 8468 36436 8477 36476
rect 4012 36392 4052 36436
rect 10156 36392 10196 36688
rect 14288 36663 14328 36772
rect 14860 36728 14900 36772
rect 14851 36688 14860 36728
rect 14900 36688 14947 36728
rect 12172 36644 12212 36653
rect 13228 36644 13268 36653
rect 10243 36604 10252 36644
rect 10292 36604 10301 36644
rect 10361 36604 10370 36644
rect 10410 36604 10444 36644
rect 10484 36604 10550 36644
rect 10793 36604 10924 36644
rect 10964 36604 10973 36644
rect 11683 36604 11692 36644
rect 11732 36604 11884 36644
rect 11924 36604 12172 36644
rect 12259 36604 12268 36644
rect 12308 36604 12739 36644
rect 12779 36604 12788 36644
rect 13268 36604 13612 36644
rect 13652 36604 13661 36644
rect 13795 36604 13804 36644
rect 13844 36604 13975 36644
rect 14179 36604 14188 36644
rect 14228 36604 14237 36644
rect 14288 36623 14301 36663
rect 14341 36623 14350 36663
rect 15340 36644 15380 37024
rect 15715 36940 15724 36980
rect 15764 36940 20852 36980
rect 15811 36856 15820 36896
rect 15860 36856 18364 36896
rect 18404 36856 18413 36896
rect 20131 36856 20140 36896
rect 20180 36856 20524 36896
rect 20564 36856 20573 36896
rect 16012 36772 17548 36812
rect 17588 36772 17597 36812
rect 17740 36772 18548 36812
rect 16012 36728 16052 36772
rect 17260 36728 17300 36772
rect 17740 36728 17780 36772
rect 15820 36688 16012 36728
rect 16052 36688 16061 36728
rect 17260 36688 17396 36728
rect 17731 36688 17740 36728
rect 17780 36688 17789 36728
rect 14537 36604 14668 36644
rect 14708 36604 14717 36644
rect 15340 36604 15523 36644
rect 15563 36604 15572 36644
rect 15619 36604 15628 36644
rect 15668 36604 15677 36644
rect 4012 36352 6988 36392
rect 7028 36352 7037 36392
rect 7267 36352 7276 36392
rect 7316 36352 10196 36392
rect 10252 36308 10292 36604
rect 12172 36595 12212 36604
rect 13228 36595 13268 36604
rect 14188 36560 14228 36604
rect 15628 36560 15668 36604
rect 14188 36520 14956 36560
rect 14996 36520 15668 36560
rect 12067 36436 12076 36476
rect 12116 36436 12556 36476
rect 12596 36436 12605 36476
rect 12931 36436 12940 36476
rect 12980 36436 14524 36476
rect 14564 36436 14573 36476
rect 15091 36436 15100 36476
rect 15140 36436 15244 36476
rect 15284 36436 15293 36476
rect 15820 36392 15860 36688
rect 16588 36644 16628 36653
rect 17356 36644 17396 36688
rect 18220 36644 18260 36653
rect 18508 36644 18548 36772
rect 20812 36728 20852 36940
rect 21510 36728 21600 36748
rect 18595 36688 18604 36728
rect 18644 36688 18653 36728
rect 20812 36688 21600 36728
rect 18604 36644 18644 36688
rect 21510 36668 21600 36688
rect 19948 36644 19988 36653
rect 15907 36604 15916 36644
rect 15956 36604 16108 36644
rect 16148 36604 16157 36644
rect 16291 36604 16300 36644
rect 16340 36604 16588 36644
rect 17098 36604 17107 36644
rect 17147 36604 17260 36644
rect 17300 36604 17309 36644
rect 17356 36604 17399 36644
rect 17439 36604 17448 36644
rect 17530 36604 17539 36644
rect 17579 36604 17588 36644
rect 17635 36604 17644 36644
rect 17684 36604 17740 36644
rect 17780 36604 17815 36644
rect 18089 36604 18220 36644
rect 18260 36604 18269 36644
rect 18499 36604 18508 36644
rect 18548 36604 18557 36644
rect 18604 36604 18700 36644
rect 18740 36604 18749 36644
rect 18883 36604 18892 36644
rect 18932 36604 19948 36644
rect 16588 36595 16628 36604
rect 17548 36560 17588 36604
rect 18220 36595 18260 36604
rect 17155 36520 17164 36560
rect 17204 36520 17444 36560
rect 17501 36520 17548 36560
rect 17588 36520 17597 36560
rect 17909 36520 17918 36560
rect 17958 36520 17967 36560
rect 17404 36476 17444 36520
rect 17918 36476 17958 36520
rect 17251 36436 17260 36476
rect 17300 36436 17309 36476
rect 17404 36436 17958 36476
rect 18010 36436 18019 36476
rect 18059 36436 18068 36476
rect 18115 36436 18124 36476
rect 18164 36436 18212 36476
rect 12835 36352 12844 36392
rect 12884 36352 15860 36392
rect 4919 36268 4928 36308
rect 4968 36268 5010 36308
rect 5050 36268 5092 36308
rect 5132 36268 5174 36308
rect 5214 36268 5256 36308
rect 5296 36268 5305 36308
rect 8803 36268 8812 36308
rect 8852 36268 10292 36308
rect 17260 36308 17300 36436
rect 17260 36268 17836 36308
rect 17876 36268 17885 36308
rect 2860 36184 4148 36224
rect 4483 36184 4492 36224
rect 4532 36184 5644 36224
rect 5684 36184 10540 36224
rect 10580 36184 10924 36224
rect 10964 36184 10973 36224
rect 13987 36184 13996 36224
rect 14036 36184 14860 36224
rect 14900 36184 14909 36224
rect 15052 36184 16588 36224
rect 16628 36184 16637 36224
rect 4108 36140 4148 36184
rect 3043 36100 3052 36140
rect 3092 36100 3340 36140
rect 3380 36100 3389 36140
rect 3881 36100 4012 36140
rect 4052 36100 4061 36140
rect 4108 36100 5972 36140
rect 6691 36100 6700 36140
rect 6740 36100 10196 36140
rect 11587 36100 11596 36140
rect 11636 36100 12268 36140
rect 12308 36100 12317 36140
rect 12730 36100 12739 36140
rect 12779 36100 13612 36140
rect 13652 36100 13661 36140
rect 0 36056 90 36076
rect 5932 36056 5972 36100
rect 10156 36056 10196 36100
rect 0 36016 1228 36056
rect 1268 36016 1277 36056
rect 1699 36016 1708 36056
rect 1748 36016 4108 36056
rect 4148 36016 4157 36056
rect 4579 36016 4588 36056
rect 4628 36016 4637 36056
rect 5644 36016 5865 36056
rect 5932 36016 7276 36056
rect 7316 36016 7325 36056
rect 7747 36016 7756 36056
rect 7796 36016 9812 36056
rect 0 35996 90 36016
rect 4588 35972 4628 36016
rect 5644 35972 5684 36016
rect 5825 35972 5865 36016
rect 835 35932 844 35972
rect 884 35932 1652 35972
rect 2153 35932 2188 35972
rect 2228 35932 2275 35972
rect 2315 35932 2333 35972
rect 2376 35932 2385 35972
rect 2425 35932 2434 35972
rect 2633 35932 2764 35972
rect 2804 35932 2813 35972
rect 3340 35963 3380 35972
rect 1612 35888 1652 35932
rect 2380 35888 2420 35932
rect 3427 35932 3436 35972
rect 3476 35963 3860 35972
rect 3476 35932 3820 35963
rect 3340 35888 3380 35923
rect 4361 35932 4492 35972
rect 4532 35932 4541 35972
rect 4588 35932 5684 35972
rect 5740 35963 5780 35972
rect 3820 35914 3860 35923
rect 5825 35932 6124 35972
rect 6164 35932 6173 35972
rect 6298 35932 6307 35972
rect 6356 35932 6487 35972
rect 6604 35932 6892 35972
rect 6932 35932 6941 35972
rect 8140 35963 8180 36016
rect 9772 35972 9812 36016
rect 10156 36016 11500 36056
rect 11540 36016 11549 36056
rect 11866 36016 11875 36056
rect 11915 36016 12307 36056
rect 10156 35972 10196 36016
rect 12267 35972 12307 36016
rect 12364 36016 13420 36056
rect 13460 36016 13469 36056
rect 5740 35888 5780 35923
rect 6604 35888 6644 35932
rect 8227 35932 8236 35972
rect 8276 35932 8524 35972
rect 8564 35932 8573 35972
rect 9641 35932 9772 35972
rect 9812 35932 9821 35972
rect 10147 35932 10156 35972
rect 10196 35932 10205 35972
rect 11107 35932 11116 35972
rect 11156 35963 11444 35972
rect 11156 35932 11404 35963
rect 8140 35914 8180 35923
rect 9772 35914 9812 35923
rect 11657 35932 11788 35972
rect 11828 35932 11837 35972
rect 11962 35932 11971 35972
rect 12011 35932 12020 35972
rect 11404 35914 11444 35923
rect 11980 35888 12020 35932
rect 12074 35900 12083 35940
rect 12123 35900 12132 35940
rect 12250 35932 12259 35972
rect 12299 35932 12308 35972
rect 12364 35963 12404 36016
rect 15052 35972 15092 36184
rect 12364 35914 12404 35923
rect 12503 35963 12548 35972
rect 12503 35923 12508 35963
rect 12630 35932 12639 35972
rect 12679 35932 12692 35972
rect 12739 35932 12748 35972
rect 12817 35932 12919 35972
rect 13027 35932 13036 35972
rect 13076 35932 13085 35972
rect 13315 35932 13324 35972
rect 13364 35963 15092 35972
rect 13364 35932 14284 35963
rect 12503 35914 12548 35923
rect 739 35848 748 35888
rect 788 35848 1228 35888
rect 1268 35848 1277 35888
rect 1603 35848 1612 35888
rect 1652 35848 1661 35888
rect 2275 35848 2284 35888
rect 2324 35848 2420 35888
rect 2851 35848 2860 35888
rect 2900 35848 2909 35888
rect 3340 35848 3628 35888
rect 3668 35848 3677 35888
rect 5740 35848 6068 35888
rect 6115 35848 6124 35888
rect 6164 35848 6644 35888
rect 6691 35848 6700 35888
rect 6740 35848 6796 35888
rect 6836 35848 6871 35888
rect 11849 35848 11980 35888
rect 12020 35848 12029 35888
rect 2860 35804 2900 35848
rect 2860 35764 3340 35804
rect 3380 35764 3820 35804
rect 3860 35764 3869 35804
rect 5731 35764 5740 35804
rect 5780 35764 5932 35804
rect 5972 35764 5981 35804
rect 0 35720 90 35740
rect 0 35680 844 35720
rect 884 35680 893 35720
rect 1459 35680 1468 35720
rect 1508 35680 1748 35720
rect 1843 35680 1852 35720
rect 1892 35680 2380 35720
rect 2420 35680 2429 35720
rect 0 35660 90 35680
rect 1708 35468 1748 35680
rect 6028 35552 6068 35848
rect 6298 35764 6307 35804
rect 6347 35764 8044 35804
rect 8084 35764 8093 35804
rect 6451 35680 6460 35720
rect 6500 35680 6509 35720
rect 8323 35680 8332 35720
rect 8372 35680 9908 35720
rect 9955 35680 9964 35720
rect 10004 35680 10924 35720
rect 10964 35680 10973 35720
rect 6460 35636 6500 35680
rect 9868 35636 9908 35680
rect 11980 35636 12020 35848
rect 6460 35596 9004 35636
rect 9044 35596 9053 35636
rect 9868 35596 12020 35636
rect 12076 35804 12116 35900
rect 12503 35804 12543 35914
rect 12652 35888 12692 35932
rect 12652 35848 12940 35888
rect 12980 35848 12989 35888
rect 12076 35764 12543 35804
rect 12076 35552 12116 35764
rect 13036 35720 13076 35932
rect 14324 35932 15092 35963
rect 15148 36100 15724 36140
rect 15764 36100 15773 36140
rect 17635 36100 17644 36140
rect 17684 36100 17827 36140
rect 17867 36100 17876 36140
rect 14284 35914 14324 35923
rect 15148 35888 15188 36100
rect 15235 36016 15244 36056
rect 15284 36016 16244 36056
rect 16291 36016 16300 36056
rect 16340 36016 17932 36056
rect 17972 36016 17981 36056
rect 16204 35972 16244 36016
rect 15427 35932 15436 35972
rect 15476 35932 15572 35972
rect 15689 35932 15724 35972
rect 15764 35932 15820 35972
rect 15860 35932 15869 35972
rect 16099 35932 16108 35972
rect 16148 35932 16157 35972
rect 16204 35963 17396 35972
rect 16204 35932 17356 35963
rect 15532 35888 15572 35932
rect 15955 35890 15964 35930
rect 16004 35890 16052 35930
rect 14813 35848 14860 35888
rect 14900 35848 14909 35888
rect 15091 35848 15100 35888
rect 15140 35848 15188 35888
rect 15427 35848 15436 35888
rect 15476 35848 15485 35888
rect 15532 35848 15628 35888
rect 15668 35848 15677 35888
rect 15834 35848 15843 35888
rect 15883 35848 15892 35888
rect 14860 35804 14900 35848
rect 14563 35764 14572 35804
rect 14612 35764 14621 35804
rect 14851 35764 14860 35804
rect 14900 35764 14909 35804
rect 14572 35720 14612 35764
rect 12547 35680 12556 35720
rect 12596 35680 13076 35720
rect 14467 35680 14476 35720
rect 14516 35680 14525 35720
rect 14572 35680 15196 35720
rect 15236 35680 15245 35720
rect 3679 35512 3688 35552
rect 3728 35512 3770 35552
rect 3810 35512 3852 35552
rect 3892 35512 3934 35552
rect 3974 35512 4016 35552
rect 4056 35512 4065 35552
rect 5155 35512 5164 35552
rect 5204 35512 7276 35552
rect 7316 35512 7325 35552
rect 10060 35512 12116 35552
rect 10060 35468 10100 35512
rect 1708 35428 4492 35468
rect 4532 35428 4541 35468
rect 6787 35428 6796 35468
rect 6836 35428 9620 35468
rect 0 35384 90 35404
rect 0 35344 172 35384
rect 212 35344 221 35384
rect 3401 35344 3532 35384
rect 3572 35344 3581 35384
rect 4195 35344 4204 35384
rect 4244 35344 5356 35384
rect 5396 35344 5405 35384
rect 6595 35344 6604 35384
rect 6644 35344 6988 35384
rect 7028 35344 7037 35384
rect 8035 35344 8044 35384
rect 8084 35344 9292 35384
rect 9332 35344 9341 35384
rect 0 35324 90 35344
rect 9580 35300 9620 35428
rect 9676 35428 10100 35468
rect 9676 35384 9716 35428
rect 9667 35344 9676 35384
rect 9716 35344 9725 35384
rect 11273 35344 11404 35384
rect 11444 35344 11453 35384
rect 12844 35344 13324 35384
rect 13364 35344 13373 35384
rect 2371 35260 2380 35300
rect 2420 35260 3956 35300
rect 643 35176 652 35216
rect 692 35176 1228 35216
rect 1268 35176 1277 35216
rect 1411 35176 1420 35216
rect 1460 35176 1612 35216
rect 1652 35176 1661 35216
rect 3340 35132 3380 35141
rect 3916 35132 3956 35260
rect 6892 35260 9484 35300
rect 9524 35260 9533 35300
rect 9580 35260 12556 35300
rect 12596 35260 12605 35300
rect 5164 35132 5204 35141
rect 6796 35132 6836 35141
rect 1961 35092 2092 35132
rect 2132 35092 2900 35132
rect 0 35048 90 35068
rect 0 35008 1324 35048
rect 1364 35008 1373 35048
rect 1459 35008 1468 35048
rect 1508 35008 2380 35048
rect 2420 35008 2429 35048
rect 0 34988 90 35008
rect 2860 34964 2900 35092
rect 3881 35092 3916 35132
rect 3956 35092 4012 35132
rect 4052 35092 4061 35132
rect 5033 35092 5164 35132
rect 5204 35092 5213 35132
rect 5539 35092 5548 35132
rect 5588 35092 5836 35132
rect 5876 35092 5885 35132
rect 3340 35048 3380 35092
rect 5164 35083 5204 35092
rect 6796 35048 6836 35092
rect 2947 35008 2956 35048
rect 2996 35008 3380 35048
rect 5347 35008 5356 35048
rect 5396 35008 6836 35048
rect 6892 34964 6932 35260
rect 7315 35176 7324 35216
rect 7364 35176 7652 35216
rect 7747 35176 7756 35216
rect 7796 35176 7808 35216
rect 7612 35132 7652 35176
rect 7768 35132 7808 35176
rect 9484 35132 9524 35141
rect 11212 35132 11252 35141
rect 12844 35132 12884 35344
rect 14476 35300 14516 35680
rect 15436 35552 15476 35848
rect 15843 35804 15883 35848
rect 16012 35804 16052 35890
rect 16108 35888 16148 35932
rect 17539 35932 17548 35972
rect 17588 35932 17726 35972
rect 17766 35932 17775 35972
rect 18028 35963 18068 36436
rect 18172 36392 18212 36436
rect 18115 36352 18124 36392
rect 18164 36352 18212 36392
rect 19948 36140 19988 36604
rect 20039 36268 20048 36308
rect 20088 36268 20130 36308
rect 20170 36268 20212 36308
rect 20252 36268 20294 36308
rect 20334 36268 20376 36308
rect 20416 36268 20425 36308
rect 21510 36224 21600 36244
rect 20899 36184 20908 36224
rect 20948 36184 21600 36224
rect 21510 36164 21600 36184
rect 19948 36100 20044 36140
rect 20084 36100 20093 36140
rect 18403 36016 18412 36056
rect 18452 36016 18740 36056
rect 19171 36016 19180 36056
rect 19220 36016 19700 36056
rect 18700 35972 18740 36016
rect 17356 35914 17396 35923
rect 18307 35932 18316 35972
rect 18356 35932 18365 35972
rect 18586 35932 18595 35972
rect 18635 35932 18644 35972
rect 18691 35932 18700 35972
rect 18740 35932 18749 35972
rect 19075 35932 19084 35972
rect 19124 35932 19276 35972
rect 19316 35932 19325 35972
rect 19660 35963 19700 36016
rect 18028 35914 18068 35923
rect 16108 35848 16780 35888
rect 16820 35848 16829 35888
rect 18316 35804 18356 35932
rect 18604 35888 18644 35932
rect 19660 35914 19700 35923
rect 20140 35963 20276 35972
rect 20180 35932 20276 35963
rect 20362 35932 20371 35972
rect 20411 35932 20812 35972
rect 20852 35932 20861 35972
rect 20140 35914 20180 35923
rect 18604 35848 18700 35888
rect 18740 35848 18749 35888
rect 19075 35848 19084 35888
rect 19124 35848 19180 35888
rect 19220 35848 19255 35888
rect 15843 35764 15956 35804
rect 16012 35764 16300 35804
rect 16340 35764 16349 35804
rect 17251 35764 17260 35804
rect 17300 35764 17548 35804
rect 17588 35764 17597 35804
rect 18019 35764 18028 35804
rect 18068 35764 18356 35804
rect 15916 35636 15956 35764
rect 18124 35680 18172 35720
rect 18212 35680 18221 35720
rect 15907 35596 15916 35636
rect 15956 35596 15965 35636
rect 14851 35512 14860 35552
rect 14900 35512 15476 35552
rect 18124 35468 18164 35680
rect 18799 35512 18808 35552
rect 18848 35512 18890 35552
rect 18930 35512 18972 35552
rect 19012 35512 19054 35552
rect 19094 35512 19136 35552
rect 19176 35512 19185 35552
rect 16108 35428 16300 35468
rect 16340 35428 18164 35468
rect 14755 35344 14764 35384
rect 14804 35344 15244 35384
rect 15284 35344 15572 35384
rect 13027 35260 13036 35300
rect 13076 35260 13085 35300
rect 14476 35260 14996 35300
rect 13036 35216 13076 35260
rect 13036 35176 13844 35216
rect 14249 35176 14284 35216
rect 14324 35176 14380 35216
rect 14420 35176 14429 35216
rect 13804 35132 13844 35176
rect 14860 35132 14900 35141
rect 7049 35092 7180 35132
rect 7220 35092 7229 35132
rect 7370 35092 7468 35132
rect 7532 35092 7550 35132
rect 7612 35092 7651 35132
rect 7691 35092 7700 35132
rect 7759 35092 7768 35132
rect 7808 35092 7843 35132
rect 7930 35092 7939 35132
rect 7979 35092 7988 35132
rect 8032 35092 8041 35132
rect 8084 35092 8215 35132
rect 8259 35092 8268 35132
rect 8308 35092 8317 35132
rect 7180 35048 7220 35092
rect 7948 35048 7988 35092
rect 8277 35048 8317 35092
rect 9524 35092 9772 35132
rect 9812 35092 9821 35132
rect 9955 35092 9964 35132
rect 10004 35092 10013 35132
rect 10339 35092 10348 35132
rect 10388 35092 11212 35132
rect 11587 35092 11596 35132
rect 11636 35092 11645 35132
rect 13027 35092 13036 35132
rect 13076 35092 13228 35132
rect 13268 35092 13277 35132
rect 13324 35092 13367 35132
rect 13407 35092 13416 35132
rect 13786 35092 13795 35132
rect 13835 35092 13844 35132
rect 13891 35092 13900 35132
rect 13940 35092 13949 35132
rect 14371 35092 14380 35132
rect 14420 35092 14764 35132
rect 14804 35092 14813 35132
rect 14956 35132 14996 35260
rect 15532 35132 15572 35344
rect 16108 35300 16148 35428
rect 20236 35384 20276 35932
rect 21510 35720 21600 35740
rect 21091 35680 21100 35720
rect 21140 35680 21600 35720
rect 21510 35660 21600 35680
rect 17923 35344 17932 35384
rect 17972 35344 18220 35384
rect 18260 35344 18269 35384
rect 20227 35344 20236 35384
rect 20276 35344 20285 35384
rect 16012 35260 16148 35300
rect 16675 35260 16684 35300
rect 16724 35260 17644 35300
rect 17684 35260 18644 35300
rect 19555 35260 19564 35300
rect 19604 35260 21100 35300
rect 21140 35260 21149 35300
rect 16012 35132 16052 35260
rect 16156 35176 16300 35216
rect 16340 35176 16349 35216
rect 16483 35176 16492 35216
rect 16532 35176 16771 35216
rect 16811 35176 16820 35216
rect 17129 35176 17260 35216
rect 17300 35176 17684 35216
rect 17827 35176 17836 35216
rect 17876 35176 18316 35216
rect 18356 35176 18365 35216
rect 16156 35132 16196 35176
rect 17260 35132 17300 35176
rect 17644 35132 17684 35176
rect 18604 35132 18644 35260
rect 21510 35216 21600 35236
rect 20515 35176 20524 35216
rect 20564 35176 21600 35216
rect 21510 35156 21600 35176
rect 20044 35132 20084 35141
rect 14956 35092 15348 35132
rect 15388 35092 15397 35132
rect 15532 35092 15820 35132
rect 15860 35092 15869 35132
rect 16003 35092 16012 35132
rect 16052 35092 16061 35132
rect 16147 35092 16156 35132
rect 16196 35092 16205 35132
rect 16282 35092 16291 35132
rect 16331 35092 16340 35132
rect 16387 35092 16396 35132
rect 16436 35092 16445 35132
rect 16500 35092 16588 35132
rect 16628 35092 16631 35132
rect 16671 35092 16680 35132
rect 16771 35092 16780 35132
rect 16820 35092 16876 35132
rect 16916 35092 16951 35132
rect 17251 35092 17260 35132
rect 17300 35092 17309 35132
rect 17530 35092 17539 35132
rect 17579 35092 17588 35132
rect 17644 35092 18028 35132
rect 18068 35092 18077 35132
rect 18595 35092 18604 35132
rect 18644 35092 18653 35132
rect 18761 35092 18796 35132
rect 18836 35092 18892 35132
rect 18932 35092 18941 35132
rect 9484 35083 9524 35092
rect 7180 35008 7892 35048
rect 7939 35008 7948 35048
rect 7988 35008 8035 35048
rect 8227 35008 8236 35048
rect 8276 35008 8317 35048
rect 7852 34964 7892 35008
rect 9964 34964 10004 35092
rect 11212 35083 11252 35092
rect 11596 34964 11636 35092
rect 12844 35083 12884 35092
rect 13324 35048 13364 35092
rect 13900 35048 13940 35092
rect 14860 35048 14900 35092
rect 13315 35008 13324 35048
rect 13364 35008 13373 35048
rect 13900 35008 14284 35048
rect 14324 35008 14333 35048
rect 14659 35008 14668 35048
rect 14708 35008 15860 35048
rect 15907 35008 15916 35048
rect 15956 35008 16087 35048
rect 15820 34964 15860 35008
rect 16300 34964 16340 35092
rect 16396 35048 16436 35092
rect 17548 35048 17588 35092
rect 20044 35048 20084 35092
rect 16396 35008 16684 35048
rect 16724 35008 16733 35048
rect 16780 35008 17588 35048
rect 17635 35008 17644 35048
rect 17684 35008 17693 35048
rect 17884 35008 18076 35048
rect 18116 35008 18125 35048
rect 18211 35008 18220 35048
rect 18260 35008 20084 35048
rect 1843 34924 1852 34964
rect 1892 34924 1901 34964
rect 2860 34924 6124 34964
rect 6164 34924 6173 34964
rect 6220 34924 6932 34964
rect 7546 34924 7555 34964
rect 7595 34924 7604 34964
rect 7843 34924 7852 34964
rect 7892 34924 7901 34964
rect 9091 34924 9100 34964
rect 9140 34924 10004 34964
rect 10060 34924 11636 34964
rect 13385 34924 13420 34964
rect 13460 34924 13516 34964
rect 13556 34924 13565 34964
rect 15497 34924 15532 34964
rect 15572 34924 15628 34964
rect 15668 34924 15677 34964
rect 15820 34924 16340 34964
rect 0 34712 90 34732
rect 1852 34712 1892 34924
rect 6220 34880 6260 34924
rect 7564 34880 7604 34924
rect 10060 34880 10100 34924
rect 16780 34880 16820 35008
rect 16954 34924 16963 34964
rect 17003 34924 17452 34964
rect 17492 34924 17501 34964
rect 2755 34840 2764 34880
rect 2804 34840 6260 34880
rect 6307 34840 6316 34880
rect 6356 34840 7604 34880
rect 8899 34840 8908 34880
rect 8948 34840 10100 34880
rect 12547 34840 12556 34880
rect 12596 34840 13324 34880
rect 13364 34840 13373 34880
rect 14947 34840 14956 34880
rect 14996 34840 16820 34880
rect 17644 34880 17684 35008
rect 17884 34964 17924 35008
rect 17827 34924 17836 34964
rect 17876 34924 17924 34964
rect 18115 34924 18124 34964
rect 18164 34924 18460 34964
rect 18500 34924 18509 34964
rect 19948 34924 20044 34964
rect 20084 34924 20093 34964
rect 17644 34840 18316 34880
rect 18356 34840 18365 34880
rect 4919 34756 4928 34796
rect 4968 34756 5010 34796
rect 5050 34756 5092 34796
rect 5132 34756 5174 34796
rect 5214 34756 5256 34796
rect 5296 34756 5305 34796
rect 6691 34756 6700 34796
rect 6740 34756 8660 34796
rect 15235 34756 15244 34796
rect 15284 34756 15628 34796
rect 15668 34756 15677 34796
rect 8620 34712 8660 34756
rect 17644 34712 17684 34840
rect 0 34672 1612 34712
rect 1652 34672 1661 34712
rect 1852 34672 5836 34712
rect 5876 34672 5885 34712
rect 8620 34672 17684 34712
rect 0 34652 90 34672
rect 18412 34628 18452 34924
rect 2659 34588 2668 34628
rect 2708 34588 2717 34628
rect 7276 34588 9196 34628
rect 9236 34588 9245 34628
rect 12067 34588 12076 34628
rect 12116 34588 12980 34628
rect 17242 34588 17251 34628
rect 17291 34588 18452 34628
rect 19948 34628 19988 34924
rect 20039 34756 20048 34796
rect 20088 34756 20130 34796
rect 20170 34756 20212 34796
rect 20252 34756 20294 34796
rect 20334 34756 20376 34796
rect 20416 34756 20425 34796
rect 21510 34712 21600 34732
rect 20995 34672 21004 34712
rect 21044 34672 21600 34712
rect 21510 34652 21600 34672
rect 19948 34588 20044 34628
rect 20084 34588 20093 34628
rect 2668 34544 2708 34588
rect 2668 34504 2996 34544
rect 2956 34460 2996 34504
rect 3340 34504 5740 34544
rect 5780 34504 5789 34544
rect 3340 34460 3380 34504
rect 7276 34460 7316 34588
rect 12940 34544 12980 34588
rect 8803 34504 8812 34544
rect 8852 34504 10348 34544
rect 10388 34504 10397 34544
rect 11004 34504 11116 34544
rect 11195 34504 11596 34544
rect 11636 34504 11645 34544
rect 12307 34504 12316 34544
rect 12356 34504 12460 34544
rect 12500 34504 12509 34544
rect 12931 34504 12940 34544
rect 12980 34504 12989 34544
rect 13891 34504 13900 34544
rect 13940 34504 13949 34544
rect 14220 34504 14284 34544
rect 14324 34504 14764 34544
rect 14804 34504 14956 34544
rect 14996 34504 15005 34544
rect 16627 34504 16636 34544
rect 16676 34504 17300 34544
rect 17443 34504 17452 34544
rect 17503 34504 17623 34544
rect 18691 34504 18700 34544
rect 18740 34504 19084 34544
rect 19124 34504 19133 34544
rect 19529 34504 19612 34544
rect 19652 34504 19660 34544
rect 19700 34504 19709 34544
rect 19843 34504 19852 34544
rect 19892 34504 19996 34544
rect 20036 34504 20045 34544
rect 20371 34504 20380 34544
rect 20420 34504 20620 34544
rect 20660 34504 20669 34544
rect 13900 34460 13940 34504
rect 14380 34460 14420 34504
rect 835 34420 844 34460
rect 884 34420 1652 34460
rect 2153 34420 2275 34460
rect 2324 34420 2333 34460
rect 2537 34420 2572 34460
rect 2612 34420 2668 34460
rect 2708 34420 2717 34460
rect 2842 34420 2851 34460
rect 2891 34420 2900 34460
rect 2947 34420 2956 34460
rect 2996 34420 3005 34460
rect 3331 34420 3340 34460
rect 3380 34420 3389 34460
rect 3523 34420 3532 34460
rect 3572 34451 3956 34460
rect 3572 34420 3916 34451
rect 0 34376 90 34396
rect 1612 34376 1652 34420
rect 2860 34376 2900 34420
rect 0 34336 460 34376
rect 500 34336 509 34376
rect 1097 34336 1228 34376
rect 1268 34336 1277 34376
rect 1603 34336 1612 34376
rect 1652 34336 1661 34376
rect 1843 34336 1852 34376
rect 1892 34336 2476 34376
rect 2516 34336 2525 34376
rect 2860 34336 2956 34376
rect 2996 34336 3005 34376
rect 0 34316 90 34336
rect 3340 34292 3380 34420
rect 4265 34420 4396 34460
rect 4436 34420 4445 34460
rect 5251 34420 5260 34460
rect 5300 34420 5309 34460
rect 6019 34420 6028 34460
rect 6068 34420 6077 34460
rect 7145 34420 7276 34460
rect 7316 34420 7325 34460
rect 7555 34420 7564 34460
rect 7604 34420 7660 34460
rect 7700 34420 7735 34460
rect 8777 34420 8908 34460
rect 8948 34420 8957 34460
rect 9370 34420 9379 34460
rect 9419 34420 9428 34460
rect 9475 34420 9484 34460
rect 9524 34420 9580 34460
rect 9620 34420 9655 34460
rect 9859 34420 9868 34460
rect 9908 34420 10060 34460
rect 10100 34420 10109 34460
rect 10313 34420 10444 34460
rect 10484 34420 10493 34460
rect 10793 34420 10924 34460
rect 10964 34420 10973 34460
rect 11971 34420 11980 34460
rect 12020 34420 12460 34460
rect 12500 34420 12509 34460
rect 13708 34451 13844 34460
rect 3916 34402 3956 34411
rect 4396 34402 4436 34411
rect 5260 34376 5300 34420
rect 6028 34376 6068 34420
rect 7276 34402 7316 34411
rect 8908 34402 8948 34411
rect 3427 34336 3436 34376
rect 3476 34336 3860 34376
rect 4618 34336 4627 34376
rect 4667 34336 4780 34376
rect 4820 34336 4829 34376
rect 4963 34336 4972 34376
rect 5012 34336 5164 34376
rect 5204 34336 5213 34376
rect 5260 34336 5404 34376
rect 5444 34336 5453 34376
rect 5801 34336 5836 34376
rect 5876 34336 5932 34376
rect 5972 34336 6068 34376
rect 2083 34252 2092 34292
rect 2132 34252 3380 34292
rect 3820 34292 3860 34336
rect 9388 34292 9428 34420
rect 10444 34402 10484 34411
rect 10924 34402 10964 34411
rect 13748 34420 13844 34451
rect 13900 34420 14275 34460
rect 14315 34420 14324 34460
rect 14371 34420 14380 34460
rect 14420 34420 14429 34460
rect 14476 34420 14764 34460
rect 14804 34420 14813 34460
rect 15235 34420 15244 34460
rect 15284 34451 15415 34460
rect 15284 34420 15340 34451
rect 13708 34402 13748 34411
rect 9955 34336 9964 34376
rect 10004 34336 10252 34376
rect 10292 34336 10301 34376
rect 11945 34336 12076 34376
rect 12116 34336 12556 34376
rect 12596 34336 12605 34376
rect 3820 34252 4780 34292
rect 4820 34252 4829 34292
rect 5011 34252 5020 34292
rect 5060 34252 5740 34292
rect 5780 34252 5789 34292
rect 9004 34252 9428 34292
rect 13804 34292 13844 34420
rect 14476 34376 14516 34420
rect 15380 34420 15415 34451
rect 15820 34451 15860 34460
rect 15340 34402 15380 34411
rect 16003 34420 16012 34460
rect 16052 34420 16820 34460
rect 14371 34336 14380 34376
rect 14420 34336 14516 34376
rect 14729 34336 14860 34376
rect 14900 34336 14909 34376
rect 13804 34252 15436 34292
rect 15476 34252 15485 34292
rect 1459 34168 1468 34208
rect 1508 34168 1996 34208
rect 2036 34168 2045 34208
rect 2563 34168 2572 34208
rect 2612 34168 3340 34208
rect 3380 34168 3389 34208
rect 5587 34168 5596 34208
rect 5636 34168 5645 34208
rect 7337 34168 7468 34208
rect 7508 34168 7517 34208
rect 5596 34124 5636 34168
rect 4291 34084 4300 34124
rect 4340 34084 5932 34124
rect 5972 34084 5981 34124
rect 0 34040 90 34060
rect 0 34000 1612 34040
rect 1652 34000 1661 34040
rect 3679 34000 3688 34040
rect 3728 34000 3770 34040
rect 3810 34000 3852 34040
rect 3892 34000 3934 34040
rect 3974 34000 4016 34040
rect 4056 34000 4065 34040
rect 4771 34000 4780 34040
rect 4820 34000 6604 34040
rect 6644 34000 6653 34040
rect 0 33980 90 34000
rect 6211 33916 6220 33956
rect 6260 33916 8428 33956
rect 8468 33916 8477 33956
rect 2563 33832 2572 33872
rect 2612 33832 2668 33872
rect 2708 33832 2743 33872
rect 5827 33832 5836 33872
rect 5876 33832 6412 33872
rect 6452 33832 6461 33872
rect 7459 33832 7468 33872
rect 7508 33832 7756 33872
rect 7796 33832 7805 33872
rect 1315 33748 1324 33788
rect 1364 33748 4052 33788
rect 0 33704 90 33724
rect 4012 33704 4052 33748
rect 4396 33748 6220 33788
rect 6260 33748 7700 33788
rect 0 33664 1996 33704
rect 2036 33664 2045 33704
rect 3148 33664 3532 33704
rect 3572 33664 3581 33704
rect 4003 33664 4012 33704
rect 4052 33664 4061 33704
rect 0 33644 90 33664
rect 3148 33662 3188 33664
rect 3136 33653 3188 33662
rect 2476 33620 2516 33629
rect 1123 33580 1132 33620
rect 1172 33580 1228 33620
rect 1268 33580 1303 33620
rect 2516 33580 2764 33620
rect 2804 33580 2813 33620
rect 3018 33580 3027 33620
rect 3067 33580 3092 33620
rect 3136 33613 3137 33653
rect 3177 33622 3188 33653
rect 3177 33613 3186 33622
rect 3820 33620 3860 33629
rect 4396 33620 4436 33748
rect 5644 33620 5684 33629
rect 7276 33620 7316 33629
rect 7660 33620 7700 33748
rect 8908 33620 8948 33629
rect 3136 33604 3186 33613
rect 3239 33580 3248 33620
rect 3288 33580 3820 33620
rect 4387 33580 4396 33620
rect 4436 33580 4445 33620
rect 6019 33580 6028 33620
rect 6068 33580 6796 33620
rect 6836 33580 6845 33620
rect 7145 33580 7276 33620
rect 7316 33580 7325 33620
rect 7651 33580 7660 33620
rect 7700 33580 7709 33620
rect 8777 33580 8812 33620
rect 8852 33580 8908 33620
rect 2476 33571 2516 33580
rect 3052 33536 3092 33580
rect 2659 33496 2668 33536
rect 2708 33496 2996 33536
rect 3043 33496 3052 33536
rect 3092 33496 3123 33536
rect 2956 33452 2996 33496
rect 3244 33452 3284 33580
rect 3820 33571 3860 33580
rect 5644 33536 5684 33580
rect 7276 33571 7316 33580
rect 8908 33571 8948 33580
rect 9004 33536 9044 34252
rect 9091 34168 9100 34208
rect 9140 34168 9149 34208
rect 9100 33620 9140 34168
rect 15820 33872 15860 34411
rect 16780 34376 16820 34420
rect 16876 34420 17155 34460
rect 17195 34420 17204 34460
rect 15907 34336 15916 34376
rect 15956 34336 16396 34376
rect 16436 34336 16445 34376
rect 16771 34336 16780 34376
rect 16820 34336 16829 34376
rect 16042 34168 16051 34208
rect 16091 34168 16820 34208
rect 15619 33832 15628 33872
rect 15668 33832 15860 33872
rect 16780 33788 16820 34168
rect 16876 33872 16916 34420
rect 17260 34376 17300 34504
rect 17635 34420 17644 34460
rect 17684 34420 17932 34460
rect 17972 34420 17981 34460
rect 18892 34451 20044 34460
rect 18932 34420 20044 34451
rect 20084 34420 20093 34460
rect 18892 34402 18932 34411
rect 17011 34336 17020 34376
rect 17060 34336 17068 34376
rect 17108 34336 17191 34376
rect 17260 34336 18836 34376
rect 18979 34336 18988 34376
rect 19028 34336 19372 34376
rect 19412 34336 19421 34376
rect 19625 34336 19660 34376
rect 19700 34336 19756 34376
rect 19796 34336 19805 34376
rect 20009 34336 20140 34376
rect 20180 34336 20189 34376
rect 18796 34292 18836 34336
rect 18796 34252 21292 34292
rect 21332 34252 21341 34292
rect 21510 34208 21600 34228
rect 17417 34168 17452 34208
rect 17492 34168 17548 34208
rect 17588 34168 17597 34208
rect 18307 34168 18316 34208
rect 18356 34168 19180 34208
rect 19220 34168 19229 34208
rect 21091 34168 21100 34208
rect 21140 34168 21600 34208
rect 21510 34148 21600 34168
rect 19843 34084 19852 34124
rect 19892 34084 20140 34124
rect 20180 34084 20189 34124
rect 18799 34000 18808 34040
rect 18848 34000 18890 34040
rect 18930 34000 18972 34040
rect 19012 34000 19054 34040
rect 19094 34000 19136 34040
rect 19176 34000 19185 34040
rect 16867 33832 16876 33872
rect 16916 33832 16925 33872
rect 10435 33748 10444 33788
rect 10484 33748 10493 33788
rect 11155 33748 11164 33788
rect 11204 33748 14092 33788
rect 14132 33748 14141 33788
rect 16780 33748 20620 33788
rect 20660 33748 20669 33788
rect 10444 33704 10484 33748
rect 21510 33704 21600 33724
rect 9859 33664 9868 33704
rect 9908 33664 10060 33704
rect 10100 33664 10109 33704
rect 10444 33664 10828 33704
rect 10868 33664 10877 33704
rect 15305 33664 15436 33704
rect 15476 33664 18356 33704
rect 10444 33620 10484 33664
rect 13804 33620 13844 33629
rect 15436 33620 15476 33664
rect 18316 33620 18356 33664
rect 21388 33664 21600 33704
rect 19948 33620 19988 33629
rect 9100 33580 9379 33620
rect 9419 33580 9428 33620
rect 9475 33580 9484 33620
rect 9524 33580 9580 33620
rect 9620 33580 9908 33620
rect 9955 33580 9964 33620
rect 10004 33580 10252 33620
rect 10292 33580 10301 33620
rect 10810 33580 10924 33620
rect 10972 33580 10990 33620
rect 12547 33580 12556 33620
rect 12596 33580 12605 33620
rect 13673 33580 13804 33620
rect 13844 33580 13853 33620
rect 14179 33580 14188 33620
rect 14228 33580 14237 33620
rect 16169 33580 16204 33620
rect 16244 33580 16300 33620
rect 16340 33580 16349 33620
rect 16457 33580 16483 33620
rect 16523 33580 16588 33620
rect 16628 33580 16637 33620
rect 16771 33580 16780 33620
rect 16820 33580 17068 33620
rect 17108 33580 17117 33620
rect 18356 33580 18508 33620
rect 18548 33580 18557 33620
rect 18691 33580 18700 33620
rect 18740 33580 18796 33620
rect 18836 33580 18871 33620
rect 9868 33536 9908 33580
rect 10444 33571 10484 33580
rect 3331 33496 3340 33536
rect 3380 33496 3518 33536
rect 3558 33496 3567 33536
rect 5644 33496 7220 33536
rect 9004 33496 9100 33536
rect 9140 33496 9149 33536
rect 9859 33496 9868 33536
rect 9908 33496 9917 33536
rect 7180 33452 7220 33496
rect 12556 33452 12596 33580
rect 13804 33571 13844 33580
rect 14188 33536 14228 33580
rect 15436 33571 15476 33580
rect 18316 33571 18356 33580
rect 18508 33536 18548 33580
rect 19948 33536 19988 33580
rect 13900 33496 14228 33536
rect 15715 33496 15724 33536
rect 15764 33496 16588 33536
rect 16628 33496 17452 33536
rect 17492 33496 17501 33536
rect 18508 33496 19988 33536
rect 21388 33536 21428 33664
rect 21510 33644 21600 33664
rect 21388 33496 21575 33536
rect 13900 33452 13940 33496
rect 2851 33412 2860 33452
rect 2900 33412 2909 33452
rect 2956 33412 3284 33452
rect 3610 33412 3619 33452
rect 3659 33412 3668 33452
rect 3715 33412 3724 33452
rect 3764 33412 3895 33452
rect 4243 33412 4252 33452
rect 4292 33412 7124 33452
rect 7180 33412 8908 33452
rect 8948 33412 8957 33452
rect 9571 33412 9580 33452
rect 9620 33412 11116 33452
rect 11156 33412 11165 33452
rect 12556 33412 13940 33452
rect 13987 33412 13996 33452
rect 14036 33412 15244 33452
rect 15284 33412 15293 33452
rect 18377 33412 18508 33452
rect 18548 33412 18557 33452
rect 19555 33412 19564 33452
rect 19604 33412 19613 33452
rect 19939 33412 19948 33452
rect 19988 33412 20140 33452
rect 20180 33412 20189 33452
rect 0 33368 90 33388
rect 2860 33368 2900 33412
rect 3628 33368 3668 33412
rect 0 33328 268 33368
rect 308 33328 317 33368
rect 2860 33328 2956 33368
rect 2996 33328 3005 33368
rect 3139 33328 3148 33368
rect 3188 33328 3668 33368
rect 7084 33368 7124 33412
rect 7084 33328 11692 33368
rect 11732 33328 11741 33368
rect 0 33308 90 33328
rect 12556 33284 12596 33412
rect 1123 33244 1132 33284
rect 1172 33244 4868 33284
rect 4919 33244 4928 33284
rect 4968 33244 5010 33284
rect 5050 33244 5092 33284
rect 5132 33244 5174 33284
rect 5214 33244 5256 33284
rect 5296 33244 5305 33284
rect 5923 33244 5932 33284
rect 5972 33244 8756 33284
rect 8995 33244 9004 33284
rect 9044 33244 12596 33284
rect 1411 33160 1420 33200
rect 1460 33160 1708 33200
rect 1748 33160 1757 33200
rect 4828 33116 4868 33244
rect 8716 33200 8756 33244
rect 19564 33200 19604 33412
rect 21535 33368 21575 33496
rect 19843 33328 19852 33368
rect 19892 33328 21575 33368
rect 20039 33244 20048 33284
rect 20088 33244 20130 33284
rect 20170 33244 20212 33284
rect 20252 33244 20294 33284
rect 20334 33244 20376 33284
rect 20416 33244 20425 33284
rect 21510 33200 21600 33220
rect 6892 33160 8236 33200
rect 8276 33160 8285 33200
rect 8419 33160 8428 33200
rect 8468 33160 8620 33200
rect 8660 33160 8669 33200
rect 8716 33160 11980 33200
rect 12020 33160 12029 33200
rect 19564 33160 19756 33200
rect 19796 33160 19805 33200
rect 20611 33160 20620 33200
rect 20660 33160 21600 33200
rect 6892 33116 6932 33160
rect 21510 33140 21600 33160
rect 3043 33076 3052 33116
rect 3092 33076 3436 33116
rect 3476 33076 3485 33116
rect 4387 33076 4396 33116
rect 4436 33076 4684 33116
rect 4724 33076 4733 33116
rect 4828 33076 6932 33116
rect 7817 33076 7948 33116
rect 7988 33076 7997 33116
rect 10147 33076 10156 33116
rect 10196 33076 10924 33116
rect 10964 33076 10973 33116
rect 13324 33076 13804 33116
rect 13844 33076 13853 33116
rect 15427 33076 15436 33116
rect 15476 33076 15485 33116
rect 16291 33076 16300 33116
rect 16340 33076 17164 33116
rect 17204 33076 17213 33116
rect 20131 33076 20140 33116
rect 20180 33076 20189 33116
rect 0 33032 90 33052
rect 0 32992 76 33032
rect 116 32992 125 33032
rect 1612 32992 4300 33032
rect 4340 32992 4349 33032
rect 0 32972 90 32992
rect 1612 32948 1652 32992
rect 931 32908 940 32948
rect 980 32908 1612 32948
rect 1652 32908 1661 32948
rect 1891 32908 1900 32948
rect 1940 32908 2092 32948
rect 2132 32908 2141 32948
rect 2467 32908 2476 32948
rect 2516 32939 2900 32948
rect 2516 32908 2860 32939
rect 3235 32908 3244 32948
rect 3284 32908 3293 32948
rect 3811 32908 3820 32948
rect 3860 32908 4492 32948
rect 4532 32908 4541 32948
rect 4963 32908 4972 32948
rect 5012 32908 5021 32948
rect 5129 32908 5164 32948
rect 5204 32908 5251 32948
rect 5291 32908 5309 32948
rect 5352 32908 5361 32948
rect 5401 32908 5410 32948
rect 5539 32908 5548 32948
rect 5588 32908 5740 32948
rect 5780 32908 5789 32948
rect 6185 32908 6316 32948
rect 6356 32908 6365 32948
rect 6665 32908 6796 32948
rect 6836 32908 6845 32948
rect 2860 32890 2900 32899
rect 3244 32864 3284 32908
rect 4492 32890 4532 32899
rect 163 32824 172 32864
rect 212 32824 1228 32864
rect 1268 32824 1277 32864
rect 3244 32824 3764 32864
rect 1891 32740 1900 32780
rect 1940 32740 3628 32780
rect 3668 32740 3677 32780
rect 0 32696 90 32716
rect 0 32656 76 32696
rect 116 32656 125 32696
rect 1459 32656 1468 32696
rect 1508 32656 1708 32696
rect 1748 32656 1757 32696
rect 0 32636 90 32656
rect 3724 32612 3764 32824
rect 4972 32780 5012 32908
rect 5361 32864 5401 32908
rect 6316 32890 6356 32899
rect 6796 32890 6836 32899
rect 6892 32864 6932 33076
rect 7747 32992 7756 33032
rect 7796 32992 8180 33032
rect 8140 32948 8180 32992
rect 13324 32948 13364 33076
rect 15436 33032 15476 33076
rect 20140 33032 20180 33076
rect 13411 32992 13420 33032
rect 13460 32992 13748 33032
rect 15436 32992 17108 33032
rect 13708 32948 13748 32992
rect 7459 32908 7468 32948
rect 7508 32908 7660 32948
rect 7700 32908 7709 32948
rect 7793 32908 7802 32948
rect 7842 32908 7948 32948
rect 7988 32908 7997 32948
rect 8131 32908 8140 32948
rect 8180 32908 8189 32948
rect 8246 32908 8255 32948
rect 8295 32908 8304 32948
rect 8419 32908 8428 32948
rect 8468 32908 8599 32948
rect 8707 32908 8716 32948
rect 8756 32908 9388 32948
rect 9428 32908 9437 32948
rect 9964 32939 10004 32948
rect 7660 32864 7700 32908
rect 8253 32864 8293 32908
rect 9964 32864 10004 32899
rect 10540 32939 11212 32948
rect 10580 32908 11212 32939
rect 11252 32908 11261 32948
rect 11683 32908 11692 32948
rect 11732 32908 11788 32948
rect 11828 32908 11863 32948
rect 11971 32908 11980 32948
rect 12020 32908 12151 32948
rect 13228 32939 13364 32948
rect 10540 32890 10580 32899
rect 13268 32908 13364 32939
rect 13690 32908 13699 32948
rect 13739 32908 13748 32948
rect 13795 32908 13804 32948
rect 13844 32908 13975 32948
rect 14179 32908 14188 32948
rect 14228 32908 14237 32948
rect 14764 32939 14900 32948
rect 13228 32890 13268 32899
rect 14188 32864 14228 32908
rect 14804 32908 14900 32939
rect 15113 32908 15244 32948
rect 15284 32908 15293 32948
rect 15715 32908 15724 32948
rect 15764 32908 16588 32948
rect 16628 32908 16780 32948
rect 16820 32908 16829 32948
rect 16972 32939 17012 32948
rect 14764 32890 14804 32899
rect 5251 32824 5260 32864
rect 5300 32824 5401 32864
rect 5705 32824 5836 32864
rect 5876 32824 5885 32864
rect 6883 32824 6892 32864
rect 6932 32824 7276 32864
rect 7316 32824 7325 32864
rect 7660 32824 8293 32864
rect 8803 32824 8812 32864
rect 8852 32824 9580 32864
rect 9620 32824 10004 32864
rect 13699 32824 13708 32864
rect 13748 32824 14228 32864
rect 14275 32824 14284 32864
rect 14324 32824 14455 32864
rect 4291 32740 4300 32780
rect 4340 32740 5012 32780
rect 8009 32740 8044 32780
rect 8084 32740 8140 32780
rect 8180 32740 8189 32780
rect 14860 32696 14900 32908
rect 15244 32890 15284 32899
rect 16972 32864 17012 32899
rect 15811 32824 15820 32864
rect 15860 32824 17012 32864
rect 17068 32864 17108 32992
rect 18412 32992 18508 33032
rect 18548 32992 18557 33032
rect 20140 32992 21388 33032
rect 21428 32992 21437 33032
rect 18412 32948 18452 32992
rect 18394 32908 18403 32948
rect 18443 32908 18452 32948
rect 18499 32908 18508 32948
rect 18548 32908 18557 32948
rect 18604 32908 18892 32948
rect 18932 32908 18941 32948
rect 19468 32939 19508 32948
rect 18508 32864 18548 32908
rect 17068 32824 17548 32864
rect 17588 32824 17597 32864
rect 17801 32824 17932 32864
rect 17972 32824 17981 32864
rect 18461 32824 18508 32864
rect 18548 32824 18557 32864
rect 18604 32780 18644 32908
rect 19817 32908 19948 32948
rect 19988 32908 19997 32948
rect 18691 32824 18700 32864
rect 18740 32824 18988 32864
rect 19028 32824 19037 32864
rect 18076 32740 18644 32780
rect 19468 32780 19508 32899
rect 19948 32890 19988 32899
rect 19468 32740 19948 32780
rect 19988 32740 19997 32780
rect 4579 32656 4588 32696
rect 4628 32656 4828 32696
rect 4868 32656 4877 32696
rect 6953 32656 7027 32696
rect 7067 32656 7084 32696
rect 7124 32656 7133 32696
rect 7459 32656 7468 32696
rect 7508 32656 7516 32696
rect 7556 32656 7639 32696
rect 7939 32656 7948 32696
rect 7988 32656 8332 32696
rect 8372 32656 9676 32696
rect 9716 32656 9725 32696
rect 10339 32656 10348 32696
rect 10388 32656 10519 32696
rect 14755 32656 14764 32696
rect 14804 32656 14900 32696
rect 17299 32656 17308 32696
rect 17348 32656 17356 32696
rect 17396 32656 17479 32696
rect 17548 32656 17692 32696
rect 17732 32656 17741 32696
rect 17548 32612 17588 32656
rect 3724 32572 8812 32612
rect 8852 32572 8861 32612
rect 16771 32572 16780 32612
rect 16820 32572 17164 32612
rect 17204 32572 17588 32612
rect 3679 32488 3688 32528
rect 3728 32488 3770 32528
rect 3810 32488 3852 32528
rect 3892 32488 3934 32528
rect 3974 32488 4016 32528
rect 4056 32488 4065 32528
rect 6988 32404 7084 32444
rect 7124 32404 7133 32444
rect 0 32360 90 32380
rect 0 32320 3532 32360
rect 3572 32320 3581 32360
rect 4771 32320 4780 32360
rect 4820 32320 5164 32360
rect 5204 32320 5213 32360
rect 6403 32320 6412 32360
rect 6452 32320 6796 32360
rect 6836 32320 6845 32360
rect 0 32300 90 32320
rect 2179 32236 2188 32276
rect 2228 32236 2668 32276
rect 2708 32236 2717 32276
rect 6988 32192 7028 32404
rect 7756 32360 7796 32572
rect 7939 32488 7948 32528
rect 7988 32488 10540 32528
rect 10580 32488 11404 32528
rect 11444 32488 11453 32528
rect 8035 32404 8044 32444
rect 8084 32404 8756 32444
rect 9091 32404 9100 32444
rect 9140 32404 12556 32444
rect 12596 32404 12605 32444
rect 14371 32404 14380 32444
rect 14420 32404 17452 32444
rect 17492 32404 17501 32444
rect 7363 32320 7372 32360
rect 7412 32320 7660 32360
rect 7700 32320 7709 32360
rect 7756 32320 7900 32360
rect 7940 32320 7949 32360
rect 7075 32236 7084 32276
rect 7124 32236 7412 32276
rect 7372 32192 7412 32236
rect 8716 32192 8756 32404
rect 8803 32320 8812 32360
rect 8852 32320 11692 32360
rect 11732 32320 11741 32360
rect 12019 32320 12028 32360
rect 12068 32320 12460 32360
rect 12500 32320 12509 32360
rect 16675 32320 16684 32360
rect 16724 32320 17068 32360
rect 17108 32320 17117 32360
rect 18076 32276 18116 32740
rect 21510 32696 21600 32716
rect 18787 32656 18796 32696
rect 18836 32656 19468 32696
rect 19508 32656 19517 32696
rect 20611 32656 20620 32696
rect 20660 32656 21600 32696
rect 21510 32636 21600 32656
rect 18799 32488 18808 32528
rect 18848 32488 18890 32528
rect 18930 32488 18972 32528
rect 19012 32488 19054 32528
rect 19094 32488 19136 32528
rect 19176 32488 19185 32528
rect 18172 32404 20428 32444
rect 20468 32404 20477 32444
rect 18172 32360 18212 32404
rect 18163 32320 18172 32360
rect 18212 32320 18221 32360
rect 9475 32236 9484 32276
rect 9524 32236 13708 32276
rect 13748 32236 14228 32276
rect 14851 32236 14860 32276
rect 14900 32236 18932 32276
rect 14188 32192 14228 32236
rect 18892 32192 18932 32236
rect 19468 32236 19948 32276
rect 19988 32236 19997 32276
rect 3082 32183 3148 32192
rect 3082 32143 3091 32183
rect 3131 32152 3148 32183
rect 3188 32152 3271 32192
rect 6403 32152 6412 32192
rect 6452 32152 6604 32192
rect 6644 32152 6653 32192
rect 6979 32152 6988 32192
rect 7028 32152 7037 32192
rect 7363 32152 7372 32192
rect 7412 32152 7421 32192
rect 7555 32152 7564 32192
rect 7604 32152 8140 32192
rect 8180 32152 8189 32192
rect 8323 32152 8332 32192
rect 8372 32152 8381 32192
rect 8707 32152 8716 32192
rect 8756 32152 8765 32192
rect 8899 32152 8908 32192
rect 8948 32152 8956 32192
rect 8996 32152 9079 32192
rect 9187 32152 9196 32192
rect 9236 32152 9388 32192
rect 9428 32152 9437 32192
rect 9763 32152 9772 32192
rect 9812 32152 9908 32192
rect 10051 32152 10060 32192
rect 10100 32152 10252 32192
rect 10292 32152 10301 32192
rect 11753 32152 11788 32192
rect 11828 32152 11884 32192
rect 11924 32152 11933 32192
rect 12067 32152 12076 32192
rect 12116 32152 12364 32192
rect 12404 32152 12413 32192
rect 14179 32152 14188 32192
rect 14228 32152 14237 32192
rect 17129 32152 17260 32192
rect 17300 32152 17309 32192
rect 17801 32152 17932 32192
rect 17972 32152 17981 32192
rect 18220 32152 18508 32192
rect 18548 32152 18557 32192
rect 18883 32152 18892 32192
rect 18932 32152 18941 32192
rect 3131 32143 3140 32152
rect 3082 32142 3140 32143
rect 2476 32108 2516 32117
rect 4588 32108 4628 32117
rect 6220 32108 6260 32117
rect 8332 32108 8372 32152
rect 9868 32108 9908 32152
rect 10828 32108 10868 32117
rect 14764 32108 14804 32117
rect 16876 32108 16916 32117
rect 18220 32108 18260 32152
rect 18508 32108 18548 32152
rect 19468 32108 19508 32236
rect 21510 32192 21600 32212
rect 19555 32152 19564 32192
rect 19604 32152 21600 32192
rect 21510 32132 21600 32152
rect 1027 32068 1036 32108
rect 1076 32068 1228 32108
rect 1268 32068 1277 32108
rect 2345 32068 2476 32108
rect 2516 32068 2525 32108
rect 2851 32068 2860 32108
rect 2900 32068 2955 32108
rect 2995 32068 3031 32108
rect 3184 32068 3193 32108
rect 3233 32068 3284 32108
rect 3331 32068 3340 32108
rect 3380 32068 3389 32108
rect 4628 32068 4780 32108
rect 4820 32068 4829 32108
rect 4963 32068 4972 32108
rect 5012 32068 5452 32108
rect 5492 32068 5501 32108
rect 7267 32068 7276 32108
rect 7316 32068 8372 32108
rect 9754 32068 9763 32108
rect 9803 32068 9812 32108
rect 9859 32068 9868 32108
rect 9908 32068 9917 32108
rect 10313 32068 10348 32108
rect 10388 32068 10444 32108
rect 10484 32068 10493 32108
rect 10697 32068 10828 32108
rect 10868 32068 10877 32108
rect 11338 32068 11347 32108
rect 11387 32068 11500 32108
rect 11540 32068 11549 32108
rect 13507 32068 13516 32108
rect 13556 32068 13699 32108
rect 13739 32068 13748 32108
rect 13795 32068 13804 32108
rect 13844 32068 13975 32108
rect 14179 32068 14188 32108
rect 14228 32068 14284 32108
rect 14324 32068 14359 32108
rect 14633 32068 14764 32108
rect 14804 32068 14813 32108
rect 15235 32068 15244 32108
rect 15292 32068 15415 32108
rect 15619 32068 15628 32108
rect 15668 32068 16300 32108
rect 16340 32068 16349 32108
rect 17443 32068 17452 32108
rect 17492 32068 18260 32108
rect 18394 32068 18403 32108
rect 18443 32068 18452 32108
rect 18499 32068 18508 32108
rect 18548 32068 18557 32108
rect 18691 32068 18700 32108
rect 18740 32068 18988 32108
rect 19028 32068 19037 32108
rect 19084 32068 19468 32108
rect 19947 32068 19956 32108
rect 19996 32068 20005 32108
rect 2476 32059 2516 32068
rect 0 32024 90 32044
rect 3244 32024 3284 32068
rect 0 31984 1228 32024
rect 1268 31984 1277 32024
rect 3043 31984 3052 32024
rect 3092 31984 3284 32024
rect 3340 32024 3380 32068
rect 4588 32059 4628 32068
rect 4780 32024 4820 32068
rect 6220 32024 6260 32068
rect 9772 32024 9812 32068
rect 10828 32059 10868 32068
rect 14188 32024 14228 32068
rect 14764 32059 14804 32068
rect 16876 32024 16916 32068
rect 18412 32024 18452 32068
rect 3340 31984 3476 32024
rect 4780 31984 6260 32024
rect 8247 31984 9668 32024
rect 9772 31984 9964 32024
rect 10004 31984 10013 32024
rect 10924 31984 12980 32024
rect 13699 31984 13708 32024
rect 13748 31984 14228 32024
rect 15244 31984 15820 32024
rect 15860 31984 16916 32024
rect 17827 31984 17836 32024
rect 17876 31984 17885 32024
rect 18412 31984 18508 32024
rect 18548 31984 18557 32024
rect 0 31964 90 31984
rect 2851 31900 2860 31940
rect 2900 31900 3340 31940
rect 3380 31900 3389 31940
rect 3436 31856 3476 31984
rect 6835 31900 6844 31940
rect 6884 31900 6988 31940
rect 7028 31900 7037 31940
rect 7219 31900 7228 31940
rect 7268 31900 7508 31940
rect 7603 31900 7612 31940
rect 7652 31900 7660 31940
rect 7700 31900 7783 31940
rect 6988 31856 7028 31900
rect 7468 31856 7508 31900
rect 3436 31816 6892 31856
rect 6932 31816 6941 31856
rect 6988 31816 7372 31856
rect 7412 31816 7421 31856
rect 7468 31816 8140 31856
rect 8180 31816 8189 31856
rect 8247 31772 8287 31984
rect 9628 31940 9668 31984
rect 10924 31940 10964 31984
rect 12940 31940 12980 31984
rect 15244 31940 15284 31984
rect 17836 31940 17876 31984
rect 8563 31900 8572 31940
rect 8612 31900 9332 31940
rect 9379 31900 9388 31940
rect 9428 31900 9436 31940
rect 9476 31900 9559 31940
rect 9628 31900 10964 31940
rect 11491 31900 11500 31940
rect 11540 31900 11549 31940
rect 12115 31900 12124 31940
rect 12164 31900 12556 31940
rect 12596 31900 12605 31940
rect 12940 31900 15284 31940
rect 15401 31900 15436 31940
rect 15476 31900 15532 31940
rect 15572 31900 15581 31940
rect 17491 31900 17500 31940
rect 17540 31900 17644 31940
rect 17684 31900 17876 31940
rect 9292 31856 9332 31900
rect 11500 31856 11540 31900
rect 18700 31856 18740 32068
rect 19084 32024 19124 32068
rect 19468 32059 19508 32068
rect 19075 31984 19084 32024
rect 19124 31984 19133 32024
rect 9292 31816 10484 31856
rect 11500 31816 12268 31856
rect 12308 31816 12460 31856
rect 12500 31816 12509 31856
rect 13699 31816 13708 31856
rect 13748 31816 18740 31856
rect 10444 31772 10484 31816
rect 3139 31732 3148 31772
rect 3188 31732 4204 31772
rect 4244 31732 4253 31772
rect 4919 31732 4928 31772
rect 4968 31732 5010 31772
rect 5050 31732 5092 31772
rect 5132 31732 5174 31772
rect 5214 31732 5256 31772
rect 5296 31732 5305 31772
rect 5539 31732 5548 31772
rect 5588 31732 8287 31772
rect 10435 31732 10444 31772
rect 10484 31732 11308 31772
rect 11348 31732 11357 31772
rect 16291 31732 16300 31772
rect 16340 31732 19468 31772
rect 19508 31732 19517 31772
rect 0 31688 90 31708
rect 19948 31688 19988 32068
rect 20131 31900 20140 31940
rect 20180 31900 21196 31940
rect 21236 31900 21245 31940
rect 20039 31732 20048 31772
rect 20088 31732 20130 31772
rect 20170 31732 20212 31772
rect 20252 31732 20294 31772
rect 20334 31732 20376 31772
rect 20416 31732 20425 31772
rect 21510 31688 21600 31708
rect 0 31648 172 31688
rect 212 31648 221 31688
rect 2668 31648 4492 31688
rect 4532 31648 4541 31688
rect 5644 31648 5876 31688
rect 19948 31648 20276 31688
rect 0 31628 90 31648
rect 1289 31396 1420 31436
rect 1460 31396 1469 31436
rect 2668 31427 2708 31648
rect 5644 31604 5684 31648
rect 4291 31564 4300 31604
rect 4340 31564 5684 31604
rect 5836 31604 5876 31648
rect 20236 31604 20276 31648
rect 20812 31648 21600 31688
rect 5836 31564 6111 31604
rect 6394 31564 6403 31604
rect 6452 31564 6583 31604
rect 9833 31564 9964 31604
rect 10004 31564 10013 31604
rect 11491 31564 11500 31604
rect 11540 31564 11596 31604
rect 11636 31564 11671 31604
rect 12940 31564 16340 31604
rect 18377 31564 18508 31604
rect 18548 31564 18557 31604
rect 20227 31564 20236 31604
rect 20276 31564 20285 31604
rect 3043 31480 3052 31520
rect 3092 31480 3223 31520
rect 4962 31480 4971 31520
rect 5011 31480 5260 31520
rect 5300 31480 5309 31520
rect 5361 31436 5401 31564
rect 5827 31480 5836 31520
rect 5876 31480 6007 31520
rect 6071 31436 6111 31564
rect 12940 31520 12980 31564
rect 8707 31480 8716 31520
rect 8756 31480 10196 31520
rect 10531 31480 10540 31520
rect 10580 31480 12980 31520
rect 13411 31480 13420 31520
rect 13460 31480 13940 31520
rect 2668 31378 2708 31387
rect 3052 31427 3284 31436
rect 3052 31396 3244 31427
rect 0 31352 90 31372
rect 3052 31352 3092 31396
rect 4195 31396 4204 31436
rect 4244 31396 4492 31436
rect 4532 31396 4541 31436
rect 5033 31396 5101 31436
rect 5141 31396 5164 31436
rect 5204 31396 5213 31436
rect 5347 31396 5356 31436
rect 5396 31396 5405 31436
rect 5624 31403 5633 31436
rect 5547 31396 5633 31403
rect 5673 31396 5684 31436
rect 3244 31378 3284 31387
rect 5547 31363 5684 31396
rect 5921 31363 5930 31403
rect 5970 31363 5979 31403
rect 6062 31396 6071 31436
rect 6111 31396 6120 31436
rect 6307 31396 6316 31436
rect 6356 31396 6495 31436
rect 6665 31396 6796 31436
rect 6836 31396 6845 31436
rect 7267 31396 7276 31436
rect 7316 31427 8084 31436
rect 7316 31396 8044 31427
rect 0 31312 652 31352
rect 692 31312 701 31352
rect 3043 31312 3052 31352
rect 3092 31312 3101 31352
rect 0 31292 90 31312
rect 5547 31268 5587 31363
rect 4588 31228 5587 31268
rect 4588 31184 4628 31228
rect 2851 31144 2860 31184
rect 2900 31144 3031 31184
rect 3523 31144 3532 31184
rect 3572 31144 4628 31184
rect 4675 31144 4684 31184
rect 4724 31144 4733 31184
rect 5626 31144 5635 31184
rect 5675 31144 5740 31184
rect 5780 31144 5815 31184
rect 0 31016 90 31036
rect 0 30976 2188 31016
rect 2228 30976 2237 31016
rect 3679 30976 3688 31016
rect 3728 30976 3770 31016
rect 3810 30976 3852 31016
rect 3892 30976 3934 31016
rect 3974 30976 4016 31016
rect 4056 30976 4065 31016
rect 0 30956 90 30976
rect 2537 30808 2668 30848
rect 2708 30808 2717 30848
rect 4361 30808 4483 30848
rect 4532 30808 4541 30848
rect 3331 30724 3340 30764
rect 3380 30724 4300 30764
rect 4340 30724 4349 30764
rect 0 30680 90 30700
rect 4684 30680 4724 31144
rect 5932 31100 5972 31363
rect 6202 31312 6211 31352
rect 6260 31312 6391 31352
rect 4867 31060 4876 31100
rect 4916 31060 5972 31100
rect 6455 30932 6495 31396
rect 8515 31396 8524 31436
rect 8564 31396 8948 31436
rect 8044 31378 8084 31387
rect 8908 31184 8948 31396
rect 9484 31268 9524 31480
rect 10156 31436 10196 31480
rect 13900 31436 13940 31480
rect 14361 31480 14572 31520
rect 14612 31480 14860 31520
rect 14900 31480 14909 31520
rect 15235 31480 15244 31520
rect 15284 31480 15436 31520
rect 15476 31480 15485 31520
rect 15532 31480 16108 31520
rect 16148 31480 16157 31520
rect 9612 31396 9676 31436
rect 9716 31427 9964 31436
rect 9716 31396 9772 31427
rect 9812 31396 9964 31427
rect 10004 31396 10100 31436
rect 10147 31396 10156 31436
rect 10196 31396 10205 31436
rect 11404 31427 11444 31436
rect 9772 31378 9812 31387
rect 10060 31352 10100 31396
rect 11945 31396 11980 31436
rect 12020 31396 12076 31436
rect 12116 31396 12125 31436
rect 12739 31396 12748 31436
rect 12788 31427 13268 31436
rect 12788 31396 13228 31427
rect 11404 31352 11444 31387
rect 13769 31396 13900 31436
rect 13940 31396 14188 31436
rect 14228 31396 14237 31436
rect 13228 31378 13268 31387
rect 14361 31352 14401 31480
rect 14458 31396 14467 31436
rect 14507 31396 14516 31436
rect 14907 31396 14956 31436
rect 14996 31396 15038 31436
rect 15078 31396 15087 31436
rect 15340 31427 15380 31436
rect 10060 31312 11444 31352
rect 13429 31312 14401 31352
rect 9484 31228 13132 31268
rect 13172 31228 13181 31268
rect 8105 31144 8236 31184
rect 8276 31144 8285 31184
rect 8908 31144 10252 31184
rect 10292 31144 12076 31184
rect 12116 31144 12125 31184
rect 6787 31060 6796 31100
rect 6836 31060 12268 31100
rect 12308 31060 12317 31100
rect 5059 30892 5068 30932
rect 5108 30892 6495 30932
rect 9484 30892 13132 30932
rect 13172 30892 13181 30932
rect 5260 30808 5740 30848
rect 5780 30808 9100 30848
rect 9140 30808 9149 30848
rect 0 30640 748 30680
rect 788 30640 797 30680
rect 2476 30640 3052 30680
rect 3092 30640 3101 30680
rect 4684 30640 4820 30680
rect 0 30620 90 30640
rect 2476 30596 2516 30640
rect 4108 30596 4148 30605
rect 4780 30596 4820 30640
rect 5260 30596 5300 30808
rect 9484 30764 9524 30892
rect 13429 30848 13469 31312
rect 14476 31268 14516 31396
rect 15340 31352 15380 31387
rect 15532 31352 15572 31480
rect 15916 31396 16204 31436
rect 16244 31396 16253 31436
rect 15916 31352 15956 31396
rect 16300 31352 16340 31564
rect 20812 31520 20852 31648
rect 21510 31628 21600 31648
rect 16531 31480 16540 31520
rect 16580 31480 20852 31520
rect 17059 31396 17068 31436
rect 17108 31396 17117 31436
rect 17443 31396 17452 31436
rect 17492 31396 18220 31436
rect 18260 31427 18391 31436
rect 18260 31396 18316 31427
rect 14563 31312 14572 31352
rect 14612 31312 15380 31352
rect 15523 31312 15532 31352
rect 15572 31312 15581 31352
rect 15907 31312 15916 31352
rect 15956 31312 15965 31352
rect 16291 31312 16300 31352
rect 16340 31312 16349 31352
rect 16579 31312 16588 31352
rect 16628 31312 16704 31352
rect 16841 31312 16876 31352
rect 16916 31312 16972 31352
rect 17012 31312 17021 31352
rect 16588 31268 16628 31312
rect 17068 31268 17108 31396
rect 18356 31396 18391 31427
rect 18787 31396 18796 31436
rect 18836 31396 19468 31436
rect 19508 31396 19517 31436
rect 19913 31396 20044 31436
rect 20084 31396 20093 31436
rect 18316 31378 18356 31387
rect 20044 31378 20084 31387
rect 14476 31228 14764 31268
rect 14804 31228 15820 31268
rect 15860 31228 15869 31268
rect 16099 31228 16108 31268
rect 16148 31228 17108 31268
rect 21510 31184 21600 31204
rect 13747 31144 13756 31184
rect 13796 31144 14188 31184
rect 14228 31144 14237 31184
rect 14729 31144 14860 31184
rect 14900 31144 14909 31184
rect 15034 31144 15043 31184
rect 15092 31144 15223 31184
rect 15763 31144 15772 31184
rect 15812 31144 15821 31184
rect 16147 31144 16156 31184
rect 16196 31144 16532 31184
rect 16579 31144 16588 31184
rect 16628 31144 16636 31184
rect 16676 31144 16759 31184
rect 18892 31144 21600 31184
rect 15772 30932 15812 31144
rect 16492 31100 16532 31144
rect 18892 31100 18932 31144
rect 21510 31124 21600 31144
rect 16492 31060 18932 31100
rect 18799 30976 18808 31016
rect 18848 30976 18890 31016
rect 18930 30976 18972 31016
rect 19012 30976 19054 31016
rect 19094 30976 19136 31016
rect 19176 30976 19185 31016
rect 15772 30892 21236 30932
rect 10697 30808 10780 30848
rect 10820 30808 10828 30848
rect 10868 30808 10877 30848
rect 11155 30808 11164 30848
rect 11204 30808 13469 30848
rect 14563 30808 14572 30848
rect 14612 30808 14743 30848
rect 18835 30808 18844 30848
rect 18884 30808 19564 30848
rect 19604 30808 19613 30848
rect 19747 30808 19756 30848
rect 19796 30808 19996 30848
rect 20036 30808 20045 30848
rect 20371 30808 20380 30848
rect 20420 30808 20908 30848
rect 20948 30808 20957 30848
rect 6796 30724 9524 30764
rect 9571 30724 9580 30764
rect 9620 30724 12940 30764
rect 12980 30724 12989 30764
rect 16012 30724 18124 30764
rect 18164 30724 18173 30764
rect 19603 30724 19612 30764
rect 19652 30724 21100 30764
rect 21140 30724 21149 30764
rect 6508 30596 6548 30605
rect 6796 30596 6836 30724
rect 6883 30640 6892 30680
rect 6932 30640 7124 30680
rect 7433 30640 7468 30680
rect 7508 30640 7564 30680
rect 7604 30640 7613 30680
rect 7084 30596 7124 30640
rect 8044 30596 8084 30605
rect 9100 30596 9140 30605
rect 9484 30596 9524 30724
rect 10348 30640 10540 30680
rect 10580 30640 10636 30680
rect 10676 30640 10685 30680
rect 10915 30640 10924 30680
rect 10964 30640 11444 30680
rect 10348 30596 10388 30640
rect 10636 30596 10676 30640
rect 355 30556 364 30596
rect 404 30556 1228 30596
rect 1268 30556 1420 30596
rect 1460 30556 1469 30596
rect 2345 30556 2476 30596
rect 2516 30556 2525 30596
rect 2851 30556 2860 30596
rect 2900 30556 4052 30596
rect 2476 30547 2516 30556
rect 0 30344 90 30364
rect 0 30304 2668 30344
rect 2708 30304 2717 30344
rect 2764 30304 3916 30344
rect 3956 30304 3965 30344
rect 0 30284 90 30304
rect 2764 30092 2804 30304
rect 4012 30260 4052 30556
rect 4148 30556 4492 30596
rect 4532 30556 4541 30596
rect 4937 30556 5068 30596
rect 5108 30556 5117 30596
rect 5251 30556 5260 30596
rect 5300 30556 5309 30596
rect 6548 30556 6836 30596
rect 6970 30556 6979 30596
rect 7019 30556 7028 30596
rect 7075 30556 7084 30596
rect 7124 30556 7133 30596
rect 7459 30556 7468 30596
rect 7508 30556 7564 30596
rect 7604 30556 7639 30596
rect 8554 30556 8563 30596
rect 8603 30556 8948 30596
rect 4108 30547 4148 30556
rect 4780 30547 4820 30556
rect 6508 30547 6548 30556
rect 6988 30512 7028 30556
rect 8044 30512 8084 30556
rect 8908 30512 8948 30556
rect 9140 30556 9524 30596
rect 10339 30556 10348 30596
rect 10388 30556 10397 30596
rect 10636 30556 11308 30596
rect 11348 30556 11357 30596
rect 9100 30547 9140 30556
rect 4195 30472 4204 30512
rect 4244 30472 4478 30512
rect 4518 30472 4527 30512
rect 6691 30472 6700 30512
rect 6740 30472 7028 30512
rect 7363 30472 7372 30512
rect 7412 30472 8084 30512
rect 8899 30472 8908 30512
rect 8948 30472 8957 30512
rect 11404 30428 11444 30640
rect 12748 30640 13469 30680
rect 12556 30596 12596 30605
rect 12355 30556 12364 30596
rect 12404 30556 12556 30596
rect 12556 30547 12596 30556
rect 12748 30512 12788 30640
rect 13429 30596 13469 30640
rect 13546 30671 13940 30680
rect 13546 30631 13555 30671
rect 13595 30640 13940 30671
rect 13595 30631 13604 30640
rect 13546 30630 13604 30631
rect 13900 30596 13940 30640
rect 14188 30640 15916 30680
rect 15956 30640 15965 30680
rect 14188 30596 14228 30640
rect 16012 30596 16052 30724
rect 21196 30680 21236 30892
rect 21510 30680 21600 30700
rect 16963 30640 16972 30680
rect 17012 30640 17164 30680
rect 17204 30640 17213 30680
rect 17548 30640 18412 30680
rect 18452 30640 18461 30680
rect 18595 30640 18604 30680
rect 18644 30640 18653 30680
rect 18787 30640 18796 30680
rect 18836 30640 18988 30680
rect 19028 30640 19037 30680
rect 19241 30640 19372 30680
rect 19412 30640 19421 30680
rect 19625 30640 19756 30680
rect 19796 30640 19805 30680
rect 20009 30640 20140 30680
rect 20180 30640 20189 30680
rect 21196 30640 21600 30680
rect 17548 30596 17588 30640
rect 18604 30596 18644 30640
rect 21510 30620 21600 30640
rect 13027 30556 13036 30596
rect 13076 30556 13324 30596
rect 13364 30556 13373 30596
rect 13420 30556 13429 30596
rect 13469 30556 13478 30596
rect 13648 30556 13657 30596
rect 13697 30556 13708 30596
rect 13748 30556 13837 30596
rect 13891 30556 13900 30596
rect 13940 30556 14071 30596
rect 14170 30556 14179 30596
rect 14219 30556 14228 30596
rect 14371 30556 14380 30596
rect 14420 30556 14764 30596
rect 14804 30556 14813 30596
rect 14188 30512 14228 30556
rect 12739 30472 12748 30512
rect 12788 30472 12797 30512
rect 13049 30472 13132 30512
rect 13172 30472 13180 30512
rect 13220 30472 13229 30512
rect 13324 30472 14228 30512
rect 14275 30472 14284 30512
rect 14324 30472 14572 30512
rect 14612 30472 15724 30512
rect 15764 30472 15773 30512
rect 4675 30388 4684 30428
rect 4724 30388 4924 30428
rect 4964 30388 4973 30428
rect 8585 30388 8716 30428
rect 8756 30388 8765 30428
rect 8899 30388 8908 30428
rect 8948 30388 11444 30428
rect 12748 30428 12788 30472
rect 12748 30388 13076 30428
rect 4684 30344 4724 30388
rect 4291 30304 4300 30344
rect 4340 30304 4724 30344
rect 4780 30304 12844 30344
rect 12884 30304 12893 30344
rect 4780 30260 4820 30304
rect 4012 30220 4820 30260
rect 4919 30220 4928 30260
rect 4968 30220 5010 30260
rect 5050 30220 5092 30260
rect 5132 30220 5174 30260
rect 5214 30220 5256 30260
rect 5296 30220 5305 30260
rect 2851 30136 2860 30176
rect 2900 30136 12940 30176
rect 12980 30136 12989 30176
rect 1420 30052 2668 30092
rect 2708 30052 2717 30092
rect 2764 30052 2860 30092
rect 2900 30052 2964 30092
rect 3043 30052 3052 30092
rect 3092 30052 3148 30092
rect 3188 30052 4204 30092
rect 4244 30052 4253 30092
rect 4972 30052 6316 30092
rect 6356 30052 6365 30092
rect 8620 30052 10636 30092
rect 10676 30052 10685 30092
rect 0 30008 90 30028
rect 0 29968 844 30008
rect 884 29968 893 30008
rect 0 29948 90 29968
rect 1420 29924 1460 30052
rect 3244 29968 4876 30008
rect 4916 29968 4925 30008
rect 3244 29924 3284 29968
rect 4972 29924 5012 30052
rect 6403 29968 6412 30008
rect 6452 29968 6461 30008
rect 7660 29968 7756 30008
rect 7796 29968 7805 30008
rect 6412 29924 6452 29968
rect 1315 29884 1324 29924
rect 1364 29884 1420 29924
rect 1460 29884 1495 29924
rect 2668 29915 3284 29924
rect 2708 29884 3244 29915
rect 2668 29866 2708 29875
rect 4483 29884 4492 29924
rect 4532 29884 4541 29924
rect 4649 29884 4780 29924
rect 4820 29884 4829 29924
rect 4963 29884 4972 29924
rect 5012 29884 5021 29924
rect 6089 29884 6220 29924
rect 6260 29884 6269 29924
rect 6412 29884 6691 29924
rect 6731 29884 6740 29924
rect 6787 29884 6796 29924
rect 6836 29884 6892 29924
rect 6932 29884 6967 29924
rect 7171 29884 7180 29924
rect 7220 29884 7564 29924
rect 7604 29884 7613 29924
rect 3244 29866 3284 29875
rect 4492 29840 4532 29884
rect 6220 29866 6260 29875
rect 7660 29840 7700 29968
rect 7756 29915 7948 29924
rect 7796 29884 7948 29915
rect 7988 29884 7997 29924
rect 8105 29884 8236 29924
rect 8276 29884 8285 29924
rect 7756 29866 7796 29875
rect 8236 29866 8276 29875
rect 8620 29840 8660 30052
rect 13036 30008 13076 30388
rect 13324 30344 13364 30472
rect 13420 30388 14188 30428
rect 14228 30388 14237 30428
rect 13315 30304 13324 30344
rect 13364 30304 13373 30344
rect 13420 30008 13460 30388
rect 16012 30344 16052 30556
rect 16204 30556 16483 30596
rect 16523 30556 16532 30596
rect 16579 30556 16588 30596
rect 16628 30556 16637 30596
rect 16937 30556 17068 30596
rect 17108 30556 17117 30596
rect 17731 30556 17740 30596
rect 17780 30556 18036 30596
rect 18076 30556 18085 30596
rect 18604 30556 20908 30596
rect 20948 30556 20957 30596
rect 16204 30512 16244 30556
rect 16588 30512 16628 30556
rect 17548 30547 17588 30556
rect 16195 30472 16204 30512
rect 16244 30472 16253 30512
rect 16387 30472 16396 30512
rect 16436 30472 16628 30512
rect 19219 30472 19228 30512
rect 19268 30472 20428 30512
rect 20468 30472 20477 30512
rect 16963 30388 16972 30428
rect 17012 30388 18220 30428
rect 18260 30388 18269 30428
rect 13996 30304 14708 30344
rect 15715 30304 15724 30344
rect 15764 30304 16052 30344
rect 8851 29968 8860 30008
rect 8900 29968 9196 30008
rect 9236 29968 9245 30008
rect 9676 29968 10348 30008
rect 10388 29968 10397 30008
rect 10540 29968 12652 30008
rect 12692 29968 12701 30008
rect 12835 29968 12844 30008
rect 12884 29968 13076 30008
rect 9676 29924 9716 29968
rect 8899 29884 8908 29924
rect 8948 29884 9004 29924
rect 9044 29884 9079 29924
rect 9187 29884 9196 29924
rect 9236 29884 9245 29924
rect 9658 29884 9667 29924
rect 9707 29884 9716 29924
rect 9763 29884 9772 29924
rect 9812 29884 9821 29924
rect 10147 29884 10156 29924
rect 10196 29884 10444 29924
rect 10484 29884 10493 29924
rect 9196 29840 9236 29884
rect 9772 29840 9812 29884
rect 4492 29800 5740 29840
rect 5780 29800 5789 29840
rect 7267 29800 7276 29840
rect 7316 29800 7700 29840
rect 8611 29800 8620 29840
rect 8660 29800 8669 29840
rect 8812 29800 9236 29840
rect 9571 29800 9580 29840
rect 9620 29800 10060 29840
rect 10100 29800 10109 29840
rect 10243 29800 10252 29840
rect 10292 29800 10301 29840
rect 4483 29716 4492 29756
rect 4532 29716 8372 29756
rect 8467 29716 8476 29756
rect 8516 29716 8716 29756
rect 8756 29716 8765 29756
rect 0 29672 90 29692
rect 8332 29672 8372 29716
rect 8812 29672 8852 29800
rect 10252 29756 10292 29800
rect 9091 29716 9100 29756
rect 9140 29716 9236 29756
rect 9379 29716 9388 29756
rect 9428 29716 10292 29756
rect 0 29632 76 29672
rect 116 29632 125 29672
rect 2851 29632 2860 29672
rect 2900 29632 3031 29672
rect 3148 29632 4012 29672
rect 4052 29632 4061 29672
rect 4505 29632 4588 29672
rect 4628 29632 4636 29672
rect 4676 29632 4685 29672
rect 8332 29632 8852 29672
rect 8995 29632 9004 29672
rect 9044 29632 9140 29672
rect 0 29612 90 29632
rect 3148 29420 3188 29632
rect 2092 29380 3188 29420
rect 3292 29548 6412 29588
rect 6452 29548 6461 29588
rect 0 29336 90 29356
rect 2092 29336 2132 29380
rect 0 29296 1324 29336
rect 1364 29296 1373 29336
rect 1459 29296 1468 29336
rect 1508 29296 2132 29336
rect 2227 29296 2236 29336
rect 2276 29296 3052 29336
rect 3092 29296 3101 29336
rect 0 29276 90 29296
rect 3292 29168 3332 29548
rect 3679 29464 3688 29504
rect 3728 29464 3770 29504
rect 3810 29464 3852 29504
rect 3892 29464 3934 29504
rect 3974 29464 4016 29504
rect 4056 29464 4065 29504
rect 6019 29464 6028 29504
rect 6068 29464 6316 29504
rect 6356 29464 8908 29504
rect 8948 29464 8957 29504
rect 9100 29420 9140 29632
rect 9196 29588 9236 29716
rect 10540 29672 10580 29968
rect 13036 29924 13076 29968
rect 13324 29968 13460 30008
rect 13612 30136 13900 30176
rect 13940 30136 13949 30176
rect 13324 29924 13364 29968
rect 13612 29924 13652 30136
rect 13996 30092 14036 30304
rect 14371 30220 14380 30260
rect 14420 30220 14612 30260
rect 14361 30136 14476 30176
rect 14516 30136 14525 30176
rect 13978 30052 13987 30092
rect 14027 30052 14036 30092
rect 14179 30052 14188 30092
rect 14228 30052 14237 30092
rect 14188 29924 14228 30052
rect 14361 29924 14401 30136
rect 14572 30092 14612 30220
rect 14458 30052 14467 30092
rect 14507 30052 14612 30092
rect 14668 30008 14708 30304
rect 16771 30220 16780 30260
rect 16820 30220 19892 30260
rect 20039 30220 20048 30260
rect 20088 30220 20130 30260
rect 20170 30220 20212 30260
rect 20252 30220 20294 30260
rect 20334 30220 20376 30260
rect 20416 30220 20425 30260
rect 19852 30176 19892 30220
rect 21510 30176 21600 30196
rect 16291 30136 16300 30176
rect 16340 30136 19756 30176
rect 19796 30136 19805 30176
rect 19852 30136 20180 30176
rect 21091 30136 21100 30176
rect 21140 30136 21600 30176
rect 14825 30052 14947 30092
rect 14996 30052 15005 30092
rect 15305 30052 15340 30092
rect 15380 30052 15436 30092
rect 15476 30052 15485 30092
rect 15820 30052 17836 30092
rect 17876 30052 17885 30092
rect 18691 30052 18700 30092
rect 18740 30052 18892 30092
rect 18932 30052 18941 30092
rect 19843 30052 19852 30092
rect 19892 30052 19996 30092
rect 20036 30052 20045 30092
rect 14668 29968 14804 30008
rect 14851 29968 14860 30008
rect 14900 29968 15476 30008
rect 14764 29924 14804 29968
rect 10627 29884 10636 29924
rect 10676 29915 10807 29924
rect 10676 29884 10732 29915
rect 10772 29884 10807 29915
rect 11081 29884 11212 29924
rect 11252 29884 11261 29924
rect 13027 29884 13036 29924
rect 13076 29884 13085 29924
rect 13315 29884 13324 29924
rect 13364 29884 13373 29924
rect 13498 29884 13507 29924
rect 13547 29884 13556 29924
rect 13612 29884 13655 29924
rect 13695 29884 13704 29924
rect 13889 29884 13898 29924
rect 13938 29884 13947 29924
rect 14146 29884 14155 29924
rect 14195 29884 14228 29924
rect 14352 29884 14361 29924
rect 14401 29884 14410 29924
rect 14611 29884 14620 29924
rect 14660 29884 14669 29924
rect 14746 29884 14755 29924
rect 14795 29884 14804 29924
rect 14851 29884 14860 29924
rect 14900 29884 15134 29924
rect 15174 29884 15183 29924
rect 15436 29915 15476 29968
rect 10732 29866 10772 29875
rect 11212 29866 11252 29875
rect 11434 29800 11443 29840
rect 11483 29800 11788 29840
rect 11828 29800 11837 29840
rect 12233 29800 12268 29840
rect 12308 29800 12364 29840
rect 12404 29800 12413 29840
rect 13516 29756 13556 29884
rect 13900 29840 13940 29884
rect 14620 29840 14660 29884
rect 14860 29840 14900 29884
rect 15436 29866 15476 29875
rect 15820 29840 15860 30052
rect 16204 29968 18260 30008
rect 18979 29968 18988 30008
rect 19028 29968 19180 30008
rect 19220 29968 19229 30008
rect 16204 29840 16244 29968
rect 18220 29924 18260 29968
rect 16378 29884 16387 29924
rect 16436 29884 16567 29924
rect 16675 29884 16684 29924
rect 16724 29884 16855 29924
rect 17146 29884 17155 29924
rect 17195 29884 17204 29924
rect 17251 29884 17260 29924
rect 17300 29884 17431 29924
rect 17548 29884 17644 29924
rect 17684 29884 17693 29924
rect 18220 29915 18412 29924
rect 17164 29840 17204 29884
rect 13786 29800 13795 29840
rect 13835 29800 13844 29840
rect 13891 29800 13900 29840
rect 13940 29800 13985 29840
rect 14179 29800 14188 29840
rect 14228 29800 14275 29840
rect 14315 29800 14359 29840
rect 14580 29800 14660 29840
rect 14764 29800 14900 29840
rect 15811 29800 15820 29840
rect 15860 29800 15869 29840
rect 16195 29800 16204 29840
rect 16244 29800 16253 29840
rect 17164 29800 17452 29840
rect 17492 29800 17501 29840
rect 13516 29716 13708 29756
rect 13748 29716 13757 29756
rect 13804 29672 13844 29800
rect 9283 29632 9292 29672
rect 9332 29632 10580 29672
rect 11539 29632 11548 29672
rect 11588 29632 11788 29672
rect 11828 29632 11837 29672
rect 12499 29632 12508 29672
rect 12548 29632 12748 29672
rect 12788 29632 12797 29672
rect 13171 29632 13180 29672
rect 13220 29632 13229 29672
rect 13498 29632 13507 29672
rect 13547 29632 13556 29672
rect 13804 29632 14476 29672
rect 14516 29632 14525 29672
rect 9196 29548 11980 29588
rect 12020 29548 12029 29588
rect 13180 29420 13220 29632
rect 13516 29504 13556 29632
rect 14580 29504 14620 29800
rect 14764 29756 14804 29800
rect 17548 29756 17588 29884
rect 18260 29884 18412 29915
rect 18452 29884 18461 29924
rect 18700 29915 18740 29924
rect 18220 29866 18260 29875
rect 19066 29884 19075 29924
rect 19115 29884 19124 29924
rect 19377 29884 19386 29924
rect 19426 29884 19948 29924
rect 19988 29884 19997 29924
rect 17731 29800 17740 29840
rect 17780 29800 17789 29840
rect 14755 29716 14764 29756
rect 14804 29716 14813 29756
rect 14947 29716 14956 29756
rect 14996 29716 15820 29756
rect 15860 29716 15869 29756
rect 16387 29716 16396 29756
rect 16436 29716 17588 29756
rect 17740 29672 17780 29800
rect 18700 29756 18740 29875
rect 19084 29840 19124 29884
rect 20140 29840 20180 30136
rect 21510 30116 21600 30136
rect 20371 30052 20380 30092
rect 20420 30052 21004 30092
rect 21044 30052 21053 30092
rect 19084 29800 19276 29840
rect 19316 29800 19325 29840
rect 19625 29800 19756 29840
rect 19796 29800 19805 29840
rect 20131 29800 20140 29840
rect 20180 29800 20189 29840
rect 18700 29716 19124 29756
rect 14851 29632 14860 29672
rect 14900 29632 15139 29672
rect 15179 29632 15188 29672
rect 15427 29632 15436 29672
rect 15476 29632 15580 29672
rect 15620 29632 15629 29672
rect 15907 29632 15916 29672
rect 15956 29632 15964 29672
rect 16004 29632 16087 29672
rect 16675 29632 16684 29672
rect 16724 29632 16733 29672
rect 17059 29632 17068 29672
rect 17108 29632 17932 29672
rect 17972 29632 17981 29672
rect 13516 29464 14620 29504
rect 3484 29380 9140 29420
rect 9283 29380 9292 29420
rect 9332 29380 11636 29420
rect 13180 29380 13748 29420
rect 3484 29252 3524 29380
rect 11596 29336 11636 29380
rect 13708 29336 13748 29380
rect 14381 29380 16108 29420
rect 16148 29380 16157 29420
rect 4003 29296 4012 29336
rect 4052 29296 4340 29336
rect 4435 29296 4444 29336
rect 4484 29296 4876 29336
rect 4916 29296 4925 29336
rect 6307 29296 6316 29336
rect 6356 29296 6508 29336
rect 6548 29296 6557 29336
rect 6604 29296 11308 29336
rect 11348 29296 11357 29336
rect 11596 29296 12940 29336
rect 12980 29296 12989 29336
rect 13385 29296 13516 29336
rect 13556 29296 13565 29336
rect 13699 29296 13708 29336
rect 13748 29296 13757 29336
rect 451 29128 460 29168
rect 500 29128 1228 29168
rect 1268 29128 1277 29168
rect 1481 29128 1612 29168
rect 1652 29128 1661 29168
rect 1865 29128 1996 29168
rect 2036 29128 2045 29168
rect 2467 29128 2476 29168
rect 2516 29128 2787 29168
rect 2827 29128 2836 29168
rect 3139 29128 3148 29168
rect 3188 29128 3197 29168
rect 3274 29159 3332 29168
rect 3148 29084 3188 29128
rect 3274 29119 3283 29159
rect 3323 29119 3332 29159
rect 3388 29212 3524 29252
rect 4300 29252 4340 29296
rect 6604 29252 6644 29296
rect 14381 29252 14421 29380
rect 14467 29296 14476 29336
rect 14516 29296 14525 29336
rect 15187 29296 15196 29336
rect 15236 29296 16244 29336
rect 4300 29212 6644 29252
rect 9235 29212 9244 29252
rect 9284 29212 14421 29252
rect 3388 29126 3428 29212
rect 14476 29168 14516 29296
rect 15436 29212 15628 29252
rect 15668 29212 15677 29252
rect 15436 29168 15476 29212
rect 4291 29128 4300 29168
rect 4340 29128 4349 29168
rect 4675 29128 4684 29168
rect 4724 29128 5548 29168
rect 5588 29128 5597 29168
rect 7267 29128 7276 29168
rect 7316 29128 7564 29168
rect 7604 29128 7613 29168
rect 8873 29128 9004 29168
rect 9044 29128 9292 29168
rect 9332 29128 9388 29168
rect 9428 29128 9437 29168
rect 9484 29128 9772 29168
rect 9812 29128 10004 29168
rect 10217 29128 10348 29168
rect 10388 29128 10397 29168
rect 10627 29128 10636 29168
rect 10676 29128 10828 29168
rect 10868 29128 10877 29168
rect 14476 29128 14668 29168
rect 14708 29128 14717 29168
rect 15427 29128 15436 29168
rect 15476 29128 15485 29168
rect 3274 29118 3332 29119
rect 3379 29086 3388 29126
rect 3428 29086 3437 29126
rect 4300 29084 4340 29128
rect 6124 29084 6164 29093
rect 7852 29084 7892 29093
rect 9484 29084 9524 29128
rect 9964 29084 10004 29128
rect 15628 29117 15764 29126
rect 10924 29084 10964 29093
rect 13324 29084 13364 29093
rect 15628 29086 15724 29117
rect 2537 29044 2668 29084
rect 2708 29044 2717 29084
rect 2851 29044 2860 29084
rect 2925 29044 3031 29084
rect 3148 29044 3157 29084
rect 3197 29044 3235 29084
rect 3619 29044 3628 29084
rect 3668 29044 3724 29084
rect 3764 29044 3799 29084
rect 3898 29044 3907 29084
rect 3947 29044 3956 29084
rect 4300 29044 4876 29084
rect 4916 29044 4925 29084
rect 6778 29044 6787 29084
rect 6827 29044 6836 29084
rect 6883 29044 6892 29084
rect 6932 29044 7316 29084
rect 7363 29044 7372 29084
rect 7412 29044 7468 29084
rect 7508 29044 7543 29084
rect 8362 29044 8371 29084
rect 8411 29044 8908 29084
rect 8948 29044 8957 29084
rect 9475 29044 9484 29084
rect 9524 29044 9533 29084
rect 9850 29044 9859 29084
rect 9899 29044 9908 29084
rect 9955 29044 9964 29084
rect 10004 29044 10013 29084
rect 10313 29044 10444 29084
rect 10484 29044 10493 29084
rect 10793 29044 10924 29084
rect 10964 29044 10973 29084
rect 11299 29044 11308 29084
rect 11348 29044 11412 29084
rect 11452 29044 11479 29084
rect 11971 29044 11980 29084
rect 12020 29044 12076 29084
rect 12116 29044 12151 29084
rect 13193 29044 13324 29084
rect 13364 29044 13373 29084
rect 14170 29044 14179 29084
rect 14219 29044 14860 29084
rect 14900 29044 14909 29084
rect 0 29000 90 29020
rect 3916 29000 3956 29044
rect 0 28960 2996 29000
rect 3523 28960 3532 29000
rect 3572 28960 3956 29000
rect 4003 28960 4012 29000
rect 4052 28960 4061 29000
rect 4217 28960 4300 29000
rect 4340 28960 4348 29000
rect 4388 28960 4397 29000
rect 0 28940 90 28960
rect 1843 28876 1852 28916
rect 1892 28876 2132 28916
rect 2441 28876 2572 28916
rect 2612 28876 2621 28916
rect 2092 28832 2132 28876
rect 2956 28832 2996 28960
rect 4012 28916 4052 28960
rect 3043 28876 3052 28916
rect 3092 28876 3916 28916
rect 3956 28876 3965 28916
rect 4012 28876 4876 28916
rect 4916 28876 4925 28916
rect 6124 28832 6164 29044
rect 6796 29000 6836 29044
rect 7276 29000 7316 29044
rect 7852 29000 7892 29044
rect 6787 28960 6796 29000
rect 6836 28960 6883 29000
rect 7267 28960 7276 29000
rect 7316 28960 7325 29000
rect 7367 28960 7376 29000
rect 7416 28960 7892 29000
rect 9868 29000 9908 29044
rect 10924 29035 10964 29044
rect 13324 29035 13364 29044
rect 9868 28960 10828 29000
rect 10868 28960 10877 29000
rect 11020 28960 12844 29000
rect 12884 28960 12893 29000
rect 14249 28960 14284 29000
rect 14324 28960 14380 29000
rect 14420 28960 14429 29000
rect 14481 28960 14490 29000
rect 14530 28960 15052 29000
rect 15092 28960 15101 29000
rect 11020 28916 11060 28960
rect 15628 28916 15668 29086
rect 15724 29068 15764 29077
rect 15835 29084 15875 29093
rect 15944 29044 15953 29084
rect 15993 29044 16002 29084
rect 15835 29000 15875 29044
rect 15715 28960 15724 29000
rect 15764 28960 15875 29000
rect 15962 29000 16002 29044
rect 16204 29000 16244 29296
rect 16684 29252 16724 29632
rect 19084 29588 19124 29716
rect 21510 29672 21600 29692
rect 19363 29632 19372 29672
rect 19412 29632 20428 29672
rect 20468 29632 20477 29672
rect 21187 29632 21196 29672
rect 21236 29632 21600 29672
rect 21510 29612 21600 29632
rect 19084 29548 19892 29588
rect 18799 29464 18808 29504
rect 18848 29464 18890 29504
rect 18930 29464 18972 29504
rect 19012 29464 19054 29504
rect 19094 29464 19136 29504
rect 19176 29464 19185 29504
rect 19852 29336 19892 29548
rect 17609 29296 17740 29336
rect 17780 29296 17789 29336
rect 19843 29296 19852 29336
rect 19892 29296 19901 29336
rect 20371 29296 20380 29336
rect 20420 29296 20620 29336
rect 20660 29296 20669 29336
rect 16684 29212 17684 29252
rect 16291 29128 16300 29168
rect 16340 29128 16349 29168
rect 16300 29084 16340 29128
rect 17548 29084 17588 29093
rect 16291 29044 16300 29084
rect 16340 29044 16387 29084
rect 17251 29044 17260 29084
rect 17300 29044 17309 29084
rect 17644 29084 17684 29212
rect 21510 29168 21600 29188
rect 17923 29128 17932 29168
rect 17972 29128 18164 29168
rect 20131 29128 20140 29168
rect 20180 29128 20524 29168
rect 20564 29128 20573 29168
rect 20995 29128 21004 29168
rect 21044 29128 21600 29168
rect 18124 29084 18164 29128
rect 21510 29108 21600 29128
rect 18220 29084 18260 29093
rect 19660 29084 19700 29093
rect 17644 29044 17918 29084
rect 17958 29044 17967 29084
rect 18115 29044 18124 29084
rect 18164 29044 18173 29084
rect 18403 29044 18412 29084
rect 18452 29044 18583 29084
rect 19529 29044 19660 29084
rect 19700 29044 19709 29084
rect 17260 29000 17300 29044
rect 15962 28960 16108 29000
rect 16148 28960 16157 29000
rect 16204 28960 17300 29000
rect 17548 29000 17588 29044
rect 17548 28960 18124 29000
rect 18164 28960 18173 29000
rect 8393 28876 8524 28916
rect 8564 28876 8573 28916
rect 9091 28876 9100 28916
rect 9140 28876 9628 28916
rect 9668 28876 9677 28916
rect 10051 28876 10060 28916
rect 10100 28876 11060 28916
rect 11587 28876 11596 28916
rect 11636 28876 12172 28916
rect 12212 28876 12556 28916
rect 12596 28876 12605 28916
rect 14899 28876 14908 28916
rect 14948 28876 15092 28916
rect 15628 28876 15820 28916
rect 15860 28876 15869 28916
rect 16099 28876 16108 28916
rect 16148 28876 17068 28916
rect 17108 28876 17117 28916
rect 17251 28876 17260 28916
rect 17300 28876 18019 28916
rect 18059 28876 18068 28916
rect 15052 28832 15092 28876
rect 18220 28832 18260 29044
rect 19660 29035 19700 29044
rect 20035 28876 20044 28916
rect 20084 28876 20093 28916
rect 20044 28832 20084 28876
rect 2092 28792 2860 28832
rect 2900 28792 2909 28832
rect 2956 28792 6068 28832
rect 6124 28792 9004 28832
rect 9044 28792 9053 28832
rect 9571 28792 9580 28832
rect 9620 28792 10348 28832
rect 10388 28792 10397 28832
rect 15052 28792 15532 28832
rect 15572 28792 15581 28832
rect 16675 28792 16684 28832
rect 16724 28792 18260 28832
rect 19948 28792 20084 28832
rect 1315 28708 1324 28748
rect 1364 28708 4820 28748
rect 4919 28708 4928 28748
rect 4968 28708 5010 28748
rect 5050 28708 5092 28748
rect 5132 28708 5174 28748
rect 5214 28708 5256 28748
rect 5296 28708 5305 28748
rect 0 28664 90 28684
rect 0 28624 1132 28664
rect 1172 28624 1181 28664
rect 3628 28624 4012 28664
rect 4052 28624 4061 28664
rect 0 28604 90 28624
rect 3628 28580 3668 28624
rect 2851 28540 2860 28580
rect 2900 28540 3284 28580
rect 3610 28540 3619 28580
rect 3659 28540 3668 28580
rect 4073 28540 4204 28580
rect 4244 28540 4253 28580
rect 3244 28496 3284 28540
rect 4780 28496 4820 28708
rect 6028 28664 6068 28792
rect 19948 28748 19988 28792
rect 8812 28708 18028 28748
rect 18068 28708 18077 28748
rect 18124 28708 19988 28748
rect 20039 28708 20048 28748
rect 20088 28708 20130 28748
rect 20170 28708 20212 28748
rect 20252 28708 20294 28748
rect 20334 28708 20376 28748
rect 20416 28708 20425 28748
rect 4876 28624 5972 28664
rect 6028 28624 8716 28664
rect 8756 28624 8765 28664
rect 4876 28580 4916 28624
rect 5932 28580 5972 28624
rect 8812 28580 8852 28708
rect 18124 28664 18164 28708
rect 21510 28664 21600 28684
rect 10444 28624 13940 28664
rect 10444 28580 10484 28624
rect 4867 28540 4876 28580
rect 4916 28540 4925 28580
rect 5129 28540 5212 28580
rect 5252 28540 5260 28580
rect 5300 28540 5309 28580
rect 5932 28540 6412 28580
rect 6452 28540 6461 28580
rect 6665 28540 6796 28580
rect 6836 28540 6845 28580
rect 8803 28540 8812 28580
rect 8852 28540 8861 28580
rect 8995 28540 9004 28580
rect 9044 28540 9244 28580
rect 9284 28540 9524 28580
rect 9619 28540 9628 28580
rect 9668 28540 10156 28580
rect 10196 28540 10205 28580
rect 10387 28540 10396 28580
rect 10436 28540 10484 28580
rect 10531 28540 10540 28580
rect 10580 28540 11308 28580
rect 11348 28540 11357 28580
rect 11683 28540 11692 28580
rect 11732 28540 12748 28580
rect 12788 28540 12980 28580
rect 2860 28456 3148 28496
rect 3188 28456 3197 28496
rect 3244 28456 3572 28496
rect 3907 28456 3916 28496
rect 3956 28456 3998 28496
rect 4038 28456 4087 28496
rect 4291 28456 4300 28496
rect 4340 28456 4349 28496
rect 4780 28456 9428 28496
rect 2860 28412 2900 28456
rect 3532 28412 3572 28456
rect 4300 28412 4340 28456
rect 1481 28372 1516 28412
rect 1556 28372 1612 28412
rect 1652 28372 1661 28412
rect 2633 28372 2764 28412
rect 2804 28372 2900 28412
rect 3043 28372 3052 28412
rect 3092 28372 3287 28412
rect 3327 28372 3336 28412
rect 3523 28372 3532 28412
rect 3572 28372 3581 28412
rect 4300 28403 4387 28412
rect 2764 28354 2804 28363
rect 4340 28372 4387 28403
rect 4457 28372 4588 28412
rect 4628 28372 4637 28412
rect 4771 28372 4780 28412
rect 4845 28372 4951 28412
rect 5059 28372 5068 28412
rect 5108 28372 5356 28412
rect 5396 28372 5405 28412
rect 6604 28403 6796 28412
rect 4300 28354 4340 28363
rect 6644 28372 6796 28403
rect 6836 28372 6845 28412
rect 7066 28372 7075 28412
rect 7115 28372 7124 28412
rect 7171 28372 7180 28412
rect 7220 28372 7276 28412
rect 7316 28372 7351 28412
rect 7433 28372 7564 28412
rect 7604 28372 7613 28412
rect 7939 28372 7948 28412
rect 7988 28403 8180 28412
rect 7988 28372 8140 28403
rect 6604 28354 6644 28363
rect 0 28328 90 28348
rect 7084 28328 7124 28372
rect 8323 28372 8332 28412
rect 8372 28403 8660 28412
rect 8372 28372 8620 28403
rect 0 28288 460 28328
rect 500 28288 509 28328
rect 3276 28288 3340 28328
rect 3380 28288 3427 28328
rect 3467 28288 3724 28328
rect 3764 28288 3773 28328
rect 4483 28288 4492 28328
rect 4532 28288 4541 28328
rect 4684 28288 4707 28328
rect 4747 28288 4756 28328
rect 4963 28288 4972 28328
rect 5012 28288 5644 28328
rect 5684 28288 5693 28328
rect 7084 28288 7468 28328
rect 7508 28288 7517 28328
rect 7651 28288 7660 28328
rect 7700 28288 7756 28328
rect 7796 28288 7860 28328
rect 0 28268 90 28288
rect 2467 28204 2476 28244
rect 2516 28204 2956 28244
rect 2996 28204 3005 28244
rect 4492 28160 4532 28288
rect 4684 28160 4724 28288
rect 7660 28244 7700 28288
rect 7267 28204 7276 28244
rect 7316 28204 7700 28244
rect 8140 28160 8180 28363
rect 8620 28354 8660 28363
rect 9388 28328 9428 28456
rect 9484 28412 9524 28540
rect 10627 28456 10636 28496
rect 10676 28456 12596 28496
rect 12556 28412 12596 28456
rect 12940 28412 12980 28540
rect 13900 28496 13940 28624
rect 14860 28624 18164 28664
rect 19843 28624 19852 28664
rect 19892 28624 21600 28664
rect 13987 28540 13996 28580
rect 14036 28540 14764 28580
rect 14804 28540 14813 28580
rect 14860 28496 14900 28624
rect 21510 28604 21600 28624
rect 15689 28540 15820 28580
rect 15860 28540 15869 28580
rect 17321 28540 17452 28580
rect 17492 28540 17501 28580
rect 19075 28540 19084 28580
rect 19124 28540 19276 28580
rect 19316 28540 19325 28580
rect 19939 28540 19948 28580
rect 19988 28540 20035 28580
rect 20075 28540 20119 28580
rect 19276 28496 19316 28540
rect 13900 28456 14900 28496
rect 16291 28456 16300 28496
rect 16340 28456 16684 28496
rect 16724 28456 17684 28496
rect 17644 28412 17684 28456
rect 19276 28456 19988 28496
rect 19276 28412 19316 28456
rect 19948 28412 19988 28456
rect 9484 28372 9772 28412
rect 9812 28372 9964 28412
rect 10004 28403 10772 28412
rect 10004 28372 10732 28403
rect 11587 28372 11596 28412
rect 11636 28372 11980 28412
rect 12020 28372 12029 28412
rect 12547 28372 12556 28412
rect 12596 28372 12605 28412
rect 12940 28403 13844 28412
rect 12940 28372 13804 28403
rect 10732 28354 10772 28363
rect 13987 28372 13996 28412
rect 14036 28372 14380 28412
rect 14420 28372 14668 28412
rect 14708 28372 14717 28412
rect 15628 28403 15820 28412
rect 13804 28354 13844 28363
rect 15668 28372 15820 28403
rect 15860 28372 15869 28412
rect 16003 28372 16012 28412
rect 16052 28372 16204 28412
rect 16244 28372 16588 28412
rect 16628 28372 16637 28412
rect 17155 28372 17164 28412
rect 17204 28403 17335 28412
rect 17204 28372 17260 28403
rect 15628 28354 15668 28363
rect 17300 28372 17335 28403
rect 17635 28372 17644 28412
rect 17684 28372 17693 28412
rect 18019 28372 18028 28412
rect 18068 28403 18932 28412
rect 18068 28372 18892 28403
rect 17260 28354 17300 28363
rect 19276 28403 19412 28412
rect 19276 28372 19372 28403
rect 18892 28354 18932 28363
rect 19372 28354 19412 28363
rect 19462 28352 19471 28392
rect 19511 28352 19520 28392
rect 19939 28372 19948 28412
rect 19988 28372 19997 28412
rect 20131 28372 20140 28412
rect 20180 28372 20236 28412
rect 20276 28372 20311 28412
rect 8873 28288 9004 28328
rect 9044 28288 9053 28328
rect 9379 28288 9388 28328
rect 9428 28288 9437 28328
rect 9763 28288 9772 28328
rect 9812 28288 9821 28328
rect 9996 28288 10060 28328
rect 10100 28288 10156 28328
rect 10196 28288 10205 28328
rect 11299 28288 11308 28328
rect 11348 28288 12364 28328
rect 12404 28288 12413 28328
rect 9772 28244 9812 28288
rect 19468 28244 19508 28352
rect 19592 28330 19601 28370
rect 19641 28330 19700 28370
rect 8707 28204 8716 28244
rect 8756 28204 9812 28244
rect 10003 28204 10012 28244
rect 10052 28204 12980 28244
rect 17923 28204 17932 28244
rect 17972 28204 19508 28244
rect 19660 28244 19700 28330
rect 19660 28204 19892 28244
rect 12940 28160 12980 28204
rect 3619 28120 3628 28160
rect 3668 28120 4003 28160
rect 4043 28120 4052 28160
rect 4492 28120 4588 28160
rect 4628 28120 4637 28160
rect 4684 28120 8180 28160
rect 10147 28120 10156 28160
rect 10196 28120 11788 28160
rect 11828 28120 11837 28160
rect 12115 28120 12124 28160
rect 12164 28120 12844 28160
rect 12884 28120 12893 28160
rect 12940 28120 19564 28160
rect 19604 28120 19613 28160
rect 19747 28120 19756 28160
rect 19796 28120 19805 28160
rect 4684 28076 4724 28120
rect 3043 28036 3052 28076
rect 3092 28036 4724 28076
rect 9955 28036 9964 28076
rect 10004 28036 13612 28076
rect 13652 28036 13661 28076
rect 0 27992 90 28012
rect 0 27952 1996 27992
rect 2036 27952 2045 27992
rect 3679 27952 3688 27992
rect 3728 27952 3770 27992
rect 3810 27952 3852 27992
rect 3892 27952 3934 27992
rect 3974 27952 4016 27992
rect 4056 27952 4065 27992
rect 10051 27952 10060 27992
rect 10100 27952 12980 27992
rect 0 27932 90 27952
rect 6019 27868 6028 27908
rect 6068 27868 10100 27908
rect 10060 27824 10100 27868
rect 10636 27868 11540 27908
rect 10636 27824 10676 27868
rect 1459 27784 1468 27824
rect 1508 27784 1804 27824
rect 1844 27784 1853 27824
rect 2659 27784 2668 27824
rect 2708 27784 3052 27824
rect 3092 27784 5204 27824
rect 7555 27784 7564 27824
rect 7604 27784 8332 27824
rect 8372 27784 8381 27824
rect 10060 27784 10636 27824
rect 10676 27784 10685 27824
rect 11011 27784 11020 27824
rect 11060 27784 11212 27824
rect 11252 27784 11261 27824
rect 172 27700 1364 27740
rect 2467 27700 2476 27740
rect 2516 27700 3188 27740
rect 0 27656 90 27676
rect 172 27656 212 27700
rect 1324 27656 1364 27700
rect 2668 27656 2708 27700
rect 0 27616 212 27656
rect 259 27616 268 27656
rect 308 27616 1228 27656
rect 1268 27616 1277 27656
rect 1324 27616 2516 27656
rect 2659 27616 2668 27656
rect 2708 27616 2717 27656
rect 0 27596 90 27616
rect 2476 27572 2516 27616
rect 2860 27572 2900 27581
rect 1603 27532 1612 27572
rect 1652 27532 2420 27572
rect 2467 27532 2476 27572
rect 2516 27532 2525 27572
rect 2729 27532 2764 27572
rect 2804 27532 2860 27572
rect 2900 27532 2964 27572
rect 2380 27404 2420 27532
rect 2860 27523 2900 27532
rect 3148 27488 3188 27700
rect 3244 27572 3284 27784
rect 3331 27700 3340 27740
rect 3380 27700 3532 27740
rect 3572 27700 3916 27740
rect 3956 27700 3965 27740
rect 4291 27700 4300 27740
rect 4340 27700 4349 27740
rect 3628 27616 4148 27656
rect 3628 27572 3668 27616
rect 3235 27532 3244 27572
rect 3284 27532 3293 27572
rect 3468 27532 3532 27572
rect 3572 27532 3628 27572
rect 3668 27532 3677 27572
rect 3785 27532 3907 27572
rect 3956 27532 3965 27572
rect 3532 27488 3572 27532
rect 4108 27488 4148 27616
rect 4300 27572 4340 27700
rect 4579 27616 4588 27656
rect 4628 27616 4876 27656
rect 4916 27616 5059 27656
rect 5099 27616 5108 27656
rect 5164 27572 5204 27784
rect 5251 27700 5260 27740
rect 5300 27700 5780 27740
rect 10819 27700 10828 27740
rect 10868 27700 11212 27740
rect 11252 27700 11261 27740
rect 5740 27656 5780 27700
rect 5251 27616 5260 27656
rect 5300 27616 5539 27656
rect 5579 27616 5588 27656
rect 5731 27616 5740 27656
rect 5780 27616 5789 27656
rect 9283 27616 9292 27656
rect 9332 27616 9341 27656
rect 9763 27616 9772 27656
rect 9812 27616 11444 27656
rect 7372 27572 7412 27581
rect 7948 27572 7988 27581
rect 9292 27572 9332 27616
rect 11404 27572 11444 27616
rect 4300 27532 4483 27572
rect 4523 27532 4532 27572
rect 4588 27532 4919 27572
rect 4959 27532 4968 27572
rect 5155 27532 5164 27572
rect 5204 27532 5213 27572
rect 5410 27532 5419 27572
rect 5459 27532 5588 27572
rect 5635 27532 5644 27572
rect 5684 27532 5815 27572
rect 6115 27532 6124 27572
rect 6164 27532 6892 27572
rect 6932 27532 6941 27572
rect 7788 27532 7852 27572
rect 7892 27532 7948 27572
rect 7988 27532 8332 27572
rect 8372 27532 8381 27572
rect 9065 27532 9196 27572
rect 9236 27532 9245 27572
rect 9292 27532 9580 27572
rect 9620 27532 9629 27572
rect 10827 27532 10836 27572
rect 10876 27532 11308 27572
rect 11348 27532 11357 27572
rect 11500 27572 11540 27868
rect 12940 27824 12980 27952
rect 13036 27952 14860 27992
rect 14900 27952 14909 27992
rect 18799 27952 18808 27992
rect 18848 27952 18890 27992
rect 18930 27952 18972 27992
rect 19012 27952 19054 27992
rect 19094 27952 19136 27992
rect 19176 27952 19185 27992
rect 13036 27824 13076 27952
rect 12940 27784 13076 27824
rect 13804 27868 16780 27908
rect 16820 27868 16829 27908
rect 13804 27740 13844 27868
rect 14563 27784 14572 27824
rect 14612 27784 15244 27824
rect 15284 27784 15293 27824
rect 16099 27784 16108 27824
rect 16148 27784 16492 27824
rect 16532 27784 16541 27824
rect 12739 27700 12748 27740
rect 12788 27700 13844 27740
rect 14380 27572 14420 27581
rect 16300 27572 16340 27581
rect 16780 27572 16820 27868
rect 17443 27700 17452 27740
rect 17492 27700 18508 27740
rect 18548 27700 18557 27740
rect 19756 27656 19796 28120
rect 19852 27824 19892 28204
rect 21510 28160 21600 28180
rect 19939 28120 19948 28160
rect 19988 28120 21600 28160
rect 21510 28100 21600 28120
rect 19843 27784 19852 27824
rect 19892 27784 19901 27824
rect 20035 27700 20044 27740
rect 20084 27700 20372 27740
rect 20332 27656 20372 27700
rect 21510 27656 21600 27676
rect 19756 27616 20276 27656
rect 20332 27616 21600 27656
rect 18028 27572 18068 27581
rect 19660 27572 19700 27581
rect 20236 27572 20276 27616
rect 21510 27596 21600 27616
rect 11500 27532 12268 27572
rect 12308 27532 12652 27572
rect 12692 27532 12701 27572
rect 13001 27532 13132 27572
rect 13172 27532 13181 27572
rect 13795 27532 13804 27572
rect 13844 27532 14380 27572
rect 15043 27532 15052 27572
rect 15092 27532 15436 27572
rect 15476 27532 15485 27572
rect 15811 27532 15820 27572
rect 15860 27532 16300 27572
rect 16771 27532 16780 27572
rect 16820 27532 16829 27572
rect 17155 27532 17164 27572
rect 17204 27532 18028 27572
rect 18377 27532 18412 27572
rect 18452 27532 18508 27572
rect 18548 27532 18557 27572
rect 19171 27532 19180 27572
rect 19220 27532 19660 27572
rect 4588 27488 4628 27532
rect 3148 27448 3572 27488
rect 3881 27448 4012 27488
rect 4052 27448 4061 27488
rect 4108 27448 4628 27488
rect 4785 27448 4794 27488
rect 4834 27448 5260 27488
rect 5300 27448 5309 27488
rect 5548 27404 5588 27532
rect 7372 27488 7412 27532
rect 7948 27523 7988 27532
rect 9196 27488 9236 27532
rect 11404 27523 11444 27532
rect 14380 27523 14420 27532
rect 7372 27448 7756 27488
rect 7796 27448 7805 27488
rect 8044 27448 8908 27488
rect 8948 27448 8957 27488
rect 9196 27448 10444 27488
rect 10484 27448 10493 27488
rect 11500 27448 12652 27488
rect 12692 27448 12701 27488
rect 8044 27404 8084 27448
rect 11500 27404 11540 27448
rect 15052 27404 15092 27532
rect 16300 27523 16340 27532
rect 18028 27523 18068 27532
rect 19660 27523 19700 27532
rect 19852 27532 19991 27572
rect 20031 27532 20040 27572
rect 20122 27532 20131 27572
rect 20171 27532 20180 27572
rect 20227 27532 20236 27572
rect 20276 27532 20285 27572
rect 19852 27488 19892 27532
rect 20140 27488 20180 27532
rect 19843 27448 19852 27488
rect 19892 27448 19901 27488
rect 20140 27448 20524 27488
rect 20564 27448 20573 27488
rect 2380 27364 2956 27404
rect 2996 27364 3005 27404
rect 3379 27364 3388 27404
rect 3428 27364 4204 27404
rect 4244 27364 4579 27404
rect 4619 27364 4628 27404
rect 4675 27364 4684 27404
rect 4724 27364 4855 27404
rect 5548 27364 5740 27404
rect 5780 27364 5789 27404
rect 6019 27364 6028 27404
rect 6068 27364 7700 27404
rect 7747 27364 7756 27404
rect 7796 27364 8084 27404
rect 8140 27364 9964 27404
rect 10004 27364 10013 27404
rect 11011 27364 11020 27404
rect 11060 27364 11540 27404
rect 11971 27364 11980 27404
rect 12020 27364 15092 27404
rect 16483 27364 16492 27404
rect 16532 27364 16780 27404
rect 16820 27364 16829 27404
rect 18089 27364 18220 27404
rect 18260 27364 18269 27404
rect 19267 27364 19276 27404
rect 19316 27364 20044 27404
rect 20084 27364 20093 27404
rect 20314 27364 20323 27404
rect 20363 27364 21292 27404
rect 21332 27364 21341 27404
rect 0 27320 90 27340
rect 7660 27320 7700 27364
rect 8140 27320 8180 27364
rect 0 27280 6508 27320
rect 6548 27280 6557 27320
rect 7660 27280 8180 27320
rect 9772 27280 11692 27320
rect 11732 27280 11741 27320
rect 0 27260 90 27280
rect 1315 27196 1324 27236
rect 1364 27196 2900 27236
rect 4919 27196 4928 27236
rect 4968 27196 5010 27236
rect 5050 27196 5092 27236
rect 5132 27196 5174 27236
rect 5214 27196 5256 27236
rect 5296 27196 5305 27236
rect 6595 27196 6604 27236
rect 6644 27196 9292 27236
rect 9332 27196 9341 27236
rect 2860 27152 2900 27196
rect 9772 27152 9812 27280
rect 10051 27196 10060 27236
rect 10100 27196 19468 27236
rect 19508 27196 19517 27236
rect 20039 27196 20048 27236
rect 20088 27196 20130 27236
rect 20170 27196 20212 27236
rect 20252 27196 20294 27236
rect 20334 27196 20376 27236
rect 20416 27196 20425 27236
rect 21510 27152 21600 27172
rect 2860 27112 9812 27152
rect 10060 27112 15724 27152
rect 15764 27112 17740 27152
rect 17780 27112 17789 27152
rect 18700 27112 19564 27152
rect 19604 27112 19613 27152
rect 19747 27112 19756 27152
rect 19796 27112 21600 27152
rect 10060 27068 10100 27112
rect 2947 27028 2956 27068
rect 2996 27028 3628 27068
rect 3668 27028 5644 27068
rect 5684 27028 5693 27068
rect 7337 27028 7468 27068
rect 7508 27028 7517 27068
rect 7817 27028 7900 27068
rect 7940 27028 7948 27068
rect 7988 27028 7997 27068
rect 8323 27028 8332 27068
rect 8372 27028 10100 27068
rect 10579 27028 10588 27068
rect 10628 27028 10828 27068
rect 10868 27028 10877 27068
rect 11177 27028 11260 27068
rect 11300 27028 11308 27068
rect 11348 27028 11357 27068
rect 0 26984 90 27004
rect 0 26944 460 26984
rect 500 26944 509 26984
rect 2563 26944 2572 26984
rect 2612 26944 2900 26984
rect 3907 26944 3916 26984
rect 3956 26944 4588 26984
rect 4628 26944 4637 26984
rect 4972 26944 5932 26984
rect 5972 26944 5981 26984
rect 6499 26944 6508 26984
rect 6548 26944 10196 26984
rect 0 26924 90 26944
rect 2860 26900 2900 26944
rect 4972 26900 5012 26944
rect 1507 26860 1516 26900
rect 1556 26860 1804 26900
rect 1844 26860 1853 26900
rect 2633 26860 2764 26900
rect 2804 26860 2813 26900
rect 2860 26860 3148 26900
rect 3188 26860 3197 26900
rect 3401 26860 3532 26900
rect 3572 26860 3581 26900
rect 3689 26860 3811 26900
rect 3860 26860 3869 26900
rect 4387 26860 4396 26900
rect 4436 26860 5012 26900
rect 5644 26891 5684 26900
rect 2764 26842 2804 26851
rect 6019 26860 6028 26900
rect 6068 26860 6988 26900
rect 7028 26860 7124 26900
rect 5644 26816 5684 26851
rect 5644 26776 6796 26816
rect 6836 26776 6845 26816
rect 7084 26732 7124 26860
rect 7276 26891 7468 26900
rect 7316 26860 7468 26891
rect 7508 26860 7756 26900
rect 7796 26860 7805 26900
rect 7939 26860 7948 26900
rect 7988 26860 8227 26900
rect 8267 26860 8276 26900
rect 8323 26860 8332 26900
rect 8372 26860 8381 26900
rect 8515 26860 8524 26900
rect 8564 26860 8716 26900
rect 8756 26860 8765 26900
rect 8899 26860 8908 26900
rect 8948 26891 9332 26900
rect 8948 26860 9292 26891
rect 7276 26842 7316 26851
rect 8332 26816 8372 26860
rect 9641 26860 9772 26900
rect 9812 26860 9821 26900
rect 9929 26860 10003 26900
rect 10043 26860 10060 26900
rect 10100 26860 10109 26900
rect 9292 26842 9332 26851
rect 9772 26842 9812 26851
rect 10156 26816 10196 26944
rect 11596 26891 11636 27112
rect 18700 27068 18740 27112
rect 21510 27092 21600 27112
rect 16579 27028 16588 27068
rect 16628 27028 18740 27068
rect 18787 27028 18796 27068
rect 18836 27028 20140 27068
rect 20180 27028 20189 27068
rect 18700 26984 18740 27028
rect 12748 26944 12980 26984
rect 14371 26944 14380 26984
rect 14420 26944 17884 26984
rect 17924 26944 17933 26984
rect 18700 26944 18932 26984
rect 19555 26944 19564 26984
rect 19604 26944 21575 26984
rect 12748 26900 12788 26944
rect 12940 26900 12980 26944
rect 18892 26900 18932 26944
rect 12259 26860 12268 26900
rect 12308 26860 12788 26900
rect 12835 26860 12844 26900
rect 12884 26860 12893 26900
rect 12940 26860 13612 26900
rect 13652 26860 13661 26900
rect 14659 26860 14668 26900
rect 14708 26891 14900 26900
rect 14708 26860 14860 26891
rect 11596 26842 11636 26851
rect 12844 26816 12884 26860
rect 15235 26860 15244 26900
rect 15284 26860 15293 26900
rect 16361 26860 16492 26900
rect 16532 26860 16541 26900
rect 16771 26860 16780 26900
rect 16820 26860 16823 26900
rect 16863 26860 16951 26900
rect 17059 26860 17068 26900
rect 17108 26860 17239 26900
rect 18211 26860 18220 26900
rect 18260 26860 18403 26900
rect 18443 26860 18452 26900
rect 18499 26860 18508 26900
rect 18548 26860 18679 26900
rect 18883 26860 18892 26900
rect 18932 26860 18941 26900
rect 19363 26860 19372 26900
rect 19412 26891 19660 26900
rect 19412 26860 19468 26891
rect 14860 26842 14900 26851
rect 7651 26776 7660 26816
rect 7700 26776 7892 26816
rect 8131 26776 8140 26816
rect 8180 26776 8372 26816
rect 8681 26776 8812 26816
rect 8852 26776 8861 26816
rect 10147 26776 10156 26816
rect 10196 26776 10205 26816
rect 10627 26776 10636 26816
rect 10676 26776 10828 26816
rect 10868 26776 10877 26816
rect 11011 26776 11020 26816
rect 11060 26776 11540 26816
rect 12163 26776 12172 26816
rect 12212 26776 13036 26816
rect 13076 26776 13085 26816
rect 2179 26692 2188 26732
rect 2228 26692 4820 26732
rect 0 26648 90 26668
rect 0 26608 268 26648
rect 308 26608 317 26648
rect 3283 26608 3292 26648
rect 3332 26608 3572 26648
rect 4195 26608 4204 26648
rect 4244 26608 4253 26648
rect 0 26588 90 26608
rect 0 26312 90 26332
rect 0 26272 3148 26312
rect 3188 26272 3197 26312
rect 0 26252 90 26272
rect 3043 26104 3052 26144
rect 3092 26104 3427 26144
rect 3467 26104 3476 26144
rect 2668 26060 2708 26069
rect 3532 26060 3572 26608
rect 3679 26440 3688 26480
rect 3728 26440 3770 26480
rect 3810 26440 3852 26480
rect 3892 26440 3934 26480
rect 3974 26440 4016 26480
rect 4056 26440 4065 26480
rect 4204 26396 4244 26608
rect 4012 26356 4244 26396
rect 3619 26104 3628 26144
rect 3668 26104 3677 26144
rect 3628 26060 3668 26104
rect 4012 26060 4052 26356
rect 4291 26272 4300 26312
rect 4340 26272 4588 26312
rect 4628 26272 4637 26312
rect 4780 26144 4820 26692
rect 5068 26692 7028 26732
rect 7084 26692 7756 26732
rect 7796 26692 7805 26732
rect 5068 26312 5108 26692
rect 6988 26648 7028 26692
rect 7852 26648 7892 26776
rect 11500 26732 11540 26776
rect 12172 26732 12212 26776
rect 15244 26732 15284 26860
rect 16492 26842 16532 26851
rect 19508 26860 19660 26891
rect 19700 26860 19709 26900
rect 19948 26891 20276 26900
rect 19468 26842 19508 26851
rect 19988 26860 20276 26891
rect 19948 26842 19988 26851
rect 16954 26776 16963 26816
rect 17003 26776 17012 26816
rect 10387 26692 10396 26732
rect 10436 26692 11308 26732
rect 11348 26692 11357 26732
rect 11500 26692 12212 26732
rect 14659 26692 14668 26732
rect 14708 26692 15284 26732
rect 16972 26648 17012 26776
rect 17068 26776 17164 26816
rect 17204 26776 17213 26816
rect 17609 26776 17740 26816
rect 17780 26776 17789 26816
rect 18115 26776 18124 26816
rect 18164 26776 18700 26816
rect 18740 26776 18749 26816
rect 18796 26776 18892 26816
rect 18932 26776 18988 26816
rect 19028 26776 19063 26816
rect 17068 26732 17108 26776
rect 17059 26692 17068 26732
rect 17108 26692 17117 26732
rect 5827 26608 5836 26648
rect 5876 26608 6796 26648
rect 6836 26608 6845 26648
rect 6988 26608 7276 26648
rect 7316 26608 7325 26648
rect 7756 26608 7892 26648
rect 9187 26608 9196 26648
rect 9236 26608 11404 26648
rect 11444 26608 11453 26648
rect 12163 26608 12172 26648
rect 12212 26608 13276 26648
rect 13316 26608 13996 26648
rect 14036 26608 14045 26648
rect 14563 26608 14572 26648
rect 14612 26608 15052 26648
rect 15092 26608 15101 26648
rect 16649 26608 16684 26648
rect 16724 26608 16780 26648
rect 16820 26608 16829 26648
rect 16972 26608 17260 26648
rect 17300 26608 17309 26648
rect 17491 26608 17500 26648
rect 17540 26608 17740 26648
rect 17780 26608 17789 26648
rect 7756 26564 7796 26608
rect 18796 26564 18836 26776
rect 6691 26524 6700 26564
rect 6740 26524 7796 26564
rect 7843 26524 7852 26564
rect 7892 26524 10060 26564
rect 10100 26524 10109 26564
rect 13027 26524 13036 26564
rect 13076 26524 18836 26564
rect 10819 26440 10828 26480
rect 10868 26440 11308 26480
rect 11348 26440 11357 26480
rect 18799 26440 18808 26480
rect 18848 26440 18890 26480
rect 18930 26440 18972 26480
rect 19012 26440 19054 26480
rect 19094 26440 19136 26480
rect 19176 26440 19185 26480
rect 9091 26356 9100 26396
rect 9140 26356 18836 26396
rect 18796 26312 18836 26356
rect 20236 26312 20276 26860
rect 21535 26816 21575 26944
rect 21388 26776 21575 26816
rect 21388 26648 21428 26776
rect 21510 26648 21600 26668
rect 21388 26608 21600 26648
rect 21510 26588 21600 26608
rect 5011 26272 5020 26312
rect 5060 26272 5108 26312
rect 5225 26272 5308 26312
rect 5348 26272 5356 26312
rect 5396 26272 5405 26312
rect 7145 26272 7276 26312
rect 7316 26272 7325 26312
rect 9209 26272 9292 26312
rect 9371 26272 9389 26312
rect 11683 26272 11692 26312
rect 11732 26272 13132 26312
rect 13172 26272 13181 26312
rect 13865 26272 13948 26312
rect 13988 26272 13996 26312
rect 14036 26272 14045 26312
rect 18787 26272 18796 26312
rect 18836 26272 18845 26312
rect 20227 26272 20236 26312
rect 20276 26272 20285 26312
rect 6787 26188 6796 26228
rect 6836 26188 7604 26228
rect 4771 26104 4780 26144
rect 4820 26104 4829 26144
rect 5539 26104 5548 26144
rect 5588 26104 6028 26144
rect 6068 26104 6077 26144
rect 7276 26104 7468 26144
rect 7508 26104 7517 26144
rect 4110 26060 4150 26069
rect 7084 26060 7124 26069
rect 7276 26060 7316 26104
rect 7564 26060 7604 26188
rect 9676 26188 9964 26228
rect 10004 26188 10013 26228
rect 11587 26188 11596 26228
rect 11636 26188 14668 26228
rect 14708 26188 14717 26228
rect 14995 26188 15004 26228
rect 15044 26188 20524 26228
rect 20564 26188 20573 26228
rect 7913 26104 7948 26144
rect 7988 26104 8044 26144
rect 8084 26104 8093 26144
rect 8140 26104 8812 26144
rect 8852 26104 8861 26144
rect 9187 26104 9196 26144
rect 9236 26104 9620 26144
rect 8140 26060 8180 26104
rect 9580 26060 9620 26104
rect 9676 26060 9716 26188
rect 14284 26144 14324 26188
rect 21510 26144 21600 26164
rect 9929 26104 10060 26144
rect 10100 26104 10109 26144
rect 11338 26104 11347 26144
rect 11387 26104 11500 26144
rect 11540 26104 11549 26144
rect 11683 26104 11692 26144
rect 11732 26104 11863 26144
rect 11923 26104 11932 26144
rect 11972 26104 11980 26144
rect 12020 26104 12103 26144
rect 13699 26104 13708 26144
rect 13748 26104 13757 26144
rect 14275 26104 14284 26144
rect 14324 26104 14333 26144
rect 14467 26104 14476 26144
rect 14516 26104 14764 26144
rect 14804 26104 14813 26144
rect 15427 26104 15436 26144
rect 15476 26104 15485 26144
rect 15715 26104 15724 26144
rect 15764 26104 16204 26144
rect 16244 26104 16253 26144
rect 20140 26104 21600 26144
rect 10636 26060 10676 26069
rect 12268 26060 12308 26069
rect 13708 26060 13748 26104
rect 15436 26060 15476 26104
rect 16300 26060 16340 26069
rect 17356 26060 17396 26069
rect 20044 26060 20084 26069
rect 1411 26020 1420 26060
rect 1460 26020 1900 26060
rect 1940 26020 1949 26060
rect 2371 26020 2380 26060
rect 2420 26020 2668 26060
rect 2755 26020 2764 26060
rect 2804 26020 3052 26060
rect 3092 26020 3101 26060
rect 3244 26020 3287 26060
rect 3327 26020 3336 26060
rect 3523 26020 3532 26060
rect 3572 26020 3581 26060
rect 3628 26020 3806 26060
rect 3846 26020 3855 26060
rect 4012 26020 4110 26060
rect 4280 26059 4289 26060
rect 0 25976 90 25996
rect 2668 25976 2708 26020
rect 3244 25976 3284 26020
rect 4110 26011 4150 26020
rect 4252 26020 4289 26059
rect 4329 26020 4340 26060
rect 4387 26020 4396 26060
rect 4436 26020 4445 26060
rect 4675 26020 4684 26060
rect 4724 26020 4733 26060
rect 5705 26020 5836 26060
rect 5876 26020 5885 26060
rect 7124 26020 7276 26060
rect 7316 26020 7325 26060
rect 7546 26020 7555 26060
rect 7595 26020 7604 26060
rect 7651 26020 7660 26060
rect 7700 26020 7709 26060
rect 8131 26020 8140 26060
rect 8180 26020 8189 26060
rect 8614 26020 8623 26060
rect 8663 26020 8908 26060
rect 8948 26020 8957 26060
rect 9130 26020 9139 26060
rect 9179 26020 9188 26060
rect 9562 26020 9571 26060
rect 9611 26020 9620 26060
rect 9667 26020 9676 26060
rect 9716 26020 9725 26060
rect 9955 26020 9964 26060
rect 10004 26020 10156 26060
rect 10196 26020 10205 26060
rect 10339 26020 10348 26060
rect 10388 26020 10636 26060
rect 11146 26020 11155 26060
rect 11195 26020 12116 26060
rect 12259 26020 12268 26060
rect 12308 26020 12439 26060
rect 13123 26020 13132 26060
rect 13172 26020 13516 26060
rect 13556 26020 13748 26060
rect 14563 26020 14572 26060
rect 14612 26020 15214 26060
rect 15254 26020 15263 26060
rect 15329 26020 15338 26060
rect 15378 26020 15387 26060
rect 15436 26020 15820 26060
rect 15860 26020 15869 26060
rect 16340 26020 16588 26060
rect 16628 26020 16637 26060
rect 16771 26020 16780 26060
rect 16828 26020 16951 26060
rect 17251 26020 17260 26060
rect 17300 26020 17356 26060
rect 17396 26020 17431 26060
rect 18473 26020 18604 26060
rect 18644 26020 18653 26060
rect 18787 26020 18796 26060
rect 18836 26020 18967 26060
rect 19913 26020 20044 26060
rect 20084 26020 20093 26060
rect 4252 26019 4340 26020
rect 0 25936 1324 25976
rect 1364 25936 1373 25976
rect 2668 25936 3092 25976
rect 3187 25936 3196 25976
rect 3236 25936 3532 25976
rect 3572 25936 3581 25976
rect 0 25916 90 25936
rect 3052 25892 3092 25936
rect 2729 25852 2764 25892
rect 2804 25852 2860 25892
rect 2900 25852 2964 25892
rect 3052 25852 3188 25892
rect 3610 25852 3619 25892
rect 3659 25852 3668 25892
rect 3898 25852 3907 25892
rect 3947 25852 3956 25892
rect 4003 25852 4012 25892
rect 4052 25852 4183 25892
rect 0 25640 90 25660
rect 3148 25640 3188 25852
rect 3628 25724 3668 25852
rect 3916 25808 3956 25852
rect 4252 25808 4292 26019
rect 4396 25976 4436 26020
rect 4684 25976 4724 26020
rect 7084 26011 7124 26020
rect 7660 25976 7700 26020
rect 9148 25976 9188 26020
rect 10636 26011 10676 26020
rect 12076 25976 12116 26020
rect 12268 26011 12308 26020
rect 15340 25976 15380 26020
rect 16300 26011 16340 26020
rect 17356 26011 17396 26020
rect 20044 26011 20084 26020
rect 4396 25936 4532 25976
rect 4593 25936 4602 25976
rect 4642 25936 4724 25976
rect 7459 25936 7468 25976
rect 7508 25936 8140 25976
rect 8180 25936 8189 25976
rect 9148 25936 10580 25976
rect 11299 25936 11308 25976
rect 11348 25936 11500 25976
rect 11540 25936 11549 25976
rect 12067 25936 12076 25976
rect 12116 25936 12125 25976
rect 13795 25936 13804 25976
rect 13844 25936 13996 25976
rect 14036 25936 14044 25976
rect 14084 25936 14093 25976
rect 15331 25936 15340 25976
rect 15380 25936 15425 25976
rect 17155 25936 17164 25976
rect 17204 25936 17300 25976
rect 3916 25768 4292 25808
rect 4492 25724 4532 25936
rect 9667 25852 9676 25892
rect 9716 25852 10100 25892
rect 10060 25808 10100 25852
rect 10540 25808 10580 25936
rect 17260 25892 17300 25936
rect 20140 25892 20180 26104
rect 21510 26084 21600 26104
rect 10627 25852 10636 25892
rect 10676 25852 11980 25892
rect 12020 25852 12029 25892
rect 16963 25852 16972 25892
rect 17012 25852 17021 25892
rect 17260 25852 17740 25892
rect 17780 25852 17789 25892
rect 19363 25852 19372 25892
rect 19412 25852 20180 25892
rect 16972 25808 17012 25852
rect 6019 25768 6028 25808
rect 6068 25768 9004 25808
rect 9044 25768 9053 25808
rect 10051 25768 10060 25808
rect 10100 25768 10109 25808
rect 10540 25768 11308 25808
rect 11348 25768 11357 25808
rect 16972 25768 19796 25808
rect 3628 25684 4532 25724
rect 4919 25684 4928 25724
rect 4968 25684 5010 25724
rect 5050 25684 5092 25724
rect 5132 25684 5174 25724
rect 5214 25684 5256 25724
rect 5296 25684 5305 25724
rect 5356 25684 15436 25724
rect 15476 25684 15485 25724
rect 5356 25640 5396 25684
rect 0 25600 556 25640
rect 596 25600 605 25640
rect 3148 25600 5396 25640
rect 9868 25600 10388 25640
rect 0 25580 90 25600
rect 1459 25432 1468 25472
rect 1508 25432 2092 25472
rect 2132 25432 2141 25472
rect 1769 25348 1804 25388
rect 1844 25348 1900 25388
rect 1940 25348 1949 25388
rect 3148 25379 3188 25600
rect 3331 25516 3340 25556
rect 3380 25516 4300 25556
rect 4340 25516 4349 25556
rect 5203 25516 5212 25556
rect 5252 25516 7852 25556
rect 7892 25516 7901 25556
rect 9091 25516 9100 25556
rect 9140 25516 9772 25556
rect 9812 25516 9821 25556
rect 9868 25472 9908 25600
rect 9955 25516 9964 25556
rect 10004 25516 10013 25556
rect 3689 25432 3772 25472
rect 3812 25432 3820 25472
rect 3860 25432 3869 25472
rect 4147 25432 4156 25472
rect 4196 25432 9908 25472
rect 9964 25388 10004 25516
rect 10348 25472 10388 25600
rect 10531 25516 10540 25556
rect 10580 25516 11116 25556
rect 11156 25516 11165 25556
rect 11299 25516 11308 25556
rect 11348 25516 11404 25556
rect 11444 25516 11479 25556
rect 16195 25516 16204 25556
rect 16244 25516 16724 25556
rect 10348 25432 12980 25472
rect 15907 25432 15916 25472
rect 15956 25432 16244 25472
rect 5347 25348 5356 25388
rect 5396 25348 5405 25388
rect 6604 25379 7276 25388
rect 3148 25330 3188 25339
rect 0 25304 90 25324
rect 5356 25304 5396 25348
rect 6644 25348 7276 25379
rect 7316 25348 7325 25388
rect 7651 25348 7660 25388
rect 7700 25348 7852 25388
rect 7892 25348 7901 25388
rect 8908 25379 9100 25388
rect 6604 25330 6644 25339
rect 8948 25348 9100 25379
rect 9140 25348 9149 25388
rect 9227 25348 9292 25388
rect 9332 25348 9358 25388
rect 9398 25348 9407 25388
rect 9472 25348 9481 25388
rect 9521 25348 9620 25388
rect 9730 25348 9772 25388
rect 9812 25348 9861 25388
rect 9901 25348 9910 25388
rect 9955 25348 9964 25388
rect 10004 25348 10013 25388
rect 10339 25348 10348 25388
rect 10388 25379 10519 25388
rect 10388 25348 10444 25379
rect 8908 25330 8948 25339
rect 9580 25304 9620 25348
rect 10484 25348 10519 25379
rect 10924 25379 11308 25388
rect 10444 25330 10484 25339
rect 10964 25348 11308 25379
rect 11348 25348 11357 25388
rect 11596 25379 12268 25388
rect 10924 25330 10964 25339
rect 11636 25348 12268 25379
rect 12308 25348 12317 25388
rect 12748 25348 12844 25388
rect 12884 25348 12893 25388
rect 11596 25330 11636 25339
rect 0 25264 76 25304
rect 116 25264 125 25304
rect 1097 25264 1228 25304
rect 1268 25264 1277 25304
rect 3523 25264 3532 25304
rect 3572 25264 3628 25304
rect 3668 25264 3703 25304
rect 3907 25264 3916 25304
rect 3956 25264 3965 25304
rect 4579 25264 4588 25304
rect 4628 25264 4637 25304
rect 4867 25264 4876 25304
rect 4916 25264 4972 25304
rect 5012 25264 5047 25304
rect 5203 25264 5212 25304
rect 5252 25264 5396 25304
rect 7049 25264 7180 25304
rect 7220 25264 7229 25304
rect 9580 25264 9964 25304
rect 10004 25264 10013 25304
rect 0 25244 90 25264
rect 3916 25220 3956 25264
rect 643 25180 652 25220
rect 692 25180 3956 25220
rect 4588 25220 4628 25264
rect 12748 25220 12788 25348
rect 12940 25220 12980 25432
rect 16204 25388 16244 25432
rect 16684 25388 16724 25516
rect 17260 25432 18316 25472
rect 18356 25432 18365 25472
rect 18787 25432 18796 25472
rect 18836 25432 19508 25472
rect 14179 25348 14188 25388
rect 14228 25348 14420 25388
rect 14467 25348 14476 25388
rect 14516 25348 14668 25388
rect 14708 25348 14956 25388
rect 14996 25348 15005 25388
rect 15593 25348 15724 25388
rect 15764 25348 15773 25388
rect 16186 25348 16195 25388
rect 16235 25348 16244 25388
rect 16291 25348 16300 25388
rect 16340 25348 16349 25388
rect 16553 25348 16684 25388
rect 16724 25348 16733 25388
rect 17260 25379 17300 25432
rect 13795 25264 13804 25304
rect 13844 25264 13900 25304
rect 13940 25264 13975 25304
rect 14380 25220 14420 25348
rect 15724 25330 15764 25339
rect 16300 25304 16340 25348
rect 17609 25348 17740 25388
rect 17780 25348 17789 25388
rect 18115 25348 18124 25388
rect 18164 25348 18604 25388
rect 18644 25348 18653 25388
rect 19372 25379 19412 25388
rect 17260 25330 17300 25339
rect 17740 25330 17780 25339
rect 19372 25304 19412 25339
rect 16195 25264 16204 25304
rect 16244 25264 16340 25304
rect 16771 25264 16780 25304
rect 16820 25264 16972 25304
rect 17012 25264 17021 25304
rect 18115 25264 18124 25304
rect 18164 25264 19412 25304
rect 19468 25304 19508 25432
rect 19756 25388 19796 25768
rect 20039 25684 20048 25724
rect 20088 25684 20130 25724
rect 20170 25684 20212 25724
rect 20252 25684 20294 25724
rect 20334 25684 20376 25724
rect 20416 25684 20425 25724
rect 21510 25640 21600 25660
rect 20515 25600 20524 25640
rect 20564 25600 21600 25640
rect 21510 25580 21600 25600
rect 20371 25516 20380 25556
rect 20420 25516 21100 25556
rect 21140 25516 21149 25556
rect 19987 25432 19996 25472
rect 20036 25432 21196 25472
rect 21236 25432 21245 25472
rect 19756 25348 20180 25388
rect 20140 25304 20180 25348
rect 19468 25264 19756 25304
rect 19796 25264 19805 25304
rect 20131 25264 20140 25304
rect 20180 25264 20189 25304
rect 20707 25264 20716 25304
rect 20756 25264 20765 25304
rect 16780 25220 16820 25264
rect 20716 25220 20756 25264
rect 4588 25180 5932 25220
rect 5972 25180 5981 25220
rect 6691 25180 6700 25220
rect 6740 25180 6940 25220
rect 6980 25180 6989 25220
rect 12739 25180 12748 25220
rect 12788 25180 12797 25220
rect 12940 25180 16820 25220
rect 17971 25180 17980 25220
rect 18020 25180 20756 25220
rect 21510 25136 21600 25156
rect 4339 25096 4348 25136
rect 4388 25096 5108 25136
rect 6499 25096 6508 25136
rect 6548 25096 6796 25136
rect 6836 25096 6845 25136
rect 9091 25096 9100 25136
rect 9140 25096 11020 25136
rect 11060 25096 11069 25136
rect 13507 25096 13516 25136
rect 13556 25096 13564 25136
rect 13604 25096 13687 25136
rect 14323 25096 14332 25136
rect 14372 25096 14572 25136
rect 14612 25096 14621 25136
rect 19555 25096 19564 25136
rect 19604 25096 19613 25136
rect 20707 25096 20716 25136
rect 20756 25096 21600 25136
rect 5068 25052 5108 25096
rect 3532 25012 4148 25052
rect 5068 25012 5836 25052
rect 5876 25012 5885 25052
rect 12940 25012 13228 25052
rect 13268 25012 13277 25052
rect 0 24968 90 24988
rect 3532 24968 3572 25012
rect 4108 24968 4148 25012
rect 12940 24968 12980 25012
rect 0 24928 3572 24968
rect 3679 24928 3688 24968
rect 3728 24928 3770 24968
rect 3810 24928 3852 24968
rect 3892 24928 3934 24968
rect 3974 24928 4016 24968
rect 4056 24928 4065 24968
rect 4108 24928 6644 24968
rect 6979 24928 6988 24968
rect 7028 24928 12980 24968
rect 16108 24928 17876 24968
rect 18799 24928 18808 24968
rect 18848 24928 18890 24968
rect 18930 24928 18972 24968
rect 19012 24928 19054 24968
rect 19094 24928 19136 24968
rect 19176 24928 19185 24968
rect 0 24908 90 24928
rect 6604 24884 6644 24928
rect 6499 24844 6508 24884
rect 6548 24844 6557 24884
rect 6604 24844 7604 24884
rect 7843 24844 7852 24884
rect 7892 24844 12748 24884
rect 12788 24844 12797 24884
rect 6508 24800 6548 24844
rect 7564 24800 7604 24844
rect 16108 24800 16148 24928
rect 17836 24884 17876 24928
rect 16963 24844 16972 24884
rect 17012 24844 17588 24884
rect 17827 24844 17836 24884
rect 17876 24844 17885 24884
rect 4579 24760 4588 24800
rect 4628 24760 5212 24800
rect 5252 24760 5261 24800
rect 5923 24760 5932 24800
rect 5972 24760 5980 24800
rect 6020 24760 6124 24800
rect 6164 24760 6180 24800
rect 6508 24760 6644 24800
rect 2755 24676 2764 24716
rect 2804 24676 3724 24716
rect 3764 24676 3773 24716
rect 5299 24676 5308 24716
rect 5348 24676 5452 24716
rect 5492 24676 5501 24716
rect 0 24632 90 24652
rect 6604 24632 6644 24760
rect 0 24592 652 24632
rect 692 24592 701 24632
rect 3331 24592 3340 24632
rect 3380 24592 3532 24632
rect 3572 24592 3581 24632
rect 4841 24592 4972 24632
rect 5012 24592 5021 24632
rect 5251 24592 5260 24632
rect 5300 24592 5548 24632
rect 5588 24592 5597 24632
rect 5731 24592 5740 24632
rect 5780 24592 5932 24632
rect 5972 24592 6316 24632
rect 6356 24592 6365 24632
rect 6412 24592 6644 24632
rect 6700 24760 7468 24800
rect 7508 24760 7517 24800
rect 7564 24760 9236 24800
rect 9379 24760 9388 24800
rect 9428 24760 9724 24800
rect 9764 24760 9773 24800
rect 11177 24760 11308 24800
rect 11348 24760 11357 24800
rect 15187 24760 15196 24800
rect 15236 24760 16148 24800
rect 16195 24760 16204 24800
rect 16244 24760 17156 24800
rect 0 24572 90 24592
rect 2572 24548 2612 24557
rect 4108 24548 4148 24557
rect 6412 24548 6452 24592
rect 6700 24548 6740 24760
rect 8035 24676 8044 24716
rect 8084 24676 8756 24716
rect 8873 24676 8956 24716
rect 8996 24676 9004 24716
rect 9044 24676 9053 24716
rect 8716 24632 8756 24676
rect 9196 24632 9236 24760
rect 9331 24676 9340 24716
rect 9380 24676 14476 24716
rect 14516 24676 14525 24716
rect 14755 24676 14764 24716
rect 14804 24676 15340 24716
rect 15380 24676 15389 24716
rect 16771 24676 16780 24716
rect 16820 24676 16829 24716
rect 6857 24592 6892 24632
rect 6932 24592 6988 24632
rect 7028 24592 7037 24632
rect 8170 24592 8179 24632
rect 8219 24592 8332 24632
rect 8372 24592 8381 24632
rect 8441 24592 8524 24632
rect 8564 24592 8572 24632
rect 8612 24592 8621 24632
rect 8707 24592 8716 24632
rect 8756 24592 8765 24632
rect 8812 24592 9100 24632
rect 9140 24592 9149 24632
rect 9196 24592 9484 24632
rect 9524 24592 9533 24632
rect 14825 24592 14956 24632
rect 14996 24592 15005 24632
rect 15427 24592 15436 24632
rect 15476 24592 16628 24632
rect 7468 24548 7508 24557
rect 1027 24508 1036 24548
rect 1076 24508 1324 24548
rect 1364 24508 1373 24548
rect 2441 24508 2572 24548
rect 2612 24508 2621 24548
rect 2851 24508 2860 24548
rect 2900 24508 3043 24548
rect 3083 24508 3092 24548
rect 3139 24508 3148 24548
rect 3188 24508 3197 24548
rect 3497 24508 3628 24548
rect 3668 24508 3677 24548
rect 4291 24508 4300 24548
rect 4340 24508 4596 24548
rect 4636 24508 4645 24548
rect 6394 24508 6403 24548
rect 6443 24508 6452 24548
rect 6499 24508 6508 24548
rect 6548 24508 6740 24548
rect 6828 24508 6892 24548
rect 6932 24508 6988 24548
rect 7028 24508 7084 24548
rect 7124 24508 7133 24548
rect 7337 24508 7468 24548
rect 7508 24508 7517 24548
rect 7843 24508 7852 24548
rect 7892 24508 7956 24548
rect 7996 24508 8023 24548
rect 2572 24499 2612 24508
rect 3148 24464 3188 24508
rect 3043 24424 3052 24464
rect 3092 24424 3188 24464
rect 4108 24464 4148 24508
rect 6508 24464 6548 24508
rect 7468 24499 7508 24508
rect 4108 24424 4876 24464
rect 4916 24424 4925 24464
rect 6307 24424 6316 24464
rect 6356 24424 6548 24464
rect 8716 24380 8756 24592
rect 8812 24464 8852 24592
rect 11116 24548 11156 24557
rect 12748 24548 12788 24557
rect 14572 24548 14612 24557
rect 16588 24548 16628 24592
rect 9859 24508 9868 24548
rect 9908 24508 10636 24548
rect 10676 24508 10685 24548
rect 11011 24508 11020 24548
rect 11060 24508 11116 24548
rect 11156 24508 11191 24548
rect 11465 24508 11500 24548
rect 11540 24508 11596 24548
rect 11636 24508 11645 24548
rect 11875 24508 11884 24548
rect 11924 24508 12748 24548
rect 13219 24508 13228 24548
rect 13268 24508 13324 24548
rect 13364 24508 13399 24548
rect 13507 24508 13516 24548
rect 13556 24508 14572 24548
rect 14659 24508 14668 24548
rect 14708 24508 15340 24548
rect 15380 24508 15628 24548
rect 15668 24508 15677 24548
rect 16780 24548 16820 24676
rect 17116 24632 17156 24760
rect 17548 24716 17588 24844
rect 19145 24760 19228 24800
rect 19268 24760 19276 24800
rect 19316 24760 19325 24800
rect 19564 24716 19604 25096
rect 21510 25076 21600 25096
rect 20131 24844 20140 24884
rect 20180 24844 21100 24884
rect 21140 24844 21149 24884
rect 19843 24760 19852 24800
rect 19892 24760 19996 24800
rect 20036 24760 20045 24800
rect 20371 24760 20380 24800
rect 20420 24760 21004 24800
rect 21044 24760 21053 24800
rect 17548 24676 17684 24716
rect 17116 24592 17204 24632
rect 17251 24592 17260 24632
rect 17300 24592 17548 24632
rect 17588 24592 17597 24632
rect 17164 24548 17204 24592
rect 17644 24548 17684 24676
rect 18604 24676 19604 24716
rect 19756 24676 21388 24716
rect 21428 24676 21437 24716
rect 18604 24581 18644 24676
rect 19756 24632 19796 24676
rect 21510 24632 21600 24652
rect 18979 24592 18988 24632
rect 19028 24592 19124 24632
rect 19241 24592 19276 24632
rect 19316 24592 19372 24632
rect 19412 24592 19421 24632
rect 19603 24592 19612 24632
rect 19652 24592 19700 24632
rect 19747 24592 19756 24632
rect 19796 24592 19805 24632
rect 20131 24592 20140 24632
rect 20180 24592 20189 24632
rect 21091 24592 21100 24632
rect 21140 24592 21600 24632
rect 18124 24548 18164 24557
rect 16780 24508 17059 24548
rect 17099 24508 17108 24548
rect 17155 24508 17164 24548
rect 17204 24508 17213 24548
rect 17635 24508 17644 24548
rect 17684 24508 17693 24548
rect 18164 24508 18316 24548
rect 18356 24508 18365 24548
rect 18604 24532 18644 24541
rect 19084 24548 19124 24592
rect 19660 24548 19700 24592
rect 20140 24548 20180 24592
rect 21510 24572 21600 24592
rect 19084 24508 19468 24548
rect 19508 24508 19517 24548
rect 19660 24508 19948 24548
rect 19988 24508 19997 24548
rect 20140 24508 21388 24548
rect 21428 24508 21437 24548
rect 11116 24499 11156 24508
rect 12748 24499 12788 24508
rect 14572 24499 14612 24508
rect 16588 24464 16628 24508
rect 18124 24499 18164 24508
rect 8803 24424 8812 24464
rect 8852 24424 8861 24464
rect 16588 24424 18028 24464
rect 18068 24424 18077 24464
rect 19843 24424 19852 24464
rect 19892 24424 20812 24464
rect 20852 24424 20861 24464
rect 4291 24340 4300 24380
rect 4340 24340 4780 24380
rect 4820 24340 4829 24380
rect 8716 24340 9388 24380
rect 9428 24340 9437 24380
rect 12931 24340 12940 24380
rect 12980 24340 12989 24380
rect 18665 24340 18796 24380
rect 18836 24340 18845 24380
rect 0 24296 90 24316
rect 0 24256 10100 24296
rect 0 24236 90 24256
rect 4919 24172 4928 24212
rect 4968 24172 5010 24212
rect 5050 24172 5092 24212
rect 5132 24172 5174 24212
rect 5214 24172 5256 24212
rect 5296 24172 5305 24212
rect 1603 24088 1612 24128
rect 1652 24088 4628 24128
rect 8035 24088 8044 24128
rect 8084 24088 9764 24128
rect 0 23960 90 23980
rect 4588 23960 4628 24088
rect 9724 24044 9764 24088
rect 4771 24004 4780 24044
rect 4820 24004 7180 24044
rect 7220 24004 7229 24044
rect 7459 24004 7468 24044
rect 7508 24004 7852 24044
rect 7892 24004 7901 24044
rect 9161 24004 9292 24044
rect 9332 24004 9341 24044
rect 9715 24004 9724 24044
rect 9764 24004 9773 24044
rect 0 23920 1036 23960
rect 1076 23920 1085 23960
rect 2755 23920 2764 23960
rect 2804 23920 3092 23960
rect 3715 23920 3724 23960
rect 3764 23920 4244 23960
rect 4588 23920 6796 23960
rect 6836 23920 6845 23960
rect 8611 23920 8620 23960
rect 8660 23920 9820 23960
rect 9860 23920 9869 23960
rect 0 23900 90 23920
rect 3052 23876 3092 23920
rect 4204 23876 4244 23920
rect 931 23836 940 23876
rect 980 23836 1324 23876
rect 1364 23836 1373 23876
rect 2441 23836 2572 23876
rect 2612 23836 2621 23876
rect 3034 23836 3043 23876
rect 3083 23836 3092 23876
rect 3139 23836 3148 23876
rect 3188 23836 3197 23876
rect 3523 23836 3532 23876
rect 3572 23836 4012 23876
rect 4052 23836 4061 23876
rect 4108 23867 4148 23876
rect 2572 23818 2612 23827
rect 3148 23792 3188 23836
rect 4204 23867 4628 23876
rect 4204 23836 4588 23867
rect 4108 23792 4148 23827
rect 4675 23836 4684 23876
rect 4724 23836 5396 23876
rect 5827 23836 5836 23876
rect 5876 23836 6028 23876
rect 6068 23836 6988 23876
rect 7028 23836 7037 23876
rect 7145 23836 7276 23876
rect 7316 23836 7325 23876
rect 7843 23836 7852 23876
rect 7892 23836 8852 23876
rect 8969 23836 9100 23876
rect 9140 23836 9149 23876
rect 4588 23818 4628 23827
rect 5356 23792 5396 23836
rect 7276 23818 7316 23827
rect 3043 23752 3052 23792
rect 3092 23752 3188 23792
rect 3497 23752 3628 23792
rect 3668 23752 3677 23792
rect 4108 23752 4340 23792
rect 4841 23752 4972 23792
rect 5012 23752 5021 23792
rect 5347 23752 5356 23792
rect 5396 23752 5452 23792
rect 5492 23752 5556 23792
rect 5923 23752 5932 23792
rect 5972 23752 5981 23792
rect 0 23624 90 23644
rect 4300 23624 4340 23752
rect 5932 23708 5972 23752
rect 5068 23668 5972 23708
rect 8812 23708 8852 23836
rect 9100 23818 9140 23827
rect 10060 23792 10100 24256
rect 12940 24044 12980 24340
rect 18979 24256 18988 24296
rect 19028 24256 19756 24296
rect 19796 24256 19805 24296
rect 17740 24172 19372 24212
rect 19412 24172 19421 24212
rect 20039 24172 20048 24212
rect 20088 24172 20130 24212
rect 20170 24172 20212 24212
rect 20252 24172 20294 24212
rect 20334 24172 20376 24212
rect 20416 24172 20425 24212
rect 17740 24044 17780 24172
rect 21510 24128 21600 24148
rect 17827 24088 17836 24128
rect 17876 24088 21600 24128
rect 21510 24068 21600 24088
rect 12940 24004 15188 24044
rect 15593 24004 15724 24044
rect 15764 24004 15773 24044
rect 16579 24004 16588 24044
rect 16628 24004 16732 24044
rect 16772 24004 16781 24044
rect 17491 24004 17500 24044
rect 17540 24004 17780 24044
rect 19084 24004 19372 24044
rect 19412 24004 19421 24044
rect 19546 24004 19555 24044
rect 19595 24004 20180 24044
rect 11971 23920 11980 23960
rect 12020 23920 14036 23960
rect 13996 23876 14036 23920
rect 15148 23876 15188 24004
rect 17827 23920 17836 23960
rect 17876 23920 18700 23960
rect 18740 23920 18749 23960
rect 18835 23920 18844 23960
rect 18884 23920 18988 23960
rect 19028 23920 19037 23960
rect 19084 23876 19124 24004
rect 20140 23960 20180 24004
rect 19258 23920 19267 23960
rect 19307 23920 19767 23960
rect 19807 23920 19816 23960
rect 20131 23920 20140 23960
rect 20180 23920 21196 23960
rect 21236 23920 21245 23960
rect 10435 23836 10444 23876
rect 10484 23836 10540 23876
rect 10580 23836 10615 23876
rect 11753 23867 11884 23876
rect 11753 23836 11788 23867
rect 11828 23836 11884 23867
rect 11924 23836 11933 23876
rect 11980 23836 12172 23876
rect 12212 23836 12652 23876
rect 12692 23836 12701 23876
rect 13385 23867 13516 23876
rect 13385 23836 13420 23867
rect 11788 23818 11828 23827
rect 11980 23792 12020 23836
rect 13460 23836 13516 23867
rect 13556 23836 13565 23876
rect 13978 23836 13987 23876
rect 14027 23836 14036 23876
rect 14083 23836 14092 23876
rect 14132 23836 14188 23876
rect 14228 23836 14263 23876
rect 14345 23836 14476 23876
rect 14516 23836 14525 23876
rect 14659 23836 14668 23876
rect 14708 23867 15092 23876
rect 14708 23836 15052 23867
rect 13420 23818 13460 23827
rect 15148 23867 15572 23876
rect 15148 23836 15532 23867
rect 15052 23818 15092 23827
rect 15532 23818 15572 23827
rect 17260 23836 18796 23876
rect 18836 23836 18845 23876
rect 18946 23836 18955 23876
rect 18995 23836 19124 23876
rect 19169 23836 19178 23876
rect 19218 23836 19227 23876
rect 19450 23836 19459 23876
rect 19499 23836 19660 23876
rect 19700 23836 19709 23876
rect 19925 23836 19934 23876
rect 19974 23836 19983 23876
rect 20236 23867 20524 23876
rect 17260 23792 17300 23836
rect 19178 23792 19218 23836
rect 19934 23792 19974 23836
rect 20276 23836 20524 23867
rect 20564 23836 20573 23876
rect 20236 23818 20276 23827
rect 9379 23752 9388 23792
rect 9428 23752 9484 23792
rect 9524 23752 9559 23792
rect 10051 23752 10060 23792
rect 10100 23752 10109 23792
rect 11971 23752 11980 23792
rect 12020 23752 12029 23792
rect 13987 23752 13996 23792
rect 14036 23752 14572 23792
rect 14612 23752 14956 23792
rect 14996 23752 15005 23792
rect 15715 23752 15724 23792
rect 15764 23752 16108 23792
rect 16148 23752 16157 23792
rect 16361 23752 16396 23792
rect 16436 23752 16492 23792
rect 16532 23752 16541 23792
rect 16867 23752 16876 23792
rect 16916 23752 16925 23792
rect 17251 23752 17260 23792
rect 17300 23752 17309 23792
rect 17705 23752 17836 23792
rect 17876 23752 17885 23792
rect 17971 23752 17980 23792
rect 18020 23752 18028 23792
rect 18068 23752 18151 23792
rect 18211 23752 18220 23792
rect 18260 23752 18269 23792
rect 18473 23752 18604 23792
rect 18644 23752 18653 23792
rect 18700 23752 19075 23792
rect 19115 23752 19124 23792
rect 19178 23752 19372 23792
rect 19412 23752 19974 23792
rect 8812 23668 12172 23708
rect 12212 23668 12221 23708
rect 5068 23624 5108 23668
rect 0 23584 3724 23624
rect 3764 23584 3773 23624
rect 3907 23584 3916 23624
rect 3956 23584 3965 23624
rect 4300 23584 5108 23624
rect 5203 23584 5212 23624
rect 5252 23584 5261 23624
rect 5587 23584 5596 23624
rect 5636 23584 7084 23624
rect 7124 23584 7133 23624
rect 7939 23584 7948 23624
rect 7988 23584 10828 23624
rect 10868 23584 10877 23624
rect 13481 23584 13612 23624
rect 13652 23584 13661 23624
rect 15859 23584 15868 23624
rect 15908 23584 16012 23624
rect 16052 23584 16061 23624
rect 0 23564 90 23584
rect 3916 23540 3956 23584
rect 5212 23540 5252 23584
rect 3916 23500 4163 23540
rect 5212 23500 14284 23540
rect 14324 23500 14333 23540
rect 4123 23456 4163 23500
rect 16876 23456 16916 23752
rect 18220 23708 18260 23752
rect 18700 23708 18740 23752
rect 18115 23668 18124 23708
rect 18164 23668 18260 23708
rect 18691 23668 18700 23708
rect 18740 23668 18749 23708
rect 21510 23624 21600 23644
rect 17107 23584 17116 23624
rect 17156 23584 17260 23624
rect 17300 23584 17309 23624
rect 17587 23584 17596 23624
rect 17636 23584 17836 23624
rect 17876 23584 17885 23624
rect 17932 23584 18220 23624
rect 18260 23584 18269 23624
rect 19625 23584 19756 23624
rect 19796 23584 19805 23624
rect 19930 23584 19939 23624
rect 19988 23584 20119 23624
rect 20803 23584 20812 23624
rect 20852 23584 21600 23624
rect 3679 23416 3688 23456
rect 3728 23416 3770 23456
rect 3810 23416 3852 23456
rect 3892 23416 3934 23456
rect 3974 23416 4016 23456
rect 4056 23416 4065 23456
rect 4123 23416 6796 23456
rect 6836 23416 6845 23456
rect 12940 23416 16916 23456
rect 1603 23332 1612 23372
rect 1652 23332 1661 23372
rect 2947 23332 2956 23372
rect 2996 23332 3005 23372
rect 0 23288 90 23308
rect 0 23228 116 23288
rect 76 23204 116 23228
rect 1612 23204 1652 23332
rect 2956 23288 2996 23332
rect 4123 23288 4163 23416
rect 4675 23332 4684 23372
rect 4724 23332 10676 23372
rect 2956 23248 3284 23288
rect 3331 23248 3340 23288
rect 3380 23248 3628 23288
rect 3668 23248 3677 23288
rect 4123 23248 4156 23288
rect 4196 23248 4205 23288
rect 4396 23248 5740 23288
rect 5780 23248 5789 23288
rect 7084 23248 10060 23288
rect 10100 23248 10109 23288
rect 10339 23248 10348 23288
rect 10388 23248 10483 23288
rect 10523 23248 10532 23288
rect 76 23164 1364 23204
rect 1459 23164 1468 23204
rect 1508 23164 1652 23204
rect 2860 23164 3148 23204
rect 3188 23164 3197 23204
rect 1324 23120 1364 23164
rect 2860 23120 2900 23164
rect 739 23080 748 23120
rect 788 23080 1228 23120
rect 1268 23080 1277 23120
rect 1324 23080 2900 23120
rect 3244 23120 3284 23248
rect 4396 23204 4436 23248
rect 7084 23204 7124 23248
rect 3706 23164 3715 23204
rect 3755 23164 4436 23204
rect 4531 23164 4540 23204
rect 4580 23164 7124 23204
rect 7180 23164 9236 23204
rect 7180 23120 7220 23164
rect 9196 23120 9236 23164
rect 10636 23120 10676 23332
rect 12940 23288 12980 23416
rect 17932 23288 17972 23584
rect 21510 23564 21600 23584
rect 18799 23416 18808 23456
rect 18848 23416 18890 23456
rect 18930 23416 18972 23456
rect 19012 23416 19054 23456
rect 19094 23416 19136 23456
rect 19176 23416 19185 23456
rect 10819 23248 10828 23288
rect 10868 23248 10972 23288
rect 11012 23248 11021 23288
rect 11635 23248 11644 23288
rect 11684 23248 11884 23288
rect 11924 23248 12980 23288
rect 15562 23248 15571 23288
rect 15611 23248 15724 23288
rect 15764 23248 15773 23288
rect 16579 23248 16588 23288
rect 16628 23248 16780 23288
rect 16820 23248 16829 23288
rect 17674 23248 17683 23288
rect 17723 23248 17972 23288
rect 18028 23332 20044 23372
rect 20084 23332 20093 23372
rect 10867 23164 10876 23204
rect 10916 23164 13036 23204
rect 13076 23164 13085 23204
rect 14284 23164 14996 23204
rect 14284 23120 14324 23164
rect 14956 23120 14996 23164
rect 18028 23120 18068 23332
rect 18451 23248 18460 23288
rect 18500 23248 19564 23288
rect 19604 23248 19613 23288
rect 19171 23164 19180 23204
rect 19220 23164 20188 23204
rect 20228 23164 20237 23204
rect 21510 23120 21600 23140
rect 3244 23080 3340 23120
rect 3380 23080 3389 23120
rect 3785 23080 3916 23120
rect 3956 23080 3965 23120
rect 4169 23080 4300 23120
rect 4340 23080 4349 23120
rect 7171 23080 7180 23120
rect 7220 23080 7229 23120
rect 7756 23080 7852 23120
rect 7892 23080 7901 23120
rect 7948 23080 8428 23120
rect 8468 23080 8852 23120
rect 8995 23080 9004 23120
rect 9044 23080 9053 23120
rect 9187 23080 9196 23120
rect 9236 23080 9388 23120
rect 9428 23080 9437 23120
rect 9667 23080 9676 23120
rect 9716 23080 9725 23120
rect 10627 23080 10636 23120
rect 10676 23080 10685 23120
rect 11203 23080 11212 23120
rect 11252 23080 11261 23120
rect 11875 23080 11884 23120
rect 11924 23080 12268 23120
rect 12308 23080 12317 23120
rect 14153 23080 14284 23120
rect 14324 23080 14333 23120
rect 14956 23080 16292 23120
rect 16387 23080 16396 23120
rect 16436 23080 16684 23120
rect 16724 23080 16788 23120
rect 17779 23080 17788 23120
rect 17828 23080 17836 23120
rect 17876 23080 17959 23120
rect 18019 23080 18028 23120
rect 18068 23080 18077 23120
rect 18211 23080 18220 23120
rect 18260 23080 18796 23120
rect 18836 23080 18845 23120
rect 21091 23080 21100 23120
rect 21140 23080 21600 23120
rect 3148 23036 3188 23045
rect 5932 23036 5972 23045
rect 7756 23036 7796 23080
rect 1891 22996 1900 23036
rect 1940 22996 1949 23036
rect 2371 22996 2380 23036
rect 2420 22996 3148 23036
rect 3401 22996 3532 23036
rect 3572 22996 3581 23036
rect 3706 22996 3715 23036
rect 3755 22996 3764 23036
rect 4675 22996 4684 23036
rect 4724 22996 4733 23036
rect 5897 22996 5932 23036
rect 5972 22996 6028 23036
rect 6068 22996 6077 23036
rect 6124 22996 6691 23036
rect 6731 22996 6740 23036
rect 6787 22996 6796 23036
rect 6836 22996 6845 23036
rect 7241 22996 7276 23036
rect 7316 22996 7372 23036
rect 7412 22996 7421 23036
rect 0 22952 90 22972
rect 0 22912 1132 22952
rect 1172 22912 1181 22952
rect 0 22892 90 22912
rect 1900 22868 1940 22996
rect 3148 22987 3188 22996
rect 3724 22952 3764 22996
rect 4684 22952 4724 22996
rect 5932 22987 5972 22996
rect 6124 22952 6164 22996
rect 3235 22912 3244 22952
rect 3284 22912 3764 22952
rect 4003 22912 4012 22952
rect 4052 22912 4300 22952
rect 4340 22912 4724 22952
rect 6115 22912 6124 22952
rect 6164 22912 6173 22952
rect 1900 22828 3532 22868
rect 3572 22828 3581 22868
rect 3724 22784 3764 22912
rect 6796 22868 6836 22996
rect 7756 22987 7796 22996
rect 7948 22868 7988 23080
rect 8812 23036 8852 23080
rect 9004 23036 9044 23080
rect 9676 23036 9716 23080
rect 9772 23036 9812 23045
rect 6796 22828 7564 22868
rect 7604 22828 7988 22868
rect 8044 22996 8244 23036
rect 8284 22996 8293 23036
rect 8668 22996 8707 23036
rect 8747 22996 8756 23036
rect 8803 22996 8812 23036
rect 8852 22996 8861 23036
rect 9004 22996 9292 23036
rect 9332 22996 9341 23036
rect 9676 22996 9772 23036
rect 10282 22996 10291 23036
rect 10331 22996 10348 23036
rect 10388 22996 10471 23036
rect 3724 22744 4204 22784
rect 4244 22744 4253 22784
rect 4919 22660 4928 22700
rect 4968 22660 5010 22700
rect 5050 22660 5092 22700
rect 5132 22660 5174 22700
rect 5214 22660 5256 22700
rect 5296 22660 5305 22700
rect 0 22616 90 22636
rect 0 22576 5836 22616
rect 5876 22576 5885 22616
rect 0 22556 90 22576
rect 8044 22532 8084 22996
rect 8668 22952 8708 22996
rect 9772 22987 9812 22996
rect 8668 22912 9004 22952
rect 9044 22912 9053 22952
rect 11212 22868 11252 23080
rect 13324 23036 13364 23045
rect 14860 23036 14900 23045
rect 16252 23036 16292 23080
rect 12067 22996 12076 23036
rect 12116 22996 12308 23036
rect 12268 22952 12308 22996
rect 12940 22996 13324 23036
rect 13603 22996 13612 23036
rect 13652 22996 13795 23036
rect 13835 22996 13844 23036
rect 13891 22996 13900 23036
rect 13940 22996 14188 23036
rect 14228 22996 14237 23036
rect 14371 22996 14380 23036
rect 14420 22996 14476 23036
rect 14516 22996 14580 23036
rect 14659 22996 14668 23036
rect 14708 22996 14860 23036
rect 15331 22996 15340 23036
rect 15388 22996 15511 23036
rect 15898 22996 15907 23036
rect 15947 22996 15956 23036
rect 16003 22996 16012 23036
rect 16052 22996 16108 23036
rect 16148 22996 16183 23036
rect 16252 22996 16492 23036
rect 16532 22996 16541 23036
rect 12259 22912 12268 22952
rect 12308 22912 12317 22952
rect 12940 22868 12980 22996
rect 13324 22987 13364 22996
rect 14380 22868 14420 22996
rect 14860 22987 14900 22996
rect 8323 22828 8332 22868
rect 8372 22828 8428 22868
rect 8468 22828 8503 22868
rect 9955 22828 9964 22868
rect 10004 22828 11252 22868
rect 12835 22828 12844 22868
rect 12884 22828 12980 22868
rect 13507 22828 13516 22868
rect 13556 22828 13900 22868
rect 13940 22828 13949 22868
rect 14380 22828 15340 22868
rect 15380 22828 15389 22868
rect 11491 22744 11500 22784
rect 11540 22744 15052 22784
rect 15092 22744 15101 22784
rect 12940 22660 15860 22700
rect 12940 22616 12980 22660
rect 8323 22576 8332 22616
rect 8372 22576 12980 22616
rect 3427 22492 3436 22532
rect 3476 22492 3764 22532
rect 5321 22492 5356 22532
rect 5396 22492 5452 22532
rect 5492 22492 5501 22532
rect 5779 22492 5788 22532
rect 5828 22492 6412 22532
rect 6452 22492 6461 22532
rect 8035 22492 8044 22532
rect 8084 22492 8093 22532
rect 10339 22492 10348 22532
rect 10388 22492 10828 22532
rect 10868 22492 10877 22532
rect 13891 22492 13900 22532
rect 13940 22492 14516 22532
rect 14650 22492 14659 22532
rect 14708 22492 14839 22532
rect 3724 22448 3764 22492
rect 14476 22448 14516 22492
rect 3331 22408 3340 22448
rect 3380 22408 3668 22448
rect 3724 22408 5492 22448
rect 5539 22408 5548 22448
rect 5588 22408 6644 22448
rect 7939 22408 7948 22448
rect 7988 22408 8332 22448
rect 8372 22408 8381 22448
rect 8611 22408 8620 22448
rect 8660 22408 8672 22448
rect 8986 22408 8995 22448
rect 9035 22408 12940 22448
rect 12980 22408 12989 22448
rect 13786 22408 13795 22448
rect 13835 22408 14228 22448
rect 3628 22364 3668 22408
rect 1769 22324 1900 22364
rect 1940 22324 1949 22364
rect 3148 22355 3436 22364
rect 3188 22324 3436 22355
rect 3476 22324 3485 22364
rect 3610 22324 3619 22364
rect 3659 22324 3668 22364
rect 3715 22324 3724 22364
rect 3764 22324 3773 22364
rect 3977 22324 4108 22364
rect 4148 22324 4157 22364
rect 4579 22324 4588 22364
rect 4628 22355 4759 22364
rect 4628 22324 4684 22355
rect 3148 22306 3188 22315
rect 0 22280 90 22300
rect 0 22240 172 22280
rect 212 22240 221 22280
rect 835 22240 844 22280
rect 884 22240 1228 22280
rect 1268 22240 1277 22280
rect 0 22220 90 22240
rect 3724 22196 3764 22324
rect 4724 22324 4759 22355
rect 5164 22355 5356 22364
rect 4684 22306 4724 22315
rect 5204 22324 5356 22355
rect 5396 22324 5405 22364
rect 5164 22306 5204 22315
rect 5452 22280 5492 22408
rect 6604 22364 6644 22408
rect 8632 22364 8672 22408
rect 14188 22364 14228 22408
rect 14458 22439 14516 22448
rect 14458 22399 14467 22439
rect 14507 22399 14516 22439
rect 15820 22448 15860 22660
rect 15916 22532 15956 22996
rect 16588 22952 16628 23080
rect 21510 23060 21600 23080
rect 16972 23036 17012 23045
rect 19852 23036 19892 23045
rect 16812 22996 16876 23036
rect 16916 22996 16972 23036
rect 17012 22996 17260 23036
rect 17300 22996 17309 23036
rect 17482 22996 17491 23036
rect 17531 22996 18028 23036
rect 18068 22996 18077 23036
rect 18595 22996 18604 23036
rect 18644 22996 18892 23036
rect 18932 22996 18941 23036
rect 19721 22996 19852 23036
rect 19892 22996 19901 23036
rect 20323 22996 20332 23036
rect 20372 22996 20381 23036
rect 16972 22987 17012 22996
rect 19852 22987 19892 22996
rect 16483 22912 16492 22952
rect 16532 22912 16628 22952
rect 19555 22828 19564 22868
rect 19604 22828 20044 22868
rect 20084 22828 20093 22868
rect 20332 22784 20372 22996
rect 19843 22744 19852 22784
rect 19892 22744 20372 22784
rect 19276 22660 19796 22700
rect 20039 22660 20048 22700
rect 20088 22660 20130 22700
rect 20170 22660 20212 22700
rect 20252 22660 20294 22700
rect 20334 22660 20376 22700
rect 20416 22660 20425 22700
rect 18508 22576 18892 22616
rect 18932 22576 18941 22616
rect 15916 22492 16492 22532
rect 16532 22492 16541 22532
rect 18019 22492 18028 22532
rect 18068 22492 18124 22532
rect 18164 22492 18199 22532
rect 18508 22448 18548 22576
rect 19276 22532 19316 22660
rect 19756 22616 19796 22660
rect 21510 22616 21600 22636
rect 19756 22576 20180 22616
rect 20995 22576 21004 22616
rect 21044 22576 21600 22616
rect 20140 22532 20180 22576
rect 21510 22556 21600 22576
rect 18691 22492 18700 22532
rect 18740 22492 18787 22532
rect 18827 22492 18871 22532
rect 19258 22492 19267 22532
rect 19307 22492 19316 22532
rect 19738 22492 19747 22532
rect 19787 22492 19852 22532
rect 19892 22492 19927 22532
rect 20131 22492 20140 22532
rect 20180 22492 20189 22532
rect 15820 22408 18548 22448
rect 18604 22408 19564 22448
rect 19604 22408 19613 22448
rect 19939 22408 19948 22448
rect 19988 22408 20276 22448
rect 14458 22398 14516 22399
rect 18604 22364 18644 22408
rect 19564 22364 19604 22408
rect 6028 22355 6068 22364
rect 6250 22355 6412 22364
rect 6028 22280 6068 22315
rect 6118 22304 6127 22344
rect 6167 22304 6176 22344
rect 6250 22315 6259 22355
rect 6299 22324 6412 22355
rect 6452 22324 6461 22364
rect 6595 22324 6604 22364
rect 6644 22324 6653 22364
rect 7459 22324 7468 22364
rect 7508 22355 8044 22364
rect 7508 22324 7852 22355
rect 6299 22315 6308 22324
rect 6250 22314 6308 22315
rect 7892 22324 8044 22355
rect 8084 22324 8093 22364
rect 8218 22324 8227 22364
rect 8267 22324 8276 22364
rect 8323 22324 8332 22364
rect 8372 22324 8535 22364
rect 8575 22324 8584 22364
rect 8632 22324 8663 22364
rect 8703 22324 8712 22364
rect 8899 22324 8908 22364
rect 8948 22324 8957 22364
rect 9091 22324 9100 22364
rect 9140 22324 9388 22364
rect 9428 22324 9437 22364
rect 10636 22355 10676 22364
rect 7892 22321 7896 22324
rect 7852 22306 7892 22315
rect 4195 22240 4204 22280
rect 4244 22240 4396 22280
rect 4436 22240 4445 22280
rect 5452 22240 5548 22280
rect 5588 22240 5597 22280
rect 5981 22240 6028 22280
rect 6068 22240 6077 22280
rect 6127 22196 6167 22304
rect 8236 22280 8276 22324
rect 8236 22240 8428 22280
rect 8468 22240 8477 22280
rect 8681 22240 8716 22280
rect 8756 22240 8803 22280
rect 8843 22240 8861 22280
rect 8908 22196 8948 22324
rect 11491 22324 11500 22364
rect 11540 22324 11692 22364
rect 11732 22324 11741 22364
rect 12780 22324 12844 22364
rect 12884 22355 12980 22364
rect 12884 22324 12940 22355
rect 10636 22196 10676 22315
rect 13123 22324 13132 22364
rect 13172 22324 13708 22364
rect 13748 22324 13757 22364
rect 13882 22324 13891 22364
rect 13931 22324 13940 22364
rect 13987 22324 13996 22364
rect 14036 22324 14083 22364
rect 14170 22324 14179 22364
rect 14219 22324 14228 22364
rect 14284 22355 14324 22364
rect 11011 22240 11020 22280
rect 11060 22240 12076 22280
rect 12116 22240 12125 22280
rect 12940 22196 12980 22315
rect 13900 22280 13940 22324
rect 13996 22280 14036 22324
rect 14562 22324 14571 22364
rect 14611 22324 14620 22364
rect 14284 22280 14324 22315
rect 14572 22280 14612 22324
rect 14668 22313 14689 22353
rect 14729 22313 14738 22353
rect 14921 22324 15052 22364
rect 15092 22324 15101 22364
rect 16300 22355 16340 22364
rect 16553 22324 16684 22364
rect 16724 22324 16876 22364
rect 16916 22324 16925 22364
rect 17827 22324 17836 22364
rect 17876 22355 18007 22364
rect 17876 22324 17932 22355
rect 13132 22240 13940 22280
rect 13987 22240 13996 22280
rect 14036 22240 14045 22280
rect 14284 22240 14380 22280
rect 14420 22240 14429 22280
rect 14533 22240 14572 22280
rect 14612 22240 14621 22280
rect 13132 22196 13172 22240
rect 13900 22196 13940 22240
rect 14668 22196 14708 22313
rect 16300 22280 16340 22315
rect 17836 22280 17876 22324
rect 17972 22324 18007 22355
rect 18466 22324 18475 22364
rect 18515 22324 18644 22364
rect 18691 22324 18700 22364
rect 18740 22324 18836 22364
rect 18883 22324 18892 22364
rect 18932 22324 18935 22364
rect 18975 22324 19063 22364
rect 19171 22324 19180 22364
rect 19220 22324 19351 22364
rect 19546 22324 19555 22364
rect 19595 22324 19604 22364
rect 19651 22324 19660 22364
rect 19700 22324 19709 22364
rect 19843 22324 19852 22364
rect 19892 22324 19934 22364
rect 19974 22324 20023 22364
rect 20236 22355 20276 22408
rect 17932 22306 17972 22315
rect 16300 22240 17876 22280
rect 18499 22240 18508 22280
rect 18548 22240 18595 22280
rect 18635 22240 18679 22280
rect 18796 22196 18836 22324
rect 19411 22282 19420 22322
rect 19460 22282 19469 22322
rect 18892 22240 19075 22280
rect 19115 22240 19124 22280
rect 3043 22156 3052 22196
rect 3092 22156 3764 22196
rect 3811 22156 3820 22196
rect 3860 22156 4588 22196
rect 4628 22156 4637 22196
rect 5923 22156 5932 22196
rect 5972 22156 6167 22196
rect 6403 22156 6412 22196
rect 6452 22156 8948 22196
rect 10147 22156 10156 22196
rect 10196 22156 11308 22196
rect 11348 22156 12980 22196
rect 13123 22156 13132 22196
rect 13172 22156 13181 22196
rect 13891 22156 13900 22196
rect 13940 22156 14708 22196
rect 17251 22156 17260 22196
rect 17300 22156 18028 22196
rect 18068 22156 18077 22196
rect 18787 22156 18796 22196
rect 18836 22156 18845 22196
rect 18892 22112 18932 22240
rect 19415 22196 19455 22282
rect 19660 22280 19700 22324
rect 20236 22306 20276 22315
rect 19660 22240 19948 22280
rect 19988 22240 20180 22280
rect 20140 22196 20180 22240
rect 19075 22156 19084 22196
rect 19124 22156 19852 22196
rect 19892 22156 19901 22196
rect 20140 22156 20236 22196
rect 20276 22156 20285 22196
rect 21510 22112 21600 22132
rect 1459 22072 1468 22112
rect 1508 22072 5828 22112
rect 8515 22072 8524 22112
rect 8564 22072 8716 22112
rect 8756 22072 8765 22112
rect 11251 22072 11260 22112
rect 11300 22072 11500 22112
rect 11540 22072 11549 22112
rect 18307 22072 18316 22112
rect 18356 22072 18932 22112
rect 19651 22072 19660 22112
rect 19700 22072 19939 22112
rect 19979 22072 19988 22112
rect 21283 22072 21292 22112
rect 21332 22072 21600 22112
rect 5788 22028 5828 22072
rect 21510 22052 21600 22072
rect 1411 21988 1420 22028
rect 1460 21988 4148 22028
rect 5788 21988 19412 22028
rect 0 21944 90 21964
rect 4108 21944 4148 21988
rect 19372 21944 19412 21988
rect 0 21904 1460 21944
rect 3679 21904 3688 21944
rect 3728 21904 3770 21944
rect 3810 21904 3852 21944
rect 3892 21904 3934 21944
rect 3974 21904 4016 21944
rect 4056 21904 4065 21944
rect 4108 21904 11212 21944
rect 11252 21904 11261 21944
rect 18799 21904 18808 21944
rect 18848 21904 18890 21944
rect 18930 21904 18972 21944
rect 19012 21904 19054 21944
rect 19094 21904 19136 21944
rect 19176 21904 19185 21944
rect 19372 21904 20044 21944
rect 20084 21904 20093 21944
rect 0 21884 90 21904
rect 1420 21860 1460 21904
rect 1411 21820 1420 21860
rect 1460 21820 1469 21860
rect 5260 21820 8332 21860
rect 8372 21820 8381 21860
rect 11299 21820 11308 21860
rect 11348 21820 11500 21860
rect 11540 21820 11549 21860
rect 18124 21820 19372 21860
rect 19412 21820 19421 21860
rect 5260 21776 5300 21820
rect 18124 21776 18164 21820
rect 1843 21736 1852 21776
rect 1892 21736 2860 21776
rect 2900 21736 2909 21776
rect 4265 21736 4348 21776
rect 4388 21736 4396 21776
rect 4436 21736 4445 21776
rect 5251 21736 5260 21776
rect 5300 21736 5309 21776
rect 6403 21736 6412 21776
rect 6452 21736 6892 21776
rect 6932 21736 8620 21776
rect 8660 21736 8669 21776
rect 8873 21736 9004 21776
rect 9044 21736 9053 21776
rect 14620 21736 15284 21776
rect 18115 21736 18124 21776
rect 18164 21736 18173 21776
rect 19363 21736 19372 21776
rect 19412 21736 19756 21776
rect 19796 21736 19805 21776
rect 20323 21736 20332 21776
rect 20372 21736 20524 21776
rect 20564 21736 20573 21776
rect 3811 21652 3820 21692
rect 3860 21652 9100 21692
rect 9140 21652 9149 21692
rect 0 21608 90 21628
rect 0 21568 980 21608
rect 1097 21568 1228 21608
rect 1268 21568 1277 21608
rect 1481 21568 1612 21608
rect 1652 21568 1661 21608
rect 1987 21568 1996 21608
rect 2036 21568 2380 21608
rect 2420 21568 2429 21608
rect 2947 21568 2956 21608
rect 2996 21568 3127 21608
rect 3907 21568 3916 21608
rect 3956 21568 4163 21608
rect 4291 21568 4300 21608
rect 4340 21568 4588 21608
rect 4628 21568 4637 21608
rect 5260 21568 6028 21608
rect 6068 21568 6077 21608
rect 7171 21568 7180 21608
rect 7220 21568 7948 21608
rect 7988 21568 8660 21608
rect 0 21548 90 21568
rect 940 21524 980 21568
rect 3532 21524 3572 21533
rect 4123 21524 4163 21568
rect 5260 21524 5300 21568
rect 6700 21524 6740 21533
rect 8620 21524 8660 21568
rect 940 21484 1132 21524
rect 1172 21484 1181 21524
rect 2458 21484 2467 21524
rect 2507 21484 2516 21524
rect 2563 21484 2572 21524
rect 2612 21484 2621 21524
rect 3043 21484 3052 21524
rect 3092 21484 3476 21524
rect 76 21316 212 21356
rect 1459 21316 1468 21356
rect 1508 21316 1612 21356
rect 1652 21316 1661 21356
rect 2227 21316 2236 21356
rect 2276 21316 2380 21356
rect 2420 21316 2429 21356
rect 76 21292 116 21316
rect 0 21232 116 21292
rect 172 21272 212 21316
rect 172 21232 1460 21272
rect 0 21212 90 21232
rect 0 20936 90 20956
rect 1420 20936 1460 21232
rect 2476 21020 2516 21484
rect 2572 21440 2612 21484
rect 2572 21400 3052 21440
rect 3092 21400 3101 21440
rect 3436 21356 3476 21484
rect 3619 21484 3628 21524
rect 3668 21484 4020 21524
rect 4060 21484 4069 21524
rect 4123 21484 4243 21524
rect 4283 21484 4292 21524
rect 4954 21484 4963 21524
rect 5003 21484 5012 21524
rect 5251 21484 5260 21524
rect 5300 21484 5309 21524
rect 5443 21484 5452 21524
rect 5492 21484 6412 21524
rect 6452 21484 6461 21524
rect 6740 21484 6988 21524
rect 7028 21484 7037 21524
rect 7363 21484 7372 21524
rect 7412 21484 7796 21524
rect 3532 21440 3572 21484
rect 4972 21440 5012 21484
rect 6700 21475 6740 21484
rect 7756 21440 7796 21484
rect 3532 21400 4204 21440
rect 4244 21400 4253 21440
rect 4972 21400 6508 21440
rect 6548 21400 6557 21440
rect 7756 21400 8332 21440
rect 8372 21400 8381 21440
rect 6508 21356 6548 21400
rect 8620 21356 8660 21484
rect 9196 21524 9236 21533
rect 10828 21524 10868 21533
rect 13708 21524 13748 21533
rect 14620 21524 14660 21736
rect 14794 21599 15044 21608
rect 14794 21559 14803 21599
rect 14843 21568 15044 21599
rect 14843 21559 14852 21568
rect 14794 21558 14852 21559
rect 15004 21524 15044 21568
rect 15244 21524 15284 21736
rect 16291 21652 16300 21692
rect 16340 21652 16436 21692
rect 16396 21608 16436 21652
rect 21510 21608 21600 21628
rect 15331 21568 15340 21608
rect 15380 21568 15619 21608
rect 15659 21568 15668 21608
rect 16396 21568 16724 21608
rect 16300 21524 16340 21533
rect 16684 21524 16724 21568
rect 18700 21568 19604 21608
rect 19747 21568 19756 21608
rect 19796 21568 21600 21608
rect 17932 21524 17972 21533
rect 18700 21524 18740 21568
rect 19564 21524 19604 21568
rect 21510 21548 21600 21568
rect 9236 21484 10156 21524
rect 10196 21484 10205 21524
rect 10273 21484 10348 21524
rect 10388 21484 10404 21524
rect 10444 21484 10453 21524
rect 11945 21484 12076 21524
rect 12116 21484 12125 21524
rect 12451 21484 12460 21524
rect 12500 21484 12509 21524
rect 13507 21484 13516 21524
rect 13556 21484 13708 21524
rect 13891 21484 13900 21524
rect 13940 21484 14092 21524
rect 14132 21484 14141 21524
rect 14225 21484 14234 21524
rect 14274 21484 14284 21524
rect 14324 21484 14414 21524
rect 14476 21484 14667 21524
rect 14707 21484 14716 21524
rect 14899 21484 14908 21524
rect 14948 21484 14957 21524
rect 15004 21484 15013 21524
rect 15053 21484 15062 21524
rect 15130 21484 15139 21524
rect 15179 21484 15188 21524
rect 15235 21484 15244 21524
rect 15284 21484 15293 21524
rect 15427 21484 15436 21524
rect 15476 21484 15479 21524
rect 15519 21484 15607 21524
rect 15715 21484 15724 21524
rect 15764 21484 15895 21524
rect 16169 21484 16300 21524
rect 16340 21484 16349 21524
rect 16675 21484 16684 21524
rect 16724 21484 17260 21524
rect 17300 21484 17309 21524
rect 17731 21484 17740 21524
rect 17780 21484 17932 21524
rect 17972 21484 18124 21524
rect 18164 21484 18173 21524
rect 18403 21484 18412 21524
rect 18452 21484 18700 21524
rect 18740 21484 18749 21524
rect 18857 21484 18979 21524
rect 19028 21484 19037 21524
rect 19171 21484 19180 21524
rect 19220 21484 19229 21524
rect 19555 21484 19564 21524
rect 19604 21484 19660 21524
rect 19700 21484 19735 21524
rect 19906 21484 19915 21524
rect 19955 21484 19964 21524
rect 20026 21484 20035 21524
rect 20084 21484 20215 21524
rect 9196 21475 9236 21484
rect 10828 21440 10868 21484
rect 8803 21400 8812 21440
rect 8852 21400 9100 21440
rect 9140 21400 9149 21440
rect 10492 21400 12364 21440
rect 12404 21400 12413 21440
rect 10492 21356 10532 21400
rect 12460 21356 12500 21484
rect 13708 21475 13748 21484
rect 14476 21440 14516 21484
rect 14908 21440 14948 21484
rect 13996 21400 14516 21440
rect 14659 21400 14668 21440
rect 14708 21400 14948 21440
rect 13996 21356 14036 21400
rect 3436 21316 3532 21356
rect 3572 21316 3581 21356
rect 5251 21316 5260 21356
rect 5300 21316 5548 21356
rect 5588 21316 5597 21356
rect 6508 21316 6892 21356
rect 6932 21316 6941 21356
rect 8620 21316 10532 21356
rect 10627 21316 10636 21356
rect 10676 21316 11020 21356
rect 11060 21316 11069 21356
rect 11203 21316 11212 21356
rect 11252 21316 12980 21356
rect 13865 21316 13900 21356
rect 13940 21316 13996 21356
rect 14036 21316 14045 21356
rect 14249 21316 14380 21356
rect 14420 21316 14429 21356
rect 14563 21316 14572 21356
rect 14612 21316 14743 21356
rect 12940 21272 12980 21316
rect 15004 21272 15044 21484
rect 15148 21440 15188 21484
rect 16300 21475 16340 21484
rect 17932 21475 17972 21484
rect 19180 21440 19220 21484
rect 19924 21440 19964 21484
rect 15148 21400 15340 21440
rect 15380 21400 15389 21440
rect 15802 21400 15811 21440
rect 15851 21400 15998 21440
rect 16038 21400 16047 21440
rect 16195 21400 16204 21440
rect 16244 21400 16253 21440
rect 19075 21400 19084 21440
rect 19124 21400 19133 21440
rect 19180 21400 19964 21440
rect 16204 21356 16244 21400
rect 15977 21316 16012 21356
rect 16052 21316 16099 21356
rect 16139 21316 16157 21356
rect 16204 21316 16588 21356
rect 16628 21316 16637 21356
rect 18259 21316 18268 21356
rect 18308 21316 18700 21356
rect 18740 21316 18749 21356
rect 19084 21272 19124 21400
rect 20227 21316 20236 21356
rect 20276 21316 20564 21356
rect 7660 21232 12844 21272
rect 12884 21232 12893 21272
rect 12940 21232 14476 21272
rect 14516 21232 14525 21272
rect 14659 21232 14668 21272
rect 14708 21232 15044 21272
rect 18115 21232 18124 21272
rect 18164 21232 19124 21272
rect 7660 21188 7700 21232
rect 4919 21148 4928 21188
rect 4968 21148 5010 21188
rect 5050 21148 5092 21188
rect 5132 21148 5174 21188
rect 5214 21148 5256 21188
rect 5296 21148 5305 21188
rect 6403 21148 6412 21188
rect 6452 21148 7700 21188
rect 8899 21148 8908 21188
rect 8948 21148 8957 21188
rect 9283 21148 9292 21188
rect 9332 21148 9341 21188
rect 10723 21148 10732 21188
rect 10772 21148 13324 21188
rect 13364 21148 13373 21188
rect 13603 21148 13612 21188
rect 13652 21148 17164 21188
rect 17204 21148 17213 21188
rect 20039 21148 20048 21188
rect 20088 21148 20130 21188
rect 20170 21148 20212 21188
rect 20252 21148 20294 21188
rect 20334 21148 20376 21188
rect 20416 21148 20425 21188
rect 8908 21020 8948 21148
rect 9292 21104 9332 21148
rect 20524 21104 20564 21316
rect 21510 21104 21600 21124
rect 9292 21064 15340 21104
rect 15380 21064 15389 21104
rect 20236 21064 20564 21104
rect 21475 21064 21484 21104
rect 21524 21064 21600 21104
rect 2476 20980 2668 21020
rect 2708 20980 2717 21020
rect 3475 20980 3484 21020
rect 3524 20980 4012 21020
rect 4052 20980 4061 21020
rect 5225 20980 5356 21020
rect 5396 20980 5405 21020
rect 5836 20980 8716 21020
rect 8756 20980 8765 21020
rect 8908 20980 9100 21020
rect 9140 20980 9292 21020
rect 9332 20980 9341 21020
rect 12940 20980 13460 21020
rect 15139 20980 15148 21020
rect 15188 20980 15724 21020
rect 15764 20980 15773 21020
rect 5836 20936 5876 20980
rect 0 20896 940 20936
rect 980 20896 989 20936
rect 1420 20896 5876 20936
rect 7075 20896 7084 20936
rect 7124 20896 7412 20936
rect 9091 20896 9100 20936
rect 9140 20896 9428 20936
rect 0 20876 90 20896
rect 7372 20852 7412 20896
rect 9388 20852 9428 20896
rect 1219 20812 1228 20852
rect 1268 20812 1900 20852
rect 1940 20812 1949 20852
rect 2371 20812 2380 20852
rect 2420 20843 2764 20852
rect 2420 20812 2476 20843
rect 2516 20812 2764 20843
rect 2804 20812 2813 20852
rect 3785 20812 3820 20852
rect 3860 20812 3916 20852
rect 3956 20812 3965 20852
rect 5033 20812 5164 20852
rect 5204 20812 5213 20852
rect 5635 20812 5644 20852
rect 5684 20812 5693 20852
rect 6115 20812 6124 20852
rect 6164 20843 7180 20852
rect 6164 20812 6892 20843
rect 2476 20794 2516 20803
rect 5164 20794 5204 20803
rect 5644 20768 5684 20812
rect 6932 20812 7180 20843
rect 7220 20812 7229 20852
rect 7354 20812 7363 20852
rect 7403 20812 7412 20852
rect 7459 20812 7468 20852
rect 7508 20812 7564 20852
rect 7604 20812 7639 20852
rect 7843 20812 7852 20852
rect 7892 20812 7901 20852
rect 8428 20843 8620 20852
rect 6892 20794 6932 20803
rect 2659 20728 2668 20768
rect 2708 20728 2860 20768
rect 2900 20728 2909 20768
rect 3235 20728 3244 20768
rect 3284 20728 3293 20768
rect 5251 20728 5260 20768
rect 5300 20728 5684 20768
rect 3244 20684 3284 20728
rect 5644 20684 5684 20728
rect 7852 20684 7892 20812
rect 8468 20812 8620 20843
rect 8660 20812 8669 20852
rect 8908 20843 9004 20852
rect 8428 20794 8468 20803
rect 8948 20812 9004 20843
rect 9044 20812 9079 20852
rect 9370 20812 9379 20852
rect 9419 20812 9428 20852
rect 9475 20812 9484 20852
rect 9524 20812 9580 20852
rect 9620 20812 9655 20852
rect 9859 20812 9868 20852
rect 9908 20812 10156 20852
rect 10196 20812 10205 20852
rect 10409 20843 10540 20852
rect 10409 20812 10444 20843
rect 8908 20794 8948 20803
rect 10484 20812 10540 20843
rect 10580 20812 10589 20852
rect 10889 20843 11020 20852
rect 10889 20812 10924 20843
rect 10444 20794 10484 20803
rect 10964 20812 11020 20843
rect 11060 20812 11069 20852
rect 11779 20812 11788 20852
rect 11828 20812 12076 20852
rect 12116 20812 12748 20852
rect 12788 20812 12797 20852
rect 10924 20794 10964 20803
rect 7939 20728 7948 20768
rect 7988 20728 8140 20768
rect 8180 20728 8189 20768
rect 9955 20728 9964 20768
rect 10004 20728 10013 20768
rect 11146 20728 11155 20768
rect 11195 20728 11500 20768
rect 11540 20728 11549 20768
rect 9964 20684 10004 20728
rect 12940 20684 12980 20980
rect 13420 20852 13460 20980
rect 13507 20896 13516 20936
rect 13556 20896 13612 20936
rect 13652 20896 13687 20936
rect 14659 20896 14668 20936
rect 14708 20896 16052 20936
rect 16243 20896 16252 20936
rect 16292 20896 16492 20936
rect 16532 20896 16541 20936
rect 17635 20896 17644 20936
rect 17684 20896 18412 20936
rect 18452 20896 18548 20936
rect 16012 20852 16052 20896
rect 18508 20852 18548 20896
rect 13328 20810 13368 20819
rect 13420 20812 13708 20852
rect 13748 20812 14380 20852
rect 14420 20812 14429 20852
rect 14960 20810 15000 20819
rect 15619 20812 15628 20852
rect 15668 20812 15677 20852
rect 15748 20812 15757 20852
rect 15797 20812 15820 20852
rect 15860 20812 15937 20852
rect 16003 20812 16012 20852
rect 16052 20812 16061 20852
rect 16195 20812 16204 20852
rect 16244 20812 16684 20852
rect 16724 20812 16733 20852
rect 17731 20812 17740 20852
rect 17780 20843 17972 20852
rect 17780 20812 17932 20843
rect 13324 20770 13328 20810
rect 13324 20768 13368 20770
rect 14956 20770 14960 20810
rect 14956 20768 15000 20770
rect 13324 20728 13516 20768
rect 13556 20761 15000 20768
rect 15628 20768 15668 20812
rect 18499 20812 18508 20852
rect 18548 20812 18557 20852
rect 19555 20812 19564 20852
rect 19604 20843 19796 20852
rect 19604 20812 19756 20843
rect 17932 20794 17972 20803
rect 19756 20794 19796 20803
rect 13556 20728 14996 20761
rect 15628 20728 16108 20768
rect 16148 20728 16157 20768
rect 16361 20728 16492 20768
rect 16532 20728 16541 20768
rect 20009 20728 20140 20768
rect 20180 20728 20189 20768
rect 15628 20684 15668 20728
rect 20236 20684 20276 21064
rect 21510 21044 21600 21064
rect 20371 20980 20380 21020
rect 20420 20980 20716 21020
rect 20756 20980 20765 21020
rect 3244 20644 3628 20684
rect 3668 20644 3677 20684
rect 5644 20644 6892 20684
rect 6932 20644 6941 20684
rect 7852 20644 8812 20684
rect 8852 20644 9388 20684
rect 9428 20644 9437 20684
rect 9964 20644 10924 20684
rect 10964 20644 10973 20684
rect 11020 20644 12980 20684
rect 13612 20644 15668 20684
rect 18115 20644 18124 20684
rect 18164 20644 20332 20684
rect 20372 20644 20436 20684
rect 0 20600 90 20620
rect 11020 20600 11060 20644
rect 0 20560 2860 20600
rect 2900 20560 2909 20600
rect 3091 20560 3100 20600
rect 3140 20560 3149 20600
rect 8035 20560 8044 20600
rect 8084 20560 11060 20600
rect 11251 20560 11260 20600
rect 11300 20560 11308 20600
rect 11348 20560 11431 20600
rect 0 20540 90 20560
rect 3100 20516 3140 20560
rect 3100 20476 10732 20516
rect 10772 20476 10781 20516
rect 13612 20432 13652 20644
rect 21510 20600 21600 20620
rect 15209 20560 15340 20600
rect 15380 20560 15389 20600
rect 18979 20560 18988 20600
rect 19028 20560 19316 20600
rect 19817 20560 19948 20600
rect 19988 20560 19997 20600
rect 20515 20560 20524 20600
rect 20564 20560 21600 20600
rect 14467 20476 14476 20516
rect 14516 20476 16108 20516
rect 16148 20476 16157 20516
rect 3679 20392 3688 20432
rect 3728 20392 3770 20432
rect 3810 20392 3852 20432
rect 3892 20392 3934 20432
rect 3974 20392 4016 20432
rect 4056 20392 4065 20432
rect 5539 20392 5548 20432
rect 5588 20392 11212 20432
rect 11252 20392 11261 20432
rect 13603 20392 13612 20432
rect 13652 20392 13661 20432
rect 13891 20392 13900 20432
rect 13940 20392 17260 20432
rect 17300 20392 17309 20432
rect 18799 20392 18808 20432
rect 18848 20392 18890 20432
rect 18930 20392 18972 20432
rect 19012 20392 19054 20432
rect 19094 20392 19136 20432
rect 19176 20392 19185 20432
rect 2860 20308 9676 20348
rect 9716 20308 9725 20348
rect 14371 20308 14380 20348
rect 14420 20308 18412 20348
rect 18452 20308 18461 20348
rect 0 20264 90 20284
rect 2860 20264 2900 20308
rect 19276 20264 19316 20560
rect 21510 20540 21600 20560
rect 0 20224 2900 20264
rect 6019 20224 6028 20264
rect 6068 20224 6604 20264
rect 6644 20224 6653 20264
rect 6883 20224 6892 20264
rect 6932 20224 11980 20264
rect 12020 20224 12029 20264
rect 13516 20224 14668 20264
rect 14708 20224 14717 20264
rect 15907 20224 15916 20264
rect 15956 20224 16492 20264
rect 16532 20224 16541 20264
rect 19171 20224 19180 20264
rect 19220 20224 19316 20264
rect 0 20204 90 20224
rect 13516 20180 13556 20224
rect 1603 20140 1612 20180
rect 1652 20140 10348 20180
rect 10388 20140 10397 20180
rect 13440 20140 13516 20180
rect 13556 20140 13565 20180
rect 13961 20140 14044 20180
rect 14084 20140 14092 20180
rect 14132 20140 14141 20180
rect 14188 20140 14516 20180
rect 15427 20140 15436 20180
rect 15476 20140 16300 20180
rect 16340 20140 16349 20180
rect 17836 20140 19564 20180
rect 19604 20140 19613 20180
rect 20179 20140 20188 20180
rect 20228 20140 21196 20180
rect 21236 20140 21245 20180
rect 259 20056 268 20096
rect 308 20056 2860 20096
rect 2900 20056 2909 20096
rect 3091 20056 3100 20096
rect 3140 20056 3340 20096
rect 3380 20056 3389 20096
rect 6508 20056 6988 20096
rect 7028 20056 7037 20096
rect 7171 20056 7180 20096
rect 7220 20056 8564 20096
rect 4780 20012 4820 20021
rect 6412 20012 6452 20021
rect 1097 19972 1228 20012
rect 1268 19972 1804 20012
rect 1844 19972 1853 20012
rect 2441 19972 2484 20012
rect 2524 19972 2572 20012
rect 2612 19972 2621 20012
rect 2860 19972 3532 20012
rect 3572 19972 4396 20012
rect 4436 19972 4445 20012
rect 5155 19972 5164 20012
rect 5204 19972 5356 20012
rect 5396 19972 5405 20012
rect 6281 19972 6316 20012
rect 6356 19972 6412 20012
rect 0 19928 90 19948
rect 2860 19928 2900 19972
rect 0 19888 844 19928
rect 884 19888 893 19928
rect 2572 19888 2900 19928
rect 4780 19928 4820 19972
rect 6316 19928 6356 19972
rect 6412 19963 6452 19972
rect 4780 19888 6356 19928
rect 0 19868 90 19888
rect 2572 19844 2612 19888
rect 6508 19844 6548 20056
rect 8524 20012 8564 20056
rect 10156 20056 10924 20096
rect 10964 20056 10973 20096
rect 11107 20056 11116 20096
rect 11156 20056 11165 20096
rect 12394 20056 12403 20096
rect 12443 20056 12748 20096
rect 12788 20056 12797 20096
rect 12931 20056 12940 20096
rect 12980 20056 12989 20096
rect 13171 20056 13180 20096
rect 13220 20056 13324 20096
rect 13364 20056 13373 20096
rect 10156 20012 10196 20056
rect 7075 19972 7084 20012
rect 7124 19972 7276 20012
rect 7316 19972 7325 20012
rect 8777 19972 8908 20012
rect 8948 19972 8957 20012
rect 10060 19972 10156 20012
rect 8524 19963 8564 19972
rect 8707 19888 8716 19928
rect 8756 19888 9004 19928
rect 9044 19888 9053 19928
rect 1891 19804 1900 19844
rect 1940 19804 2612 19844
rect 2659 19804 2668 19844
rect 2708 19804 2717 19844
rect 4387 19804 4396 19844
rect 4436 19804 4972 19844
rect 5012 19804 5021 19844
rect 5443 19804 5452 19844
rect 5492 19804 6548 19844
rect 6604 19804 6748 19844
rect 6788 19804 6797 19844
rect 0 19592 90 19612
rect 0 19552 460 19592
rect 500 19552 509 19592
rect 0 19532 90 19552
rect 2668 19340 2708 19804
rect 6604 19760 6644 19804
rect 10060 19760 10100 19972
rect 10156 19963 10196 19972
rect 10348 19972 10627 20012
rect 10667 19972 10676 20012
rect 10723 19972 10732 20012
rect 10772 19972 10781 20012
rect 10348 19928 10388 19972
rect 10732 19928 10772 19972
rect 10339 19888 10348 19928
rect 10388 19888 10397 19928
rect 10636 19888 10772 19928
rect 10636 19844 10676 19888
rect 10147 19804 10156 19844
rect 10196 19804 10676 19844
rect 11116 19844 11156 20056
rect 11692 20012 11732 20021
rect 12940 20012 12980 20056
rect 13516 20012 13556 20140
rect 14188 20096 14228 20140
rect 13795 20056 13804 20096
rect 13844 20056 14228 20096
rect 14476 20096 14516 20140
rect 14476 20056 16340 20096
rect 16387 20056 16396 20096
rect 16436 20056 17740 20096
rect 17780 20056 17789 20096
rect 11203 19972 11212 20012
rect 11252 19972 11383 20012
rect 11561 19972 11692 20012
rect 11732 19972 11741 20012
rect 11971 19972 11980 20012
rect 12020 19972 12180 20012
rect 12220 19972 12229 20012
rect 12451 19972 12460 20012
rect 12500 19972 12980 20012
rect 13507 19972 13516 20012
rect 13556 19972 13565 20012
rect 13651 19972 13660 20012
rect 13700 19972 14135 20012
rect 14175 19972 14184 20012
rect 14266 20007 14275 20012
rect 14236 19972 14275 20007
rect 14315 19972 14324 20012
rect 14371 19972 14380 20012
rect 14420 19972 14551 20012
rect 14755 19972 14764 20012
rect 14804 19972 14935 20012
rect 15034 19972 15043 20012
rect 15083 19972 15092 20012
rect 15235 19972 15244 20012
rect 15284 19972 15619 20012
rect 15659 19972 15668 20012
rect 15881 19972 15930 20012
rect 15970 19972 16012 20012
rect 16052 19972 16061 20012
rect 11692 19963 11732 19972
rect 12172 19888 13516 19928
rect 13556 19888 13708 19928
rect 13748 19888 13757 19928
rect 12172 19844 12212 19888
rect 13900 19844 13940 19972
rect 14236 19967 14324 19972
rect 11116 19804 12212 19844
rect 12355 19804 12364 19844
rect 12404 19804 12508 19844
rect 12548 19804 12557 19844
rect 13891 19804 13900 19844
rect 13940 19804 13949 19844
rect 5923 19720 5932 19760
rect 5972 19720 6644 19760
rect 7843 19720 7852 19760
rect 7892 19720 10100 19760
rect 14236 19760 14276 19967
rect 15052 19928 15092 19972
rect 14685 19888 15092 19928
rect 15139 19888 15148 19928
rect 15188 19888 16052 19928
rect 14685 19844 14725 19888
rect 16012 19844 16052 19888
rect 14458 19804 14467 19844
rect 14507 19804 14516 19844
rect 14659 19804 14668 19844
rect 14708 19804 14725 19844
rect 14860 19804 15715 19844
rect 15755 19804 15764 19844
rect 16003 19804 16012 19844
rect 16052 19804 16061 19844
rect 16147 19804 16156 19844
rect 16196 19804 16244 19844
rect 14476 19760 14516 19804
rect 14236 19720 14380 19760
rect 14420 19720 14429 19760
rect 14476 19720 14612 19760
rect 14572 19676 14612 19720
rect 14860 19676 14900 19804
rect 4919 19636 4928 19676
rect 4968 19636 5010 19676
rect 5050 19636 5092 19676
rect 5132 19636 5174 19676
rect 5214 19636 5256 19676
rect 5296 19636 5305 19676
rect 6211 19636 6220 19676
rect 6260 19636 8084 19676
rect 8899 19636 8908 19676
rect 8948 19636 10444 19676
rect 10484 19636 11212 19676
rect 11252 19636 11261 19676
rect 14572 19636 14900 19676
rect 16204 19676 16244 19804
rect 16300 19760 16340 20056
rect 17836 20012 17876 20140
rect 21510 20096 21600 20116
rect 18019 20056 18028 20096
rect 18068 20056 18452 20096
rect 18499 20056 18508 20096
rect 18548 20056 18796 20096
rect 18836 20056 18845 20096
rect 21196 20056 21600 20096
rect 18412 20012 18452 20056
rect 19371 20012 19411 20021
rect 21196 20012 21236 20056
rect 21510 20036 21600 20056
rect 16553 19972 16588 20012
rect 16628 19972 16684 20012
rect 16724 19972 16733 20012
rect 17705 19972 17836 20012
rect 17876 19972 17885 20012
rect 18028 19972 18307 20012
rect 18347 19972 18356 20012
rect 18403 19972 18412 20012
rect 18452 19972 18461 20012
rect 18761 19972 18892 20012
rect 18932 19972 18941 20012
rect 19075 19972 19084 20012
rect 19124 19972 19371 20012
rect 19817 19972 19891 20012
rect 19931 19972 19948 20012
rect 19988 19972 19997 20012
rect 20201 19972 20332 20012
rect 20372 19972 20381 20012
rect 21187 19972 21196 20012
rect 21236 19972 21245 20012
rect 17836 19963 17876 19972
rect 18028 19928 18068 19972
rect 19371 19963 19411 19972
rect 18019 19888 18028 19928
rect 18068 19888 18077 19928
rect 19913 19804 20044 19844
rect 20084 19804 20093 19844
rect 16300 19720 20948 19760
rect 16204 19636 17164 19676
rect 17204 19636 17213 19676
rect 20039 19636 20048 19676
rect 20088 19636 20130 19676
rect 20170 19636 20212 19676
rect 20252 19636 20294 19676
rect 20334 19636 20376 19676
rect 20416 19636 20425 19676
rect 5923 19552 5932 19592
rect 5972 19552 7508 19592
rect 7468 19508 7508 19552
rect 8044 19508 8084 19636
rect 20908 19592 20948 19720
rect 21510 19592 21600 19612
rect 14860 19552 15436 19592
rect 15476 19552 15485 19592
rect 16003 19552 16012 19592
rect 16052 19552 18124 19592
rect 18164 19552 18173 19592
rect 18796 19552 20524 19592
rect 20564 19552 20573 19592
rect 20908 19552 21600 19592
rect 14860 19508 14900 19552
rect 18796 19508 18836 19552
rect 21510 19532 21600 19552
rect 4195 19468 4204 19508
rect 4244 19468 4724 19508
rect 4771 19468 4780 19508
rect 4820 19468 5260 19508
rect 5300 19468 5309 19508
rect 7363 19468 7372 19508
rect 7412 19468 7421 19508
rect 7468 19468 7900 19508
rect 7940 19468 7949 19508
rect 8044 19468 8668 19508
rect 8708 19468 8717 19508
rect 10099 19468 10108 19508
rect 10148 19468 10252 19508
rect 10292 19468 10301 19508
rect 11107 19468 11116 19508
rect 11156 19468 11828 19508
rect 11971 19468 11980 19508
rect 12020 19468 12268 19508
rect 12308 19468 12317 19508
rect 14227 19468 14236 19508
rect 14276 19468 14476 19508
rect 14516 19468 14525 19508
rect 14659 19468 14668 19508
rect 14708 19468 14900 19508
rect 15113 19468 15244 19508
rect 15284 19468 15293 19508
rect 15955 19468 15964 19508
rect 16004 19468 18836 19508
rect 20009 19468 20140 19508
rect 20180 19468 20189 19508
rect 4684 19424 4724 19468
rect 7372 19424 7412 19468
rect 11788 19424 11828 19468
rect 2755 19384 2764 19424
rect 2804 19384 4628 19424
rect 4684 19384 5012 19424
rect 5539 19384 5548 19424
rect 5588 19384 5876 19424
rect 7372 19384 8180 19424
rect 10435 19384 10444 19424
rect 10484 19384 11596 19424
rect 11636 19384 11645 19424
rect 11788 19384 13228 19424
rect 13268 19384 13277 19424
rect 14380 19384 14572 19424
rect 14612 19384 14621 19424
rect 14755 19384 14764 19424
rect 14804 19384 14900 19424
rect 15139 19384 15148 19424
rect 15188 19384 16588 19424
rect 16628 19384 16637 19424
rect 17923 19384 17932 19424
rect 17972 19384 18452 19424
rect 1315 19300 1324 19340
rect 1364 19300 1612 19340
rect 1652 19300 1996 19340
rect 2036 19300 2045 19340
rect 2441 19300 2572 19340
rect 2612 19300 2621 19340
rect 2668 19300 3043 19340
rect 3083 19300 3092 19340
rect 3139 19300 3148 19340
rect 3188 19300 3197 19340
rect 3340 19300 3532 19340
rect 3572 19300 3581 19340
rect 4073 19331 4204 19340
rect 4073 19300 4108 19331
rect 2572 19282 2612 19291
rect 0 19256 90 19276
rect 3148 19256 3188 19300
rect 0 19216 748 19256
rect 788 19216 797 19256
rect 2956 19216 3188 19256
rect 0 19196 90 19216
rect 2956 19088 2996 19216
rect 3340 19172 3380 19300
rect 4148 19300 4204 19331
rect 4244 19300 4253 19340
rect 4588 19331 4628 19384
rect 4108 19282 4148 19291
rect 4588 19282 4628 19291
rect 4972 19256 5012 19384
rect 5836 19340 5876 19384
rect 5356 19300 5635 19340
rect 5675 19300 5684 19340
rect 5731 19300 5740 19340
rect 5780 19300 5789 19340
rect 5836 19331 6740 19340
rect 5836 19300 6700 19331
rect 3497 19216 3628 19256
rect 3668 19216 3677 19256
rect 4963 19216 4972 19256
rect 5012 19216 5021 19256
rect 5356 19172 5396 19300
rect 3043 19132 3052 19172
rect 3092 19132 3380 19172
rect 4387 19132 4396 19172
rect 4436 19132 5396 19172
rect 2956 19048 3436 19088
rect 3476 19048 3485 19088
rect 4195 19048 4204 19088
rect 4244 19048 5212 19088
rect 5252 19048 5261 19088
rect 0 18920 90 18940
rect 0 18880 3532 18920
rect 3572 18880 3581 18920
rect 3679 18880 3688 18920
rect 3728 18880 3770 18920
rect 3810 18880 3852 18920
rect 3892 18880 3934 18920
rect 3974 18880 4016 18920
rect 4056 18880 4065 18920
rect 0 18860 90 18880
rect 5740 18752 5780 19300
rect 6700 19282 6740 19291
rect 7180 19331 7220 19340
rect 7180 19256 7220 19291
rect 8140 19256 8180 19384
rect 10828 19340 10868 19384
rect 14380 19340 14420 19384
rect 14860 19340 14900 19384
rect 8323 19300 8332 19340
rect 8372 19300 9908 19340
rect 10051 19300 10060 19340
rect 10100 19300 10484 19340
rect 10819 19300 10828 19340
rect 10868 19300 10877 19340
rect 12076 19331 12460 19340
rect 9868 19256 9908 19300
rect 10444 19256 10484 19300
rect 12116 19300 12460 19331
rect 12500 19300 12652 19340
rect 12692 19300 12701 19340
rect 13865 19300 13996 19340
rect 14036 19300 14045 19340
rect 14371 19300 14380 19340
rect 14420 19300 14429 19340
rect 14563 19300 14572 19340
rect 14612 19300 14621 19340
rect 14746 19300 14755 19340
rect 14795 19300 14804 19340
rect 14860 19300 15043 19340
rect 15083 19300 15092 19340
rect 12076 19282 12116 19291
rect 14572 19256 14612 19300
rect 5993 19216 6124 19256
rect 6164 19216 6173 19256
rect 6250 19216 6259 19256
rect 6299 19216 6308 19256
rect 7171 19216 7180 19256
rect 7220 19216 7267 19256
rect 7721 19216 7756 19256
rect 7796 19216 7852 19256
rect 7892 19216 7901 19256
rect 8131 19216 8140 19256
rect 8180 19216 8189 19256
rect 8393 19216 8428 19256
rect 8468 19216 8524 19256
rect 8564 19216 8573 19256
rect 8707 19216 8716 19256
rect 8756 19216 8908 19256
rect 8948 19216 8957 19256
rect 9091 19216 9100 19256
rect 9140 19216 9271 19256
rect 9545 19216 9676 19256
rect 9716 19216 9725 19256
rect 9859 19216 9868 19256
rect 9908 19216 9917 19256
rect 9964 19216 10388 19256
rect 10435 19216 10444 19256
rect 10484 19216 10493 19256
rect 13891 19216 13900 19256
rect 13940 19216 14612 19256
rect 14764 19256 14804 19300
rect 14764 19216 15052 19256
rect 15092 19216 15101 19256
rect 6268 19172 6308 19216
rect 9964 19172 10004 19216
rect 6211 19132 6220 19172
rect 6260 19132 8044 19172
rect 8084 19132 8093 19172
rect 9331 19132 9340 19172
rect 9380 19132 10004 19172
rect 10348 19172 10388 19216
rect 15148 19172 15188 19384
rect 18412 19340 18452 19384
rect 18988 19384 19852 19424
rect 19892 19384 19901 19424
rect 15345 19300 15354 19340
rect 15394 19300 15724 19340
rect 15764 19300 15773 19340
rect 16099 19300 16108 19340
rect 16148 19300 16492 19340
rect 16532 19300 16541 19340
rect 17705 19331 17836 19340
rect 17705 19300 17740 19331
rect 17780 19300 17836 19331
rect 17876 19300 17885 19340
rect 18394 19300 18403 19340
rect 18443 19300 18452 19340
rect 18499 19300 18508 19340
rect 18548 19300 18679 19340
rect 18761 19300 18892 19340
rect 18932 19300 18941 19340
rect 17740 19282 17780 19291
rect 18988 19256 19028 19384
rect 19116 19300 19180 19340
rect 19220 19331 19508 19340
rect 19220 19300 19468 19331
rect 10348 19132 13804 19172
rect 13844 19132 13853 19172
rect 14131 19132 14140 19172
rect 14180 19132 15188 19172
rect 15532 19216 15676 19256
rect 15716 19216 15725 19256
rect 15811 19216 15820 19256
rect 15860 19216 16300 19256
rect 16340 19216 16349 19256
rect 18700 19216 18988 19256
rect 19028 19216 19037 19256
rect 15532 19088 15572 19216
rect 15820 19132 16012 19172
rect 16052 19132 16061 19172
rect 15820 19088 15860 19132
rect 6307 19048 6316 19088
rect 6356 19048 7516 19088
rect 7556 19048 7565 19088
rect 8275 19048 8284 19088
rect 8324 19048 8333 19088
rect 8620 19048 9436 19088
rect 9476 19048 9485 19088
rect 9667 19048 9676 19088
rect 9716 19048 10204 19088
rect 10244 19048 10253 19088
rect 13027 19048 13036 19088
rect 13076 19048 15572 19088
rect 15811 19048 15820 19088
rect 15860 19048 15869 19088
rect 16012 19048 16060 19088
rect 16100 19048 16109 19088
rect 8284 18920 8324 19048
rect 6787 18880 6796 18920
rect 6836 18880 8324 18920
rect 8620 18836 8660 19048
rect 16012 19004 16052 19048
rect 15043 18964 15052 19004
rect 15092 18964 16012 19004
rect 16052 18964 16061 19004
rect 8899 18880 8908 18920
rect 8948 18880 12364 18920
rect 12404 18880 12413 18920
rect 18700 18836 18740 19216
rect 18799 18880 18808 18920
rect 18848 18880 18890 18920
rect 18930 18880 18972 18920
rect 19012 18880 19054 18920
rect 19094 18880 19136 18920
rect 19176 18880 19185 18920
rect 19276 18836 19316 19300
rect 19817 19300 19948 19340
rect 19988 19300 19997 19340
rect 19468 19282 19508 19291
rect 19948 19282 19988 19291
rect 21510 19088 21600 19108
rect 20707 19048 20716 19088
rect 20756 19048 21600 19088
rect 21510 19028 21600 19048
rect 6499 18796 6508 18836
rect 6548 18796 8660 18836
rect 11395 18796 11404 18836
rect 11444 18796 18508 18836
rect 18548 18796 18557 18836
rect 18700 18796 18836 18836
rect 18796 18752 18836 18796
rect 19180 18796 19316 18836
rect 19180 18752 19220 18796
rect 1459 18712 1468 18752
rect 1508 18712 1804 18752
rect 1844 18712 1853 18752
rect 3523 18712 3532 18752
rect 3572 18712 9004 18752
rect 9044 18712 9053 18752
rect 18787 18712 18796 18752
rect 18836 18712 18845 18752
rect 19171 18712 19180 18752
rect 19220 18712 19229 18752
rect 19555 18712 19564 18752
rect 19604 18712 19613 18752
rect 19817 18712 19948 18752
rect 19988 18712 19997 18752
rect 19564 18668 19604 18712
rect 1132 18628 9676 18668
rect 9716 18628 9725 18668
rect 13420 18628 14284 18668
rect 14324 18628 14333 18668
rect 15532 18628 17012 18668
rect 17059 18628 17068 18668
rect 17108 18628 17780 18668
rect 18115 18628 18124 18668
rect 18164 18628 19468 18668
rect 19508 18628 19517 18668
rect 19564 18628 19796 18668
rect 20371 18628 20380 18668
rect 20420 18628 20812 18668
rect 20852 18628 20861 18668
rect 0 18584 90 18604
rect 1132 18584 1172 18628
rect 0 18544 1172 18584
rect 1219 18544 1228 18584
rect 1268 18544 1324 18584
rect 1364 18544 1399 18584
rect 1603 18544 1612 18584
rect 1652 18544 1661 18584
rect 1987 18544 1996 18584
rect 2036 18544 2045 18584
rect 2825 18544 2956 18584
rect 2996 18544 3005 18584
rect 4169 18544 4243 18584
rect 4283 18544 4300 18584
rect 4340 18544 4349 18584
rect 4457 18544 4588 18584
rect 4628 18544 4637 18584
rect 4771 18544 4780 18584
rect 4820 18544 4951 18584
rect 5033 18544 5068 18584
rect 5108 18544 5164 18584
rect 5204 18544 5213 18584
rect 5395 18544 5404 18584
rect 5444 18544 5740 18584
rect 5780 18544 5789 18584
rect 6499 18544 6508 18584
rect 6548 18544 6557 18584
rect 7180 18544 7852 18584
rect 7892 18544 7901 18584
rect 8035 18544 8044 18584
rect 8084 18544 8716 18584
rect 8756 18544 8765 18584
rect 9322 18544 9331 18584
rect 9371 18544 9676 18584
rect 9716 18544 9725 18584
rect 12931 18544 12940 18584
rect 12980 18544 13324 18584
rect 13364 18544 13373 18584
rect 0 18524 90 18544
rect 1612 18500 1652 18544
rect 1996 18500 2036 18544
rect 3532 18500 3572 18509
rect 6508 18500 6548 18544
rect 6988 18500 7028 18509
rect 7180 18500 7220 18544
rect 11980 18500 12020 18509
rect 13420 18500 13460 18628
rect 15532 18584 15572 18628
rect 547 18460 556 18500
rect 596 18460 1652 18500
rect 1708 18460 2036 18500
rect 2315 18460 2380 18500
rect 2420 18460 2446 18500
rect 2486 18460 2495 18500
rect 2563 18460 2572 18500
rect 2612 18460 2860 18500
rect 2900 18460 2996 18500
rect 3043 18460 3052 18500
rect 3092 18460 3340 18500
rect 3380 18460 3389 18500
rect 4003 18460 4012 18500
rect 4060 18460 4183 18500
rect 5731 18460 5740 18500
rect 5780 18460 6548 18500
rect 6979 18460 6988 18500
rect 7028 18460 7220 18500
rect 7267 18460 7276 18500
rect 7316 18460 7555 18500
rect 7595 18460 7604 18500
rect 7651 18460 7660 18500
rect 7700 18460 7831 18500
rect 8009 18460 8140 18500
rect 8180 18460 8189 18500
rect 8614 18460 8623 18500
rect 8663 18460 9044 18500
rect 9091 18460 9100 18500
rect 9148 18460 9271 18500
rect 10572 18460 10636 18500
rect 10676 18460 10732 18500
rect 10772 18460 10924 18500
rect 10964 18460 10973 18500
rect 11683 18460 11692 18500
rect 11732 18460 11980 18500
rect 1708 18416 1748 18460
rect 2956 18416 2996 18460
rect 3532 18416 3572 18460
rect 6988 18451 7028 18460
rect 7660 18416 7700 18460
rect 9004 18416 9044 18460
rect 11980 18451 12020 18460
rect 12172 18460 12451 18500
rect 12491 18460 12500 18500
rect 12547 18460 12556 18500
rect 12596 18460 12605 18500
rect 13027 18460 13036 18500
rect 13076 18460 13460 18500
rect 13516 18544 15572 18584
rect 16972 18584 17012 18628
rect 17740 18584 17780 18628
rect 16972 18544 17164 18584
rect 17204 18544 17213 18584
rect 17731 18544 17740 18584
rect 17780 18544 17789 18584
rect 17923 18544 17932 18584
rect 17972 18544 18124 18584
rect 18164 18544 18173 18584
rect 18316 18544 18700 18584
rect 18740 18544 18749 18584
rect 13516 18500 13556 18544
rect 15628 18500 15668 18509
rect 17260 18500 17300 18509
rect 18316 18500 18356 18544
rect 19756 18500 19796 18628
rect 21510 18584 21600 18604
rect 20009 18544 20140 18584
rect 20180 18544 20189 18584
rect 20236 18544 21600 18584
rect 20236 18500 20276 18544
rect 21510 18524 21600 18544
rect 13891 18460 13900 18500
rect 13940 18460 14004 18500
rect 14044 18460 14071 18500
rect 14284 18460 14380 18500
rect 14420 18460 14429 18500
rect 15331 18460 15340 18500
rect 15380 18460 15628 18500
rect 15977 18460 16012 18500
rect 16052 18460 16108 18500
rect 16148 18460 16300 18500
rect 16340 18460 16349 18500
rect 17827 18460 17836 18500
rect 17876 18460 18124 18500
rect 18164 18460 18173 18500
rect 18307 18460 18316 18500
rect 18356 18460 18365 18500
rect 18412 18460 18508 18500
rect 18548 18460 18557 18500
rect 19939 18460 19948 18500
rect 19988 18460 20276 18500
rect 12172 18416 12212 18460
rect 12556 18416 12596 18460
rect 13516 18451 13556 18460
rect 14284 18416 14324 18460
rect 67 18376 76 18416
rect 116 18376 1748 18416
rect 1843 18376 1852 18416
rect 1892 18376 2668 18416
rect 2708 18376 2717 18416
rect 2956 18376 3052 18416
rect 3092 18376 3101 18416
rect 3235 18376 3244 18416
rect 3284 18376 3572 18416
rect 3619 18376 3628 18416
rect 3668 18376 4348 18416
rect 4388 18376 4397 18416
rect 4889 18376 4972 18416
rect 5012 18376 5020 18416
rect 5060 18376 5069 18416
rect 5155 18376 5164 18416
rect 5204 18376 6508 18416
rect 6548 18376 6557 18416
rect 7171 18376 7180 18416
rect 7220 18376 7351 18416
rect 7660 18376 8428 18416
rect 8468 18376 8477 18416
rect 8995 18376 9004 18416
rect 9044 18376 9053 18416
rect 12163 18376 12172 18416
rect 12212 18376 12221 18416
rect 12556 18376 12940 18416
rect 12980 18376 13132 18416
rect 13172 18376 13181 18416
rect 14092 18376 14324 18416
rect 15628 18416 15668 18460
rect 17260 18416 17300 18460
rect 18412 18416 18452 18460
rect 19756 18451 19796 18460
rect 15628 18376 17300 18416
rect 18307 18376 18316 18416
rect 18356 18376 18452 18416
rect 355 18292 364 18332
rect 404 18292 2236 18332
rect 2276 18292 2285 18332
rect 7555 18292 7564 18332
rect 7604 18292 9436 18332
rect 9476 18292 9485 18332
rect 12067 18292 12076 18332
rect 12116 18292 12268 18332
rect 12308 18292 12317 18332
rect 0 18248 90 18268
rect 14092 18248 14132 18376
rect 14179 18292 14188 18332
rect 14228 18292 14237 18332
rect 0 18208 556 18248
rect 596 18208 605 18248
rect 4771 18208 4780 18248
rect 4820 18208 7660 18248
rect 7700 18208 14132 18248
rect 0 18188 90 18208
rect 1795 18124 1804 18164
rect 1844 18124 2900 18164
rect 4919 18124 4928 18164
rect 4968 18124 5010 18164
rect 5050 18124 5092 18164
rect 5132 18124 5174 18164
rect 5214 18124 5256 18164
rect 5296 18124 5305 18164
rect 8035 18124 8044 18164
rect 8084 18124 10156 18164
rect 10196 18124 10205 18164
rect 12940 18124 13612 18164
rect 13652 18124 13661 18164
rect 2860 18080 2900 18124
rect 2860 18040 9236 18080
rect 9196 17996 9236 18040
rect 12940 17996 12980 18124
rect 1385 17956 1468 17996
rect 1508 17956 1516 17996
rect 1556 17956 1565 17996
rect 3043 17956 3052 17996
rect 3092 17956 4012 17996
rect 4052 17956 4061 17996
rect 5155 17956 5164 17996
rect 5204 17956 5836 17996
rect 5876 17956 5885 17996
rect 8131 17956 8140 17996
rect 8180 17956 9100 17996
rect 9140 17956 9149 17996
rect 9196 17956 12980 17996
rect 13315 17956 13324 17996
rect 13364 17956 13900 17996
rect 13940 17956 13949 17996
rect 0 17912 90 17932
rect 0 17872 1804 17912
rect 1844 17872 1853 17912
rect 4492 17872 5492 17912
rect 5539 17872 5548 17912
rect 5588 17872 5692 17912
rect 5732 17872 5741 17912
rect 6499 17872 6508 17912
rect 6548 17872 6740 17912
rect 8419 17872 8428 17912
rect 8468 17872 8564 17912
rect 8611 17872 8620 17912
rect 8660 17872 9524 17912
rect 0 17852 90 17872
rect 4492 17828 4532 17872
rect 5452 17828 5492 17872
rect 6700 17828 6740 17872
rect 8524 17828 8564 17872
rect 9484 17828 9524 17872
rect 9580 17872 12268 17912
rect 12308 17872 12317 17912
rect 1481 17788 1612 17828
rect 1652 17788 1661 17828
rect 2851 17788 2860 17828
rect 2900 17788 3031 17828
rect 3235 17788 3244 17828
rect 3284 17788 3427 17828
rect 3467 17788 3476 17828
rect 3523 17788 3532 17828
rect 3572 17788 3703 17828
rect 3907 17788 3916 17828
rect 3956 17788 4087 17828
rect 4361 17788 4492 17828
rect 4532 17788 4541 17828
rect 4675 17788 4684 17828
rect 4724 17819 5012 17828
rect 4724 17788 4972 17819
rect 2860 17770 2900 17779
rect 4492 17770 4532 17779
rect 5452 17788 6028 17828
rect 6068 17788 6077 17828
rect 6691 17788 6700 17828
rect 6740 17788 7372 17828
rect 7412 17788 7421 17828
rect 7843 17788 7852 17828
rect 7892 17819 8023 17828
rect 7892 17788 7948 17819
rect 4972 17770 5012 17779
rect 7988 17788 8023 17819
rect 8131 17788 8140 17828
rect 8180 17788 8419 17828
rect 8459 17788 8468 17828
rect 8515 17788 8524 17828
rect 8564 17788 8573 17828
rect 8748 17788 8812 17828
rect 8852 17788 8908 17828
rect 8948 17788 9100 17828
rect 9140 17788 9149 17828
rect 9353 17788 9484 17828
rect 9524 17788 9533 17828
rect 7948 17770 7988 17779
rect 9484 17770 9524 17779
rect 643 17704 652 17744
rect 692 17704 1228 17744
rect 1268 17704 1277 17744
rect 4003 17704 4012 17744
rect 4052 17704 4183 17744
rect 5225 17704 5356 17744
rect 5396 17704 5405 17744
rect 5731 17704 5740 17744
rect 5780 17704 5932 17744
rect 5972 17704 5981 17744
rect 6115 17704 6124 17744
rect 6164 17704 6508 17744
rect 6548 17704 7892 17744
rect 8515 17704 8524 17744
rect 8564 17704 9004 17744
rect 9044 17704 9053 17744
rect 7852 17660 7892 17704
rect 9580 17660 9620 17872
rect 9964 17819 10636 17828
rect 10004 17788 10636 17819
rect 10676 17788 10685 17828
rect 11849 17788 11884 17828
rect 11924 17788 11980 17828
rect 12020 17788 12556 17828
rect 12596 17788 12605 17828
rect 12940 17819 13172 17828
rect 12940 17788 13132 17819
rect 9964 17770 10004 17779
rect 12940 17744 12980 17788
rect 13132 17770 13172 17779
rect 10147 17704 10156 17744
rect 10235 17704 10327 17744
rect 10627 17704 10636 17744
rect 10676 17704 11020 17744
rect 11060 17704 11069 17744
rect 11683 17704 11692 17744
rect 11732 17704 12980 17744
rect 14188 17744 14228 18292
rect 14284 18164 14324 18376
rect 15235 18292 15244 18332
rect 15284 18292 15820 18332
rect 15860 18292 15869 18332
rect 17443 18292 17452 18332
rect 17492 18292 17501 18332
rect 17971 18292 17980 18332
rect 18020 18292 18260 18332
rect 14284 18124 16108 18164
rect 16148 18124 16876 18164
rect 16916 18124 16925 18164
rect 14956 18040 15244 18080
rect 15284 18040 15293 18080
rect 14956 17828 14996 18040
rect 15043 17872 15052 17912
rect 15092 17872 16492 17912
rect 16532 17872 16541 17912
rect 15724 17828 15764 17872
rect 17452 17828 17492 18292
rect 18220 18248 18260 18292
rect 18220 18208 21484 18248
rect 21524 18208 21533 18248
rect 17923 18124 17932 18164
rect 17972 18124 18412 18164
rect 18452 18124 18461 18164
rect 20039 18124 20048 18164
rect 20088 18124 20130 18164
rect 20170 18124 20212 18164
rect 20252 18124 20294 18164
rect 20334 18124 20376 18164
rect 20416 18124 20425 18164
rect 21510 18080 21600 18100
rect 19363 18040 19372 18080
rect 19412 18040 21600 18080
rect 21510 18020 21600 18040
rect 20371 17956 20380 17996
rect 20420 17956 21100 17996
rect 21140 17956 21149 17996
rect 14956 17788 15139 17828
rect 15179 17788 15188 17828
rect 15235 17788 15244 17828
rect 15284 17788 15415 17828
rect 15715 17788 15724 17828
rect 15764 17788 15773 17828
rect 16204 17819 16244 17828
rect 16553 17788 16684 17828
rect 16724 17788 16733 17828
rect 17251 17788 17260 17828
rect 17300 17788 17396 17828
rect 17452 17788 17539 17828
rect 17579 17788 17588 17828
rect 17635 17788 17644 17828
rect 17684 17788 17693 17828
rect 17932 17788 18028 17828
rect 18068 17788 18077 17828
rect 18604 17819 18691 17828
rect 16204 17744 16244 17779
rect 16684 17770 16724 17779
rect 17356 17744 17396 17788
rect 17644 17744 17684 17788
rect 14188 17704 14380 17744
rect 14420 17704 14429 17744
rect 14851 17704 14860 17744
rect 14900 17704 15284 17744
rect 15497 17704 15628 17744
rect 15668 17704 15677 17744
rect 16204 17704 16492 17744
rect 16532 17704 16541 17744
rect 16906 17704 16915 17744
rect 16955 17704 17260 17744
rect 17300 17704 17309 17744
rect 17356 17704 17836 17744
rect 17876 17704 17885 17744
rect 4867 17620 4876 17660
rect 4916 17620 7564 17660
rect 7604 17620 7613 17660
rect 7852 17620 9620 17660
rect 9955 17620 9964 17660
rect 10004 17620 14668 17660
rect 14708 17620 14717 17660
rect 0 17576 90 17596
rect 15244 17576 15284 17704
rect 15628 17660 15668 17704
rect 17932 17660 17972 17788
rect 18644 17788 18691 17819
rect 19084 17819 19276 17828
rect 18604 17744 18644 17779
rect 19124 17788 19276 17819
rect 19316 17788 19325 17828
rect 19084 17770 19124 17779
rect 18019 17704 18028 17744
rect 18068 17704 18124 17744
rect 18164 17704 18199 17744
rect 18595 17704 18604 17744
rect 18644 17704 18653 17744
rect 19529 17704 19660 17744
rect 19700 17704 19709 17744
rect 20009 17704 20140 17744
rect 20180 17704 20189 17744
rect 15628 17620 19180 17660
rect 19220 17620 19700 17660
rect 19660 17576 19700 17620
rect 21510 17576 21600 17596
rect 0 17536 1364 17576
rect 3043 17536 3052 17576
rect 3092 17536 4148 17576
rect 5587 17536 5596 17576
rect 5636 17536 6260 17576
rect 6355 17536 6364 17576
rect 6404 17536 7180 17576
rect 7220 17536 7229 17576
rect 10265 17536 10348 17576
rect 10388 17536 10396 17576
rect 10436 17536 10445 17576
rect 14009 17536 14092 17576
rect 14132 17536 14140 17576
rect 14180 17536 14189 17576
rect 14371 17536 14380 17576
rect 14420 17536 14620 17576
rect 14660 17536 14669 17576
rect 15244 17536 15380 17576
rect 15811 17536 15820 17576
rect 15860 17536 17020 17576
rect 17060 17536 17069 17576
rect 19306 17536 19315 17576
rect 19355 17536 19364 17576
rect 19411 17536 19420 17576
rect 19460 17536 19468 17576
rect 19508 17536 19591 17576
rect 19651 17536 19660 17576
rect 19700 17536 19709 17576
rect 20899 17536 20908 17576
rect 20948 17536 21600 17576
rect 0 17516 90 17536
rect 1324 17492 1364 17536
rect 1324 17452 3532 17492
rect 3572 17452 3581 17492
rect 4108 17408 4148 17536
rect 6220 17492 6260 17536
rect 15340 17492 15380 17536
rect 19324 17492 19364 17536
rect 21510 17516 21600 17536
rect 6220 17452 7084 17492
rect 7124 17452 7133 17492
rect 8707 17452 8716 17492
rect 8756 17452 15244 17492
rect 15284 17452 15293 17492
rect 15340 17452 19364 17492
rect 3679 17368 3688 17408
rect 3728 17368 3770 17408
rect 3810 17368 3852 17408
rect 3892 17368 3934 17408
rect 3974 17368 4016 17408
rect 4056 17368 4065 17408
rect 4108 17368 13324 17408
rect 13364 17368 13373 17408
rect 17740 17368 18124 17408
rect 18164 17368 18604 17408
rect 18644 17368 18653 17408
rect 18799 17368 18808 17408
rect 18848 17368 18890 17408
rect 18930 17368 18972 17408
rect 19012 17368 19054 17408
rect 19094 17368 19136 17408
rect 19176 17368 19185 17408
rect 17740 17324 17780 17368
rect 3331 17284 3340 17324
rect 3380 17284 4876 17324
rect 4916 17284 4925 17324
rect 6211 17284 6220 17324
rect 6260 17284 6508 17324
rect 6548 17284 6557 17324
rect 11011 17284 11020 17324
rect 11060 17284 17780 17324
rect 17827 17284 17836 17324
rect 17876 17284 18028 17324
rect 18068 17284 18077 17324
rect 0 17240 90 17260
rect 0 17200 4588 17240
rect 4628 17200 4637 17240
rect 6499 17200 6508 17240
rect 6548 17200 7276 17240
rect 7316 17200 7325 17240
rect 8009 17200 8140 17240
rect 8180 17200 8189 17240
rect 16675 17200 16684 17240
rect 16724 17200 16972 17240
rect 17012 17200 17021 17240
rect 17251 17200 17260 17240
rect 17300 17200 17308 17240
rect 17348 17200 17431 17240
rect 19171 17200 19180 17240
rect 19220 17200 19276 17240
rect 19316 17200 19351 17240
rect 19603 17200 19612 17240
rect 19652 17200 19756 17240
rect 19796 17200 19805 17240
rect 19852 17200 20044 17240
rect 20084 17200 20093 17240
rect 20371 17200 20380 17240
rect 20420 17200 21004 17240
rect 21044 17200 21053 17240
rect 0 17180 90 17200
rect 19852 17156 19892 17200
rect 2371 17116 2380 17156
rect 2420 17116 2668 17156
rect 2708 17116 2717 17156
rect 2851 17116 2860 17156
rect 2900 17116 2909 17156
rect 4195 17116 4204 17156
rect 4244 17116 8284 17156
rect 8324 17116 8333 17156
rect 10156 17116 10732 17156
rect 10772 17116 11404 17156
rect 11444 17116 11453 17156
rect 12643 17116 12652 17156
rect 12692 17116 16244 17156
rect 2860 17072 2900 17116
rect 2476 17032 3476 17072
rect 3523 17032 3532 17072
rect 3572 17032 4012 17072
rect 4052 17032 4061 17072
rect 6316 17032 7852 17072
rect 7892 17032 7901 17072
rect 8323 17032 8332 17072
rect 8372 17032 8524 17072
rect 8564 17032 8573 17072
rect 9353 17032 9484 17072
rect 9524 17032 9533 17072
rect 2476 16988 2516 17032
rect 3436 16988 3476 17032
rect 4108 16988 4148 16997
rect 6316 16988 6356 17032
rect 7948 16988 7988 16997
rect 10060 16988 10100 16997
rect 10156 16988 10196 17116
rect 10762 17032 10771 17072
rect 10811 17032 11116 17072
rect 11156 17032 11165 17072
rect 11491 17032 11500 17072
rect 11540 17032 12788 17072
rect 13603 17032 13612 17072
rect 13652 17032 14092 17072
rect 14132 17032 14141 17072
rect 12748 16988 12788 17032
rect 14668 16988 14708 16997
rect 16204 16988 16244 17116
rect 17548 17116 19700 17156
rect 17548 17072 17588 17116
rect 17539 17032 17548 17072
rect 17588 17032 17597 17072
rect 19363 17032 19372 17072
rect 19412 17032 19421 17072
rect 16780 16988 16820 16997
rect 18988 16988 19028 16997
rect 1097 16948 1228 16988
rect 1268 16948 1277 16988
rect 2851 16948 2860 16988
rect 2900 16948 3043 16988
rect 3083 16948 3092 16988
rect 3139 16948 3148 16988
rect 3188 16948 3197 16988
rect 3427 16948 3436 16988
rect 3476 16948 3485 16988
rect 3619 16948 3628 16988
rect 3668 16948 3799 16988
rect 4148 16948 4300 16988
rect 4340 16948 4349 16988
rect 4587 16948 4596 16988
rect 4636 16948 4645 16988
rect 4937 16948 5068 16988
rect 5108 16948 5117 16988
rect 6499 16948 6508 16988
rect 6548 16948 6700 16988
rect 6740 16948 6749 16988
rect 7459 16948 7468 16988
rect 7508 16948 7948 16988
rect 7988 16948 7997 16988
rect 8986 16948 8995 16988
rect 9035 16948 9044 16988
rect 9091 16948 9100 16988
rect 9140 16948 9271 16988
rect 9571 16948 9580 16988
rect 9620 16948 9868 16988
rect 9908 16948 9917 16988
rect 10100 16948 10196 16988
rect 10570 16948 10579 16988
rect 10619 16948 10732 16988
rect 10772 16948 10781 16988
rect 11491 16948 11500 16988
rect 11540 16948 12268 16988
rect 12308 16948 12317 16988
rect 12788 16948 12884 16988
rect 13594 16948 13603 16988
rect 13643 16948 13652 16988
rect 13699 16948 13708 16988
rect 13748 16948 13879 16988
rect 14153 16948 14188 16988
rect 14228 16948 14284 16988
rect 14324 16948 14333 16988
rect 14537 16948 14668 16988
rect 14708 16948 14717 16988
rect 15178 16948 15187 16988
rect 15227 16948 15284 16988
rect 15427 16948 15436 16988
rect 15476 16948 15532 16988
rect 15572 16948 15607 16988
rect 16204 16948 16780 16988
rect 17731 16948 17740 16988
rect 17780 16948 18316 16988
rect 18356 16948 18365 16988
rect 2476 16939 2516 16948
rect 0 16904 90 16924
rect 3148 16904 3188 16948
rect 4108 16939 4148 16948
rect 0 16864 1460 16904
rect 3148 16864 3820 16904
rect 3860 16864 3869 16904
rect 0 16844 90 16864
rect 1420 16820 1460 16864
rect 4588 16820 4628 16948
rect 6316 16939 6356 16948
rect 7948 16939 7988 16948
rect 1420 16780 4300 16820
rect 4340 16780 4349 16820
rect 4540 16780 4628 16820
rect 4684 16864 4916 16904
rect 1516 16612 4204 16652
rect 4244 16612 4253 16652
rect 0 16568 90 16588
rect 1516 16568 1556 16612
rect 4540 16568 4580 16780
rect 0 16528 1556 16568
rect 1603 16528 1612 16568
rect 1652 16528 2900 16568
rect 3715 16528 3724 16568
rect 3764 16528 4580 16568
rect 0 16508 90 16528
rect 2860 16484 2900 16528
rect 4684 16484 4724 16864
rect 4876 16820 4916 16864
rect 4771 16780 4780 16820
rect 4820 16780 4829 16820
rect 4876 16780 6604 16820
rect 6644 16780 6653 16820
rect 4780 16568 4820 16780
rect 4919 16612 4928 16652
rect 4968 16612 5010 16652
rect 5050 16612 5092 16652
rect 5132 16612 5174 16652
rect 5214 16612 5256 16652
rect 5296 16612 5305 16652
rect 4780 16528 6028 16568
rect 6068 16528 6077 16568
rect 9004 16484 9044 16948
rect 9100 16904 9140 16948
rect 10060 16939 10100 16948
rect 12748 16939 12788 16948
rect 9100 16864 9964 16904
rect 10004 16864 10013 16904
rect 12844 16820 12884 16948
rect 13612 16904 13652 16948
rect 14668 16939 14708 16948
rect 12931 16864 12940 16904
rect 12980 16864 13652 16904
rect 10243 16780 10252 16820
rect 10292 16780 10876 16820
rect 10916 16780 10925 16820
rect 12844 16780 14228 16820
rect 1459 16444 1468 16484
rect 1508 16444 1708 16484
rect 1748 16444 1757 16484
rect 2860 16444 4724 16484
rect 5443 16444 5452 16484
rect 5492 16444 6124 16484
rect 6164 16444 6173 16484
rect 7049 16444 7132 16484
rect 7172 16444 7180 16484
rect 7220 16444 7229 16484
rect 8899 16444 8908 16484
rect 8948 16444 9044 16484
rect 10505 16444 10636 16484
rect 10676 16444 10685 16484
rect 14188 16400 14228 16780
rect 15244 16484 15284 16948
rect 16780 16904 16820 16948
rect 18988 16904 19028 16948
rect 16780 16864 19028 16904
rect 19372 16820 19412 17032
rect 19660 16904 19700 17116
rect 19756 17116 19892 17156
rect 19987 17116 19996 17156
rect 20036 17116 21292 17156
rect 21332 17116 21341 17156
rect 19756 17072 19796 17116
rect 21510 17072 21600 17092
rect 19747 17032 19756 17072
rect 19796 17032 19805 17072
rect 20009 17032 20140 17072
rect 20180 17032 20189 17072
rect 21292 17032 21600 17072
rect 19660 16864 21196 16904
rect 21236 16864 21245 16904
rect 15331 16780 15340 16820
rect 15380 16780 16492 16820
rect 16532 16780 16541 16820
rect 19372 16780 20524 16820
rect 20564 16780 20573 16820
rect 21292 16736 21332 17032
rect 21510 17012 21600 17032
rect 19843 16696 19852 16736
rect 19892 16696 21332 16736
rect 20039 16612 20048 16652
rect 20088 16612 20130 16652
rect 20170 16612 20212 16652
rect 20252 16612 20294 16652
rect 20334 16612 20376 16652
rect 20416 16612 20425 16652
rect 21510 16568 21600 16588
rect 20995 16528 21004 16568
rect 21044 16528 21600 16568
rect 21510 16508 21600 16528
rect 14921 16444 15052 16484
rect 15092 16444 15101 16484
rect 15235 16444 15244 16484
rect 15284 16444 15293 16484
rect 16867 16444 16876 16484
rect 16916 16444 17116 16484
rect 17156 16444 17165 16484
rect 17827 16444 17836 16484
rect 17876 16444 17884 16484
rect 17924 16444 18007 16484
rect 19555 16444 19564 16484
rect 19604 16444 20140 16484
rect 20180 16444 20189 16484
rect 6595 16360 6604 16400
rect 6644 16360 6653 16400
rect 7939 16360 7948 16400
rect 7988 16360 10484 16400
rect 12643 16360 12652 16400
rect 12692 16360 13364 16400
rect 6604 16316 6644 16360
rect 1699 16276 1708 16316
rect 1748 16276 2380 16316
rect 2420 16276 2429 16316
rect 2947 16276 2956 16316
rect 2996 16276 3127 16316
rect 3331 16276 3340 16316
rect 3380 16276 3715 16316
rect 3755 16276 3764 16316
rect 3811 16276 3820 16316
rect 3860 16276 3991 16316
rect 4099 16276 4108 16316
rect 4148 16276 4204 16316
rect 4244 16276 4279 16316
rect 4780 16307 4972 16316
rect 2956 16258 2996 16267
rect 4820 16276 4972 16307
rect 5012 16276 5021 16316
rect 5129 16276 5260 16316
rect 5300 16276 5309 16316
rect 6316 16276 6644 16316
rect 7459 16276 7468 16316
rect 7508 16276 7517 16316
rect 8585 16276 8716 16316
rect 8756 16276 8765 16316
rect 9065 16276 9196 16316
rect 9236 16276 9245 16316
rect 10444 16307 10484 16360
rect 13324 16316 13364 16360
rect 13420 16360 13708 16400
rect 13748 16360 13757 16400
rect 14188 16360 15476 16400
rect 13420 16316 13460 16360
rect 4780 16258 4820 16267
rect 5260 16258 5300 16267
rect 0 16232 90 16252
rect 0 16192 268 16232
rect 308 16192 317 16232
rect 1027 16192 1036 16232
rect 1076 16192 1228 16232
rect 1268 16192 1277 16232
rect 3619 16192 3628 16232
rect 3668 16192 4300 16232
rect 4340 16192 4492 16232
rect 4532 16192 4541 16232
rect 5705 16192 5836 16232
rect 5876 16192 5885 16232
rect 6019 16192 6028 16232
rect 6068 16192 6220 16232
rect 6260 16192 6269 16232
rect 0 16172 90 16192
rect 6316 16148 6356 16276
rect 7468 16232 7508 16276
rect 8716 16258 8756 16267
rect 10627 16276 10636 16316
rect 10676 16276 11212 16316
rect 11252 16276 11261 16316
rect 12259 16276 12268 16316
rect 12308 16307 12500 16316
rect 12308 16276 12460 16307
rect 10444 16232 10484 16267
rect 13306 16276 13315 16316
rect 13355 16276 13364 16316
rect 13411 16276 13420 16316
rect 13460 16276 13469 16316
rect 13603 16276 13612 16316
rect 13652 16276 13804 16316
rect 13844 16276 13853 16316
rect 14345 16307 14476 16316
rect 14345 16276 14380 16307
rect 12460 16258 12500 16267
rect 13420 16232 13460 16276
rect 14420 16276 14476 16307
rect 14516 16276 14525 16316
rect 14729 16276 14860 16316
rect 14900 16276 14909 16316
rect 15436 16307 15476 16360
rect 17356 16360 19372 16400
rect 19412 16360 19421 16400
rect 14380 16258 14420 16267
rect 14860 16258 14900 16267
rect 16675 16276 16684 16316
rect 16724 16276 16972 16316
rect 17012 16276 17021 16316
rect 15436 16258 15476 16267
rect 17356 16232 17396 16360
rect 18115 16276 18124 16316
rect 18164 16276 18403 16316
rect 18443 16276 18452 16316
rect 18499 16276 18508 16316
rect 18548 16276 18679 16316
rect 18761 16276 18892 16316
rect 18932 16276 18941 16316
rect 19468 16307 19660 16316
rect 19508 16276 19660 16307
rect 19700 16276 19709 16316
rect 19948 16307 20524 16316
rect 19468 16258 19508 16267
rect 19988 16276 20524 16307
rect 20564 16276 20573 16316
rect 19948 16258 19988 16267
rect 6403 16192 6412 16232
rect 6452 16192 6604 16232
rect 6644 16192 6653 16232
rect 6857 16192 6892 16232
rect 6932 16192 6988 16232
rect 7028 16192 7037 16232
rect 7337 16192 7468 16232
rect 7508 16192 8620 16232
rect 8660 16192 8669 16232
rect 10444 16192 10828 16232
rect 10868 16192 12364 16232
rect 12404 16192 12413 16232
rect 12931 16192 12940 16232
rect 12980 16192 13460 16232
rect 13740 16192 13804 16232
rect 13844 16192 13900 16232
rect 13940 16192 14284 16232
rect 14324 16192 14333 16232
rect 17347 16192 17356 16232
rect 17396 16192 17405 16232
rect 17731 16192 17740 16232
rect 17780 16192 17789 16232
rect 18115 16192 18124 16232
rect 18164 16192 18173 16232
rect 18691 16192 18700 16232
rect 18740 16192 18988 16232
rect 19028 16192 19037 16232
rect 17740 16148 17780 16192
rect 18124 16148 18164 16192
rect 3139 16108 3148 16148
rect 3188 16108 3724 16148
rect 3764 16108 3773 16148
rect 4780 16108 6356 16148
rect 10627 16108 10636 16148
rect 10676 16108 16204 16148
rect 16244 16108 16253 16148
rect 17251 16108 17260 16148
rect 17300 16108 17500 16148
rect 17540 16108 17549 16148
rect 17740 16108 18068 16148
rect 18124 16108 20716 16148
rect 20756 16108 20765 16148
rect 4780 16064 4820 16108
rect 18028 16064 18068 16108
rect 21510 16064 21600 16084
rect 355 16024 364 16064
rect 404 16024 4820 16064
rect 5587 16024 5596 16064
rect 5636 16024 5644 16064
rect 5684 16024 5767 16064
rect 5971 16024 5980 16064
rect 6020 16024 6028 16064
rect 6068 16024 6151 16064
rect 6508 16024 6652 16064
rect 6692 16024 8716 16064
rect 8756 16024 8765 16064
rect 11059 16024 11068 16064
rect 11108 16024 12172 16064
rect 12212 16024 12221 16064
rect 15082 16024 15091 16064
rect 15131 16024 17836 16064
rect 17876 16024 17885 16064
rect 18028 16024 19948 16064
rect 19988 16024 19997 16064
rect 21379 16024 21388 16064
rect 21428 16024 21600 16064
rect 6508 15980 6548 16024
rect 21510 16004 21600 16024
rect 2563 15940 2572 15980
rect 2612 15940 6548 15980
rect 6595 15940 6604 15980
rect 6644 15940 6988 15980
rect 7028 15940 7037 15980
rect 7468 15940 10636 15980
rect 10676 15940 10685 15980
rect 0 15896 90 15916
rect 7468 15896 7508 15940
rect 0 15856 1324 15896
rect 1364 15856 1373 15896
rect 3679 15856 3688 15896
rect 3728 15856 3770 15896
rect 3810 15856 3852 15896
rect 3892 15856 3934 15896
rect 3974 15856 4016 15896
rect 4056 15856 4065 15896
rect 4291 15856 4300 15896
rect 4340 15856 5780 15896
rect 5827 15856 5836 15896
rect 5876 15856 7508 15896
rect 18799 15856 18808 15896
rect 18848 15856 18890 15896
rect 18930 15856 18972 15896
rect 19012 15856 19054 15896
rect 19094 15856 19136 15896
rect 19176 15856 19185 15896
rect 0 15836 90 15856
rect 5740 15728 5780 15856
rect 6892 15772 14380 15812
rect 14420 15772 14429 15812
rect 2633 15688 2764 15728
rect 2804 15688 2813 15728
rect 4553 15688 4684 15728
rect 4724 15688 4733 15728
rect 5740 15688 6652 15728
rect 6692 15688 6701 15728
rect 172 15604 4204 15644
rect 4244 15604 4253 15644
rect 4483 15604 4492 15644
rect 4532 15604 5260 15644
rect 5300 15604 5309 15644
rect 6595 15604 6604 15644
rect 6644 15604 6653 15644
rect 0 15560 90 15580
rect 172 15560 212 15604
rect 0 15520 212 15560
rect 6377 15520 6508 15560
rect 6548 15520 6557 15560
rect 0 15500 90 15520
rect 2572 15476 2612 15485
rect 4300 15476 4340 15485
rect 4876 15476 4916 15485
rect 6604 15476 6644 15604
rect 6892 15560 6932 15772
rect 6979 15688 6988 15728
rect 7028 15688 10348 15728
rect 10388 15688 10397 15728
rect 10601 15688 10732 15728
rect 10772 15688 10781 15728
rect 11020 15688 12460 15728
rect 12500 15688 12509 15728
rect 13219 15688 13228 15728
rect 13268 15688 13748 15728
rect 14563 15688 14572 15728
rect 14612 15688 14860 15728
rect 14900 15688 14909 15728
rect 17993 15688 18124 15728
rect 18164 15688 18173 15728
rect 11020 15644 11060 15688
rect 13708 15644 13748 15688
rect 7180 15604 9292 15644
rect 9332 15604 9341 15644
rect 10444 15604 11060 15644
rect 12451 15604 12460 15644
rect 12500 15604 12980 15644
rect 13708 15604 15092 15644
rect 16291 15604 16300 15644
rect 16340 15604 16436 15644
rect 7180 15560 7220 15604
rect 10444 15560 10484 15604
rect 6883 15520 6892 15560
rect 6932 15520 6941 15560
rect 7171 15520 7180 15560
rect 7220 15520 7229 15560
rect 9292 15520 10484 15560
rect 7180 15476 7220 15520
rect 8908 15476 8948 15485
rect 9292 15476 9332 15520
rect 10540 15476 10580 15485
rect 11020 15476 11060 15604
rect 12940 15560 12980 15604
rect 12355 15520 12364 15560
rect 12404 15520 12652 15560
rect 12692 15520 12701 15560
rect 12940 15520 14284 15560
rect 14324 15520 14333 15560
rect 12268 15476 12308 15485
rect 14380 15476 14420 15485
rect 15052 15476 15092 15604
rect 16300 15476 16340 15485
rect 16396 15476 16436 15604
rect 21510 15560 21600 15580
rect 18499 15520 18508 15560
rect 18548 15520 18892 15560
rect 18932 15520 18941 15560
rect 21187 15520 21196 15560
rect 21236 15520 21600 15560
rect 21510 15500 21600 15520
rect 17932 15476 17972 15485
rect 19468 15476 19508 15485
rect 355 15436 364 15476
rect 404 15436 1324 15476
rect 1364 15436 1373 15476
rect 2612 15436 2764 15476
rect 2804 15436 2813 15476
rect 3043 15436 3052 15476
rect 3092 15436 3628 15476
rect 3668 15436 3677 15476
rect 4169 15436 4300 15476
rect 4340 15436 4349 15476
rect 4916 15436 5740 15476
rect 5780 15436 5789 15476
rect 6115 15436 6124 15476
rect 6164 15436 6644 15476
rect 7171 15436 7180 15476
rect 7220 15436 7296 15476
rect 7529 15436 7660 15476
rect 7700 15436 7709 15476
rect 8777 15436 8908 15476
rect 8948 15436 8957 15476
rect 9004 15436 9292 15476
rect 9332 15436 9341 15476
rect 10580 15436 10676 15476
rect 11011 15436 11020 15476
rect 11060 15436 11069 15476
rect 12137 15436 12268 15476
rect 12308 15436 12317 15476
rect 13027 15436 13036 15476
rect 13076 15436 13132 15476
rect 13172 15436 13207 15476
rect 14179 15436 14188 15476
rect 14228 15436 14380 15476
rect 15043 15436 15052 15476
rect 15092 15436 15436 15476
rect 15476 15436 15485 15476
rect 16169 15436 16300 15476
rect 16340 15436 16349 15476
rect 16396 15436 16684 15476
rect 16724 15436 16972 15476
rect 17012 15436 17021 15476
rect 17443 15436 17452 15476
rect 17492 15436 17932 15476
rect 17972 15436 18124 15476
rect 18164 15436 18173 15476
rect 18394 15436 18403 15476
rect 18443 15436 18452 15476
rect 18499 15436 18508 15476
rect 18548 15436 18644 15476
rect 18691 15436 18700 15476
rect 18740 15436 18988 15476
rect 19028 15436 19037 15476
rect 19363 15436 19372 15476
rect 19412 15436 19468 15476
rect 19508 15436 19543 15476
rect 19978 15436 19987 15476
rect 20027 15436 20620 15476
rect 20660 15436 20669 15476
rect 2572 15427 2612 15436
rect 4300 15427 4340 15436
rect 4876 15427 4916 15436
rect 8908 15427 8948 15436
rect 3139 15268 3148 15308
rect 3188 15268 6268 15308
rect 6308 15268 6317 15308
rect 7411 15268 7420 15308
rect 7460 15268 8620 15308
rect 8660 15268 8669 15308
rect 0 15224 90 15244
rect 9004 15224 9044 15436
rect 10540 15427 10580 15436
rect 10636 15392 10676 15436
rect 12268 15392 12308 15436
rect 14380 15427 14420 15436
rect 16300 15427 16340 15436
rect 17932 15427 17972 15436
rect 18412 15392 18452 15436
rect 10627 15352 10636 15392
rect 10676 15352 10685 15392
rect 12268 15352 12892 15392
rect 12932 15352 13556 15392
rect 9091 15268 9100 15308
rect 9140 15268 9149 15308
rect 9283 15268 9292 15308
rect 9332 15268 13228 15308
rect 13268 15268 13277 15308
rect 0 15184 364 15224
rect 404 15184 413 15224
rect 7267 15184 7276 15224
rect 7316 15184 9044 15224
rect 9100 15224 9140 15268
rect 13516 15224 13556 15352
rect 16396 15352 17164 15392
rect 17204 15352 17213 15392
rect 18412 15352 18508 15392
rect 18548 15352 18557 15392
rect 9100 15184 9868 15224
rect 9908 15184 9917 15224
rect 13516 15184 14188 15224
rect 14228 15184 14237 15224
rect 0 15164 90 15184
rect 16396 15140 16436 15352
rect 18604 15308 18644 15436
rect 19468 15427 19508 15436
rect 16483 15268 16492 15308
rect 16532 15268 16541 15308
rect 17443 15268 17452 15308
rect 17492 15268 18220 15308
rect 18260 15268 18644 15308
rect 20131 15268 20140 15308
rect 20180 15268 20812 15308
rect 20852 15268 20861 15308
rect 4919 15100 4928 15140
rect 4968 15100 5010 15140
rect 5050 15100 5092 15140
rect 5132 15100 5174 15140
rect 5214 15100 5256 15140
rect 5296 15100 5305 15140
rect 9187 15100 9196 15140
rect 9236 15100 16436 15140
rect 3619 15016 3628 15056
rect 3668 15016 7412 15056
rect 9475 15016 9484 15056
rect 9524 15016 11636 15056
rect 13027 15016 13036 15056
rect 13076 15016 13996 15056
rect 14036 15016 14045 15056
rect 14092 15016 16436 15056
rect 7372 14972 7412 15016
rect 11596 14972 11636 15016
rect 14092 14972 14132 15016
rect 2851 14932 2860 14972
rect 2900 14932 3340 14972
rect 3380 14932 3389 14972
rect 4204 14932 4300 14972
rect 4340 14932 4349 14972
rect 7171 14932 7180 14972
rect 7220 14932 7229 14972
rect 7363 14932 7372 14972
rect 7412 14932 11060 14972
rect 11587 14932 11596 14972
rect 11636 14932 14132 14972
rect 14275 14932 14284 14972
rect 14324 14932 14420 14972
rect 14537 14932 14572 14972
rect 14612 14932 14668 14972
rect 14708 14932 14717 14972
rect 15139 14932 15148 14972
rect 15188 14932 15292 14972
rect 15332 14932 15341 14972
rect 0 14888 90 14908
rect 4204 14888 4244 14932
rect 0 14848 1516 14888
rect 1556 14848 1565 14888
rect 2860 14848 4244 14888
rect 4300 14848 5740 14888
rect 5780 14848 6988 14888
rect 7028 14848 7037 14888
rect 0 14828 90 14848
rect 2860 14804 2900 14848
rect 1219 14764 1228 14804
rect 1268 14764 1420 14804
rect 1460 14764 1996 14804
rect 2036 14764 2045 14804
rect 2668 14795 2900 14804
rect 2708 14764 2900 14795
rect 3043 14764 3052 14804
rect 3092 14764 3628 14804
rect 3668 14764 3677 14804
rect 4300 14795 4340 14848
rect 2668 14746 2708 14755
rect 3052 14636 3092 14764
rect 4553 14764 4684 14804
rect 4724 14764 4733 14804
rect 5932 14795 5972 14848
rect 7180 14804 7220 14932
rect 7747 14848 7756 14888
rect 7796 14848 8468 14888
rect 8803 14848 8812 14888
rect 8852 14848 8861 14888
rect 8428 14804 8468 14848
rect 8812 14804 8852 14848
rect 11020 14804 11060 14932
rect 4300 14746 4340 14755
rect 6307 14764 6316 14804
rect 6356 14764 7220 14804
rect 7276 14795 7604 14804
rect 7276 14764 7564 14795
rect 5932 14746 5972 14755
rect 7276 14636 7316 14764
rect 8410 14764 8419 14804
rect 8459 14764 8468 14804
rect 8515 14764 8524 14804
rect 8564 14764 8852 14804
rect 8899 14764 8908 14804
rect 8948 14764 9196 14804
rect 9236 14764 9245 14804
rect 9292 14764 9484 14804
rect 9524 14764 9533 14804
rect 9859 14764 9868 14804
rect 9908 14795 10039 14804
rect 9908 14764 9964 14795
rect 7564 14746 7604 14755
rect 8131 14680 8140 14720
rect 8180 14680 8189 14720
rect 8995 14680 9004 14720
rect 9044 14680 9053 14720
rect 1987 14596 1996 14636
rect 2036 14596 3092 14636
rect 4291 14596 4300 14636
rect 4340 14596 7316 14636
rect 0 14552 90 14572
rect 0 14512 2572 14552
rect 2612 14512 2621 14552
rect 4361 14512 4492 14552
rect 4532 14512 4541 14552
rect 6115 14512 6124 14552
rect 6164 14512 7084 14552
rect 7124 14512 7133 14552
rect 7180 14512 7900 14552
rect 7940 14512 7949 14552
rect 0 14492 90 14512
rect 3679 14344 3688 14384
rect 3728 14344 3770 14384
rect 3810 14344 3852 14384
rect 3892 14344 3934 14384
rect 3974 14344 4016 14384
rect 4056 14344 4065 14384
rect 3331 14260 3340 14300
rect 3380 14260 6220 14300
rect 6260 14260 6269 14300
rect 0 14216 90 14236
rect 7180 14216 7220 14512
rect 8140 14468 8180 14680
rect 9004 14552 9044 14680
rect 9292 14636 9332 14764
rect 9484 14746 9524 14755
rect 10004 14764 10039 14795
rect 11011 14764 11020 14804
rect 11060 14764 11069 14804
rect 12137 14764 12172 14804
rect 12212 14795 12308 14804
rect 12212 14764 12268 14795
rect 9964 14746 10004 14755
rect 12355 14764 12364 14804
rect 12404 14764 12835 14804
rect 12875 14764 12884 14804
rect 12931 14764 12940 14804
rect 12980 14764 13111 14804
rect 13315 14764 13324 14804
rect 13364 14764 13612 14804
rect 13652 14764 13661 14804
rect 13865 14795 13996 14804
rect 13865 14764 13900 14795
rect 12268 14746 12308 14755
rect 13940 14764 13996 14795
rect 14036 14764 14284 14804
rect 14324 14764 14333 14804
rect 14380 14795 14420 14932
rect 16090 14848 16099 14888
rect 16139 14848 16148 14888
rect 13900 14746 13940 14755
rect 14380 14746 14420 14755
rect 16108 14720 16148 14848
rect 16396 14804 16436 15016
rect 16492 14888 16532 15268
rect 16867 15100 16876 15140
rect 16916 15100 18412 15140
rect 18452 15100 18604 15140
rect 18644 15100 18653 15140
rect 20039 15100 20048 15140
rect 20088 15100 20130 15140
rect 20170 15100 20212 15140
rect 20252 15100 20294 15140
rect 20334 15100 20376 15140
rect 20416 15100 20425 15140
rect 21510 15056 21600 15076
rect 20803 15016 20812 15056
rect 20852 15016 21600 15056
rect 21510 14996 21600 15016
rect 18211 14932 18220 14972
rect 18260 14932 18268 14972
rect 18308 14932 18391 14972
rect 20131 14932 20140 14972
rect 20180 14932 20524 14972
rect 20564 14932 20573 14972
rect 16492 14848 17876 14888
rect 18115 14848 18124 14888
rect 18164 14848 19988 14888
rect 17836 14824 17876 14848
rect 16282 14764 16291 14804
rect 16331 14764 16340 14804
rect 16396 14795 16876 14804
rect 16396 14764 16780 14795
rect 10339 14680 10348 14720
rect 10388 14680 10636 14720
rect 10676 14680 10685 14720
rect 13411 14680 13420 14720
rect 13460 14680 13804 14720
rect 13844 14680 13853 14720
rect 15523 14680 15532 14720
rect 15572 14680 15581 14720
rect 15907 14680 15916 14720
rect 15956 14680 16148 14720
rect 15532 14636 15572 14680
rect 16300 14636 16340 14764
rect 16820 14764 16876 14795
rect 16916 14764 16925 14804
rect 17129 14764 17260 14804
rect 17300 14764 17309 14804
rect 17731 14764 17740 14804
rect 17780 14764 17789 14804
rect 17836 14784 17853 14824
rect 17893 14784 17902 14824
rect 18220 14764 18700 14804
rect 18740 14764 18749 14804
rect 19948 14795 19988 14848
rect 16780 14746 16820 14755
rect 17740 14720 17780 14764
rect 18220 14720 18260 14764
rect 19948 14746 19988 14755
rect 17155 14680 17164 14720
rect 17204 14680 17356 14720
rect 17396 14680 17405 14720
rect 17740 14680 18028 14720
rect 18068 14680 18077 14720
rect 18211 14680 18220 14720
rect 18260 14680 18269 14720
rect 18499 14680 18508 14720
rect 18548 14680 19852 14720
rect 19892 14680 19901 14720
rect 9283 14596 9292 14636
rect 9332 14596 9341 14636
rect 10147 14596 10156 14636
rect 10196 14596 10204 14636
rect 10244 14596 10327 14636
rect 10627 14596 10636 14636
rect 10676 14596 10876 14636
rect 10916 14596 15052 14636
rect 15092 14596 15101 14636
rect 15532 14596 16244 14636
rect 16300 14596 17356 14636
rect 17396 14596 17405 14636
rect 19660 14596 20812 14636
rect 20852 14596 20861 14636
rect 16204 14552 16244 14596
rect 19660 14552 19700 14596
rect 21510 14552 21600 14572
rect 9004 14512 10444 14552
rect 10484 14512 11020 14552
rect 11060 14512 11069 14552
rect 12329 14512 12460 14552
rect 12500 14512 12509 14552
rect 14371 14512 14380 14552
rect 14420 14512 15676 14552
rect 15716 14512 15725 14552
rect 16204 14512 19700 14552
rect 19747 14512 19756 14552
rect 19796 14512 21600 14552
rect 21510 14492 21600 14512
rect 8140 14428 16588 14468
rect 16628 14428 16637 14468
rect 8131 14344 8140 14384
rect 8180 14344 11404 14384
rect 11444 14344 11453 14384
rect 16003 14344 16012 14384
rect 16052 14344 17260 14384
rect 17300 14344 17309 14384
rect 18799 14344 18808 14384
rect 18848 14344 18890 14384
rect 18930 14344 18972 14384
rect 19012 14344 19054 14384
rect 19094 14344 19136 14384
rect 19176 14344 19185 14384
rect 7747 14260 7756 14300
rect 7796 14260 9620 14300
rect 9580 14216 9620 14260
rect 0 14176 7220 14216
rect 7459 14176 7468 14216
rect 7508 14176 9436 14216
rect 9476 14176 9485 14216
rect 9580 14176 10012 14216
rect 10052 14176 10061 14216
rect 12233 14176 12364 14216
rect 12404 14176 12413 14216
rect 13987 14176 13996 14216
rect 14036 14176 15628 14216
rect 15668 14176 15677 14216
rect 18377 14176 18508 14216
rect 18548 14176 18557 14216
rect 20227 14176 20236 14216
rect 20276 14176 20620 14216
rect 20660 14176 20669 14216
rect 0 14156 90 14176
rect 1769 14092 1852 14132
rect 1892 14092 1900 14132
rect 1940 14092 1949 14132
rect 2153 14092 2236 14132
rect 2276 14092 2284 14132
rect 2324 14092 2333 14132
rect 4723 14092 4732 14132
rect 4772 14092 10004 14132
rect 10339 14092 10348 14132
rect 10388 14092 10397 14132
rect 13481 14092 13612 14132
rect 13652 14092 14284 14132
rect 14324 14092 14333 14132
rect 14851 14092 14860 14132
rect 14900 14092 15764 14132
rect 163 14008 172 14048
rect 212 14008 1228 14048
rect 1268 14008 1277 14048
rect 1411 14008 1420 14048
rect 1460 14008 1612 14048
rect 1652 14008 1661 14048
rect 1987 14008 1996 14048
rect 2036 14008 2045 14048
rect 2371 14008 2380 14048
rect 2420 14008 2708 14048
rect 3043 14008 3052 14048
rect 3092 14008 3340 14048
rect 3380 14008 3389 14048
rect 4361 14008 4396 14048
rect 4436 14008 4492 14048
rect 4532 14008 4541 14048
rect 5059 14008 5068 14048
rect 5108 14008 5836 14048
rect 5876 14008 5885 14048
rect 6019 14008 6028 14048
rect 6068 14008 6220 14048
rect 6260 14008 6269 14048
rect 7363 14008 7372 14048
rect 7412 14008 7700 14048
rect 8035 14008 8044 14048
rect 8084 14008 8524 14048
rect 8564 14008 8573 14048
rect 9322 14008 9331 14048
rect 9371 14008 9676 14048
rect 9716 14008 9725 14048
rect 1996 13964 2036 14008
rect 2668 13964 2708 14008
rect 3628 13964 3668 13973
rect 6604 13964 6644 13973
rect 7660 13964 7700 14008
rect 8620 13964 8660 13973
rect 1123 13924 1132 13964
rect 1172 13924 2036 13964
rect 2554 13924 2563 13964
rect 2603 13924 2612 13964
rect 2659 13924 2668 13964
rect 2708 13924 2717 13964
rect 2851 13924 2860 13964
rect 2900 13924 3148 13964
rect 3188 13924 3197 13964
rect 3497 13924 3628 13964
rect 3668 13924 3677 13964
rect 3994 13924 4108 13964
rect 4156 13924 4174 13964
rect 4483 13924 4492 13964
rect 4532 13924 5539 13964
rect 5579 13924 5588 13964
rect 5635 13924 5644 13964
rect 5684 13924 5876 13964
rect 6115 13924 6124 13964
rect 6164 13924 6173 13964
rect 7075 13924 7084 13964
rect 7132 13924 7255 13964
rect 7546 13924 7555 13964
rect 7595 13924 7604 13964
rect 7651 13924 7660 13964
rect 7700 13924 7709 13964
rect 7843 13924 7852 13964
rect 7892 13924 7901 13964
rect 8009 13924 8140 13964
rect 8180 13924 8189 13964
rect 8986 13924 9100 13964
rect 9148 13924 9166 13964
rect 0 13880 90 13900
rect 2572 13880 2612 13924
rect 0 13840 76 13880
rect 116 13840 125 13880
rect 1459 13840 1468 13880
rect 1508 13840 2476 13880
rect 2516 13840 2525 13880
rect 2572 13840 2668 13880
rect 2708 13840 2717 13880
rect 0 13820 90 13840
rect 3148 13712 3188 13924
rect 3628 13915 3668 13924
rect 4579 13840 4588 13880
rect 4628 13840 4828 13880
rect 4868 13840 4877 13880
rect 5836 13796 5876 13924
rect 6124 13880 6164 13924
rect 5923 13840 5932 13880
rect 5972 13840 6164 13880
rect 4291 13756 4300 13796
rect 4340 13756 4492 13796
rect 4532 13756 4541 13796
rect 5827 13756 5836 13796
rect 5876 13756 5885 13796
rect 6604 13712 6644 13924
rect 7564 13880 7604 13924
rect 7852 13880 7892 13924
rect 8620 13880 8660 13924
rect 7564 13840 7660 13880
rect 7700 13840 7709 13880
rect 7852 13840 8660 13880
rect 7267 13756 7276 13796
rect 7316 13756 7852 13796
rect 7892 13756 7901 13796
rect 3148 13672 6644 13712
rect 9964 13712 10004 14092
rect 10348 14048 10388 14092
rect 13612 14048 13652 14092
rect 14284 14048 14324 14092
rect 10121 14008 10156 14048
rect 10196 14008 10252 14048
rect 10292 14008 10301 14048
rect 10348 14008 10540 14048
rect 10580 14008 10589 14048
rect 13603 14008 13612 14048
rect 13652 14008 13661 14048
rect 14284 14008 15284 14048
rect 15497 14008 15628 14048
rect 15668 14008 15677 14048
rect 12172 13964 12212 13973
rect 14188 13964 14228 13973
rect 15244 13964 15284 14008
rect 15724 13964 15764 14092
rect 21510 14048 21600 14068
rect 16483 14008 16492 14048
rect 16532 14008 16780 14048
rect 16820 14008 17108 14048
rect 16204 13964 16244 13973
rect 17068 13964 17108 14008
rect 18316 14008 20084 14048
rect 20803 14008 20812 14048
rect 20852 14008 21600 14048
rect 18316 13964 18356 14008
rect 20044 13964 20084 14008
rect 21510 13988 21600 14008
rect 10915 13924 10924 13964
rect 10964 13924 11404 13964
rect 11444 13924 11453 13964
rect 11587 13924 11596 13964
rect 11636 13924 12172 13964
rect 12212 13924 12221 13964
rect 12451 13924 12460 13964
rect 12500 13924 13123 13964
rect 13163 13924 13172 13964
rect 13219 13924 13228 13964
rect 13268 13924 13277 13964
rect 13673 13924 13708 13964
rect 13748 13924 13804 13964
rect 13844 13924 13853 13964
rect 13987 13924 13996 13964
rect 14036 13924 14188 13964
rect 12172 13915 12212 13924
rect 13228 13880 13268 13924
rect 14188 13915 14228 13924
rect 14380 13924 14676 13964
rect 14716 13924 14725 13964
rect 15130 13924 15139 13964
rect 15179 13924 15188 13964
rect 15235 13924 15244 13964
rect 15284 13924 15293 13964
rect 15715 13924 15724 13964
rect 15764 13924 15773 13964
rect 16073 13924 16204 13964
rect 16244 13924 16396 13964
rect 16436 13924 16445 13964
rect 16714 13924 16723 13964
rect 16763 13924 16876 13964
rect 16916 13924 16925 13964
rect 17059 13924 17068 13964
rect 17108 13924 17117 13964
rect 18115 13924 18124 13964
rect 18164 13924 18316 13964
rect 18787 13924 18796 13964
rect 18836 13924 18845 13964
rect 12931 13840 12940 13880
rect 12980 13840 13612 13880
rect 13652 13840 13661 13880
rect 10771 13756 10780 13796
rect 10820 13756 12748 13796
rect 12788 13756 12797 13796
rect 9964 13672 12980 13712
rect 4919 13588 4928 13628
rect 4968 13588 5010 13628
rect 5050 13588 5092 13628
rect 5132 13588 5174 13628
rect 5214 13588 5256 13628
rect 5296 13588 5305 13628
rect 5923 13588 5932 13628
rect 5972 13588 6124 13628
rect 6164 13588 12844 13628
rect 12884 13588 12893 13628
rect 0 13544 90 13564
rect 12940 13544 12980 13672
rect 0 13504 1804 13544
rect 1844 13504 1853 13544
rect 5347 13504 5356 13544
rect 5396 13504 5548 13544
rect 5588 13504 7276 13544
rect 7316 13504 7325 13544
rect 8611 13504 8620 13544
rect 8660 13504 11212 13544
rect 11252 13504 11261 13544
rect 12940 13504 13036 13544
rect 13076 13504 13085 13544
rect 0 13484 90 13504
rect 14380 13460 14420 13924
rect 15148 13880 15188 13924
rect 16204 13915 16244 13924
rect 18316 13915 18356 13924
rect 15148 13840 15244 13880
rect 15284 13840 15293 13880
rect 18796 13796 18836 13924
rect 20044 13915 20084 13924
rect 14851 13756 14860 13796
rect 14900 13756 15436 13796
rect 15476 13756 15485 13796
rect 16867 13756 16876 13796
rect 16916 13756 16925 13796
rect 17635 13756 17644 13796
rect 17684 13756 18836 13796
rect 1459 13420 1468 13460
rect 1508 13420 1612 13460
rect 1652 13420 1661 13460
rect 3043 13420 3052 13460
rect 3092 13420 3244 13460
rect 3284 13420 3293 13460
rect 3523 13420 3532 13460
rect 3572 13420 3580 13460
rect 3620 13420 3703 13460
rect 4291 13420 4300 13460
rect 4340 13420 5164 13460
rect 5204 13420 6068 13460
rect 7363 13420 7372 13460
rect 7412 13420 7421 13460
rect 14371 13420 14380 13460
rect 14420 13420 14429 13460
rect 15427 13420 15436 13460
rect 15476 13420 15484 13460
rect 15524 13420 15607 13460
rect 67 13336 76 13376
rect 116 13336 3148 13376
rect 3188 13336 3197 13376
rect 4108 13336 5932 13376
rect 5972 13336 5981 13376
rect 4108 13292 4148 13336
rect 6028 13292 6068 13420
rect 7372 13376 7412 13420
rect 16876 13376 16916 13756
rect 20039 13588 20048 13628
rect 20088 13588 20130 13628
rect 20170 13588 20212 13628
rect 20252 13588 20294 13628
rect 20334 13588 20376 13628
rect 20416 13588 20425 13628
rect 21510 13544 21600 13564
rect 16963 13504 16972 13544
rect 17012 13504 18700 13544
rect 18740 13504 18749 13544
rect 19267 13504 19276 13544
rect 19316 13504 21600 13544
rect 21510 13484 21600 13504
rect 17225 13420 17356 13460
rect 17396 13420 17405 13460
rect 17827 13420 17836 13460
rect 17876 13420 18740 13460
rect 19721 13420 19852 13460
rect 19892 13420 19901 13460
rect 20083 13420 20092 13460
rect 20132 13420 21292 13460
rect 21332 13420 21341 13460
rect 7372 13336 9620 13376
rect 10627 13336 10636 13376
rect 10676 13336 11252 13376
rect 16876 13336 17780 13376
rect 9580 13292 9620 13336
rect 11212 13292 11252 13336
rect 931 13252 940 13292
rect 980 13252 1268 13292
rect 1411 13252 1420 13292
rect 1460 13252 1612 13292
rect 1652 13252 1661 13292
rect 1891 13252 1900 13292
rect 1940 13283 2900 13292
rect 1940 13252 2860 13283
rect 0 13208 90 13228
rect 1228 13208 1268 13252
rect 2860 13234 2900 13243
rect 3244 13252 3436 13292
rect 3476 13252 3485 13292
rect 4099 13252 4108 13292
rect 4148 13252 4157 13292
rect 5356 13283 5396 13292
rect 3244 13208 3284 13252
rect 5539 13252 5548 13292
rect 5588 13252 5836 13292
rect 5876 13252 5885 13292
rect 6028 13283 7124 13292
rect 6028 13252 7084 13283
rect 5356 13208 5396 13243
rect 7363 13252 7372 13292
rect 7412 13252 8372 13292
rect 9571 13252 9580 13292
rect 9620 13252 9629 13292
rect 10697 13252 10828 13292
rect 10868 13252 10877 13292
rect 11203 13252 11212 13292
rect 11252 13252 11788 13292
rect 11828 13252 11837 13292
rect 12460 13283 12500 13292
rect 7084 13234 7124 13243
rect 8332 13208 8372 13252
rect 10828 13208 10868 13243
rect 12931 13252 12940 13292
rect 12980 13252 13132 13292
rect 13172 13252 13181 13292
rect 14057 13252 14188 13292
rect 14228 13252 14237 13292
rect 15907 13252 15916 13292
rect 15956 13252 16108 13292
rect 16148 13252 16157 13292
rect 16291 13252 16300 13292
rect 16340 13252 16684 13292
rect 16724 13283 17204 13292
rect 16724 13252 17164 13283
rect 12460 13208 12500 13243
rect 14188 13234 14228 13243
rect 17164 13234 17204 13243
rect 17740 13208 17780 13336
rect 18124 13336 18316 13376
rect 18356 13336 18365 13376
rect 18124 13292 18164 13336
rect 18106 13252 18115 13292
rect 18155 13252 18164 13292
rect 18211 13252 18220 13292
rect 18260 13252 18269 13292
rect 18403 13252 18412 13292
rect 18452 13252 18604 13292
rect 18644 13252 18653 13292
rect 18220 13208 18260 13252
rect 18700 13208 18740 13420
rect 19180 13283 19220 13292
rect 19529 13252 19660 13292
rect 19700 13252 19709 13292
rect 0 13168 1172 13208
rect 1219 13168 1228 13208
rect 1268 13168 1277 13208
rect 3235 13168 3244 13208
rect 3284 13168 3293 13208
rect 3436 13168 3668 13208
rect 3811 13168 3820 13208
rect 3860 13168 5260 13208
rect 5300 13168 5309 13208
rect 5356 13168 6316 13208
rect 6356 13168 6365 13208
rect 7276 13168 7660 13208
rect 7700 13168 7709 13208
rect 7843 13168 7852 13208
rect 7892 13168 7948 13208
rect 7988 13168 8023 13208
rect 8323 13168 8332 13208
rect 8372 13168 8381 13208
rect 8707 13168 8716 13208
rect 8756 13168 10444 13208
rect 10484 13168 10493 13208
rect 10828 13168 12500 13208
rect 15715 13168 15724 13208
rect 15764 13168 16972 13208
rect 17012 13168 17021 13208
rect 17731 13168 17740 13208
rect 17780 13168 17789 13208
rect 18115 13168 18124 13208
rect 18164 13168 18260 13208
rect 18691 13168 18700 13208
rect 18740 13168 18749 13208
rect 0 13148 90 13168
rect 1132 13124 1172 13168
rect 3436 13124 3476 13168
rect 1132 13084 3476 13124
rect 3628 13124 3668 13168
rect 7276 13124 7316 13168
rect 19180 13124 19220 13243
rect 19660 13234 19700 13243
rect 20323 13168 20332 13208
rect 20372 13168 20908 13208
rect 20948 13168 20957 13208
rect 3628 13084 5684 13124
rect 7267 13084 7276 13124
rect 7316 13084 7325 13124
rect 7372 13084 8092 13124
rect 8132 13084 8141 13124
rect 11491 13084 11500 13124
rect 11540 13084 17500 13124
rect 17540 13084 17549 13124
rect 17644 13084 19220 13124
rect 5644 13040 5684 13084
rect 7372 13040 7412 13084
rect 1411 13000 1420 13040
rect 1460 13000 1708 13040
rect 1748 13000 1757 13040
rect 2851 13000 2860 13040
rect 2900 13000 3484 13040
rect 3524 13000 4300 13040
rect 4340 13000 4349 13040
rect 5417 13000 5548 13040
rect 5588 13000 5597 13040
rect 5644 13000 7412 13040
rect 7577 13000 7660 13040
rect 7700 13000 7708 13040
rect 7748 13000 7757 13040
rect 7852 13000 8476 13040
rect 8516 13000 8525 13040
rect 11011 13000 11020 13040
rect 11060 13000 11788 13040
rect 11828 13000 11837 13040
rect 12643 13000 12652 13040
rect 12692 13000 13420 13040
rect 13460 13000 13469 13040
rect 16579 13000 16588 13040
rect 16628 13000 17356 13040
rect 17396 13000 17405 13040
rect 7852 12956 7892 13000
rect 17644 12956 17684 13084
rect 21510 13040 21600 13060
rect 20899 13000 20908 13040
rect 20948 13000 21600 13040
rect 21510 12980 21600 13000
rect 643 12916 652 12956
rect 692 12916 7892 12956
rect 8044 12916 14996 12956
rect 17251 12916 17260 12956
rect 17300 12916 17684 12956
rect 0 12872 90 12892
rect 0 12832 76 12872
rect 116 12832 125 12872
rect 3679 12832 3688 12872
rect 3728 12832 3770 12872
rect 3810 12832 3852 12872
rect 3892 12832 3934 12872
rect 3974 12832 4016 12872
rect 4056 12832 4065 12872
rect 0 12812 90 12832
rect 8044 12788 8084 12916
rect 14956 12872 14996 12916
rect 8515 12832 8524 12872
rect 8564 12832 14764 12872
rect 14804 12832 14813 12872
rect 14956 12832 17452 12872
rect 17492 12832 17501 12872
rect 18799 12832 18808 12872
rect 18848 12832 18890 12872
rect 18930 12832 18972 12872
rect 19012 12832 19054 12872
rect 19094 12832 19136 12872
rect 19176 12832 19185 12872
rect 2236 12748 8084 12788
rect 8131 12748 8140 12788
rect 8180 12748 15820 12788
rect 15860 12748 15869 12788
rect 17260 12748 18644 12788
rect 18691 12748 18700 12788
rect 18740 12748 21140 12788
rect 2236 12704 2276 12748
rect 2227 12664 2236 12704
rect 2276 12664 2285 12704
rect 5251 12664 5260 12704
rect 5300 12664 7228 12704
rect 7268 12664 7277 12704
rect 7843 12664 7852 12704
rect 7892 12664 14380 12704
rect 14420 12664 14429 12704
rect 15113 12664 15244 12704
rect 15284 12664 15293 12704
rect 16745 12664 16876 12704
rect 16916 12664 16925 12704
rect 163 12580 172 12620
rect 212 12580 7612 12620
rect 7652 12580 7661 12620
rect 8035 12580 8044 12620
rect 8084 12580 8524 12620
rect 8564 12580 8573 12620
rect 8899 12580 8908 12620
rect 8948 12580 8957 12620
rect 9763 12580 9772 12620
rect 9812 12580 12076 12620
rect 12116 12580 12125 12620
rect 12364 12580 13516 12620
rect 13556 12580 13565 12620
rect 16963 12580 16972 12620
rect 17012 12580 17020 12620
rect 17060 12580 17143 12620
rect 0 12536 90 12556
rect 8908 12536 8948 12580
rect 12364 12536 12404 12580
rect 17260 12536 17300 12748
rect 18604 12704 18644 12748
rect 17347 12664 17356 12704
rect 17396 12664 17404 12704
rect 17444 12664 17527 12704
rect 18604 12664 19852 12704
rect 19892 12664 19901 12704
rect 17644 12580 19276 12620
rect 19316 12580 19325 12620
rect 17644 12536 17684 12580
rect 21100 12536 21140 12748
rect 21510 12536 21600 12556
rect 0 12496 652 12536
rect 692 12496 701 12536
rect 835 12496 844 12536
rect 884 12496 1228 12536
rect 1268 12496 1277 12536
rect 1603 12496 1612 12536
rect 1652 12496 1661 12536
rect 1987 12496 1996 12536
rect 2036 12496 2045 12536
rect 2371 12496 2380 12536
rect 2420 12496 2612 12536
rect 2947 12496 2956 12536
rect 2996 12496 3052 12536
rect 3092 12496 3127 12536
rect 3532 12496 3724 12536
rect 3764 12496 3773 12536
rect 4265 12496 4300 12536
rect 4340 12496 4396 12536
rect 4436 12496 4445 12536
rect 4627 12496 4636 12536
rect 4676 12496 4876 12536
rect 4916 12496 4925 12536
rect 5033 12496 5116 12536
rect 5156 12496 5164 12536
rect 5204 12496 5213 12536
rect 5356 12496 5548 12536
rect 5588 12496 5597 12536
rect 5705 12496 5836 12536
rect 5876 12496 5885 12536
rect 6412 12496 6604 12536
rect 6644 12496 6653 12536
rect 7114 12496 7123 12536
rect 7163 12496 7468 12536
rect 7508 12496 7517 12536
rect 7721 12496 7852 12536
rect 7892 12496 7901 12536
rect 8419 12496 8428 12536
rect 8468 12496 9196 12536
rect 9236 12496 9245 12536
rect 11779 12496 11788 12536
rect 11828 12496 11837 12536
rect 12355 12496 12364 12536
rect 12404 12496 12413 12536
rect 12460 12496 12844 12536
rect 12884 12496 12893 12536
rect 17251 12496 17260 12536
rect 17300 12496 17309 12536
rect 17635 12496 17644 12536
rect 17684 12496 17693 12536
rect 18281 12496 18412 12536
rect 18452 12496 18461 12536
rect 18595 12496 18604 12536
rect 18644 12496 18653 12536
rect 20323 12496 20332 12536
rect 20372 12496 21004 12536
rect 21044 12496 21053 12536
rect 21100 12496 21600 12536
rect 0 12476 90 12496
rect 1612 12452 1652 12496
rect 451 12412 460 12452
rect 500 12412 1652 12452
rect 1996 12368 2036 12496
rect 2572 12452 2612 12496
rect 3532 12452 3572 12496
rect 5356 12452 5396 12496
rect 6412 12452 6452 12496
rect 9868 12452 9908 12461
rect 11788 12452 11828 12496
rect 12460 12452 12500 12496
rect 12940 12452 12980 12461
rect 15052 12452 15092 12461
rect 16684 12452 16724 12461
rect 18604 12452 18644 12496
rect 21510 12476 21600 12496
rect 18988 12452 19028 12461
rect 2458 12412 2467 12452
rect 2507 12412 2516 12452
rect 2563 12412 2572 12452
rect 2612 12412 2621 12452
rect 3043 12412 3052 12452
rect 3092 12412 3244 12452
rect 3284 12412 3293 12452
rect 3619 12412 3628 12452
rect 3668 12412 4020 12452
rect 4060 12412 4069 12452
rect 5338 12412 5347 12452
rect 5387 12412 5396 12452
rect 5443 12412 5452 12452
rect 5492 12412 5684 12452
rect 5923 12412 5932 12452
rect 5972 12412 6124 12452
rect 6164 12412 6173 12452
rect 6895 12451 6904 12452
rect 739 12328 748 12368
rect 788 12328 2036 12368
rect 2476 12368 2516 12412
rect 3532 12403 3572 12412
rect 2476 12328 2572 12368
rect 2612 12328 2621 12368
rect 5644 12284 5684 12412
rect 6412 12403 6452 12412
rect 6892 12412 6904 12451
rect 6944 12412 6953 12452
rect 8611 12412 8620 12452
rect 8660 12412 9004 12452
rect 9044 12412 9053 12452
rect 9737 12412 9868 12452
rect 9908 12412 9917 12452
rect 11788 12412 11854 12452
rect 11894 12412 11903 12452
rect 11968 12412 11977 12452
rect 12017 12412 12076 12452
rect 12116 12412 12157 12452
rect 12329 12412 12460 12452
rect 12500 12412 12509 12452
rect 12809 12412 12940 12452
rect 12980 12412 12989 12452
rect 13411 12412 13420 12452
rect 13468 12412 13591 12452
rect 13795 12412 13804 12452
rect 13844 12412 14764 12452
rect 14804 12412 14813 12452
rect 14921 12412 15052 12452
rect 15092 12412 15188 12452
rect 15305 12412 15436 12452
rect 15476 12412 15485 12452
rect 15619 12412 15628 12452
rect 15668 12412 16684 12452
rect 16724 12412 16733 12452
rect 17771 12412 17836 12452
rect 17876 12412 17902 12452
rect 17942 12412 17951 12452
rect 18019 12412 18028 12452
rect 18068 12412 18124 12452
rect 18164 12412 18228 12452
rect 18377 12412 18508 12452
rect 18548 12412 18557 12452
rect 18604 12412 18988 12452
rect 19363 12412 19372 12452
rect 19412 12412 19476 12452
rect 19516 12412 19543 12452
rect 6892 12411 6949 12412
rect 6892 12368 6932 12411
rect 9868 12403 9908 12412
rect 12940 12403 12980 12412
rect 15052 12403 15092 12412
rect 6595 12328 6604 12368
rect 6644 12328 6932 12368
rect 15148 12368 15188 12412
rect 16684 12403 16724 12412
rect 18028 12368 18068 12412
rect 18988 12403 19028 12412
rect 15148 12328 16340 12368
rect 17443 12328 17452 12368
rect 17492 12328 18068 12368
rect 19084 12328 20092 12368
rect 20132 12328 20141 12368
rect 16300 12284 16340 12328
rect 19084 12284 19124 12328
rect 1459 12244 1468 12284
rect 1508 12244 1748 12284
rect 1843 12244 1852 12284
rect 1892 12244 2764 12284
rect 2804 12244 2813 12284
rect 4195 12244 4204 12284
rect 4244 12244 4300 12284
rect 4340 12244 4375 12284
rect 5155 12244 5164 12284
rect 5204 12244 5548 12284
rect 5588 12244 5597 12284
rect 5644 12244 5932 12284
rect 5972 12244 6124 12284
rect 6164 12244 6173 12284
rect 8057 12244 8140 12284
rect 8180 12244 8188 12284
rect 8228 12244 8237 12284
rect 10051 12244 10060 12284
rect 10100 12244 10231 12284
rect 13603 12244 13612 12284
rect 13652 12244 16204 12284
rect 16244 12244 16253 12284
rect 16300 12244 17164 12284
rect 17204 12244 17213 12284
rect 18220 12244 19124 12284
rect 19651 12244 19660 12284
rect 19700 12244 19709 12284
rect 0 12200 90 12220
rect 1708 12200 1748 12244
rect 0 12160 748 12200
rect 788 12160 797 12200
rect 1708 12160 6412 12200
rect 6452 12160 6461 12200
rect 9187 12160 9196 12200
rect 9236 12160 16108 12200
rect 16148 12160 16157 12200
rect 16483 12160 16492 12200
rect 16532 12160 16972 12200
rect 17012 12160 17021 12200
rect 0 12140 90 12160
rect 1804 12076 4588 12116
rect 4628 12076 4637 12116
rect 4919 12076 4928 12116
rect 4968 12076 5010 12116
rect 5050 12076 5092 12116
rect 5132 12076 5174 12116
rect 5214 12076 5256 12116
rect 5296 12076 5305 12116
rect 547 11908 556 11948
rect 596 11908 1180 11948
rect 1220 11908 1229 11948
rect 1481 11908 1564 11948
rect 1604 11908 1612 11948
rect 1652 11908 1661 11948
rect 0 11864 90 11884
rect 0 11824 940 11864
rect 980 11824 989 11864
rect 0 11804 90 11824
rect 1804 11696 1844 12076
rect 18220 12032 18260 12244
rect 2188 11992 4684 12032
rect 4724 11992 4733 12032
rect 7267 11992 7276 12032
rect 7316 11992 9236 12032
rect 12931 11992 12940 12032
rect 12980 11992 14188 12032
rect 14228 11992 14237 12032
rect 14947 11992 14956 12032
rect 14996 11992 18260 12032
rect 2188 11780 2228 11992
rect 9196 11948 9236 11992
rect 3619 11908 3628 11948
rect 3668 11908 4108 11948
rect 4148 11908 4157 11948
rect 4291 11908 4300 11948
rect 4340 11908 4349 11948
rect 6499 11908 6508 11948
rect 6548 11908 6604 11948
rect 6644 11908 6679 11948
rect 8419 11908 8428 11948
rect 8468 11908 9100 11948
rect 9140 11908 9149 11948
rect 9196 11908 16444 11948
rect 16484 11908 16493 11948
rect 16588 11908 17452 11948
rect 17492 11908 17501 11948
rect 18185 11908 18316 11948
rect 18356 11908 18365 11948
rect 4300 11864 4340 11908
rect 16588 11864 16628 11908
rect 19660 11864 19700 12244
rect 20039 12076 20048 12116
rect 20088 12076 20130 12116
rect 20170 12076 20212 12116
rect 20252 12076 20294 12116
rect 20334 12076 20376 12116
rect 20416 12076 20425 12116
rect 21510 12032 21600 12052
rect 20995 11992 21004 12032
rect 21044 11992 21600 12032
rect 21510 11972 21600 11992
rect 3763 11824 3772 11864
rect 3812 11824 4012 11864
rect 4052 11824 4061 11864
rect 4300 11824 4916 11864
rect 4963 11824 4972 11864
rect 5012 11824 8044 11864
rect 8084 11824 8093 11864
rect 9283 11824 9292 11864
rect 9332 11824 9812 11864
rect 10051 11824 10060 11864
rect 10100 11824 10292 11864
rect 13123 11824 13132 11864
rect 13172 11824 13181 11864
rect 14371 11824 14380 11864
rect 14420 11824 14516 11864
rect 14659 11824 14668 11864
rect 14708 11824 15436 11864
rect 15476 11824 15485 11864
rect 16339 11824 16348 11864
rect 16388 11824 16628 11864
rect 16684 11824 19700 11864
rect 19843 11824 19852 11864
rect 19892 11824 20092 11864
rect 20132 11824 20141 11864
rect 2179 11740 2188 11780
rect 2228 11740 2237 11780
rect 2851 11740 2860 11780
rect 2900 11771 3480 11780
rect 2900 11740 3440 11771
rect 3440 11722 3480 11731
rect 4012 11740 4820 11780
rect 4012 11696 4052 11740
rect 1411 11656 1420 11696
rect 1460 11656 1469 11696
rect 1795 11656 1804 11696
rect 1844 11656 1853 11696
rect 4003 11656 4012 11696
rect 4052 11656 4061 11696
rect 4361 11656 4492 11696
rect 4532 11656 4541 11696
rect 1420 11612 1460 11656
rect 4780 11612 4820 11740
rect 4876 11696 4916 11824
rect 9772 11780 9812 11824
rect 5059 11740 5068 11780
rect 5108 11740 5740 11780
rect 5780 11740 5789 11780
rect 6185 11740 6316 11780
rect 6356 11740 6365 11780
rect 6499 11740 6508 11780
rect 6548 11740 6988 11780
rect 7028 11740 7037 11780
rect 8131 11740 8140 11780
rect 8180 11771 8311 11780
rect 8180 11740 8236 11771
rect 6316 11722 6356 11731
rect 8276 11740 8311 11771
rect 8515 11740 8524 11780
rect 8564 11740 8707 11780
rect 8747 11740 8756 11780
rect 8803 11740 8812 11780
rect 8852 11740 8983 11780
rect 9187 11740 9196 11780
rect 9236 11740 9388 11780
rect 9428 11740 9437 11780
rect 9641 11740 9772 11780
rect 9812 11740 9821 11780
rect 10252 11771 10292 11824
rect 13132 11780 13172 11824
rect 8236 11722 8276 11731
rect 9772 11722 9812 11731
rect 11561 11740 11692 11780
rect 11732 11740 11741 11780
rect 12809 11740 12940 11780
rect 12980 11740 12989 11780
rect 13132 11740 13411 11780
rect 13451 11740 13460 11780
rect 13507 11740 13516 11780
rect 13556 11740 13687 11780
rect 13795 11740 13804 11780
rect 13844 11740 13900 11780
rect 13940 11740 13975 11780
rect 14476 11771 14516 11824
rect 10252 11722 10292 11731
rect 12940 11722 12980 11731
rect 14825 11740 14956 11780
rect 14996 11740 15005 11780
rect 14476 11722 14516 11731
rect 14956 11722 14996 11731
rect 16684 11696 16724 11824
rect 16841 11740 16876 11780
rect 16916 11740 16972 11780
rect 17012 11740 17021 11780
rect 17155 11740 17164 11780
rect 17204 11771 18164 11780
rect 17204 11740 18124 11771
rect 18377 11740 18508 11780
rect 18548 11740 18557 11780
rect 19756 11771 19796 11780
rect 18124 11696 18164 11731
rect 19756 11696 19796 11731
rect 4867 11656 4876 11696
rect 4916 11656 4925 11696
rect 9161 11656 9292 11696
rect 9332 11656 9341 11696
rect 10474 11656 10483 11696
rect 10523 11656 10828 11696
rect 10868 11656 10877 11696
rect 13987 11656 13996 11696
rect 14036 11656 14380 11696
rect 14420 11656 14429 11696
rect 15178 11656 15187 11696
rect 15227 11656 15532 11696
rect 15572 11656 15581 11696
rect 15977 11656 16108 11696
rect 16148 11656 16628 11696
rect 16675 11656 16684 11696
rect 16724 11656 16733 11696
rect 18124 11656 19796 11696
rect 20323 11656 20332 11696
rect 20372 11656 21388 11696
rect 21428 11656 21437 11696
rect 16588 11612 16628 11656
rect 1420 11572 2860 11612
rect 2900 11572 2909 11612
rect 2956 11572 4252 11612
rect 4292 11572 4301 11612
rect 4387 11572 4396 11612
rect 4436 11572 4636 11612
rect 4676 11572 4685 11612
rect 4780 11572 15292 11612
rect 15332 11572 15341 11612
rect 16588 11572 18700 11612
rect 18740 11572 18749 11612
rect 19651 11572 19660 11612
rect 19700 11572 19948 11612
rect 19988 11572 19997 11612
rect 0 11528 90 11548
rect 0 11488 1996 11528
rect 2036 11488 2045 11528
rect 0 11468 90 11488
rect 2956 11444 2996 11572
rect 21510 11528 21600 11548
rect 2371 11404 2380 11444
rect 2420 11404 2996 11444
rect 9484 11488 10292 11528
rect 10339 11488 10348 11528
rect 10388 11488 10588 11528
rect 10628 11488 10637 11528
rect 10723 11488 10732 11528
rect 10772 11488 16972 11528
rect 17012 11488 17021 11528
rect 17635 11488 17644 11528
rect 17684 11488 18124 11528
rect 18164 11488 18508 11528
rect 18548 11488 18557 11528
rect 20716 11488 21600 11528
rect 3679 11320 3688 11360
rect 3728 11320 3770 11360
rect 3810 11320 3852 11360
rect 3892 11320 3934 11360
rect 3974 11320 4016 11360
rect 4056 11320 4065 11360
rect 1228 11236 1900 11276
rect 1940 11236 3284 11276
rect 0 11192 90 11212
rect 0 11152 460 11192
rect 500 11152 509 11192
rect 0 11132 90 11152
rect 1228 10940 1268 11236
rect 2537 11152 2668 11192
rect 2708 11152 2717 11192
rect 1315 11068 1324 11108
rect 1364 11068 2812 11108
rect 2852 11068 2861 11108
rect 3244 11024 3284 11236
rect 3427 11152 3436 11192
rect 3476 11152 3484 11192
rect 3524 11152 3607 11192
rect 3820 11152 6412 11192
rect 6452 11152 6461 11192
rect 8035 11152 8044 11192
rect 8084 11152 8524 11192
rect 8564 11152 8573 11192
rect 3820 11024 3860 11152
rect 9484 11108 9524 11488
rect 10252 11444 10292 11488
rect 17644 11444 17684 11488
rect 20716 11444 20756 11488
rect 21510 11468 21600 11488
rect 10252 11404 11692 11444
rect 11732 11404 15340 11444
rect 15380 11404 15389 11444
rect 15811 11404 15820 11444
rect 15860 11404 17684 11444
rect 20035 11404 20044 11444
rect 20084 11404 20756 11444
rect 4012 11068 9524 11108
rect 4012 11024 4052 11068
rect 2921 10984 2956 11024
rect 2996 10984 3052 11024
rect 3092 10984 3101 11024
rect 3235 10984 3244 11024
rect 3284 10984 3293 11024
rect 3811 10984 3820 11024
rect 3860 10984 3869 11024
rect 4003 10984 4012 11024
rect 4052 10984 4061 11024
rect 6403 10984 6412 11024
rect 6452 10984 6604 11024
rect 6644 10984 6653 11024
rect 7180 10984 7372 11024
rect 7412 10984 7948 11024
rect 7988 10984 7997 11024
rect 2476 10940 2516 10949
rect 5644 10940 5684 10949
rect 7180 10940 7220 10984
rect 8236 10940 8276 10949
rect 9484 10940 9524 11068
rect 9772 11320 13996 11360
rect 14036 11320 14045 11360
rect 14188 11320 18316 11360
rect 18356 11320 18365 11360
rect 18799 11320 18808 11360
rect 18848 11320 18890 11360
rect 18930 11320 18972 11360
rect 19012 11320 19054 11360
rect 19094 11320 19136 11360
rect 19176 11320 19185 11360
rect 9772 10940 9812 11320
rect 14188 11276 14228 11320
rect 9859 11236 9868 11276
rect 9908 11236 11788 11276
rect 11828 11236 11837 11276
rect 12940 11236 14228 11276
rect 14284 11236 17740 11276
rect 17780 11236 17789 11276
rect 11020 11152 11500 11192
rect 11540 11152 11884 11192
rect 11924 11152 11933 11192
rect 11020 10940 11060 11152
rect 12940 11108 12980 11236
rect 11980 11068 12980 11108
rect 11980 11024 12020 11068
rect 1219 10900 1228 10940
rect 1268 10900 1277 10940
rect 2516 10900 2764 10940
rect 2804 10900 2813 10940
rect 4387 10900 4396 10940
rect 4436 10900 5356 10940
rect 5396 10900 5405 10940
rect 2476 10891 2516 10900
rect 0 10856 90 10876
rect 0 10816 1612 10856
rect 1652 10816 1661 10856
rect 2668 10816 2900 10856
rect 0 10796 90 10816
rect 2668 10772 2708 10816
rect 2467 10732 2476 10772
rect 2516 10732 2708 10772
rect 2860 10772 2900 10816
rect 5644 10772 5684 10900
rect 5836 10900 6115 10940
rect 6155 10900 6164 10940
rect 6211 10900 6220 10940
rect 6260 10900 6269 10940
rect 6569 10900 6700 10940
rect 6740 10900 6749 10940
rect 7690 10900 7699 10940
rect 7739 10900 8044 10940
rect 8084 10900 8093 10940
rect 9475 10900 9484 10940
rect 9524 10900 9533 10940
rect 9763 10900 9772 10940
rect 9812 10900 9821 10940
rect 5836 10856 5876 10900
rect 6220 10856 6260 10900
rect 7180 10891 7220 10900
rect 8236 10856 8276 10900
rect 11020 10891 11060 10900
rect 11116 10984 11980 11024
rect 12020 10984 12029 11024
rect 12652 10984 13652 11024
rect 5827 10816 5836 10856
rect 5876 10816 5885 10856
rect 6060 10816 6124 10856
rect 6164 10816 6892 10856
rect 6932 10816 6941 10856
rect 7612 10816 9868 10856
rect 9908 10816 9917 10856
rect 7612 10772 7652 10816
rect 2860 10732 3580 10772
rect 3620 10732 3629 10772
rect 4243 10732 4252 10772
rect 4292 10732 4300 10772
rect 4340 10732 4423 10772
rect 5644 10732 7564 10772
rect 7604 10732 7652 10772
rect 7721 10732 7852 10772
rect 7892 10732 7901 10772
rect 8515 10732 8524 10772
rect 8564 10732 10252 10772
rect 10292 10732 10301 10772
rect 11116 10688 11156 10984
rect 12556 10940 12596 10949
rect 11482 10900 11491 10940
rect 11531 10900 11540 10940
rect 11587 10900 11596 10940
rect 11636 10900 11645 10940
rect 12067 10900 12076 10940
rect 12116 10900 12460 10940
rect 12500 10900 12509 10940
rect 11500 10856 11540 10900
rect 11203 10816 11212 10856
rect 11252 10816 11540 10856
rect 11596 10856 11636 10900
rect 11596 10816 12076 10856
rect 12116 10816 12125 10856
rect 12556 10688 12596 10900
rect 2659 10648 2668 10688
rect 2708 10648 5492 10688
rect 6883 10648 6892 10688
rect 6932 10648 11156 10688
rect 11299 10648 11308 10688
rect 11348 10648 12596 10688
rect 1795 10564 1804 10604
rect 1844 10564 4820 10604
rect 4919 10564 4928 10604
rect 4968 10564 5010 10604
rect 5050 10564 5092 10604
rect 5132 10564 5174 10604
rect 5214 10564 5256 10604
rect 5296 10564 5305 10604
rect 0 10520 90 10540
rect 0 10480 652 10520
rect 692 10480 701 10520
rect 0 10460 90 10480
rect 259 10396 268 10436
rect 308 10396 1180 10436
rect 1220 10396 1229 10436
rect 1507 10396 1516 10436
rect 1556 10396 2236 10436
rect 2276 10396 2285 10436
rect 2947 10396 2956 10436
rect 2996 10396 3005 10436
rect 4457 10396 4588 10436
rect 4628 10396 4637 10436
rect 2956 10310 2996 10396
rect 4780 10352 4820 10564
rect 5452 10436 5492 10648
rect 12652 10604 12692 10984
rect 13612 10940 13652 10984
rect 14284 10940 14324 11236
rect 14921 11152 14956 11192
rect 14996 11152 15052 11192
rect 15092 11152 15101 11192
rect 19241 11152 19372 11192
rect 19412 11152 19421 11192
rect 19555 11152 19564 11192
rect 19604 11152 19708 11192
rect 19748 11152 19757 11192
rect 19939 11152 19948 11192
rect 19988 11152 20092 11192
rect 20132 11152 20141 11192
rect 14371 11068 14380 11108
rect 14420 11068 16052 11108
rect 15907 10984 15916 11024
rect 15956 10984 15965 11024
rect 14860 10940 14900 10949
rect 8995 10564 9004 10604
rect 9044 10564 12692 10604
rect 12940 10900 13044 10940
rect 13084 10900 13093 10940
rect 13603 10900 13612 10940
rect 13652 10900 14324 10940
rect 14467 10900 14476 10940
rect 14516 10900 14860 10940
rect 15418 10900 15427 10940
rect 15467 10900 15476 10940
rect 15523 10900 15532 10940
rect 15572 10900 15860 10940
rect 12940 10520 12980 10900
rect 14860 10891 14900 10900
rect 13219 10732 13228 10772
rect 13268 10732 14380 10772
rect 14420 10732 14429 10772
rect 15436 10604 15476 10900
rect 15820 10604 15860 10900
rect 15916 10688 15956 10984
rect 16012 10940 16052 11068
rect 21510 11024 21600 11044
rect 17194 10984 17203 11024
rect 17243 10984 17548 11024
rect 17588 10984 17597 11024
rect 19747 10984 19756 11024
rect 19796 10984 19948 11024
rect 19988 10984 19997 11024
rect 20323 10984 20332 11024
rect 20372 10984 21196 11024
rect 21236 10984 21245 11024
rect 21379 10984 21388 11024
rect 21428 10984 21600 11024
rect 21510 10964 21600 10984
rect 16492 10940 16532 10949
rect 19180 10940 19220 10949
rect 16003 10900 16012 10940
rect 16052 10900 16061 10940
rect 16361 10900 16492 10940
rect 16532 10900 16541 10940
rect 16867 10900 16876 10940
rect 16916 10900 16980 10940
rect 17020 10900 17047 10940
rect 17731 10900 17740 10940
rect 17780 10900 17932 10940
rect 17972 10900 17981 10940
rect 18691 10900 18700 10940
rect 18740 10900 19180 10940
rect 16492 10891 16532 10900
rect 19180 10891 19220 10900
rect 16387 10732 16396 10772
rect 16436 10732 17308 10772
rect 17348 10732 17357 10772
rect 15916 10648 17260 10688
rect 17300 10648 17309 10688
rect 15436 10564 15668 10604
rect 15820 10564 18028 10604
rect 18068 10564 18077 10604
rect 20039 10564 20048 10604
rect 20088 10564 20130 10604
rect 20170 10564 20212 10604
rect 20252 10564 20294 10604
rect 20334 10564 20376 10604
rect 20416 10564 20425 10604
rect 12172 10480 12980 10520
rect 12172 10436 12212 10480
rect 15628 10436 15668 10564
rect 21510 10520 21600 10540
rect 19555 10480 19564 10520
rect 19604 10480 21600 10520
rect 21510 10460 21600 10480
rect 5452 10396 7220 10436
rect 7939 10396 7948 10436
rect 7988 10396 8044 10436
rect 8084 10396 8119 10436
rect 12163 10396 12172 10436
rect 12212 10396 12221 10436
rect 12451 10396 12460 10436
rect 12500 10396 12844 10436
rect 12884 10396 13076 10436
rect 13699 10396 13708 10436
rect 13748 10396 14188 10436
rect 14228 10396 14237 10436
rect 15628 10396 15820 10436
rect 15860 10396 15869 10436
rect 17635 10396 17644 10436
rect 17684 10396 17836 10436
rect 17876 10396 17885 10436
rect 18019 10396 18028 10436
rect 18068 10396 18604 10436
rect 18644 10396 19604 10436
rect 20083 10396 20092 10436
rect 20132 10396 20524 10436
rect 20564 10396 20573 10436
rect 3235 10312 3244 10352
rect 3284 10312 3860 10352
rect 2946 10301 2996 10310
rect 2699 10228 2764 10268
rect 2804 10228 2830 10268
rect 2870 10228 2879 10268
rect 2946 10261 2947 10301
rect 2987 10261 2996 10301
rect 3820 10268 3860 10312
rect 4780 10312 7084 10352
rect 7124 10312 7133 10352
rect 4780 10268 4820 10312
rect 2946 10252 2996 10261
rect 3331 10228 3340 10268
rect 3380 10228 3628 10268
rect 3668 10228 3677 10268
rect 3820 10259 3956 10268
rect 3820 10228 3916 10259
rect 4195 10228 4204 10268
rect 4244 10259 4436 10268
rect 4244 10228 4396 10259
rect 3916 10210 3956 10219
rect 4771 10228 4780 10268
rect 4820 10228 4829 10268
rect 6028 10259 6068 10268
rect 4396 10210 4436 10219
rect 6377 10228 6508 10268
rect 6548 10228 6557 10268
rect 0 10184 90 10204
rect 6028 10184 6068 10219
rect 0 10144 172 10184
rect 212 10144 221 10184
rect 1411 10144 1420 10184
rect 1460 10144 1469 10184
rect 1699 10144 1708 10184
rect 1748 10144 1900 10184
rect 1940 10144 1949 10184
rect 2131 10144 2140 10184
rect 2180 10144 2284 10184
rect 2324 10144 2333 10184
rect 2467 10144 2476 10184
rect 2516 10144 2860 10184
rect 2900 10144 2909 10184
rect 3305 10144 3436 10184
rect 3476 10144 3485 10184
rect 6028 10144 6316 10184
rect 6356 10144 6365 10184
rect 0 10124 90 10144
rect 1420 10016 1460 10144
rect 7180 10100 7220 10396
rect 10828 10312 11116 10352
rect 11156 10312 11165 10352
rect 12163 10312 12172 10352
rect 12212 10312 12364 10352
rect 12404 10312 12596 10352
rect 7555 10228 7564 10268
rect 7604 10259 7796 10268
rect 7604 10228 7756 10259
rect 10601 10228 10732 10268
rect 10772 10228 10781 10268
rect 7756 10210 7796 10219
rect 7843 10144 7852 10184
rect 7892 10144 8332 10184
rect 8372 10144 8381 10184
rect 9283 10144 9292 10184
rect 9332 10144 10060 10184
rect 10100 10144 10109 10184
rect 10828 10100 10868 10312
rect 12556 10268 12596 10312
rect 7180 10060 8092 10100
rect 8132 10060 8141 10100
rect 10723 10060 10732 10100
rect 10772 10060 10868 10100
rect 10924 10228 11404 10268
rect 11444 10228 11453 10268
rect 11779 10228 11788 10268
rect 11828 10259 12020 10268
rect 11828 10228 11980 10259
rect 10924 10016 10964 10228
rect 12067 10228 12076 10268
rect 12116 10228 12451 10268
rect 12491 10228 12500 10268
rect 12547 10228 12556 10268
rect 12596 10228 12605 10268
rect 12931 10228 12940 10268
rect 12980 10228 12989 10268
rect 11980 10184 12020 10219
rect 11933 10144 11980 10184
rect 12020 10144 12029 10184
rect 12940 10100 12980 10228
rect 13036 10184 13076 10396
rect 13516 10312 13804 10352
rect 13844 10312 13853 10352
rect 14380 10312 16300 10352
rect 16340 10312 16349 10352
rect 17635 10312 17644 10352
rect 17684 10312 17923 10352
rect 17963 10312 17972 10352
rect 18403 10312 18412 10352
rect 18452 10312 19220 10352
rect 13516 10259 13556 10312
rect 14380 10268 14420 10312
rect 13865 10228 13996 10268
rect 14036 10228 14045 10268
rect 14371 10228 14380 10268
rect 14420 10228 14429 10268
rect 15497 10228 15628 10268
rect 15668 10228 15677 10268
rect 16195 10228 16204 10268
rect 16244 10228 16253 10268
rect 17321 10228 17452 10268
rect 17492 10228 17501 10268
rect 18106 10228 18115 10268
rect 18155 10228 18508 10268
rect 18548 10228 18557 10268
rect 18604 10259 18644 10268
rect 13516 10210 13556 10219
rect 13996 10210 14036 10219
rect 15628 10184 15668 10219
rect 13027 10144 13036 10184
rect 13076 10144 13085 10184
rect 14467 10144 14476 10184
rect 14516 10144 15668 10184
rect 16204 10100 16244 10228
rect 17452 10210 17492 10219
rect 18604 10184 18644 10219
rect 18892 10228 19084 10268
rect 19124 10228 19133 10268
rect 12739 10060 12748 10100
rect 12788 10060 13516 10100
rect 13556 10060 13565 10100
rect 15331 10060 15340 10100
rect 15380 10060 16244 10100
rect 17068 10144 17396 10184
rect 17068 10016 17108 10144
rect 17356 10100 17396 10144
rect 17548 10144 18700 10184
rect 18740 10144 18804 10184
rect 17548 10100 17588 10144
rect 17356 10060 17588 10100
rect 18892 10016 18932 10228
rect 19180 10184 19220 10312
rect 19564 10268 19604 10396
rect 19555 10228 19564 10268
rect 19604 10228 19613 10268
rect 19660 10209 19677 10249
rect 19717 10209 19726 10249
rect 19171 10144 19180 10184
rect 19220 10144 19229 10184
rect 19660 10100 19700 10209
rect 20323 10144 20332 10184
rect 20372 10144 20812 10184
rect 20852 10144 20861 10184
rect 19267 10060 19276 10100
rect 19316 10060 19700 10100
rect 21510 10016 21600 10036
rect 1420 9976 1708 10016
rect 1748 9976 1757 10016
rect 6089 9976 6220 10016
rect 6260 9976 6269 10016
rect 6316 9976 10964 10016
rect 11107 9976 11116 10016
rect 11156 9976 13900 10016
rect 13940 9976 13949 10016
rect 15907 9976 15916 10016
rect 15956 9976 17108 10016
rect 18508 9976 18932 10016
rect 21091 9976 21100 10016
rect 21140 9976 21600 10016
rect 6316 9932 6356 9976
rect 2860 9892 6356 9932
rect 0 9848 90 9868
rect 0 9808 1228 9848
rect 1268 9808 1277 9848
rect 0 9788 90 9808
rect 355 9640 364 9680
rect 404 9640 1180 9680
rect 1220 9640 1229 9680
rect 2275 9556 2284 9596
rect 2324 9556 2476 9596
rect 2516 9556 2525 9596
rect 0 9512 90 9532
rect 2860 9512 2900 9892
rect 3679 9808 3688 9848
rect 3728 9808 3770 9848
rect 3810 9808 3852 9848
rect 3892 9808 3934 9848
rect 3974 9808 4016 9848
rect 4056 9808 4065 9848
rect 8899 9808 8908 9848
rect 8948 9808 18124 9848
rect 18164 9808 18173 9848
rect 18508 9764 18548 9976
rect 21510 9956 21600 9976
rect 18799 9808 18808 9848
rect 18848 9808 18890 9848
rect 18930 9808 18972 9848
rect 19012 9808 19054 9848
rect 19094 9808 19136 9848
rect 19176 9808 19185 9848
rect 3427 9724 3436 9764
rect 3476 9724 9004 9764
rect 9044 9724 9053 9764
rect 10243 9724 10252 9764
rect 10292 9724 10732 9764
rect 10772 9724 11444 9764
rect 11491 9724 11500 9764
rect 11540 9724 15820 9764
rect 15860 9724 15869 9764
rect 16483 9724 16492 9764
rect 16532 9724 18548 9764
rect 11404 9680 11444 9724
rect 3139 9640 3148 9680
rect 3188 9640 3484 9680
rect 3524 9640 3533 9680
rect 3628 9640 5548 9680
rect 5588 9640 5597 9680
rect 5827 9640 5836 9680
rect 5876 9640 6076 9680
rect 6116 9640 6125 9680
rect 9859 9640 9868 9680
rect 9908 9640 11348 9680
rect 11404 9640 14227 9680
rect 14267 9640 14276 9680
rect 15209 9640 15292 9680
rect 15332 9640 15340 9680
rect 15380 9640 15389 9680
rect 16745 9640 16876 9680
rect 16916 9640 16925 9680
rect 16972 9640 18220 9680
rect 18260 9640 18269 9680
rect 3331 9556 3340 9596
rect 3380 9556 3532 9596
rect 3572 9556 3581 9596
rect 0 9472 1076 9512
rect 1411 9472 1420 9512
rect 1460 9472 2900 9512
rect 0 9452 90 9472
rect 1036 9428 1076 9472
rect 3148 9428 3188 9437
rect 3628 9428 3668 9640
rect 11308 9596 11348 9640
rect 16972 9596 17012 9640
rect 3724 9556 11164 9596
rect 11204 9556 11213 9596
rect 11308 9556 16300 9596
rect 16340 9556 16349 9596
rect 16588 9556 17012 9596
rect 17635 9556 17644 9596
rect 17684 9556 17693 9596
rect 3724 9512 3764 9556
rect 3715 9472 3724 9512
rect 3764 9472 3773 9512
rect 4003 9472 4012 9512
rect 4052 9472 4340 9512
rect 4553 9472 4684 9512
rect 4724 9472 4733 9512
rect 5962 9472 5971 9512
rect 6011 9472 6316 9512
rect 6356 9472 6365 9512
rect 6883 9472 6892 9512
rect 6932 9472 6941 9512
rect 9187 9472 9196 9512
rect 9236 9472 9772 9512
rect 9812 9472 9868 9512
rect 9908 9472 9917 9512
rect 9964 9472 10252 9512
rect 10292 9472 10301 9512
rect 11050 9472 11059 9512
rect 11099 9472 11404 9512
rect 11444 9472 11453 9512
rect 12739 9472 12748 9512
rect 12788 9472 12940 9512
rect 12980 9472 12989 9512
rect 14371 9472 14380 9512
rect 14420 9472 14572 9512
rect 14612 9472 14621 9512
rect 14755 9472 14764 9512
rect 14804 9472 15052 9512
rect 15092 9472 15101 9512
rect 4300 9428 4340 9472
rect 5260 9428 5300 9437
rect 1036 9388 1708 9428
rect 1748 9388 1757 9428
rect 1891 9388 1900 9428
rect 1940 9388 2284 9428
rect 2324 9388 2333 9428
rect 2467 9388 2476 9428
rect 2516 9388 3148 9428
rect 3188 9388 3668 9428
rect 4186 9388 4195 9428
rect 4235 9388 4244 9428
rect 4291 9388 4300 9428
rect 4340 9388 4349 9428
rect 4771 9388 4780 9428
rect 4820 9388 5164 9428
rect 5204 9388 5213 9428
rect 5770 9388 5779 9428
rect 5819 9388 6220 9428
rect 6260 9388 6269 9428
rect 3148 9379 3188 9388
rect 4204 9344 4244 9388
rect 4780 9344 4820 9388
rect 4204 9304 4492 9344
rect 4532 9304 4541 9344
rect 4675 9304 4684 9344
rect 4724 9304 4820 9344
rect 5260 9344 5300 9388
rect 5260 9304 6796 9344
rect 6836 9304 6845 9344
rect 4099 9220 4108 9260
rect 4148 9220 6164 9260
rect 6595 9220 6604 9260
rect 6644 9220 6652 9260
rect 6692 9220 6775 9260
rect 0 9176 90 9196
rect 0 9136 3532 9176
rect 3572 9136 3581 9176
rect 0 9116 90 9136
rect 6124 9092 6164 9220
rect 6892 9176 6932 9472
rect 8812 9428 8852 9437
rect 9964 9428 10004 9472
rect 10348 9428 10388 9437
rect 13516 9428 13556 9437
rect 16588 9428 16628 9556
rect 17644 9512 17684 9556
rect 17251 9472 17260 9512
rect 17300 9472 17309 9512
rect 17635 9472 17644 9512
rect 17684 9472 17731 9512
rect 18281 9472 18412 9512
rect 18452 9472 18461 9512
rect 7433 9388 7564 9428
rect 7604 9388 7613 9428
rect 8777 9388 8812 9428
rect 8852 9388 8908 9428
rect 8948 9388 8957 9428
rect 9004 9388 9283 9428
rect 9323 9388 9332 9428
rect 9379 9388 9388 9428
rect 9428 9388 9437 9428
rect 9859 9388 9868 9428
rect 9908 9388 10004 9428
rect 10051 9388 10060 9428
rect 10100 9388 10348 9428
rect 8812 9379 8852 9388
rect 9004 9344 9044 9388
rect 9388 9344 9428 9388
rect 10348 9379 10388 9388
rect 10444 9388 10836 9428
rect 10876 9388 10885 9428
rect 11875 9388 11884 9428
rect 11924 9388 12451 9428
rect 12491 9388 12500 9428
rect 12547 9388 12556 9428
rect 12596 9388 12605 9428
rect 12835 9388 12844 9428
rect 12884 9388 13036 9428
rect 13076 9388 13085 9428
rect 13315 9388 13324 9428
rect 13364 9388 13516 9428
rect 13556 9388 13804 9428
rect 13844 9388 13853 9428
rect 14026 9388 14035 9428
rect 14075 9388 14284 9428
rect 14324 9388 14333 9428
rect 15427 9388 15436 9428
rect 15476 9388 16628 9428
rect 16684 9428 16724 9437
rect 8995 9304 9004 9344
rect 9044 9304 9053 9344
rect 9388 9304 10156 9344
rect 10196 9304 10205 9344
rect 10444 9260 10484 9388
rect 12556 9344 12596 9388
rect 13516 9379 13556 9388
rect 16684 9344 16724 9388
rect 12355 9304 12364 9344
rect 12404 9304 12596 9344
rect 14467 9304 14476 9344
rect 14516 9304 16724 9344
rect 10243 9220 10252 9260
rect 10292 9220 10484 9260
rect 13603 9220 13612 9260
rect 13652 9220 14332 9260
rect 14372 9220 14381 9260
rect 16579 9220 16588 9260
rect 16628 9220 17020 9260
rect 17060 9220 17069 9260
rect 17260 9176 17300 9472
rect 18508 9428 18548 9724
rect 20035 9640 20044 9680
rect 20084 9640 20092 9680
rect 20132 9640 20215 9680
rect 21510 9512 21600 9532
rect 20323 9472 20332 9512
rect 20372 9472 20908 9512
rect 20948 9472 20957 9512
rect 21187 9472 21196 9512
rect 21236 9472 21600 9512
rect 21510 9452 21600 9472
rect 18988 9428 19028 9437
rect 17731 9388 17740 9428
rect 17780 9388 17923 9428
rect 17963 9388 17972 9428
rect 18019 9388 18028 9428
rect 18068 9388 18077 9428
rect 18499 9388 18508 9428
rect 18548 9388 18557 9428
rect 18691 9388 18700 9428
rect 18740 9388 18988 9428
rect 19498 9388 19507 9428
rect 19547 9388 19756 9428
rect 19796 9388 19805 9428
rect 18028 9344 18068 9388
rect 18988 9379 19028 9388
rect 18028 9304 18604 9344
rect 18644 9304 18653 9344
rect 17395 9220 17404 9260
rect 17444 9220 17548 9260
rect 17588 9220 17597 9260
rect 18115 9220 18124 9260
rect 18164 9220 19180 9260
rect 19220 9220 19229 9260
rect 19529 9220 19660 9260
rect 19700 9220 19709 9260
rect 6211 9136 6220 9176
rect 6260 9136 6932 9176
rect 7171 9136 7180 9176
rect 7220 9136 13132 9176
rect 13172 9136 14188 9176
rect 14228 9136 14237 9176
rect 17260 9136 19508 9176
rect 4919 9052 4928 9092
rect 4968 9052 5010 9092
rect 5050 9052 5092 9092
rect 5132 9052 5174 9092
rect 5214 9052 5256 9092
rect 5296 9052 5305 9092
rect 6124 9052 7796 9092
rect 16291 9052 16300 9092
rect 16340 9052 18700 9092
rect 18740 9052 18749 9092
rect 7756 9008 7796 9052
rect 19468 9008 19508 9136
rect 20039 9052 20048 9092
rect 20088 9052 20130 9092
rect 20170 9052 20212 9092
rect 20252 9052 20294 9092
rect 20334 9052 20376 9092
rect 20416 9052 20425 9092
rect 21510 9008 21600 9028
rect 3052 8968 7660 9008
rect 7700 8968 7709 9008
rect 7756 8968 19412 9008
rect 19468 8968 21600 9008
rect 2563 8884 2572 8924
rect 2612 8884 2668 8924
rect 2708 8884 2743 8924
rect 0 8840 90 8860
rect 0 8800 1132 8840
rect 1172 8800 1181 8840
rect 1891 8800 1900 8840
rect 1940 8800 2812 8840
rect 2852 8800 2861 8840
rect 0 8780 90 8800
rect 1219 8716 1228 8756
rect 1268 8716 1420 8756
rect 1460 8716 1804 8756
rect 1844 8716 1853 8756
rect 2345 8716 2476 8756
rect 2516 8716 2525 8756
rect 2476 8698 2516 8707
rect 3052 8672 3092 8968
rect 19372 8924 19412 8968
rect 21510 8948 21600 8968
rect 4003 8884 4012 8924
rect 4052 8884 5068 8924
rect 5108 8884 5117 8924
rect 5260 8884 7372 8924
rect 7412 8884 7421 8924
rect 10051 8884 10060 8924
rect 10100 8884 11404 8924
rect 11444 8884 11453 8924
rect 11753 8884 11884 8924
rect 11924 8884 11933 8924
rect 13123 8884 13132 8924
rect 13172 8884 13996 8924
rect 14036 8884 14860 8924
rect 14900 8884 14909 8924
rect 15139 8884 15148 8924
rect 15188 8884 15292 8924
rect 15332 8884 15341 8924
rect 15907 8884 15916 8924
rect 15956 8884 16684 8924
rect 16724 8884 16916 8924
rect 16963 8884 16972 8924
rect 17012 8884 17492 8924
rect 17539 8884 17548 8924
rect 17588 8884 18124 8924
rect 18164 8884 18173 8924
rect 19145 8884 19180 8924
rect 19220 8884 19276 8924
rect 19316 8884 19325 8924
rect 19372 8884 20092 8924
rect 20132 8884 20141 8924
rect 3331 8800 3340 8840
rect 3380 8800 3772 8840
rect 3812 8800 3821 8840
rect 4396 8756 4436 8884
rect 4675 8800 4684 8840
rect 4724 8800 4916 8840
rect 3244 8716 3436 8756
rect 3476 8716 3485 8756
rect 4099 8716 4108 8756
rect 4148 8716 4291 8756
rect 4331 8716 4340 8756
rect 4387 8716 4396 8756
rect 4436 8716 4445 8756
rect 4771 8716 4780 8756
rect 4820 8716 4829 8756
rect 3244 8672 3284 8716
rect 3043 8632 3052 8672
rect 3092 8632 3101 8672
rect 3235 8632 3244 8672
rect 3284 8632 3293 8672
rect 3475 8632 3484 8672
rect 3524 8632 3820 8672
rect 3860 8632 3869 8672
rect 4003 8632 4012 8672
rect 4052 8632 4588 8672
rect 4628 8632 4637 8672
rect 4780 8588 4820 8716
rect 4876 8672 4916 8800
rect 5260 8756 5300 8884
rect 6115 8800 6124 8840
rect 6164 8800 6452 8840
rect 6691 8800 6700 8840
rect 6740 8800 8188 8840
rect 8228 8800 8237 8840
rect 8620 8800 10924 8840
rect 10964 8800 10973 8840
rect 11971 8800 11980 8840
rect 12020 8800 14668 8840
rect 14708 8800 15100 8840
rect 15140 8800 15149 8840
rect 15619 8800 15628 8840
rect 15668 8800 15956 8840
rect 16099 8800 16108 8840
rect 16148 8800 16436 8840
rect 6412 8756 6452 8800
rect 8620 8756 8660 8800
rect 15916 8756 15956 8800
rect 5260 8747 5396 8756
rect 5260 8716 5356 8747
rect 5705 8716 5836 8756
rect 5876 8716 5885 8756
rect 6298 8716 6307 8756
rect 6347 8716 6356 8756
rect 6403 8716 6412 8756
rect 6452 8716 6461 8756
rect 6787 8716 6796 8756
rect 6836 8716 7084 8756
rect 7124 8716 7133 8756
rect 7241 8716 7372 8756
rect 7412 8716 7421 8756
rect 7721 8716 7852 8756
rect 7892 8716 7901 8756
rect 8489 8716 8620 8756
rect 8660 8716 8669 8756
rect 8899 8716 8908 8756
rect 8948 8747 9908 8756
rect 8948 8716 9868 8747
rect 5356 8698 5396 8707
rect 5836 8698 5876 8707
rect 6312 8672 6352 8716
rect 4867 8632 4876 8672
rect 4916 8632 4925 8672
rect 6058 8632 6067 8672
rect 6107 8632 6220 8672
rect 6260 8632 6269 8672
rect 6312 8632 6700 8672
rect 6740 8632 6749 8672
rect 6796 8588 6836 8716
rect 7372 8698 7412 8707
rect 7852 8698 7892 8707
rect 10409 8716 10444 8756
rect 10484 8716 10540 8756
rect 10580 8716 10589 8756
rect 11561 8716 11596 8756
rect 11636 8747 11732 8756
rect 11636 8716 11692 8747
rect 9868 8698 9908 8707
rect 11779 8716 11788 8756
rect 11828 8716 12259 8756
rect 12299 8716 12308 8756
rect 12355 8716 12364 8756
rect 12404 8716 12535 8756
rect 12617 8716 12748 8756
rect 12788 8716 12797 8756
rect 13193 8716 13324 8756
rect 13364 8716 13373 8756
rect 13673 8716 13804 8756
rect 13844 8716 13853 8756
rect 14179 8716 14188 8756
rect 14228 8716 15572 8756
rect 15802 8716 15811 8756
rect 15851 8716 15860 8756
rect 15907 8716 15916 8756
rect 15956 8716 15965 8756
rect 16169 8716 16300 8756
rect 16340 8716 16349 8756
rect 11692 8698 11732 8707
rect 12364 8672 12404 8716
rect 13324 8698 13364 8707
rect 13804 8698 13844 8707
rect 15532 8672 15572 8716
rect 15820 8672 15860 8716
rect 16396 8672 16436 8800
rect 16876 8747 16916 8884
rect 17452 8756 17492 8884
rect 18403 8800 18412 8840
rect 18452 8800 19708 8840
rect 19748 8800 19757 8840
rect 17225 8716 17356 8756
rect 17396 8716 17405 8756
rect 17452 8716 17740 8756
rect 17780 8716 17789 8756
rect 18988 8747 19372 8756
rect 16876 8698 16916 8707
rect 17356 8698 17396 8707
rect 19028 8716 19372 8747
rect 19412 8716 19421 8756
rect 18988 8672 19028 8707
rect 6883 8632 6892 8672
rect 6932 8632 7063 8672
rect 8074 8632 8083 8672
rect 8123 8632 8428 8672
rect 8468 8632 8477 8672
rect 11971 8632 11980 8672
rect 12020 8632 12404 8672
rect 12713 8632 12844 8672
rect 12884 8632 12893 8672
rect 14851 8632 14860 8672
rect 14900 8632 15476 8672
rect 15523 8632 15532 8672
rect 15572 8632 15581 8672
rect 15820 8632 16108 8672
rect 16148 8632 16157 8672
rect 16387 8632 16396 8672
rect 16436 8632 16445 8672
rect 17443 8632 17452 8672
rect 17492 8632 19028 8672
rect 19171 8632 19180 8672
rect 19220 8632 19324 8672
rect 19364 8632 19373 8672
rect 19433 8632 19564 8672
rect 19604 8632 19613 8672
rect 19817 8632 19948 8672
rect 19988 8632 19997 8672
rect 20323 8632 20332 8672
rect 20372 8632 21004 8672
rect 21044 8632 21053 8672
rect 15436 8588 15476 8632
rect 4780 8548 6412 8588
rect 6452 8548 6836 8588
rect 7555 8548 7564 8588
rect 7604 8548 12556 8588
rect 12596 8548 12605 8588
rect 15436 8548 15820 8588
rect 15860 8548 16492 8588
rect 16532 8548 16541 8588
rect 0 8504 90 8524
rect 21510 8504 21600 8524
rect 0 8464 844 8504
rect 884 8464 893 8504
rect 10051 8464 10060 8504
rect 10100 8464 10252 8504
rect 10292 8464 10301 8504
rect 20899 8464 20908 8504
rect 20948 8464 21600 8504
rect 0 8444 90 8464
rect 21510 8444 21600 8464
rect 11011 8380 11020 8420
rect 11060 8380 13324 8420
rect 13364 8380 13373 8420
rect 3679 8296 3688 8336
rect 3728 8296 3770 8336
rect 3810 8296 3852 8336
rect 3892 8296 3934 8336
rect 3974 8296 4016 8336
rect 4056 8296 4065 8336
rect 10348 8296 15052 8336
rect 15092 8296 15101 8336
rect 18799 8296 18808 8336
rect 18848 8296 18890 8336
rect 18930 8296 18972 8336
rect 19012 8296 19054 8336
rect 19094 8296 19136 8336
rect 19176 8296 19185 8336
rect 6403 8212 6412 8252
rect 6452 8212 9676 8252
rect 9716 8212 9725 8252
rect 0 8168 90 8188
rect 0 8128 364 8168
rect 404 8128 413 8168
rect 2851 8128 2860 8168
rect 2900 8128 3031 8168
rect 4361 8128 4492 8168
rect 4532 8128 4541 8168
rect 5827 8128 5836 8168
rect 5876 8128 6220 8168
rect 6260 8128 6269 8168
rect 7817 8128 7852 8168
rect 7892 8128 7948 8168
rect 7988 8128 7997 8168
rect 0 8108 90 8128
rect 2275 8044 2284 8084
rect 2324 8044 3092 8084
rect 1507 7960 1516 8000
rect 1556 7960 2708 8000
rect 2668 7916 2708 7960
rect 3052 7916 3092 8044
rect 4300 8044 6316 8084
rect 6356 8044 6365 8084
rect 4300 7916 4340 8044
rect 8140 7960 9908 8000
rect 6028 7916 6068 7925
rect 7756 7916 7796 7925
rect 8140 7916 8180 7960
rect 9868 7916 9908 7960
rect 10348 7916 10388 8296
rect 10915 8212 10924 8252
rect 10964 8212 15476 8252
rect 11657 8128 11788 8168
rect 11828 8128 11837 8168
rect 13673 8128 13804 8168
rect 13844 8128 13853 8168
rect 13987 8128 13996 8168
rect 14036 8128 14167 8168
rect 12364 8044 15340 8084
rect 15380 8044 15389 8084
rect 11596 7916 11636 7925
rect 12364 7916 12404 8044
rect 12940 7960 13652 8000
rect 1289 7876 1420 7916
rect 1460 7876 1469 7916
rect 2633 7876 2668 7916
rect 2708 7876 2764 7916
rect 2804 7876 2813 7916
rect 3043 7876 3052 7916
rect 3092 7876 3101 7916
rect 4771 7876 4780 7916
rect 4820 7876 4829 7916
rect 6068 7876 6220 7916
rect 6260 7876 6269 7916
rect 6412 7876 6508 7916
rect 6548 7876 7180 7916
rect 7220 7876 7229 7916
rect 7796 7876 8140 7916
rect 8180 7876 8189 7916
rect 8489 7876 8620 7916
rect 8660 7876 8669 7916
rect 10339 7876 10348 7916
rect 10388 7876 10397 7916
rect 11465 7876 11596 7916
rect 11636 7876 11645 7916
rect 12355 7876 12364 7916
rect 12404 7876 12413 7916
rect 2668 7867 2708 7876
rect 4300 7867 4340 7876
rect 0 7832 90 7852
rect 0 7792 1652 7832
rect 0 7772 90 7792
rect 1612 7748 1652 7792
rect 4780 7748 4820 7876
rect 6028 7867 6068 7876
rect 6412 7748 6452 7876
rect 7756 7867 7796 7876
rect 9868 7867 9908 7876
rect 11596 7832 11636 7876
rect 12940 7832 12980 7960
rect 13612 7916 13652 7960
rect 14188 7916 14228 7925
rect 15436 7916 15476 8212
rect 16147 8128 16156 8168
rect 16196 8128 16300 8168
rect 16340 8128 16349 8168
rect 17609 8128 17740 8168
rect 17780 8128 17789 8168
rect 18499 8128 18508 8168
rect 18548 8128 19948 8168
rect 19988 8128 19997 8168
rect 18691 8044 18700 8084
rect 18740 8044 20092 8084
rect 20132 8044 20141 8084
rect 21510 8000 21600 8020
rect 15907 7960 15916 8000
rect 15956 7960 16012 8000
rect 16052 7960 16087 8000
rect 17993 7960 18124 8000
rect 18164 7960 18173 8000
rect 20323 7960 20332 8000
rect 20372 7960 21388 8000
rect 21428 7960 21437 8000
rect 21484 7940 21600 8000
rect 17548 7916 17588 7925
rect 19756 7916 19796 7925
rect 21484 7916 21524 7940
rect 13652 7876 14188 7916
rect 15427 7876 15436 7916
rect 15476 7876 15485 7916
rect 16195 7876 16204 7916
rect 16244 7876 16300 7916
rect 16340 7876 16375 7916
rect 17443 7876 17452 7916
rect 17492 7876 17548 7916
rect 17588 7876 17623 7916
rect 18019 7876 18028 7916
rect 18068 7876 18508 7916
rect 18548 7876 18557 7916
rect 19363 7876 19372 7916
rect 19412 7876 19756 7916
rect 20707 7876 20716 7916
rect 20756 7876 21524 7916
rect 13612 7867 13652 7876
rect 11596 7792 12980 7832
rect 1612 7708 3148 7748
rect 3188 7708 3197 7748
rect 4780 7708 6452 7748
rect 10051 7708 10060 7748
rect 10100 7708 10109 7748
rect 4919 7540 4928 7580
rect 4968 7540 5010 7580
rect 5050 7540 5092 7580
rect 5132 7540 5174 7580
rect 5214 7540 5256 7580
rect 5296 7540 5305 7580
rect 0 7496 90 7516
rect 0 7456 1036 7496
rect 1076 7456 1085 7496
rect 0 7436 90 7456
rect 3811 7372 3820 7412
rect 3860 7372 4204 7412
rect 4244 7372 4253 7412
rect 6569 7372 6700 7412
rect 6740 7372 6749 7412
rect 3628 7288 6220 7328
rect 6260 7288 6269 7328
rect 6508 7288 8180 7328
rect 8652 7288 8716 7328
rect 8756 7288 9908 7328
rect 3628 7244 3668 7288
rect 4204 7244 4244 7288
rect 2275 7204 2284 7244
rect 2324 7204 2380 7244
rect 2420 7204 2455 7244
rect 2755 7204 2764 7244
rect 2804 7235 3668 7244
rect 2804 7204 3628 7235
rect 4195 7204 4204 7244
rect 4244 7204 4320 7244
rect 5251 7204 5260 7244
rect 5300 7204 5740 7244
rect 5780 7204 5789 7244
rect 6508 7235 6548 7288
rect 8140 7244 8180 7288
rect 8812 7244 8852 7288
rect 3628 7186 3668 7195
rect 6979 7204 6988 7244
rect 7028 7204 7564 7244
rect 7604 7204 7613 7244
rect 8131 7204 8140 7244
rect 8180 7235 8311 7244
rect 8180 7204 8236 7235
rect 6508 7186 6548 7195
rect 8276 7204 8311 7235
rect 8698 7204 8707 7244
rect 8747 7204 8756 7244
rect 8803 7204 8812 7244
rect 8852 7204 8861 7244
rect 9065 7204 9196 7244
rect 9236 7204 9245 7244
rect 9641 7204 9772 7244
rect 9812 7204 9821 7244
rect 8236 7186 8276 7195
rect 0 7160 90 7180
rect 0 7120 692 7160
rect 739 7120 748 7160
rect 788 7120 1180 7160
rect 1220 7120 1229 7160
rect 1411 7120 1420 7160
rect 1460 7120 1591 7160
rect 1673 7120 1804 7160
rect 1844 7120 1853 7160
rect 1939 7120 1948 7160
rect 1988 7120 1996 7160
rect 2036 7120 2119 7160
rect 2179 7120 2188 7160
rect 2228 7120 2860 7160
rect 2900 7120 2909 7160
rect 4195 7120 4204 7160
rect 4244 7120 4396 7160
rect 4436 7120 4445 7160
rect 4579 7120 4588 7160
rect 4628 7120 4759 7160
rect 4963 7120 4972 7160
rect 5012 7120 5356 7160
rect 5396 7120 5405 7160
rect 0 7100 90 7120
rect 652 7076 692 7120
rect 8716 7076 8756 7204
rect 9772 7186 9812 7195
rect 9868 7160 9908 7288
rect 10060 7244 10100 7708
rect 10636 7288 12556 7328
rect 12596 7288 12605 7328
rect 10636 7244 10676 7288
rect 10060 7235 10292 7244
rect 10060 7204 10252 7235
rect 10627 7204 10636 7244
rect 10676 7204 10685 7244
rect 11587 7204 11596 7244
rect 11636 7235 11924 7244
rect 11636 7204 11884 7235
rect 10252 7186 10292 7195
rect 12835 7204 12844 7244
rect 12884 7204 13324 7244
rect 13364 7204 13373 7244
rect 14092 7235 14132 7876
rect 14188 7867 14228 7876
rect 17548 7867 17588 7876
rect 19756 7867 19796 7876
rect 15811 7708 15820 7748
rect 15860 7708 17884 7748
rect 17924 7708 17933 7748
rect 15331 7624 15340 7664
rect 15380 7624 18700 7664
rect 18740 7624 18749 7664
rect 20039 7540 20048 7580
rect 20088 7540 20130 7580
rect 20170 7540 20212 7580
rect 20252 7540 20294 7580
rect 20334 7540 20376 7580
rect 20416 7540 20425 7580
rect 21510 7496 21600 7516
rect 17443 7456 17452 7496
rect 17492 7456 17972 7496
rect 20515 7456 20524 7496
rect 20564 7456 21600 7496
rect 15043 7372 15052 7412
rect 15092 7372 17588 7412
rect 15916 7244 15956 7372
rect 16300 7288 17452 7328
rect 17492 7288 17501 7328
rect 16300 7244 16340 7288
rect 17548 7244 17588 7372
rect 11884 7186 11924 7195
rect 14537 7204 14668 7244
rect 14708 7204 14717 7244
rect 15907 7204 15916 7244
rect 15956 7204 15965 7244
rect 16169 7204 16300 7244
rect 16340 7204 16349 7244
rect 17539 7204 17548 7244
rect 17588 7204 17597 7244
rect 17932 7235 17972 7456
rect 21510 7436 21600 7456
rect 14092 7186 14132 7195
rect 14668 7186 14708 7195
rect 16300 7186 16340 7195
rect 18691 7204 18700 7244
rect 18740 7204 19180 7244
rect 19220 7204 19229 7244
rect 17932 7186 17972 7195
rect 9283 7120 9292 7160
rect 9332 7120 9341 7160
rect 9868 7120 10196 7160
rect 652 7036 4348 7076
rect 4388 7036 4397 7076
rect 8419 7036 8428 7076
rect 8468 7036 8756 7076
rect 9292 7076 9332 7120
rect 10156 7076 10196 7120
rect 10348 7120 11308 7160
rect 11348 7120 11357 7160
rect 15977 7120 16099 7160
rect 16148 7120 16157 7160
rect 17347 7120 17356 7160
rect 17396 7120 17731 7160
rect 17771 7120 17780 7160
rect 19529 7120 19660 7160
rect 19700 7120 19709 7160
rect 20323 7120 20332 7160
rect 20372 7120 21100 7160
rect 21140 7120 21149 7160
rect 10348 7076 10388 7120
rect 9292 7036 9868 7076
rect 9908 7036 9917 7076
rect 10156 7036 10388 7076
rect 10483 7036 10492 7076
rect 10532 7036 10732 7076
rect 10772 7036 10781 7076
rect 11945 7036 12076 7076
rect 12116 7036 12125 7076
rect 14153 7036 14284 7076
rect 14324 7036 14333 7076
rect 14380 7036 20092 7076
rect 20132 7036 20141 7076
rect 14380 6992 14420 7036
rect 21510 6992 21600 7012
rect 931 6952 940 6992
rect 980 6952 1564 6992
rect 1604 6952 1613 6992
rect 3523 6952 3532 6992
rect 3572 6952 3964 6992
rect 4004 6952 4013 6992
rect 4108 6952 4732 6992
rect 4772 6952 4781 6992
rect 6211 6952 6220 6992
rect 6260 6952 12172 6992
rect 12212 6952 12221 6992
rect 12355 6952 12364 6992
rect 12404 6952 14420 6992
rect 14467 6952 14476 6992
rect 14516 6952 15340 6992
rect 15380 6952 15389 6992
rect 17347 6952 17356 6992
rect 17396 6952 19420 6992
rect 19460 6952 19469 6992
rect 19555 6952 19564 6992
rect 19604 6952 21600 6992
rect 4108 6908 4148 6952
rect 21510 6932 21600 6952
rect 2860 6868 4148 6908
rect 6115 6868 6124 6908
rect 6164 6868 12980 6908
rect 0 6824 90 6844
rect 2860 6824 2900 6868
rect 12940 6824 12980 6868
rect 0 6784 2900 6824
rect 3679 6784 3688 6824
rect 3728 6784 3770 6824
rect 3810 6784 3852 6824
rect 3892 6784 3934 6824
rect 3974 6784 4016 6824
rect 4056 6784 4065 6824
rect 4387 6784 4396 6824
rect 4436 6784 6028 6824
rect 6068 6784 6077 6824
rect 12940 6784 16396 6824
rect 16436 6784 16445 6824
rect 18799 6784 18808 6824
rect 18848 6784 18890 6824
rect 18930 6784 18972 6824
rect 19012 6784 19054 6824
rect 19094 6784 19136 6824
rect 19176 6784 19185 6824
rect 0 6764 90 6784
rect 2572 6700 12980 6740
rect 451 6616 460 6656
rect 500 6616 1180 6656
rect 1220 6616 1229 6656
rect 1555 6616 1564 6656
rect 1604 6616 1612 6656
rect 1652 6616 1735 6656
rect 1219 6532 1228 6572
rect 1268 6532 2332 6572
rect 2372 6532 2381 6572
rect 0 6488 90 6508
rect 2572 6488 2612 6700
rect 12940 6656 12980 6700
rect 2755 6616 2764 6656
rect 2804 6616 2812 6656
rect 2852 6616 2935 6656
rect 3065 6616 3148 6656
rect 3188 6616 3196 6656
rect 3236 6616 3245 6656
rect 3907 6616 3916 6656
rect 3956 6616 4108 6656
rect 4148 6616 4157 6656
rect 7939 6616 7948 6656
rect 7988 6616 12364 6656
rect 12404 6616 12413 6656
rect 12940 6616 15820 6656
rect 15860 6616 15869 6656
rect 19625 6616 19756 6656
rect 19796 6616 19805 6656
rect 2860 6532 3340 6572
rect 3380 6532 3389 6572
rect 3436 6532 6988 6572
rect 7028 6532 7037 6572
rect 8611 6532 8620 6572
rect 8660 6532 10300 6572
rect 10340 6532 10349 6572
rect 15916 6532 16588 6572
rect 16628 6532 16637 6572
rect 17251 6532 17260 6572
rect 17300 6532 20092 6572
rect 20132 6532 20141 6572
rect 20332 6532 21196 6572
rect 21236 6532 21245 6572
rect 0 6448 556 6488
rect 596 6448 605 6488
rect 1411 6448 1420 6488
rect 1460 6448 1612 6488
rect 1652 6448 1661 6488
rect 1795 6448 1804 6488
rect 1844 6448 1853 6488
rect 1987 6448 1996 6488
rect 2036 6448 2284 6488
rect 2324 6448 2333 6488
rect 2563 6448 2572 6488
rect 2612 6448 2621 6488
rect 0 6428 90 6448
rect 1804 6404 1844 6448
rect 2860 6404 2900 6532
rect 3436 6488 3476 6532
rect 15916 6488 15956 6532
rect 20332 6488 20372 6532
rect 21510 6488 21600 6508
rect 3043 6448 3052 6488
rect 3092 6448 3101 6488
rect 3427 6448 3436 6488
rect 3476 6448 3485 6488
rect 8899 6448 8908 6488
rect 8948 6448 9196 6488
rect 9236 6448 9245 6488
rect 9388 6448 9868 6488
rect 9908 6448 9917 6488
rect 10531 6448 10540 6488
rect 10580 6448 10732 6488
rect 10772 6448 10781 6488
rect 14921 6448 15052 6488
rect 15092 6448 15101 6488
rect 15785 6448 15916 6488
rect 15956 6448 15965 6488
rect 17194 6448 17203 6488
rect 17243 6448 17548 6488
rect 17588 6448 17597 6488
rect 20323 6448 20332 6488
rect 20372 6448 20381 6488
rect 20716 6448 21600 6488
rect 1804 6364 2900 6404
rect 3052 6320 3092 6448
rect 4108 6404 4148 6413
rect 7756 6404 7796 6413
rect 9388 6404 9428 6448
rect 4073 6364 4108 6404
rect 4148 6364 4204 6404
rect 4244 6364 4253 6404
rect 5347 6364 5356 6404
rect 5396 6364 5740 6404
rect 5780 6364 5789 6404
rect 6499 6364 6508 6404
rect 6548 6364 6892 6404
rect 6932 6364 6941 6404
rect 8035 6364 8044 6404
rect 8084 6364 8419 6404
rect 8459 6364 8468 6404
rect 8515 6364 8524 6404
rect 8564 6364 8716 6404
rect 8756 6364 8765 6404
rect 8995 6364 9004 6404
rect 9044 6364 9428 6404
rect 9478 6364 9487 6404
rect 9527 6364 9772 6404
rect 9812 6364 9821 6404
rect 4108 6355 4148 6364
rect 7756 6320 7796 6364
rect 9868 6320 9908 6448
rect 12364 6404 12404 6413
rect 14476 6404 14516 6413
rect 16492 6404 16532 6413
rect 19564 6404 19604 6413
rect 20716 6404 20756 6448
rect 21510 6428 21600 6448
rect 9955 6364 9964 6404
rect 10012 6364 10135 6404
rect 10531 6364 10540 6404
rect 10580 6364 11116 6404
rect 11156 6364 11165 6404
rect 12163 6364 12172 6404
rect 12212 6364 12364 6404
rect 13193 6364 13228 6404
rect 13268 6364 13324 6404
rect 13364 6364 13373 6404
rect 14345 6364 14476 6404
rect 14516 6364 14525 6404
rect 15275 6364 15340 6404
rect 15380 6364 15406 6404
rect 15446 6364 15455 6404
rect 15523 6364 15532 6404
rect 15572 6364 15581 6404
rect 15881 6364 16012 6404
rect 16052 6364 16061 6404
rect 16532 6364 16684 6404
rect 16724 6364 16733 6404
rect 16963 6364 16972 6404
rect 17020 6364 17143 6404
rect 18211 6364 18220 6404
rect 18260 6364 18316 6404
rect 18356 6364 18391 6404
rect 19363 6364 19372 6404
rect 19412 6364 19564 6404
rect 19939 6364 19948 6404
rect 19988 6364 20756 6404
rect 12364 6355 12404 6364
rect 14476 6355 14516 6364
rect 15532 6320 15572 6364
rect 16492 6355 16532 6364
rect 19564 6355 19604 6364
rect 2227 6280 2236 6320
rect 2276 6280 2860 6320
rect 2900 6280 2909 6320
rect 3052 6280 4052 6320
rect 6307 6280 6316 6320
rect 6356 6280 7796 6320
rect 7852 6280 8908 6320
rect 8948 6280 8957 6320
rect 9868 6280 11500 6320
rect 11540 6280 11549 6320
rect 15497 6280 15628 6320
rect 15668 6280 16396 6320
rect 16436 6280 16445 6320
rect 4012 6236 4052 6280
rect 7852 6236 7892 6280
rect 4012 6196 7892 6236
rect 7939 6196 7948 6236
rect 7988 6196 9868 6236
rect 9908 6196 9917 6236
rect 10025 6196 10156 6236
rect 10196 6196 10205 6236
rect 12547 6196 12556 6236
rect 12596 6196 13036 6236
rect 13076 6196 13085 6236
rect 14467 6196 14476 6236
rect 14516 6196 14668 6236
rect 14708 6196 14717 6236
rect 14764 6196 14812 6236
rect 14852 6196 14861 6236
rect 17177 6196 17260 6236
rect 17300 6196 17308 6236
rect 17348 6196 17357 6236
rect 0 6152 90 6172
rect 0 6112 1324 6152
rect 1364 6112 1373 6152
rect 10051 6112 10060 6152
rect 10100 6112 13132 6152
rect 13172 6112 13181 6152
rect 0 6092 90 6112
rect 14764 6068 14804 6196
rect 4919 6028 4928 6068
rect 4968 6028 5010 6068
rect 5050 6028 5092 6068
rect 5132 6028 5174 6068
rect 5214 6028 5256 6068
rect 5296 6028 5305 6068
rect 9379 6028 9388 6068
rect 9428 6028 9964 6068
rect 10004 6028 10013 6068
rect 10435 6028 10444 6068
rect 10484 6028 14804 6068
rect 20039 6028 20048 6068
rect 20088 6028 20130 6068
rect 20170 6028 20212 6068
rect 20252 6028 20294 6068
rect 20334 6028 20376 6068
rect 20416 6028 20425 6068
rect 21510 5984 21600 6004
rect 4492 5944 6604 5984
rect 6644 5944 6653 5984
rect 13315 5944 13324 5984
rect 13364 5944 14764 5984
rect 14804 5944 14813 5984
rect 19180 5944 21600 5984
rect 4492 5900 4532 5944
rect 1411 5860 1420 5900
rect 1460 5860 4532 5900
rect 4579 5860 4588 5900
rect 4628 5860 14612 5900
rect 14659 5860 14668 5900
rect 14708 5860 15052 5900
rect 15092 5860 15101 5900
rect 15619 5860 15628 5900
rect 15668 5860 16300 5900
rect 16340 5860 16349 5900
rect 16483 5860 16492 5900
rect 16532 5860 16972 5900
rect 17012 5860 17021 5900
rect 0 5816 90 5836
rect 14572 5816 14612 5860
rect 0 5776 268 5816
rect 308 5776 317 5816
rect 2092 5776 2332 5816
rect 2372 5776 2381 5816
rect 3244 5776 3340 5816
rect 3380 5776 3389 5816
rect 6220 5776 6508 5816
rect 6548 5776 6557 5816
rect 9676 5776 10540 5816
rect 10580 5776 10589 5816
rect 10860 5776 10924 5816
rect 10964 5776 11308 5816
rect 11348 5776 12596 5816
rect 0 5756 90 5776
rect 2092 5732 2132 5776
rect 3244 5732 3284 5776
rect 6220 5732 6260 5776
rect 9676 5732 9716 5776
rect 11020 5732 11060 5776
rect 355 5692 364 5732
rect 404 5692 2132 5732
rect 2188 5692 3284 5732
rect 3340 5692 4300 5732
rect 4340 5692 4349 5732
rect 4588 5692 5260 5732
rect 5300 5692 6260 5732
rect 6307 5692 6316 5732
rect 6356 5723 6548 5732
rect 6356 5692 6508 5723
rect 2188 5648 2228 5692
rect 3340 5648 3380 5692
rect 4588 5648 4628 5692
rect 6761 5692 6892 5732
rect 6932 5692 6941 5732
rect 8009 5692 8140 5732
rect 8180 5692 8189 5732
rect 8515 5692 8524 5732
rect 8564 5692 9716 5732
rect 9772 5723 9812 5732
rect 6508 5674 6548 5683
rect 8140 5648 8180 5683
rect 9772 5648 9812 5683
rect 643 5608 652 5648
rect 692 5608 1180 5648
rect 1220 5608 1229 5648
rect 1411 5608 1420 5648
rect 1460 5608 1469 5648
rect 1795 5608 1804 5648
rect 1844 5608 1996 5648
rect 2036 5608 2045 5648
rect 2179 5608 2188 5648
rect 2228 5608 2237 5648
rect 2371 5608 2380 5648
rect 2420 5608 2572 5648
rect 2612 5608 2621 5648
rect 2755 5608 2764 5648
rect 2804 5608 3284 5648
rect 3331 5608 3340 5648
rect 3380 5608 3389 5648
rect 4291 5608 4300 5648
rect 4340 5608 4628 5648
rect 4675 5608 4684 5648
rect 4724 5608 4733 5648
rect 4867 5608 4876 5648
rect 4916 5608 4924 5648
rect 4964 5608 5047 5648
rect 8140 5608 9812 5648
rect 10060 5692 10484 5732
rect 10723 5692 10732 5732
rect 10772 5692 10915 5732
rect 10955 5692 10964 5732
rect 11011 5692 11020 5732
rect 11060 5692 11069 5732
rect 11395 5692 11404 5732
rect 11444 5692 11453 5732
rect 11587 5692 11596 5732
rect 11636 5723 12020 5732
rect 11636 5692 11980 5723
rect 1420 5564 1460 5608
rect 163 5524 172 5564
rect 212 5524 1172 5564
rect 1420 5524 2092 5564
rect 2132 5524 2141 5564
rect 2995 5524 3004 5564
rect 3044 5524 3148 5564
rect 3188 5524 3197 5564
rect 0 5480 90 5500
rect 1132 5480 1172 5524
rect 0 5440 1076 5480
rect 1132 5440 1564 5480
rect 1604 5440 1613 5480
rect 1699 5440 1708 5480
rect 1748 5440 1948 5480
rect 1988 5440 1997 5480
rect 2860 5440 3100 5480
rect 3140 5440 3149 5480
rect 0 5420 90 5440
rect 1036 5396 1076 5440
rect 2860 5396 2900 5440
rect 1036 5356 2900 5396
rect 3244 5396 3284 5608
rect 4684 5564 4724 5608
rect 10060 5564 10100 5692
rect 10444 5648 10484 5692
rect 10147 5608 10156 5648
rect 10196 5608 10348 5648
rect 10388 5608 10397 5648
rect 10444 5608 11348 5648
rect 4684 5524 7948 5564
rect 7988 5524 7997 5564
rect 8323 5524 8332 5564
rect 8372 5524 9388 5564
rect 9428 5524 9437 5564
rect 9484 5524 10100 5564
rect 9484 5480 9524 5524
rect 4531 5440 4540 5480
rect 4580 5440 4780 5480
rect 4820 5440 4829 5480
rect 6569 5440 6700 5480
rect 6740 5440 6749 5480
rect 7075 5440 7084 5480
rect 7124 5440 9524 5480
rect 9955 5440 9964 5480
rect 10004 5440 10013 5480
rect 10099 5440 10108 5480
rect 10148 5440 10156 5480
rect 10196 5440 10279 5480
rect 3244 5356 7372 5396
rect 7412 5356 7421 5396
rect 3679 5272 3688 5312
rect 3728 5272 3770 5312
rect 3810 5272 3852 5312
rect 3892 5272 3934 5312
rect 3974 5272 4016 5312
rect 4056 5272 4065 5312
rect 6499 5272 6508 5312
rect 6548 5272 9004 5312
rect 9044 5272 9053 5312
rect 9964 5228 10004 5440
rect 11308 5396 11348 5608
rect 11404 5480 11444 5692
rect 12329 5692 12460 5732
rect 12500 5692 12509 5732
rect 11980 5674 12020 5683
rect 12460 5674 12500 5683
rect 12556 5648 12596 5776
rect 12940 5776 13036 5816
rect 13076 5776 13085 5816
rect 14380 5776 14476 5816
rect 14516 5776 14525 5816
rect 14572 5776 15820 5816
rect 15860 5776 15869 5816
rect 16012 5776 16820 5816
rect 12940 5732 12980 5776
rect 14380 5732 14420 5776
rect 16012 5732 16052 5776
rect 12922 5692 12931 5732
rect 12971 5692 12980 5732
rect 13027 5692 13036 5732
rect 13076 5692 13085 5732
rect 13289 5692 13420 5732
rect 13460 5692 13469 5732
rect 13865 5692 13996 5732
rect 14036 5692 14045 5732
rect 14380 5723 14516 5732
rect 14380 5692 14476 5723
rect 11491 5608 11500 5648
rect 11540 5608 11549 5648
rect 12556 5608 12980 5648
rect 11500 5564 11540 5608
rect 12940 5564 12980 5608
rect 13036 5564 13076 5692
rect 13996 5674 14036 5683
rect 14729 5692 14764 5732
rect 14804 5692 14860 5732
rect 14900 5692 14909 5732
rect 15043 5692 15052 5732
rect 15092 5692 16052 5732
rect 16108 5723 16300 5732
rect 14476 5674 14516 5683
rect 16148 5692 16300 5723
rect 16340 5692 16349 5732
rect 16483 5692 16492 5732
rect 16532 5723 16724 5732
rect 16532 5692 16684 5723
rect 16108 5674 16148 5683
rect 16684 5674 16724 5683
rect 16780 5648 16820 5776
rect 17923 5692 17932 5732
rect 17972 5692 18700 5732
rect 18740 5692 18749 5732
rect 19180 5648 19220 5944
rect 21510 5924 21600 5944
rect 19948 5692 20716 5732
rect 20756 5692 20765 5732
rect 19948 5648 19988 5692
rect 13507 5608 13516 5648
rect 13556 5608 13900 5648
rect 13940 5608 13949 5648
rect 16780 5608 18940 5648
rect 18980 5608 18989 5648
rect 19171 5608 19180 5648
rect 19220 5608 19229 5648
rect 19433 5608 19564 5648
rect 19604 5608 19613 5648
rect 19939 5608 19948 5648
rect 19988 5608 19997 5648
rect 20323 5608 20332 5648
rect 20372 5608 20908 5648
rect 20948 5608 20957 5648
rect 11491 5524 11500 5564
rect 11540 5524 12844 5564
rect 12884 5524 12893 5564
rect 12940 5524 13460 5564
rect 13987 5524 13996 5564
rect 14036 5524 19708 5564
rect 19748 5524 19757 5564
rect 13420 5480 13460 5524
rect 21510 5480 21600 5500
rect 11404 5440 12076 5480
rect 12116 5440 12125 5480
rect 12682 5440 12691 5480
rect 12731 5440 13324 5480
rect 13364 5440 13373 5480
rect 13420 5440 19324 5480
rect 19364 5440 19373 5480
rect 20083 5440 20092 5480
rect 20132 5440 20141 5480
rect 21283 5440 21292 5480
rect 21332 5440 21600 5480
rect 20092 5396 20132 5440
rect 21510 5420 21600 5440
rect 11308 5356 20132 5396
rect 11395 5272 11404 5312
rect 11444 5272 16340 5312
rect 18799 5272 18808 5312
rect 18848 5272 18890 5312
rect 18930 5272 18972 5312
rect 19012 5272 19054 5312
rect 19094 5272 19136 5312
rect 19176 5272 19185 5312
rect 835 5188 844 5228
rect 884 5188 1460 5228
rect 0 5144 90 5164
rect 1420 5144 1460 5188
rect 1804 5188 8620 5228
rect 8660 5188 8669 5228
rect 9964 5188 10060 5228
rect 10100 5188 10164 5228
rect 12067 5188 12076 5228
rect 12116 5188 13420 5228
rect 13460 5188 13469 5228
rect 0 5104 940 5144
rect 980 5104 989 5144
rect 1123 5104 1132 5144
rect 1172 5104 1180 5144
rect 1220 5104 1303 5144
rect 1420 5104 1564 5144
rect 1604 5104 1613 5144
rect 0 5084 90 5104
rect 259 5020 268 5060
rect 308 5020 1556 5060
rect 1289 4936 1420 4976
rect 1460 4936 1469 4976
rect 1516 4892 1556 5020
rect 1804 4976 1844 5188
rect 1987 5104 1996 5144
rect 2036 5104 3148 5144
rect 3188 5104 3197 5144
rect 3331 5104 3340 5144
rect 3380 5104 7468 5144
rect 7508 5104 7517 5144
rect 7913 5104 8044 5144
rect 8084 5104 8093 5144
rect 10531 5104 10540 5144
rect 10580 5104 10732 5144
rect 10772 5104 10781 5144
rect 13001 5104 13084 5144
rect 13124 5104 13132 5144
rect 13172 5104 13181 5144
rect 15811 5104 15820 5144
rect 15860 5104 15868 5144
rect 15908 5104 15991 5144
rect 16300 5060 16340 5272
rect 18595 5188 18604 5228
rect 18644 5188 19604 5228
rect 19564 5144 19604 5188
rect 16387 5104 16396 5144
rect 16436 5104 19324 5144
rect 19364 5104 19373 5144
rect 19564 5104 20092 5144
rect 20132 5104 20141 5144
rect 1948 5020 2332 5060
rect 2372 5020 2381 5060
rect 2860 5020 10156 5060
rect 10196 5020 10205 5060
rect 10444 5020 11404 5060
rect 11444 5020 11453 5060
rect 14659 5020 14668 5060
rect 14708 5020 15092 5060
rect 16300 5020 19708 5060
rect 19748 5020 19757 5060
rect 1795 4936 1804 4976
rect 1844 4936 1853 4976
rect 1948 4892 1988 5020
rect 2860 4976 2900 5020
rect 10444 4976 10484 5020
rect 2179 4936 2188 4976
rect 2228 4936 2380 4976
rect 2420 4936 2429 4976
rect 2563 4936 2572 4976
rect 2612 4936 2900 4976
rect 2947 4936 2956 4976
rect 2996 4936 7412 4976
rect 1516 4852 1988 4892
rect 6499 4852 6508 4892
rect 6548 4852 6604 4892
rect 6644 4852 6679 4892
rect 0 4808 90 4828
rect 0 4768 2716 4808
rect 2756 4768 2765 4808
rect 3139 4768 3148 4808
rect 3188 4768 7276 4808
rect 7316 4768 7325 4808
rect 0 4748 90 4768
rect 7372 4724 7412 4936
rect 10348 4936 10484 4976
rect 11299 4936 11308 4976
rect 11348 4936 11500 4976
rect 11540 4936 11549 4976
rect 12586 4936 12595 4976
rect 12635 4936 12940 4976
rect 12980 4936 12989 4976
rect 13193 4936 13324 4976
rect 13364 4936 13373 4976
rect 14467 4936 14476 4976
rect 14516 4936 14525 4976
rect 7852 4892 7892 4901
rect 10348 4892 10388 4936
rect 11884 4892 11924 4901
rect 7892 4852 8140 4892
rect 8180 4852 8189 4892
rect 8995 4852 9004 4892
rect 9044 4852 9100 4892
rect 9140 4852 9175 4892
rect 7852 4843 7892 4852
rect 10348 4843 10388 4852
rect 10444 4852 10819 4892
rect 10859 4852 10868 4892
rect 10915 4852 10924 4892
rect 10964 4852 11095 4892
rect 11395 4852 11404 4892
rect 11444 4852 11453 4892
rect 11753 4852 11884 4892
rect 11924 4852 11933 4892
rect 12067 4852 12076 4892
rect 12116 4852 12372 4892
rect 12412 4852 12421 4892
rect 12547 4852 12556 4892
rect 12596 4852 13987 4892
rect 14027 4852 14036 4892
rect 14083 4852 14092 4892
rect 14132 4852 14188 4892
rect 14228 4852 14263 4892
rect 7948 4768 10252 4808
rect 10292 4768 10301 4808
rect 7948 4724 7988 4768
rect 10444 4724 10484 4852
rect 1027 4684 1036 4724
rect 1076 4684 1948 4724
rect 1988 4684 1997 4724
rect 2083 4684 2092 4724
rect 2132 4684 4492 4724
rect 4532 4684 4541 4724
rect 7372 4684 7988 4724
rect 9859 4684 9868 4724
rect 9908 4684 10484 4724
rect 11404 4724 11444 4852
rect 11884 4843 11924 4852
rect 12172 4768 13900 4808
rect 13940 4768 13949 4808
rect 12172 4724 12212 4768
rect 14476 4724 14516 4936
rect 15052 4892 15092 5020
rect 21510 4976 21600 4996
rect 15754 4936 15763 4976
rect 15803 4936 16108 4976
rect 16148 4936 16157 4976
rect 19555 4936 19564 4976
rect 19604 4936 19613 4976
rect 19817 4936 19948 4976
rect 19988 4936 19997 4976
rect 20323 4936 20332 4976
rect 20372 4936 20428 4976
rect 20468 4936 20503 4976
rect 20620 4936 21600 4976
rect 19564 4892 19604 4936
rect 20620 4892 20660 4936
rect 21510 4916 21600 4936
rect 14563 4852 14572 4892
rect 14612 4852 14668 4892
rect 14708 4852 14743 4892
rect 15562 4852 15571 4892
rect 15611 4852 15628 4892
rect 15668 4852 15751 4892
rect 19564 4852 20660 4892
rect 15052 4808 15092 4852
rect 15052 4768 16684 4808
rect 16724 4768 16733 4808
rect 11404 4684 12212 4724
rect 12547 4684 12556 4724
rect 12596 4684 12700 4724
rect 12740 4684 12749 4724
rect 13411 4684 13420 4724
rect 13460 4684 15916 4724
rect 15956 4684 15965 4724
rect 1411 4600 1420 4640
rect 1460 4600 17548 4640
rect 17588 4600 17597 4640
rect 4919 4516 4928 4556
rect 4968 4516 5010 4556
rect 5050 4516 5092 4556
rect 5132 4516 5174 4556
rect 5214 4516 5256 4556
rect 5296 4516 5305 4556
rect 6883 4516 6892 4556
rect 6932 4516 10636 4556
rect 10676 4516 10685 4556
rect 11875 4516 11884 4556
rect 11924 4516 14668 4556
rect 14708 4516 16012 4556
rect 16052 4516 16061 4556
rect 20039 4516 20048 4556
rect 20088 4516 20130 4556
rect 20170 4516 20212 4556
rect 20252 4516 20294 4556
rect 20334 4516 20376 4556
rect 20416 4516 20425 4556
rect 0 4472 90 4492
rect 21510 4472 21600 4492
rect 0 4432 364 4472
rect 404 4432 413 4472
rect 2371 4432 2380 4472
rect 2420 4432 5300 4472
rect 6691 4432 6700 4472
rect 6740 4432 12076 4472
rect 12116 4432 12125 4472
rect 19948 4432 21600 4472
rect 0 4412 90 4432
rect 5260 4388 5300 4432
rect 1708 4348 3052 4388
rect 3092 4348 3101 4388
rect 5260 4348 7756 4388
rect 7796 4348 7805 4388
rect 8323 4348 8332 4388
rect 8372 4348 12556 4388
rect 12596 4348 12605 4388
rect 547 4264 556 4304
rect 596 4264 1180 4304
rect 1220 4264 1229 4304
rect 1315 4264 1324 4304
rect 1364 4264 1564 4304
rect 1604 4264 1613 4304
rect 0 4136 90 4156
rect 1708 4136 1748 4348
rect 1804 4264 17356 4304
rect 17396 4264 17405 4304
rect 18307 4264 18316 4304
rect 18356 4264 19708 4304
rect 19748 4264 19757 4304
rect 1804 4136 1844 4264
rect 2572 4180 2900 4220
rect 10627 4180 10636 4220
rect 10676 4180 10924 4220
rect 10964 4180 10973 4220
rect 11491 4180 11500 4220
rect 11540 4180 12172 4220
rect 12212 4180 12221 4220
rect 2572 4136 2612 4180
rect 2860 4136 2900 4180
rect 12172 4162 12212 4171
rect 19948 4136 19988 4432
rect 21510 4412 21600 4432
rect 0 4096 788 4136
rect 1411 4096 1420 4136
rect 1460 4096 1748 4136
rect 1795 4096 1804 4136
rect 1844 4096 1853 4136
rect 2057 4096 2188 4136
rect 2228 4096 2237 4136
rect 2563 4096 2572 4136
rect 2612 4096 2621 4136
rect 2755 4096 2764 4136
rect 2804 4096 2813 4136
rect 2860 4096 10828 4136
rect 10868 4096 10877 4136
rect 19939 4096 19948 4136
rect 19988 4096 19997 4136
rect 20323 4096 20332 4136
rect 20372 4096 21292 4136
rect 21332 4096 21341 4136
rect 0 4076 90 4096
rect 748 4052 788 4096
rect 2764 4052 2804 4096
rect 748 4012 1516 4052
rect 1556 4012 1565 4052
rect 1987 4012 1996 4052
rect 2036 4012 2804 4052
rect 2995 4012 3004 4052
rect 3044 4012 12980 4052
rect 17827 4012 17836 4052
rect 17876 4012 20092 4052
rect 20132 4012 20141 4052
rect 12940 3968 12980 4012
rect 21510 3968 21600 3988
rect 1939 3928 1948 3968
rect 1988 3928 1997 3968
rect 2092 3928 2332 3968
rect 2372 3928 2381 3968
rect 12329 3928 12364 3968
rect 12404 3928 12460 3968
rect 12500 3928 12509 3968
rect 12940 3928 13516 3968
rect 13556 3928 13565 3968
rect 20323 3928 20332 3968
rect 20372 3928 21600 3968
rect 1948 3884 1988 3928
rect 931 3844 940 3884
rect 980 3844 1988 3884
rect 0 3800 90 3820
rect 2092 3800 2132 3928
rect 21510 3908 21600 3928
rect 0 3760 2132 3800
rect 3679 3760 3688 3800
rect 3728 3760 3770 3800
rect 3810 3760 3852 3800
rect 3892 3760 3934 3800
rect 3974 3760 4016 3800
rect 4056 3760 4065 3800
rect 18799 3760 18808 3800
rect 18848 3760 18890 3800
rect 18930 3760 18972 3800
rect 19012 3760 19054 3800
rect 19094 3760 19136 3800
rect 19176 3760 19185 3800
rect 0 3740 90 3760
rect 1420 3676 17260 3716
rect 17300 3676 17309 3716
rect 355 3592 364 3632
rect 404 3592 1180 3632
rect 1220 3592 1229 3632
rect 0 3464 90 3484
rect 1420 3464 1460 3676
rect 1507 3592 1516 3632
rect 1556 3592 1564 3632
rect 1604 3592 1687 3632
rect 2179 3592 2188 3632
rect 2228 3592 3188 3632
rect 3763 3592 3772 3632
rect 3812 3592 8428 3632
rect 8468 3592 8477 3632
rect 8611 3592 8620 3632
rect 8660 3592 17644 3632
rect 17684 3592 17693 3632
rect 1804 3508 2668 3548
rect 2708 3508 2717 3548
rect 2956 3508 3052 3548
rect 3092 3508 3101 3548
rect 1804 3464 1844 3508
rect 2956 3464 2996 3508
rect 3148 3464 3188 3592
rect 3379 3508 3388 3548
rect 3428 3508 11980 3548
rect 12020 3508 12029 3548
rect 12940 3508 13612 3548
rect 13652 3508 13661 3548
rect 0 3424 212 3464
rect 1411 3424 1420 3464
rect 1460 3424 1469 3464
rect 1795 3424 1804 3464
rect 1844 3424 1853 3464
rect 2179 3424 2188 3464
rect 2228 3424 2237 3464
rect 2371 3424 2380 3464
rect 2420 3424 2551 3464
rect 2947 3424 2956 3464
rect 2996 3424 3005 3464
rect 3139 3424 3148 3464
rect 3188 3424 3197 3464
rect 3401 3424 3532 3464
rect 3572 3424 3581 3464
rect 0 3404 90 3424
rect 172 3296 212 3424
rect 2188 3380 2228 3424
rect 12940 3380 12980 3508
rect 20201 3424 20332 3464
rect 20372 3424 20381 3464
rect 2188 3340 12980 3380
rect 172 3256 1948 3296
rect 1988 3256 1997 3296
rect 2611 3256 2620 3296
rect 2660 3256 12748 3296
rect 12788 3256 12797 3296
rect 1795 3172 1804 3212
rect 1844 3172 2716 3212
rect 2756 3172 2765 3212
rect 18691 3172 18700 3212
rect 18740 3172 20092 3212
rect 20132 3172 20141 3212
rect 0 3128 90 3148
rect 0 3088 76 3128
rect 116 3088 125 3128
rect 1891 3088 1900 3128
rect 1940 3088 3532 3128
rect 3572 3088 3581 3128
rect 0 3068 90 3088
rect 4919 3004 4928 3044
rect 4968 3004 5010 3044
rect 5050 3004 5092 3044
rect 5132 3004 5174 3044
rect 5214 3004 5256 3044
rect 5296 3004 5305 3044
rect 8332 3004 13804 3044
rect 13844 3004 13853 3044
rect 20039 3004 20048 3044
rect 20088 3004 20130 3044
rect 20170 3004 20212 3044
rect 20252 3004 20294 3044
rect 20334 3004 20376 3044
rect 20416 3004 20425 3044
rect 67 2920 76 2960
rect 116 2920 500 2960
rect 460 2876 500 2920
rect 4492 2920 5204 2960
rect 4492 2876 4532 2920
rect 460 2836 1180 2876
rect 1220 2836 1229 2876
rect 3859 2836 3868 2876
rect 3908 2836 4108 2876
rect 4148 2836 4157 2876
rect 4243 2836 4252 2876
rect 4292 2836 4532 2876
rect 4627 2836 4636 2876
rect 4676 2836 4684 2876
rect 4724 2836 4807 2876
rect 0 2792 90 2812
rect 5164 2792 5204 2920
rect 8332 2876 8372 3004
rect 10051 2920 10060 2960
rect 10100 2920 11156 2960
rect 11116 2876 11156 2920
rect 5705 2836 5788 2876
rect 5828 2836 5836 2876
rect 5876 2836 5885 2876
rect 6163 2836 6172 2876
rect 6212 2836 8372 2876
rect 8419 2836 8428 2876
rect 8468 2836 8476 2876
rect 8516 2836 8599 2876
rect 11116 2836 14284 2876
rect 14324 2836 14333 2876
rect 0 2752 1804 2792
rect 1844 2752 1853 2792
rect 3401 2752 3484 2792
rect 3524 2752 3532 2792
rect 3572 2752 3581 2792
rect 4867 2752 4876 2792
rect 4916 2752 5020 2792
rect 5060 2752 5069 2792
rect 5164 2752 5740 2792
rect 5780 2752 5789 2792
rect 9964 2752 17164 2792
rect 17204 2752 17213 2792
rect 0 2732 90 2752
rect 9964 2624 10004 2752
rect 10147 2668 10156 2708
rect 10196 2668 11020 2708
rect 11060 2668 11069 2708
rect 11683 2668 11692 2708
rect 11732 2668 12844 2708
rect 12884 2668 12893 2708
rect 13228 2668 13420 2708
rect 13460 2668 13469 2708
rect 13699 2668 13708 2708
rect 13748 2668 15188 2708
rect 13228 2624 13268 2668
rect 15148 2624 15188 2668
rect 1289 2584 1420 2624
rect 1460 2584 1469 2624
rect 1577 2584 1708 2624
rect 1748 2584 1757 2624
rect 1961 2584 2092 2624
rect 2132 2584 2141 2624
rect 2563 2584 2572 2624
rect 2612 2584 2621 2624
rect 2755 2584 2764 2624
rect 2804 2584 2812 2624
rect 2852 2584 2935 2624
rect 3113 2584 3148 2624
rect 3188 2584 3244 2624
rect 3284 2584 3293 2624
rect 3497 2584 3628 2624
rect 3668 2584 3677 2624
rect 4003 2584 4012 2624
rect 4052 2584 4108 2624
rect 4148 2584 4183 2624
rect 4265 2584 4300 2624
rect 4340 2584 4396 2624
rect 4436 2584 4445 2624
rect 4649 2584 4684 2624
rect 4724 2584 4780 2624
rect 4820 2584 4829 2624
rect 5155 2584 5164 2624
rect 5204 2584 5356 2624
rect 5396 2584 5405 2624
rect 5452 2584 5548 2624
rect 5588 2584 5597 2624
rect 5801 2584 5836 2624
rect 5876 2584 5932 2624
rect 5972 2584 5981 2624
rect 8227 2584 8236 2624
rect 8276 2584 8285 2624
rect 9065 2584 9196 2624
rect 9236 2584 9245 2624
rect 9571 2584 9580 2624
rect 9620 2584 9676 2624
rect 9716 2584 9751 2624
rect 9955 2584 9964 2624
rect 10004 2584 10013 2624
rect 10217 2584 10348 2624
rect 10388 2584 10397 2624
rect 10601 2584 10732 2624
rect 10772 2584 10781 2624
rect 10985 2584 11116 2624
rect 11156 2584 11165 2624
rect 12259 2584 12268 2624
rect 12308 2584 12844 2624
rect 12884 2584 12893 2624
rect 13219 2584 13228 2624
rect 13268 2584 13277 2624
rect 13481 2584 13612 2624
rect 13652 2584 13661 2624
rect 13865 2584 13996 2624
rect 14036 2584 14045 2624
rect 14249 2584 14380 2624
rect 14420 2584 14429 2624
rect 14633 2584 14764 2624
rect 14804 2584 14813 2624
rect 15139 2584 15148 2624
rect 15188 2584 15197 2624
rect 15401 2584 15532 2624
rect 15572 2584 15581 2624
rect 2572 2540 2612 2584
rect 5452 2540 5492 2584
rect 8236 2540 8276 2584
rect 1939 2500 1948 2540
rect 1988 2500 2476 2540
rect 2516 2500 2525 2540
rect 2572 2500 4436 2540
rect 5443 2500 5452 2540
rect 5492 2500 5501 2540
rect 8236 2500 18700 2540
rect 18740 2500 18749 2540
rect 2323 2416 2332 2456
rect 2372 2416 4340 2456
rect 3679 2248 3688 2288
rect 3728 2248 3770 2288
rect 3810 2248 3852 2288
rect 3892 2248 3934 2288
rect 3974 2248 4016 2288
rect 4056 2248 4065 2288
rect 4300 2204 4340 2416
rect 4396 2288 4436 2500
rect 5251 2416 5260 2456
rect 5300 2416 5404 2456
rect 5444 2416 5453 2456
rect 5635 2416 5644 2456
rect 5684 2416 7276 2456
rect 7316 2416 7325 2456
rect 8825 2416 8908 2456
rect 8948 2416 8956 2456
rect 8996 2416 9005 2456
rect 9209 2416 9292 2456
rect 9332 2416 9340 2456
rect 9380 2416 9389 2456
rect 9593 2416 9676 2456
rect 9716 2416 9724 2456
rect 9764 2416 9773 2456
rect 9977 2416 10060 2456
rect 10100 2416 10108 2456
rect 10148 2416 10157 2456
rect 10361 2416 10444 2456
rect 10484 2416 10492 2456
rect 10532 2416 10541 2456
rect 10745 2416 10828 2456
rect 10868 2416 10876 2456
rect 10916 2416 10925 2456
rect 12473 2416 12556 2456
rect 12596 2416 12604 2456
rect 12644 2416 12653 2456
rect 12828 2416 12940 2456
rect 12980 2416 12988 2456
rect 13028 2416 13037 2456
rect 13241 2416 13324 2456
rect 13364 2416 13372 2456
rect 13412 2416 13421 2456
rect 13625 2416 13708 2456
rect 13748 2416 13756 2456
rect 13796 2416 13805 2456
rect 14009 2416 14092 2456
rect 14132 2416 14140 2456
rect 14180 2416 14189 2456
rect 14393 2416 14476 2456
rect 14516 2416 14524 2456
rect 14564 2416 14573 2456
rect 14777 2416 14860 2456
rect 14900 2416 14908 2456
rect 14948 2416 14957 2456
rect 15161 2416 15244 2456
rect 15284 2416 15292 2456
rect 15332 2416 15341 2456
rect 6019 2332 6028 2372
rect 6068 2332 14188 2372
rect 14228 2332 14237 2372
rect 4396 2248 17300 2288
rect 18799 2248 18808 2288
rect 18848 2248 18890 2288
rect 18930 2248 18972 2288
rect 19012 2248 19054 2288
rect 19094 2248 19136 2288
rect 19176 2248 19185 2288
rect 17260 2204 17300 2248
rect 3043 2164 3052 2204
rect 3092 2164 4052 2204
rect 4300 2164 12596 2204
rect 17260 2164 17740 2204
rect 17780 2164 17789 2204
rect 1939 2080 1948 2120
rect 1988 2080 2284 2120
rect 2324 2080 2333 2120
rect 2563 2080 2572 2120
rect 2612 2080 2812 2120
rect 2852 2080 2861 2120
rect 3331 2080 3340 2120
rect 3380 2080 3868 2120
rect 3908 2080 3917 2120
rect 4012 2036 4052 2164
rect 4195 2080 4204 2120
rect 4244 2080 4252 2120
rect 4292 2080 4375 2120
rect 5011 2080 5020 2120
rect 5060 2080 5548 2120
rect 5588 2080 5597 2120
rect 6163 2080 6172 2120
rect 6212 2080 6316 2120
rect 6356 2080 6365 2120
rect 6547 2080 6556 2120
rect 6596 2080 6700 2120
rect 6740 2080 6749 2120
rect 6883 2080 6892 2120
rect 6932 2080 7036 2120
rect 7076 2080 7085 2120
rect 7625 2080 7708 2120
rect 7748 2080 7756 2120
rect 7796 2080 7805 2120
rect 12556 2036 12596 2164
rect 12739 2080 12748 2120
rect 12788 2080 14996 2120
rect 17347 2080 17356 2120
rect 17396 2080 17404 2120
rect 17444 2080 17527 2120
rect 1324 1996 2380 2036
rect 2420 1996 2429 2036
rect 3244 1996 3724 2036
rect 3764 1996 3773 2036
rect 4012 1996 4348 2036
rect 4388 1996 4397 2036
rect 5164 1996 5644 2036
rect 5684 1996 5693 2036
rect 6931 1996 6940 2036
rect 6980 1996 7084 2036
rect 7124 1996 7133 2036
rect 7267 1996 7276 2036
rect 7316 1996 11308 2036
rect 11348 1996 11357 2036
rect 11884 1996 12460 2036
rect 12500 1996 12509 2036
rect 12556 1996 13844 2036
rect 13891 1996 13900 2036
rect 13940 1996 14716 2036
rect 14756 1996 14765 2036
rect 1324 1952 1364 1996
rect 3244 1952 3284 1996
rect 5164 1952 5204 1996
rect 11884 1952 11924 1996
rect 13804 1952 13844 1996
rect 14956 1952 14996 2080
rect 16108 1996 19468 2036
rect 19508 1996 19517 2036
rect 16108 1952 16148 1996
rect 1315 1912 1324 1952
rect 1364 1912 1373 1952
rect 1699 1912 1708 1952
rect 1748 1912 1757 1952
rect 2083 1912 2092 1952
rect 2132 1912 2141 1952
rect 2467 1912 2476 1952
rect 2516 1912 2996 1952
rect 3043 1912 3052 1952
rect 3092 1912 3101 1952
rect 3235 1912 3244 1952
rect 3284 1912 3293 1952
rect 3619 1912 3628 1952
rect 3668 1912 3677 1952
rect 4003 1912 4012 1952
rect 4052 1912 4532 1952
rect 4579 1912 4588 1952
rect 4628 1912 4637 1952
rect 4771 1912 4780 1952
rect 4820 1912 5108 1952
rect 5155 1912 5164 1952
rect 5204 1912 5213 1952
rect 5539 1912 5548 1952
rect 5588 1912 5876 1952
rect 5923 1912 5932 1952
rect 5972 1912 6260 1952
rect 6307 1912 6316 1952
rect 6356 1912 6412 1952
rect 6452 1912 6487 1952
rect 6569 1912 6604 1952
rect 6644 1912 6700 1952
rect 6740 1912 6749 1952
rect 6979 1912 6988 1952
rect 7028 1912 7276 1952
rect 7316 1912 7325 1952
rect 7459 1912 7468 1952
rect 7508 1912 7517 1952
rect 8105 1912 8236 1952
rect 8276 1912 8285 1952
rect 8489 1912 8620 1952
rect 8660 1912 8669 1952
rect 8873 1912 9004 1952
rect 9044 1912 9053 1952
rect 9257 1912 9388 1952
rect 9428 1912 9437 1952
rect 9641 1912 9772 1952
rect 9812 1912 9821 1952
rect 10025 1912 10156 1952
rect 10196 1912 10205 1952
rect 10531 1912 10540 1952
rect 10580 1912 10589 1952
rect 10793 1912 10924 1952
rect 10964 1912 10973 1952
rect 11369 1912 11500 1952
rect 11540 1912 11549 1952
rect 11875 1912 11884 1952
rect 11924 1912 11933 1952
rect 12137 1912 12268 1952
rect 12308 1912 12317 1952
rect 12521 1912 12652 1952
rect 12692 1912 12701 1952
rect 12905 1912 13036 1952
rect 13076 1912 13085 1952
rect 13289 1912 13420 1952
rect 13460 1912 13469 1952
rect 13795 1912 13804 1952
rect 13844 1912 13853 1952
rect 14057 1912 14188 1952
rect 14228 1912 14237 1952
rect 14441 1912 14572 1952
rect 14612 1912 14621 1952
rect 14947 1912 14956 1952
rect 14996 1912 15005 1952
rect 15209 1912 15340 1952
rect 15380 1912 15389 1952
rect 15593 1912 15724 1952
rect 15764 1912 15773 1952
rect 16099 1912 16108 1952
rect 16148 1912 16157 1952
rect 16361 1912 16492 1952
rect 16532 1912 16541 1952
rect 17347 1912 17356 1952
rect 17396 1912 17644 1952
rect 17684 1912 17693 1952
rect 1708 1784 1748 1912
rect 2092 1868 2132 1912
rect 2956 1868 2996 1912
rect 3052 1868 3092 1912
rect 3628 1868 3668 1912
rect 4492 1868 4532 1912
rect 4588 1868 4628 1912
rect 5068 1868 5108 1912
rect 5836 1868 5876 1912
rect 6220 1868 6260 1912
rect 7468 1868 7508 1912
rect 10540 1868 10580 1912
rect 2092 1828 2764 1868
rect 2804 1828 2813 1868
rect 2947 1828 2956 1868
rect 2996 1828 3005 1868
rect 3052 1828 3340 1868
rect 3380 1828 3389 1868
rect 3628 1828 4204 1868
rect 4244 1828 4253 1868
rect 4483 1828 4492 1868
rect 4532 1828 4541 1868
rect 4588 1828 4780 1868
rect 4820 1828 4829 1868
rect 5068 1828 5548 1868
rect 5588 1828 5597 1868
rect 5836 1828 6028 1868
rect 6068 1828 6077 1868
rect 6211 1828 6220 1868
rect 6260 1828 6269 1868
rect 6787 1828 6796 1868
rect 6836 1828 7508 1868
rect 8803 1828 8812 1868
rect 8852 1828 10580 1868
rect 1708 1744 2572 1784
rect 2612 1744 2621 1784
rect 2707 1744 2716 1784
rect 2756 1744 3244 1784
rect 3284 1744 3293 1784
rect 5395 1744 5404 1784
rect 5444 1744 9196 1784
rect 9236 1744 9245 1784
rect 11155 1744 11164 1784
rect 11204 1744 11212 1784
rect 11252 1744 11335 1784
rect 11779 1744 11788 1784
rect 11828 1744 12412 1784
rect 12452 1744 12461 1784
rect 12739 1744 12748 1784
rect 12788 1744 13564 1784
rect 13604 1744 13613 1784
rect 14659 1744 14668 1784
rect 14708 1744 15484 1784
rect 15524 1744 15533 1784
rect 1555 1660 1564 1700
rect 1604 1660 1844 1700
rect 2323 1660 2332 1700
rect 2372 1660 2476 1700
rect 2516 1660 2525 1700
rect 3475 1660 3484 1700
rect 3524 1660 3956 1700
rect 5779 1660 5788 1700
rect 5828 1660 8372 1700
rect 8467 1660 8476 1700
rect 8516 1660 8716 1700
rect 8756 1660 8765 1700
rect 8851 1660 8860 1700
rect 8900 1660 9100 1700
rect 9140 1660 9149 1700
rect 9235 1660 9244 1700
rect 9284 1660 9484 1700
rect 9524 1660 9533 1700
rect 9619 1660 9628 1700
rect 9668 1660 9868 1700
rect 9908 1660 9917 1700
rect 10003 1660 10012 1700
rect 10052 1660 10252 1700
rect 10292 1660 10301 1700
rect 10387 1660 10396 1700
rect 10436 1660 10636 1700
rect 10676 1660 10685 1700
rect 10771 1660 10780 1700
rect 10820 1660 11020 1700
rect 11060 1660 11069 1700
rect 11251 1660 11260 1700
rect 11300 1660 11404 1700
rect 11444 1660 11453 1700
rect 11513 1660 11596 1700
rect 11636 1660 11644 1700
rect 11684 1660 11693 1700
rect 11897 1660 11980 1700
rect 12020 1660 12028 1700
rect 12068 1660 12077 1700
rect 12163 1660 12172 1700
rect 12212 1660 12796 1700
rect 12836 1660 12845 1700
rect 12940 1660 13180 1700
rect 13220 1660 13229 1700
rect 13324 1660 13948 1700
rect 13988 1660 13997 1700
rect 14092 1660 14332 1700
rect 14372 1660 14381 1700
rect 14572 1660 15100 1700
rect 15140 1660 15149 1700
rect 15244 1660 15868 1700
rect 15908 1660 15917 1700
rect 16012 1660 16252 1700
rect 16292 1660 16301 1700
rect 1804 1616 1844 1660
rect 3916 1616 3956 1660
rect 8332 1616 8372 1660
rect 12940 1616 12980 1660
rect 13324 1616 13364 1660
rect 14092 1616 14132 1660
rect 14572 1616 14612 1660
rect 15244 1616 15284 1660
rect 16012 1616 16052 1660
rect 1804 1576 2900 1616
rect 3916 1576 4396 1616
rect 4436 1576 4445 1616
rect 4492 1576 6452 1616
rect 8332 1576 11692 1616
rect 11732 1576 11741 1616
rect 12355 1576 12364 1616
rect 12404 1576 12980 1616
rect 13123 1576 13132 1616
rect 13172 1576 13364 1616
rect 13507 1576 13516 1616
rect 13556 1576 14132 1616
rect 14275 1576 14284 1616
rect 14324 1576 14612 1616
rect 15043 1576 15052 1616
rect 15092 1576 15284 1616
rect 15427 1576 15436 1616
rect 15476 1576 16052 1616
rect 2860 1532 2900 1576
rect 4492 1532 4532 1576
rect 6412 1532 6452 1576
rect 2860 1492 4532 1532
rect 4919 1492 4928 1532
rect 4968 1492 5010 1532
rect 5050 1492 5092 1532
rect 5132 1492 5174 1532
rect 5214 1492 5256 1532
rect 5296 1492 5305 1532
rect 6412 1492 9964 1532
rect 10004 1492 10013 1532
rect 10723 1492 10732 1532
rect 10772 1492 17644 1532
rect 17684 1492 17693 1532
rect 20039 1492 20048 1532
rect 20088 1492 20130 1532
rect 20170 1492 20212 1532
rect 20252 1492 20294 1532
rect 20334 1492 20376 1532
rect 20416 1492 20425 1532
<< via2 >>
rect 4928 95236 4968 95276
rect 5010 95236 5050 95276
rect 5092 95236 5132 95276
rect 5174 95236 5214 95276
rect 5256 95236 5296 95276
rect 20048 95236 20088 95276
rect 20130 95236 20170 95276
rect 20212 95236 20252 95276
rect 20294 95236 20334 95276
rect 20376 95236 20416 95276
rect 13516 95068 13556 95108
rect 2572 94984 2612 95024
rect 3340 94984 3380 95024
rect 4204 94984 4244 95024
rect 4588 94984 4628 95024
rect 5644 94984 5684 95024
rect 6412 94984 6452 95024
rect 7564 94984 7604 95024
rect 7852 94984 7892 95024
rect 8332 94984 8372 95024
rect 11308 94984 11348 95024
rect 12748 94984 12788 95024
rect 15628 94984 15668 95024
rect 15916 94984 15956 95024
rect 16204 94984 16244 95024
rect 17356 94984 17396 95024
rect 8716 94900 8756 94940
rect 9100 94900 9140 94940
rect 9484 94900 9524 94940
rect 9868 94900 9908 94940
rect 10252 94900 10292 94940
rect 10636 94900 10676 94940
rect 11020 94900 11060 94940
rect 11212 94900 11252 94940
rect 11980 94900 12020 94940
rect 12172 94900 12212 94940
rect 13132 94900 13172 94940
rect 1324 94816 1364 94856
rect 1708 94816 1748 94856
rect 2092 94816 2132 94856
rect 2476 94816 2516 94856
rect 3244 94816 3284 94856
rect 3628 94816 3668 94856
rect 4012 94816 4052 94856
rect 4396 94816 4436 94856
rect 5548 94816 5588 94856
rect 5932 94816 5972 94856
rect 6316 94816 6356 94856
rect 6700 94816 6740 94856
rect 7084 94816 7124 94856
rect 11404 94816 11444 94856
rect 11596 94816 11636 94856
rect 2956 94732 2996 94772
rect 3724 94732 3764 94772
rect 4492 94732 4532 94772
rect 3148 94564 3188 94604
rect 4780 94564 4820 94604
rect 3688 94480 3728 94520
rect 3770 94480 3810 94520
rect 3852 94480 3892 94520
rect 3934 94480 3974 94520
rect 4016 94480 4056 94520
rect 6028 94732 6068 94772
rect 6796 94732 6836 94772
rect 7180 94648 7220 94688
rect 7564 94732 7604 94772
rect 8140 94732 8180 94772
rect 10732 94732 10772 94772
rect 11500 94732 11540 94772
rect 11788 94732 11828 94772
rect 12364 94732 12404 94772
rect 13228 94732 13268 94772
rect 8428 94648 8468 94688
rect 8812 94648 8852 94688
rect 9388 94648 9428 94688
rect 9772 94648 9812 94688
rect 10540 94648 10580 94688
rect 11212 94648 11252 94688
rect 11596 94648 11636 94688
rect 12172 94648 12212 94688
rect 13036 94648 13076 94688
rect 16396 94900 16436 94940
rect 17164 94900 17204 94940
rect 18124 94900 18164 94940
rect 19948 94900 19988 94940
rect 16300 94816 16340 94856
rect 16492 94816 16532 94856
rect 17068 94816 17108 94856
rect 17452 94816 17492 94856
rect 17644 94816 17684 94856
rect 18220 94816 18260 94856
rect 18604 94816 18644 94856
rect 18796 94816 18836 94856
rect 19756 94816 19796 94856
rect 14380 94732 14420 94772
rect 11788 94564 11828 94604
rect 12460 94564 12500 94604
rect 14572 94648 14612 94688
rect 14764 94648 14804 94688
rect 13420 94480 13460 94520
rect 2668 94396 2708 94436
rect 2380 94312 2420 94352
rect 2764 94312 2804 94352
rect 3532 94312 3572 94352
rect 4108 94312 4148 94352
rect 4300 94312 4340 94352
rect 4684 94312 4724 94352
rect 5356 94312 5396 94352
rect 5836 94312 5876 94352
rect 19660 94732 19700 94772
rect 16012 94648 16052 94688
rect 16588 94648 16628 94688
rect 18124 94648 18164 94688
rect 13900 94564 13940 94604
rect 15340 94564 15380 94604
rect 16492 94564 16532 94604
rect 16780 94564 16820 94604
rect 17836 94564 17876 94604
rect 17452 94480 17492 94520
rect 18220 94480 18260 94520
rect 18604 94480 18644 94520
rect 18808 94480 18848 94520
rect 18890 94480 18930 94520
rect 18972 94480 19012 94520
rect 19054 94480 19094 94520
rect 19136 94480 19176 94520
rect 6220 94312 6260 94352
rect 6604 94312 6644 94352
rect 6988 94312 7028 94352
rect 7372 94312 7412 94352
rect 7756 94312 7796 94352
rect 8524 94312 8564 94352
rect 17740 94396 17780 94436
rect 2188 94228 2228 94268
rect 5452 94228 5492 94268
rect 8908 94228 8948 94268
rect 9676 94228 9716 94268
rect 10444 94228 10484 94268
rect 12940 94228 12980 94268
rect 13708 94228 13748 94268
rect 1228 94144 1268 94184
rect 2764 94144 2804 94184
rect 3148 94144 3188 94184
rect 4588 94144 4628 94184
rect 4972 94144 5012 94184
rect 5356 94144 5396 94184
rect 5740 94144 5780 94184
rect 76 93808 116 93848
rect 2860 94060 2900 94100
rect 6124 94144 6164 94184
rect 6892 94144 6932 94184
rect 7276 94144 7316 94184
rect 8044 94144 8084 94184
rect 8236 94144 8276 94184
rect 9292 94144 9332 94184
rect 10060 94144 10100 94184
rect 10828 94144 10868 94184
rect 12556 94144 12596 94184
rect 13324 94144 13364 94184
rect 4684 94060 4724 94100
rect 7180 94060 7220 94100
rect 14476 94228 14516 94268
rect 15052 94228 15092 94268
rect 14092 94144 14132 94184
rect 15244 94144 15284 94184
rect 16204 94144 16244 94184
rect 16972 94144 17012 94184
rect 17356 94144 17396 94184
rect 17740 94144 17780 94184
rect 18124 94144 18164 94184
rect 18604 94144 18644 94184
rect 19852 94144 19892 94184
rect 20236 94144 20276 94184
rect 9484 94060 9524 94100
rect 11692 94060 11732 94100
rect 14860 94060 14900 94100
rect 18028 94060 18068 94100
rect 8140 93976 8180 94016
rect 9580 93976 9620 94016
rect 9964 93976 10004 94016
rect 11020 93976 11060 94016
rect 12076 93976 12116 94016
rect 13420 93976 13460 94016
rect 7468 93892 7508 93932
rect 7660 93892 7700 93932
rect 10156 93892 10196 93932
rect 10828 93892 10868 93932
rect 12652 93892 12692 93932
rect 12940 93892 12980 93932
rect 13900 93892 13940 93932
rect 14284 93892 14324 93932
rect 14668 93892 14708 93932
rect 15148 93892 15188 93932
rect 16588 93892 16628 93932
rect 17452 93892 17492 93932
rect 17740 93892 17780 93932
rect 19564 93892 19604 93932
rect 19756 93892 19796 93932
rect 8620 93808 8660 93848
rect 14476 93808 14516 93848
rect 17548 93808 17588 93848
rect 18316 93808 18356 93848
rect 18796 93808 18836 93848
rect 4928 93724 4968 93764
rect 5010 93724 5050 93764
rect 5092 93724 5132 93764
rect 5174 93724 5214 93764
rect 5256 93724 5296 93764
rect 7468 93724 7508 93764
rect 12268 93724 12308 93764
rect 14956 93724 14996 93764
rect 16396 93724 16436 93764
rect 18220 93724 18260 93764
rect 18988 93724 19028 93764
rect 19852 93724 19892 93764
rect 20048 93724 20088 93764
rect 20130 93724 20170 93764
rect 20212 93724 20252 93764
rect 20294 93724 20334 93764
rect 20376 93724 20416 93764
rect 76 93640 116 93680
rect 6028 93640 6068 93680
rect 14572 93640 14612 93680
rect 15436 93640 15476 93680
rect 18316 93640 18356 93680
rect 19948 93640 19988 93680
rect 172 93556 212 93596
rect 1996 93556 2036 93596
rect 18508 93556 18548 93596
rect 19660 93556 19700 93596
rect 2476 93472 2516 93512
rect 18700 93472 18740 93512
rect 172 93388 212 93428
rect 460 93304 500 93344
rect 1612 93304 1652 93344
rect 19756 93388 19796 93428
rect 18796 93304 18836 93344
rect 18988 93304 19028 93344
rect 19948 93304 19988 93344
rect 20140 93304 20180 93344
rect 4780 93220 4820 93260
rect 1228 93136 1268 93176
rect 1708 93136 1748 93176
rect 4108 93136 4148 93176
rect 3688 92968 3728 93008
rect 3770 92968 3810 93008
rect 3852 92968 3892 93008
rect 3934 92968 3974 93008
rect 4016 92968 4056 93008
rect 8716 92884 8756 92924
rect 2188 92800 2228 92840
rect 13612 92716 13652 92756
rect 1228 92632 1268 92672
rect 1420 92632 1460 92672
rect 1996 92632 2036 92672
rect 2956 92632 2996 92672
rect 1900 92548 1940 92588
rect 19084 93220 19124 93260
rect 19564 93220 19604 93260
rect 18700 93136 18740 93176
rect 21004 93136 21044 93176
rect 18808 92968 18848 93008
rect 18890 92968 18930 93008
rect 18972 92968 19012 93008
rect 19054 92968 19094 93008
rect 19136 92968 19176 93008
rect 19276 92800 19316 92840
rect 19468 92800 19508 92840
rect 19180 92632 19220 92672
rect 19468 92632 19508 92672
rect 19756 92632 19796 92672
rect 20524 92632 20564 92672
rect 21004 92632 21044 92672
rect 19660 92548 19700 92588
rect 15532 92464 15572 92504
rect 2668 92380 2708 92420
rect 6796 92380 6836 92420
rect 16012 92380 16052 92420
rect 19180 92380 19220 92420
rect 21004 92380 21044 92420
rect 3148 92296 3188 92336
rect 2956 92212 2996 92252
rect 4928 92212 4968 92252
rect 5010 92212 5050 92252
rect 5092 92212 5132 92252
rect 5174 92212 5214 92252
rect 5256 92212 5296 92252
rect 20048 92212 20088 92252
rect 20130 92212 20170 92252
rect 20212 92212 20252 92252
rect 20294 92212 20334 92252
rect 20376 92212 20416 92252
rect 1612 92128 1652 92168
rect 5932 92044 5972 92084
rect 19372 92044 19412 92084
rect 1324 91960 1364 92000
rect 1132 91876 1172 91916
rect 460 91792 500 91832
rect 748 91792 788 91832
rect 1516 91792 1556 91832
rect 8044 91792 8084 91832
rect 19564 91792 19604 91832
rect 19756 91792 19796 91832
rect 20908 91792 20948 91832
rect 1612 91624 1652 91664
rect 2188 91624 2228 91664
rect 2476 91624 2516 91664
rect 9676 91624 9716 91664
rect 20812 91624 20852 91664
rect 21004 91624 21044 91664
rect 18508 91540 18548 91580
rect 3688 91456 3728 91496
rect 3770 91456 3810 91496
rect 3852 91456 3892 91496
rect 3934 91456 3974 91496
rect 4016 91456 4056 91496
rect 18808 91456 18848 91496
rect 18890 91456 18930 91496
rect 18972 91456 19012 91496
rect 19054 91456 19094 91496
rect 19136 91456 19176 91496
rect 2572 91372 2612 91412
rect 10828 91372 10868 91412
rect 76 91288 116 91328
rect 6892 91288 6932 91328
rect 1996 91204 2036 91244
rect 7276 91204 7316 91244
rect 844 91120 884 91160
rect 2572 91120 2612 91160
rect 7948 91120 7988 91160
rect 8332 91120 8372 91160
rect 19660 91120 19700 91160
rect 20140 91120 20180 91160
rect 2380 91036 2420 91076
rect 268 90952 308 90992
rect 9964 90952 10004 90992
rect 20716 90952 20756 90992
rect 1804 90868 1844 90908
rect 3052 90868 3092 90908
rect 21004 90868 21044 90908
rect 1324 90784 1364 90824
rect 4684 90784 4724 90824
rect 6028 90784 6068 90824
rect 4928 90700 4968 90740
rect 5010 90700 5050 90740
rect 5092 90700 5132 90740
rect 5174 90700 5214 90740
rect 5256 90700 5296 90740
rect 20048 90700 20088 90740
rect 20130 90700 20170 90740
rect 20212 90700 20252 90740
rect 20294 90700 20334 90740
rect 20376 90700 20416 90740
rect 20812 90616 20852 90656
rect 4492 90532 4532 90572
rect 17068 90532 17108 90572
rect 1420 90448 1460 90488
rect 14188 90448 14228 90488
rect 652 90280 692 90320
rect 1420 90280 1460 90320
rect 2092 90280 2132 90320
rect 11404 90364 11444 90404
rect 2668 90280 2708 90320
rect 13132 90364 13172 90404
rect 15340 90364 15380 90404
rect 15628 90395 15668 90404
rect 15628 90364 15668 90395
rect 3340 90280 3380 90320
rect 3532 90280 3572 90320
rect 17260 90280 17300 90320
rect 19276 90280 19316 90320
rect 20140 90280 20180 90320
rect 1036 90196 1076 90236
rect 11020 90196 11060 90236
rect 21292 90196 21332 90236
rect 1228 90112 1268 90152
rect 2284 90112 2324 90152
rect 1420 90028 1460 90068
rect 3148 90112 3188 90152
rect 4012 90112 4052 90152
rect 4204 90112 4244 90152
rect 5740 90112 5780 90152
rect 13036 90112 13076 90152
rect 16108 90112 16148 90152
rect 20716 90112 20756 90152
rect 20812 90028 20852 90068
rect 3688 89944 3728 89984
rect 3770 89944 3810 89984
rect 3852 89944 3892 89984
rect 3934 89944 3974 89984
rect 4016 89944 4056 89984
rect 18808 89944 18848 89984
rect 18890 89944 18930 89984
rect 18972 89944 19012 89984
rect 19054 89944 19094 89984
rect 19136 89944 19176 89984
rect 1324 89860 1364 89900
rect 2668 89860 2708 89900
rect 11596 89860 11636 89900
rect 3628 89776 3668 89816
rect 11500 89776 11540 89816
rect 2092 89692 2132 89732
rect 2668 89692 2708 89732
rect 2860 89692 2900 89732
rect 10636 89692 10676 89732
rect 13228 89692 13268 89732
rect 17164 89692 17204 89732
rect 21196 89692 21236 89732
rect 940 89608 980 89648
rect 1996 89608 2036 89648
rect 2476 89608 2516 89648
rect 3436 89608 3476 89648
rect 3820 89608 3860 89648
rect 13036 89608 13076 89648
rect 13516 89608 13556 89648
rect 15340 89608 15380 89648
rect 18028 89608 18068 89648
rect 19468 89608 19508 89648
rect 19756 89608 19796 89648
rect 20140 89608 20180 89648
rect 172 89524 212 89564
rect 2092 89524 2132 89564
rect 1420 89440 1460 89480
rect 2860 89524 2900 89564
rect 4684 89524 4724 89564
rect 9292 89524 9332 89564
rect 11404 89524 11444 89564
rect 12748 89524 12788 89564
rect 13708 89524 13748 89564
rect 16780 89524 16820 89564
rect 18124 89524 18164 89564
rect 19564 89524 19604 89564
rect 3244 89440 3284 89480
rect 4012 89440 4052 89480
rect 6220 89440 6260 89480
rect 10060 89440 10100 89480
rect 12844 89440 12884 89480
rect 13804 89440 13844 89480
rect 17260 89440 17300 89480
rect 20620 89440 20660 89480
rect 1612 89356 1652 89396
rect 3052 89356 3092 89396
rect 3628 89356 3668 89396
rect 6412 89356 6452 89396
rect 14380 89356 14420 89396
rect 14860 89356 14900 89396
rect 1420 89272 1460 89312
rect 12556 89272 12596 89312
rect 17644 89356 17684 89396
rect 21100 89356 21140 89396
rect 13132 89272 13172 89312
rect 20716 89272 20756 89312
rect 3820 89188 3860 89228
rect 4928 89188 4968 89228
rect 5010 89188 5050 89228
rect 5092 89188 5132 89228
rect 5174 89188 5214 89228
rect 5256 89188 5296 89228
rect 6220 89188 6260 89228
rect 13900 89188 13940 89228
rect 20048 89188 20088 89228
rect 20130 89188 20170 89228
rect 20212 89188 20252 89228
rect 20294 89188 20334 89228
rect 20376 89188 20416 89228
rect 3532 89104 3572 89144
rect 12844 89104 12884 89144
rect 21004 89104 21044 89144
rect 5356 89020 5396 89060
rect 11692 89020 11732 89060
rect 13132 89020 13172 89060
rect 14284 89020 14324 89060
rect 3532 88936 3572 88976
rect 76 88768 116 88808
rect 1228 88852 1268 88892
rect 2764 88852 2804 88892
rect 3052 88852 3092 88892
rect 4012 88883 4052 88892
rect 4012 88852 4052 88883
rect 4396 88852 4436 88892
rect 364 88768 404 88808
rect 8716 88852 8756 88892
rect 10732 88852 10772 88892
rect 11980 88852 12020 88892
rect 460 88684 500 88724
rect 2956 88684 2996 88724
rect 12172 88852 12212 88892
rect 12844 88852 12884 88892
rect 13516 88852 13556 88892
rect 13996 88852 14036 88892
rect 16300 89020 16340 89060
rect 21484 88936 21524 88976
rect 14380 88852 14420 88892
rect 16108 88883 16148 88892
rect 16108 88852 16148 88883
rect 16780 88852 16820 88892
rect 17260 88852 17300 88892
rect 9292 88768 9332 88808
rect 10636 88768 10676 88808
rect 13132 88768 13172 88808
rect 14284 88768 14324 88808
rect 10924 88684 10964 88724
rect 13708 88684 13748 88724
rect 18604 88768 18644 88808
rect 18988 88768 19028 88808
rect 19372 88768 19412 88808
rect 19756 88768 19796 88808
rect 20140 88768 20180 88808
rect 21388 88768 21428 88808
rect 20236 88684 20276 88724
rect 76 88600 116 88640
rect 4780 88600 4820 88640
rect 6220 88600 6260 88640
rect 7084 88600 7124 88640
rect 9868 88600 9908 88640
rect 10540 88600 10580 88640
rect 13804 88600 13844 88640
rect 18700 88600 18740 88640
rect 20332 88600 20372 88640
rect 20620 88600 20660 88640
rect 1132 88432 1172 88472
rect 4396 88516 4436 88556
rect 8524 88516 8564 88556
rect 13132 88516 13172 88556
rect 13516 88516 13556 88556
rect 14284 88516 14324 88556
rect 21004 88516 21044 88556
rect 3688 88432 3728 88472
rect 3770 88432 3810 88472
rect 3852 88432 3892 88472
rect 3934 88432 3974 88472
rect 4016 88432 4056 88472
rect 10348 88432 10388 88472
rect 18808 88432 18848 88472
rect 18890 88432 18930 88472
rect 18972 88432 19012 88472
rect 19054 88432 19094 88472
rect 19136 88432 19176 88472
rect 2476 88264 2516 88304
rect 8620 88264 8660 88304
rect 12172 88264 12212 88304
rect 12748 88264 12788 88304
rect 18796 88264 18836 88304
rect 556 88180 596 88220
rect 3340 88180 3380 88220
rect 13132 88180 13172 88220
rect 4396 88096 4436 88136
rect 5452 88096 5492 88136
rect 8908 88096 8948 88136
rect 10636 88096 10676 88136
rect 10924 88096 10964 88136
rect 2764 88012 2804 88052
rect 2476 87928 2516 87968
rect 2092 87844 2132 87884
rect 2764 87844 2804 87884
rect 2572 87760 2612 87800
rect 13516 88096 13556 88136
rect 17932 88180 17972 88220
rect 3532 88012 3572 88052
rect 4012 88012 4052 88052
rect 5356 88012 5396 88052
rect 5644 88012 5684 88052
rect 5836 88012 5876 88052
rect 6220 88012 6260 88052
rect 8716 88012 8756 88052
rect 9292 88012 9332 88052
rect 10540 88012 10580 88052
rect 11980 88012 11988 88052
rect 11988 88012 12020 88052
rect 12556 88012 12596 88052
rect 13132 88012 13172 88052
rect 5548 87928 5588 87968
rect 8620 87928 8660 87968
rect 14092 88012 14132 88052
rect 11116 87928 11156 87968
rect 18220 88096 18260 88136
rect 20812 88096 20852 88136
rect 16588 88012 16628 88052
rect 18124 88012 18164 88052
rect 18508 88012 18548 88052
rect 15628 87928 15668 87968
rect 19276 87928 19316 87968
rect 20236 87928 20276 87968
rect 5356 87844 5396 87884
rect 5932 87844 5972 87884
rect 7372 87844 7412 87884
rect 9292 87844 9332 87884
rect 11308 87844 11348 87884
rect 12748 87844 12788 87884
rect 15340 87844 15380 87884
rect 19852 87844 19892 87884
rect 4492 87760 4532 87800
rect 9196 87760 9236 87800
rect 12844 87760 12884 87800
rect 4928 87676 4968 87716
rect 5010 87676 5050 87716
rect 5092 87676 5132 87716
rect 5174 87676 5214 87716
rect 5256 87676 5296 87716
rect 10060 87676 10100 87716
rect 10444 87676 10484 87716
rect 17836 87676 17876 87716
rect 9868 87592 9908 87632
rect 12940 87592 12980 87632
rect 6604 87508 6644 87548
rect 8716 87508 8756 87548
rect 1516 87424 1556 87464
rect 2476 87424 2516 87464
rect 5548 87424 5588 87464
rect 7084 87424 7124 87464
rect 2860 87371 2900 87380
rect 2860 87340 2900 87371
rect 3052 87340 3092 87380
rect 4780 87340 4820 87380
rect 5164 87340 5204 87380
rect 5452 87340 5492 87380
rect 5836 87340 5876 87380
rect 1324 87256 1364 87296
rect 3340 87256 3380 87296
rect 3628 87256 3668 87296
rect 1612 87172 1652 87212
rect 6412 87371 6452 87380
rect 6412 87340 6452 87371
rect 7948 87340 7988 87380
rect 5644 87256 5684 87296
rect 7084 87256 7124 87296
rect 5260 87172 5300 87212
rect 12364 87508 12404 87548
rect 13036 87508 13076 87548
rect 13324 87508 13364 87548
rect 13132 87424 13172 87464
rect 20048 87676 20088 87716
rect 20130 87676 20170 87716
rect 20212 87676 20252 87716
rect 20294 87676 20334 87716
rect 20376 87676 20416 87716
rect 20236 87508 20276 87548
rect 17452 87424 17483 87464
rect 17483 87424 17492 87464
rect 12172 87340 12212 87380
rect 10732 87256 10772 87296
rect 16588 87340 16628 87380
rect 17260 87340 17300 87380
rect 17644 87340 17675 87380
rect 17675 87340 17684 87380
rect 18316 87340 18356 87380
rect 18604 87340 18644 87380
rect 19276 87340 19316 87380
rect 18412 87256 18452 87296
rect 19756 87256 19796 87296
rect 20140 87256 20180 87296
rect 21484 87256 21524 87296
rect 8812 87172 8852 87212
rect 13324 87172 13364 87212
rect 17740 87172 17780 87212
rect 748 87088 788 87128
rect 1516 87088 1556 87128
rect 3052 87088 3092 87128
rect 3340 87088 3380 87128
rect 3532 87088 3572 87128
rect 5452 87088 5492 87128
rect 6412 87088 6452 87128
rect 9388 87088 9428 87128
rect 11308 87088 11348 87128
rect 13228 87088 13268 87128
rect 17644 87088 17684 87128
rect 17836 87088 17876 87128
rect 18124 87088 18164 87128
rect 18604 87088 18644 87128
rect 20716 87088 20756 87128
rect 9100 87004 9140 87044
rect 3688 86920 3728 86960
rect 3770 86920 3810 86960
rect 3852 86920 3892 86960
rect 3934 86920 3974 86960
rect 4016 86920 4056 86960
rect 10732 86836 10772 86876
rect 1420 86752 1460 86792
rect 2764 86752 2804 86792
rect 5644 86752 5684 86792
rect 8908 86752 8948 86792
rect 10060 86752 10100 86792
rect 10444 86752 10484 86792
rect 11212 86752 11252 86792
rect 12364 86752 12404 86792
rect 1612 86668 1652 86708
rect 3436 86668 3476 86708
rect 4492 86668 4532 86708
rect 5548 86668 5588 86708
rect 6124 86668 6164 86708
rect 11692 86668 11732 86708
rect 2860 86584 2900 86624
rect 5164 86584 5204 86624
rect 6028 86584 6068 86624
rect 7180 86584 7220 86624
rect 7852 86584 7892 86624
rect 1132 86080 1172 86120
rect 1612 86500 1652 86540
rect 4012 86500 4052 86540
rect 5260 86500 5300 86540
rect 5644 86500 5684 86540
rect 5836 86500 5876 86540
rect 7372 86500 7412 86540
rect 7948 86500 7988 86540
rect 9292 86584 9332 86624
rect 8236 86500 8276 86540
rect 8620 86500 8660 86540
rect 13036 86668 13076 86708
rect 12940 86584 12980 86624
rect 13228 86584 13268 86624
rect 18808 86920 18848 86960
rect 18890 86920 18930 86960
rect 18972 86920 19012 86960
rect 19054 86920 19094 86960
rect 19136 86920 19176 86960
rect 20908 86752 20948 86792
rect 17260 86584 17300 86624
rect 18412 86584 18452 86624
rect 19756 86584 19796 86624
rect 20140 86584 20180 86624
rect 21292 86584 21332 86624
rect 10636 86500 10676 86540
rect 12172 86500 12212 86540
rect 13612 86500 13652 86540
rect 15532 86500 15572 86540
rect 17740 86500 17780 86540
rect 18124 86500 18164 86540
rect 18316 86500 18356 86540
rect 18700 86500 18740 86540
rect 6124 86416 6164 86456
rect 7084 86416 7124 86456
rect 8716 86416 8756 86456
rect 13036 86416 13076 86456
rect 13228 86416 13268 86456
rect 15340 86416 15380 86456
rect 16972 86416 17012 86456
rect 17452 86416 17492 86456
rect 17932 86416 17972 86456
rect 18796 86416 18836 86456
rect 20716 86416 20756 86456
rect 5452 86332 5492 86372
rect 6412 86332 6452 86372
rect 6700 86332 6740 86372
rect 12556 86332 12596 86372
rect 19948 86332 19988 86372
rect 20236 86332 20276 86372
rect 21292 86332 21332 86372
rect 3244 86248 3284 86288
rect 4012 86248 4052 86288
rect 4780 86248 4820 86288
rect 15724 86248 15764 86288
rect 4928 86164 4968 86204
rect 5010 86164 5050 86204
rect 5092 86164 5132 86204
rect 5174 86164 5214 86204
rect 5256 86164 5296 86204
rect 1420 86080 1460 86120
rect 2476 86080 2516 86120
rect 4396 86080 4436 86120
rect 12460 86164 12500 86204
rect 15244 86164 15284 86204
rect 20048 86164 20088 86204
rect 20130 86164 20170 86204
rect 20212 86164 20252 86204
rect 20294 86164 20334 86204
rect 20376 86164 20416 86204
rect 12844 86080 12884 86120
rect 17932 86080 17972 86120
rect 18124 86080 18164 86120
rect 21004 86080 21044 86120
rect 1228 85996 1268 86036
rect 2380 85996 2420 86036
rect 5836 85996 5876 86036
rect 8620 85996 8660 86036
rect 12556 85996 12596 86036
rect 14284 85996 14324 86036
rect 12748 85912 12788 85952
rect 13612 85912 13652 85952
rect 16492 85912 16532 85952
rect 2380 85828 2420 85868
rect 2860 85828 2900 85868
rect 4780 85828 4820 85868
rect 1228 85744 1268 85784
rect 2476 85660 2516 85700
rect 7180 85828 7220 85868
rect 6508 85744 6548 85784
rect 4492 85660 4532 85700
rect 6700 85660 6740 85700
rect 8812 85828 8852 85868
rect 10252 85828 10292 85868
rect 9004 85744 9044 85784
rect 11884 85828 11924 85868
rect 12364 85828 12404 85868
rect 14092 85828 14132 85868
rect 15052 85859 15092 85868
rect 15052 85828 15092 85859
rect 15532 85828 15572 85868
rect 8812 85660 8852 85700
rect 18508 85828 18548 85868
rect 13036 85744 13076 85784
rect 13612 85744 13652 85784
rect 17452 85744 17492 85784
rect 17836 85744 17876 85784
rect 18412 85744 18452 85784
rect 15820 85660 15860 85700
rect 16684 85660 16724 85700
rect 18220 85660 18260 85700
rect 2572 85576 2612 85616
rect 8908 85576 8948 85616
rect 10444 85576 10484 85616
rect 12556 85576 12596 85616
rect 12844 85576 12875 85616
rect 12875 85576 12884 85616
rect 20044 85828 20084 85868
rect 14380 85576 14420 85616
rect 18124 85576 18164 85616
rect 19372 85576 19412 85616
rect 21196 85576 21236 85616
rect 4300 85492 4340 85532
rect 14860 85492 14900 85532
rect 268 85408 308 85448
rect 3688 85408 3728 85448
rect 3770 85408 3810 85448
rect 3852 85408 3892 85448
rect 3934 85408 3974 85448
rect 4016 85408 4056 85448
rect 4396 85408 4436 85448
rect 10636 85408 10676 85448
rect 12364 85408 12404 85448
rect 12748 85408 12788 85448
rect 1420 85324 1460 85364
rect 2860 85240 2900 85280
rect 5452 85240 5492 85280
rect 3244 85156 3284 85196
rect 844 85072 884 85112
rect 4780 85156 4820 85196
rect 8716 85240 8756 85280
rect 9868 85240 9908 85280
rect 10540 85240 10580 85280
rect 8524 85156 8564 85196
rect 13132 85156 13172 85196
rect 4396 85072 4436 85112
rect 7180 85072 7220 85112
rect 7468 85072 7508 85112
rect 7756 85072 7796 85112
rect 9004 85072 9044 85112
rect 12364 85072 12404 85112
rect 12748 85072 12788 85112
rect 13996 85072 14036 85112
rect 15628 85072 15668 85112
rect 15820 85072 15860 85112
rect 18604 85492 18644 85532
rect 18808 85408 18848 85448
rect 18890 85408 18930 85448
rect 18972 85408 19012 85448
rect 19054 85408 19094 85448
rect 19136 85408 19176 85448
rect 17068 85156 17108 85196
rect 21292 85072 21332 85112
rect 1612 84988 1652 85028
rect 2860 84988 2900 85028
rect 3340 84988 3380 85028
rect 4108 84988 4148 85028
rect 5548 84988 5588 85028
rect 7564 84988 7604 85028
rect 7852 84988 7892 85028
rect 8044 84988 8084 85028
rect 9292 84988 9332 85028
rect 10252 84988 10292 85028
rect 10636 84988 10676 85028
rect 11884 84988 11924 85028
rect 12460 84988 12500 85028
rect 12940 84988 12980 85028
rect 15244 84988 15284 85028
rect 15724 84988 15764 85028
rect 18124 84988 18164 85028
rect 20044 84988 20084 85028
rect 3628 84904 3668 84944
rect 7660 84904 7700 84944
rect 8332 84904 8372 84944
rect 2956 84820 2996 84860
rect 6700 84820 6740 84860
rect 6892 84820 6932 84860
rect 1420 84736 1460 84776
rect 14188 84904 14228 84944
rect 8140 84820 8180 84860
rect 9292 84820 9332 84860
rect 10444 84820 10484 84860
rect 12940 84820 12980 84860
rect 13612 84820 13652 84860
rect 14668 84820 14708 84860
rect 16108 84820 16148 84860
rect 16876 84820 16916 84860
rect 18508 84820 18548 84860
rect 20716 84820 20756 84860
rect 8524 84736 8564 84776
rect 8908 84736 8948 84776
rect 11692 84736 11732 84776
rect 12460 84736 12500 84776
rect 3628 84652 3668 84692
rect 4928 84652 4968 84692
rect 5010 84652 5050 84692
rect 5092 84652 5132 84692
rect 5174 84652 5214 84692
rect 5256 84652 5296 84692
rect 15628 84652 15668 84692
rect 17932 84652 17972 84692
rect 20048 84652 20088 84692
rect 20130 84652 20170 84692
rect 20212 84652 20252 84692
rect 20294 84652 20334 84692
rect 20376 84652 20416 84692
rect 6028 84568 6068 84608
rect 7468 84568 7508 84608
rect 20908 84568 20948 84608
rect 5548 84484 5588 84524
rect 5740 84484 5780 84524
rect 7852 84484 7892 84524
rect 11980 84484 12020 84524
rect 12364 84484 12404 84524
rect 14380 84484 14420 84524
rect 14860 84484 14900 84524
rect 16876 84484 16916 84524
rect 2188 84400 2228 84440
rect 2764 84400 2804 84440
rect 3340 84400 3380 84440
rect 3436 84316 3476 84356
rect 268 84232 308 84272
rect 1420 84232 1460 84272
rect 2188 84232 2228 84272
rect 2764 84232 2804 84272
rect 3244 84232 3284 84272
rect 3724 84316 3764 84356
rect 4300 84347 4340 84356
rect 4300 84316 4340 84347
rect 844 84148 884 84188
rect 5644 84400 5684 84440
rect 6700 84400 6740 84440
rect 4684 84316 4724 84356
rect 8332 84400 8372 84440
rect 12940 84400 12980 84440
rect 13708 84400 13748 84440
rect 14284 84400 14315 84440
rect 14315 84400 14324 84440
rect 14668 84400 14708 84440
rect 15340 84400 15380 84440
rect 16588 84400 16628 84440
rect 18508 84400 18548 84440
rect 5836 84316 5876 84356
rect 6028 84316 6068 84356
rect 6988 84347 7028 84356
rect 6988 84316 7028 84347
rect 7468 84347 7508 84356
rect 7468 84316 7508 84347
rect 7852 84316 7892 84356
rect 8524 84316 8564 84356
rect 8908 84316 8948 84356
rect 9772 84316 9812 84356
rect 10252 84316 10292 84356
rect 4492 84232 4532 84272
rect 7660 84232 7700 84272
rect 5644 84148 5684 84188
rect 10636 84316 10676 84356
rect 11500 84316 11540 84356
rect 11884 84316 11924 84356
rect 12556 84316 12596 84356
rect 13132 84316 13172 84356
rect 14380 84316 14420 84356
rect 14860 84316 14900 84356
rect 15244 84316 15284 84356
rect 15628 84316 15668 84356
rect 15820 84316 15860 84356
rect 10828 84232 10868 84272
rect 13036 84232 13076 84272
rect 15724 84232 15764 84272
rect 16972 84316 17012 84356
rect 17932 84316 17972 84356
rect 18700 84316 18740 84356
rect 19372 84347 19412 84356
rect 19372 84316 19412 84347
rect 18124 84232 18164 84272
rect 20140 84232 20180 84272
rect 8332 84148 8372 84188
rect 14668 84148 14708 84188
rect 16300 84148 16340 84188
rect 17740 84148 17780 84188
rect 19372 84148 19412 84188
rect 1612 84064 1652 84104
rect 1900 84064 1940 84104
rect 3628 84064 3668 84104
rect 8524 84064 8564 84104
rect 2668 83980 2708 84020
rect 2860 83980 2900 84020
rect 11212 84064 11252 84104
rect 13708 84064 13748 84104
rect 14188 84064 14228 84104
rect 20044 84064 20084 84104
rect 20908 84064 20948 84104
rect 21100 84064 21140 84104
rect 3688 83896 3728 83936
rect 3770 83896 3810 83936
rect 3852 83896 3892 83936
rect 3934 83896 3974 83936
rect 4016 83896 4056 83936
rect 16972 83980 17012 84020
rect 17260 83980 17300 84020
rect 21292 83980 21332 84020
rect 9292 83896 9332 83936
rect 12556 83896 12596 83936
rect 18808 83896 18848 83936
rect 18890 83896 18930 83936
rect 18972 83896 19012 83936
rect 19054 83896 19094 83936
rect 19136 83896 19176 83936
rect 7756 83812 7796 83852
rect 11404 83812 11444 83852
rect 13420 83812 13460 83852
rect 15724 83812 15764 83852
rect 18124 83812 18164 83852
rect 2764 83728 2804 83768
rect 3244 83728 3284 83768
rect 3820 83728 3860 83768
rect 4396 83728 4436 83768
rect 5260 83728 5300 83768
rect 6892 83728 6932 83768
rect 7564 83728 7604 83768
rect 12748 83728 12788 83768
rect 13996 83728 14036 83768
rect 16300 83728 16340 83768
rect 17836 83728 17876 83768
rect 3052 83644 3092 83684
rect 8044 83644 8084 83684
rect 10636 83644 10676 83684
rect 12844 83644 12884 83684
rect 14284 83644 14324 83684
rect 16684 83644 16724 83684
rect 16972 83644 17012 83684
rect 18124 83644 18164 83684
rect 1900 83476 1940 83516
rect 2764 83476 2804 83516
rect 3436 83560 3476 83600
rect 6988 83560 7028 83600
rect 8524 83560 8564 83600
rect 3724 83476 3764 83516
rect 4396 83476 4436 83516
rect 4780 83476 4820 83516
rect 5836 83476 5876 83516
rect 6796 83476 6836 83516
rect 7468 83476 7508 83516
rect 1036 83392 1076 83432
rect 3340 83392 3380 83432
rect 8332 83476 8372 83516
rect 7372 83392 7412 83432
rect 7660 83392 7700 83432
rect 8524 83392 8564 83432
rect 2956 83308 2996 83348
rect 11212 83560 11252 83600
rect 11980 83560 12020 83600
rect 9964 83476 10004 83516
rect 10828 83476 10868 83516
rect 11404 83476 11444 83516
rect 11692 83476 11732 83516
rect 12076 83476 12116 83516
rect 12556 83560 12596 83600
rect 13900 83560 13940 83600
rect 15052 83560 15092 83600
rect 15916 83560 15956 83600
rect 17836 83560 17876 83600
rect 652 83140 692 83180
rect 4928 83140 4968 83180
rect 5010 83140 5050 83180
rect 5092 83140 5132 83180
rect 5174 83140 5214 83180
rect 5256 83140 5296 83180
rect 5644 83140 5684 83180
rect 18988 83728 19028 83768
rect 21196 83728 21236 83768
rect 18700 83644 18740 83684
rect 19564 83644 19604 83684
rect 19852 83560 19892 83600
rect 20140 83560 20180 83600
rect 21196 83560 21236 83600
rect 15820 83476 15860 83516
rect 16012 83476 16052 83516
rect 17260 83476 17300 83516
rect 17932 83476 17972 83516
rect 12268 83392 12308 83432
rect 8044 83140 8084 83180
rect 8428 83140 8468 83180
rect 4396 83056 4436 83096
rect 4684 83056 4724 83096
rect 13804 83056 13844 83096
rect 4972 82972 5012 83012
rect 7564 82972 7604 83012
rect 8332 82972 8372 83012
rect 14284 82972 14324 83012
rect 14764 83056 14804 83096
rect 15052 83392 15092 83432
rect 19084 83392 19124 83432
rect 19852 83392 19892 83432
rect 15340 83308 15380 83348
rect 20048 83140 20088 83180
rect 20130 83140 20170 83180
rect 20212 83140 20252 83180
rect 20294 83140 20334 83180
rect 20376 83140 20416 83180
rect 21388 83056 21428 83096
rect 17740 82972 17780 83012
rect 2764 82888 2804 82928
rect 2860 82804 2900 82844
rect 3340 82804 3380 82844
rect 4300 82835 4340 82844
rect 4300 82804 4340 82835
rect 3532 82720 3572 82760
rect 4204 82720 4244 82760
rect 6220 82804 6260 82844
rect 7372 82804 7412 82844
rect 2764 82636 2804 82676
rect 3244 82636 3284 82676
rect 3820 82636 3860 82676
rect 8524 82720 8564 82760
rect 10252 82804 10292 82844
rect 10444 82804 10484 82844
rect 11788 82804 11828 82844
rect 11980 82804 12020 82844
rect 12268 82804 12308 82844
rect 12748 82804 12788 82844
rect 11404 82720 11444 82760
rect 11692 82720 11732 82760
rect 14764 82888 14804 82928
rect 13804 82804 13844 82844
rect 15628 82804 15668 82844
rect 15916 82804 15956 82844
rect 16972 82804 17012 82844
rect 17740 82804 17780 82844
rect 18508 82804 18548 82844
rect 14092 82720 14132 82760
rect 14668 82720 14691 82760
rect 14691 82720 14708 82760
rect 15148 82720 15188 82760
rect 15340 82720 15380 82760
rect 16204 82720 16244 82760
rect 8428 82636 8468 82676
rect 13036 82636 13076 82676
rect 14284 82636 14324 82676
rect 16012 82636 16052 82676
rect 21100 82636 21140 82676
rect 4300 82552 4340 82592
rect 6124 82552 6164 82592
rect 6796 82552 6836 82592
rect 12556 82552 12596 82592
rect 18316 82552 18356 82592
rect 18508 82552 18548 82592
rect 6508 82468 6548 82508
rect 3688 82384 3728 82424
rect 3770 82384 3810 82424
rect 3852 82384 3892 82424
rect 3934 82384 3974 82424
rect 4016 82384 4056 82424
rect 6892 82384 6932 82424
rect 14956 82384 14996 82424
rect 18808 82384 18848 82424
rect 18890 82384 18930 82424
rect 18972 82384 19012 82424
rect 19054 82384 19094 82424
rect 19136 82384 19176 82424
rect 652 82300 692 82340
rect 1420 82300 1460 82340
rect 1900 82300 1940 82340
rect 16492 82300 16532 82340
rect 1036 82216 1076 82256
rect 4396 82216 4436 82256
rect 8140 82216 8180 82256
rect 13036 82216 13076 82256
rect 14380 82216 14420 82256
rect 15148 82216 15188 82256
rect 2764 82132 2804 82172
rect 7468 82132 7508 82172
rect 13804 82132 13844 82172
rect 1420 82048 1460 82088
rect 2860 82048 2900 82088
rect 3628 82048 3668 82088
rect 4012 82048 4052 82088
rect 6508 82048 6548 82088
rect 1996 81964 2036 82004
rect 2476 81964 2516 82004
rect 2956 81964 2996 82004
rect 3340 81964 3380 82004
rect 3820 81964 3860 82004
rect 4396 81964 4436 82004
rect 5356 81964 5396 82004
rect 6700 81964 6740 82004
rect 7276 81964 7316 82004
rect 7564 81964 7604 82004
rect 8428 82048 8468 82088
rect 8908 82048 8948 82088
rect 9100 82048 9140 82088
rect 11788 82048 11828 82088
rect 13516 82048 13556 82088
rect 14380 82048 14420 82088
rect 15052 82048 15092 82088
rect 18124 82048 18164 82088
rect 18892 82048 18932 82088
rect 9964 81964 10004 82004
rect 10252 81964 10292 82004
rect 3148 81880 3188 81920
rect 3724 81880 3764 81920
rect 6988 81880 7028 81920
rect 7180 81880 7220 81920
rect 3436 81796 3476 81836
rect 4972 81796 5012 81836
rect 7084 81796 7115 81836
rect 7115 81796 7124 81836
rect 76 81712 116 81752
rect 8428 81880 8468 81920
rect 8332 81796 8372 81836
rect 7852 81712 7892 81752
rect 11404 81964 11444 82004
rect 11692 81964 11732 82004
rect 12364 81964 12404 82004
rect 12556 81964 12596 82004
rect 13036 81964 13076 82004
rect 13804 81964 13844 82004
rect 14092 81964 14132 82004
rect 14476 81964 14516 82004
rect 14956 81964 14996 82004
rect 15340 81964 15380 82004
rect 15628 81964 15668 82004
rect 16012 81964 16052 82004
rect 16684 81964 16724 82004
rect 16972 81964 17012 82004
rect 18316 81964 18356 82004
rect 18988 81964 19028 82004
rect 19180 81964 19220 82004
rect 19660 81964 19700 82004
rect 13996 81880 14036 81920
rect 16780 81880 16820 81920
rect 17068 81880 17108 81920
rect 11884 81796 11924 81836
rect 15916 81796 15956 81836
rect 18316 81796 18356 81836
rect 21388 81796 21428 81836
rect 10732 81712 10772 81752
rect 4928 81628 4968 81668
rect 5010 81628 5050 81668
rect 5092 81628 5132 81668
rect 5174 81628 5214 81668
rect 5256 81628 5296 81668
rect 7468 81628 7508 81668
rect 4684 81460 4724 81500
rect 7180 81460 7220 81500
rect 7852 81460 7883 81500
rect 7883 81460 7892 81500
rect 9484 81460 9524 81500
rect 10828 81460 10868 81500
rect 172 81376 212 81416
rect 2476 81376 2516 81416
rect 4108 81376 4148 81416
rect 5836 81376 5876 81416
rect 6412 81376 6452 81416
rect 7660 81376 7700 81416
rect 2860 81323 2900 81332
rect 2860 81292 2900 81323
rect 3532 81292 3572 81332
rect 3820 81292 3860 81332
rect 4972 81292 5012 81332
rect 5356 81292 5396 81332
rect 5932 81323 5972 81332
rect 5932 81292 5972 81323
rect 6124 81292 6164 81332
rect 6700 81292 6740 81332
rect 7180 81292 7211 81332
rect 7211 81292 7220 81332
rect 7372 81292 7412 81332
rect 7852 81292 7892 81332
rect 8428 81292 8459 81332
rect 8459 81292 8468 81332
rect 8812 81292 8852 81332
rect 13516 81712 13556 81752
rect 15724 81712 15764 81752
rect 18028 81712 18068 81752
rect 18604 81712 18644 81752
rect 20048 81628 20088 81668
rect 20130 81628 20170 81668
rect 20212 81628 20252 81668
rect 20294 81628 20334 81668
rect 20376 81628 20416 81668
rect 18220 81544 18260 81584
rect 14860 81460 14900 81500
rect 15820 81460 15860 81500
rect 17548 81460 17588 81500
rect 19084 81460 19124 81500
rect 14668 81376 14708 81416
rect 16204 81376 16244 81416
rect 18220 81376 18260 81416
rect 18508 81376 18548 81416
rect 76 81208 116 81248
rect 3244 81208 3284 81248
rect 3628 81208 3668 81248
rect 4108 81208 4148 81248
rect 4396 81208 4436 81248
rect 11404 81292 11444 81332
rect 11788 81292 11828 81332
rect 12364 81323 12404 81332
rect 12364 81292 12404 81323
rect 10444 81208 10484 81248
rect 11692 81208 11732 81248
rect 3724 81124 3764 81164
rect 13708 81292 13748 81332
rect 14764 81323 14804 81332
rect 14764 81292 14804 81323
rect 15724 81292 15764 81332
rect 18604 81292 18644 81332
rect 18892 81292 18932 81332
rect 19180 81292 19220 81332
rect 14380 81124 14420 81164
rect 17260 81208 17300 81248
rect 17932 81208 17972 81248
rect 18508 81208 18548 81248
rect 18988 81208 19028 81248
rect 16780 81124 16820 81164
rect 19372 81124 19412 81164
rect 20716 81292 20756 81332
rect 940 81040 980 81080
rect 1996 81040 2036 81080
rect 3052 81040 3092 81080
rect 7564 81040 7604 81080
rect 15148 81040 15188 81080
rect 18604 81040 18644 81080
rect 21004 81040 21044 81080
rect 17932 80956 17972 80996
rect 18316 80956 18356 80996
rect 3688 80872 3728 80912
rect 3770 80872 3810 80912
rect 3852 80872 3892 80912
rect 3934 80872 3974 80912
rect 4016 80872 4056 80912
rect 7276 80872 7316 80912
rect 8908 80872 8948 80912
rect 18808 80872 18848 80912
rect 18890 80872 18930 80912
rect 18972 80872 19012 80912
rect 19054 80872 19094 80912
rect 19136 80872 19176 80912
rect 1420 80788 1460 80828
rect 2188 80788 2228 80828
rect 14284 80788 14324 80828
rect 1132 80704 1172 80744
rect 6700 80704 6740 80744
rect 6028 80620 6068 80660
rect 748 80536 788 80576
rect 3628 80536 3668 80576
rect 11212 80620 11252 80660
rect 7084 80536 7124 80576
rect 18988 80704 19028 80744
rect 18316 80620 18356 80660
rect 20716 80620 20756 80660
rect 21388 80620 21428 80660
rect 10444 80536 10484 80576
rect 12748 80536 12788 80576
rect 13708 80536 13748 80576
rect 15532 80536 15572 80576
rect 16972 80536 17012 80576
rect 17548 80536 17588 80576
rect 18124 80536 18164 80576
rect 21484 80536 21524 80576
rect 1132 80452 1172 80492
rect 2476 80452 2516 80492
rect 2860 80452 2900 80492
rect 3148 80452 3188 80492
rect 4300 80452 4340 80492
rect 10732 80452 10772 80492
rect 11980 80452 12020 80492
rect 13324 80452 13364 80492
rect 14764 80452 14804 80492
rect 15916 80452 15956 80492
rect 652 80368 692 80408
rect 4204 80284 4244 80324
rect 652 80200 692 80240
rect 6028 80368 6068 80408
rect 7852 80368 7892 80408
rect 10060 80368 10100 80408
rect 10636 80368 10676 80408
rect 11788 80368 11828 80408
rect 12268 80368 12308 80408
rect 15340 80368 15380 80408
rect 16780 80452 16820 80492
rect 6508 80284 6548 80324
rect 7468 80284 7508 80324
rect 12172 80284 12212 80324
rect 12364 80284 12404 80324
rect 12748 80284 12788 80324
rect 14284 80284 14324 80324
rect 16300 80284 16340 80324
rect 16780 80284 16820 80324
rect 1612 80200 1652 80240
rect 4684 80200 4724 80240
rect 7564 80200 7604 80240
rect 4928 80116 4968 80156
rect 5010 80116 5050 80156
rect 5092 80116 5132 80156
rect 5174 80116 5214 80156
rect 5256 80116 5296 80156
rect 460 80032 500 80072
rect 5260 79948 5300 79988
rect 7468 79948 7508 79988
rect 3052 79864 3092 79904
rect 3340 79864 3380 79904
rect 5452 79864 5492 79904
rect 5836 79864 5876 79904
rect 18028 80452 18068 80492
rect 18796 80452 18836 80492
rect 20044 80368 20084 80408
rect 17836 80284 17876 80324
rect 18412 80284 18452 80324
rect 9292 80116 9332 80156
rect 10636 80116 10676 80156
rect 13228 80116 13268 80156
rect 9580 79948 9620 79988
rect 11788 79948 11828 79988
rect 1804 79780 1844 79820
rect 2764 79811 2804 79820
rect 2764 79780 2804 79811
rect 3148 79780 3179 79820
rect 3179 79780 3188 79820
rect 364 79696 404 79736
rect 3052 79696 3092 79736
rect 3532 79696 3572 79736
rect 6028 79780 6068 79820
rect 7372 79780 7412 79820
rect 7852 79780 7892 79820
rect 8236 79780 8276 79820
rect 8812 79811 8852 79820
rect 8812 79780 8852 79811
rect 9676 79864 9716 79904
rect 12844 79864 12884 79904
rect 14188 79864 14228 79904
rect 7468 79696 7508 79736
rect 10732 79780 10772 79820
rect 11692 79780 11732 79820
rect 11980 79780 12020 79820
rect 13324 79780 13364 79820
rect 14092 79780 14132 79820
rect 14380 79811 14420 79820
rect 14380 79780 14420 79811
rect 15340 79780 15380 79820
rect 9676 79696 9716 79736
rect 11212 79696 11252 79736
rect 11788 79696 11828 79736
rect 9292 79612 9332 79652
rect 556 79360 596 79400
rect 2956 79528 2996 79568
rect 7276 79528 7316 79568
rect 12556 79696 12596 79736
rect 12940 79696 12980 79736
rect 13228 79696 13268 79736
rect 15820 79780 15860 79820
rect 16492 79780 16532 79820
rect 18796 79780 18836 79820
rect 20048 80116 20088 80156
rect 20130 80116 20170 80156
rect 20212 80116 20252 80156
rect 20294 80116 20334 80156
rect 20376 80116 20416 80156
rect 19948 79780 19988 79820
rect 16300 79696 16340 79736
rect 17260 79696 17300 79736
rect 20140 79696 20180 79736
rect 21388 79696 21428 79736
rect 11404 79612 11444 79652
rect 12748 79612 12788 79652
rect 14188 79612 14228 79652
rect 21004 79612 21044 79652
rect 11212 79528 11252 79568
rect 14572 79528 14612 79568
rect 15820 79528 15860 79568
rect 18508 79528 18548 79568
rect 19372 79528 19412 79568
rect 20428 79528 20468 79568
rect 8524 79444 8564 79484
rect 3688 79360 3728 79400
rect 3770 79360 3810 79400
rect 3852 79360 3892 79400
rect 3934 79360 3974 79400
rect 4016 79360 4056 79400
rect 6412 79360 6452 79400
rect 9292 79360 9332 79400
rect 13324 79360 13364 79400
rect 18808 79360 18848 79400
rect 18890 79360 18930 79400
rect 18972 79360 19012 79400
rect 19054 79360 19094 79400
rect 19136 79360 19176 79400
rect 10636 79276 10676 79316
rect 11212 79276 11252 79316
rect 13036 79276 13076 79316
rect 20140 79276 20180 79316
rect 556 79192 596 79232
rect 2764 79192 2804 79232
rect 3148 79192 3188 79232
rect 12844 79192 12884 79232
rect 15628 79192 15668 79232
rect 19180 79192 19220 79232
rect 19948 79192 19988 79232
rect 1036 79108 1076 79148
rect 172 79024 212 79064
rect 4300 79108 4340 79148
rect 5452 79108 5492 79148
rect 8812 79108 8852 79148
rect 9676 79108 9716 79148
rect 11212 79108 11252 79148
rect 3340 79024 3380 79064
rect 1612 78940 1652 78980
rect 2188 78940 2228 78980
rect 3244 78940 3284 78980
rect 3532 78940 3572 78980
rect 4300 78940 4340 78980
rect 5836 78940 5876 78980
rect 2188 78772 2228 78812
rect 3340 78772 3380 78812
rect 7468 79024 7508 79064
rect 8140 79024 8180 79064
rect 10732 79024 10772 79064
rect 12556 79024 12596 79064
rect 12748 79024 12788 79064
rect 7852 78940 7892 78980
rect 8908 78940 8948 78980
rect 11788 78940 11828 78980
rect 7660 78856 7700 78896
rect 1900 78688 1940 78728
rect 3148 78688 3188 78728
rect 4108 78688 4148 78728
rect 4928 78604 4968 78644
rect 5010 78604 5050 78644
rect 5092 78604 5132 78644
rect 5174 78604 5214 78644
rect 5256 78604 5296 78644
rect 9292 78856 9332 78896
rect 10540 78856 10580 78896
rect 3532 78520 3572 78560
rect 3052 78436 3083 78476
rect 3083 78436 3092 78476
rect 844 78352 884 78392
rect 2092 78268 2132 78308
rect 2380 78268 2420 78308
rect 4012 78268 4052 78308
rect 3436 78184 3476 78224
rect 3724 78184 3764 78224
rect 4108 78184 4148 78224
rect 17164 79108 17204 79148
rect 19660 79108 19700 79148
rect 12940 79024 12980 79064
rect 14476 79024 14516 79064
rect 13228 78940 13257 78980
rect 13257 78940 13268 78980
rect 12172 78772 12212 78812
rect 12748 78772 12788 78812
rect 13228 78772 13259 78812
rect 13259 78772 13268 78812
rect 9484 78688 9524 78728
rect 13036 78688 13076 78728
rect 10636 78604 10676 78644
rect 10540 78520 10580 78560
rect 7180 78436 7220 78476
rect 13804 78856 13844 78896
rect 20812 79024 20852 79064
rect 14764 78940 14804 78980
rect 15148 78940 15188 78980
rect 15628 78940 15668 78980
rect 17740 78940 17780 78980
rect 18220 78940 18260 78980
rect 19084 78940 19124 78980
rect 13900 78772 13940 78812
rect 18988 78772 19028 78812
rect 19564 78772 19604 78812
rect 19180 78520 19220 78560
rect 10348 78436 10388 78476
rect 10924 78436 10964 78476
rect 11980 78436 12020 78476
rect 12940 78436 12980 78476
rect 10252 78352 10292 78392
rect 16492 78436 16532 78476
rect 16972 78436 17012 78476
rect 17932 78436 17972 78476
rect 18028 78352 18068 78392
rect 18796 78352 18836 78392
rect 4396 78268 4436 78308
rect 4588 78268 4628 78308
rect 6700 78268 6740 78308
rect 6892 78268 6932 78308
rect 7468 78268 7508 78308
rect 8428 78268 8468 78308
rect 10060 78268 10100 78308
rect 10348 78268 10388 78308
rect 11884 78268 11924 78308
rect 12364 78268 12404 78308
rect 12556 78268 12596 78308
rect 14380 78268 14420 78308
rect 5260 78184 5300 78224
rect 9964 78184 10004 78224
rect 14092 78184 14132 78224
rect 1324 78016 1364 78056
rect 3148 78016 3188 78056
rect 6412 77932 6452 77972
rect 9100 78100 9140 78140
rect 12364 78100 12404 78140
rect 15628 78184 15668 78224
rect 13612 78100 13652 78140
rect 9868 78016 9908 78056
rect 13324 78016 13364 78056
rect 13900 78016 13940 78056
rect 16492 78268 16532 78308
rect 16108 78184 16148 78224
rect 18892 78268 18932 78308
rect 19180 78268 19220 78308
rect 17164 78184 17204 78224
rect 18796 78184 18836 78224
rect 19564 78184 19604 78224
rect 17932 78100 17972 78140
rect 17164 78016 17204 78056
rect 18988 78016 19028 78056
rect 8524 77932 8564 77972
rect 15724 77932 15764 77972
rect 20044 78856 20084 78896
rect 19948 78772 19988 78812
rect 20048 78604 20088 78644
rect 20130 78604 20170 78644
rect 20212 78604 20252 78644
rect 20294 78604 20334 78644
rect 20376 78604 20416 78644
rect 20044 78352 20084 78392
rect 20140 78268 20180 78308
rect 20044 78100 20084 78140
rect 20140 78016 20180 78056
rect 20908 78016 20948 78056
rect 3688 77848 3728 77888
rect 3770 77848 3810 77888
rect 3852 77848 3892 77888
rect 3934 77848 3974 77888
rect 4016 77848 4056 77888
rect 12844 77848 12884 77888
rect 16492 77848 16532 77888
rect 18808 77848 18848 77888
rect 18890 77848 18930 77888
rect 18972 77848 19012 77888
rect 19054 77848 19094 77888
rect 19136 77848 19176 77888
rect 19276 77848 19316 77888
rect 20908 77848 20948 77888
rect 2284 77680 2324 77720
rect 14476 77764 14516 77804
rect 16108 77764 16148 77804
rect 16684 77764 16724 77804
rect 17164 77764 17204 77804
rect 9100 77680 9140 77720
rect 19852 77680 19892 77720
rect 21292 77680 21332 77720
rect 13516 77596 13556 77636
rect 14476 77596 14516 77636
rect 15724 77596 15764 77636
rect 19372 77596 19412 77636
rect 460 77512 500 77552
rect 7852 77512 7892 77552
rect 9868 77512 9908 77552
rect 12748 77512 12788 77552
rect 15052 77512 15092 77552
rect 15820 77512 15860 77552
rect 17836 77512 17876 77552
rect 1324 77428 1364 77468
rect 2284 77428 2324 77468
rect 3436 77428 3476 77468
rect 3820 77428 3860 77468
rect 4300 77428 4340 77468
rect 7756 77428 7796 77468
rect 8524 77428 8564 77468
rect 10348 77428 10388 77468
rect 10540 77428 10580 77468
rect 12172 77428 12212 77468
rect 15628 77428 15668 77468
rect 16108 77428 16148 77468
rect 16684 77428 16724 77468
rect 17644 77428 17684 77468
rect 18892 77428 18932 77468
rect 3148 77344 3188 77384
rect 1900 77260 1940 77300
rect 4588 77260 4628 77300
rect 5356 77260 5396 77300
rect 21196 77512 21236 77552
rect 19372 77428 19412 77468
rect 19948 77428 19988 77468
rect 9868 77344 9908 77384
rect 11500 77344 11540 77384
rect 12940 77344 12980 77384
rect 16300 77344 16340 77384
rect 19852 77344 19892 77384
rect 7180 77260 7220 77300
rect 8044 77260 8084 77300
rect 10444 77260 10484 77300
rect 12172 77260 12212 77300
rect 17260 77260 17300 77300
rect 2476 77176 2516 77216
rect 6316 77176 6356 77216
rect 12364 77176 12404 77216
rect 15532 77176 15572 77216
rect 2668 77092 2708 77132
rect 4928 77092 4968 77132
rect 5010 77092 5050 77132
rect 5092 77092 5132 77132
rect 5174 77092 5214 77132
rect 5256 77092 5296 77132
rect 10252 77092 10292 77132
rect 10732 77092 10772 77132
rect 14860 77092 14900 77132
rect 4492 77008 4532 77048
rect 4780 76924 4820 76964
rect 5836 76924 5876 76964
rect 6316 76924 6356 76964
rect 8140 76924 8180 76964
rect 10252 76924 10292 76964
rect 1036 76840 1076 76880
rect 1612 76756 1652 76796
rect 2860 76756 2900 76796
rect 3532 76756 3572 76796
rect 1228 76672 1268 76712
rect 2956 76672 2996 76712
rect 4396 76756 4436 76796
rect 4684 76787 4724 76796
rect 4684 76756 4724 76787
rect 5068 76756 5108 76796
rect 5356 76756 5396 76796
rect 8044 76840 8084 76880
rect 8908 76840 8948 76880
rect 9388 76840 9428 76880
rect 6604 76756 6644 76796
rect 7756 76756 7796 76796
rect 4012 76672 4052 76712
rect 6316 76672 6356 76712
rect 8812 76756 8852 76796
rect 9868 76787 9908 76796
rect 9868 76756 9908 76787
rect 10636 76756 10676 76796
rect 8332 76672 8372 76712
rect 9100 76672 9140 76712
rect 9388 76672 9428 76712
rect 3628 76588 3668 76628
rect 4300 76588 4340 76628
rect 4684 76588 4724 76628
rect 8236 76588 8276 76628
rect 9964 76588 10004 76628
rect 10444 76588 10484 76628
rect 10924 76588 10964 76628
rect 14476 77008 14516 77048
rect 14092 76924 14132 76964
rect 15148 76924 15188 76964
rect 20048 77092 20088 77132
rect 20130 77092 20170 77132
rect 20212 77092 20252 77132
rect 20294 77092 20334 77132
rect 20376 77092 20416 77132
rect 15820 76924 15860 76964
rect 18892 76924 18932 76964
rect 18604 76840 18644 76880
rect 12940 76756 12980 76796
rect 13804 76756 13844 76796
rect 14668 76756 14708 76796
rect 16972 76756 17012 76796
rect 18220 76756 18260 76796
rect 19948 76756 19988 76796
rect 20140 76756 20180 76796
rect 14092 76672 14132 76712
rect 15340 76672 15380 76712
rect 2668 76504 2708 76544
rect 4492 76504 4532 76544
rect 6412 76504 6452 76544
rect 6604 76504 6644 76544
rect 17644 76504 17684 76544
rect 10060 76420 10100 76460
rect 10444 76420 10484 76460
rect 15628 76420 15668 76460
rect 20428 76588 20468 76628
rect 21388 76588 21428 76628
rect 18508 76420 18548 76460
rect 19852 76420 19892 76460
rect 3688 76336 3728 76376
rect 3770 76336 3810 76376
rect 3852 76336 3892 76376
rect 3934 76336 3974 76376
rect 4016 76336 4056 76376
rect 12364 76336 12404 76376
rect 18808 76336 18848 76376
rect 18890 76336 18930 76376
rect 18972 76336 19012 76376
rect 19054 76336 19094 76376
rect 19136 76336 19176 76376
rect 14092 76252 14132 76292
rect 14764 76252 14804 76292
rect 17068 76252 17108 76292
rect 18220 76252 18260 76292
rect 8332 76168 8372 76208
rect 9868 76168 9908 76208
rect 12364 76168 12404 76208
rect 7948 76084 7988 76124
rect 8908 76084 8948 76124
rect 10732 76084 10772 76124
rect 12844 76084 12884 76124
rect 1420 76000 1460 76040
rect 2860 76000 2900 76040
rect 3532 76000 3572 76040
rect 4300 76000 4340 76040
rect 5548 76000 5588 76040
rect 5932 76000 5972 76040
rect 7468 76000 7508 76040
rect 1228 75916 1268 75956
rect 2380 75916 2420 75956
rect 3340 75916 3380 75956
rect 3628 75916 3668 75956
rect 4396 75916 4436 75956
rect 5068 75916 5108 75956
rect 5260 75916 5300 75956
rect 6988 75916 7028 75956
rect 7852 75916 7892 75956
rect 15052 76168 15092 76208
rect 18124 76168 18164 76208
rect 15340 76084 15380 76124
rect 10924 76000 10964 76040
rect 13708 76000 13748 76040
rect 9484 75916 9524 75956
rect 6124 75832 6164 75872
rect 6892 75832 6932 75872
rect 11500 75916 11540 75956
rect 12172 75916 12203 75956
rect 12203 75916 12212 75956
rect 13036 75916 13076 75956
rect 13324 75916 13364 75956
rect 13612 75916 13652 75956
rect 14380 75916 14420 75956
rect 19276 76084 19316 76124
rect 17644 76000 17684 76040
rect 18892 76000 18932 76040
rect 20140 76000 20180 76040
rect 17068 75916 17108 75956
rect 17836 75916 17865 75956
rect 17865 75916 17876 75956
rect 18220 75916 18260 75956
rect 12460 75832 12500 75872
rect 12844 75832 12884 75872
rect 16972 75832 17012 75872
rect 2764 75748 2804 75788
rect 5452 75748 5492 75788
rect 6508 75748 6548 75788
rect 6988 75748 7028 75788
rect 7372 75748 7412 75788
rect 13708 75748 13748 75788
rect 13996 75748 14036 75788
rect 15532 75748 15572 75788
rect 17740 75832 17780 75872
rect 18508 75832 18548 75872
rect 17260 75748 17300 75788
rect 17548 75748 17588 75788
rect 19948 75748 19988 75788
rect 20908 75748 20948 75788
rect 940 75664 980 75704
rect 15340 75664 15380 75704
rect 1612 75580 1652 75620
rect 4684 75580 4724 75620
rect 4928 75580 4968 75620
rect 5010 75580 5050 75620
rect 5092 75580 5132 75620
rect 5174 75580 5214 75620
rect 5256 75580 5296 75620
rect 15052 75580 15092 75620
rect 20048 75580 20088 75620
rect 20130 75580 20170 75620
rect 20212 75580 20252 75620
rect 20294 75580 20334 75620
rect 20376 75580 20416 75620
rect 8908 75496 8948 75536
rect 13612 75496 13652 75536
rect 17548 75496 17588 75536
rect 21100 75496 21140 75536
rect 7948 75412 7988 75452
rect 8428 75412 8468 75452
rect 10060 75412 10100 75452
rect 13036 75412 13076 75452
rect 13420 75412 13460 75452
rect 268 75328 308 75368
rect 2476 75328 2516 75368
rect 6412 75328 6452 75368
rect 16588 75412 16628 75452
rect 16204 75328 16244 75368
rect 18796 75328 18836 75368
rect 2284 75244 2324 75284
rect 4876 75244 4916 75284
rect 6124 75244 6164 75284
rect 6988 75244 7028 75284
rect 7756 75244 7796 75284
rect 8620 75244 8660 75284
rect 8908 75244 8948 75284
rect 10252 75244 10292 75284
rect 652 75160 692 75200
rect 1420 75160 1460 75200
rect 2380 75160 2420 75200
rect 4684 75160 4724 75200
rect 8044 75160 8084 75200
rect 9196 75160 9236 75200
rect 844 75076 884 75116
rect 3340 75076 3380 75116
rect 4876 75076 4916 75116
rect 8428 75076 8468 75116
rect 11500 75244 11540 75284
rect 13420 75244 13460 75284
rect 13708 75244 13748 75284
rect 14284 75244 14324 75284
rect 15340 75244 15380 75284
rect 16012 75275 16052 75284
rect 16012 75244 16052 75275
rect 16396 75244 16436 75284
rect 16780 75244 16820 75284
rect 17068 75244 17108 75284
rect 18508 75244 18548 75284
rect 18892 75244 18932 75284
rect 11884 75160 11924 75200
rect 12748 75160 12788 75200
rect 13996 75160 14036 75200
rect 14188 75160 14228 75200
rect 14860 75160 14900 75200
rect 15628 75160 15668 75200
rect 16108 75160 16148 75200
rect 16972 75160 17012 75200
rect 18316 75160 18356 75200
rect 10252 75076 10292 75116
rect 10924 75076 10964 75116
rect 13324 75076 13364 75116
rect 20332 75076 20372 75116
rect 1612 74992 1652 75032
rect 4108 74992 4148 75032
rect 5740 74992 5780 75032
rect 7756 74992 7796 75032
rect 7948 74992 7979 75032
rect 7979 74992 7988 75032
rect 12172 74992 12212 75032
rect 18028 74992 18068 75032
rect 19276 74992 19316 75032
rect 20044 74992 20084 75032
rect 21292 74992 21332 75032
rect 940 74908 980 74948
rect 13804 74908 13844 74948
rect 17068 74908 17108 74948
rect 21100 74908 21140 74948
rect 268 74824 308 74864
rect 3688 74824 3728 74864
rect 3770 74824 3810 74864
rect 3852 74824 3892 74864
rect 3934 74824 3974 74864
rect 4016 74824 4056 74864
rect 12460 74824 12500 74864
rect 18316 74824 18356 74864
rect 18808 74824 18848 74864
rect 18890 74824 18930 74864
rect 18972 74824 19012 74864
rect 19054 74824 19094 74864
rect 19136 74824 19176 74864
rect 4300 74740 4340 74780
rect 8908 74740 8948 74780
rect 556 74656 596 74696
rect 2860 74488 2900 74528
rect 3532 74488 3572 74528
rect 3916 74488 3956 74528
rect 5260 74656 5300 74696
rect 8428 74656 8468 74696
rect 9484 74656 9524 74696
rect 12748 74656 12788 74696
rect 15340 74656 15380 74696
rect 17068 74656 17108 74696
rect 17356 74656 17396 74696
rect 17836 74656 17876 74696
rect 1228 74404 1268 74444
rect 2476 74404 2516 74444
rect 2668 74404 2708 74444
rect 4012 74404 4052 74444
rect 1804 74320 1844 74360
rect 3532 74320 3572 74360
rect 5068 74572 5108 74612
rect 5740 74488 5780 74528
rect 6220 74488 6260 74528
rect 6700 74488 6740 74528
rect 7948 74488 7988 74528
rect 10252 74488 10292 74528
rect 13324 74488 13364 74528
rect 14572 74488 14612 74528
rect 15628 74488 15668 74528
rect 4396 74404 4436 74444
rect 4780 74404 4820 74444
rect 5068 74404 5108 74444
rect 7084 74404 7124 74444
rect 8716 74404 8756 74444
rect 9100 74404 9140 74444
rect 11500 74404 11540 74444
rect 12748 74404 12788 74444
rect 13804 74404 13844 74444
rect 14476 74404 14516 74444
rect 5836 74320 5876 74360
rect 7372 74320 7412 74360
rect 8044 74320 8084 74360
rect 2668 74236 2708 74276
rect 4876 74236 4916 74276
rect 5164 74236 5204 74276
rect 7468 74236 7508 74276
rect 7660 74236 7700 74276
rect 364 73984 404 74024
rect 1996 73900 2036 73940
rect 4396 73900 4436 73940
rect 3244 73816 3284 73856
rect 3532 73816 3572 73856
rect 17260 74488 17300 74528
rect 17644 74488 17684 74528
rect 17836 74488 17876 74528
rect 18028 74488 18068 74528
rect 20332 74488 20372 74528
rect 15340 74404 15380 74444
rect 15532 74404 15572 74444
rect 16396 74404 16436 74444
rect 18412 74404 18452 74444
rect 18892 74404 18932 74444
rect 19948 74404 19988 74444
rect 14572 74320 14612 74360
rect 15628 74320 15668 74360
rect 17932 74320 17972 74360
rect 13036 74236 13076 74276
rect 13804 74236 13844 74276
rect 17740 74236 17780 74276
rect 17068 74152 17108 74192
rect 4928 74068 4968 74108
rect 5010 74068 5050 74108
rect 5092 74068 5132 74108
rect 5174 74068 5214 74108
rect 5256 74068 5296 74108
rect 8236 74068 8276 74108
rect 15820 74068 15860 74108
rect 19084 74236 19124 74276
rect 21292 74236 21332 74276
rect 20048 74068 20088 74108
rect 20130 74068 20170 74108
rect 20212 74068 20252 74108
rect 20294 74068 20334 74108
rect 20376 74068 20416 74108
rect 6988 73984 7028 74024
rect 8140 73984 8180 74024
rect 14668 73984 14708 74024
rect 15628 73984 15668 74024
rect 17836 73984 17876 74024
rect 21196 73984 21236 74024
rect 5548 73900 5588 73940
rect 5356 73816 5396 73856
rect 7084 73816 7124 73856
rect 2284 73732 2324 73772
rect 2476 73732 2516 73772
rect 268 73648 308 73688
rect 4300 73732 4340 73772
rect 4588 73763 4628 73772
rect 4588 73732 4628 73763
rect 5164 73732 5204 73772
rect 6220 73732 6260 73772
rect 7180 73732 7220 73772
rect 7372 73732 7412 73772
rect 7756 73816 7796 73856
rect 4012 73648 4052 73688
rect 7564 73648 7604 73688
rect 8140 73648 8180 73688
rect 4300 73480 4340 73520
rect 11500 73900 11540 73940
rect 11884 73900 11924 73940
rect 15436 73900 15476 73940
rect 16492 73900 16532 73940
rect 17644 73900 17684 73940
rect 19276 73900 19316 73940
rect 11116 73816 11156 73856
rect 13708 73816 13748 73856
rect 17548 73816 17588 73856
rect 18508 73816 18548 73856
rect 18892 73816 18932 73856
rect 10252 73732 10292 73772
rect 11500 73732 11540 73772
rect 13516 73732 13556 73772
rect 13804 73763 13844 73772
rect 13804 73732 13844 73763
rect 14188 73732 14228 73772
rect 14380 73732 14420 73772
rect 15820 73732 15860 73772
rect 16396 73732 16436 73772
rect 12460 73648 12500 73688
rect 12748 73648 12788 73688
rect 13132 73648 13172 73688
rect 13420 73648 13460 73688
rect 14668 73648 14708 73688
rect 15052 73648 15092 73688
rect 10924 73564 10964 73604
rect 8428 73480 8468 73520
rect 18124 73732 18164 73772
rect 18604 73732 18644 73772
rect 15916 73648 15956 73688
rect 12076 73564 12116 73604
rect 19660 73564 19700 73604
rect 20812 73564 20852 73604
rect 8908 73480 8948 73520
rect 9100 73480 9140 73520
rect 15628 73480 15668 73520
rect 16396 73480 16436 73520
rect 17836 73480 17876 73520
rect 19756 73480 19796 73520
rect 3340 73396 3380 73436
rect 364 73312 404 73352
rect 3688 73312 3728 73352
rect 3770 73312 3810 73352
rect 3852 73312 3892 73352
rect 3934 73312 3974 73352
rect 4016 73312 4056 73352
rect 5260 73312 5300 73352
rect 10060 73312 10100 73352
rect 13804 73312 13844 73352
rect 17068 73312 17108 73352
rect 18808 73312 18848 73352
rect 18890 73312 18930 73352
rect 18972 73312 19012 73352
rect 19054 73312 19094 73352
rect 19136 73312 19176 73352
rect 20908 73312 20948 73352
rect 3340 73144 3380 73184
rect 5932 73144 5972 73184
rect 76 72976 116 73016
rect 2572 72892 2612 72932
rect 2956 72892 2996 72932
rect 6796 73228 6836 73268
rect 14188 73228 14228 73268
rect 7084 73144 7124 73184
rect 8140 73144 8180 73184
rect 10828 73144 10868 73184
rect 19276 73144 19307 73184
rect 19307 73144 19316 73184
rect 11020 73060 11060 73100
rect 8140 72976 8180 73016
rect 9100 72976 9140 73016
rect 11500 72976 11540 73016
rect 13324 72976 13364 73016
rect 15244 72976 15284 73016
rect 15628 72976 15668 73016
rect 76 72808 116 72848
rect 4972 72892 5012 72932
rect 5548 72892 5588 72932
rect 6220 72892 6260 72932
rect 6508 72808 6548 72848
rect 8620 72892 8660 72932
rect 8908 72892 8948 72932
rect 10828 72892 10868 72932
rect 11020 72892 11060 72932
rect 11980 72892 12020 72932
rect 12172 72892 12212 72932
rect 13132 72892 13172 72932
rect 13804 72892 13844 72932
rect 15916 72892 15956 72932
rect 18412 72892 18452 72932
rect 11308 72808 11348 72848
rect 3052 72724 3092 72764
rect 3436 72724 3476 72764
rect 4396 72724 4436 72764
rect 6124 72724 6164 72764
rect 9772 72724 9812 72764
rect 14668 72724 14708 72764
rect 748 72640 788 72680
rect 9388 72640 9428 72680
rect 11020 72640 11060 72680
rect 4928 72556 4968 72596
rect 5010 72556 5050 72596
rect 5092 72556 5132 72596
rect 5174 72556 5214 72596
rect 5256 72556 5296 72596
rect 7276 72556 7316 72596
rect 10636 72556 10676 72596
rect 17164 72808 17204 72848
rect 17932 72808 17972 72848
rect 18316 72808 18356 72848
rect 18508 72808 18548 72848
rect 19084 72892 19124 72932
rect 19660 72976 19700 73016
rect 19180 72808 19220 72848
rect 17260 72724 17300 72764
rect 17644 72724 17684 72764
rect 19084 72724 19124 72764
rect 21484 73144 21524 73184
rect 21100 72976 21140 73016
rect 21484 72724 21524 72764
rect 14668 72556 14708 72596
rect 20048 72556 20088 72596
rect 20130 72556 20170 72596
rect 20212 72556 20252 72596
rect 20294 72556 20334 72596
rect 20376 72556 20416 72596
rect 940 72472 980 72512
rect 1708 72472 1748 72512
rect 13132 72472 13172 72512
rect 6796 72388 6836 72428
rect 6988 72388 7028 72428
rect 9196 72388 9236 72428
rect 11500 72388 11540 72428
rect 14668 72388 14708 72428
rect 940 72304 980 72344
rect 3532 72304 3572 72344
rect 5644 72304 5684 72344
rect 1708 72220 1748 72260
rect 2668 72220 2708 72260
rect 2956 72220 2996 72260
rect 3340 72220 3380 72260
rect 4300 72220 4340 72260
rect 6124 72220 6164 72260
rect 6700 72220 6740 72260
rect 7372 72251 7412 72260
rect 7372 72220 7412 72251
rect 7852 72251 7892 72260
rect 7852 72220 7892 72251
rect 8620 72304 8660 72344
rect 11980 72304 12020 72344
rect 9772 72220 9812 72260
rect 10828 72220 10868 72260
rect 12844 72220 12884 72260
rect 14668 72220 14708 72260
rect 18604 72472 18644 72512
rect 21004 72472 21044 72512
rect 17260 72388 17300 72428
rect 17548 72304 17588 72344
rect 20332 72304 20372 72344
rect 14956 72220 14996 72260
rect 15820 72220 15860 72260
rect 16396 72220 16436 72260
rect 17644 72220 17684 72260
rect 18316 72220 18356 72260
rect 18796 72220 18836 72260
rect 19084 72220 19124 72260
rect 268 72136 308 72176
rect 3628 72136 3668 72176
rect 4204 72136 4244 72176
rect 4588 72136 4628 72176
rect 5164 72136 5204 72176
rect 5740 72136 5780 72176
rect 5932 72136 5972 72176
rect 6892 72136 6932 72176
rect 9196 72136 9236 72176
rect 9388 72136 9428 72176
rect 9964 72136 10004 72176
rect 10636 72136 10676 72176
rect 11212 72136 11252 72176
rect 364 72052 404 72092
rect 1708 72052 1748 72092
rect 8620 72052 8660 72092
rect 8908 72052 8948 72092
rect 9100 72052 9140 72092
rect 17164 72052 17204 72092
rect 19948 72251 19988 72260
rect 19948 72220 19988 72251
rect 18124 72136 18164 72176
rect 18892 72052 18932 72092
rect 556 71968 596 72008
rect 2380 71968 2420 72008
rect 6604 71968 6644 72008
rect 13420 71968 13460 72008
rect 14668 71968 14708 72008
rect 14956 71968 14996 72008
rect 16684 71968 16724 72008
rect 19084 71968 19124 72008
rect 21100 71968 21140 72008
rect 2188 71884 2228 71924
rect 9292 71884 9332 71924
rect 18412 71884 18452 71924
rect 3688 71800 3728 71840
rect 3770 71800 3810 71840
rect 3852 71800 3892 71840
rect 3934 71800 3974 71840
rect 4016 71800 4056 71840
rect 12076 71800 12116 71840
rect 15628 71800 15668 71840
rect 18808 71800 18848 71840
rect 18890 71800 18930 71840
rect 18972 71800 19012 71840
rect 19054 71800 19094 71840
rect 19136 71800 19176 71840
rect 1228 71632 1268 71672
rect 7660 71632 7700 71672
rect 7852 71632 7892 71672
rect 15532 71632 15572 71672
rect 12172 71548 12212 71588
rect 14572 71548 14612 71588
rect 15436 71548 15476 71588
rect 16396 71548 16436 71588
rect 1708 71464 1748 71504
rect 2476 71464 2516 71504
rect 2860 71464 2900 71504
rect 3340 71464 3380 71504
rect 4588 71464 4628 71504
rect 5260 71464 5300 71504
rect 10348 71464 10388 71504
rect 2764 71380 2804 71420
rect 3820 71380 3860 71420
rect 4108 71380 4148 71420
rect 5548 71380 5588 71420
rect 2284 71296 2324 71336
rect 3724 71296 3764 71336
rect 5932 71296 5972 71336
rect 556 71212 596 71252
rect 5740 71212 5780 71252
rect 15532 71464 15572 71504
rect 17260 71464 17300 71504
rect 18508 71464 18548 71504
rect 19948 71464 19988 71504
rect 20332 71464 20372 71504
rect 6604 71380 6644 71420
rect 8044 71380 8084 71420
rect 8716 71380 8756 71420
rect 10252 71380 10292 71420
rect 10636 71380 10676 71420
rect 11500 71380 11540 71420
rect 12076 71380 12116 71420
rect 12844 71380 12884 71420
rect 13036 71380 13076 71420
rect 13420 71380 13460 71420
rect 15340 71380 15380 71420
rect 15820 71380 15860 71420
rect 16108 71380 16148 71420
rect 16684 71380 16724 71420
rect 17836 71380 17876 71420
rect 18412 71380 18452 71420
rect 19756 71380 19796 71420
rect 6220 71296 6260 71336
rect 13324 71296 13364 71336
rect 12844 71212 12884 71252
rect 13420 71212 13460 71252
rect 14572 71212 14612 71252
rect 2572 71044 2612 71084
rect 7660 71128 7700 71168
rect 13804 71128 13844 71168
rect 15532 71296 15572 71336
rect 18124 71296 18164 71336
rect 18988 71212 19028 71252
rect 4928 71044 4968 71084
rect 5010 71044 5050 71084
rect 5092 71044 5132 71084
rect 5174 71044 5214 71084
rect 5256 71044 5296 71084
rect 6028 71044 6068 71084
rect 1228 70960 1268 71000
rect 2092 70960 2132 71000
rect 13036 70960 13076 71000
rect 1132 70876 1172 70916
rect 7468 70876 7508 70916
rect 11980 70876 12020 70916
rect 748 70708 788 70748
rect 2764 70708 2804 70748
rect 3436 70708 3476 70748
rect 1420 70624 1460 70664
rect 2668 70624 2708 70664
rect 20044 71212 20084 71252
rect 21100 71212 21140 71252
rect 19756 71128 19796 71168
rect 20048 71044 20088 71084
rect 20130 71044 20170 71084
rect 20212 71044 20252 71084
rect 20294 71044 20334 71084
rect 20376 71044 20416 71084
rect 19276 70960 19316 71000
rect 17548 70876 17588 70916
rect 20332 70876 20372 70916
rect 4396 70792 4436 70832
rect 6796 70792 6836 70832
rect 7180 70792 7220 70832
rect 4876 70708 4916 70748
rect 12076 70792 12116 70832
rect 12460 70792 12500 70832
rect 18988 70792 19028 70832
rect 20428 70792 20468 70832
rect 4300 70624 4340 70664
rect 748 70540 788 70580
rect 4108 70540 4148 70580
rect 1420 70456 1460 70496
rect 4300 70456 4340 70496
rect 6028 70708 6068 70748
rect 7372 70708 7412 70748
rect 9292 70708 9332 70748
rect 9772 70708 9812 70748
rect 10348 70708 10388 70748
rect 7276 70624 7316 70664
rect 12172 70708 12212 70748
rect 13132 70708 13172 70748
rect 13612 70708 13652 70748
rect 14572 70708 14612 70748
rect 15724 70708 15764 70748
rect 17068 70708 17108 70748
rect 17260 70708 17300 70748
rect 17932 70708 17972 70748
rect 18220 70708 18260 70748
rect 19276 70708 19316 70748
rect 11212 70624 11252 70664
rect 12844 70624 12884 70664
rect 18028 70624 18068 70664
rect 18604 70624 18644 70664
rect 6604 70540 6644 70580
rect 13036 70540 13076 70580
rect 18508 70540 18548 70580
rect 19852 70540 19892 70580
rect 5740 70456 5780 70496
rect 6028 70456 6068 70496
rect 7180 70456 7220 70496
rect 13228 70456 13268 70496
rect 17548 70456 17588 70496
rect 17836 70456 17876 70496
rect 4876 70372 4916 70412
rect 9004 70372 9044 70412
rect 11500 70372 11540 70412
rect 14764 70372 14804 70412
rect 15436 70372 15476 70412
rect 17356 70372 17396 70412
rect 172 70288 212 70328
rect 3688 70288 3728 70328
rect 3770 70288 3810 70328
rect 3852 70288 3892 70328
rect 3934 70288 3974 70328
rect 4016 70288 4056 70328
rect 16396 70288 16436 70328
rect 18808 70288 18848 70328
rect 18890 70288 18930 70328
rect 18972 70288 19012 70328
rect 19054 70288 19094 70328
rect 19136 70288 19176 70328
rect 19660 70288 19700 70328
rect 9196 70204 9236 70244
rect 16108 70204 16148 70244
rect 17164 70204 17204 70244
rect 8140 70120 8180 70160
rect 16012 70120 16052 70160
rect 17452 70120 17492 70160
rect 18796 70120 18836 70160
rect 19756 70120 19796 70160
rect 4492 70036 4532 70076
rect 4684 70036 4724 70076
rect 7564 70036 7604 70076
rect 13708 70036 13748 70076
rect 19660 70036 19700 70076
rect 1708 69868 1748 69908
rect 2572 69868 2612 69908
rect 2860 69868 2900 69908
rect 4972 69868 5012 69908
rect 6892 69868 6932 69908
rect 7180 69868 7211 69908
rect 7211 69868 7220 69908
rect 7372 69868 7412 69908
rect 8236 69952 8276 69992
rect 8716 69952 8756 69992
rect 10348 69952 10388 69992
rect 10828 69952 10868 69992
rect 12076 69952 12116 69992
rect 12652 69952 12692 69992
rect 14572 69952 14612 69992
rect 17164 69952 17204 69992
rect 17932 69952 17972 69992
rect 18316 69952 18356 69992
rect 19756 69952 19796 69992
rect 20140 69952 20180 69992
rect 8620 69868 8660 69908
rect 9772 69868 9812 69908
rect 10540 69868 10580 69908
rect 11308 69868 11348 69908
rect 12748 69868 12788 69908
rect 14092 69868 14132 69908
rect 16012 69868 16052 69908
rect 1324 69616 1364 69656
rect 460 69280 500 69320
rect 4012 69784 4052 69824
rect 4876 69784 4916 69824
rect 6124 69784 6164 69824
rect 8140 69784 8180 69824
rect 12556 69784 12596 69824
rect 2956 69700 2996 69740
rect 4588 69700 4628 69740
rect 7180 69700 7220 69740
rect 8236 69700 8276 69740
rect 11308 69700 11348 69740
rect 2092 69616 2132 69656
rect 4928 69532 4968 69572
rect 5010 69532 5050 69572
rect 5092 69532 5132 69572
rect 5174 69532 5214 69572
rect 5256 69532 5296 69572
rect 5740 69532 5780 69572
rect 1708 69364 1748 69404
rect 7372 69448 7412 69488
rect 7564 69364 7595 69404
rect 7595 69364 7604 69404
rect 13516 69700 13556 69740
rect 15532 69700 15572 69740
rect 8044 69364 8084 69404
rect 6988 69280 7028 69320
rect 1228 68944 1268 68984
rect 76 68608 116 68648
rect 1324 68356 1364 68396
rect 1036 68272 1076 68312
rect 2764 69196 2804 69236
rect 3052 69196 3092 69236
rect 3628 69196 3668 69236
rect 4012 69196 4052 69236
rect 2860 69112 2900 69152
rect 4300 69196 4340 69236
rect 5260 69196 5300 69236
rect 6892 69196 6932 69236
rect 7372 69196 7412 69236
rect 8236 69280 8276 69320
rect 8044 69196 8073 69236
rect 8073 69196 8084 69236
rect 11020 69280 11060 69320
rect 17548 69868 17588 69908
rect 18412 69868 18452 69908
rect 18796 69868 18836 69908
rect 19276 69868 19316 69908
rect 21196 69868 21236 69908
rect 18124 69784 18164 69824
rect 21004 69784 21044 69824
rect 18892 69700 18932 69740
rect 19756 69700 19796 69740
rect 20044 69700 20084 69740
rect 21196 69700 21236 69740
rect 19084 69616 19124 69656
rect 14764 69448 14804 69488
rect 15052 69448 15092 69488
rect 20048 69532 20088 69572
rect 20130 69532 20170 69572
rect 20212 69532 20252 69572
rect 20294 69532 20334 69572
rect 20376 69532 20416 69572
rect 17932 69448 17972 69488
rect 21388 69448 21428 69488
rect 18412 69280 18452 69320
rect 18796 69280 18836 69320
rect 20236 69280 20276 69320
rect 5548 69112 5588 69152
rect 11500 69196 11540 69236
rect 11788 69196 11828 69236
rect 14572 69196 14612 69236
rect 10252 69112 10292 69152
rect 10540 69112 10580 69152
rect 13324 69112 13364 69152
rect 13804 69112 13844 69152
rect 15244 69196 15284 69236
rect 15532 69196 15572 69236
rect 14764 69112 14804 69152
rect 3052 69028 3092 69068
rect 3340 69028 3380 69068
rect 7276 69028 7316 69068
rect 8236 69028 8276 69068
rect 9772 69028 9812 69068
rect 10348 69028 10388 69068
rect 13228 69028 13268 69068
rect 2860 68944 2900 68984
rect 6700 68944 6740 68984
rect 7564 68944 7604 68984
rect 9868 68944 9908 68984
rect 12460 68944 12500 68984
rect 3688 68776 3728 68816
rect 3770 68776 3810 68816
rect 3852 68776 3892 68816
rect 3934 68776 3974 68816
rect 4016 68776 4056 68816
rect 7372 68776 7412 68816
rect 16972 69196 17012 69236
rect 17836 69227 17876 69236
rect 17836 69196 17876 69227
rect 19852 69227 19892 69236
rect 19852 69196 19892 69227
rect 16012 69112 16052 69152
rect 16588 69112 16628 69152
rect 18124 69112 18164 69152
rect 18892 69112 18932 69152
rect 18412 69028 18452 69068
rect 14956 68944 14996 68984
rect 20812 68944 20852 68984
rect 13804 68860 13844 68900
rect 17548 68860 17588 68900
rect 14572 68776 14612 68816
rect 18808 68776 18848 68816
rect 18890 68776 18930 68816
rect 18972 68776 19012 68816
rect 19054 68776 19094 68816
rect 19136 68776 19176 68816
rect 10924 68692 10964 68732
rect 12460 68692 12500 68732
rect 2188 68608 2228 68648
rect 2476 68608 2516 68648
rect 1804 68272 1844 68312
rect 1612 68188 1652 68228
rect 4972 68608 5012 68648
rect 6220 68608 6260 68648
rect 10060 68608 10100 68648
rect 15244 68608 15284 68648
rect 16492 68608 16532 68648
rect 19276 68608 19316 68648
rect 7468 68524 7508 68564
rect 8716 68524 8756 68564
rect 12652 68524 12692 68564
rect 12940 68524 12980 68564
rect 4012 68440 4052 68480
rect 6124 68440 6164 68480
rect 7180 68440 7220 68480
rect 7564 68440 7604 68480
rect 8236 68440 8276 68480
rect 9484 68440 9524 68480
rect 20908 68524 20948 68564
rect 1996 68356 2036 68396
rect 2956 68356 2996 68396
rect 3916 68356 3956 68396
rect 5932 68356 5972 68396
rect 7372 68356 7412 68396
rect 9868 68356 9908 68396
rect 11788 68356 11828 68396
rect 12460 68356 12500 68396
rect 13228 68356 13268 68396
rect 2572 68188 2612 68228
rect 4300 68272 4340 68312
rect 7468 68272 7508 68312
rect 10252 68272 10292 68312
rect 12940 68272 12980 68312
rect 4972 68188 5012 68228
rect 5548 68188 5588 68228
rect 7180 68188 7220 68228
rect 8236 68188 8276 68228
rect 15532 68440 15572 68480
rect 19852 68440 19892 68480
rect 13804 68356 13812 68396
rect 13812 68356 13844 68396
rect 14380 68356 14420 68396
rect 15820 68356 15860 68396
rect 16204 68356 16244 68396
rect 17548 68356 17588 68396
rect 18796 68356 18836 68396
rect 13996 68272 14036 68312
rect 14572 68272 14612 68312
rect 16108 68272 16148 68312
rect 4204 68104 4244 68144
rect 10060 68104 10100 68144
rect 10252 68104 10292 68144
rect 16588 68188 16628 68228
rect 17260 68188 17300 68228
rect 20236 68188 20276 68228
rect 21388 68188 21428 68228
rect 14860 68104 14900 68144
rect 16492 68104 16532 68144
rect 1324 68020 1364 68060
rect 4928 68020 4968 68060
rect 5010 68020 5050 68060
rect 5092 68020 5132 68060
rect 5174 68020 5214 68060
rect 5256 68020 5296 68060
rect 7564 68020 7604 68060
rect 13996 68020 14036 68060
rect 844 67936 884 67976
rect 7084 67936 7124 67976
rect 10636 67936 10676 67976
rect 11116 67936 11156 67976
rect 11884 67936 11924 67976
rect 10540 67852 10580 67892
rect 12748 67852 12788 67892
rect 13036 67852 13076 67892
rect 15532 67852 15572 67892
rect 16204 67852 16244 67892
rect 3916 67768 3956 67808
rect 7180 67768 7220 67808
rect 9484 67768 9524 67808
rect 844 67684 884 67724
rect 2476 67684 2516 67724
rect 2668 67684 2708 67724
rect 2860 67684 2900 67724
rect 4108 67715 4148 67724
rect 4108 67684 4148 67715
rect 4588 67715 4628 67724
rect 4588 67684 4628 67715
rect 5740 67684 5780 67724
rect 6892 67715 6932 67724
rect 6892 67684 6932 67715
rect 8236 67684 8276 67724
rect 8428 67684 8468 67724
rect 9292 67684 9332 67724
rect 10348 67684 10388 67724
rect 1420 67600 1460 67640
rect 3340 67600 3380 67640
rect 4780 67600 4820 67640
rect 9004 67600 9044 67640
rect 9676 67600 9716 67640
rect 15436 67768 15476 67808
rect 11116 67684 11156 67724
rect 12172 67684 12212 67724
rect 20048 68020 20088 68060
rect 20130 68020 20170 68060
rect 20212 68020 20252 68060
rect 20294 68020 20334 68060
rect 20376 68020 20416 68060
rect 12748 67684 12788 67724
rect 4300 67516 4340 67556
rect 4876 67516 4916 67556
rect 8044 67516 8084 67556
rect 14092 67684 14132 67724
rect 15244 67684 15284 67724
rect 16588 67684 16628 67724
rect 20140 67684 20180 67724
rect 14860 67600 14900 67640
rect 16492 67600 16532 67640
rect 17260 67600 17300 67640
rect 13996 67516 14036 67556
rect 14380 67516 14420 67556
rect 15820 67516 15860 67556
rect 18796 67516 18836 67556
rect 2476 67432 2516 67472
rect 14668 67432 14708 67472
rect 15436 67432 15476 67472
rect 21292 67432 21332 67472
rect 652 67264 692 67304
rect 2092 67264 2132 67304
rect 3688 67264 3728 67304
rect 3770 67264 3810 67304
rect 3852 67264 3892 67304
rect 3934 67264 3974 67304
rect 4016 67264 4056 67304
rect 5836 67096 5876 67136
rect 4396 67012 4436 67052
rect 4972 67012 5012 67052
rect 1420 66928 1460 66968
rect 4108 66928 4148 66968
rect 8620 67012 8660 67052
rect 7660 66928 7700 66968
rect 8908 67096 8948 67136
rect 1996 66844 2036 66884
rect 2956 66844 2996 66884
rect 4204 66844 4244 66884
rect 4876 66844 4916 66884
rect 5836 66844 5876 66884
rect 6220 66844 6260 66884
rect 8140 66844 8180 66884
rect 7372 66760 7412 66800
rect 9484 66844 9524 66884
rect 10156 66844 10196 66884
rect 11500 66928 11540 66968
rect 11404 66844 11444 66884
rect 11692 66844 11732 66884
rect 13132 67096 13172 67136
rect 18028 67096 18068 67136
rect 12844 67012 12884 67052
rect 17164 67012 17204 67052
rect 18808 67264 18848 67304
rect 18890 67264 18930 67304
rect 18972 67264 19012 67304
rect 19054 67264 19094 67304
rect 19136 67264 19176 67304
rect 13996 66928 14036 66968
rect 15244 66928 15284 66968
rect 15820 66928 15860 66968
rect 20812 67012 20852 67052
rect 20716 66928 20756 66968
rect 13516 66844 13556 66884
rect 14092 66844 14132 66884
rect 14860 66844 14900 66884
rect 16300 66844 16340 66884
rect 16588 66844 16628 66884
rect 17740 66844 17780 66884
rect 18412 66844 18452 66884
rect 18796 66844 18836 66884
rect 7660 66760 7700 66800
rect 12748 66760 12788 66800
rect 18124 66760 18164 66800
rect 18316 66760 18356 66800
rect 652 66676 692 66716
rect 2668 66676 2708 66716
rect 4204 66676 4244 66716
rect 8332 66676 8372 66716
rect 11116 66676 11156 66716
rect 13036 66676 13076 66716
rect 15052 66676 15092 66716
rect 16108 66676 16148 66716
rect 17356 66676 17396 66716
rect 17836 66676 17876 66716
rect 19756 66676 19796 66716
rect 20428 66676 20468 66716
rect 940 66592 980 66632
rect 11884 66592 11924 66632
rect 13516 66592 13556 66632
rect 16492 66592 16532 66632
rect 4928 66508 4968 66548
rect 5010 66508 5050 66548
rect 5092 66508 5132 66548
rect 5174 66508 5214 66548
rect 5256 66508 5296 66548
rect 6412 66508 6452 66548
rect 20048 66508 20088 66548
rect 20130 66508 20170 66548
rect 20212 66508 20252 66548
rect 20294 66508 20334 66548
rect 20376 66508 20416 66548
rect 4780 66340 4820 66380
rect 6988 66340 7028 66380
rect 7276 66340 7316 66380
rect 1228 66256 1268 66296
rect 2860 66256 2900 66296
rect 4492 66256 4532 66296
rect 5356 66256 5396 66296
rect 1420 66172 1460 66212
rect 1612 66172 1652 66212
rect 2572 66172 2612 66212
rect 3628 66172 3668 66212
rect 3820 66172 3860 66212
rect 4204 66203 4244 66212
rect 4204 66172 4244 66203
rect 6220 66172 6260 66212
rect 13804 66340 13844 66380
rect 21292 66340 21332 66380
rect 12652 66256 12692 66296
rect 14668 66256 14708 66296
rect 18028 66256 18068 66296
rect 7948 66172 7988 66212
rect 9484 66172 9524 66212
rect 11788 66172 11828 66212
rect 12076 66172 12116 66212
rect 12460 66172 12500 66212
rect 14380 66172 14420 66212
rect 15340 66172 15380 66212
rect 15628 66172 15668 66212
rect 1804 66088 1844 66128
rect 1996 66088 2036 66128
rect 6604 66088 6643 66128
rect 6643 66088 6644 66128
rect 6892 66088 6932 66128
rect 11212 66088 11252 66128
rect 13036 66088 13076 66128
rect 13228 66088 13268 66128
rect 13516 66088 13556 66128
rect 16396 66203 16436 66212
rect 16396 66172 16436 66203
rect 17836 66172 17876 66212
rect 18316 66172 18356 66212
rect 19276 66203 19316 66212
rect 19276 66172 19316 66203
rect 14764 66088 14804 66128
rect 15724 66088 15764 66128
rect 17740 66088 17780 66128
rect 19180 66088 19220 66128
rect 2860 66004 2900 66044
rect 7180 66004 7220 66044
rect 15820 66004 15860 66044
rect 16780 66004 16820 66044
rect 460 65920 500 65960
rect 940 65920 980 65960
rect 1612 65920 1652 65960
rect 1996 65920 2036 65960
rect 5356 65920 5396 65960
rect 5836 65920 5876 65960
rect 9484 65920 9524 65960
rect 9964 65920 10004 65960
rect 10636 65920 10676 65960
rect 11020 65920 11060 65960
rect 11500 65920 11540 65960
rect 16492 65920 16532 65960
rect 1228 65836 1268 65876
rect 11212 65836 11252 65876
rect 13804 65836 13844 65876
rect 3688 65752 3728 65792
rect 3770 65752 3810 65792
rect 3852 65752 3892 65792
rect 3934 65752 3974 65792
rect 4016 65752 4056 65792
rect 5356 65752 5396 65792
rect 1804 65668 1844 65708
rect 8812 65668 8852 65708
rect 268 65584 308 65624
rect 1420 65584 1460 65624
rect 2956 65584 2996 65624
rect 4012 65584 4052 65624
rect 5932 65584 5972 65624
rect 6220 65584 6260 65624
rect 7948 65500 7988 65540
rect 9292 65500 9332 65540
rect 2860 65416 2900 65456
rect 3532 65416 3572 65456
rect 4300 65416 4340 65456
rect 1420 65332 1460 65372
rect 2956 65332 2996 65372
rect 5164 65332 5204 65372
rect 364 65248 404 65288
rect 1036 65248 1076 65288
rect 2956 65164 2996 65204
rect 3532 65164 3572 65204
rect 4012 65080 4052 65120
rect 9484 65416 9524 65456
rect 18604 66004 18644 66044
rect 20044 65920 20084 65960
rect 18808 65752 18848 65792
rect 18890 65752 18930 65792
rect 18972 65752 19012 65792
rect 19054 65752 19094 65792
rect 19136 65752 19176 65792
rect 21484 65920 21524 65960
rect 12652 65584 12692 65624
rect 15340 65584 15380 65624
rect 11692 65416 11732 65456
rect 12844 65416 12884 65456
rect 13132 65416 13172 65456
rect 16396 65500 16436 65540
rect 18508 65500 18548 65540
rect 13516 65416 13556 65456
rect 15628 65416 15668 65456
rect 10060 65332 10100 65372
rect 10252 65332 10292 65372
rect 10540 65332 10580 65372
rect 11020 65332 11028 65372
rect 11028 65332 11060 65372
rect 12748 65332 12788 65372
rect 13420 65332 13460 65372
rect 14092 65332 14132 65372
rect 15052 65332 15092 65372
rect 6700 65248 6740 65288
rect 7756 65248 7796 65288
rect 10156 65248 10196 65288
rect 5932 65164 5972 65204
rect 15724 65332 15764 65372
rect 16300 65332 16340 65372
rect 16684 65332 16692 65372
rect 16692 65332 16724 65372
rect 17356 65332 17396 65372
rect 18508 65332 18548 65372
rect 19084 65332 19124 65372
rect 13516 65248 13556 65288
rect 14668 65248 14708 65288
rect 16876 65248 16916 65288
rect 17644 65248 17684 65288
rect 19180 65248 19220 65288
rect 8524 65164 8564 65204
rect 9484 65164 9524 65204
rect 9964 65164 10004 65204
rect 11212 65164 11252 65204
rect 11980 65164 12020 65204
rect 14572 65164 14612 65204
rect 17740 65164 17780 65204
rect 20140 65164 20180 65204
rect 21388 65164 21428 65204
rect 11692 65080 11732 65120
rect 4928 64996 4968 65036
rect 5010 64996 5050 65036
rect 5092 64996 5132 65036
rect 5174 64996 5214 65036
rect 5256 64996 5296 65036
rect 8620 64996 8660 65036
rect 8812 64996 8852 65036
rect 12940 64996 12980 65036
rect 20048 64996 20088 65036
rect 20130 64996 20170 65036
rect 20212 64996 20252 65036
rect 20294 64996 20334 65036
rect 20376 64996 20416 65036
rect 556 64912 596 64952
rect 10156 64912 10196 64952
rect 11212 64912 11252 64952
rect 21100 64912 21140 64952
rect 4300 64828 4340 64868
rect 9292 64828 9332 64868
rect 9676 64828 9716 64868
rect 10252 64828 10292 64868
rect 14092 64828 14132 64868
rect 16684 64828 16724 64868
rect 19180 64828 19220 64868
rect 20428 64828 20468 64868
rect 4492 64744 4532 64784
rect 2668 64660 2708 64700
rect 3052 64660 3092 64700
rect 3340 64660 3380 64700
rect 3820 64660 3860 64700
rect 4684 64660 4724 64700
rect 1228 64576 1268 64616
rect 1708 64576 1748 64616
rect 3628 64576 3668 64616
rect 5836 64691 5876 64700
rect 5836 64660 5876 64691
rect 7180 64660 7220 64700
rect 7756 64660 7796 64700
rect 8140 64691 8180 64700
rect 8140 64660 8180 64691
rect 10156 64744 10196 64784
rect 12076 64744 12116 64784
rect 12652 64744 12692 64784
rect 21100 64744 21140 64784
rect 8524 64660 8555 64700
rect 8555 64660 8564 64700
rect 8812 64660 8852 64700
rect 9292 64660 9332 64700
rect 9484 64660 9524 64700
rect 10540 64660 10580 64700
rect 11116 64691 11156 64700
rect 11116 64660 11156 64691
rect 13804 64660 13844 64700
rect 15724 64660 15764 64700
rect 4876 64576 4916 64616
rect 9004 64576 9044 64616
rect 10060 64576 10100 64616
rect 11020 64576 11060 64616
rect 12076 64576 12116 64616
rect 12460 64576 12500 64616
rect 12748 64576 12788 64616
rect 2476 64492 2516 64532
rect 4300 64492 4340 64532
rect 6124 64492 6164 64532
rect 8620 64492 8660 64532
rect 556 64408 596 64448
rect 1804 64408 1844 64448
rect 3052 64408 3092 64448
rect 4012 64408 4052 64448
rect 8812 64408 8852 64448
rect 16780 64660 16820 64700
rect 16972 64660 17012 64700
rect 18220 64660 18260 64700
rect 16396 64576 16436 64616
rect 17260 64576 17300 64616
rect 20140 64576 20180 64616
rect 20908 64576 20948 64616
rect 11116 64408 11156 64448
rect 12460 64408 12500 64448
rect 18028 64408 18068 64448
rect 1420 64324 1460 64364
rect 4300 64324 4340 64364
rect 7948 64324 7988 64364
rect 1132 64240 1172 64280
rect 3688 64240 3728 64280
rect 3770 64240 3810 64280
rect 3852 64240 3892 64280
rect 3934 64240 3974 64280
rect 4016 64240 4056 64280
rect 5068 64240 5108 64280
rect 5836 64240 5876 64280
rect 7756 64240 7796 64280
rect 9868 64240 9908 64280
rect 12556 64240 12596 64280
rect 12940 64240 12980 64280
rect 15436 64240 15476 64280
rect 18808 64240 18848 64280
rect 18890 64240 18930 64280
rect 18972 64240 19012 64280
rect 19054 64240 19094 64280
rect 19136 64240 19176 64280
rect 6124 64156 6164 64196
rect 11308 64156 11348 64196
rect 4780 64072 4820 64112
rect 9196 64072 9236 64112
rect 16684 64072 16724 64112
rect 3340 63988 3380 64028
rect 6220 63988 6260 64028
rect 8620 63988 8660 64028
rect 11692 63988 11732 64028
rect 12076 63988 12116 64028
rect 748 63904 788 63944
rect 5068 63904 5108 63944
rect 6700 63904 6740 63944
rect 7756 63904 7796 63944
rect 8140 63904 8180 63944
rect 8428 63904 8468 63944
rect 9004 63904 9044 63944
rect 9676 63904 9716 63944
rect 12268 63904 12308 63944
rect 1420 63820 1460 63860
rect 2860 63820 2900 63860
rect 3916 63820 3956 63860
rect 4300 63820 4340 63860
rect 6220 63820 6260 63860
rect 7276 63820 7316 63860
rect 15052 63988 15092 64028
rect 15916 63988 15956 64028
rect 12652 63904 12692 63944
rect 15436 63904 15476 63944
rect 15724 63904 15764 63944
rect 8524 63820 8555 63860
rect 8555 63820 8564 63860
rect 9292 63820 9332 63860
rect 9484 63820 9524 63860
rect 10732 63820 10772 63860
rect 11500 63820 11540 63860
rect 11980 63820 12020 63860
rect 13132 63820 13172 63860
rect 13996 63820 14036 63860
rect 19276 63988 19316 64028
rect 17356 63904 17396 63944
rect 18508 63904 18548 63944
rect 20908 64408 20948 64448
rect 19564 63904 19604 63944
rect 20044 64072 20084 64112
rect 15916 63820 15956 63860
rect 16396 63820 16436 63860
rect 17260 63820 17300 63860
rect 18220 63820 18260 63860
rect 18796 63820 18836 63860
rect 18988 63820 19028 63860
rect 19180 63820 19220 63860
rect 20812 63988 20852 64028
rect 21100 63904 21140 63944
rect 4204 63736 4244 63776
rect 5740 63736 5780 63776
rect 9196 63736 9236 63776
rect 11788 63736 11828 63776
rect 13228 63736 13268 63776
rect 14092 63736 14132 63776
rect 1708 63652 1748 63692
rect 2092 63652 2132 63692
rect 5356 63652 5396 63692
rect 6124 63652 6164 63692
rect 7756 63652 7796 63692
rect 9004 63652 9044 63692
rect 10060 63652 10100 63692
rect 12076 63652 12116 63692
rect 14380 63652 14420 63692
rect 15244 63652 15284 63692
rect 19852 63652 19892 63692
rect 1324 63568 1364 63608
rect 7948 63568 7988 63608
rect 1708 63484 1748 63524
rect 4928 63484 4968 63524
rect 5010 63484 5050 63524
rect 5092 63484 5132 63524
rect 5174 63484 5214 63524
rect 5256 63484 5296 63524
rect 4492 63400 4532 63440
rect 11308 63568 11348 63608
rect 12652 63568 12692 63608
rect 20428 63652 20468 63692
rect 16684 63568 16724 63608
rect 18604 63568 18644 63608
rect 8620 63484 8660 63524
rect 8908 63484 8948 63524
rect 9388 63484 9428 63524
rect 11116 63484 11156 63524
rect 13612 63484 13652 63524
rect 15052 63484 15092 63524
rect 16300 63484 16340 63524
rect 17260 63484 17300 63524
rect 20048 63484 20088 63524
rect 20130 63484 20170 63524
rect 20212 63484 20252 63524
rect 20294 63484 20334 63524
rect 20376 63484 20416 63524
rect 9964 63400 10004 63440
rect 12940 63400 12980 63440
rect 13900 63400 13940 63440
rect 6700 63316 6740 63356
rect 9196 63316 9227 63356
rect 9227 63316 9236 63356
rect 9676 63316 9716 63356
rect 12556 63316 12596 63356
rect 14668 63316 14708 63356
rect 15724 63316 15764 63356
rect 15916 63316 15956 63356
rect 21196 63400 21236 63440
rect 20236 63316 20276 63356
rect 1228 63232 1268 63272
rect 8812 63232 8852 63272
rect 1420 63148 1460 63188
rect 2668 63148 2708 63188
rect 3916 63148 3956 63188
rect 4780 63148 4820 63188
rect 6604 63148 6644 63188
rect 7756 63148 7796 63188
rect 8044 63148 8084 63188
rect 1516 63064 1556 63104
rect 7564 63064 7604 63104
rect 8140 63064 8180 63104
rect 1900 62980 1940 63020
rect 4012 62980 4052 63020
rect 4972 62980 5012 63020
rect 5452 62980 5492 63020
rect 6700 62980 6740 63020
rect 9388 63148 9428 63188
rect 9676 63148 9716 63188
rect 10348 63148 10388 63188
rect 10828 63148 10868 63188
rect 11500 63148 11540 63188
rect 11692 63148 11732 63188
rect 12748 63148 12788 63188
rect 13612 63148 13652 63188
rect 9004 63064 9035 63104
rect 9035 63064 9044 63104
rect 12172 63064 12212 63104
rect 14380 63148 14420 63188
rect 14956 63148 14996 63188
rect 16972 63148 17012 63188
rect 18028 63148 18068 63188
rect 18220 63148 18258 63188
rect 18258 63148 18260 63188
rect 18508 63148 18548 63188
rect 19180 63179 19220 63188
rect 19180 63148 19220 63179
rect 14092 63064 14132 63104
rect 15052 63064 15092 63104
rect 17836 63064 17876 63104
rect 18796 63064 18836 63104
rect 19468 63064 19508 63104
rect 8524 62980 8564 63020
rect 9388 62980 9428 63020
rect 460 62896 500 62936
rect 3148 62896 3188 62936
rect 5740 62896 5780 62936
rect 11020 62896 11060 62936
rect 11692 62896 11732 62936
rect 14380 62896 14420 62936
rect 15436 62896 15476 62936
rect 15052 62812 15092 62852
rect 16012 62896 16052 62936
rect 18028 62896 18068 62936
rect 18988 62980 19028 63020
rect 15820 62812 15860 62852
rect 20812 62896 20852 62936
rect 1516 62728 1556 62768
rect 3688 62728 3728 62768
rect 3770 62728 3810 62768
rect 3852 62728 3892 62768
rect 3934 62728 3974 62768
rect 4016 62728 4056 62768
rect 4876 62728 4916 62768
rect 6604 62728 6644 62768
rect 10636 62728 10676 62768
rect 18808 62728 18848 62768
rect 18890 62728 18930 62768
rect 18972 62728 19012 62768
rect 19054 62728 19094 62768
rect 19136 62728 19176 62768
rect 2860 62644 2900 62684
rect 7756 62644 7796 62684
rect 13132 62644 13172 62684
rect 13420 62644 13460 62684
rect 17260 62644 17300 62684
rect 5740 62560 5780 62600
rect 6700 62560 6740 62600
rect 7084 62560 7124 62600
rect 8908 62560 8948 62600
rect 9388 62560 9428 62600
rect 9676 62560 9716 62600
rect 10444 62560 10484 62600
rect 13516 62560 13556 62600
rect 13996 62560 14036 62600
rect 1420 62308 1460 62348
rect 2860 62476 2900 62516
rect 5644 62476 5684 62516
rect 6316 62476 6356 62516
rect 7564 62476 7604 62516
rect 10156 62476 10196 62516
rect 4204 62392 4244 62432
rect 5932 62392 5972 62432
rect 2764 62308 2804 62348
rect 2956 62308 2996 62348
rect 3628 62308 3668 62348
rect 2284 62140 2324 62180
rect 1516 62056 1556 62096
rect 8044 62392 8084 62432
rect 8524 62392 8564 62432
rect 10060 62392 10100 62432
rect 12268 62476 12308 62516
rect 12748 62476 12788 62516
rect 13996 62392 14036 62432
rect 14380 62392 14420 62432
rect 15244 62392 15284 62432
rect 18028 62560 18068 62600
rect 18796 62560 18836 62600
rect 17260 62476 17300 62516
rect 18604 62476 18644 62516
rect 20044 62392 20084 62432
rect 4012 62308 4052 62348
rect 4492 62308 4532 62348
rect 5356 62308 5396 62348
rect 6316 62224 6356 62264
rect 7372 62308 7412 62348
rect 8716 62308 8756 62348
rect 9484 62308 9524 62348
rect 10828 62308 10868 62348
rect 11692 62308 11732 62348
rect 12172 62308 12212 62348
rect 9964 62224 10004 62264
rect 15724 62308 15764 62348
rect 16012 62308 16052 62348
rect 16684 62308 16724 62348
rect 18220 62308 18260 62348
rect 19564 62308 19604 62348
rect 15244 62224 15284 62264
rect 15916 62224 15956 62264
rect 16492 62224 16532 62264
rect 5548 62140 5588 62180
rect 6604 62140 6644 62180
rect 7756 62140 7796 62180
rect 10828 62140 10868 62180
rect 11500 62140 11540 62180
rect 14380 62140 14420 62180
rect 9964 62056 10004 62096
rect 2188 61972 2228 62012
rect 4928 61972 4968 62012
rect 5010 61972 5050 62012
rect 5092 61972 5132 62012
rect 5174 61972 5214 62012
rect 5256 61972 5296 62012
rect 7468 61972 7508 62012
rect 9484 61972 9524 62012
rect 1036 61888 1076 61928
rect 7564 61888 7604 61928
rect 14668 62140 14708 62180
rect 15820 62140 15860 62180
rect 18124 62140 18164 62180
rect 19564 62140 19604 62180
rect 20908 62140 20948 62180
rect 18796 61972 18836 62012
rect 20048 61972 20088 62012
rect 20130 61972 20170 62012
rect 20212 61972 20252 62012
rect 20294 61972 20334 62012
rect 20376 61972 20416 62012
rect 16876 61888 16916 61928
rect 17932 61888 17972 61928
rect 4780 61804 4820 61844
rect 6316 61804 6356 61844
rect 7372 61804 7412 61844
rect 10732 61804 10772 61844
rect 11116 61804 11156 61844
rect 12268 61804 12308 61844
rect 13612 61804 13652 61844
rect 17356 61804 17396 61844
rect 18508 61804 18548 61844
rect 20716 61804 20756 61844
rect 2956 61720 2996 61760
rect 5644 61720 5684 61760
rect 12844 61720 12884 61760
rect 16204 61720 16244 61760
rect 2764 61636 2804 61676
rect 3340 61636 3380 61676
rect 4204 61636 4244 61676
rect 4492 61667 4532 61676
rect 4492 61636 4532 61667
rect 4780 61636 4820 61676
rect 5452 61636 5492 61676
rect 6124 61636 6164 61676
rect 6700 61636 6740 61676
rect 9868 61636 9908 61676
rect 10156 61636 10196 61676
rect 652 61552 692 61592
rect 4012 61552 4052 61592
rect 5548 61552 5588 61592
rect 7756 61552 7796 61592
rect 172 61384 212 61424
rect 3532 61384 3572 61424
rect 1996 61216 2036 61256
rect 3688 61216 3728 61256
rect 3770 61216 3810 61256
rect 3852 61216 3892 61256
rect 3934 61216 3974 61256
rect 4016 61216 4056 61256
rect 2572 60964 2612 61004
rect 10828 61636 10868 61676
rect 12172 61636 12212 61676
rect 13420 61667 13460 61676
rect 13420 61636 13460 61667
rect 13708 61636 13748 61676
rect 15436 61636 15476 61676
rect 17068 61636 17108 61676
rect 21100 61888 21140 61928
rect 21100 61720 21140 61760
rect 11116 61552 11156 61592
rect 12844 61552 12884 61592
rect 15820 61552 15860 61592
rect 16300 61552 16340 61592
rect 18124 61636 18164 61676
rect 18604 61636 18644 61676
rect 19468 61667 19508 61676
rect 19468 61636 19508 61667
rect 16876 61552 16916 61592
rect 18028 61552 18068 61592
rect 18988 61552 19028 61592
rect 11500 61468 11540 61508
rect 12940 61468 12980 61508
rect 16396 61468 16436 61508
rect 17356 61468 17396 61508
rect 12172 61384 12212 61424
rect 14380 61384 14420 61424
rect 8812 61216 8852 61256
rect 13612 61132 13652 61172
rect 11116 61048 11156 61088
rect 14188 61048 14228 61088
rect 7564 60964 7604 61004
rect 7756 60964 7796 61004
rect 1612 60880 1652 60920
rect 3436 60880 3476 60920
rect 4012 60880 4052 60920
rect 8332 60880 8372 60920
rect 8524 60880 8564 60920
rect 18808 61216 18848 61256
rect 18890 61216 18930 61256
rect 18972 61216 19012 61256
rect 19054 61216 19094 61256
rect 19136 61216 19176 61256
rect 21388 61384 21428 61424
rect 16396 61048 16436 61088
rect 17932 60964 17972 61004
rect 11596 60880 11636 60920
rect 1996 60796 2036 60836
rect 2668 60796 2708 60836
rect 3148 60796 3188 60836
rect 3820 60796 3860 60836
rect 4588 60796 4628 60836
rect 5548 60796 5588 60836
rect 7276 60796 7316 60836
rect 8716 60796 8756 60836
rect 9484 60796 9524 60836
rect 10060 60796 10100 60836
rect 10348 60796 10388 60836
rect 12172 60796 12212 60836
rect 13996 60796 14036 60836
rect 17740 60880 17780 60920
rect 16684 60796 16724 60836
rect 18220 60880 18260 60920
rect 19180 60880 19220 60920
rect 21484 60880 21524 60920
rect 3916 60712 3956 60752
rect 2668 60628 2708 60668
rect 2956 60628 2996 60668
rect 4012 60628 4052 60668
rect 4588 60628 4628 60668
rect 940 60544 980 60584
rect 1516 60544 1556 60584
rect 12652 60712 12692 60752
rect 9772 60628 9812 60668
rect 18220 60628 18260 60668
rect 4928 60460 4968 60500
rect 5010 60460 5050 60500
rect 5092 60460 5132 60500
rect 5174 60460 5214 60500
rect 5256 60460 5296 60500
rect 7276 60460 7316 60500
rect 12652 60460 12692 60500
rect 16204 60460 16244 60500
rect 16684 60460 16724 60500
rect 20048 60460 20088 60500
rect 20130 60460 20170 60500
rect 20212 60460 20252 60500
rect 20294 60460 20334 60500
rect 20376 60460 20416 60500
rect 5356 60376 5396 60416
rect 1324 60208 1364 60248
rect 20716 60376 20756 60416
rect 1996 60292 2036 60332
rect 4396 60292 4436 60332
rect 5548 60292 5588 60332
rect 8236 60292 8276 60332
rect 12652 60292 12692 60332
rect 17260 60292 17300 60332
rect 2284 60208 2324 60248
rect 12268 60208 12308 60248
rect 16204 60208 16244 60248
rect 19468 60208 19508 60248
rect 2476 60124 2516 60164
rect 2764 60124 2804 60164
rect 3340 60124 3380 60164
rect 3532 60124 3572 60164
rect 4012 60124 4052 60164
rect 5644 60124 5684 60164
rect 5932 60124 5972 60164
rect 6124 60124 6164 60164
rect 10060 60124 10100 60164
rect 10732 60124 10772 60164
rect 15532 60124 15572 60164
rect 16396 60124 16436 60164
rect 17068 60124 17099 60164
rect 17099 60124 17108 60164
rect 17356 60124 17396 60164
rect 17836 60124 17867 60164
rect 17867 60124 17876 60164
rect 18508 60124 18548 60164
rect 19660 60124 19700 60164
rect 76 60040 116 60080
rect 2860 60040 2900 60080
rect 10924 60040 10964 60080
rect 12460 60040 12500 60080
rect 13132 60040 13172 60080
rect 14380 60040 14420 60080
rect 14668 60040 14708 60080
rect 14956 60040 14996 60080
rect 15436 60040 15476 60080
rect 15820 60040 15860 60080
rect 2092 59956 2132 59996
rect 3724 59956 3764 59996
rect 4012 59956 4052 59996
rect 268 59872 308 59912
rect 1900 59536 1940 59576
rect 1420 59368 1460 59408
rect 3688 59704 3728 59744
rect 3770 59704 3810 59744
rect 3852 59704 3892 59744
rect 3934 59704 3974 59744
rect 4016 59704 4056 59744
rect 8812 59956 8852 59996
rect 11212 59956 11252 59996
rect 5644 59872 5684 59912
rect 7276 59872 7316 59912
rect 8620 59872 8660 59912
rect 12172 59872 12212 59912
rect 12652 59872 12692 59912
rect 5740 59788 5780 59828
rect 6124 59788 6164 59828
rect 10828 59788 10868 59828
rect 20044 60124 20084 60164
rect 16204 60040 16244 60080
rect 18316 60040 18356 60080
rect 19180 60040 19220 60080
rect 17548 59956 17588 59996
rect 20428 59956 20468 59996
rect 16972 59872 17012 59912
rect 17452 59872 17492 59912
rect 18412 59872 18452 59912
rect 19660 59872 19700 59912
rect 21292 59872 21332 59912
rect 18808 59704 18848 59744
rect 18890 59704 18930 59744
rect 18972 59704 19012 59744
rect 19054 59704 19094 59744
rect 19136 59704 19176 59744
rect 6700 59620 6740 59660
rect 11116 59620 11156 59660
rect 3628 59536 3668 59576
rect 7852 59536 7892 59576
rect 8140 59536 8180 59576
rect 9292 59536 9332 59576
rect 12940 59536 12980 59576
rect 15916 59536 15956 59576
rect 16396 59536 16436 59576
rect 20044 59536 20084 59576
rect 3724 59452 3764 59492
rect 6124 59452 6164 59492
rect 6316 59452 6356 59492
rect 10828 59452 10868 59492
rect 11788 59452 11828 59492
rect 15532 59452 15572 59492
rect 18796 59452 18836 59492
rect 19468 59452 19508 59492
rect 3916 59368 3956 59408
rect 5740 59368 5780 59408
rect 5932 59368 5972 59408
rect 8044 59368 8084 59408
rect 11212 59368 11252 59408
rect 12172 59368 12212 59408
rect 18028 59368 18068 59408
rect 2284 59284 2324 59324
rect 3436 59284 3476 59324
rect 4396 59284 4436 59324
rect 6124 59284 6164 59324
rect 6604 59284 6644 59324
rect 7276 59284 7316 59324
rect 8620 59284 8660 59324
rect 9004 59284 9044 59324
rect 10348 59284 10388 59324
rect 10828 59284 10868 59324
rect 12940 59284 12980 59324
rect 14380 59284 14420 59324
rect 14956 59284 14996 59324
rect 16396 59284 16436 59324
rect 16588 59284 16628 59324
rect 18604 59284 18644 59324
rect 1804 59200 1844 59240
rect 3820 59200 3860 59240
rect 6412 59200 6452 59240
rect 7852 59200 7892 59240
rect 12268 59200 12308 59240
rect 20428 59368 20468 59408
rect 19468 59284 19508 59324
rect 21292 59200 21332 59240
rect 748 59116 788 59156
rect 3052 59116 3092 59156
rect 8620 59116 8660 59156
rect 10156 59116 10196 59156
rect 10828 59116 10868 59156
rect 18028 59116 18068 59156
rect 7564 59032 7604 59072
rect 16300 59032 16340 59072
rect 2764 58948 2804 58988
rect 4928 58948 4968 58988
rect 5010 58948 5050 58988
rect 5092 58948 5132 58988
rect 5174 58948 5214 58988
rect 5256 58948 5296 58988
rect 5932 58948 5972 58988
rect 13708 58948 13748 58988
rect 20048 58948 20088 58988
rect 20130 58948 20170 58988
rect 20212 58948 20252 58988
rect 20294 58948 20334 58988
rect 20376 58948 20416 58988
rect 556 58864 596 58904
rect 1612 58612 1652 58652
rect 3916 58780 3956 58820
rect 4876 58780 4916 58820
rect 5836 58780 5876 58820
rect 2668 58696 2708 58736
rect 2860 58696 2900 58736
rect 3436 58696 3476 58736
rect 2476 58612 2516 58652
rect 2764 58612 2804 58652
rect 3340 58643 3380 58652
rect 3340 58612 3380 58643
rect 3820 58643 3860 58652
rect 3820 58612 3860 58643
rect 4876 58612 4916 58652
rect 5644 58612 5684 58652
rect 6028 58612 6068 58652
rect 2668 58528 2708 58568
rect 3916 58528 3956 58568
rect 5548 58528 5588 58568
rect 2380 58444 2420 58484
rect 652 58360 692 58400
rect 1420 58360 1460 58400
rect 460 58192 500 58232
rect 7180 58864 7220 58904
rect 8812 58864 8852 58904
rect 9292 58864 9332 58904
rect 9484 58864 9524 58904
rect 11692 58864 11732 58904
rect 12076 58864 12116 58904
rect 14764 58864 14804 58904
rect 16012 58864 16052 58904
rect 18220 58864 18260 58904
rect 8524 58696 8564 58736
rect 9676 58696 9716 58736
rect 8620 58612 8651 58652
rect 8651 58612 8660 58652
rect 13036 58780 13076 58820
rect 16204 58780 16244 58820
rect 17836 58780 17876 58820
rect 12172 58696 12212 58736
rect 14956 58696 14996 58736
rect 15916 58696 15956 58736
rect 17260 58696 17300 58736
rect 17452 58696 17492 58736
rect 9292 58612 9332 58652
rect 10540 58612 10564 58652
rect 10564 58612 10580 58652
rect 11116 58612 11153 58652
rect 11153 58612 11156 58652
rect 11500 58612 11540 58652
rect 13996 58612 14036 58652
rect 14380 58612 14420 58652
rect 9004 58528 9044 58568
rect 9580 58528 9620 58568
rect 10156 58528 10196 58568
rect 10828 58528 10868 58568
rect 10924 58444 10964 58484
rect 11212 58444 11252 58484
rect 10444 58360 10484 58400
rect 3688 58192 3728 58232
rect 3770 58192 3810 58232
rect 3852 58192 3892 58232
rect 3934 58192 3974 58232
rect 4016 58192 4056 58232
rect 5548 58024 5588 58064
rect 11116 58108 11156 58148
rect 10540 58024 10580 58064
rect 13132 58528 13172 58568
rect 12172 58444 12212 58484
rect 13420 58444 13460 58484
rect 14476 58444 14516 58484
rect 14188 58360 14228 58400
rect 15052 58276 15092 58316
rect 12076 58192 12116 58232
rect 11788 58024 11828 58064
rect 14284 58024 14324 58064
rect 14956 58024 14996 58064
rect 6700 57940 6740 57980
rect 10924 57940 10964 57980
rect 14572 57940 14612 57980
rect 15052 57940 15092 57980
rect 3436 57856 3476 57896
rect 4204 57856 4244 57896
rect 7084 57856 7124 57896
rect 9004 57856 9044 57896
rect 11020 57856 11060 57896
rect 1324 57772 1364 57812
rect 4012 57772 4052 57812
rect 4876 57772 4916 57812
rect 14668 57856 14708 57896
rect 5644 57772 5676 57812
rect 5676 57772 5684 57812
rect 6892 57772 6932 57812
rect 7852 57772 7892 57812
rect 8140 57772 8180 57812
rect 8620 57772 8660 57812
rect 9196 57772 9236 57812
rect 10540 57772 10580 57812
rect 11116 57772 11156 57812
rect 11308 57772 11348 57812
rect 12556 57772 12596 57812
rect 13324 57772 13364 57812
rect 13900 57772 13940 57812
rect 10924 57688 10964 57728
rect 2476 57604 2516 57644
rect 6412 57604 6452 57644
rect 8044 57604 8084 57644
rect 9292 57604 9332 57644
rect 12076 57688 12116 57728
rect 16012 58612 16052 58652
rect 16876 58612 16916 58652
rect 17548 58612 17588 58652
rect 18796 58696 18836 58736
rect 18028 58612 18068 58652
rect 19564 58612 19604 58652
rect 16300 58528 16340 58568
rect 18412 58528 18452 58568
rect 17356 58360 17387 58400
rect 17387 58360 17396 58400
rect 18220 58360 18260 58400
rect 21100 58360 21140 58400
rect 19372 58276 19412 58316
rect 18808 58192 18848 58232
rect 18890 58192 18930 58232
rect 18972 58192 19012 58232
rect 19054 58192 19094 58232
rect 19136 58192 19176 58232
rect 15820 58024 15860 58064
rect 16972 57940 17012 57980
rect 16684 57856 16724 57896
rect 18796 57856 18836 57896
rect 20716 57856 20756 57896
rect 16204 57772 16244 57812
rect 16492 57772 16532 57812
rect 16780 57772 16820 57812
rect 18028 57772 18068 57812
rect 18412 57772 18452 57812
rect 18892 57772 18932 57812
rect 10156 57604 10196 57644
rect 10828 57604 10868 57644
rect 14860 57604 14900 57644
rect 1516 57520 1556 57560
rect 11308 57520 11348 57560
rect 12076 57520 12116 57560
rect 12748 57520 12788 57560
rect 19852 57520 19892 57560
rect 4928 57436 4968 57476
rect 5010 57436 5050 57476
rect 5092 57436 5132 57476
rect 5174 57436 5214 57476
rect 5256 57436 5296 57476
rect 5356 57436 5396 57476
rect 13036 57436 13076 57476
rect 20048 57436 20088 57476
rect 20130 57436 20170 57476
rect 20212 57436 20252 57476
rect 20294 57436 20334 57476
rect 20376 57436 20416 57476
rect 14188 57352 14228 57392
rect 2668 57268 2708 57308
rect 3148 57268 3188 57308
rect 10828 57268 10868 57308
rect 172 57184 212 57224
rect 3052 57184 3092 57224
rect 5932 57184 5972 57224
rect 2668 57100 2708 57140
rect 3436 57100 3476 57140
rect 5548 57100 5588 57140
rect 1804 57016 1844 57056
rect 1996 57016 2036 57056
rect 4588 57016 4628 57056
rect 9484 57184 9524 57224
rect 12556 57184 12596 57224
rect 6412 57131 6452 57140
rect 6412 57100 6452 57131
rect 7852 57100 7892 57140
rect 8524 57100 8564 57140
rect 2572 56932 2612 56972
rect 5644 56932 5684 56972
rect 6124 56932 6164 56972
rect 9292 57131 9332 57140
rect 9292 57100 9332 57131
rect 11116 57131 11156 57140
rect 11116 57100 11156 57131
rect 11788 57100 11828 57140
rect 12652 57100 12692 57140
rect 14476 57268 14516 57308
rect 15724 57268 15764 57308
rect 16300 57184 16340 57224
rect 13420 57100 13460 57140
rect 20620 57352 20660 57392
rect 16876 57268 16916 57308
rect 18508 57268 18548 57308
rect 18124 57184 18164 57224
rect 14284 57131 14324 57140
rect 14284 57100 14324 57131
rect 15436 57100 15476 57140
rect 15724 57100 15764 57140
rect 8428 57016 8468 57056
rect 13900 57016 13940 57056
rect 7852 56932 7892 56972
rect 13804 56932 13844 56972
rect 268 56848 308 56888
rect 460 56848 500 56888
rect 1324 56848 1364 56888
rect 1804 56848 1844 56888
rect 2668 56848 2708 56888
rect 9964 56848 10004 56888
rect 844 56764 884 56804
rect 3688 56680 3728 56720
rect 3770 56680 3810 56720
rect 3852 56680 3892 56720
rect 3934 56680 3974 56720
rect 4016 56680 4056 56720
rect 76 56512 116 56552
rect 3628 56512 3668 56552
rect 5932 56512 5972 56552
rect 6988 56764 7028 56804
rect 8332 56764 8372 56804
rect 13900 56764 13940 56804
rect 8332 56596 8372 56636
rect 12172 56596 12212 56636
rect 7852 56512 7892 56552
rect 10060 56512 10100 56552
rect 17164 57100 17204 57140
rect 20716 56932 20756 56972
rect 16876 56848 16916 56888
rect 18796 56848 18836 56888
rect 20812 56848 20852 56888
rect 3148 56344 3188 56384
rect 4204 56344 4244 56384
rect 6412 56344 6452 56384
rect 6604 56344 6644 56384
rect 7372 56344 7412 56384
rect 7756 56344 7796 56384
rect 844 56260 884 56300
rect 2956 56260 2996 56300
rect 3628 56260 3668 56300
rect 4492 56260 4532 56300
rect 4780 56260 4820 56300
rect 5356 56260 5396 56300
rect 5836 56260 5876 56300
rect 8332 56260 8372 56300
rect 9292 56260 9332 56300
rect 18808 56680 18848 56720
rect 18890 56680 18930 56720
rect 18972 56680 19012 56720
rect 19054 56680 19094 56720
rect 19136 56680 19176 56720
rect 9964 56344 10004 56384
rect 13420 56344 13460 56384
rect 13804 56344 13844 56384
rect 15820 56344 15860 56384
rect 16300 56344 16340 56384
rect 17068 56344 17108 56384
rect 17740 56344 17780 56384
rect 18796 56344 18836 56384
rect 10828 56260 10868 56300
rect 12076 56260 12116 56300
rect 12556 56260 12596 56300
rect 13900 56260 13940 56300
rect 14284 56260 14324 56300
rect 14860 56260 14868 56300
rect 14868 56260 14900 56300
rect 15052 56260 15092 56300
rect 15436 56260 15476 56300
rect 16012 56260 16052 56300
rect 16780 56260 16820 56300
rect 556 56176 596 56216
rect 5452 56176 5492 56216
rect 12268 56176 12308 56216
rect 12652 56176 12692 56216
rect 13420 56176 13460 56216
rect 14668 56176 14708 56216
rect 16300 56176 16340 56216
rect 17068 56176 17108 56216
rect 3052 56092 3092 56132
rect 5260 56092 5300 56132
rect 8620 56092 8660 56132
rect 9964 56092 10004 56132
rect 19852 56344 19892 56384
rect 20908 56344 20948 56384
rect 18508 56260 18548 56300
rect 19180 56260 19220 56300
rect 18220 56176 18260 56216
rect 21004 56176 21044 56216
rect 4928 55924 4968 55964
rect 5010 55924 5050 55964
rect 5092 55924 5132 55964
rect 5174 55924 5214 55964
rect 5256 55924 5296 55964
rect 20048 55924 20088 55964
rect 20130 55924 20170 55964
rect 20212 55924 20252 55964
rect 20294 55924 20334 55964
rect 20376 55924 20416 55964
rect 748 55840 788 55880
rect 4204 55840 4244 55880
rect 4492 55840 4532 55880
rect 9292 55840 9332 55880
rect 15340 55840 15380 55880
rect 19660 55840 19700 55880
rect 2284 55756 2324 55796
rect 3436 55756 3476 55796
rect 5356 55756 5396 55796
rect 6316 55756 6356 55796
rect 6892 55756 6932 55796
rect 9004 55756 9044 55796
rect 9580 55756 9620 55796
rect 2668 55672 2708 55712
rect 1996 55588 2036 55628
rect 2572 55588 2612 55628
rect 6412 55672 6452 55712
rect 7660 55672 7700 55712
rect 8908 55672 8948 55712
rect 10156 55672 10196 55712
rect 1420 55504 1460 55544
rect 2764 55336 2804 55376
rect 6700 55588 6740 55628
rect 9004 55588 9044 55628
rect 9676 55588 9716 55628
rect 9964 55619 10004 55628
rect 9964 55588 10004 55619
rect 12076 55588 12116 55628
rect 12748 55588 12788 55628
rect 13708 55588 13748 55628
rect 14188 55588 14228 55628
rect 15436 55588 15476 55628
rect 15820 55588 15860 55628
rect 16300 55588 16340 55628
rect 16876 55619 16916 55628
rect 16876 55588 16916 55619
rect 18124 55588 18164 55628
rect 18316 55588 18356 55628
rect 6508 55504 6548 55544
rect 8044 55504 8084 55544
rect 8812 55504 8852 55544
rect 12268 55504 12308 55544
rect 16012 55504 16052 55544
rect 17164 55504 17204 55544
rect 19660 55504 19700 55544
rect 14092 55420 14132 55460
rect 16588 55420 16628 55460
rect 20812 55420 20852 55460
rect 6220 55336 6260 55376
rect 7276 55336 7316 55376
rect 10924 55336 10964 55376
rect 14860 55336 14900 55376
rect 19852 55336 19892 55376
rect 20908 55336 20948 55376
rect 17068 55252 17108 55292
rect 20620 55252 20660 55292
rect 652 55168 692 55208
rect 3688 55168 3728 55208
rect 3770 55168 3810 55208
rect 3852 55168 3892 55208
rect 3934 55168 3974 55208
rect 4016 55168 4056 55208
rect 18808 55168 18848 55208
rect 18890 55168 18930 55208
rect 18972 55168 19012 55208
rect 19054 55168 19094 55208
rect 19136 55168 19176 55208
rect 2668 55084 2708 55124
rect 13324 55084 13364 55124
rect 1804 54832 1844 54872
rect 2860 54832 2900 54872
rect 3724 54832 3764 54872
rect 4204 54832 4244 54872
rect 11788 55000 11828 55040
rect 13420 55000 13460 55040
rect 15052 55000 15092 55040
rect 16780 55000 16820 55040
rect 18892 55000 18932 55040
rect 9676 54916 9716 54956
rect 12172 54916 12212 54956
rect 12844 54916 12884 54956
rect 19948 54916 19988 54956
rect 9580 54832 9620 54872
rect 10732 54832 10772 54872
rect 16300 54832 16340 54872
rect 18316 54832 18356 54872
rect 20716 54832 20756 54872
rect 2284 54748 2324 54788
rect 2572 54748 2612 54788
rect 4492 54748 4532 54788
rect 5548 54748 5588 54788
rect 6028 54748 6068 54788
rect 6892 54748 6932 54788
rect 9004 54748 9044 54788
rect 9196 54748 9236 54788
rect 9676 54748 9716 54788
rect 10444 54748 10484 54788
rect 11308 54748 11348 54788
rect 11788 54748 11828 54788
rect 13324 54748 13364 54788
rect 13708 54748 13748 54788
rect 14860 54748 14900 54788
rect 15724 54748 15764 54788
rect 17164 54748 17204 54788
rect 18412 54748 18452 54788
rect 19468 54748 19508 54788
rect 3628 54664 3659 54704
rect 3659 54664 3668 54704
rect 3916 54664 3956 54704
rect 3052 54580 3092 54620
rect 3532 54580 3572 54620
rect 4204 54580 4244 54620
rect 7756 54580 7796 54620
rect 9292 54580 9332 54620
rect 2764 54496 2804 54536
rect 3916 54496 3956 54536
rect 4928 54412 4968 54452
rect 5010 54412 5050 54452
rect 5092 54412 5132 54452
rect 5174 54412 5214 54452
rect 5256 54412 5296 54452
rect 3532 54328 3572 54368
rect 1708 54244 1748 54284
rect 3820 54244 3860 54284
rect 1324 54160 1364 54200
rect 3724 54160 3764 54200
rect 2092 54076 2132 54116
rect 2476 54076 2516 54116
rect 3628 54076 3668 54116
rect 16684 54664 16724 54704
rect 17260 54664 17300 54704
rect 18508 54580 18548 54620
rect 8812 54496 8852 54536
rect 9964 54496 10004 54536
rect 19084 54496 19124 54536
rect 13612 54412 13652 54452
rect 20048 54412 20088 54452
rect 20130 54412 20170 54452
rect 20212 54412 20252 54452
rect 20294 54412 20334 54452
rect 20376 54412 20416 54452
rect 14764 54328 14804 54368
rect 6220 54244 6260 54284
rect 7276 54244 7316 54284
rect 7948 54244 7988 54284
rect 8524 54244 8564 54284
rect 9004 54244 9044 54284
rect 11308 54244 11348 54284
rect 12940 54244 12980 54284
rect 14956 54244 14996 54284
rect 7852 54160 7892 54200
rect 9580 54160 9620 54200
rect 4204 54076 4233 54116
rect 4233 54076 4244 54116
rect 4492 54076 4532 54116
rect 5740 54107 5780 54116
rect 5740 54076 5780 54107
rect 7180 54076 7220 54116
rect 11788 54160 11828 54200
rect 18892 54328 18932 54368
rect 20620 54328 20660 54368
rect 1708 53992 1748 54032
rect 3916 53992 3956 54032
rect 460 53824 500 53864
rect 652 53824 692 53864
rect 7756 54107 7796 54116
rect 7756 54076 7796 54107
rect 9292 54076 9332 54116
rect 9676 54076 9716 54116
rect 10444 54107 10484 54116
rect 10444 54076 10484 54107
rect 10924 54107 10964 54116
rect 10924 54076 10964 54107
rect 14092 54076 14132 54116
rect 8908 53992 8948 54032
rect 9964 53992 10004 54032
rect 15244 54076 15284 54116
rect 15628 54076 15668 54116
rect 16012 54076 16052 54116
rect 16588 54076 16628 54116
rect 17932 54076 17972 54116
rect 13324 53992 13364 54032
rect 15820 53992 15860 54032
rect 4204 53908 4244 53948
rect 5932 53908 5972 53948
rect 7180 53908 7220 53948
rect 8812 53908 8852 53948
rect 15724 53908 15764 53948
rect 3724 53824 3755 53864
rect 3755 53824 3764 53864
rect 6604 53824 6644 53864
rect 10060 53824 10100 53864
rect 10348 53824 10388 53864
rect 10636 53824 10676 53864
rect 11500 53824 11540 53864
rect 1900 53656 1940 53696
rect 3688 53656 3728 53696
rect 3770 53656 3810 53696
rect 3852 53656 3892 53696
rect 3934 53656 3974 53696
rect 4016 53656 4056 53696
rect 5740 53656 5780 53696
rect 6988 53656 7028 53696
rect 12652 53656 12692 53696
rect 5932 53572 5972 53612
rect 9964 53572 10004 53612
rect 14572 53572 14612 53612
rect 556 53488 596 53528
rect 2188 53488 2228 53528
rect 12748 53488 12788 53528
rect 14380 53488 14420 53528
rect 18508 54160 18548 54200
rect 18604 54076 18644 54116
rect 18796 54076 18836 54116
rect 19084 54076 19124 54116
rect 19468 54076 19508 54116
rect 19852 54107 19892 54116
rect 19852 54076 19892 54107
rect 18892 53992 18932 54032
rect 18796 53824 18836 53864
rect 21004 53824 21044 53864
rect 18808 53656 18848 53696
rect 18890 53656 18930 53696
rect 18972 53656 19012 53696
rect 19054 53656 19094 53696
rect 19136 53656 19176 53696
rect 17164 53572 17204 53612
rect 3052 53404 3092 53444
rect 3244 53404 3284 53444
rect 6892 53404 6932 53444
rect 7276 53404 7316 53444
rect 8428 53404 8468 53444
rect 10060 53404 10100 53444
rect 10444 53404 10484 53444
rect 10636 53404 10676 53444
rect 10924 53404 10964 53444
rect 11788 53404 11828 53444
rect 556 53320 596 53360
rect 2092 53320 2132 53360
rect 1324 53152 1364 53192
rect 652 52816 692 52856
rect 7180 53320 7220 53360
rect 10348 53320 10388 53360
rect 12460 53320 12500 53360
rect 13324 53320 13364 53360
rect 16012 53320 16052 53360
rect 16972 53320 17012 53360
rect 17452 53320 17492 53360
rect 18508 53320 18548 53360
rect 20812 53320 20852 53360
rect 4012 53236 4052 53276
rect 4204 53236 4212 53276
rect 4212 53236 4244 53276
rect 5548 53236 5588 53276
rect 5740 53236 5780 53276
rect 6604 53236 6644 53276
rect 7276 53236 7316 53276
rect 7852 53236 7892 53276
rect 8236 53236 8244 53276
rect 8244 53236 8276 53276
rect 9484 53236 9524 53276
rect 12844 53236 12884 53276
rect 14380 53236 14420 53276
rect 15628 53236 15668 53276
rect 16204 53236 16244 53276
rect 16684 53236 16724 53276
rect 18604 53236 18644 53276
rect 19084 53236 19124 53276
rect 19372 53236 19412 53276
rect 19948 53236 19988 53276
rect 2860 53152 2900 53192
rect 5836 53152 5876 53192
rect 9676 53152 9716 53192
rect 4396 53068 4436 53108
rect 6028 53068 6068 53108
rect 6604 53068 6644 53108
rect 9964 53068 10004 53108
rect 5356 52984 5396 53024
rect 9292 52984 9332 53024
rect 10732 52984 10772 53024
rect 4928 52900 4968 52940
rect 5010 52900 5050 52940
rect 5092 52900 5132 52940
rect 5174 52900 5214 52940
rect 5256 52900 5296 52940
rect 9484 52816 9524 52856
rect 19660 53068 19700 53108
rect 20048 52900 20088 52940
rect 20130 52900 20170 52940
rect 20212 52900 20252 52940
rect 20294 52900 20334 52940
rect 20376 52900 20416 52940
rect 20908 52816 20948 52856
rect 5740 52732 5780 52772
rect 6604 52732 6644 52772
rect 6892 52732 6932 52772
rect 10732 52732 10772 52772
rect 12844 52732 12884 52772
rect 19084 52732 19124 52772
rect 1708 52564 1748 52604
rect 2476 52595 2516 52604
rect 2476 52564 2516 52595
rect 4108 52564 4148 52604
rect 7372 52648 7412 52688
rect 9484 52648 9524 52688
rect 10540 52648 10580 52688
rect 13708 52648 13748 52688
rect 5548 52564 5588 52604
rect 6028 52564 6068 52604
rect 6316 52564 6356 52604
rect 6892 52595 6932 52604
rect 6892 52564 6932 52595
rect 652 52480 692 52520
rect 4684 52480 4724 52520
rect 5932 52480 5972 52520
rect 9292 52564 9332 52604
rect 9676 52595 9716 52604
rect 9676 52564 9716 52595
rect 9964 52564 10004 52604
rect 10444 52564 10484 52604
rect 8428 52480 8468 52520
rect 6508 52396 6548 52436
rect 9964 52396 10004 52436
rect 12748 52595 12788 52604
rect 12748 52564 12788 52595
rect 14188 52564 14228 52604
rect 17068 52648 17108 52688
rect 10348 52480 10388 52520
rect 10636 52480 10676 52520
rect 10924 52396 10964 52436
rect 3688 52144 3728 52184
rect 3770 52144 3810 52184
rect 3852 52144 3892 52184
rect 3934 52144 3974 52184
rect 4016 52144 4056 52184
rect 15724 52564 15764 52604
rect 17260 52564 17300 52604
rect 19948 52564 19988 52604
rect 19660 52480 19700 52520
rect 20140 52480 20180 52520
rect 17452 52396 17492 52436
rect 17836 52396 17876 52436
rect 19756 52396 19796 52436
rect 17644 52312 17684 52352
rect 18412 52312 18452 52352
rect 20428 52312 20468 52352
rect 16396 52144 16436 52184
rect 17260 52144 17300 52184
rect 18808 52144 18848 52184
rect 18890 52144 18930 52184
rect 18972 52144 19012 52184
rect 19054 52144 19094 52184
rect 19136 52144 19176 52184
rect 10444 52060 10484 52100
rect 14092 52060 14132 52100
rect 6028 51976 6068 52016
rect 8236 51976 8276 52016
rect 8716 51976 8756 52016
rect 10636 51976 10676 52016
rect 10924 51976 10964 52016
rect 2860 51892 2900 51932
rect 5548 51892 5588 51932
rect 556 51808 596 51848
rect 1804 51808 1844 51848
rect 2572 51808 2612 51848
rect 4396 51808 4436 51848
rect 7084 51808 7124 51848
rect 9964 51892 10004 51932
rect 12844 51892 12884 51932
rect 17260 51892 17300 51932
rect 9676 51808 9716 51848
rect 10540 51808 10580 51848
rect 11308 51808 11348 51848
rect 18316 51808 18356 51848
rect 20140 51808 20180 51848
rect 20428 51808 20468 51848
rect 2380 51640 2420 51680
rect 3628 51724 3668 51764
rect 6508 51724 6548 51764
rect 7948 51724 7988 51764
rect 9484 51724 9524 51764
rect 10060 51724 10091 51764
rect 10091 51724 10100 51764
rect 10348 51724 10359 51764
rect 10359 51724 10388 51764
rect 556 51556 596 51596
rect 652 51220 692 51260
rect 1324 51220 1364 51260
rect 556 51136 596 51176
rect 1996 50968 2036 51008
rect 2860 51556 2900 51596
rect 2572 50968 2612 51008
rect 4492 51640 4532 51680
rect 5356 51556 5396 51596
rect 4928 51388 4968 51428
rect 5010 51388 5050 51428
rect 5092 51388 5132 51428
rect 5174 51388 5214 51428
rect 5256 51388 5296 51428
rect 6316 51640 6356 51680
rect 6988 51640 7028 51680
rect 11884 51724 11924 51764
rect 12556 51724 12596 51764
rect 12748 51724 12788 51764
rect 8428 51640 8468 51680
rect 10156 51640 10196 51680
rect 12172 51640 12212 51680
rect 13228 51640 13268 51680
rect 16492 51640 16532 51680
rect 12748 51556 12788 51596
rect 15340 51556 15380 51596
rect 13132 51472 13172 51512
rect 12460 51220 12500 51260
rect 14380 51220 14420 51260
rect 16204 51220 16244 51260
rect 17452 51220 17492 51260
rect 4108 51052 4148 51092
rect 4492 51052 4532 51092
rect 5836 51052 5876 51092
rect 6508 51052 6548 51092
rect 7948 51052 7988 51092
rect 7180 50968 7220 51008
rect 7756 50968 7796 51008
rect 10828 51052 10868 51092
rect 11692 51052 11732 51092
rect 12748 51052 12788 51092
rect 15340 51052 15380 51092
rect 16204 51052 16244 51092
rect 16780 51083 16820 51092
rect 16780 51052 16820 51083
rect 19660 51556 19700 51596
rect 20048 51388 20088 51428
rect 20130 51388 20170 51428
rect 20212 51388 20252 51428
rect 20294 51388 20334 51428
rect 20376 51388 20416 51428
rect 19756 51220 19796 51260
rect 17644 51052 17684 51092
rect 10444 50968 10484 51008
rect 11020 50968 11060 51008
rect 11884 50968 11924 51008
rect 13228 50968 13268 51008
rect 15532 50968 15572 51008
rect 16300 50968 16340 51008
rect 21196 51052 21236 51092
rect 19372 50968 19412 51008
rect 21100 50968 21140 51008
rect 2380 50800 2420 50840
rect 8716 50800 8756 50840
rect 10348 50800 10388 50840
rect 11980 50800 12020 50840
rect 20716 50800 20756 50840
rect 7564 50716 7604 50756
rect 20236 50716 20276 50756
rect 2956 50632 2996 50672
rect 3688 50632 3728 50672
rect 3770 50632 3810 50672
rect 3852 50632 3892 50672
rect 3934 50632 3974 50672
rect 4016 50632 4056 50672
rect 4492 50632 4532 50672
rect 7756 50632 7796 50672
rect 18808 50632 18848 50672
rect 18890 50632 18930 50672
rect 18972 50632 19012 50672
rect 19054 50632 19094 50672
rect 19136 50632 19176 50672
rect 8332 50464 8372 50504
rect 11020 50464 11060 50504
rect 9196 50380 9236 50420
rect 11692 50380 11732 50420
rect 15628 50380 15668 50420
rect 19660 50380 19700 50420
rect 9004 50296 9044 50336
rect 10060 50296 10100 50336
rect 11404 50296 11444 50336
rect 12268 50296 12308 50336
rect 15916 50296 15956 50336
rect 16396 50296 16436 50336
rect 19468 50296 19508 50336
rect 20236 50296 20276 50336
rect 20716 50296 20756 50336
rect 4300 50212 4340 50252
rect 8140 50212 8180 50252
rect 8524 50212 8564 50252
rect 9772 50212 9812 50252
rect 10156 50212 10196 50252
rect 10348 50212 10388 50252
rect 12556 50212 12596 50252
rect 13996 50212 14036 50252
rect 16876 50212 16916 50252
rect 19180 50212 19220 50252
rect 19756 50212 19796 50252
rect 3532 50044 3572 50084
rect 5740 50044 5780 50084
rect 3340 49624 3380 49664
rect 4928 49876 4968 49916
rect 5010 49876 5050 49916
rect 5092 49876 5132 49916
rect 5174 49876 5214 49916
rect 5256 49876 5296 49916
rect 9292 50044 9332 50084
rect 11308 50044 11348 50084
rect 11884 50044 11924 50084
rect 15340 50044 15380 50084
rect 15820 50044 15860 50084
rect 14188 49792 14228 49832
rect 16204 50128 16244 50168
rect 16300 50044 16340 50084
rect 17068 50044 17108 50084
rect 20524 50128 20564 50168
rect 10924 49708 10964 49748
rect 20048 49876 20088 49916
rect 20130 49876 20170 49916
rect 20212 49876 20252 49916
rect 20294 49876 20334 49916
rect 20376 49876 20416 49916
rect 10444 49624 10484 49664
rect 11116 49624 11156 49664
rect 16204 49624 16244 49664
rect 6124 49540 6164 49580
rect 7180 49540 7220 49580
rect 7948 49540 7988 49580
rect 9484 49540 9524 49580
rect 9772 49540 9812 49580
rect 10156 49540 10196 49580
rect 10732 49571 10772 49580
rect 10732 49540 10772 49571
rect 11212 49571 11252 49580
rect 11212 49540 11252 49571
rect 13228 49571 13268 49580
rect 13228 49540 13268 49571
rect 15628 49571 15668 49580
rect 15628 49540 15668 49571
rect 16876 49540 16916 49580
rect 6508 49456 6548 49496
rect 10252 49456 10292 49496
rect 11308 49456 11348 49496
rect 19372 49456 19412 49496
rect 19948 49456 19988 49496
rect 4108 49372 4148 49412
rect 6220 49372 6260 49412
rect 12844 49372 12884 49412
rect 16300 49372 16340 49412
rect 4684 49288 4724 49328
rect 6604 49288 6644 49328
rect 13420 49288 13460 49328
rect 17644 49288 17684 49328
rect 20428 49288 20468 49328
rect 15724 49204 15764 49244
rect 3688 49120 3728 49160
rect 3770 49120 3810 49160
rect 3852 49120 3892 49160
rect 3934 49120 3974 49160
rect 4016 49120 4056 49160
rect 18808 49120 18848 49160
rect 18890 49120 18930 49160
rect 18972 49120 19012 49160
rect 19054 49120 19094 49160
rect 19136 49120 19176 49160
rect 11212 48952 11252 48992
rect 15820 48952 15860 48992
rect 19468 48952 19508 48992
rect 4204 48868 4244 48908
rect 8620 48868 8660 48908
rect 14476 48868 14516 48908
rect 18220 48868 18260 48908
rect 19756 48868 19796 48908
rect 20428 48868 20468 48908
rect 2764 48784 2804 48824
rect 4780 48784 4820 48824
rect 8908 48784 8948 48824
rect 9196 48784 9236 48824
rect 9676 48784 9716 48824
rect 11980 48784 12020 48824
rect 12172 48784 12212 48824
rect 15532 48784 15572 48824
rect 5644 48700 5684 48740
rect 4396 48616 4436 48656
rect 4204 48532 4244 48572
rect 6124 48700 6164 48740
rect 6604 48700 6612 48740
rect 6612 48700 6644 48740
rect 7180 48700 7220 48740
rect 7948 48700 7988 48740
rect 8812 48700 8852 48740
rect 9964 48700 10004 48740
rect 10636 48700 10676 48740
rect 12268 48700 12308 48740
rect 12748 48700 12788 48740
rect 13420 48700 13460 48740
rect 15340 48700 15371 48740
rect 15371 48700 15380 48740
rect 15820 48700 15860 48740
rect 12652 48616 12692 48656
rect 6796 48532 6836 48572
rect 13516 48532 13556 48572
rect 15820 48532 15860 48572
rect 5836 48448 5876 48488
rect 8236 48448 8276 48488
rect 4928 48364 4968 48404
rect 5010 48364 5050 48404
rect 5092 48364 5132 48404
rect 5174 48364 5214 48404
rect 5256 48364 5296 48404
rect 4492 48196 4532 48236
rect 6412 48196 6452 48236
rect 1996 48112 2036 48152
rect 3244 48112 3284 48152
rect 7468 48112 7508 48152
rect 2668 48028 2708 48068
rect 3340 48028 3380 48068
rect 4108 48028 4148 48068
rect 4588 48028 4628 48068
rect 17548 48784 17588 48824
rect 18316 48784 18356 48824
rect 18604 48784 18644 48824
rect 16396 48700 16436 48740
rect 19372 48784 19412 48824
rect 20524 48784 20564 48824
rect 21100 48784 21140 48824
rect 18220 48700 18260 48740
rect 19468 48700 19508 48740
rect 16972 48616 17012 48656
rect 18316 48616 18356 48656
rect 20812 48532 20852 48572
rect 20048 48364 20088 48404
rect 20130 48364 20170 48404
rect 20212 48364 20252 48404
rect 20294 48364 20334 48404
rect 20376 48364 20416 48404
rect 17452 48196 17492 48236
rect 5740 48059 5780 48068
rect 5740 48028 5780 48059
rect 12940 48028 12980 48068
rect 13228 48028 13268 48068
rect 14284 48028 14324 48068
rect 16204 48028 16244 48068
rect 16396 48028 16436 48068
rect 2188 47944 2228 47984
rect 2764 47944 2804 47984
rect 4204 47944 4244 47984
rect 4876 47944 4916 47984
rect 8044 47944 8084 47984
rect 11308 47944 11348 47984
rect 15820 47944 15860 47984
rect 17260 48059 17300 48068
rect 17260 48028 17300 48059
rect 16300 47944 16340 47984
rect 8908 47860 8948 47900
rect 10636 47860 10676 47900
rect 16780 47860 16820 47900
rect 8140 47776 8180 47816
rect 8812 47776 8852 47816
rect 10540 47776 10580 47816
rect 10732 47776 10772 47816
rect 14956 47776 14996 47816
rect 6316 47692 6356 47732
rect 19276 48028 19316 48068
rect 19756 47944 19796 47984
rect 20140 47944 20180 47984
rect 3688 47608 3728 47648
rect 3770 47608 3810 47648
rect 3852 47608 3892 47648
rect 3934 47608 3974 47648
rect 4016 47608 4056 47648
rect 10732 47608 10772 47648
rect 18808 47608 18848 47648
rect 18890 47608 18930 47648
rect 18972 47608 19012 47648
rect 19054 47608 19094 47648
rect 19136 47608 19176 47648
rect 3340 47440 3380 47480
rect 9388 47440 9428 47480
rect 15820 47440 15860 47480
rect 17260 47440 17300 47480
rect 19468 47440 19508 47480
rect 3244 47356 3284 47396
rect 7660 47356 7700 47396
rect 10828 47356 10868 47396
rect 3532 47272 3572 47312
rect 2860 47188 2900 47228
rect 3436 47188 3476 47228
rect 3916 47188 3956 47228
rect 11500 47272 11540 47312
rect 19660 47272 19700 47312
rect 4684 47188 4724 47228
rect 4780 47020 4820 47060
rect 5644 47020 5684 47060
rect 4928 46852 4968 46892
rect 5010 46852 5050 46892
rect 5092 46852 5132 46892
rect 5174 46852 5214 46892
rect 5256 46852 5296 46892
rect 8620 47188 8660 47228
rect 9388 47188 9428 47228
rect 10444 47188 10484 47228
rect 11596 47188 11636 47228
rect 12268 47188 12308 47228
rect 12844 47188 12884 47228
rect 13996 47188 14036 47228
rect 14572 47188 14612 47228
rect 15628 47188 15668 47228
rect 15820 47188 15860 47228
rect 18028 47188 18068 47228
rect 19276 47188 19316 47228
rect 20524 47188 20564 47228
rect 8908 47020 8948 47060
rect 8524 46936 8564 46976
rect 12556 47020 12596 47060
rect 11212 46936 11252 46976
rect 14188 47020 14228 47060
rect 15820 46852 15860 46892
rect 20048 46852 20088 46892
rect 20130 46852 20170 46892
rect 20212 46852 20252 46892
rect 20294 46852 20334 46892
rect 20376 46852 20416 46892
rect 2188 46684 2228 46724
rect 3340 46684 3380 46724
rect 4684 46684 4724 46724
rect 9388 46684 9428 46724
rect 10348 46684 10388 46724
rect 11692 46768 11732 46808
rect 12076 46768 12116 46808
rect 14764 46684 14804 46724
rect 2860 46516 2900 46556
rect 5356 46516 5396 46556
rect 3436 46432 3476 46472
rect 4492 46432 4532 46472
rect 8140 46600 8180 46640
rect 13996 46600 14036 46640
rect 6700 46516 6740 46556
rect 6988 46516 7028 46556
rect 7180 46516 7220 46556
rect 7468 46516 7508 46556
rect 8908 46516 8948 46556
rect 9580 46516 9620 46556
rect 10252 46516 10292 46556
rect 11116 46516 11156 46556
rect 11308 46516 11348 46556
rect 11500 46516 11540 46556
rect 12556 46516 12596 46556
rect 13612 46516 13652 46556
rect 13900 46516 13940 46556
rect 14476 46547 14516 46556
rect 14476 46516 14516 46547
rect 14956 46547 14996 46556
rect 14956 46516 14996 46547
rect 16876 46516 16916 46556
rect 17548 46516 17588 46556
rect 9772 46432 9812 46472
rect 10444 46432 10484 46472
rect 10636 46432 10676 46472
rect 10828 46432 10868 46472
rect 13420 46432 13460 46472
rect 14380 46432 14420 46472
rect 17356 46432 17396 46472
rect 20140 46432 20180 46472
rect 4300 46348 4340 46388
rect 4972 46348 4975 46388
rect 4975 46348 5012 46388
rect 5356 46348 5396 46388
rect 11500 46348 11540 46388
rect 14476 46348 14516 46388
rect 17260 46348 17300 46388
rect 20620 46348 20660 46388
rect 4204 46264 4244 46304
rect 6604 46264 6644 46304
rect 10828 46264 10868 46304
rect 11692 46264 11732 46304
rect 12268 46264 12308 46304
rect 12556 46264 12596 46304
rect 15340 46264 15380 46304
rect 19276 46264 19316 46304
rect 17548 46180 17588 46220
rect 2284 46096 2324 46136
rect 3688 46096 3728 46136
rect 3770 46096 3810 46136
rect 3852 46096 3892 46136
rect 3934 46096 3974 46136
rect 4016 46096 4056 46136
rect 5452 46096 5492 46136
rect 6700 46096 6740 46136
rect 18808 46096 18848 46136
rect 18890 46096 18930 46136
rect 18972 46096 19012 46136
rect 19054 46096 19094 46136
rect 19136 46096 19176 46136
rect 5260 46012 5300 46052
rect 5740 46012 5780 46052
rect 6220 46012 6260 46052
rect 8236 46012 8276 46052
rect 18412 46012 18452 46052
rect 3916 45928 3956 45968
rect 5452 45928 5492 45968
rect 6412 45928 6452 45968
rect 7852 45928 7892 45968
rect 9772 45928 9812 45968
rect 10156 45928 10196 45968
rect 10636 45928 10676 45968
rect 13420 45928 13460 45968
rect 15052 45928 15092 45968
rect 19564 45928 19604 45968
rect 4780 45844 4820 45884
rect 5164 45844 5204 45884
rect 76 45760 116 45800
rect 4012 45760 4052 45800
rect 4492 45760 4532 45800
rect 4684 45760 4724 45800
rect 76 45424 116 45464
rect 5260 45760 5300 45800
rect 7180 45844 7220 45884
rect 8140 45844 8180 45884
rect 20524 45844 20564 45884
rect 6796 45760 6836 45800
rect 8428 45760 8468 45800
rect 10156 45760 10196 45800
rect 11788 45760 11828 45800
rect 12940 45760 12980 45800
rect 14188 45760 14228 45800
rect 14380 45760 14420 45800
rect 17548 45760 17588 45800
rect 18316 45760 18356 45800
rect 19564 45760 19604 45800
rect 20620 45760 20660 45800
rect 3916 45676 3956 45716
rect 4108 45676 4148 45716
rect 5068 45676 5108 45716
rect 5932 45676 5972 45716
rect 6412 45676 6452 45716
rect 6604 45676 6644 45716
rect 8236 45676 8276 45716
rect 9388 45676 9428 45716
rect 11596 45676 11636 45716
rect 13228 45676 13268 45716
rect 13516 45676 13556 45716
rect 14860 45676 14900 45716
rect 15340 45676 15380 45716
rect 18124 45676 18164 45716
rect 18412 45676 18452 45716
rect 18892 45676 18932 45716
rect 19276 45676 19316 45716
rect 6700 45592 6740 45632
rect 6988 45592 7028 45632
rect 7180 45592 7220 45632
rect 4972 45508 5012 45548
rect 4492 45424 4532 45464
rect 4780 45424 4820 45464
rect 4928 45340 4968 45380
rect 5010 45340 5050 45380
rect 5092 45340 5132 45380
rect 5174 45340 5214 45380
rect 5256 45340 5296 45380
rect 4108 45172 4148 45212
rect 5452 45172 5492 45212
rect 5740 45172 5771 45212
rect 5771 45172 5780 45212
rect 3916 45088 3956 45128
rect 5356 45088 5396 45128
rect 5644 45088 5673 45128
rect 5673 45088 5684 45128
rect 76 44920 116 44960
rect 1612 44920 1652 44960
rect 4108 45004 4148 45044
rect 4492 44920 4532 44960
rect 4684 44920 4724 44960
rect 2572 44836 2612 44876
rect 76 44752 116 44792
rect 1420 44752 1460 44792
rect 2380 44752 2420 44792
rect 5452 45004 5492 45044
rect 7660 45424 7700 45464
rect 8332 45592 8372 45632
rect 6412 45340 6452 45380
rect 6892 45340 6932 45380
rect 7564 45340 7604 45380
rect 11500 45592 11540 45632
rect 13900 45592 13940 45632
rect 17260 45592 17300 45632
rect 15340 45508 15380 45548
rect 17740 45508 17780 45548
rect 14572 45424 14612 45464
rect 15244 45424 15284 45464
rect 6220 45256 6260 45296
rect 6700 45256 6740 45296
rect 7084 45256 7124 45296
rect 7948 45256 7988 45296
rect 6028 45172 6068 45212
rect 6892 45172 6932 45212
rect 9196 45172 9236 45212
rect 10444 45172 10484 45212
rect 11212 45172 11252 45212
rect 6316 45088 6356 45128
rect 6796 45088 6836 45128
rect 6988 45088 7028 45128
rect 7660 45088 7700 45128
rect 7948 45088 7988 45128
rect 8620 45088 8660 45128
rect 10348 45088 10388 45128
rect 5164 44836 5204 44876
rect 6028 45004 6068 45044
rect 6700 45004 6740 45044
rect 7468 45004 7508 45044
rect 7852 45004 7892 45044
rect 8140 45004 8180 45044
rect 8428 45004 8453 45044
rect 8453 45004 8468 45044
rect 10156 45004 10196 45044
rect 6892 44920 6932 44960
rect 7276 44920 7316 44960
rect 6700 44836 6740 44876
rect 7180 44836 7220 44876
rect 10828 45004 10859 45044
rect 10859 45004 10868 45044
rect 16492 45256 16532 45296
rect 15052 45172 15092 45212
rect 21004 45592 21044 45632
rect 21484 45592 21524 45632
rect 20524 45424 20564 45464
rect 20048 45340 20088 45380
rect 20130 45340 20170 45380
rect 20212 45340 20252 45380
rect 20294 45340 20334 45380
rect 20376 45340 20416 45380
rect 18412 45172 18452 45212
rect 18892 45172 18932 45212
rect 13420 45004 13460 45044
rect 13900 45004 13940 45044
rect 14476 45004 14516 45044
rect 15052 45035 15092 45044
rect 15052 45004 15092 45035
rect 17260 45035 17300 45044
rect 17260 45004 17300 45035
rect 8908 44920 8948 44960
rect 9292 44920 9332 44960
rect 10636 44920 10676 44960
rect 11500 44920 11540 44960
rect 13612 44920 13652 44960
rect 14188 44920 14228 44960
rect 14860 44920 14900 44960
rect 5932 44752 5972 44792
rect 6316 44752 6356 44792
rect 17644 45004 17684 45044
rect 18124 45004 18164 45044
rect 18412 45004 18452 45044
rect 18988 45004 19028 45044
rect 19276 45004 19316 45044
rect 20140 45004 20180 45044
rect 21292 44920 21332 44960
rect 19948 44836 19988 44876
rect 11212 44752 11252 44792
rect 12844 44752 12884 44792
rect 16204 44752 16244 44792
rect 10828 44668 10868 44708
rect 19564 44668 19604 44708
rect 3688 44584 3728 44624
rect 3770 44584 3810 44624
rect 3852 44584 3892 44624
rect 3934 44584 3974 44624
rect 4016 44584 4056 44624
rect 8716 44584 8756 44624
rect 11308 44584 11348 44624
rect 11500 44584 11540 44624
rect 18808 44584 18848 44624
rect 18890 44584 18930 44624
rect 18972 44584 19012 44624
rect 19054 44584 19094 44624
rect 19136 44584 19176 44624
rect 1612 44416 1652 44456
rect 4012 44416 4052 44456
rect 3916 44332 3956 44372
rect 76 44248 116 44288
rect 3052 44248 3092 44288
rect 4204 44248 4244 44288
rect 76 44080 116 44120
rect 2476 44164 2516 44204
rect 3340 44164 3380 44204
rect 3532 44164 3572 44204
rect 2668 44080 2708 44120
rect 3244 44080 3284 44120
rect 3436 43996 3476 44036
rect 6028 44500 6068 44540
rect 6700 44500 6740 44540
rect 9388 44500 9428 44540
rect 9868 44500 9908 44540
rect 14188 44500 14228 44540
rect 19276 44500 19316 44540
rect 5260 44416 5300 44456
rect 7276 44416 7316 44456
rect 13420 44416 13460 44456
rect 15052 44416 15092 44456
rect 17644 44416 17684 44456
rect 18028 44416 18068 44456
rect 20140 44416 20180 44456
rect 4492 44363 4532 44372
rect 4492 44332 4500 44363
rect 4500 44332 4532 44363
rect 5068 44332 5108 44372
rect 5740 44332 5780 44372
rect 6508 44332 6548 44372
rect 15916 44332 15956 44372
rect 16492 44332 16532 44372
rect 4876 44248 4916 44288
rect 5260 44248 5300 44288
rect 5932 44248 5972 44288
rect 6412 44248 6452 44288
rect 9772 44248 9803 44288
rect 9803 44248 9812 44288
rect 10348 44248 10388 44288
rect 10540 44248 10580 44288
rect 11308 44248 11348 44288
rect 11788 44248 11828 44288
rect 4684 44164 4724 44204
rect 18412 44248 18452 44288
rect 21004 44248 21044 44288
rect 6316 44164 6341 44204
rect 6341 44164 6356 44204
rect 5452 44080 5492 44120
rect 4684 43996 4724 44036
rect 5164 43996 5204 44036
rect 7564 44164 7604 44204
rect 8236 44164 8276 44204
rect 8908 44164 8948 44204
rect 9196 44164 9227 44204
rect 9227 44164 9236 44204
rect 9868 44164 9908 44204
rect 15052 44164 15092 44204
rect 15628 44164 15659 44204
rect 15659 44164 15668 44204
rect 16204 44164 16244 44204
rect 17740 44164 17780 44204
rect 17932 44164 17972 44204
rect 5932 44080 5972 44120
rect 1228 43744 1268 43784
rect 4928 43828 4968 43868
rect 5010 43828 5050 43868
rect 5092 43828 5132 43868
rect 5174 43828 5214 43868
rect 5256 43828 5296 43868
rect 5356 43828 5396 43868
rect 4492 43744 4532 43784
rect 2764 43660 2804 43700
rect 4204 43576 4244 43616
rect 3628 43492 3668 43532
rect 4108 43492 4148 43532
rect 6700 44080 6740 44120
rect 7948 44080 7988 44120
rect 9388 44080 9428 44120
rect 17644 44080 17684 44120
rect 7180 43996 7220 44036
rect 7468 43996 7508 44036
rect 8332 43996 8372 44036
rect 10252 43996 10292 44036
rect 6796 43828 6836 43868
rect 9868 43828 9908 43868
rect 14956 43996 14996 44036
rect 18316 43996 18356 44036
rect 14284 43828 14324 43868
rect 18124 43828 18164 43868
rect 20048 43828 20088 43868
rect 20130 43828 20170 43868
rect 20212 43828 20252 43868
rect 20294 43828 20334 43868
rect 20376 43828 20416 43868
rect 12844 43744 12884 43784
rect 8236 43660 8276 43700
rect 5260 43576 5300 43616
rect 5836 43576 5865 43616
rect 5865 43576 5876 43616
rect 6700 43576 6740 43616
rect 8716 43576 8756 43616
rect 8908 43576 8948 43616
rect 5740 43492 5780 43532
rect 6028 43492 6068 43532
rect 13228 43744 13268 43784
rect 12460 43660 12500 43700
rect 15052 43660 15092 43700
rect 12172 43576 12212 43616
rect 16780 43660 16820 43700
rect 19756 43660 19796 43700
rect 4012 43408 4052 43448
rect 2188 43324 2228 43364
rect 2092 43240 2132 43280
rect 3688 43072 3728 43112
rect 3770 43072 3810 43112
rect 3852 43072 3892 43112
rect 3934 43072 3974 43112
rect 4016 43072 4056 43112
rect 6988 43492 7028 43532
rect 6508 43408 6548 43448
rect 7756 43492 7796 43532
rect 7948 43492 7988 43532
rect 9292 43492 9332 43532
rect 10732 43492 10772 43532
rect 11020 43492 11060 43532
rect 11404 43492 11444 43532
rect 12364 43492 12404 43532
rect 14572 43492 14612 43532
rect 15052 43492 15092 43532
rect 15340 43492 15371 43532
rect 15371 43492 15380 43532
rect 17260 43492 17300 43532
rect 7084 43408 7124 43448
rect 11500 43408 11540 43448
rect 18124 43492 18164 43532
rect 18508 43492 18548 43532
rect 12844 43408 12884 43448
rect 13420 43408 13460 43448
rect 14476 43408 14516 43448
rect 15628 43408 15668 43448
rect 16300 43408 16340 43448
rect 19276 43492 19316 43532
rect 19564 43523 19604 43532
rect 19564 43492 19604 43523
rect 18604 43408 18644 43448
rect 20524 43408 20564 43448
rect 4972 43324 5012 43364
rect 5260 43324 5300 43364
rect 11404 43324 11444 43364
rect 13036 43324 13076 43364
rect 13708 43324 13748 43364
rect 14188 43324 14228 43364
rect 15340 43324 15380 43364
rect 16108 43324 16148 43364
rect 18700 43324 18740 43364
rect 4780 43240 4820 43280
rect 9868 43240 9908 43280
rect 11788 43240 11828 43280
rect 14380 43240 14420 43280
rect 11116 43156 11156 43196
rect 12844 43156 12884 43196
rect 15052 43156 15092 43196
rect 6316 42988 6356 43028
rect 11500 43072 11540 43112
rect 13324 43072 13364 43112
rect 15436 43072 15476 43112
rect 18808 43072 18848 43112
rect 18890 43072 18930 43112
rect 18972 43072 19012 43112
rect 19054 43072 19094 43112
rect 19136 43072 19176 43112
rect 4684 42904 4724 42944
rect 4972 42904 5012 42944
rect 5932 42904 5972 42944
rect 6124 42904 6164 42944
rect 9772 42904 9812 42944
rect 11980 42904 12020 42944
rect 15628 42904 15668 42944
rect 1036 42820 1076 42860
rect 5164 42820 5204 42860
rect 6028 42820 6068 42860
rect 4108 42736 4148 42776
rect 6508 42736 6548 42776
rect 3148 42652 3188 42692
rect 4684 42652 4724 42692
rect 5356 42652 5385 42692
rect 5385 42652 5396 42692
rect 5644 42652 5684 42692
rect 6124 42652 6164 42692
rect 6412 42652 6452 42692
rect 1804 42568 1844 42608
rect 1708 42484 1748 42524
rect 5260 42568 5300 42608
rect 6028 42568 6068 42608
rect 6892 42568 6932 42608
rect 2476 42484 2516 42524
rect 4684 42484 4724 42524
rect 6988 42484 7028 42524
rect 6892 42400 6932 42440
rect 8236 42736 8276 42776
rect 12652 42736 12692 42776
rect 13804 42736 13844 42776
rect 15436 42736 15476 42776
rect 18508 42736 18548 42776
rect 20524 42736 20564 42776
rect 7948 42652 7988 42692
rect 8332 42652 8372 42692
rect 9868 42652 9908 42692
rect 11212 42652 11252 42692
rect 13324 42652 13355 42692
rect 13355 42652 13364 42692
rect 14188 42652 14228 42692
rect 15244 42652 15284 42692
rect 15628 42652 15668 42692
rect 16300 42652 16340 42692
rect 13804 42568 13844 42608
rect 4780 42316 4820 42356
rect 4928 42316 4968 42356
rect 5010 42316 5050 42356
rect 5092 42316 5132 42356
rect 5174 42316 5214 42356
rect 5256 42316 5296 42356
rect 14284 42484 14324 42524
rect 15052 42484 15092 42524
rect 7372 42232 7412 42272
rect 2956 42148 2996 42188
rect 3628 42148 3668 42188
rect 7948 42148 7988 42188
rect 10444 42148 10484 42188
rect 10732 42148 10772 42188
rect 3532 42064 3572 42104
rect 11212 42400 11252 42440
rect 12940 42400 12980 42440
rect 15820 42484 15860 42524
rect 14476 42400 14516 42440
rect 13036 42232 13076 42272
rect 13420 42148 13460 42188
rect 11788 42064 11828 42104
rect 13036 42064 13076 42104
rect 15436 42064 15476 42104
rect 18124 42652 18164 42692
rect 18604 42652 18644 42692
rect 19276 42652 19316 42692
rect 20812 42652 20852 42692
rect 17836 42484 17876 42524
rect 16204 42232 16244 42272
rect 20048 42316 20088 42356
rect 20130 42316 20170 42356
rect 20212 42316 20252 42356
rect 20294 42316 20334 42356
rect 20376 42316 20416 42356
rect 20620 42232 20660 42272
rect 15628 42148 15668 42188
rect 19564 42148 19604 42188
rect 20524 42148 20564 42188
rect 2476 41980 2516 42020
rect 2860 41980 2900 42020
rect 4588 41980 4628 42020
rect 6220 41980 6260 42020
rect 3148 41896 3188 41936
rect 5356 41896 5396 41936
rect 5644 41896 5684 41936
rect 5932 41896 5972 41936
rect 8428 41980 8468 42020
rect 8716 41980 8756 42020
rect 9868 41980 9908 42020
rect 10636 41980 10676 42020
rect 12460 41980 12500 42020
rect 13708 41980 13748 42020
rect 14188 41980 14228 42020
rect 7948 41896 7988 41936
rect 9772 41896 9812 41936
rect 11596 41896 11636 41936
rect 15052 41980 15092 42020
rect 16108 42064 16148 42104
rect 15820 41980 15845 42020
rect 15845 41980 15860 42020
rect 15436 41896 15476 41936
rect 16684 41980 16724 42020
rect 17836 42011 17876 42020
rect 17836 41980 17876 42011
rect 18412 41980 18452 42020
rect 18700 41980 18740 42020
rect 21388 41896 21428 41936
rect 4108 41812 4148 41852
rect 4780 41812 4820 41852
rect 5836 41812 5876 41852
rect 6796 41812 6836 41852
rect 7180 41812 7220 41852
rect 7852 41812 7892 41852
rect 11500 41812 11540 41852
rect 12268 41812 12308 41852
rect 13804 41812 13844 41852
rect 15820 41812 15860 41852
rect 16300 41812 16340 41852
rect 16684 41812 16724 41852
rect 172 41728 212 41768
rect 1900 41728 1940 41768
rect 14188 41728 14228 41768
rect 18412 41728 18452 41768
rect 7852 41644 7892 41684
rect 13804 41644 13844 41684
rect 16108 41644 16148 41684
rect 16492 41644 16532 41684
rect 18508 41644 18548 41684
rect 3688 41560 3728 41600
rect 3770 41560 3810 41600
rect 3852 41560 3892 41600
rect 3934 41560 3974 41600
rect 4016 41560 4056 41600
rect 7180 41560 7220 41600
rect 8044 41560 8084 41600
rect 13996 41560 14036 41600
rect 15628 41560 15668 41600
rect 17836 41560 17876 41600
rect 18808 41560 18848 41600
rect 18890 41560 18930 41600
rect 18972 41560 19012 41600
rect 19054 41560 19094 41600
rect 19136 41560 19176 41600
rect 21004 41560 21044 41600
rect 1612 41392 1652 41432
rect 2668 41392 2708 41432
rect 4108 41392 4148 41432
rect 4588 41392 4628 41432
rect 6508 41392 6548 41432
rect 9484 41392 9524 41432
rect 12460 41392 12500 41432
rect 14188 41392 14228 41432
rect 16204 41392 16244 41432
rect 16492 41392 16532 41432
rect 18028 41392 18068 41432
rect 21100 41476 21140 41516
rect 1516 41308 1556 41348
rect 4492 41224 4532 41264
rect 5356 41224 5396 41264
rect 6508 41224 6548 41264
rect 11308 41224 11348 41264
rect 12460 41224 12500 41264
rect 13324 41308 13364 41348
rect 15244 41308 15284 41348
rect 16012 41308 16052 41348
rect 18700 41308 18740 41348
rect 14572 41224 14612 41264
rect 15820 41224 15860 41264
rect 18988 41224 19028 41264
rect 460 41140 500 41180
rect 1228 41140 1268 41180
rect 2476 41140 2516 41180
rect 2668 41140 2708 41180
rect 3052 41140 3092 41180
rect 4108 41140 4148 41180
rect 5164 41140 5204 41180
rect 6028 41140 6059 41180
rect 6059 41140 6068 41180
rect 6796 41140 6836 41180
rect 7180 41140 7220 41180
rect 7468 41140 7508 41180
rect 8716 41140 8756 41180
rect 10156 41140 10196 41180
rect 10636 41140 10676 41180
rect 76 41056 116 41096
rect 5260 41056 5300 41096
rect 4012 40972 4052 41012
rect 5356 40972 5387 41012
rect 5387 40972 5396 41012
rect 11500 41140 11540 41180
rect 12364 41140 12372 41180
rect 12372 41140 12404 41180
rect 13708 41140 13748 41180
rect 15436 41140 15476 41180
rect 15916 41140 15956 41180
rect 16108 41140 16148 41180
rect 6124 41056 6164 41096
rect 6604 41056 6644 41096
rect 10732 41056 10772 41096
rect 10924 41056 10964 41096
rect 14188 41056 14228 41096
rect 15244 41056 15284 41096
rect 5932 40972 5972 41012
rect 6220 40972 6260 41012
rect 6508 40972 6548 41012
rect 7180 40972 7220 41012
rect 12652 40972 12692 41012
rect 13804 40972 13844 41012
rect 15436 40972 15476 41012
rect 16204 40972 16244 41012
rect 17740 41140 17780 41180
rect 18220 41140 18260 41180
rect 18508 41140 18548 41180
rect 18892 41140 18932 41180
rect 17644 41056 17684 41096
rect 1420 40888 1460 40928
rect 4108 40888 4148 40928
rect 6604 40888 6644 40928
rect 7468 40888 7508 40928
rect 16492 40888 16532 40928
rect 1228 40720 1268 40760
rect 1900 40636 1940 40676
rect 2284 40636 2324 40676
rect 76 40552 116 40592
rect 1516 40552 1556 40592
rect 2668 40552 2708 40592
rect 2284 40468 2324 40508
rect 2572 40468 2612 40508
rect 172 40384 212 40424
rect 1612 40384 1652 40424
rect 2668 40384 2708 40424
rect 4928 40804 4968 40844
rect 5010 40804 5050 40844
rect 5092 40804 5132 40844
rect 5174 40804 5214 40844
rect 5256 40804 5296 40844
rect 6028 40804 6068 40844
rect 12940 40804 12980 40844
rect 16012 40804 16052 40844
rect 6796 40720 6836 40760
rect 8716 40720 8756 40760
rect 9964 40720 10004 40760
rect 13420 40720 13460 40760
rect 15436 40720 15476 40760
rect 4492 40636 4532 40676
rect 4972 40636 5012 40676
rect 6220 40636 6260 40676
rect 7180 40636 7220 40676
rect 6124 40552 6164 40592
rect 7084 40552 7124 40592
rect 9484 40636 9524 40676
rect 7756 40552 7787 40592
rect 7787 40552 7796 40592
rect 3148 40468 3188 40508
rect 3340 40468 3380 40508
rect 4012 40468 4052 40508
rect 5164 40468 5204 40508
rect 6028 40468 6068 40508
rect 5260 40384 5300 40424
rect 1420 40300 1460 40340
rect 1708 40300 1748 40340
rect 2476 40300 2516 40340
rect 4876 40300 4916 40340
rect 5644 40300 5684 40340
rect 6220 40468 6260 40508
rect 7660 40468 7698 40484
rect 7698 40468 7700 40484
rect 7660 40444 7700 40468
rect 12364 40636 12404 40676
rect 13612 40636 13652 40676
rect 15628 40636 15668 40676
rect 14572 40552 14612 40592
rect 9772 40468 9812 40508
rect 10252 40468 10292 40508
rect 10828 40468 10868 40508
rect 20524 41392 20564 41432
rect 20620 41308 20660 41348
rect 20044 41140 20084 41180
rect 17836 40972 17876 41012
rect 20048 40804 20088 40844
rect 20130 40804 20170 40844
rect 20212 40804 20252 40844
rect 20294 40804 20334 40844
rect 20376 40804 20416 40844
rect 18412 40636 18452 40676
rect 20044 40636 20084 40676
rect 21100 40636 21140 40676
rect 21292 40552 21332 40592
rect 13324 40468 13364 40508
rect 13804 40468 13844 40508
rect 6316 40384 6356 40424
rect 7372 40384 7412 40424
rect 8044 40384 8084 40424
rect 8620 40384 8660 40424
rect 9004 40384 9044 40424
rect 9484 40384 9524 40424
rect 13132 40384 13172 40424
rect 12844 40300 12884 40340
rect 2956 40216 2996 40256
rect 6316 40216 6356 40256
rect 8908 40216 8948 40256
rect 1900 40132 1940 40172
rect 9964 40132 10004 40172
rect 14668 40468 14708 40508
rect 15628 40468 15668 40508
rect 16492 40468 16532 40508
rect 16876 40468 16916 40508
rect 17548 40468 17588 40508
rect 17836 40468 17876 40508
rect 19276 40468 19316 40508
rect 19564 40468 19604 40508
rect 20140 40499 20180 40508
rect 20140 40468 20180 40499
rect 14188 40384 14228 40424
rect 15436 40384 15476 40424
rect 15820 40384 15860 40424
rect 18124 40384 18164 40424
rect 18604 40384 18644 40424
rect 18988 40384 19028 40424
rect 14092 40300 14132 40340
rect 19852 40300 19892 40340
rect 14092 40132 14132 40172
rect 364 40048 404 40088
rect 3688 40048 3728 40088
rect 3770 40048 3810 40088
rect 3852 40048 3892 40088
rect 3934 40048 3974 40088
rect 4016 40048 4056 40088
rect 8620 40048 8660 40088
rect 8812 40048 8852 40088
rect 16492 40048 16532 40088
rect 18808 40048 18848 40088
rect 18890 40048 18930 40088
rect 18972 40048 19012 40088
rect 19054 40048 19094 40088
rect 19136 40048 19176 40088
rect 11980 39964 12020 40004
rect 12556 39964 12596 40004
rect 1900 39880 1940 39920
rect 6124 39880 6164 39920
rect 6412 39880 6443 39920
rect 6443 39880 6452 39920
rect 8428 39880 8468 39920
rect 12364 39880 12404 39920
rect 13900 39880 13940 39920
rect 2860 39796 2900 39836
rect 5164 39796 5204 39836
rect 5836 39796 5876 39836
rect 9772 39796 9812 39836
rect 10060 39796 10100 39836
rect 11020 39796 11060 39836
rect 1228 39712 1268 39752
rect 1420 39712 1460 39752
rect 2668 39712 2708 39752
rect 3148 39712 3188 39752
rect 4396 39712 4436 39752
rect 4780 39712 4820 39752
rect 1612 39628 1652 39668
rect 5356 39712 5396 39752
rect 6604 39712 6644 39752
rect 10348 39712 10388 39752
rect 10924 39712 10964 39752
rect 12940 39712 12980 39752
rect 13516 39712 13556 39752
rect 1804 39628 1844 39668
rect 2956 39628 2996 39668
rect 1708 39544 1748 39584
rect 1900 39544 1940 39584
rect 2668 39544 2708 39584
rect 940 39460 980 39500
rect 3148 39460 3188 39500
rect 1228 39040 1268 39080
rect 3724 39124 3764 39164
rect 4492 39628 4532 39668
rect 5932 39628 5953 39668
rect 5953 39628 5972 39668
rect 6316 39628 6356 39668
rect 4204 39460 4244 39500
rect 4876 39460 4916 39500
rect 5164 39460 5204 39500
rect 4928 39292 4968 39332
rect 5010 39292 5050 39332
rect 5092 39292 5132 39332
rect 5174 39292 5214 39332
rect 5256 39292 5296 39332
rect 14092 39796 14132 39836
rect 7084 39628 7124 39668
rect 7852 39628 7892 39668
rect 8236 39628 8276 39668
rect 9484 39628 9524 39668
rect 10828 39628 10868 39668
rect 6028 39544 6068 39584
rect 6220 39544 6260 39584
rect 6412 39544 6441 39584
rect 6441 39544 6452 39584
rect 5836 39460 5876 39500
rect 6988 39460 7028 39500
rect 12268 39628 12308 39650
rect 12268 39610 12308 39628
rect 12556 39628 12596 39668
rect 13420 39628 13460 39668
rect 17740 39880 17780 39920
rect 19948 39880 19988 39920
rect 20140 39880 20180 39920
rect 14476 39796 14516 39836
rect 20044 39796 20084 39836
rect 12652 39544 12692 39584
rect 13036 39544 13076 39584
rect 14668 39544 14708 39584
rect 9292 39460 9332 39500
rect 10636 39460 10676 39500
rect 13132 39460 13172 39500
rect 15820 39712 15860 39752
rect 18124 39712 18164 39752
rect 18508 39712 18548 39752
rect 17548 39628 17588 39668
rect 18892 39628 18932 39668
rect 6700 39376 6740 39416
rect 9484 39376 9524 39416
rect 10060 39376 10100 39416
rect 11500 39376 11540 39416
rect 8524 39292 8564 39332
rect 10924 39292 10964 39332
rect 13228 39292 13268 39332
rect 6988 39208 7028 39248
rect 8620 39208 8660 39248
rect 8812 39208 8852 39248
rect 13036 39208 13076 39248
rect 13420 39208 13460 39248
rect 4876 39124 4916 39164
rect 5548 39124 5588 39164
rect 6028 39124 6068 39164
rect 8908 39124 8948 39164
rect 9292 39124 9332 39164
rect 12652 39124 12692 39164
rect 6220 39040 6260 39080
rect 6796 39040 6836 39080
rect 8332 39040 8372 39080
rect 11116 39040 11156 39080
rect 2476 38956 2516 38996
rect 4012 38956 4052 38996
rect 4300 38956 4340 38996
rect 4684 38956 4724 38996
rect 5452 38956 5492 38996
rect 5740 38987 5780 38996
rect 5740 38956 5780 38987
rect 6124 38956 6164 38996
rect 6988 38956 7028 38996
rect 7276 38956 7316 38996
rect 364 38872 404 38912
rect 1612 38872 1652 38912
rect 4204 38872 4244 38912
rect 4780 38872 4820 38912
rect 6700 38872 6740 38912
rect 6892 38872 6932 38912
rect 7180 38872 7220 38912
rect 8812 38956 8852 38996
rect 17644 39544 17684 39584
rect 21292 39460 21332 39500
rect 20048 39292 20088 39332
rect 20130 39292 20170 39332
rect 20212 39292 20252 39332
rect 20294 39292 20334 39332
rect 20376 39292 20416 39332
rect 20620 39208 20660 39248
rect 14188 39124 14228 39164
rect 18508 39124 18548 39164
rect 21004 39040 21044 39080
rect 10924 38956 10964 38996
rect 11884 38956 11924 38996
rect 13228 38956 13268 38996
rect 13516 38956 13547 38996
rect 13547 38956 13556 38996
rect 13708 38956 13748 38996
rect 15820 38956 15860 38996
rect 16876 38956 16916 38996
rect 18028 38956 18068 38996
rect 8428 38788 8468 38828
rect 10636 38872 10676 38912
rect 10828 38872 10868 38912
rect 11116 38872 11156 38912
rect 12460 38872 12500 38912
rect 13036 38872 13076 38912
rect 13996 38872 14036 38912
rect 16300 38872 16340 38912
rect 18508 38872 18548 38912
rect 11020 38788 11060 38828
rect 15436 38788 15476 38828
rect 18124 38788 18164 38828
rect 1612 38704 1652 38744
rect 1900 38704 1940 38744
rect 10444 38704 10484 38744
rect 16012 38704 16052 38744
rect 18412 38704 18452 38744
rect 19948 38704 19988 38744
rect 3688 38536 3728 38576
rect 3770 38536 3810 38576
rect 3852 38536 3892 38576
rect 3934 38536 3974 38576
rect 4016 38536 4056 38576
rect 3532 38452 3572 38492
rect 2572 38368 2612 38408
rect 2764 38284 2804 38324
rect 3052 38200 3092 38240
rect 4300 38368 4340 38408
rect 12652 38620 12692 38660
rect 19852 38620 19892 38660
rect 5452 38536 5492 38576
rect 16780 38536 16820 38576
rect 18808 38536 18848 38576
rect 18890 38536 18930 38576
rect 18972 38536 19012 38576
rect 19054 38536 19094 38576
rect 19136 38536 19176 38576
rect 6700 38452 6740 38492
rect 11596 38452 11636 38492
rect 12268 38452 12308 38492
rect 12748 38452 12788 38492
rect 12460 38368 12500 38408
rect 14668 38368 14708 38408
rect 15724 38368 15764 38408
rect 18508 38368 18548 38408
rect 5836 38284 5876 38324
rect 6124 38284 6164 38324
rect 6508 38284 6548 38324
rect 8620 38284 8660 38324
rect 9964 38284 10004 38324
rect 12172 38284 12212 38324
rect 13228 38284 13268 38324
rect 4300 38200 4340 38240
rect 5548 38200 5588 38240
rect 5932 38200 5972 38240
rect 7756 38200 7796 38240
rect 8428 38200 8468 38240
rect 9196 38200 9236 38240
rect 9484 38200 9524 38240
rect 12844 38200 12884 38240
rect 15052 38200 15092 38240
rect 15436 38200 15476 38240
rect 16012 38200 16052 38240
rect 16876 38200 16916 38240
rect 18412 38284 18452 38324
rect 19276 38200 19316 38240
rect 19660 38200 19700 38240
rect 1324 38116 1364 38156
rect 4108 38116 4148 38156
rect 748 38032 788 38072
rect 5836 38032 5876 38072
rect 6124 38032 6164 38072
rect 6316 38032 6356 38072
rect 5452 37948 5492 37988
rect 7372 38116 7412 38156
rect 11884 38116 11924 38156
rect 12172 38116 12212 38156
rect 12748 38116 12788 38156
rect 13804 38116 13844 38156
rect 2860 37864 2900 37904
rect 6892 38032 6932 38072
rect 7084 38032 7124 38072
rect 10828 38032 10868 38072
rect 11596 38032 11636 38072
rect 13516 38032 13556 38072
rect 19084 38116 19124 38156
rect 20524 38116 20564 38156
rect 15436 38032 15476 38072
rect 15820 38032 15860 38072
rect 16492 38032 16532 38072
rect 18412 38032 18452 38072
rect 18604 38032 18644 38072
rect 6796 37948 6827 37988
rect 6827 37948 6836 37988
rect 7372 37948 7412 37988
rect 8620 37948 8660 37988
rect 10540 37948 10580 37988
rect 12748 37948 12788 37988
rect 14860 37948 14900 37988
rect 15244 37948 15284 37988
rect 11500 37864 11540 37904
rect 12268 37864 12308 37904
rect 4928 37780 4968 37820
rect 5010 37780 5050 37820
rect 5092 37780 5132 37820
rect 5174 37780 5214 37820
rect 5256 37780 5296 37820
rect 9484 37780 9524 37820
rect 10540 37780 10580 37820
rect 11596 37780 11636 37820
rect 12844 37780 12884 37820
rect 844 37696 884 37736
rect 12556 37696 12596 37736
rect 2092 37612 2132 37652
rect 5452 37612 5492 37652
rect 5836 37612 5876 37652
rect 12172 37612 12212 37652
rect 13132 37612 13172 37652
rect 13420 37612 13460 37652
rect 3436 37528 3476 37568
rect 8044 37528 8084 37568
rect 10060 37528 10100 37568
rect 11884 37528 11924 37568
rect 12844 37528 12884 37568
rect 1708 37444 1748 37484
rect 2860 37444 2900 37484
rect 3820 37444 3860 37484
rect 4780 37444 4820 37484
rect 5932 37444 5972 37484
rect 6124 37444 6164 37484
rect 6700 37444 6740 37484
rect 7660 37444 7700 37484
rect 9964 37444 10004 37484
rect 10540 37444 10580 37484
rect 11500 37444 11540 37484
rect 13324 37528 13364 37568
rect 17836 37528 17876 37568
rect 20908 37948 20948 37988
rect 20048 37780 20088 37820
rect 20130 37780 20170 37820
rect 20212 37780 20252 37820
rect 20294 37780 20334 37820
rect 20376 37780 20416 37820
rect 21004 37696 21044 37736
rect 18412 37528 18452 37568
rect 18892 37528 18932 37568
rect 2764 37360 2804 37400
rect 2668 37276 2708 37316
rect 3340 37192 3380 37232
rect 12652 37444 12659 37484
rect 12659 37444 12692 37484
rect 13516 37444 13556 37484
rect 13804 37444 13844 37484
rect 15052 37475 15092 37484
rect 15052 37444 15092 37475
rect 15244 37444 15284 37484
rect 16588 37444 16628 37484
rect 19276 37444 19316 37484
rect 19948 37444 19988 37484
rect 7756 37360 7796 37400
rect 8620 37360 8660 37400
rect 12748 37360 12779 37400
rect 12779 37360 12788 37400
rect 13612 37360 13652 37400
rect 16876 37360 16916 37400
rect 17356 37360 17396 37400
rect 17644 37360 17684 37400
rect 18124 37360 18164 37400
rect 18604 37360 18644 37400
rect 19084 37360 19124 37400
rect 7276 37276 7316 37316
rect 8812 37276 8852 37316
rect 10348 37276 10388 37316
rect 4108 37192 4148 37232
rect 6316 37192 6356 37232
rect 17164 37276 17204 37316
rect 17548 37276 17588 37316
rect 8236 37192 8276 37232
rect 14860 37192 14900 37232
rect 17260 37192 17300 37232
rect 18124 37192 18164 37232
rect 21292 37192 21332 37232
rect 3688 37024 3728 37064
rect 3770 37024 3810 37064
rect 3852 37024 3892 37064
rect 3934 37024 3974 37064
rect 4016 37024 4056 37064
rect 5452 36940 5492 36980
rect 7948 36856 7988 36896
rect 3052 36772 3092 36812
rect 6796 36772 6836 36812
rect 652 36688 692 36728
rect 1228 36688 1268 36728
rect 1612 36688 1652 36728
rect 2572 36688 2612 36728
rect 3628 36688 3668 36728
rect 8236 36688 8267 36728
rect 8267 36688 8276 36728
rect 18220 37108 18260 37148
rect 19948 37108 19988 37148
rect 18808 37024 18848 37064
rect 18890 37024 18930 37064
rect 18972 37024 19012 37064
rect 19054 37024 19094 37064
rect 19136 37024 19176 37064
rect 14860 36772 14900 36812
rect 9484 36688 9524 36728
rect 11788 36688 11828 36728
rect 13708 36688 13748 36728
rect 2380 36604 2420 36644
rect 1420 36352 1460 36392
rect 3532 36604 3572 36644
rect 6124 36604 6164 36644
rect 6700 36604 6740 36644
rect 7756 36604 7796 36644
rect 9292 36604 9332 36644
rect 9964 36604 10004 36644
rect 3820 36520 3860 36560
rect 4684 36520 4724 36560
rect 9100 36520 9140 36560
rect 6124 36436 6164 36476
rect 7660 36436 7700 36476
rect 8428 36436 8459 36476
rect 8459 36436 8468 36476
rect 10444 36604 10484 36644
rect 10924 36604 10964 36644
rect 11692 36604 11732 36644
rect 11884 36604 11924 36644
rect 12268 36604 12308 36644
rect 13612 36604 13652 36644
rect 13804 36604 13844 36644
rect 15724 36940 15764 36980
rect 15820 36856 15860 36896
rect 20524 36856 20564 36896
rect 17548 36772 17588 36812
rect 14668 36604 14708 36644
rect 6988 36352 7028 36392
rect 7276 36352 7316 36392
rect 14956 36520 14996 36560
rect 12076 36436 12116 36476
rect 12940 36436 12980 36476
rect 15244 36436 15284 36476
rect 18604 36688 18644 36728
rect 15916 36604 15956 36644
rect 16300 36604 16340 36644
rect 17260 36604 17300 36644
rect 17740 36604 17780 36644
rect 18220 36604 18260 36644
rect 18892 36604 18932 36644
rect 17164 36520 17204 36560
rect 17548 36520 17588 36560
rect 12844 36352 12884 36392
rect 4928 36268 4968 36308
rect 5010 36268 5050 36308
rect 5092 36268 5132 36308
rect 5174 36268 5214 36308
rect 5256 36268 5296 36308
rect 8812 36268 8852 36308
rect 17836 36268 17876 36308
rect 4492 36184 4532 36224
rect 5644 36184 5684 36224
rect 10540 36184 10580 36224
rect 10924 36184 10964 36224
rect 13996 36184 14036 36224
rect 14860 36184 14900 36224
rect 16588 36184 16628 36224
rect 3052 36100 3092 36140
rect 3340 36100 3380 36140
rect 4012 36100 4052 36140
rect 6700 36100 6740 36140
rect 12268 36100 12308 36140
rect 13612 36100 13652 36140
rect 1228 36016 1268 36056
rect 1708 36016 1748 36056
rect 4108 36016 4148 36056
rect 4588 36016 4628 36056
rect 7276 36016 7316 36056
rect 7756 36016 7796 36056
rect 844 35932 884 35972
rect 2188 35932 2228 35972
rect 2764 35932 2804 35972
rect 3436 35932 3476 35972
rect 4492 35932 4532 35972
rect 6316 35932 6347 35972
rect 6347 35932 6356 35972
rect 11500 36016 11540 36056
rect 13420 36016 13460 36056
rect 8236 35932 8276 35972
rect 9772 35963 9812 35972
rect 9772 35932 9812 35963
rect 11116 35932 11156 35972
rect 11788 35932 11828 35972
rect 12748 35932 12777 35972
rect 12777 35932 12788 35972
rect 13324 35932 13364 35972
rect 748 35848 788 35888
rect 2284 35848 2324 35888
rect 3628 35848 3668 35888
rect 6124 35848 6164 35888
rect 6796 35848 6836 35888
rect 11980 35848 12020 35888
rect 3340 35764 3380 35804
rect 3820 35764 3860 35804
rect 5740 35764 5780 35804
rect 844 35680 884 35720
rect 2380 35680 2420 35720
rect 8044 35764 8084 35804
rect 10924 35680 10964 35720
rect 9004 35596 9044 35636
rect 12940 35848 12980 35888
rect 15724 36100 15764 36140
rect 17644 36100 17684 36140
rect 15244 36016 15284 36056
rect 16300 36016 16340 36056
rect 15436 35932 15476 35972
rect 15820 35932 15860 35972
rect 14572 35764 14612 35804
rect 14860 35764 14900 35804
rect 12556 35680 12596 35720
rect 3688 35512 3728 35552
rect 3770 35512 3810 35552
rect 3852 35512 3892 35552
rect 3934 35512 3974 35552
rect 4016 35512 4056 35552
rect 5164 35512 5204 35552
rect 7276 35512 7316 35552
rect 4492 35428 4532 35468
rect 6796 35428 6836 35468
rect 172 35344 212 35384
rect 3532 35344 3572 35384
rect 4204 35344 4244 35384
rect 6604 35344 6644 35384
rect 9292 35344 9332 35384
rect 11404 35344 11444 35384
rect 13324 35344 13364 35384
rect 2380 35260 2420 35300
rect 652 35176 692 35216
rect 1420 35176 1460 35216
rect 9484 35260 9524 35300
rect 12556 35260 12596 35300
rect 2092 35092 2132 35132
rect 1324 35008 1364 35048
rect 2380 35008 2420 35048
rect 4012 35092 4052 35132
rect 5164 35092 5204 35132
rect 5836 35092 5876 35132
rect 2956 35008 2996 35048
rect 5356 35008 5396 35048
rect 7756 35176 7796 35216
rect 17548 35932 17588 35972
rect 18124 36352 18164 36392
rect 20048 36268 20088 36308
rect 20130 36268 20170 36308
rect 20212 36268 20252 36308
rect 20294 36268 20334 36308
rect 20376 36268 20416 36308
rect 20908 36184 20948 36224
rect 20044 36100 20084 36140
rect 18412 36016 18452 36056
rect 19180 36016 19220 36056
rect 19276 35932 19316 35972
rect 16780 35848 16820 35888
rect 20812 35932 20852 35972
rect 18700 35848 18740 35888
rect 19084 35848 19124 35888
rect 16300 35764 16340 35804
rect 17260 35764 17300 35804
rect 18028 35764 18068 35804
rect 15916 35596 15956 35636
rect 14860 35512 14900 35552
rect 18808 35512 18848 35552
rect 18890 35512 18930 35552
rect 18972 35512 19012 35552
rect 19054 35512 19094 35552
rect 19136 35512 19176 35552
rect 16300 35428 16340 35468
rect 14764 35344 14804 35384
rect 15244 35344 15284 35384
rect 14380 35176 14420 35216
rect 7180 35092 7220 35132
rect 7468 35092 7492 35132
rect 7492 35092 7508 35132
rect 8044 35092 8081 35132
rect 8081 35092 8084 35132
rect 9772 35092 9812 35132
rect 10348 35092 10388 35132
rect 13036 35092 13076 35132
rect 14764 35092 14804 35132
rect 21100 35680 21140 35720
rect 18220 35344 18260 35384
rect 16684 35260 16724 35300
rect 17644 35260 17684 35300
rect 19564 35260 19604 35300
rect 21100 35260 21140 35300
rect 16300 35176 16340 35216
rect 17260 35176 17300 35216
rect 17836 35176 17876 35216
rect 20524 35176 20564 35216
rect 16588 35092 16628 35132
rect 16780 35092 16820 35132
rect 18028 35092 18068 35132
rect 18892 35092 18932 35132
rect 7948 35008 7988 35048
rect 8236 35008 8276 35048
rect 13324 35008 13364 35048
rect 14284 35008 14324 35048
rect 14668 35008 14708 35048
rect 15916 35008 15956 35048
rect 16684 35008 16724 35048
rect 18220 35008 18260 35048
rect 6124 34924 6164 34964
rect 7852 34924 7892 34964
rect 9100 34924 9140 34964
rect 13420 34924 13460 34964
rect 15628 34924 15668 34964
rect 17452 34924 17492 34964
rect 2764 34840 2804 34880
rect 6316 34840 6356 34880
rect 8908 34840 8948 34880
rect 12556 34840 12596 34880
rect 13324 34840 13364 34880
rect 14956 34840 14996 34880
rect 17836 34924 17876 34964
rect 18124 34924 18164 34964
rect 20044 34924 20084 34964
rect 18316 34840 18356 34880
rect 4928 34756 4968 34796
rect 5010 34756 5050 34796
rect 5092 34756 5132 34796
rect 5174 34756 5214 34796
rect 5256 34756 5296 34796
rect 6700 34756 6740 34796
rect 15244 34756 15284 34796
rect 15628 34756 15668 34796
rect 1612 34672 1652 34712
rect 5836 34672 5876 34712
rect 2668 34588 2708 34628
rect 9196 34588 9236 34628
rect 12076 34588 12116 34628
rect 20048 34756 20088 34796
rect 20130 34756 20170 34796
rect 20212 34756 20252 34796
rect 20294 34756 20334 34796
rect 20376 34756 20416 34796
rect 21004 34672 21044 34712
rect 20044 34588 20084 34628
rect 5740 34504 5780 34544
rect 8812 34504 8852 34544
rect 10348 34504 10388 34544
rect 11116 34504 11155 34544
rect 11155 34504 11156 34544
rect 11596 34504 11636 34544
rect 12460 34504 12500 34544
rect 12940 34504 12980 34544
rect 14284 34504 14324 34544
rect 14764 34504 14804 34544
rect 14956 34504 14996 34544
rect 17452 34504 17463 34544
rect 17463 34504 17492 34544
rect 18700 34504 18740 34544
rect 19660 34504 19700 34544
rect 19852 34504 19892 34544
rect 20620 34504 20660 34544
rect 844 34420 884 34460
rect 2284 34420 2315 34460
rect 2315 34420 2324 34460
rect 2668 34420 2708 34460
rect 3532 34420 3572 34460
rect 460 34336 500 34376
rect 1228 34336 1268 34376
rect 2476 34336 2516 34376
rect 2956 34336 2996 34376
rect 4396 34451 4436 34460
rect 4396 34420 4436 34451
rect 5260 34420 5300 34460
rect 7276 34451 7316 34460
rect 7276 34420 7316 34451
rect 7564 34420 7604 34460
rect 8908 34451 8948 34460
rect 8908 34420 8948 34451
rect 9580 34420 9620 34460
rect 10060 34420 10100 34460
rect 10444 34451 10484 34460
rect 10444 34420 10484 34451
rect 10924 34451 10964 34460
rect 10924 34420 10964 34451
rect 11980 34420 12020 34460
rect 4972 34336 5012 34376
rect 5932 34336 5972 34376
rect 2092 34252 2132 34292
rect 15244 34420 15284 34460
rect 10252 34336 10292 34376
rect 12076 34336 12116 34376
rect 12556 34336 12596 34376
rect 4780 34252 4820 34292
rect 5740 34252 5780 34292
rect 16012 34420 16052 34460
rect 14380 34336 14420 34376
rect 14860 34336 14900 34376
rect 15436 34252 15476 34292
rect 1996 34168 2036 34208
rect 3340 34168 3380 34208
rect 7468 34168 7508 34208
rect 4300 34084 4340 34124
rect 5932 34084 5972 34124
rect 1612 34000 1652 34040
rect 3688 34000 3728 34040
rect 3770 34000 3810 34040
rect 3852 34000 3892 34040
rect 3934 34000 3974 34040
rect 4016 34000 4056 34040
rect 4780 34000 4820 34040
rect 6604 34000 6644 34040
rect 6220 33916 6260 33956
rect 8428 33916 8468 33956
rect 2572 33832 2612 33872
rect 6412 33832 6452 33872
rect 7756 33832 7796 33872
rect 1324 33748 1364 33788
rect 6220 33748 6260 33788
rect 1996 33664 2036 33704
rect 3532 33664 3572 33704
rect 1132 33580 1172 33620
rect 2764 33580 2804 33620
rect 6796 33580 6836 33620
rect 7276 33580 7316 33620
rect 8812 33580 8852 33620
rect 2668 33496 2708 33536
rect 3052 33496 3092 33536
rect 15916 34336 15956 34376
rect 17932 34420 17972 34460
rect 20044 34420 20084 34460
rect 17068 34336 17108 34376
rect 18988 34336 19028 34376
rect 19660 34336 19700 34376
rect 20140 34336 20180 34376
rect 21292 34252 21332 34292
rect 17548 34168 17588 34208
rect 18316 34168 18356 34208
rect 19180 34168 19220 34208
rect 21100 34168 21140 34208
rect 19852 34084 19892 34124
rect 20140 34084 20180 34124
rect 18808 34000 18848 34040
rect 18890 34000 18930 34040
rect 18972 34000 19012 34040
rect 19054 34000 19094 34040
rect 19136 34000 19176 34040
rect 10444 33748 10484 33788
rect 14092 33748 14132 33788
rect 20620 33748 20660 33788
rect 10060 33664 10100 33704
rect 10828 33664 10868 33704
rect 15436 33664 15476 33704
rect 9580 33580 9620 33620
rect 10252 33580 10292 33620
rect 10924 33580 10932 33620
rect 10932 33580 10964 33620
rect 13804 33580 13844 33620
rect 16300 33580 16340 33620
rect 16588 33580 16628 33620
rect 16780 33580 16820 33620
rect 18508 33580 18548 33620
rect 18796 33580 18836 33620
rect 3340 33496 3380 33536
rect 9868 33496 9908 33536
rect 15724 33496 15764 33536
rect 17452 33496 17492 33536
rect 3724 33412 3764 33452
rect 8908 33412 8948 33452
rect 9580 33412 9620 33452
rect 15244 33412 15284 33452
rect 18508 33412 18548 33452
rect 19564 33412 19604 33452
rect 19948 33412 19988 33452
rect 268 33328 308 33368
rect 2956 33328 2996 33368
rect 3148 33328 3188 33368
rect 11692 33328 11732 33368
rect 1132 33244 1172 33284
rect 4928 33244 4968 33284
rect 5010 33244 5050 33284
rect 5092 33244 5132 33284
rect 5174 33244 5214 33284
rect 5256 33244 5296 33284
rect 5932 33244 5972 33284
rect 9004 33244 9044 33284
rect 1420 33160 1460 33200
rect 1708 33160 1748 33200
rect 19852 33328 19892 33368
rect 20048 33244 20088 33284
rect 20130 33244 20170 33284
rect 20212 33244 20252 33284
rect 20294 33244 20334 33284
rect 20376 33244 20416 33284
rect 8236 33160 8276 33200
rect 8428 33160 8468 33200
rect 8620 33160 8660 33200
rect 11980 33160 12020 33200
rect 19756 33160 19796 33200
rect 20620 33160 20660 33200
rect 3436 33076 3476 33116
rect 4396 33076 4436 33116
rect 7948 33076 7988 33116
rect 10924 33076 10964 33116
rect 13804 33076 13844 33116
rect 16300 33076 16340 33116
rect 76 32992 116 33032
rect 4300 32992 4340 33032
rect 940 32908 980 32948
rect 1900 32908 1940 32948
rect 2092 32908 2132 32948
rect 2476 32908 2516 32948
rect 3820 32908 3860 32948
rect 4492 32939 4532 32948
rect 4492 32908 4532 32939
rect 5164 32908 5204 32948
rect 5548 32908 5588 32948
rect 6316 32939 6356 32948
rect 6316 32908 6356 32939
rect 6796 32939 6836 32948
rect 6796 32908 6836 32939
rect 172 32824 212 32864
rect 1900 32740 1940 32780
rect 3628 32740 3668 32780
rect 76 32656 116 32696
rect 1708 32656 1748 32696
rect 7756 32992 7796 33032
rect 7468 32908 7508 32948
rect 7948 32908 7988 32948
rect 8428 32908 8468 32948
rect 9388 32908 9428 32948
rect 11212 32908 11252 32948
rect 11692 32908 11732 32948
rect 11980 32908 12020 32948
rect 13804 32908 13844 32948
rect 15244 32939 15284 32948
rect 15244 32908 15284 32939
rect 16588 32908 16628 32948
rect 16780 32908 16820 32948
rect 5260 32824 5300 32864
rect 5836 32824 5876 32864
rect 6892 32824 6932 32864
rect 8812 32824 8852 32864
rect 9580 32824 9620 32864
rect 13708 32824 13748 32864
rect 14284 32824 14324 32864
rect 4300 32740 4340 32780
rect 8044 32740 8084 32780
rect 15820 32824 15860 32864
rect 18508 32992 18548 33032
rect 21388 32992 21428 33032
rect 17932 32824 17972 32864
rect 18508 32824 18548 32864
rect 19948 32939 19988 32948
rect 19948 32908 19988 32939
rect 18700 32824 18740 32864
rect 19948 32740 19988 32780
rect 4588 32656 4628 32696
rect 7084 32656 7124 32696
rect 7468 32656 7508 32696
rect 7948 32656 7988 32696
rect 8332 32656 8372 32696
rect 9676 32656 9716 32696
rect 10348 32656 10388 32696
rect 14764 32656 14804 32696
rect 17356 32656 17396 32696
rect 8812 32572 8852 32612
rect 16780 32572 16820 32612
rect 17164 32572 17204 32612
rect 3688 32488 3728 32528
rect 3770 32488 3810 32528
rect 3852 32488 3892 32528
rect 3934 32488 3974 32528
rect 4016 32488 4056 32528
rect 7084 32404 7124 32444
rect 3532 32320 3572 32360
rect 5164 32320 5204 32360
rect 6796 32320 6836 32360
rect 2188 32236 2228 32276
rect 7948 32488 7988 32528
rect 10540 32488 10580 32528
rect 11404 32488 11444 32528
rect 8044 32404 8084 32444
rect 9100 32404 9140 32444
rect 12556 32404 12596 32444
rect 14380 32404 14420 32444
rect 17452 32404 17492 32444
rect 7372 32320 7412 32360
rect 7660 32320 7700 32360
rect 7084 32236 7124 32276
rect 8812 32320 8852 32360
rect 11692 32320 11732 32360
rect 12460 32320 12500 32360
rect 16684 32320 16724 32360
rect 18796 32656 18836 32696
rect 19468 32656 19508 32696
rect 20620 32656 20660 32696
rect 18808 32488 18848 32528
rect 18890 32488 18930 32528
rect 18972 32488 19012 32528
rect 19054 32488 19094 32528
rect 19136 32488 19176 32528
rect 20428 32404 20468 32444
rect 9484 32236 9524 32276
rect 13708 32236 13748 32276
rect 14860 32236 14900 32276
rect 19948 32236 19988 32276
rect 3148 32152 3188 32192
rect 6412 32152 6452 32192
rect 7564 32152 7604 32192
rect 8908 32152 8948 32192
rect 9388 32152 9428 32192
rect 9772 32152 9812 32192
rect 10060 32152 10100 32192
rect 11884 32152 11924 32192
rect 12076 32152 12116 32192
rect 17260 32152 17300 32192
rect 17932 32152 17972 32192
rect 18508 32152 18548 32192
rect 19564 32152 19604 32192
rect 1036 32068 1076 32108
rect 2476 32068 2516 32108
rect 2860 32068 2900 32108
rect 4780 32068 4820 32108
rect 5452 32068 5492 32108
rect 7276 32068 7316 32108
rect 10444 32068 10484 32108
rect 10828 32068 10868 32108
rect 11500 32068 11540 32108
rect 13516 32068 13556 32108
rect 13804 32068 13844 32108
rect 14188 32068 14228 32108
rect 14764 32068 14804 32108
rect 15244 32068 15252 32108
rect 15252 32068 15284 32108
rect 16300 32068 16340 32108
rect 17452 32068 17492 32108
rect 18700 32068 18740 32108
rect 1228 31984 1268 32024
rect 3052 31984 3092 32024
rect 9964 31984 10004 32024
rect 13708 31984 13748 32024
rect 15820 31984 15860 32024
rect 17836 31984 17876 32024
rect 18508 31984 18548 32024
rect 3340 31900 3380 31940
rect 6988 31900 7028 31940
rect 7660 31900 7700 31940
rect 6892 31816 6932 31856
rect 7372 31816 7412 31856
rect 8140 31816 8180 31856
rect 9388 31900 9428 31940
rect 12556 31900 12596 31940
rect 15532 31900 15572 31940
rect 17644 31900 17684 31940
rect 19084 31984 19124 32024
rect 12268 31816 12308 31856
rect 12460 31816 12500 31856
rect 13708 31816 13748 31856
rect 3148 31732 3188 31772
rect 4204 31732 4244 31772
rect 4928 31732 4968 31772
rect 5010 31732 5050 31772
rect 5092 31732 5132 31772
rect 5174 31732 5214 31772
rect 5256 31732 5296 31772
rect 5548 31732 5588 31772
rect 10444 31732 10484 31772
rect 11308 31732 11348 31772
rect 16300 31732 16340 31772
rect 19468 31732 19508 31772
rect 21196 31900 21236 31940
rect 20048 31732 20088 31772
rect 20130 31732 20170 31772
rect 20212 31732 20252 31772
rect 20294 31732 20334 31772
rect 20376 31732 20416 31772
rect 172 31648 212 31688
rect 4492 31648 4532 31688
rect 1420 31396 1460 31436
rect 4300 31564 4340 31604
rect 6412 31564 6443 31604
rect 6443 31564 6452 31604
rect 9964 31564 10004 31604
rect 11500 31564 11540 31604
rect 18508 31564 18548 31604
rect 3052 31480 3092 31520
rect 5260 31480 5300 31520
rect 5836 31480 5876 31520
rect 8716 31480 8756 31520
rect 10540 31480 10580 31520
rect 4204 31396 4244 31436
rect 5164 31396 5204 31436
rect 6796 31396 6836 31436
rect 7276 31396 7316 31436
rect 652 31312 692 31352
rect 3052 31312 3092 31352
rect 2860 31144 2900 31184
rect 3532 31144 3572 31184
rect 5740 31144 5780 31184
rect 2188 30976 2228 31016
rect 3688 30976 3728 31016
rect 3770 30976 3810 31016
rect 3852 30976 3892 31016
rect 3934 30976 3974 31016
rect 4016 30976 4056 31016
rect 2668 30808 2708 30848
rect 4492 30808 4523 30848
rect 4523 30808 4532 30848
rect 3340 30724 3380 30764
rect 4300 30724 4340 30764
rect 6220 31312 6251 31352
rect 6251 31312 6260 31352
rect 4876 31060 4916 31100
rect 14860 31480 14900 31520
rect 15436 31480 15476 31520
rect 16108 31480 16148 31520
rect 9676 31396 9716 31436
rect 9964 31396 10004 31436
rect 12076 31396 12116 31436
rect 12748 31396 12788 31436
rect 13900 31396 13940 31436
rect 14956 31396 14996 31436
rect 13132 31228 13172 31268
rect 8236 31144 8276 31184
rect 10252 31144 10292 31184
rect 12076 31144 12116 31184
rect 6796 31060 6836 31100
rect 12268 31060 12308 31100
rect 5068 30892 5108 30932
rect 13132 30892 13172 30932
rect 5740 30808 5780 30848
rect 9100 30808 9140 30848
rect 748 30640 788 30680
rect 3052 30640 3092 30680
rect 16204 31396 16244 31436
rect 17452 31396 17492 31436
rect 18220 31396 18260 31436
rect 14572 31312 14612 31352
rect 16588 31312 16628 31352
rect 16972 31312 17012 31352
rect 19468 31396 19508 31436
rect 20044 31427 20084 31436
rect 20044 31396 20084 31427
rect 14764 31228 14804 31268
rect 15820 31228 15860 31268
rect 16108 31228 16148 31268
rect 14188 31144 14228 31184
rect 14860 31144 14900 31184
rect 15052 31144 15083 31184
rect 15083 31144 15092 31184
rect 16588 31144 16628 31184
rect 18808 30976 18848 31016
rect 18890 30976 18930 31016
rect 18972 30976 19012 31016
rect 19054 30976 19094 31016
rect 19136 30976 19176 31016
rect 10828 30808 10868 30848
rect 14572 30808 14612 30848
rect 19564 30808 19604 30848
rect 19756 30808 19796 30848
rect 20908 30808 20948 30848
rect 9580 30724 9620 30764
rect 12940 30724 12980 30764
rect 18124 30724 18164 30764
rect 21100 30724 21140 30764
rect 6892 30640 6932 30680
rect 7564 30640 7604 30680
rect 10636 30640 10676 30680
rect 364 30556 404 30596
rect 1420 30556 1460 30596
rect 2476 30556 2516 30596
rect 2668 30304 2708 30344
rect 3916 30304 3956 30344
rect 4492 30556 4532 30596
rect 5068 30556 5108 30596
rect 7468 30556 7508 30596
rect 4204 30472 4244 30512
rect 7372 30472 7412 30512
rect 12364 30556 12404 30596
rect 15916 30640 15956 30680
rect 17164 30640 17204 30680
rect 18412 30640 18452 30680
rect 18796 30640 18836 30680
rect 19372 30640 19412 30680
rect 19756 30640 19796 30680
rect 20140 30640 20180 30680
rect 13708 30556 13748 30596
rect 13900 30556 13940 30596
rect 14380 30556 14420 30596
rect 13132 30472 13172 30512
rect 14572 30472 14612 30512
rect 15724 30472 15764 30512
rect 8716 30388 8756 30428
rect 8908 30388 8948 30428
rect 4300 30304 4340 30344
rect 12844 30304 12884 30344
rect 4928 30220 4968 30260
rect 5010 30220 5050 30260
rect 5092 30220 5132 30260
rect 5174 30220 5214 30260
rect 5256 30220 5296 30260
rect 2860 30136 2900 30176
rect 12940 30136 12980 30176
rect 2668 30052 2708 30092
rect 3148 30052 3188 30092
rect 4204 30052 4244 30092
rect 6316 30052 6356 30092
rect 10636 30052 10676 30092
rect 844 29968 884 30008
rect 4876 29968 4916 30008
rect 7756 29968 7796 30008
rect 1324 29884 1364 29924
rect 4780 29884 4820 29924
rect 6220 29915 6260 29924
rect 6220 29884 6260 29915
rect 6892 29884 6932 29924
rect 7564 29884 7604 29924
rect 7948 29884 7988 29924
rect 8236 29915 8276 29924
rect 8236 29884 8276 29915
rect 14188 30388 14228 30428
rect 13324 30304 13364 30344
rect 17068 30556 17108 30596
rect 17740 30556 17780 30596
rect 20908 30556 20948 30596
rect 16396 30472 16436 30512
rect 20428 30472 20468 30512
rect 16972 30388 17012 30428
rect 15724 30304 15764 30344
rect 9196 29968 9236 30008
rect 10348 29968 10388 30008
rect 12652 29968 12692 30008
rect 12844 29968 12884 30008
rect 8908 29884 8948 29924
rect 10444 29884 10484 29924
rect 5740 29800 5780 29840
rect 9580 29800 9620 29840
rect 10060 29800 10100 29840
rect 4492 29716 4532 29756
rect 8716 29716 8756 29756
rect 9100 29716 9140 29756
rect 9388 29716 9428 29756
rect 76 29632 116 29672
rect 2860 29632 2900 29672
rect 4012 29632 4052 29672
rect 4588 29632 4628 29672
rect 6412 29548 6452 29588
rect 1324 29296 1364 29336
rect 3052 29296 3092 29336
rect 3688 29464 3728 29504
rect 3770 29464 3810 29504
rect 3852 29464 3892 29504
rect 3934 29464 3974 29504
rect 4016 29464 4056 29504
rect 6028 29464 6068 29504
rect 6316 29464 6356 29504
rect 8908 29464 8948 29504
rect 13900 30136 13940 30176
rect 14380 30220 14420 30260
rect 14476 30136 14516 30176
rect 14188 30052 14228 30092
rect 16780 30220 16820 30260
rect 20048 30220 20088 30260
rect 20130 30220 20170 30260
rect 20212 30220 20252 30260
rect 20294 30220 20334 30260
rect 20376 30220 20416 30260
rect 16300 30136 16340 30176
rect 19756 30136 19796 30176
rect 21100 30136 21140 30176
rect 14956 30052 14987 30092
rect 14987 30052 14996 30092
rect 15436 30052 15476 30092
rect 17836 30052 17876 30092
rect 18700 30052 18740 30092
rect 19852 30052 19892 30092
rect 14860 29968 14900 30008
rect 10636 29884 10676 29924
rect 11212 29915 11252 29924
rect 11212 29884 11252 29915
rect 12364 29800 12404 29840
rect 18988 29968 19028 30008
rect 16396 29884 16427 29924
rect 16427 29884 16436 29924
rect 16684 29884 16724 29924
rect 17260 29884 17300 29924
rect 13900 29800 13940 29840
rect 14188 29800 14228 29840
rect 17452 29800 17492 29840
rect 13708 29716 13748 29756
rect 9292 29632 9332 29672
rect 11788 29632 11828 29672
rect 12748 29632 12788 29672
rect 14476 29632 14516 29672
rect 11980 29548 12020 29588
rect 18412 29884 18452 29924
rect 19948 29884 19988 29924
rect 14764 29716 14804 29756
rect 14956 29716 14996 29756
rect 15820 29716 15860 29756
rect 16396 29716 16436 29756
rect 21004 30052 21044 30092
rect 19276 29800 19316 29840
rect 19756 29800 19796 29840
rect 14860 29632 14900 29672
rect 15436 29632 15476 29672
rect 15916 29632 15956 29672
rect 17068 29632 17108 29672
rect 17932 29632 17972 29672
rect 9292 29380 9332 29420
rect 16108 29380 16148 29420
rect 4012 29296 4052 29336
rect 4876 29296 4916 29336
rect 6508 29296 6548 29336
rect 11308 29296 11348 29336
rect 12940 29296 12980 29336
rect 13516 29296 13556 29336
rect 13708 29296 13748 29336
rect 460 29128 500 29168
rect 1612 29128 1652 29168
rect 1996 29128 2036 29168
rect 2476 29128 2516 29168
rect 3148 29128 3188 29168
rect 15628 29212 15668 29252
rect 4300 29128 4340 29168
rect 5548 29128 5588 29168
rect 7564 29128 7604 29168
rect 9004 29128 9044 29168
rect 9292 29128 9332 29168
rect 9772 29128 9812 29168
rect 10348 29128 10388 29168
rect 10636 29128 10676 29168
rect 10828 29128 10868 29168
rect 2668 29044 2708 29084
rect 2860 29044 2885 29084
rect 2885 29044 2900 29084
rect 3724 29044 3764 29084
rect 6892 29044 6932 29084
rect 7468 29044 7508 29084
rect 8908 29044 8948 29084
rect 9484 29044 9524 29084
rect 10444 29044 10484 29084
rect 10924 29044 10964 29084
rect 11308 29044 11348 29084
rect 11980 29044 12020 29084
rect 13324 29044 13364 29084
rect 14860 29044 14900 29084
rect 3532 28960 3572 29000
rect 4300 28960 4340 29000
rect 2572 28876 2612 28916
rect 3916 28876 3956 28916
rect 4876 28876 4916 28916
rect 6796 28960 6836 29000
rect 7276 28960 7316 29000
rect 7376 28960 7416 29000
rect 10828 28960 10868 29000
rect 12844 28960 12884 29000
rect 14380 28960 14420 29000
rect 15052 28960 15092 29000
rect 15724 28960 15764 29000
rect 20428 29632 20468 29672
rect 21196 29632 21236 29672
rect 18808 29464 18848 29504
rect 18890 29464 18930 29504
rect 18972 29464 19012 29504
rect 19054 29464 19094 29504
rect 19136 29464 19176 29504
rect 17740 29296 17780 29336
rect 20620 29296 20660 29336
rect 16300 29128 16340 29168
rect 17260 29044 17300 29084
rect 17932 29128 17972 29168
rect 20524 29128 20564 29168
rect 21004 29128 21044 29168
rect 18412 29044 18452 29084
rect 19660 29044 19700 29084
rect 16108 28960 16148 29000
rect 18124 28960 18164 29000
rect 8524 28876 8564 28916
rect 9100 28876 9140 28916
rect 10060 28876 10100 28916
rect 12172 28876 12212 28916
rect 12556 28876 12596 28916
rect 15820 28876 15860 28916
rect 17068 28876 17108 28916
rect 17260 28876 17300 28916
rect 20044 28876 20084 28916
rect 2860 28792 2900 28832
rect 9004 28792 9044 28832
rect 9580 28792 9620 28832
rect 10348 28792 10388 28832
rect 15532 28792 15572 28832
rect 16684 28792 16724 28832
rect 1324 28708 1364 28748
rect 4928 28708 4968 28748
rect 5010 28708 5050 28748
rect 5092 28708 5132 28748
rect 5174 28708 5214 28748
rect 5256 28708 5296 28748
rect 1132 28624 1172 28664
rect 4012 28624 4052 28664
rect 2860 28540 2900 28580
rect 4204 28540 4244 28580
rect 18028 28708 18068 28748
rect 20048 28708 20088 28748
rect 20130 28708 20170 28748
rect 20212 28708 20252 28748
rect 20294 28708 20334 28748
rect 20376 28708 20416 28748
rect 8716 28624 8756 28664
rect 4876 28540 4916 28580
rect 5260 28540 5300 28580
rect 6412 28540 6452 28580
rect 6796 28540 6836 28580
rect 9004 28540 9044 28580
rect 10156 28540 10196 28580
rect 11308 28540 11348 28580
rect 11692 28540 11732 28580
rect 12748 28540 12788 28580
rect 3148 28456 3188 28496
rect 3916 28456 3956 28496
rect 4300 28456 4340 28496
rect 1612 28372 1652 28412
rect 2764 28403 2804 28412
rect 2764 28372 2804 28403
rect 3052 28372 3092 28412
rect 4588 28372 4628 28412
rect 4780 28372 4805 28412
rect 4805 28372 4820 28412
rect 5068 28372 5108 28412
rect 6796 28372 6836 28412
rect 7276 28372 7316 28412
rect 7564 28372 7604 28412
rect 7948 28372 7988 28412
rect 8332 28372 8372 28412
rect 460 28288 500 28328
rect 3340 28288 3380 28328
rect 3724 28288 3764 28328
rect 5644 28288 5684 28328
rect 7468 28288 7508 28328
rect 7756 28288 7796 28328
rect 2476 28204 2516 28244
rect 7276 28204 7316 28244
rect 10636 28456 10676 28496
rect 19852 28624 19892 28664
rect 14764 28540 14804 28580
rect 15820 28540 15860 28580
rect 17452 28540 17492 28580
rect 19276 28540 19316 28580
rect 19948 28540 19988 28580
rect 16300 28456 16340 28496
rect 16684 28456 16724 28496
rect 9772 28372 9812 28412
rect 9964 28372 10004 28412
rect 11596 28372 11636 28412
rect 13996 28372 14036 28412
rect 14668 28372 14708 28412
rect 15820 28372 15860 28412
rect 16204 28372 16244 28412
rect 16588 28372 16628 28412
rect 17164 28372 17204 28412
rect 18028 28372 18068 28412
rect 20140 28372 20180 28412
rect 9004 28288 9044 28328
rect 10060 28288 10100 28328
rect 11308 28288 11348 28328
rect 8716 28204 8756 28244
rect 17932 28204 17972 28244
rect 3628 28120 3668 28160
rect 4588 28120 4628 28160
rect 10156 28120 10196 28160
rect 11788 28120 11828 28160
rect 12844 28120 12884 28160
rect 19564 28120 19604 28160
rect 3052 28036 3092 28076
rect 9964 28036 10004 28076
rect 13612 28036 13652 28076
rect 1996 27952 2036 27992
rect 3688 27952 3728 27992
rect 3770 27952 3810 27992
rect 3852 27952 3892 27992
rect 3934 27952 3974 27992
rect 4016 27952 4056 27992
rect 10060 27952 10100 27992
rect 6028 27868 6068 27908
rect 1804 27784 1844 27824
rect 2668 27784 2708 27824
rect 8332 27784 8372 27824
rect 10636 27784 10676 27824
rect 11212 27784 11252 27824
rect 2476 27700 2516 27740
rect 268 27616 308 27656
rect 2668 27616 2708 27656
rect 2476 27532 2516 27572
rect 2764 27532 2804 27572
rect 3340 27700 3380 27740
rect 3532 27700 3572 27740
rect 3916 27700 3956 27740
rect 3532 27532 3572 27572
rect 3916 27532 3947 27572
rect 3947 27532 3956 27572
rect 4588 27616 4628 27656
rect 4876 27616 4916 27656
rect 5260 27700 5300 27740
rect 10828 27700 10868 27740
rect 9292 27616 9332 27656
rect 9772 27616 9812 27656
rect 5644 27532 5684 27572
rect 6892 27532 6932 27572
rect 7852 27532 7892 27572
rect 8332 27532 8372 27572
rect 9196 27532 9236 27572
rect 11308 27532 11348 27572
rect 14860 27952 14900 27992
rect 18808 27952 18848 27992
rect 18890 27952 18930 27992
rect 18972 27952 19012 27992
rect 19054 27952 19094 27992
rect 19136 27952 19176 27992
rect 16780 27868 16820 27908
rect 15244 27784 15284 27824
rect 16108 27784 16148 27824
rect 12748 27700 12788 27740
rect 17452 27700 17492 27740
rect 18508 27700 18548 27740
rect 19948 28120 19988 28160
rect 20044 27700 20084 27740
rect 12268 27532 12308 27572
rect 13132 27532 13172 27572
rect 13804 27532 13844 27572
rect 15436 27532 15476 27572
rect 15820 27532 15860 27572
rect 17164 27532 17204 27572
rect 18508 27532 18548 27572
rect 19180 27532 19220 27572
rect 4012 27448 4052 27488
rect 5260 27448 5300 27488
rect 7756 27448 7796 27488
rect 8908 27448 8948 27488
rect 10444 27448 10484 27488
rect 12652 27448 12692 27488
rect 20524 27448 20564 27488
rect 2956 27364 2996 27404
rect 4204 27364 4244 27404
rect 4684 27364 4724 27404
rect 5740 27364 5780 27404
rect 6028 27364 6068 27404
rect 9964 27364 10004 27404
rect 11020 27364 11060 27404
rect 11980 27364 12020 27404
rect 16780 27364 16820 27404
rect 18220 27364 18260 27404
rect 19276 27364 19316 27404
rect 20044 27364 20084 27404
rect 21292 27364 21332 27404
rect 6508 27280 6548 27320
rect 11692 27280 11732 27320
rect 1324 27196 1364 27236
rect 4928 27196 4968 27236
rect 5010 27196 5050 27236
rect 5092 27196 5132 27236
rect 5174 27196 5214 27236
rect 5256 27196 5296 27236
rect 6604 27196 6644 27236
rect 9292 27196 9332 27236
rect 10060 27196 10100 27236
rect 19468 27196 19508 27236
rect 20048 27196 20088 27236
rect 20130 27196 20170 27236
rect 20212 27196 20252 27236
rect 20294 27196 20334 27236
rect 20376 27196 20416 27236
rect 15724 27112 15764 27152
rect 17740 27112 17780 27152
rect 19564 27112 19604 27152
rect 19756 27112 19796 27152
rect 3628 27028 3668 27068
rect 5644 27028 5684 27068
rect 7468 27028 7508 27068
rect 7948 27028 7988 27068
rect 8332 27028 8372 27068
rect 10828 27028 10868 27068
rect 11308 27028 11348 27068
rect 460 26944 500 26984
rect 2572 26944 2612 26984
rect 4588 26944 4628 26984
rect 5932 26944 5972 26984
rect 6508 26944 6548 26984
rect 1804 26860 1844 26900
rect 2764 26891 2804 26900
rect 2764 26860 2804 26891
rect 3532 26860 3572 26900
rect 3820 26860 3851 26900
rect 3851 26860 3860 26900
rect 6988 26860 7028 26900
rect 6796 26776 6836 26816
rect 7468 26860 7508 26900
rect 7756 26860 7796 26900
rect 7948 26860 7988 26900
rect 8524 26860 8564 26900
rect 8908 26860 8948 26900
rect 9772 26891 9812 26900
rect 9772 26860 9812 26891
rect 10060 26860 10100 26900
rect 16588 27028 16628 27068
rect 18796 27028 18836 27068
rect 14380 26944 14420 26984
rect 19564 26944 19604 26984
rect 12268 26860 12308 26900
rect 14668 26860 14708 26900
rect 16492 26891 16532 26900
rect 16492 26860 16532 26891
rect 16780 26860 16820 26900
rect 17068 26860 17108 26900
rect 18220 26860 18260 26900
rect 18508 26860 18548 26900
rect 19372 26860 19412 26900
rect 8140 26776 8180 26816
rect 8812 26776 8852 26816
rect 10636 26776 10676 26816
rect 12172 26776 12212 26816
rect 2188 26692 2228 26732
rect 268 26608 308 26648
rect 3148 26272 3188 26312
rect 3052 26104 3092 26144
rect 3688 26440 3728 26480
rect 3770 26440 3810 26480
rect 3852 26440 3892 26480
rect 3934 26440 3974 26480
rect 4016 26440 4056 26480
rect 3628 26104 3668 26144
rect 4300 26272 4340 26312
rect 7756 26692 7796 26732
rect 19660 26860 19700 26900
rect 11308 26692 11348 26732
rect 14668 26692 14708 26732
rect 17740 26776 17780 26816
rect 18700 26776 18740 26816
rect 18892 26776 18932 26816
rect 17068 26692 17108 26732
rect 6796 26608 6836 26648
rect 7276 26608 7316 26648
rect 9196 26608 9236 26648
rect 12172 26608 12212 26648
rect 13996 26608 14036 26648
rect 14572 26608 14612 26648
rect 16780 26608 16820 26648
rect 17260 26608 17300 26648
rect 17740 26608 17780 26648
rect 6700 26524 6740 26564
rect 7852 26524 7892 26564
rect 10060 26524 10100 26564
rect 13036 26524 13076 26564
rect 10828 26440 10868 26480
rect 11308 26440 11348 26480
rect 18808 26440 18848 26480
rect 18890 26440 18930 26480
rect 18972 26440 19012 26480
rect 19054 26440 19094 26480
rect 19136 26440 19176 26480
rect 9100 26356 9140 26396
rect 5356 26272 5396 26312
rect 7276 26272 7316 26312
rect 9292 26272 9331 26312
rect 9331 26272 9332 26312
rect 11692 26272 11732 26312
rect 13132 26272 13172 26312
rect 13996 26272 14036 26312
rect 18796 26272 18836 26312
rect 6796 26188 6836 26228
rect 6028 26104 6068 26144
rect 7468 26104 7508 26144
rect 9964 26188 10004 26228
rect 11596 26188 11636 26228
rect 14668 26188 14708 26228
rect 20524 26188 20564 26228
rect 7948 26104 7988 26144
rect 8812 26104 8852 26144
rect 9196 26104 9236 26144
rect 10060 26104 10100 26144
rect 11500 26104 11540 26144
rect 11692 26104 11732 26144
rect 11980 26104 12020 26144
rect 14476 26104 14516 26144
rect 15436 26104 15476 26144
rect 16204 26104 16244 26144
rect 1900 26020 1940 26060
rect 2380 26020 2420 26060
rect 2764 26020 2804 26060
rect 4684 26020 4724 26060
rect 5836 26020 5876 26060
rect 7276 26020 7316 26060
rect 8908 26020 8948 26060
rect 9964 26020 10004 26060
rect 10348 26020 10388 26060
rect 12268 26020 12308 26060
rect 13132 26020 13172 26060
rect 14572 26020 14612 26060
rect 16588 26020 16628 26060
rect 16780 26020 16788 26060
rect 16788 26020 16820 26060
rect 17260 26020 17300 26060
rect 18604 26020 18644 26060
rect 18796 26020 18836 26060
rect 20044 26020 20084 26060
rect 1324 25936 1364 25976
rect 3532 25936 3572 25976
rect 2764 25852 2804 25892
rect 4012 25852 4052 25892
rect 7468 25936 7508 25976
rect 8140 25936 8180 25976
rect 11308 25936 11348 25976
rect 11500 25936 11540 25976
rect 13804 25936 13844 25976
rect 13996 25936 14036 25976
rect 15340 25936 15380 25976
rect 9676 25852 9716 25892
rect 10636 25852 10676 25892
rect 11980 25852 12020 25892
rect 17740 25852 17780 25892
rect 19372 25852 19412 25892
rect 6028 25768 6068 25808
rect 9004 25768 9044 25808
rect 10060 25768 10100 25808
rect 11308 25768 11348 25808
rect 4928 25684 4968 25724
rect 5010 25684 5050 25724
rect 5092 25684 5132 25724
rect 5174 25684 5214 25724
rect 5256 25684 5296 25724
rect 15436 25684 15476 25724
rect 556 25600 596 25640
rect 2092 25432 2132 25472
rect 1804 25348 1844 25388
rect 4300 25516 4340 25556
rect 7852 25516 7892 25556
rect 9772 25516 9812 25556
rect 9964 25516 10004 25556
rect 3820 25432 3860 25472
rect 10540 25516 10580 25556
rect 11308 25516 11348 25556
rect 16204 25516 16244 25556
rect 7276 25348 7316 25388
rect 7852 25348 7892 25388
rect 9100 25348 9140 25388
rect 9292 25348 9332 25388
rect 9772 25348 9812 25388
rect 10348 25348 10388 25388
rect 11308 25348 11348 25388
rect 12268 25348 12308 25388
rect 76 25264 116 25304
rect 1228 25264 1268 25304
rect 3628 25264 3668 25304
rect 4876 25264 4916 25304
rect 7180 25264 7220 25304
rect 9964 25264 10004 25304
rect 652 25180 692 25220
rect 18316 25432 18356 25472
rect 18796 25432 18836 25472
rect 14668 25348 14708 25388
rect 14956 25348 14996 25388
rect 15724 25379 15764 25388
rect 15724 25348 15764 25379
rect 16684 25348 16724 25388
rect 13900 25264 13940 25304
rect 17740 25379 17780 25388
rect 17740 25348 17780 25379
rect 18604 25348 18644 25388
rect 16204 25264 16244 25304
rect 16972 25264 17012 25304
rect 18124 25264 18164 25304
rect 20048 25684 20088 25724
rect 20130 25684 20170 25724
rect 20212 25684 20252 25724
rect 20294 25684 20334 25724
rect 20376 25684 20416 25724
rect 20524 25600 20564 25640
rect 21100 25516 21140 25556
rect 21196 25432 21236 25472
rect 20716 25264 20756 25304
rect 5932 25180 5972 25220
rect 6700 25180 6740 25220
rect 12748 25180 12788 25220
rect 6508 25096 6548 25136
rect 9100 25096 9140 25136
rect 11020 25096 11060 25136
rect 13516 25096 13556 25136
rect 14572 25096 14612 25136
rect 20716 25096 20756 25136
rect 5836 25012 5876 25052
rect 13228 25012 13268 25052
rect 3688 24928 3728 24968
rect 3770 24928 3810 24968
rect 3852 24928 3892 24968
rect 3934 24928 3974 24968
rect 4016 24928 4056 24968
rect 6988 24928 7028 24968
rect 18808 24928 18848 24968
rect 18890 24928 18930 24968
rect 18972 24928 19012 24968
rect 19054 24928 19094 24968
rect 19136 24928 19176 24968
rect 6508 24844 6548 24884
rect 7852 24844 7892 24884
rect 12748 24844 12788 24884
rect 16972 24844 17012 24884
rect 17836 24844 17876 24884
rect 4588 24760 4628 24800
rect 5932 24760 5972 24800
rect 6124 24760 6164 24800
rect 3724 24676 3764 24716
rect 5452 24676 5492 24716
rect 652 24592 692 24632
rect 3340 24592 3380 24632
rect 4972 24592 5012 24632
rect 5260 24592 5300 24632
rect 5932 24592 5972 24632
rect 6316 24592 6356 24632
rect 7468 24760 7508 24800
rect 9388 24760 9428 24800
rect 11308 24760 11348 24800
rect 16204 24760 16244 24800
rect 8044 24676 8084 24716
rect 9004 24676 9044 24716
rect 14476 24676 14516 24716
rect 15340 24676 15380 24716
rect 6988 24592 7028 24632
rect 8524 24592 8564 24632
rect 14956 24592 14996 24632
rect 15436 24592 15476 24632
rect 1036 24508 1076 24548
rect 2572 24508 2612 24548
rect 2860 24508 2900 24548
rect 3628 24508 3668 24548
rect 4300 24508 4340 24548
rect 6892 24508 6932 24548
rect 7084 24508 7124 24548
rect 7468 24508 7508 24548
rect 7852 24508 7892 24548
rect 3052 24424 3092 24464
rect 4876 24424 4916 24464
rect 6316 24424 6356 24464
rect 10636 24508 10676 24548
rect 11020 24508 11060 24548
rect 11596 24508 11636 24548
rect 11884 24508 11924 24548
rect 13228 24508 13268 24548
rect 13516 24508 13556 24548
rect 14668 24508 14708 24548
rect 15628 24508 15668 24548
rect 19276 24760 19316 24800
rect 20140 24844 20180 24884
rect 21100 24844 21140 24884
rect 19852 24760 19892 24800
rect 21004 24760 21044 24800
rect 17260 24592 17300 24632
rect 21388 24676 21428 24716
rect 19276 24592 19316 24632
rect 21100 24592 21140 24632
rect 18316 24508 18356 24548
rect 19468 24508 19508 24548
rect 19948 24508 19988 24548
rect 21388 24508 21428 24548
rect 8812 24424 8852 24464
rect 18028 24424 18068 24464
rect 19852 24424 19892 24464
rect 20812 24424 20852 24464
rect 4300 24340 4340 24380
rect 9388 24340 9428 24380
rect 18796 24340 18836 24380
rect 4928 24172 4968 24212
rect 5010 24172 5050 24212
rect 5092 24172 5132 24212
rect 5174 24172 5214 24212
rect 5256 24172 5296 24212
rect 1612 24088 1652 24128
rect 8044 24088 8084 24128
rect 7180 24004 7220 24044
rect 7852 24004 7892 24044
rect 9292 24004 9332 24044
rect 1036 23920 1076 23960
rect 3724 23920 3764 23960
rect 6796 23920 6836 23960
rect 8620 23920 8660 23960
rect 940 23836 980 23876
rect 2572 23867 2612 23876
rect 2572 23836 2612 23867
rect 4012 23836 4052 23876
rect 4684 23836 4724 23876
rect 5836 23836 5876 23876
rect 6988 23836 7028 23876
rect 7276 23867 7316 23876
rect 7276 23836 7316 23867
rect 9100 23867 9140 23876
rect 9100 23836 9140 23867
rect 3052 23752 3092 23792
rect 3628 23752 3668 23792
rect 4972 23752 5012 23792
rect 5452 23752 5492 23792
rect 5932 23752 5972 23792
rect 18988 24256 19028 24296
rect 19756 24256 19796 24296
rect 19372 24172 19412 24212
rect 20048 24172 20088 24212
rect 20130 24172 20170 24212
rect 20212 24172 20252 24212
rect 20294 24172 20334 24212
rect 20376 24172 20416 24212
rect 17836 24088 17876 24128
rect 15724 24004 15764 24044
rect 16588 24004 16628 24044
rect 19372 24004 19412 24044
rect 17836 23920 17876 23960
rect 18700 23920 18740 23960
rect 18988 23920 19028 23960
rect 21196 23920 21236 23960
rect 10444 23836 10484 23876
rect 11884 23836 11924 23876
rect 12652 23836 12692 23876
rect 13516 23836 13556 23876
rect 14188 23836 14228 23876
rect 14476 23836 14516 23876
rect 14668 23836 14708 23876
rect 18796 23836 18836 23876
rect 19660 23836 19700 23876
rect 20524 23836 20564 23876
rect 9388 23752 9428 23792
rect 11980 23752 12020 23792
rect 13996 23752 14036 23792
rect 14956 23752 14996 23792
rect 15724 23752 15764 23792
rect 16396 23752 16436 23792
rect 17836 23752 17876 23792
rect 18028 23752 18068 23792
rect 18604 23752 18644 23792
rect 19372 23752 19412 23792
rect 12172 23668 12212 23708
rect 3724 23584 3764 23624
rect 3916 23584 3956 23624
rect 7084 23584 7124 23624
rect 7948 23584 7988 23624
rect 10828 23584 10868 23624
rect 13612 23584 13652 23624
rect 16012 23584 16052 23624
rect 14284 23500 14324 23540
rect 18124 23668 18164 23708
rect 18700 23668 18740 23708
rect 17260 23584 17300 23624
rect 17836 23584 17876 23624
rect 18220 23584 18260 23624
rect 19756 23584 19796 23624
rect 19948 23584 19979 23624
rect 19979 23584 19988 23624
rect 20812 23584 20852 23624
rect 3688 23416 3728 23456
rect 3770 23416 3810 23456
rect 3852 23416 3892 23456
rect 3934 23416 3974 23456
rect 4016 23416 4056 23456
rect 6796 23416 6836 23456
rect 1612 23332 1652 23372
rect 2956 23332 2996 23372
rect 4684 23332 4724 23372
rect 3628 23248 3668 23288
rect 5740 23248 5780 23288
rect 10060 23248 10100 23288
rect 10348 23248 10388 23288
rect 3148 23164 3188 23204
rect 748 23080 788 23120
rect 18808 23416 18848 23456
rect 18890 23416 18930 23456
rect 18972 23416 19012 23456
rect 19054 23416 19094 23456
rect 19136 23416 19176 23456
rect 10828 23248 10868 23288
rect 11884 23248 11924 23288
rect 15724 23248 15764 23288
rect 16588 23248 16628 23288
rect 16780 23248 16820 23288
rect 20044 23332 20084 23372
rect 13036 23164 13076 23204
rect 19564 23248 19604 23288
rect 19180 23164 19220 23204
rect 3340 23080 3380 23120
rect 3916 23080 3956 23120
rect 4300 23080 4340 23120
rect 7852 23080 7892 23120
rect 8428 23080 8468 23120
rect 9004 23080 9044 23120
rect 9388 23080 9428 23120
rect 9676 23080 9716 23120
rect 12268 23080 12308 23120
rect 14284 23080 14324 23120
rect 16684 23080 16724 23120
rect 17836 23080 17876 23120
rect 18796 23080 18836 23120
rect 21100 23080 21140 23120
rect 2380 22996 2420 23036
rect 3532 22996 3572 23036
rect 6028 22996 6068 23036
rect 7372 22996 7412 23036
rect 1132 22912 1172 22952
rect 3244 22912 3284 22952
rect 4012 22912 4052 22952
rect 4300 22912 4340 22952
rect 3532 22828 3572 22868
rect 7564 22828 7604 22868
rect 10348 22996 10388 23036
rect 4204 22744 4244 22784
rect 4928 22660 4968 22700
rect 5010 22660 5050 22700
rect 5092 22660 5132 22700
rect 5174 22660 5214 22700
rect 5256 22660 5296 22700
rect 5836 22576 5876 22616
rect 9004 22912 9044 22952
rect 13612 22996 13652 23036
rect 14188 22996 14228 23036
rect 14476 22996 14516 23036
rect 14668 22996 14708 23036
rect 15340 22996 15348 23036
rect 15348 22996 15380 23036
rect 16108 22996 16148 23036
rect 12268 22912 12308 22952
rect 8332 22828 8372 22868
rect 9964 22828 10004 22868
rect 12844 22828 12884 22868
rect 13900 22828 13940 22868
rect 15340 22828 15380 22868
rect 11500 22744 11540 22784
rect 15052 22744 15092 22784
rect 8332 22576 8372 22616
rect 3436 22492 3476 22532
rect 5452 22492 5492 22532
rect 6412 22492 6452 22532
rect 10348 22492 10388 22532
rect 13900 22492 13940 22532
rect 14668 22492 14699 22532
rect 14699 22492 14708 22532
rect 5548 22408 5588 22448
rect 7948 22408 7988 22448
rect 8620 22408 8660 22448
rect 12940 22408 12980 22448
rect 1900 22324 1940 22364
rect 3436 22324 3476 22364
rect 4108 22324 4148 22364
rect 4588 22324 4628 22364
rect 172 22240 212 22280
rect 844 22240 884 22280
rect 5356 22324 5396 22364
rect 16876 22996 16916 23036
rect 17260 22996 17300 23036
rect 18028 22996 18068 23036
rect 18892 22996 18932 23036
rect 19852 22996 19892 23036
rect 16492 22912 16532 22952
rect 19564 22828 19604 22868
rect 19852 22744 19892 22784
rect 20048 22660 20088 22700
rect 20130 22660 20170 22700
rect 20212 22660 20252 22700
rect 20294 22660 20334 22700
rect 20376 22660 20416 22700
rect 18892 22576 18932 22616
rect 18028 22492 18068 22532
rect 21004 22576 21044 22616
rect 18700 22492 18740 22532
rect 19852 22492 19892 22532
rect 19564 22408 19604 22448
rect 19948 22408 19988 22448
rect 6412 22324 6452 22364
rect 7468 22324 7508 22364
rect 8044 22324 8084 22364
rect 8332 22324 8372 22364
rect 9100 22324 9140 22364
rect 4396 22240 4436 22280
rect 6028 22240 6068 22280
rect 8428 22240 8468 22280
rect 8716 22240 8756 22280
rect 11500 22324 11540 22364
rect 12844 22324 12884 22364
rect 13132 22324 13172 22364
rect 12076 22240 12116 22280
rect 15052 22324 15092 22364
rect 16684 22324 16724 22364
rect 16876 22324 16916 22364
rect 17836 22324 17876 22364
rect 13996 22240 14036 22280
rect 14380 22240 14420 22280
rect 14572 22240 14612 22280
rect 18892 22324 18932 22364
rect 19180 22324 19220 22364
rect 19852 22324 19892 22364
rect 18508 22240 18548 22280
rect 3052 22156 3092 22196
rect 3820 22156 3860 22196
rect 4588 22156 4628 22196
rect 5932 22156 5972 22196
rect 10156 22156 10196 22196
rect 11308 22156 11348 22196
rect 13900 22156 13940 22196
rect 17260 22156 17300 22196
rect 18028 22156 18068 22196
rect 18796 22156 18836 22196
rect 19948 22240 19988 22280
rect 19084 22156 19124 22196
rect 19852 22156 19892 22196
rect 20236 22156 20276 22196
rect 8716 22072 8756 22112
rect 11500 22072 11540 22112
rect 18316 22072 18356 22112
rect 19660 22072 19700 22112
rect 21292 22072 21332 22112
rect 1420 21988 1460 22028
rect 3688 21904 3728 21944
rect 3770 21904 3810 21944
rect 3852 21904 3892 21944
rect 3934 21904 3974 21944
rect 4016 21904 4056 21944
rect 11212 21904 11252 21944
rect 18808 21904 18848 21944
rect 18890 21904 18930 21944
rect 18972 21904 19012 21944
rect 19054 21904 19094 21944
rect 19136 21904 19176 21944
rect 20044 21904 20084 21944
rect 1420 21820 1460 21860
rect 8332 21820 8372 21860
rect 11308 21820 11348 21860
rect 11500 21820 11540 21860
rect 19372 21820 19412 21860
rect 2860 21736 2900 21776
rect 4396 21736 4436 21776
rect 6412 21736 6452 21776
rect 8620 21736 8660 21776
rect 9004 21736 9044 21776
rect 19756 21736 19796 21776
rect 20524 21736 20564 21776
rect 3820 21652 3860 21692
rect 9100 21652 9140 21692
rect 1228 21568 1268 21608
rect 1612 21568 1652 21608
rect 2380 21568 2420 21608
rect 2956 21568 2996 21608
rect 3916 21568 3956 21608
rect 4300 21568 4340 21608
rect 6028 21568 6068 21608
rect 7180 21568 7220 21608
rect 7948 21568 7988 21608
rect 1132 21484 1172 21524
rect 1612 21316 1652 21356
rect 2380 21316 2420 21356
rect 3052 21400 3092 21440
rect 3628 21484 3668 21524
rect 6412 21484 6452 21524
rect 6988 21484 7028 21524
rect 4204 21400 4244 21440
rect 6508 21400 6548 21440
rect 8332 21400 8372 21440
rect 16300 21652 16340 21692
rect 19756 21568 19796 21608
rect 10156 21484 10196 21524
rect 10348 21484 10388 21524
rect 12076 21484 12116 21524
rect 13516 21484 13556 21524
rect 13900 21484 13940 21524
rect 14284 21484 14324 21524
rect 15436 21484 15476 21524
rect 15724 21484 15764 21524
rect 16300 21484 16340 21524
rect 17260 21484 17300 21524
rect 17740 21484 17780 21524
rect 18124 21484 18164 21524
rect 18988 21484 19019 21524
rect 19019 21484 19028 21524
rect 19180 21484 19220 21524
rect 19564 21484 19604 21524
rect 20044 21484 20075 21524
rect 20075 21484 20084 21524
rect 9100 21400 9140 21440
rect 12364 21400 12404 21440
rect 14668 21400 14708 21440
rect 3532 21316 3572 21356
rect 5260 21316 5300 21356
rect 5548 21316 5588 21356
rect 6892 21316 6932 21356
rect 11020 21316 11060 21356
rect 11212 21316 11252 21356
rect 13996 21316 14036 21356
rect 14380 21316 14420 21356
rect 14572 21316 14612 21356
rect 15340 21400 15380 21440
rect 16012 21316 16052 21356
rect 16588 21316 16628 21356
rect 18700 21316 18740 21356
rect 20236 21316 20276 21356
rect 12844 21232 12884 21272
rect 14476 21232 14516 21272
rect 14668 21232 14708 21272
rect 18124 21232 18164 21272
rect 4928 21148 4968 21188
rect 5010 21148 5050 21188
rect 5092 21148 5132 21188
rect 5174 21148 5214 21188
rect 5256 21148 5296 21188
rect 6412 21148 6452 21188
rect 8908 21148 8948 21188
rect 9292 21148 9332 21188
rect 10732 21148 10772 21188
rect 13324 21148 13364 21188
rect 13612 21148 13652 21188
rect 17164 21148 17204 21188
rect 20048 21148 20088 21188
rect 20130 21148 20170 21188
rect 20212 21148 20252 21188
rect 20294 21148 20334 21188
rect 20376 21148 20416 21188
rect 15340 21064 15380 21104
rect 21484 21064 21524 21104
rect 4012 20980 4052 21020
rect 5356 20980 5396 21020
rect 8716 20980 8756 21020
rect 9292 20980 9332 21020
rect 15724 20980 15764 21020
rect 940 20896 980 20936
rect 9100 20896 9140 20936
rect 1900 20812 1940 20852
rect 2380 20812 2420 20852
rect 2764 20812 2804 20852
rect 3820 20812 3860 20852
rect 5164 20843 5204 20852
rect 5164 20812 5204 20843
rect 6124 20812 6164 20852
rect 7180 20812 7220 20852
rect 7564 20812 7604 20852
rect 2668 20728 2708 20768
rect 5260 20728 5300 20768
rect 8620 20812 8660 20852
rect 9004 20812 9044 20852
rect 9580 20812 9620 20852
rect 10156 20812 10196 20852
rect 10540 20812 10580 20852
rect 11020 20812 11060 20852
rect 11788 20812 11828 20852
rect 12748 20812 12788 20852
rect 8140 20728 8180 20768
rect 13612 20896 13652 20936
rect 14668 20896 14708 20936
rect 16492 20896 16532 20936
rect 17644 20896 17684 20936
rect 18412 20896 18452 20936
rect 14380 20812 14420 20852
rect 15820 20812 15860 20852
rect 16204 20812 16244 20852
rect 17740 20812 17780 20852
rect 13516 20728 13556 20768
rect 19564 20812 19604 20852
rect 16108 20728 16148 20768
rect 16492 20728 16532 20768
rect 20140 20728 20180 20768
rect 20716 20980 20756 21020
rect 3628 20644 3668 20684
rect 6892 20644 6932 20684
rect 8812 20644 8852 20684
rect 9388 20644 9428 20684
rect 10924 20644 10964 20684
rect 20332 20644 20372 20684
rect 2860 20560 2900 20600
rect 8044 20560 8084 20600
rect 11308 20560 11348 20600
rect 10732 20476 10772 20516
rect 15340 20560 15380 20600
rect 18988 20560 19028 20600
rect 19948 20560 19988 20600
rect 20524 20560 20564 20600
rect 14476 20476 14516 20516
rect 16108 20476 16148 20516
rect 3688 20392 3728 20432
rect 3770 20392 3810 20432
rect 3852 20392 3892 20432
rect 3934 20392 3974 20432
rect 4016 20392 4056 20432
rect 5548 20392 5588 20432
rect 11212 20392 11252 20432
rect 13612 20392 13652 20432
rect 13900 20392 13940 20432
rect 17260 20392 17300 20432
rect 18808 20392 18848 20432
rect 18890 20392 18930 20432
rect 18972 20392 19012 20432
rect 19054 20392 19094 20432
rect 19136 20392 19176 20432
rect 9676 20308 9716 20348
rect 14380 20308 14420 20348
rect 18412 20308 18452 20348
rect 6028 20224 6068 20264
rect 6892 20224 6932 20264
rect 11980 20224 12020 20264
rect 14668 20224 14708 20264
rect 16492 20224 16532 20264
rect 19180 20224 19220 20264
rect 1612 20140 1652 20180
rect 10348 20140 10388 20180
rect 13516 20140 13556 20180
rect 14092 20140 14132 20180
rect 16300 20140 16340 20180
rect 19564 20140 19604 20180
rect 21196 20140 21236 20180
rect 268 20056 308 20096
rect 3340 20056 3380 20096
rect 7180 20056 7220 20096
rect 1228 19972 1268 20012
rect 1804 19972 1844 20012
rect 2572 19972 2612 20012
rect 4396 19972 4436 20012
rect 5356 19972 5396 20012
rect 6316 19972 6356 20012
rect 844 19888 884 19928
rect 10924 20056 10964 20096
rect 13324 20056 13364 20096
rect 7084 19972 7124 20012
rect 8908 19972 8948 20012
rect 9004 19888 9044 19928
rect 1900 19804 1940 19844
rect 4396 19804 4436 19844
rect 5452 19804 5492 19844
rect 460 19552 500 19592
rect 10156 19804 10196 19844
rect 17740 20056 17780 20096
rect 11212 19972 11252 20012
rect 11692 19972 11732 20012
rect 11980 19972 12020 20012
rect 12460 19972 12500 20012
rect 14380 19972 14420 20012
rect 14764 19972 14804 20012
rect 15244 19972 15284 20012
rect 16012 19972 16052 20012
rect 13516 19888 13556 19928
rect 13708 19888 13748 19928
rect 12364 19804 12404 19844
rect 13900 19804 13940 19844
rect 5932 19720 5972 19760
rect 7852 19720 7892 19760
rect 14668 19804 14708 19844
rect 16012 19804 16052 19844
rect 14380 19720 14420 19760
rect 4928 19636 4968 19676
rect 5010 19636 5050 19676
rect 5092 19636 5132 19676
rect 5174 19636 5214 19676
rect 5256 19636 5296 19676
rect 6220 19636 6260 19676
rect 8908 19636 8948 19676
rect 10444 19636 10484 19676
rect 11212 19636 11252 19676
rect 18028 20056 18068 20096
rect 18508 20056 18548 20096
rect 16684 19972 16724 20012
rect 17836 19972 17876 20012
rect 18892 19972 18932 20012
rect 19084 19972 19124 20012
rect 19948 19972 19988 20012
rect 20332 19972 20372 20012
rect 21196 19972 21236 20012
rect 20044 19804 20084 19844
rect 17164 19636 17204 19676
rect 20048 19636 20088 19676
rect 20130 19636 20170 19676
rect 20212 19636 20252 19676
rect 20294 19636 20334 19676
rect 20376 19636 20416 19676
rect 5932 19552 5972 19592
rect 15436 19552 15476 19592
rect 16012 19552 16052 19592
rect 18124 19552 18164 19592
rect 20524 19552 20564 19592
rect 4204 19468 4244 19508
rect 5260 19468 5300 19508
rect 10252 19468 10292 19508
rect 11116 19468 11156 19508
rect 11980 19468 12020 19508
rect 14476 19468 14516 19508
rect 15244 19468 15284 19508
rect 20140 19468 20180 19508
rect 5548 19384 5588 19424
rect 10444 19384 10484 19424
rect 11596 19384 11636 19424
rect 13228 19384 13268 19424
rect 14572 19384 14612 19424
rect 14764 19384 14804 19424
rect 16588 19384 16628 19424
rect 1612 19300 1652 19340
rect 1996 19300 2036 19340
rect 2572 19331 2612 19340
rect 2572 19300 2612 19331
rect 748 19216 788 19256
rect 4204 19300 4244 19340
rect 3628 19216 3668 19256
rect 3052 19132 3092 19172
rect 4396 19132 4436 19172
rect 3436 19048 3476 19088
rect 4204 19048 4244 19088
rect 3532 18880 3572 18920
rect 3688 18880 3728 18920
rect 3770 18880 3810 18920
rect 3852 18880 3892 18920
rect 3934 18880 3974 18920
rect 4016 18880 4056 18920
rect 8332 19300 8372 19340
rect 10060 19300 10100 19340
rect 12460 19300 12500 19340
rect 12652 19300 12692 19340
rect 13996 19300 14036 19340
rect 6124 19216 6164 19256
rect 7180 19216 7220 19256
rect 7852 19216 7892 19256
rect 8428 19216 8468 19256
rect 8716 19216 8756 19256
rect 9100 19216 9140 19256
rect 9676 19216 9716 19256
rect 13900 19216 13940 19256
rect 15052 19216 15092 19256
rect 6220 19132 6260 19172
rect 8044 19132 8084 19172
rect 19852 19384 19892 19424
rect 15724 19300 15764 19340
rect 16108 19300 16148 19340
rect 17836 19300 17876 19340
rect 18508 19300 18548 19340
rect 18892 19300 18932 19340
rect 19180 19300 19220 19340
rect 13804 19132 13844 19172
rect 15820 19216 15860 19256
rect 16012 19132 16052 19172
rect 6316 19048 6356 19088
rect 9676 19048 9716 19088
rect 13036 19048 13076 19088
rect 15820 19048 15860 19088
rect 6796 18880 6836 18920
rect 15052 18964 15092 19004
rect 16012 18964 16052 19004
rect 8908 18880 8948 18920
rect 12364 18880 12404 18920
rect 18808 18880 18848 18920
rect 18890 18880 18930 18920
rect 18972 18880 19012 18920
rect 19054 18880 19094 18920
rect 19136 18880 19176 18920
rect 19948 19331 19988 19340
rect 19948 19300 19988 19331
rect 20716 19048 20756 19088
rect 6508 18796 6548 18836
rect 11404 18796 11444 18836
rect 18508 18796 18548 18836
rect 1804 18712 1844 18752
rect 3532 18712 3572 18752
rect 9004 18712 9044 18752
rect 18796 18712 18836 18752
rect 19180 18712 19220 18752
rect 19564 18712 19604 18752
rect 19948 18712 19988 18752
rect 9676 18628 9716 18668
rect 14284 18628 14324 18668
rect 17068 18628 17108 18668
rect 19468 18628 19508 18668
rect 20812 18628 20852 18668
rect 1324 18544 1364 18584
rect 2956 18544 2996 18584
rect 4300 18544 4340 18584
rect 4588 18544 4628 18584
rect 4780 18544 4820 18584
rect 5068 18544 5108 18584
rect 5740 18544 5780 18584
rect 6508 18544 6548 18584
rect 7852 18544 7892 18584
rect 8716 18544 8756 18584
rect 13324 18544 13364 18584
rect 556 18460 596 18500
rect 2380 18460 2420 18500
rect 2860 18460 2900 18500
rect 3340 18460 3380 18500
rect 4012 18460 4020 18500
rect 4020 18460 4052 18500
rect 6988 18460 7028 18500
rect 7276 18460 7316 18500
rect 7660 18460 7700 18500
rect 8140 18460 8180 18500
rect 9100 18460 9108 18500
rect 9108 18460 9140 18500
rect 10636 18460 10676 18500
rect 10924 18460 10964 18500
rect 11692 18460 11732 18500
rect 17164 18544 17204 18584
rect 17932 18544 17972 18584
rect 18124 18544 18164 18584
rect 18700 18544 18740 18584
rect 20140 18544 20180 18584
rect 13900 18460 13940 18500
rect 15340 18460 15380 18500
rect 16108 18460 16148 18500
rect 16300 18460 16340 18500
rect 17836 18460 17876 18500
rect 19948 18460 19988 18500
rect 76 18376 116 18416
rect 2668 18376 2708 18416
rect 3052 18376 3092 18416
rect 3244 18376 3284 18416
rect 3628 18376 3668 18416
rect 4972 18376 5012 18416
rect 5164 18376 5204 18416
rect 6508 18376 6548 18416
rect 7180 18376 7220 18416
rect 8428 18376 8468 18416
rect 9004 18376 9044 18416
rect 12940 18376 12980 18416
rect 13132 18376 13172 18416
rect 18316 18376 18356 18416
rect 364 18292 404 18332
rect 7564 18292 7604 18332
rect 12076 18292 12116 18332
rect 12268 18292 12308 18332
rect 556 18208 596 18248
rect 4780 18208 4820 18248
rect 7660 18208 7700 18248
rect 1804 18124 1844 18164
rect 4928 18124 4968 18164
rect 5010 18124 5050 18164
rect 5092 18124 5132 18164
rect 5174 18124 5214 18164
rect 5256 18124 5296 18164
rect 8044 18124 8084 18164
rect 10156 18124 10196 18164
rect 13612 18124 13652 18164
rect 1516 17956 1556 17996
rect 4012 17956 4052 17996
rect 5836 17956 5876 17996
rect 9100 17956 9140 17996
rect 13900 17956 13940 17996
rect 1804 17872 1844 17912
rect 5548 17872 5588 17912
rect 6508 17872 6548 17912
rect 8428 17872 8468 17912
rect 8620 17872 8660 17912
rect 12268 17872 12308 17912
rect 1612 17788 1652 17828
rect 2860 17819 2900 17828
rect 2860 17788 2900 17819
rect 3244 17788 3284 17828
rect 3532 17788 3572 17828
rect 3916 17788 3956 17828
rect 4492 17819 4532 17828
rect 4492 17788 4532 17819
rect 4684 17788 4724 17828
rect 6028 17788 6068 17828
rect 7372 17788 7412 17828
rect 7852 17788 7892 17828
rect 8140 17788 8180 17828
rect 8812 17788 8852 17828
rect 9100 17788 9140 17828
rect 9484 17819 9524 17828
rect 9484 17788 9524 17819
rect 652 17704 692 17744
rect 4012 17704 4052 17744
rect 5356 17704 5396 17744
rect 5740 17704 5780 17744
rect 6508 17704 6548 17744
rect 8524 17704 8564 17744
rect 10636 17788 10676 17828
rect 11980 17788 12020 17828
rect 12556 17788 12596 17828
rect 10156 17704 10195 17744
rect 10195 17704 10196 17744
rect 11020 17704 11060 17744
rect 11692 17704 11732 17744
rect 15244 18292 15284 18332
rect 16108 18124 16148 18164
rect 16876 18124 16916 18164
rect 15244 18040 15284 18080
rect 15052 17872 15092 17912
rect 16492 17872 16532 17912
rect 21484 18208 21524 18248
rect 17932 18124 17972 18164
rect 18412 18124 18452 18164
rect 20048 18124 20088 18164
rect 20130 18124 20170 18164
rect 20212 18124 20252 18164
rect 20294 18124 20334 18164
rect 20376 18124 20416 18164
rect 19372 18040 19412 18080
rect 21100 17956 21140 17996
rect 15244 17788 15284 17828
rect 16684 17819 16724 17828
rect 16684 17788 16724 17819
rect 17260 17788 17300 17828
rect 15628 17704 15668 17744
rect 16492 17704 16532 17744
rect 17836 17704 17876 17744
rect 4876 17620 4916 17660
rect 7564 17620 7604 17660
rect 9964 17620 10004 17660
rect 14668 17620 14708 17660
rect 19276 17788 19316 17828
rect 18028 17704 18068 17744
rect 18604 17704 18644 17744
rect 19660 17704 19700 17744
rect 20140 17704 20180 17744
rect 19180 17620 19220 17660
rect 3052 17536 3092 17576
rect 7180 17536 7220 17576
rect 10348 17536 10388 17576
rect 14092 17536 14132 17576
rect 14380 17536 14420 17576
rect 15820 17536 15860 17576
rect 19468 17536 19508 17576
rect 19660 17536 19700 17576
rect 20908 17536 20948 17576
rect 3532 17452 3572 17492
rect 7084 17452 7124 17492
rect 8716 17452 8756 17492
rect 15244 17452 15284 17492
rect 3688 17368 3728 17408
rect 3770 17368 3810 17408
rect 3852 17368 3892 17408
rect 3934 17368 3974 17408
rect 4016 17368 4056 17408
rect 13324 17368 13364 17408
rect 18124 17368 18164 17408
rect 18604 17368 18644 17408
rect 18808 17368 18848 17408
rect 18890 17368 18930 17408
rect 18972 17368 19012 17408
rect 19054 17368 19094 17408
rect 19136 17368 19176 17408
rect 3340 17284 3380 17324
rect 4876 17284 4916 17324
rect 6220 17284 6260 17324
rect 6508 17284 6548 17324
rect 11020 17284 11060 17324
rect 17836 17284 17876 17324
rect 18028 17284 18068 17324
rect 4588 17200 4628 17240
rect 7276 17200 7316 17240
rect 8140 17200 8180 17240
rect 16684 17200 16724 17240
rect 17260 17200 17300 17240
rect 19276 17200 19316 17240
rect 19756 17200 19796 17240
rect 20044 17200 20084 17240
rect 21004 17200 21044 17240
rect 2380 17116 2420 17156
rect 2860 17116 2900 17156
rect 4204 17116 4244 17156
rect 10732 17116 10772 17156
rect 11404 17116 11444 17156
rect 12652 17116 12692 17156
rect 4012 17032 4052 17072
rect 7852 17032 7892 17072
rect 8332 17032 8372 17072
rect 9484 17032 9524 17072
rect 11500 17032 11540 17072
rect 13612 17032 13652 17072
rect 1228 16948 1268 16988
rect 2860 16948 2900 16988
rect 3436 16948 3476 16988
rect 3628 16948 3668 16988
rect 4300 16948 4340 16988
rect 5068 16948 5108 16988
rect 6508 16948 6548 16988
rect 7468 16948 7508 16988
rect 7948 16948 7988 16988
rect 9100 16948 9140 16988
rect 9868 16948 9908 16988
rect 10732 16948 10772 16988
rect 12268 16948 12308 16988
rect 13708 16948 13748 16988
rect 14284 16948 14324 16988
rect 14668 16948 14708 16988
rect 15436 16948 15476 16988
rect 18316 16948 18356 16988
rect 3820 16864 3860 16904
rect 4300 16780 4340 16820
rect 4204 16612 4244 16652
rect 1612 16528 1652 16568
rect 3724 16528 3764 16568
rect 6604 16780 6644 16820
rect 4928 16612 4968 16652
rect 5010 16612 5050 16652
rect 5092 16612 5132 16652
rect 5174 16612 5214 16652
rect 5256 16612 5296 16652
rect 6028 16528 6068 16568
rect 9964 16864 10004 16904
rect 10252 16780 10292 16820
rect 1708 16444 1748 16484
rect 6124 16444 6164 16484
rect 7180 16444 7220 16484
rect 10636 16444 10676 16484
rect 21292 17116 21332 17156
rect 20140 17032 20180 17072
rect 21196 16864 21236 16904
rect 16492 16780 16532 16820
rect 20524 16780 20564 16820
rect 19852 16696 19892 16736
rect 20048 16612 20088 16652
rect 20130 16612 20170 16652
rect 20212 16612 20252 16652
rect 20294 16612 20334 16652
rect 20376 16612 20416 16652
rect 21004 16528 21044 16568
rect 15052 16444 15092 16484
rect 16876 16444 16916 16484
rect 17836 16444 17876 16484
rect 19564 16444 19604 16484
rect 6604 16360 6644 16400
rect 7948 16360 7988 16400
rect 2380 16276 2420 16316
rect 2956 16307 2996 16316
rect 2956 16276 2996 16307
rect 3340 16276 3380 16316
rect 3820 16276 3860 16316
rect 4108 16276 4148 16316
rect 4972 16276 5012 16316
rect 5260 16307 5300 16316
rect 5260 16276 5300 16307
rect 8716 16307 8756 16316
rect 8716 16276 8756 16307
rect 9196 16276 9236 16316
rect 13708 16360 13748 16400
rect 268 16192 308 16232
rect 1036 16192 1076 16232
rect 3628 16192 3668 16232
rect 4492 16192 4532 16232
rect 5836 16192 5876 16232
rect 6028 16192 6068 16232
rect 10636 16276 10676 16316
rect 12268 16276 12308 16316
rect 13612 16276 13652 16316
rect 14476 16276 14516 16316
rect 14860 16307 14900 16316
rect 14860 16276 14900 16307
rect 19372 16360 19412 16400
rect 16972 16276 17012 16316
rect 18124 16276 18164 16316
rect 18508 16276 18548 16316
rect 18892 16276 18932 16316
rect 19660 16276 19700 16316
rect 20524 16276 20564 16316
rect 6604 16192 6644 16232
rect 6988 16192 7028 16232
rect 7468 16192 7508 16232
rect 8620 16192 8660 16232
rect 12364 16192 12404 16232
rect 12940 16192 12980 16232
rect 13804 16192 13844 16232
rect 14284 16192 14324 16232
rect 18700 16192 18740 16232
rect 3724 16108 3764 16148
rect 10636 16108 10676 16148
rect 16204 16108 16244 16148
rect 17260 16108 17300 16148
rect 20716 16108 20756 16148
rect 364 16024 404 16064
rect 5644 16024 5684 16064
rect 6028 16024 6068 16064
rect 8716 16024 8756 16064
rect 12172 16024 12212 16064
rect 17836 16024 17876 16064
rect 19948 16024 19988 16064
rect 21388 16024 21428 16064
rect 2572 15940 2612 15980
rect 6604 15940 6644 15980
rect 6988 15940 7028 15980
rect 10636 15940 10676 15980
rect 1324 15856 1364 15896
rect 3688 15856 3728 15896
rect 3770 15856 3810 15896
rect 3852 15856 3892 15896
rect 3934 15856 3974 15896
rect 4016 15856 4056 15896
rect 4300 15856 4340 15896
rect 5836 15856 5876 15896
rect 18808 15856 18848 15896
rect 18890 15856 18930 15896
rect 18972 15856 19012 15896
rect 19054 15856 19094 15896
rect 19136 15856 19176 15896
rect 14380 15772 14420 15812
rect 2764 15688 2804 15728
rect 4684 15688 4724 15728
rect 4204 15604 4244 15644
rect 5260 15604 5300 15644
rect 6604 15604 6644 15644
rect 6508 15520 6548 15560
rect 6988 15688 7028 15728
rect 10348 15688 10388 15728
rect 10732 15688 10772 15728
rect 12460 15688 12500 15728
rect 13228 15688 13268 15728
rect 14860 15688 14900 15728
rect 18124 15688 18164 15728
rect 9292 15604 9332 15644
rect 16300 15604 16340 15644
rect 12364 15520 12404 15560
rect 14284 15520 14324 15560
rect 18508 15520 18548 15560
rect 21196 15520 21236 15560
rect 364 15436 404 15476
rect 2764 15436 2804 15476
rect 3628 15436 3668 15476
rect 4300 15436 4340 15476
rect 5740 15436 5780 15476
rect 7180 15436 7220 15476
rect 7660 15436 7700 15476
rect 8908 15436 8948 15476
rect 12268 15436 12308 15476
rect 13036 15436 13076 15476
rect 14188 15436 14228 15476
rect 15436 15436 15476 15476
rect 16300 15436 16340 15476
rect 16972 15436 17012 15476
rect 17452 15436 17492 15476
rect 18124 15436 18164 15476
rect 18700 15436 18740 15476
rect 19372 15436 19412 15476
rect 20620 15436 20660 15476
rect 3148 15268 3188 15308
rect 8620 15268 8660 15308
rect 10636 15352 10676 15392
rect 9292 15268 9332 15308
rect 13228 15268 13268 15308
rect 364 15184 404 15224
rect 7276 15184 7316 15224
rect 17164 15352 17204 15392
rect 18508 15352 18548 15392
rect 9868 15184 9908 15224
rect 14188 15184 14228 15224
rect 17452 15268 17492 15308
rect 18220 15268 18260 15308
rect 20812 15268 20852 15308
rect 4928 15100 4968 15140
rect 5010 15100 5050 15140
rect 5092 15100 5132 15140
rect 5174 15100 5214 15140
rect 5256 15100 5296 15140
rect 9196 15100 9236 15140
rect 3628 15016 3668 15056
rect 9484 15016 9524 15056
rect 13036 15016 13076 15056
rect 13996 15016 14036 15056
rect 3340 14932 3380 14972
rect 4300 14932 4340 14972
rect 7180 14932 7220 14972
rect 7372 14932 7412 14972
rect 11596 14932 11636 14972
rect 14284 14932 14324 14972
rect 14668 14932 14708 14972
rect 15148 14932 15188 14972
rect 1516 14848 1556 14888
rect 5740 14848 5780 14888
rect 6988 14848 7028 14888
rect 1228 14764 1268 14804
rect 1996 14764 2036 14804
rect 3628 14764 3668 14804
rect 4684 14764 4724 14804
rect 8812 14848 8852 14888
rect 9196 14764 9236 14804
rect 9484 14795 9524 14804
rect 9484 14764 9524 14795
rect 9868 14764 9908 14804
rect 1996 14596 2036 14636
rect 4300 14596 4340 14636
rect 2572 14512 2612 14552
rect 4492 14512 4532 14552
rect 7084 14512 7124 14552
rect 3688 14344 3728 14384
rect 3770 14344 3810 14384
rect 3852 14344 3892 14384
rect 3934 14344 3974 14384
rect 4016 14344 4056 14384
rect 3340 14260 3380 14300
rect 6220 14260 6260 14300
rect 12172 14764 12212 14804
rect 12364 14764 12404 14804
rect 12940 14764 12980 14804
rect 13612 14764 13652 14804
rect 13996 14764 14036 14804
rect 14284 14764 14324 14804
rect 16876 15100 16916 15140
rect 18412 15100 18452 15140
rect 18604 15100 18644 15140
rect 20048 15100 20088 15140
rect 20130 15100 20170 15140
rect 20212 15100 20252 15140
rect 20294 15100 20334 15140
rect 20376 15100 20416 15140
rect 20812 15016 20852 15056
rect 18220 14932 18260 14972
rect 20524 14932 20564 14972
rect 18124 14848 18164 14888
rect 10348 14680 10388 14720
rect 13804 14680 13844 14720
rect 16876 14764 16916 14804
rect 17260 14764 17300 14804
rect 17164 14680 17204 14720
rect 18028 14680 18068 14720
rect 18220 14680 18260 14720
rect 19852 14680 19892 14720
rect 9292 14596 9332 14636
rect 10156 14596 10196 14636
rect 10636 14596 10676 14636
rect 15052 14596 15092 14636
rect 17356 14596 17396 14636
rect 20812 14596 20852 14636
rect 10444 14512 10484 14552
rect 11020 14512 11060 14552
rect 12460 14512 12500 14552
rect 14380 14512 14420 14552
rect 19756 14512 19796 14552
rect 16588 14428 16628 14468
rect 8140 14344 8180 14384
rect 11404 14344 11444 14384
rect 16012 14344 16052 14384
rect 17260 14344 17300 14384
rect 18808 14344 18848 14384
rect 18890 14344 18930 14384
rect 18972 14344 19012 14384
rect 19054 14344 19094 14384
rect 19136 14344 19176 14384
rect 7756 14260 7796 14300
rect 7468 14176 7508 14216
rect 12364 14176 12404 14216
rect 13996 14176 14036 14216
rect 15628 14176 15668 14216
rect 18508 14176 18548 14216
rect 20620 14176 20660 14216
rect 1900 14092 1940 14132
rect 2284 14092 2324 14132
rect 10348 14092 10388 14132
rect 13612 14092 13652 14132
rect 14284 14092 14324 14132
rect 14860 14092 14900 14132
rect 172 14008 212 14048
rect 1420 14008 1460 14048
rect 2380 14008 2420 14048
rect 3340 14008 3380 14048
rect 4396 14008 4436 14048
rect 5836 14008 5876 14048
rect 6220 14008 6260 14048
rect 7372 14008 7412 14048
rect 8524 14008 8564 14048
rect 1132 13924 1172 13964
rect 2860 13924 2900 13964
rect 3628 13924 3668 13964
rect 4108 13924 4116 13964
rect 4116 13924 4148 13964
rect 4492 13924 4532 13964
rect 7084 13924 7092 13964
rect 7092 13924 7124 13964
rect 7852 13924 7892 13964
rect 8140 13924 8180 13964
rect 9100 13924 9108 13964
rect 9108 13924 9140 13964
rect 76 13840 116 13880
rect 2476 13840 2516 13880
rect 2668 13840 2708 13880
rect 4588 13840 4628 13880
rect 5932 13840 5972 13880
rect 4492 13756 4532 13796
rect 5836 13756 5876 13796
rect 7660 13840 7700 13880
rect 7852 13756 7892 13796
rect 10156 14008 10196 14048
rect 15628 14008 15668 14048
rect 16492 14008 16532 14048
rect 16780 14008 16820 14048
rect 20812 14008 20852 14048
rect 11404 13924 11444 13964
rect 11596 13924 11636 13964
rect 12172 13924 12212 13964
rect 12460 13924 12500 13964
rect 13804 13924 13844 13964
rect 13996 13924 14036 13964
rect 16204 13924 16244 13964
rect 16396 13924 16436 13964
rect 16876 13924 16916 13964
rect 18124 13924 18164 13964
rect 12940 13840 12980 13880
rect 13612 13840 13652 13880
rect 12748 13756 12788 13796
rect 4928 13588 4968 13628
rect 5010 13588 5050 13628
rect 5092 13588 5132 13628
rect 5174 13588 5214 13628
rect 5256 13588 5296 13628
rect 5932 13588 5972 13628
rect 6124 13588 6164 13628
rect 12844 13588 12884 13628
rect 1804 13504 1844 13544
rect 5356 13504 5396 13544
rect 5548 13504 5588 13544
rect 7276 13504 7316 13544
rect 8620 13504 8660 13544
rect 11212 13504 11252 13544
rect 13036 13504 13076 13544
rect 15244 13840 15284 13880
rect 15436 13756 15476 13796
rect 17644 13756 17684 13796
rect 1612 13420 1652 13460
rect 3244 13420 3284 13460
rect 3532 13420 3572 13460
rect 4300 13420 4340 13460
rect 5164 13420 5204 13460
rect 7372 13420 7412 13460
rect 15436 13420 15476 13460
rect 76 13336 116 13376
rect 3148 13336 3188 13376
rect 5932 13336 5972 13376
rect 20048 13588 20088 13628
rect 20130 13588 20170 13628
rect 20212 13588 20252 13628
rect 20294 13588 20334 13628
rect 20376 13588 20416 13628
rect 16972 13504 17012 13544
rect 18700 13504 18740 13544
rect 19276 13504 19316 13544
rect 17356 13420 17396 13460
rect 17836 13420 17876 13460
rect 19852 13420 19892 13460
rect 21292 13420 21332 13460
rect 10636 13336 10676 13376
rect 940 13252 980 13292
rect 1420 13252 1460 13292
rect 1900 13252 1940 13292
rect 3436 13252 3476 13292
rect 5548 13252 5588 13292
rect 7372 13252 7412 13292
rect 10828 13283 10868 13292
rect 10828 13252 10868 13283
rect 11788 13252 11828 13292
rect 13132 13252 13172 13292
rect 14188 13283 14228 13292
rect 14188 13252 14228 13283
rect 16108 13252 16148 13292
rect 16300 13252 16340 13292
rect 16684 13252 16724 13292
rect 18316 13336 18356 13376
rect 18412 13252 18452 13292
rect 19660 13283 19700 13292
rect 19660 13252 19700 13283
rect 5260 13168 5300 13208
rect 6316 13168 6356 13208
rect 7660 13168 7700 13208
rect 7852 13168 7892 13208
rect 10444 13168 10484 13208
rect 16972 13168 17012 13208
rect 18124 13168 18164 13208
rect 20908 13168 20948 13208
rect 11500 13084 11540 13124
rect 1420 13000 1460 13040
rect 1708 13000 1748 13040
rect 2860 13000 2900 13040
rect 4300 13000 4340 13040
rect 5548 13000 5588 13040
rect 7660 13000 7700 13040
rect 11788 13000 11828 13040
rect 13420 13000 13460 13040
rect 16588 13000 16628 13040
rect 17356 13000 17396 13040
rect 20908 13000 20948 13040
rect 652 12916 692 12956
rect 17260 12916 17300 12956
rect 76 12832 116 12872
rect 3688 12832 3728 12872
rect 3770 12832 3810 12872
rect 3852 12832 3892 12872
rect 3934 12832 3974 12872
rect 4016 12832 4056 12872
rect 8524 12832 8564 12872
rect 14764 12832 14804 12872
rect 17452 12832 17492 12872
rect 18808 12832 18848 12872
rect 18890 12832 18930 12872
rect 18972 12832 19012 12872
rect 19054 12832 19094 12872
rect 19136 12832 19176 12872
rect 8140 12748 8180 12788
rect 15820 12748 15860 12788
rect 18700 12748 18740 12788
rect 5260 12664 5300 12704
rect 7852 12664 7892 12704
rect 14380 12664 14420 12704
rect 15244 12664 15284 12704
rect 16876 12664 16916 12704
rect 172 12580 212 12620
rect 8044 12580 8084 12620
rect 8524 12580 8564 12620
rect 8908 12580 8948 12620
rect 9772 12580 9812 12620
rect 12076 12580 12116 12620
rect 13516 12580 13556 12620
rect 16972 12580 17012 12620
rect 17356 12664 17396 12704
rect 19852 12664 19892 12704
rect 19276 12580 19316 12620
rect 652 12496 692 12536
rect 844 12496 884 12536
rect 2380 12496 2420 12536
rect 3052 12496 3092 12536
rect 3724 12496 3764 12536
rect 4300 12496 4340 12536
rect 4876 12496 4916 12536
rect 5164 12496 5204 12536
rect 5548 12496 5588 12536
rect 5836 12496 5876 12536
rect 6604 12496 6644 12536
rect 7852 12496 7892 12536
rect 9196 12496 9236 12536
rect 11788 12496 11828 12536
rect 12844 12496 12884 12536
rect 18412 12496 18452 12536
rect 18604 12496 18644 12536
rect 21004 12496 21044 12536
rect 460 12412 500 12452
rect 3244 12412 3284 12452
rect 3628 12412 3668 12452
rect 6124 12412 6164 12452
rect 748 12328 788 12368
rect 2572 12328 2612 12368
rect 9004 12412 9044 12452
rect 9868 12412 9908 12452
rect 12076 12412 12116 12452
rect 12460 12412 12500 12452
rect 12940 12412 12980 12452
rect 13420 12412 13428 12452
rect 13428 12412 13460 12452
rect 14764 12412 14804 12452
rect 15052 12412 15092 12452
rect 15436 12412 15476 12452
rect 15628 12412 15668 12452
rect 16684 12412 16724 12452
rect 17836 12412 17876 12452
rect 18124 12412 18164 12452
rect 18508 12412 18548 12452
rect 19372 12412 19412 12452
rect 6604 12328 6644 12368
rect 17452 12328 17492 12368
rect 2764 12244 2804 12284
rect 4300 12244 4340 12284
rect 5164 12244 5204 12284
rect 5548 12244 5588 12284
rect 5932 12244 5972 12284
rect 6124 12244 6164 12284
rect 8140 12244 8180 12284
rect 10060 12244 10100 12284
rect 16204 12244 16244 12284
rect 17164 12244 17204 12284
rect 748 12160 788 12200
rect 6412 12160 6452 12200
rect 9196 12160 9236 12200
rect 16108 12160 16148 12200
rect 16492 12160 16532 12200
rect 16972 12160 17012 12200
rect 4588 12076 4628 12116
rect 4928 12076 4968 12116
rect 5010 12076 5050 12116
rect 5092 12076 5132 12116
rect 5174 12076 5214 12116
rect 5256 12076 5296 12116
rect 556 11908 596 11948
rect 1612 11908 1652 11948
rect 940 11824 980 11864
rect 4684 11992 4724 12032
rect 7276 11992 7316 12032
rect 12940 11992 12980 12032
rect 14188 11992 14228 12032
rect 14956 11992 14996 12032
rect 4108 11908 4148 11948
rect 4300 11908 4340 11948
rect 6604 11908 6644 11948
rect 9100 11908 9140 11948
rect 17452 11908 17492 11948
rect 18316 11908 18356 11948
rect 20048 12076 20088 12116
rect 20130 12076 20170 12116
rect 20212 12076 20252 12116
rect 20294 12076 20334 12116
rect 20376 12076 20416 12116
rect 21004 11992 21044 12032
rect 4012 11824 4052 11864
rect 4972 11824 5012 11864
rect 8044 11824 8084 11864
rect 9292 11824 9332 11864
rect 10060 11824 10100 11864
rect 14380 11824 14420 11864
rect 14668 11824 14708 11864
rect 15436 11824 15476 11864
rect 19852 11824 19892 11864
rect 2860 11740 2900 11780
rect 4492 11656 4532 11696
rect 5740 11740 5780 11780
rect 6316 11771 6356 11780
rect 6316 11740 6356 11771
rect 6508 11740 6548 11780
rect 6988 11740 7028 11780
rect 8140 11740 8180 11780
rect 8524 11740 8564 11780
rect 8812 11740 8852 11780
rect 9388 11740 9428 11780
rect 9772 11771 9812 11780
rect 9772 11740 9812 11771
rect 11692 11740 11732 11780
rect 12940 11771 12980 11780
rect 12940 11740 12980 11771
rect 13516 11740 13556 11780
rect 13804 11740 13844 11780
rect 14956 11771 14996 11780
rect 14956 11740 14996 11771
rect 16972 11740 17012 11780
rect 17164 11740 17204 11780
rect 18508 11740 18548 11780
rect 9292 11656 9332 11696
rect 14380 11656 14420 11696
rect 16108 11656 16148 11696
rect 21388 11656 21428 11696
rect 2860 11572 2900 11612
rect 4396 11572 4436 11612
rect 18700 11572 18740 11612
rect 19660 11572 19700 11612
rect 1996 11488 2036 11528
rect 2380 11404 2420 11444
rect 10348 11488 10388 11528
rect 10732 11488 10772 11528
rect 16972 11488 17012 11528
rect 17644 11488 17684 11528
rect 18124 11488 18164 11528
rect 18508 11488 18548 11528
rect 3688 11320 3728 11360
rect 3770 11320 3810 11360
rect 3852 11320 3892 11360
rect 3934 11320 3974 11360
rect 4016 11320 4056 11360
rect 1900 11236 1940 11276
rect 460 11152 500 11192
rect 2668 11152 2708 11192
rect 1324 11068 1364 11108
rect 3436 11152 3476 11192
rect 6412 11152 6452 11192
rect 8524 11152 8564 11192
rect 11692 11404 11732 11444
rect 15340 11404 15380 11444
rect 15820 11404 15860 11444
rect 20044 11404 20084 11444
rect 2956 10984 2996 11024
rect 6412 10984 6452 11024
rect 7372 10984 7412 11024
rect 7948 10984 7988 11024
rect 13996 11320 14036 11360
rect 18316 11320 18356 11360
rect 18808 11320 18848 11360
rect 18890 11320 18930 11360
rect 18972 11320 19012 11360
rect 19054 11320 19094 11360
rect 19136 11320 19176 11360
rect 9868 11236 9908 11276
rect 11788 11236 11828 11276
rect 17740 11236 17780 11276
rect 11500 11152 11540 11192
rect 11884 11152 11924 11192
rect 2764 10900 2804 10940
rect 5356 10900 5396 10940
rect 1612 10816 1652 10856
rect 2476 10732 2516 10772
rect 6700 10900 6740 10940
rect 8044 10900 8084 10940
rect 6124 10816 6164 10856
rect 6892 10816 6932 10856
rect 9868 10816 9908 10856
rect 4300 10732 4340 10772
rect 7564 10732 7604 10772
rect 7852 10732 7892 10772
rect 8524 10732 8564 10772
rect 10252 10732 10292 10772
rect 12460 10900 12500 10940
rect 12076 10816 12116 10856
rect 2668 10648 2708 10688
rect 6892 10648 6932 10688
rect 11308 10648 11348 10688
rect 1804 10564 1844 10604
rect 4928 10564 4968 10604
rect 5010 10564 5050 10604
rect 5092 10564 5132 10604
rect 5174 10564 5214 10604
rect 5256 10564 5296 10604
rect 652 10480 692 10520
rect 268 10396 308 10436
rect 1516 10396 1556 10436
rect 2956 10396 2996 10436
rect 4588 10396 4628 10436
rect 14956 11152 14996 11192
rect 19372 11152 19412 11192
rect 19564 11152 19604 11192
rect 19948 11152 19988 11192
rect 14380 11068 14420 11108
rect 9004 10564 9044 10604
rect 14476 10900 14516 10940
rect 14380 10732 14420 10772
rect 19756 10984 19796 11024
rect 21196 10984 21236 11024
rect 21388 10984 21428 11024
rect 16492 10900 16532 10940
rect 16876 10900 16916 10940
rect 17740 10900 17780 10940
rect 18700 10900 18740 10940
rect 16396 10732 16436 10772
rect 17260 10648 17300 10688
rect 18028 10564 18068 10604
rect 20048 10564 20088 10604
rect 20130 10564 20170 10604
rect 20212 10564 20252 10604
rect 20294 10564 20334 10604
rect 20376 10564 20416 10604
rect 19564 10480 19604 10520
rect 8044 10396 8084 10436
rect 12460 10396 12500 10436
rect 12844 10396 12884 10436
rect 13708 10396 13748 10436
rect 17836 10396 17876 10436
rect 18028 10396 18068 10436
rect 18604 10396 18644 10436
rect 20524 10396 20564 10436
rect 3244 10312 3284 10352
rect 2764 10228 2804 10268
rect 7084 10312 7124 10352
rect 3628 10228 3668 10268
rect 4204 10228 4244 10268
rect 6508 10228 6548 10268
rect 172 10144 212 10184
rect 1708 10144 1748 10184
rect 2284 10144 2324 10184
rect 2860 10144 2900 10184
rect 3436 10144 3476 10184
rect 6316 10144 6356 10184
rect 11116 10312 11156 10352
rect 12172 10312 12212 10352
rect 12364 10312 12404 10352
rect 7564 10228 7604 10268
rect 10732 10228 10772 10268
rect 7852 10144 7892 10184
rect 9292 10144 9332 10184
rect 10060 10144 10100 10184
rect 10732 10060 10772 10100
rect 11404 10228 11444 10268
rect 11788 10228 11828 10268
rect 12076 10228 12116 10268
rect 11980 10144 12020 10184
rect 13804 10312 13844 10352
rect 16300 10312 16340 10352
rect 17644 10312 17684 10352
rect 18412 10312 18452 10352
rect 13996 10259 14036 10268
rect 13996 10228 14036 10259
rect 15628 10259 15668 10268
rect 15628 10228 15668 10259
rect 17452 10259 17492 10268
rect 17452 10228 17492 10259
rect 18508 10228 18548 10268
rect 14476 10144 14516 10184
rect 12748 10060 12788 10100
rect 13516 10060 13556 10100
rect 15340 10060 15380 10100
rect 18700 10144 18740 10184
rect 20812 10144 20852 10184
rect 19276 10060 19316 10100
rect 1708 9976 1748 10016
rect 6220 9976 6260 10016
rect 11116 9976 11156 10016
rect 13900 9976 13940 10016
rect 15916 9976 15956 10016
rect 21100 9976 21140 10016
rect 1228 9808 1268 9848
rect 364 9640 404 9680
rect 2284 9556 2324 9596
rect 2476 9556 2516 9596
rect 3688 9808 3728 9848
rect 3770 9808 3810 9848
rect 3852 9808 3892 9848
rect 3934 9808 3974 9848
rect 4016 9808 4056 9848
rect 8908 9808 8948 9848
rect 18124 9808 18164 9848
rect 18808 9808 18848 9848
rect 18890 9808 18930 9848
rect 18972 9808 19012 9848
rect 19054 9808 19094 9848
rect 19136 9808 19176 9848
rect 3436 9724 3476 9764
rect 9004 9724 9044 9764
rect 10252 9724 10292 9764
rect 10732 9724 10772 9764
rect 11500 9724 11540 9764
rect 15820 9724 15860 9764
rect 16492 9724 16532 9764
rect 3148 9640 3188 9680
rect 5548 9640 5588 9680
rect 5836 9640 5876 9680
rect 9868 9640 9908 9680
rect 15340 9640 15380 9680
rect 16876 9640 16916 9680
rect 18220 9640 18260 9680
rect 3532 9556 3572 9596
rect 16300 9556 16340 9596
rect 17644 9556 17684 9596
rect 4012 9472 4052 9512
rect 4684 9472 4724 9512
rect 9196 9472 9236 9512
rect 9868 9472 9908 9512
rect 10252 9472 10292 9512
rect 12748 9472 12788 9512
rect 14380 9472 14420 9512
rect 14764 9472 14804 9512
rect 15052 9472 15092 9512
rect 1708 9388 1748 9428
rect 2284 9388 2324 9428
rect 2476 9388 2516 9428
rect 5164 9388 5204 9428
rect 6220 9388 6260 9428
rect 4492 9304 4532 9344
rect 4684 9304 4724 9344
rect 6796 9304 6836 9344
rect 4108 9220 4148 9260
rect 6604 9220 6644 9260
rect 3532 9136 3572 9176
rect 18412 9472 18452 9512
rect 7564 9388 7604 9428
rect 8908 9388 8948 9428
rect 10060 9388 10100 9428
rect 11884 9388 11924 9428
rect 12844 9388 12884 9428
rect 13324 9388 13364 9428
rect 13804 9388 13844 9428
rect 14284 9388 14324 9428
rect 10156 9304 10196 9344
rect 12364 9304 12404 9344
rect 14476 9304 14516 9344
rect 10252 9220 10292 9260
rect 13612 9220 13652 9260
rect 16588 9220 16628 9260
rect 20044 9640 20084 9680
rect 20908 9472 20948 9512
rect 21196 9472 21236 9512
rect 17740 9388 17780 9428
rect 18700 9388 18740 9428
rect 19756 9388 19796 9428
rect 18604 9304 18644 9344
rect 17548 9220 17588 9260
rect 18124 9220 18164 9260
rect 19180 9220 19220 9260
rect 19660 9220 19700 9260
rect 6220 9136 6260 9176
rect 7180 9136 7220 9176
rect 13132 9136 13172 9176
rect 14188 9136 14228 9176
rect 4928 9052 4968 9092
rect 5010 9052 5050 9092
rect 5092 9052 5132 9092
rect 5174 9052 5214 9092
rect 5256 9052 5296 9092
rect 16300 9052 16340 9092
rect 18700 9052 18740 9092
rect 20048 9052 20088 9092
rect 20130 9052 20170 9092
rect 20212 9052 20252 9092
rect 20294 9052 20334 9092
rect 20376 9052 20416 9092
rect 7660 8968 7700 9008
rect 2572 8884 2612 8924
rect 1132 8800 1172 8840
rect 1900 8800 1940 8840
rect 1420 8716 1460 8756
rect 1804 8716 1844 8756
rect 2476 8747 2516 8756
rect 2476 8716 2516 8747
rect 4012 8884 4052 8924
rect 5068 8884 5108 8924
rect 7372 8884 7412 8924
rect 10060 8884 10100 8924
rect 11404 8884 11444 8924
rect 11884 8884 11924 8924
rect 13132 8884 13172 8924
rect 14860 8884 14900 8924
rect 15148 8884 15188 8924
rect 15916 8884 15956 8924
rect 16684 8884 16724 8924
rect 16972 8884 17012 8924
rect 18124 8884 18164 8924
rect 19276 8884 19316 8924
rect 3340 8800 3380 8840
rect 4684 8800 4724 8840
rect 3436 8716 3476 8756
rect 4108 8716 4148 8756
rect 3820 8632 3860 8672
rect 4588 8632 4628 8672
rect 6124 8800 6164 8840
rect 6700 8800 6740 8840
rect 10924 8800 10964 8840
rect 11980 8800 12020 8840
rect 14668 8800 14708 8840
rect 15628 8800 15668 8840
rect 16108 8800 16148 8840
rect 5836 8747 5876 8756
rect 5836 8716 5876 8747
rect 7084 8716 7124 8756
rect 7372 8747 7412 8756
rect 7372 8716 7412 8747
rect 7852 8747 7892 8756
rect 7852 8716 7892 8747
rect 8620 8716 8660 8756
rect 8908 8716 8948 8756
rect 6220 8632 6260 8672
rect 6700 8632 6740 8672
rect 10540 8716 10580 8756
rect 11596 8716 11636 8756
rect 11788 8716 11828 8756
rect 12364 8716 12404 8756
rect 12748 8716 12788 8756
rect 13324 8747 13364 8756
rect 13324 8716 13364 8747
rect 13804 8747 13844 8756
rect 13804 8716 13844 8747
rect 14188 8716 14228 8756
rect 16300 8716 16340 8756
rect 18412 8800 18452 8840
rect 17356 8747 17396 8756
rect 17356 8716 17396 8747
rect 19372 8716 19412 8756
rect 6892 8632 6932 8672
rect 11980 8632 12020 8672
rect 12844 8632 12884 8672
rect 16108 8632 16148 8672
rect 17452 8632 17492 8672
rect 19180 8632 19220 8672
rect 19564 8632 19604 8672
rect 19948 8632 19988 8672
rect 21004 8632 21044 8672
rect 6412 8548 6452 8588
rect 7564 8548 7604 8588
rect 12556 8548 12596 8588
rect 15820 8548 15860 8588
rect 16492 8548 16532 8588
rect 844 8464 884 8504
rect 10252 8464 10292 8504
rect 20908 8464 20948 8504
rect 11020 8380 11060 8420
rect 13324 8380 13364 8420
rect 3688 8296 3728 8336
rect 3770 8296 3810 8336
rect 3852 8296 3892 8336
rect 3934 8296 3974 8336
rect 4016 8296 4056 8336
rect 15052 8296 15092 8336
rect 18808 8296 18848 8336
rect 18890 8296 18930 8336
rect 18972 8296 19012 8336
rect 19054 8296 19094 8336
rect 19136 8296 19176 8336
rect 6412 8212 6452 8252
rect 9676 8212 9716 8252
rect 364 8128 404 8168
rect 2860 8128 2900 8168
rect 4492 8128 4532 8168
rect 5836 8128 5876 8168
rect 7852 8128 7892 8168
rect 2284 8044 2324 8084
rect 1516 7960 1556 8000
rect 6316 8044 6356 8084
rect 10924 8212 10964 8252
rect 11788 8128 11828 8168
rect 13804 8128 13844 8168
rect 13996 8128 14036 8168
rect 15340 8044 15380 8084
rect 1420 7876 1460 7916
rect 2764 7876 2804 7916
rect 6220 7876 6260 7916
rect 7180 7876 7220 7916
rect 8140 7876 8180 7916
rect 8620 7876 8660 7916
rect 11596 7876 11636 7916
rect 16300 8128 16340 8168
rect 17740 8128 17780 8168
rect 18508 8128 18548 8168
rect 18700 8044 18740 8084
rect 16012 7960 16052 8000
rect 18124 7960 18164 8000
rect 21388 7960 21428 8000
rect 16204 7876 16244 7916
rect 17452 7876 17492 7916
rect 18028 7876 18068 7916
rect 19372 7876 19412 7916
rect 20716 7876 20756 7916
rect 3148 7708 3188 7748
rect 4928 7540 4968 7580
rect 5010 7540 5050 7580
rect 5092 7540 5132 7580
rect 5174 7540 5214 7580
rect 5256 7540 5296 7580
rect 1036 7456 1076 7496
rect 4204 7372 4244 7412
rect 6700 7372 6740 7412
rect 6220 7288 6260 7328
rect 8716 7288 8756 7328
rect 2284 7204 2324 7244
rect 2764 7204 2804 7244
rect 4204 7204 4244 7244
rect 5740 7204 5780 7244
rect 7564 7204 7604 7244
rect 8140 7204 8180 7244
rect 9196 7204 9236 7244
rect 9772 7235 9812 7244
rect 9772 7204 9812 7235
rect 748 7120 788 7160
rect 1420 7120 1460 7160
rect 1804 7120 1844 7160
rect 1996 7120 2036 7160
rect 2860 7120 2900 7160
rect 4396 7120 4436 7160
rect 4588 7120 4628 7160
rect 5356 7120 5396 7160
rect 12556 7288 12596 7328
rect 11596 7204 11636 7244
rect 13324 7204 13364 7244
rect 15820 7708 15860 7748
rect 15340 7624 15380 7664
rect 18700 7624 18740 7664
rect 20048 7540 20088 7580
rect 20130 7540 20170 7580
rect 20212 7540 20252 7580
rect 20294 7540 20334 7580
rect 20376 7540 20416 7580
rect 17452 7456 17492 7496
rect 20524 7456 20564 7496
rect 15052 7372 15092 7412
rect 17452 7288 17492 7328
rect 14668 7235 14708 7244
rect 14668 7204 14708 7235
rect 16300 7235 16340 7244
rect 16300 7204 16340 7235
rect 18700 7204 18740 7244
rect 11308 7120 11348 7160
rect 16108 7120 16139 7160
rect 16139 7120 16148 7160
rect 17356 7120 17396 7160
rect 19660 7120 19700 7160
rect 21100 7120 21140 7160
rect 9868 7036 9908 7076
rect 10732 7036 10772 7076
rect 12076 7036 12116 7076
rect 14284 7036 14324 7076
rect 940 6952 980 6992
rect 3532 6952 3572 6992
rect 6220 6952 6260 6992
rect 12172 6952 12212 6992
rect 12364 6952 12404 6992
rect 15340 6952 15380 6992
rect 17356 6952 17396 6992
rect 19564 6952 19604 6992
rect 6124 6868 6164 6908
rect 3688 6784 3728 6824
rect 3770 6784 3810 6824
rect 3852 6784 3892 6824
rect 3934 6784 3974 6824
rect 4016 6784 4056 6824
rect 4396 6784 4436 6824
rect 6028 6784 6068 6824
rect 16396 6784 16436 6824
rect 18808 6784 18848 6824
rect 18890 6784 18930 6824
rect 18972 6784 19012 6824
rect 19054 6784 19094 6824
rect 19136 6784 19176 6824
rect 460 6616 500 6656
rect 1612 6616 1652 6656
rect 1228 6532 1268 6572
rect 2764 6616 2804 6656
rect 3148 6616 3188 6656
rect 4108 6616 4148 6656
rect 7948 6616 7988 6656
rect 12364 6616 12404 6656
rect 15820 6616 15860 6656
rect 19756 6616 19796 6656
rect 3340 6532 3380 6572
rect 6988 6532 7028 6572
rect 8620 6532 8660 6572
rect 16588 6532 16628 6572
rect 17260 6532 17300 6572
rect 21196 6532 21236 6572
rect 556 6448 596 6488
rect 1612 6448 1652 6488
rect 2284 6448 2324 6488
rect 9196 6448 9236 6488
rect 9868 6448 9908 6488
rect 10732 6448 10772 6488
rect 15052 6448 15092 6488
rect 15916 6448 15956 6488
rect 4204 6364 4244 6404
rect 5740 6364 5780 6404
rect 6892 6364 6932 6404
rect 8044 6364 8084 6404
rect 8716 6364 8756 6404
rect 9772 6364 9812 6404
rect 9964 6364 9972 6404
rect 9972 6364 10004 6404
rect 10540 6364 10580 6404
rect 12172 6364 12212 6404
rect 13324 6364 13364 6404
rect 14476 6364 14516 6404
rect 15340 6364 15380 6404
rect 16012 6364 16052 6404
rect 16684 6364 16724 6404
rect 16972 6364 16980 6404
rect 16980 6364 17012 6404
rect 18220 6364 18260 6404
rect 19372 6364 19412 6404
rect 19948 6364 19988 6404
rect 2860 6280 2900 6320
rect 6316 6280 6356 6320
rect 8908 6280 8948 6320
rect 11500 6280 11540 6320
rect 15628 6280 15668 6320
rect 16396 6280 16436 6320
rect 9868 6196 9908 6236
rect 10156 6196 10196 6236
rect 13036 6196 13076 6236
rect 14476 6196 14516 6236
rect 17260 6196 17300 6236
rect 1324 6112 1364 6152
rect 10060 6112 10100 6152
rect 13132 6112 13172 6152
rect 4928 6028 4968 6068
rect 5010 6028 5050 6068
rect 5092 6028 5132 6068
rect 5174 6028 5214 6068
rect 5256 6028 5296 6068
rect 9388 6028 9428 6068
rect 9964 6028 10004 6068
rect 10444 6028 10484 6068
rect 20048 6028 20088 6068
rect 20130 6028 20170 6068
rect 20212 6028 20252 6068
rect 20294 6028 20334 6068
rect 20376 6028 20416 6068
rect 6604 5944 6644 5984
rect 13324 5944 13364 5984
rect 14764 5944 14804 5984
rect 1420 5860 1460 5900
rect 4588 5860 4628 5900
rect 15052 5860 15092 5900
rect 15628 5860 15668 5900
rect 16972 5860 17012 5900
rect 268 5776 308 5816
rect 3340 5776 3380 5816
rect 6508 5776 6548 5816
rect 10540 5776 10580 5816
rect 10924 5776 10964 5816
rect 11308 5776 11348 5816
rect 364 5692 404 5732
rect 4300 5692 4340 5732
rect 6316 5692 6356 5732
rect 6892 5692 6932 5732
rect 8140 5723 8180 5732
rect 8140 5692 8180 5723
rect 652 5608 692 5648
rect 1996 5608 2036 5648
rect 2380 5608 2420 5648
rect 4876 5608 4916 5648
rect 10732 5692 10772 5732
rect 11596 5692 11636 5732
rect 172 5524 212 5564
rect 2092 5524 2132 5564
rect 3148 5524 3188 5564
rect 1708 5440 1748 5480
rect 10156 5608 10196 5648
rect 7948 5524 7988 5564
rect 9388 5524 9428 5564
rect 4780 5440 4820 5480
rect 6700 5440 6740 5480
rect 7084 5440 7124 5480
rect 10156 5440 10196 5480
rect 7372 5356 7412 5396
rect 3688 5272 3728 5312
rect 3770 5272 3810 5312
rect 3852 5272 3892 5312
rect 3934 5272 3974 5312
rect 4016 5272 4056 5312
rect 6508 5272 6548 5312
rect 9004 5272 9044 5312
rect 12460 5723 12500 5732
rect 12460 5692 12500 5723
rect 13036 5776 13076 5816
rect 14476 5776 14516 5816
rect 15820 5776 15860 5816
rect 13420 5692 13460 5732
rect 13996 5723 14036 5732
rect 13996 5692 14036 5723
rect 14764 5692 14804 5732
rect 15052 5692 15092 5732
rect 16300 5692 16340 5732
rect 16492 5692 16532 5732
rect 18700 5692 18740 5732
rect 20716 5692 20756 5732
rect 13900 5608 13940 5648
rect 19564 5608 19604 5648
rect 20908 5608 20948 5648
rect 11500 5524 11540 5564
rect 12844 5524 12884 5564
rect 13996 5524 14036 5564
rect 12076 5440 12116 5480
rect 13324 5440 13364 5480
rect 21292 5440 21332 5480
rect 11404 5272 11444 5312
rect 18808 5272 18848 5312
rect 18890 5272 18930 5312
rect 18972 5272 19012 5312
rect 19054 5272 19094 5312
rect 19136 5272 19176 5312
rect 844 5188 884 5228
rect 8620 5188 8660 5228
rect 10060 5188 10100 5228
rect 12076 5188 12116 5228
rect 13420 5188 13460 5228
rect 940 5104 980 5144
rect 1132 5104 1172 5144
rect 268 5020 308 5060
rect 1420 4936 1460 4976
rect 1996 5104 2036 5144
rect 3148 5104 3188 5144
rect 3340 5104 3380 5144
rect 7468 5104 7508 5144
rect 8044 5104 8084 5144
rect 10732 5104 10772 5144
rect 13132 5104 13172 5144
rect 15820 5104 15860 5144
rect 18604 5188 18644 5228
rect 16396 5104 16436 5144
rect 10156 5020 10196 5060
rect 11404 5020 11444 5060
rect 14668 5020 14708 5060
rect 2380 4936 2420 4976
rect 6508 4852 6548 4892
rect 3148 4768 3188 4808
rect 7276 4768 7316 4808
rect 11500 4936 11540 4976
rect 13324 4936 13364 4976
rect 8140 4852 8180 4892
rect 9004 4852 9044 4892
rect 10924 4852 10964 4892
rect 11884 4852 11924 4892
rect 12076 4852 12116 4892
rect 12556 4852 12596 4892
rect 14188 4852 14228 4892
rect 10252 4768 10292 4808
rect 1036 4684 1076 4724
rect 2092 4684 2132 4724
rect 4492 4684 4532 4724
rect 9868 4684 9908 4724
rect 13900 4768 13940 4808
rect 19948 4936 19988 4976
rect 20428 4936 20468 4976
rect 14668 4852 14708 4892
rect 15628 4852 15668 4892
rect 16684 4768 16724 4808
rect 12556 4684 12596 4724
rect 13420 4684 13460 4724
rect 15916 4684 15956 4724
rect 1420 4600 1460 4640
rect 17548 4600 17588 4640
rect 4928 4516 4968 4556
rect 5010 4516 5050 4556
rect 5092 4516 5132 4556
rect 5174 4516 5214 4556
rect 5256 4516 5296 4556
rect 6892 4516 6932 4556
rect 10636 4516 10676 4556
rect 11884 4516 11924 4556
rect 14668 4516 14708 4556
rect 16012 4516 16052 4556
rect 20048 4516 20088 4556
rect 20130 4516 20170 4556
rect 20212 4516 20252 4556
rect 20294 4516 20334 4556
rect 20376 4516 20416 4556
rect 364 4432 404 4472
rect 2380 4432 2420 4472
rect 6700 4432 6740 4472
rect 12076 4432 12116 4472
rect 3052 4348 3092 4388
rect 7756 4348 7796 4388
rect 8332 4348 8372 4388
rect 12556 4348 12596 4388
rect 556 4264 596 4304
rect 1324 4264 1364 4304
rect 17356 4264 17396 4304
rect 18316 4264 18356 4304
rect 10636 4180 10676 4220
rect 11500 4180 11540 4220
rect 12172 4211 12212 4220
rect 12172 4180 12212 4211
rect 2188 4096 2228 4136
rect 10828 4096 10868 4136
rect 21292 4096 21332 4136
rect 1516 4012 1556 4052
rect 1996 4012 2036 4052
rect 17836 4012 17876 4052
rect 12460 3928 12500 3968
rect 13516 3928 13556 3968
rect 20332 3928 20372 3968
rect 940 3844 980 3884
rect 3688 3760 3728 3800
rect 3770 3760 3810 3800
rect 3852 3760 3892 3800
rect 3934 3760 3974 3800
rect 4016 3760 4056 3800
rect 18808 3760 18848 3800
rect 18890 3760 18930 3800
rect 18972 3760 19012 3800
rect 19054 3760 19094 3800
rect 19136 3760 19176 3800
rect 17260 3676 17300 3716
rect 364 3592 404 3632
rect 1516 3592 1556 3632
rect 2188 3592 2228 3632
rect 8428 3592 8468 3632
rect 8620 3592 8660 3632
rect 17644 3592 17684 3632
rect 2668 3508 2708 3548
rect 3052 3508 3092 3548
rect 11980 3508 12020 3548
rect 13612 3508 13652 3548
rect 2380 3424 2420 3464
rect 3532 3424 3572 3464
rect 20332 3424 20372 3464
rect 12748 3256 12788 3296
rect 1804 3172 1844 3212
rect 18700 3172 18740 3212
rect 76 3088 116 3128
rect 1900 3088 1940 3128
rect 3532 3088 3572 3128
rect 4928 3004 4968 3044
rect 5010 3004 5050 3044
rect 5092 3004 5132 3044
rect 5174 3004 5214 3044
rect 5256 3004 5296 3044
rect 13804 3004 13844 3044
rect 20048 3004 20088 3044
rect 20130 3004 20170 3044
rect 20212 3004 20252 3044
rect 20294 3004 20334 3044
rect 20376 3004 20416 3044
rect 76 2920 116 2960
rect 4108 2836 4148 2876
rect 4684 2836 4724 2876
rect 10060 2920 10100 2960
rect 5836 2836 5876 2876
rect 8428 2836 8468 2876
rect 14284 2836 14324 2876
rect 1804 2752 1844 2792
rect 3532 2752 3572 2792
rect 4876 2752 4916 2792
rect 5740 2752 5780 2792
rect 17164 2752 17204 2792
rect 10156 2668 10196 2708
rect 11020 2668 11060 2708
rect 11692 2668 11732 2708
rect 12844 2668 12884 2708
rect 13420 2668 13460 2708
rect 13708 2668 13748 2708
rect 1420 2584 1460 2624
rect 1708 2584 1748 2624
rect 2092 2584 2132 2624
rect 2764 2584 2804 2624
rect 3148 2584 3188 2624
rect 3628 2584 3668 2624
rect 4108 2584 4148 2624
rect 4300 2584 4340 2624
rect 4684 2584 4724 2624
rect 5356 2584 5396 2624
rect 5836 2584 5876 2624
rect 9196 2584 9236 2624
rect 9676 2584 9716 2624
rect 10348 2584 10388 2624
rect 10732 2584 10772 2624
rect 11116 2584 11156 2624
rect 12268 2584 12308 2624
rect 13612 2584 13652 2624
rect 13996 2584 14036 2624
rect 14380 2584 14420 2624
rect 14764 2584 14804 2624
rect 15532 2584 15572 2624
rect 2476 2500 2516 2540
rect 5452 2500 5492 2540
rect 18700 2500 18740 2540
rect 3688 2248 3728 2288
rect 3770 2248 3810 2288
rect 3852 2248 3892 2288
rect 3934 2248 3974 2288
rect 4016 2248 4056 2288
rect 5260 2416 5300 2456
rect 5644 2416 5684 2456
rect 7276 2416 7316 2456
rect 8908 2416 8948 2456
rect 9292 2416 9332 2456
rect 9676 2416 9716 2456
rect 10060 2416 10100 2456
rect 10444 2416 10484 2456
rect 10828 2416 10868 2456
rect 12556 2416 12596 2456
rect 12940 2416 12980 2456
rect 13324 2416 13364 2456
rect 13708 2416 13748 2456
rect 14092 2416 14132 2456
rect 14476 2416 14516 2456
rect 14860 2416 14900 2456
rect 15244 2416 15284 2456
rect 6028 2332 6068 2372
rect 14188 2332 14228 2372
rect 18808 2248 18848 2288
rect 18890 2248 18930 2288
rect 18972 2248 19012 2288
rect 19054 2248 19094 2288
rect 19136 2248 19176 2288
rect 3052 2164 3092 2204
rect 17740 2164 17780 2204
rect 2284 2080 2324 2120
rect 2572 2080 2612 2120
rect 3340 2080 3380 2120
rect 4204 2080 4244 2120
rect 5548 2080 5588 2120
rect 6316 2080 6356 2120
rect 6700 2080 6740 2120
rect 6892 2080 6932 2120
rect 7756 2080 7796 2120
rect 12748 2080 12788 2120
rect 17356 2080 17396 2120
rect 2380 1996 2420 2036
rect 3724 1996 3764 2036
rect 5644 1996 5684 2036
rect 7084 1996 7124 2036
rect 7276 1996 7316 2036
rect 11308 1996 11348 2036
rect 12460 1996 12500 2036
rect 13900 1996 13940 2036
rect 19468 1996 19508 2036
rect 6412 1912 6452 1952
rect 6604 1912 6644 1952
rect 6988 1912 7028 1952
rect 8236 1912 8276 1952
rect 8620 1912 8660 1952
rect 9004 1912 9044 1952
rect 9388 1912 9428 1952
rect 9772 1912 9812 1952
rect 10156 1912 10196 1952
rect 10924 1912 10964 1952
rect 11500 1912 11540 1952
rect 12268 1912 12308 1952
rect 12652 1912 12692 1952
rect 13036 1912 13076 1952
rect 13420 1912 13460 1952
rect 14188 1912 14228 1952
rect 14572 1912 14612 1952
rect 15340 1912 15380 1952
rect 15724 1912 15764 1952
rect 16492 1912 16532 1952
rect 17356 1912 17396 1952
rect 2764 1828 2804 1868
rect 2956 1828 2996 1868
rect 3340 1828 3380 1868
rect 4204 1828 4244 1868
rect 4492 1828 4532 1868
rect 4780 1828 4820 1868
rect 5548 1828 5588 1868
rect 6028 1828 6068 1868
rect 6220 1828 6260 1868
rect 6796 1828 6836 1868
rect 8812 1828 8852 1868
rect 2572 1744 2612 1784
rect 3244 1744 3284 1784
rect 9196 1744 9236 1784
rect 11212 1744 11252 1784
rect 11788 1744 11828 1784
rect 12748 1744 12788 1784
rect 14668 1744 14708 1784
rect 2476 1660 2516 1700
rect 8716 1660 8756 1700
rect 9100 1660 9140 1700
rect 9484 1660 9524 1700
rect 9868 1660 9908 1700
rect 10252 1660 10292 1700
rect 10636 1660 10676 1700
rect 11020 1660 11060 1700
rect 11404 1660 11444 1700
rect 11596 1660 11636 1700
rect 11980 1660 12020 1700
rect 12172 1660 12212 1700
rect 4396 1576 4436 1616
rect 11692 1576 11732 1616
rect 12364 1576 12404 1616
rect 13132 1576 13172 1616
rect 13516 1576 13556 1616
rect 14284 1576 14324 1616
rect 15052 1576 15092 1616
rect 15436 1576 15476 1616
rect 4928 1492 4968 1532
rect 5010 1492 5050 1532
rect 5092 1492 5132 1532
rect 5174 1492 5214 1532
rect 5256 1492 5296 1532
rect 9964 1492 10004 1532
rect 10732 1492 10772 1532
rect 17644 1492 17684 1532
rect 20048 1492 20088 1532
rect 20130 1492 20170 1532
rect 20212 1492 20252 1532
rect 20294 1492 20334 1532
rect 20376 1492 20416 1532
<< metal3 >>
rect 1784 96688 1864 96768
rect 1976 96688 2056 96768
rect 2168 96688 2248 96768
rect 2360 96688 2440 96768
rect 2552 96688 2632 96768
rect 2744 96688 2824 96768
rect 2936 96688 3016 96768
rect 3128 96688 3208 96768
rect 3320 96688 3400 96768
rect 3512 96688 3592 96768
rect 3704 96688 3784 96768
rect 3896 96688 3976 96768
rect 4088 96688 4168 96768
rect 4280 96688 4360 96768
rect 4472 96688 4552 96768
rect 4664 96688 4744 96768
rect 4856 96688 4936 96768
rect 5048 96688 5128 96768
rect 5240 96688 5320 96768
rect 5432 96688 5512 96768
rect 5624 96688 5704 96768
rect 5816 96688 5896 96768
rect 6008 96688 6088 96768
rect 6200 96688 6280 96768
rect 6392 96688 6472 96768
rect 6584 96688 6664 96768
rect 6776 96688 6856 96768
rect 6968 96688 7048 96768
rect 7160 96688 7240 96768
rect 7352 96688 7432 96768
rect 7544 96688 7624 96768
rect 7736 96688 7816 96768
rect 7928 96688 8008 96768
rect 8120 96688 8200 96768
rect 8312 96688 8392 96768
rect 8504 96688 8584 96768
rect 8696 96688 8776 96768
rect 8888 96688 8968 96768
rect 9080 96688 9160 96768
rect 9272 96688 9352 96768
rect 9464 96688 9544 96768
rect 9656 96688 9736 96768
rect 9848 96688 9928 96768
rect 10040 96688 10120 96768
rect 10232 96688 10312 96768
rect 10424 96688 10504 96768
rect 10616 96688 10696 96768
rect 10808 96688 10888 96768
rect 11000 96688 11080 96768
rect 11192 96688 11272 96768
rect 11384 96688 11464 96768
rect 11576 96688 11656 96768
rect 11768 96688 11848 96768
rect 11960 96688 12040 96768
rect 12152 96688 12232 96768
rect 12344 96688 12424 96768
rect 12536 96688 12616 96768
rect 12728 96688 12808 96768
rect 12920 96688 13000 96768
rect 13112 96688 13192 96768
rect 13304 96688 13384 96768
rect 13496 96688 13576 96768
rect 13688 96688 13768 96768
rect 13880 96688 13960 96768
rect 14072 96688 14152 96768
rect 14264 96688 14344 96768
rect 14456 96688 14536 96768
rect 14648 96688 14728 96768
rect 14840 96688 14920 96768
rect 15032 96688 15112 96768
rect 15224 96688 15304 96768
rect 15416 96688 15496 96768
rect 15608 96688 15688 96768
rect 15800 96688 15880 96768
rect 15992 96688 16072 96768
rect 16184 96688 16264 96768
rect 16376 96688 16456 96768
rect 16568 96688 16648 96768
rect 16760 96688 16840 96768
rect 16952 96688 17032 96768
rect 17144 96688 17224 96768
rect 17336 96688 17416 96768
rect 17528 96688 17608 96768
rect 17720 96688 17800 96768
rect 17912 96688 17992 96768
rect 18104 96688 18184 96768
rect 18296 96688 18376 96768
rect 18488 96688 18568 96768
rect 18680 96688 18760 96768
rect 18872 96688 18952 96768
rect 19064 96688 19144 96768
rect 19256 96688 19336 96768
rect 19448 96688 19528 96768
rect 1324 94856 1364 94865
rect 1324 94721 1364 94816
rect 1708 94856 1748 94865
rect 1708 94721 1748 94816
rect 1228 94184 1268 94193
rect 76 93848 116 93857
rect 76 93680 116 93808
rect 76 93631 116 93640
rect 172 93596 212 93605
rect 172 93428 212 93556
rect 172 93379 212 93388
rect 460 93344 500 93353
rect 460 91832 500 93304
rect 1228 93176 1268 94144
rect 1804 93620 1844 96688
rect 1804 93580 1940 93620
rect 1228 93127 1268 93136
rect 1612 93344 1652 93353
rect 1228 92672 1268 92681
rect 1132 91916 1172 91925
rect 460 91783 500 91792
rect 748 91832 788 91841
rect 76 91328 116 91337
rect 76 88808 116 91288
rect 268 90992 308 91001
rect 76 88759 116 88768
rect 172 89564 212 89573
rect 76 88640 116 88649
rect 76 81752 116 88600
rect 76 81703 116 81712
rect 172 81416 212 89524
rect 268 85448 308 90952
rect 652 90320 692 90329
rect 268 85399 308 85408
rect 364 88808 404 88817
rect 172 81367 212 81376
rect 268 84272 308 84281
rect 76 81248 116 81257
rect 76 73016 116 81208
rect 76 72967 116 72976
rect 172 79064 212 79073
rect 76 72848 116 72857
rect 76 68648 116 72808
rect 172 70328 212 79024
rect 268 75368 308 84232
rect 364 79736 404 88768
rect 460 88724 500 88733
rect 460 80072 500 88684
rect 460 80023 500 80032
rect 556 88220 596 88229
rect 364 79687 404 79696
rect 268 75319 308 75328
rect 364 79568 404 79577
rect 268 74864 308 74873
rect 268 73688 308 74824
rect 364 74024 404 79528
rect 556 79400 596 88180
rect 652 83180 692 90280
rect 748 87128 788 91792
rect 748 87079 788 87088
rect 844 91160 884 91169
rect 652 83131 692 83140
rect 748 86204 788 86213
rect 652 82340 692 82349
rect 652 80912 692 82300
rect 652 80863 692 80872
rect 748 80744 788 86164
rect 844 85112 884 91120
rect 1036 90236 1076 90245
rect 844 85063 884 85072
rect 940 89648 980 89657
rect 652 80704 788 80744
rect 844 84188 884 84197
rect 652 80408 692 80704
rect 652 80359 692 80368
rect 748 80576 788 80585
rect 556 79351 596 79360
rect 652 80240 692 80249
rect 556 79232 596 79241
rect 364 73975 404 73984
rect 460 77552 500 77561
rect 268 73639 308 73648
rect 364 73856 404 73865
rect 364 73352 404 73816
rect 364 73303 404 73312
rect 172 70279 212 70288
rect 268 72176 308 72185
rect 76 68599 116 68608
rect 268 65624 308 72136
rect 268 65575 308 65584
rect 364 72092 404 72101
rect 364 65288 404 72052
rect 460 69320 500 77512
rect 556 75536 596 79192
rect 556 75487 596 75496
rect 652 75368 692 80200
rect 556 75328 692 75368
rect 556 74696 596 75328
rect 556 74647 596 74656
rect 652 75200 692 75209
rect 556 74444 596 74453
rect 556 72008 596 74404
rect 556 71959 596 71968
rect 460 69271 500 69280
rect 556 71252 596 71261
rect 460 69152 500 69161
rect 460 65960 500 69112
rect 460 65911 500 65920
rect 364 65239 404 65248
rect 556 64952 596 71212
rect 652 67304 692 75160
rect 748 72680 788 80536
rect 844 78392 884 84148
rect 940 81080 980 89608
rect 1036 83432 1076 90196
rect 1132 88472 1172 91876
rect 1228 90152 1268 92632
rect 1420 92672 1460 92681
rect 1324 92000 1364 92009
rect 1324 90824 1364 91960
rect 1324 90775 1364 90784
rect 1420 90488 1460 92632
rect 1612 92168 1652 93304
rect 1612 92119 1652 92128
rect 1708 93176 1748 93185
rect 1420 90439 1460 90448
rect 1516 91832 1556 91841
rect 1420 90320 1460 90329
rect 1420 90185 1460 90280
rect 1228 90103 1268 90112
rect 1420 90068 1460 90077
rect 1324 89900 1364 89909
rect 1132 88423 1172 88432
rect 1228 88892 1268 88901
rect 1132 87464 1172 87473
rect 1132 86120 1172 87424
rect 1228 86204 1268 88852
rect 1324 87464 1364 89860
rect 1420 89900 1460 90028
rect 1420 89851 1460 89860
rect 1420 89480 1460 89575
rect 1420 89431 1460 89440
rect 1324 87415 1364 87424
rect 1420 89312 1460 89321
rect 1228 86155 1268 86164
rect 1324 87296 1364 87305
rect 1132 86071 1172 86080
rect 1228 86036 1268 86045
rect 1228 85952 1268 85996
rect 1036 83383 1076 83392
rect 1132 85912 1268 85952
rect 940 81031 980 81040
rect 1036 82256 1076 82265
rect 844 78343 884 78352
rect 940 80912 980 80921
rect 844 76796 884 76805
rect 844 75284 884 76756
rect 940 75704 980 80872
rect 1036 79148 1076 82216
rect 1132 80744 1172 85912
rect 1132 80695 1172 80704
rect 1228 85784 1268 85793
rect 1036 79099 1076 79108
rect 1132 80492 1172 80501
rect 940 75655 980 75664
rect 1036 76880 1076 76889
rect 844 75244 980 75284
rect 748 72631 788 72640
rect 844 75116 884 75125
rect 748 70748 788 70843
rect 748 70699 788 70708
rect 652 67255 692 67264
rect 748 70580 788 70589
rect 556 64903 596 64912
rect 652 66716 692 66725
rect 556 64448 596 64457
rect 460 62936 500 62945
rect 172 61424 212 61433
rect 76 60080 116 60089
rect 76 56552 116 60040
rect 172 57224 212 61384
rect 172 57175 212 57184
rect 268 59912 308 59921
rect 268 56888 308 59872
rect 460 58232 500 62896
rect 556 58904 596 64408
rect 652 61592 692 66676
rect 748 63944 788 70540
rect 844 67976 884 75076
rect 940 74948 980 75244
rect 940 74899 980 74908
rect 1036 72680 1076 76840
rect 1132 76796 1172 80452
rect 1132 76747 1172 76756
rect 1228 76712 1268 85744
rect 1324 78056 1364 87256
rect 1420 86792 1460 89272
rect 1516 87464 1556 91792
rect 1612 91664 1652 91673
rect 1612 89732 1652 91624
rect 1612 89683 1652 89692
rect 1612 89396 1652 89405
rect 1612 89261 1652 89356
rect 1516 87415 1556 87424
rect 1612 87212 1652 87221
rect 1420 86743 1460 86752
rect 1516 87128 1556 87137
rect 1420 86120 1460 86129
rect 1420 85532 1460 86080
rect 1420 85483 1460 85492
rect 1420 85364 1460 85373
rect 1420 84776 1460 85324
rect 1420 84727 1460 84736
rect 1420 84272 1460 84281
rect 1420 82340 1460 84232
rect 1420 82291 1460 82300
rect 1420 82088 1460 82097
rect 1420 81953 1460 82048
rect 1324 78007 1364 78016
rect 1420 80828 1460 80837
rect 1228 76663 1268 76672
rect 1324 77468 1364 77477
rect 1228 76544 1268 76553
rect 1228 75956 1268 76504
rect 1132 75788 1172 75797
rect 1132 74192 1172 75748
rect 1228 74444 1268 75916
rect 1228 74395 1268 74404
rect 1132 74152 1268 74192
rect 940 72640 1076 72680
rect 940 72512 980 72640
rect 940 72463 980 72472
rect 1036 72512 1076 72521
rect 844 67927 884 67936
rect 940 72344 980 72353
rect 748 63895 788 63904
rect 844 67724 884 67733
rect 652 61543 692 61552
rect 556 58855 596 58864
rect 748 59156 788 59165
rect 460 58183 500 58192
rect 652 58400 692 58409
rect 268 56839 308 56848
rect 460 56888 500 56897
rect 76 56503 116 56512
rect 460 53864 500 56848
rect 460 53815 500 53824
rect 556 56216 596 56225
rect 556 53528 596 56176
rect 652 55208 692 58360
rect 748 55880 788 59116
rect 844 56804 884 67684
rect 940 66632 980 72304
rect 1036 68312 1076 72472
rect 1228 71672 1268 74152
rect 1228 71623 1268 71632
rect 1228 71000 1268 71009
rect 1036 68263 1076 68272
rect 1132 70916 1172 70925
rect 940 66583 980 66592
rect 940 65960 980 65969
rect 940 60584 980 65920
rect 1036 65288 1076 65297
rect 1036 61928 1076 65248
rect 1132 64280 1172 70876
rect 1228 70865 1268 70960
rect 1324 69656 1364 77428
rect 1420 76040 1460 80788
rect 1420 75991 1460 76000
rect 1420 75200 1460 75209
rect 1420 74360 1460 75160
rect 1420 74311 1460 74320
rect 1420 74192 1460 74201
rect 1420 70664 1460 74152
rect 1420 70615 1460 70624
rect 1324 69607 1364 69616
rect 1420 70496 1460 70505
rect 1228 68984 1268 68993
rect 1228 68849 1268 68944
rect 1420 68732 1460 70456
rect 1228 68692 1460 68732
rect 1228 66296 1268 68692
rect 1324 68396 1364 68405
rect 1324 68228 1364 68356
rect 1324 68179 1364 68188
rect 1228 66247 1268 66256
rect 1324 68060 1364 68069
rect 1228 65876 1268 65885
rect 1228 64616 1268 65836
rect 1228 64567 1268 64576
rect 1324 64448 1364 68020
rect 1420 67640 1460 67649
rect 1420 67505 1460 67600
rect 1420 66968 1460 66977
rect 1420 66833 1460 66928
rect 1420 66212 1460 66221
rect 1420 65624 1460 66172
rect 1420 65575 1460 65584
rect 1132 64231 1172 64240
rect 1228 64408 1364 64448
rect 1420 65372 1460 65381
rect 1228 63272 1268 64408
rect 1420 64364 1460 65332
rect 1420 63860 1460 64324
rect 1420 63811 1460 63820
rect 1228 63223 1268 63232
rect 1324 63608 1364 63617
rect 1036 61879 1076 61888
rect 940 60535 980 60544
rect 1324 60248 1364 63568
rect 1516 63356 1556 87088
rect 1612 86708 1652 87172
rect 1612 86659 1652 86668
rect 1612 86540 1652 86549
rect 1612 85028 1652 86500
rect 1612 84979 1652 84988
rect 1612 84104 1652 84113
rect 1612 83969 1652 84064
rect 1708 83540 1748 93136
rect 1900 92924 1940 93580
rect 1996 93596 2036 96688
rect 2092 94856 2132 94865
rect 2092 94721 2132 94816
rect 2188 94268 2228 96688
rect 2380 94352 2420 96688
rect 2572 95024 2612 96688
rect 2572 94975 2612 94984
rect 2476 94856 2516 94865
rect 2476 94721 2516 94816
rect 2380 94303 2420 94312
rect 2668 94436 2708 94445
rect 2188 94219 2228 94228
rect 1996 93547 2036 93556
rect 2572 93596 2612 93605
rect 2476 93512 2516 93521
rect 2284 93472 2476 93512
rect 1900 92884 2228 92924
rect 2188 92840 2228 92884
rect 2188 92791 2228 92800
rect 1996 92672 2036 92681
rect 1900 92588 1940 92597
rect 1612 83500 1748 83540
rect 1804 90908 1844 90917
rect 1612 80408 1652 83500
rect 1612 80359 1652 80368
rect 1708 83432 1748 83441
rect 1612 80240 1652 80249
rect 1612 79316 1652 80200
rect 1612 79267 1652 79276
rect 1612 78980 1652 78989
rect 1612 76964 1652 78940
rect 1612 76915 1652 76924
rect 1612 76796 1652 76805
rect 1612 75620 1652 76756
rect 1612 75571 1652 75580
rect 1612 75032 1652 75041
rect 1612 68396 1652 74992
rect 1708 73460 1748 83392
rect 1804 80576 1844 90868
rect 1900 84272 1940 92548
rect 1996 91244 2036 92632
rect 2284 91832 2324 93472
rect 2476 93463 2516 93472
rect 1996 91195 2036 91204
rect 2092 91792 2324 91832
rect 2092 90488 2132 91792
rect 1996 90448 2132 90488
rect 2188 91664 2228 91673
rect 1996 89816 2036 90448
rect 1996 89767 2036 89776
rect 2092 90320 2132 90329
rect 2092 89732 2132 90280
rect 2092 89683 2132 89692
rect 1996 89648 2036 89657
rect 1996 89513 2036 89608
rect 2092 89564 2132 89573
rect 2092 89396 2132 89524
rect 1900 84223 1940 84232
rect 1996 89356 2132 89396
rect 1900 84104 1940 84113
rect 1900 83969 1940 84064
rect 1900 83516 1940 83525
rect 1900 82676 1940 83476
rect 1900 82627 1940 82636
rect 1900 82340 1940 82435
rect 1900 82291 1940 82300
rect 1804 80527 1844 80536
rect 1900 82172 1940 82181
rect 1804 79904 1844 79913
rect 1804 79820 1844 79864
rect 1804 79769 1844 79780
rect 1804 79484 1844 79493
rect 1804 74360 1844 79444
rect 1900 78728 1940 82132
rect 1996 82004 2036 89356
rect 1996 81955 2036 81964
rect 2092 87884 2132 87893
rect 1900 78679 1940 78688
rect 1996 81080 2036 81089
rect 1804 74311 1844 74320
rect 1900 77300 1940 77309
rect 1708 73420 1844 73460
rect 1708 72512 1748 72521
rect 1708 72260 1748 72472
rect 1708 72211 1748 72220
rect 1708 72092 1748 72101
rect 1708 71957 1748 72052
rect 1708 71504 1748 71513
rect 1708 69908 1748 71464
rect 1708 69859 1748 69868
rect 1612 68347 1652 68356
rect 1708 69404 1748 69413
rect 1612 68228 1652 68237
rect 1612 66212 1652 68188
rect 1612 66163 1652 66172
rect 1324 60199 1364 60208
rect 1420 63272 1460 63312
rect 1516 63307 1556 63316
rect 1612 65960 1652 65969
rect 1420 63188 1460 63232
rect 1420 62348 1460 63148
rect 1516 63104 1556 63113
rect 1516 62768 1556 63064
rect 1516 62719 1556 62728
rect 1420 59576 1460 62308
rect 1516 62096 1556 62105
rect 1516 60752 1556 62056
rect 1612 60920 1652 65920
rect 1708 64616 1748 69364
rect 1804 68480 1844 73420
rect 1804 68431 1844 68440
rect 1804 68312 1844 68321
rect 1804 66296 1844 68272
rect 1804 66247 1844 66256
rect 1804 66128 1844 66137
rect 1804 65708 1844 66088
rect 1804 65659 1844 65668
rect 1708 64567 1748 64576
rect 1708 64448 1748 64457
rect 1708 63692 1748 64408
rect 1708 63643 1748 63652
rect 1804 64448 1844 64457
rect 1612 60871 1652 60880
rect 1708 63524 1748 63533
rect 1516 60712 1652 60752
rect 1324 59536 1460 59576
rect 1516 60584 1556 60593
rect 1324 57812 1364 59536
rect 1420 59408 1460 59417
rect 1420 59273 1460 59368
rect 1324 57763 1364 57772
rect 1420 58400 1460 58409
rect 844 56300 884 56764
rect 844 56251 884 56260
rect 1324 56888 1364 56897
rect 748 55831 788 55840
rect 652 55159 692 55168
rect 1324 54200 1364 56848
rect 1420 55544 1460 58360
rect 1516 57560 1556 60544
rect 1612 58652 1652 60712
rect 1612 58603 1652 58612
rect 1516 57511 1556 57520
rect 1420 55495 1460 55504
rect 1708 54284 1748 63484
rect 1804 59240 1844 64408
rect 1900 63524 1940 77260
rect 1996 77132 2036 81040
rect 2092 80660 2132 87844
rect 2188 86372 2228 91624
rect 2476 91664 2516 91673
rect 2380 91076 2420 91085
rect 2188 86323 2228 86332
rect 2284 90152 2324 90161
rect 2188 85784 2228 85793
rect 2188 84440 2228 85744
rect 2188 84391 2228 84400
rect 2188 84272 2228 84281
rect 2188 80828 2228 84232
rect 2188 80779 2228 80788
rect 2284 80744 2324 90112
rect 2380 86036 2420 91036
rect 2476 89648 2516 91624
rect 2572 91412 2612 93556
rect 2668 92420 2708 94396
rect 2764 94352 2804 96688
rect 2956 94772 2996 96688
rect 2956 94723 2996 94732
rect 3148 94604 3188 96688
rect 3340 95024 3380 96688
rect 3340 94975 3380 94984
rect 3148 94555 3188 94564
rect 3244 94856 3284 94865
rect 2764 94303 2804 94312
rect 2668 92371 2708 92380
rect 2764 94184 2804 94193
rect 2764 92336 2804 94144
rect 3148 94184 3188 94193
rect 2860 94100 2900 94109
rect 2860 93596 2900 94060
rect 3148 93848 3188 94144
rect 3148 93799 3188 93808
rect 2860 93547 2900 93556
rect 2956 92672 2996 92681
rect 2956 92537 2996 92632
rect 2764 92287 2804 92296
rect 3148 92336 3188 92345
rect 2572 91363 2612 91372
rect 2956 92252 2996 92261
rect 2476 89599 2516 89608
rect 2572 91160 2612 91169
rect 2476 89312 2516 89321
rect 2476 88304 2516 89272
rect 2476 88255 2516 88264
rect 2476 87968 2516 87977
rect 2476 87833 2516 87928
rect 2572 87800 2612 91120
rect 2956 90824 2996 92212
rect 2764 90784 2996 90824
rect 3052 90908 3092 90917
rect 2668 90320 2708 90329
rect 2668 89900 2708 90280
rect 2764 89984 2804 90784
rect 3052 90773 3092 90868
rect 3148 90488 3188 92296
rect 2764 89935 2804 89944
rect 2956 90448 3188 90488
rect 2668 89851 2708 89860
rect 2572 87751 2612 87760
rect 2668 89732 2708 89741
rect 2860 89732 2900 89741
rect 2668 87632 2708 89692
rect 2764 89692 2860 89732
rect 2764 88892 2804 89692
rect 2860 89664 2900 89692
rect 2860 89564 2900 89573
rect 2860 89480 2900 89524
rect 2860 89429 2900 89440
rect 2764 88052 2804 88852
rect 2956 88892 2996 90448
rect 3148 90152 3188 90161
rect 3052 89396 3092 89405
rect 3052 89261 3092 89356
rect 2956 88843 2996 88852
rect 3052 88892 3092 88901
rect 2764 88003 2804 88012
rect 2956 88724 2996 88733
rect 2764 87884 2804 87893
rect 2764 87749 2804 87844
rect 2572 87592 2708 87632
rect 2476 87464 2516 87473
rect 2476 86120 2516 87424
rect 2476 86071 2516 86080
rect 2380 85987 2420 85996
rect 2380 85868 2420 85877
rect 2380 80912 2420 85828
rect 2572 85784 2612 87592
rect 2956 87548 2996 88684
rect 2572 85735 2612 85744
rect 2668 87508 2996 87548
rect 2476 85700 2516 85709
rect 2476 82172 2516 85660
rect 2476 82123 2516 82132
rect 2572 85616 2612 85625
rect 2476 82004 2516 82015
rect 2476 81920 2516 81964
rect 2476 81871 2516 81880
rect 2380 80863 2420 80872
rect 2476 81416 2516 81425
rect 2284 80704 2420 80744
rect 2092 80620 2324 80660
rect 2092 80492 2132 80501
rect 2092 78308 2132 80452
rect 2188 80240 2228 80249
rect 2188 78980 2228 80200
rect 2188 78931 2228 78940
rect 2092 78259 2132 78268
rect 2188 78812 2228 78821
rect 1996 77092 2132 77132
rect 1996 76964 2036 76973
rect 1996 74108 2036 76924
rect 1996 74059 2036 74068
rect 1996 73940 2036 73949
rect 1996 73460 2036 73900
rect 1996 73411 2036 73420
rect 1996 73352 2036 73361
rect 1996 68396 2036 73312
rect 2092 71000 2132 77092
rect 2188 71924 2228 78772
rect 2284 77720 2324 80620
rect 2380 79148 2420 80704
rect 2380 79099 2420 79108
rect 2476 80492 2516 81376
rect 2284 77671 2324 77680
rect 2380 78308 2420 78317
rect 2284 77468 2324 77477
rect 2284 76964 2324 77428
rect 2284 76915 2324 76924
rect 2284 76796 2324 76805
rect 2284 75284 2324 76756
rect 2284 73772 2324 75244
rect 2284 73723 2324 73732
rect 2380 75956 2420 78268
rect 2476 77216 2516 80452
rect 2476 77167 2516 77176
rect 2380 75200 2420 75916
rect 2476 77048 2516 77057
rect 2476 75368 2516 77008
rect 2476 75319 2516 75328
rect 2284 73604 2324 73613
rect 2284 73352 2324 73564
rect 2380 73460 2420 75160
rect 2380 73411 2420 73420
rect 2476 74444 2516 74453
rect 2476 73772 2516 74404
rect 2284 73312 2420 73352
rect 2380 72512 2420 73312
rect 2476 72932 2516 73732
rect 2572 73100 2612 85576
rect 2668 85028 2708 87508
rect 2860 87380 2900 87389
rect 2668 84979 2708 84988
rect 2764 86792 2804 86801
rect 2764 84440 2804 86752
rect 2860 86624 2900 87340
rect 3052 87380 3092 88852
rect 3052 87331 3092 87340
rect 2860 85868 2900 86584
rect 2860 85280 2900 85828
rect 2860 85231 2900 85240
rect 2956 87296 2996 87305
rect 2956 85112 2996 87256
rect 2956 85063 2996 85072
rect 3052 87128 3092 87137
rect 2764 84391 2804 84400
rect 2860 85028 2900 85037
rect 2764 84272 2804 84281
rect 2668 84020 2708 84029
rect 2668 83885 2708 83980
rect 2764 83768 2804 84232
rect 2860 84020 2900 84988
rect 2860 83971 2900 83980
rect 2956 84860 2996 84869
rect 2764 83719 2804 83728
rect 2764 83516 2804 83525
rect 2956 83516 2996 84820
rect 3052 83684 3092 87088
rect 3052 83635 3092 83644
rect 2668 83432 2708 83441
rect 2668 81332 2708 83392
rect 2764 82928 2804 83476
rect 2764 82879 2804 82888
rect 2860 83476 2996 83516
rect 2860 82844 2900 83476
rect 3148 83432 3188 90112
rect 3244 89648 3284 94816
rect 3532 94352 3572 96688
rect 3628 94940 3668 94951
rect 3628 94856 3668 94900
rect 3628 94807 3668 94816
rect 3724 94772 3764 96688
rect 3916 95444 3956 96688
rect 4108 95780 4148 96688
rect 4108 95740 4244 95780
rect 3916 95404 4148 95444
rect 3724 94723 3764 94732
rect 4012 94856 4052 94865
rect 4012 94721 4052 94816
rect 3688 94520 4056 94529
rect 3728 94480 3770 94520
rect 3810 94480 3852 94520
rect 3892 94480 3934 94520
rect 3974 94480 4016 94520
rect 3688 94471 4056 94480
rect 3532 94303 3572 94312
rect 4108 94352 4148 95404
rect 4204 95024 4244 95740
rect 4204 94975 4244 94984
rect 4108 94303 4148 94312
rect 4300 94352 4340 96688
rect 4396 94856 4436 94865
rect 4396 94721 4436 94816
rect 4492 94772 4532 96688
rect 4588 95612 4628 95621
rect 4588 95024 4628 95572
rect 4588 94975 4628 94984
rect 4492 94723 4532 94732
rect 4300 94303 4340 94312
rect 4684 94352 4724 96688
rect 4876 95444 4916 96688
rect 4780 95404 4916 95444
rect 5068 95444 5108 96688
rect 5260 95612 5300 96688
rect 5260 95563 5300 95572
rect 5068 95404 5396 95444
rect 4780 94604 4820 95404
rect 4928 95276 5296 95285
rect 4968 95236 5010 95276
rect 5050 95236 5092 95276
rect 5132 95236 5174 95276
rect 5214 95236 5256 95276
rect 4928 95227 5296 95236
rect 4780 94555 4820 94564
rect 4684 94303 4724 94312
rect 5356 94352 5396 95404
rect 5356 94303 5396 94312
rect 5452 94268 5492 96688
rect 5644 95024 5684 96688
rect 5644 94975 5684 94984
rect 5548 94856 5588 94865
rect 5548 94721 5588 94816
rect 5836 94352 5876 96688
rect 5836 94303 5876 94312
rect 5932 94856 5972 94865
rect 5452 94219 5492 94228
rect 4588 94184 4628 94193
rect 4588 93932 4628 94144
rect 4972 94184 5012 94193
rect 4588 93883 4628 93892
rect 4684 94100 4724 94109
rect 4684 93620 4724 94060
rect 4972 94049 5012 94144
rect 5356 94184 5396 94193
rect 5356 94049 5396 94144
rect 5740 94184 5780 94193
rect 5740 94049 5780 94144
rect 4928 93764 5296 93773
rect 4968 93724 5010 93764
rect 5050 93724 5092 93764
rect 5132 93724 5174 93764
rect 5214 93724 5256 93764
rect 4928 93715 5296 93724
rect 4588 93580 4724 93620
rect 4108 93176 4148 93185
rect 3688 93008 4056 93017
rect 3728 92968 3770 93008
rect 3810 92968 3852 93008
rect 3892 92968 3934 93008
rect 3974 92968 4016 93008
rect 3688 92959 4056 92968
rect 3688 91496 4056 91505
rect 3728 91456 3770 91496
rect 3810 91456 3852 91496
rect 3892 91456 3934 91496
rect 3974 91456 4016 91496
rect 3688 91447 4056 91456
rect 3244 89599 3284 89608
rect 3340 90320 3380 90329
rect 3244 89480 3284 89489
rect 3244 89060 3284 89440
rect 3244 89011 3284 89020
rect 3244 88892 3284 88901
rect 3244 87548 3284 88852
rect 3340 88220 3380 90280
rect 3532 90320 3572 90329
rect 3340 88171 3380 88180
rect 3436 89648 3476 89657
rect 3244 87508 3380 87548
rect 3340 87296 3380 87508
rect 3340 87247 3380 87256
rect 3340 87128 3380 87137
rect 3244 86288 3284 86297
rect 3244 85196 3284 86248
rect 3244 85147 3284 85156
rect 3244 85028 3284 85037
rect 3244 84272 3284 84988
rect 3340 85028 3380 87088
rect 3436 86708 3476 89608
rect 3532 89144 3572 90280
rect 4012 90152 4052 90247
rect 4012 90103 4052 90112
rect 3688 89984 4056 89993
rect 3728 89944 3770 89984
rect 3810 89944 3852 89984
rect 3892 89944 3934 89984
rect 3974 89944 4016 89984
rect 3688 89935 4056 89944
rect 3628 89816 3668 89825
rect 3628 89681 3668 89776
rect 3820 89648 3860 89657
rect 3628 89396 3668 89405
rect 3628 89261 3668 89356
rect 3820 89228 3860 89608
rect 3820 89179 3860 89188
rect 4012 89480 4052 89489
rect 3532 89095 3572 89104
rect 3532 88976 3572 88985
rect 3532 88052 3572 88936
rect 4012 88892 4052 89440
rect 4012 88843 4052 88852
rect 3688 88472 4056 88481
rect 3728 88432 3770 88472
rect 3810 88432 3852 88472
rect 3892 88432 3934 88472
rect 3974 88432 4016 88472
rect 3688 88423 4056 88432
rect 3532 88003 3572 88012
rect 4012 88052 4052 88061
rect 3628 87296 3668 87305
rect 3628 87161 3668 87256
rect 3436 86659 3476 86668
rect 3532 87128 3572 87137
rect 3340 84979 3380 84988
rect 3244 83768 3284 84232
rect 3244 83719 3284 83728
rect 3340 84440 3380 84449
rect 3052 83392 3188 83432
rect 3244 83600 3284 83609
rect 2860 82795 2900 82804
rect 2956 83348 2996 83357
rect 2764 82676 2804 82685
rect 2764 82172 2804 82636
rect 2764 82123 2804 82132
rect 2860 82088 2900 82097
rect 2860 82004 2900 82048
rect 2668 81283 2708 81292
rect 2764 81964 2900 82004
rect 2956 82004 2996 83308
rect 2668 81080 2708 81089
rect 2668 80576 2708 81040
rect 2668 80527 2708 80536
rect 2764 80408 2804 81964
rect 2956 81955 2996 81964
rect 3052 81836 3092 83392
rect 2956 81796 3092 81836
rect 3148 83264 3188 83273
rect 3148 81920 3188 83224
rect 3244 82676 3284 83560
rect 3244 82627 3284 82636
rect 3340 83432 3380 84400
rect 3340 82844 3380 83392
rect 3436 84356 3476 84365
rect 3436 83600 3476 84316
rect 3436 82844 3476 83560
rect 3532 83012 3572 87088
rect 4012 87128 4052 88012
rect 4012 87079 4052 87088
rect 3688 86960 4056 86969
rect 3728 86920 3770 86960
rect 3810 86920 3852 86960
rect 3892 86920 3934 86960
rect 3974 86920 4016 86960
rect 3688 86911 4056 86920
rect 4012 86792 4052 86801
rect 4012 86540 4052 86752
rect 4012 86288 4052 86500
rect 4012 86239 4052 86248
rect 3688 85448 4056 85457
rect 3728 85408 3770 85448
rect 3810 85408 3852 85448
rect 3892 85408 3934 85448
rect 3974 85408 4016 85448
rect 3688 85399 4056 85408
rect 4108 85196 4148 93136
rect 4492 90572 4532 90581
rect 4012 85156 4148 85196
rect 4204 90152 4244 90161
rect 3628 84944 3668 85039
rect 3628 84895 3668 84904
rect 3628 84692 3668 84701
rect 3628 84104 3668 84652
rect 3724 84608 3764 84617
rect 3724 84356 3764 84568
rect 3724 84221 3764 84316
rect 3628 84055 3668 84064
rect 4012 84104 4052 85156
rect 4012 84055 4052 84064
rect 4108 85028 4148 85037
rect 3688 83936 4056 83945
rect 3728 83896 3770 83936
rect 3810 83896 3852 83936
rect 3892 83896 3934 83936
rect 3974 83896 4016 83936
rect 3688 83887 4056 83896
rect 3820 83768 3860 83777
rect 4108 83768 4148 84988
rect 3532 82963 3572 82972
rect 3724 83684 3764 83693
rect 3724 83516 3764 83644
rect 3436 82804 3572 82844
rect 2860 81332 2900 81341
rect 2860 80744 2900 81292
rect 2860 80695 2900 80704
rect 2668 80368 2804 80408
rect 2860 80492 2900 80501
rect 2668 79988 2708 80368
rect 2860 80324 2900 80452
rect 2668 79939 2708 79948
rect 2764 80284 2900 80324
rect 2764 79820 2804 80284
rect 2956 80240 2996 81796
rect 2956 80191 2996 80200
rect 3052 81080 3092 81089
rect 2764 79232 2804 79780
rect 2956 80072 2996 80081
rect 2956 79736 2996 80032
rect 3052 79904 3092 81040
rect 3148 80492 3188 81880
rect 3244 82508 3284 82517
rect 3244 81836 3284 82468
rect 3340 82004 3380 82804
rect 3532 82760 3572 82804
rect 3532 82088 3572 82720
rect 3724 82592 3764 83476
rect 3820 82676 3860 83728
rect 3820 82627 3860 82636
rect 3916 83728 4148 83768
rect 3724 82543 3764 82552
rect 3916 82592 3956 83728
rect 3916 82543 3956 82552
rect 4108 83600 4148 83609
rect 3688 82424 4056 82433
rect 3728 82384 3770 82424
rect 3810 82384 3852 82424
rect 3892 82384 3934 82424
rect 3974 82384 4016 82424
rect 3688 82375 4056 82384
rect 3628 82088 3668 82097
rect 3532 82048 3628 82088
rect 3628 82039 3668 82048
rect 4012 82088 4052 82097
rect 3340 81955 3380 81964
rect 3820 82004 3860 82013
rect 3724 81920 3764 81929
rect 3436 81836 3476 81845
rect 3244 81796 3380 81836
rect 3148 80443 3188 80452
rect 3244 81248 3284 81257
rect 3052 79855 3092 79864
rect 3148 79820 3188 79829
rect 2764 79183 2804 79192
rect 2860 79696 2996 79736
rect 3052 79736 3092 79745
rect 2668 79148 2708 79157
rect 2668 77132 2708 79108
rect 2860 79064 2900 79696
rect 2668 77083 2708 77092
rect 2764 79024 2900 79064
rect 2956 79568 2996 79577
rect 2764 76628 2804 79024
rect 2860 77216 2900 77225
rect 2860 76796 2900 77176
rect 2860 76747 2900 76756
rect 2956 76712 2996 79528
rect 3052 78476 3092 79696
rect 3148 79232 3188 79780
rect 3244 79484 3284 81208
rect 3340 80072 3380 81796
rect 3340 80023 3380 80032
rect 3244 79435 3284 79444
rect 3340 79904 3380 79913
rect 3148 79183 3188 79192
rect 3340 79064 3380 79864
rect 3340 79015 3380 79024
rect 3244 78980 3284 78989
rect 3244 78845 3284 78940
rect 3340 78812 3380 78821
rect 3052 78427 3092 78436
rect 3148 78728 3188 78737
rect 3148 78308 3188 78688
rect 2956 76663 2996 76672
rect 3052 78268 3188 78308
rect 2860 76628 2900 76637
rect 2764 76588 2860 76628
rect 2860 76560 2900 76588
rect 2668 76544 2708 76553
rect 2668 74444 2708 76504
rect 2956 76376 2996 76385
rect 2860 76040 2900 76049
rect 2860 75905 2900 76000
rect 2668 74395 2708 74404
rect 2764 75788 2804 75797
rect 2572 73051 2612 73060
rect 2668 74276 2708 74285
rect 2572 72932 2612 72941
rect 2476 72892 2572 72932
rect 2380 72472 2516 72512
rect 2188 71875 2228 71884
rect 2380 72008 2420 72017
rect 2092 70951 2132 70960
rect 2188 71756 2228 71765
rect 1996 68347 2036 68356
rect 2092 69656 2132 69665
rect 2092 67472 2132 69616
rect 2188 68648 2228 71716
rect 2284 71336 2324 71345
rect 2284 71201 2324 71296
rect 2188 68599 2228 68608
rect 2284 68480 2324 68489
rect 2092 67423 2132 67432
rect 2188 68396 2228 68405
rect 2092 67304 2132 67313
rect 1996 66884 2036 66979
rect 1996 66835 2036 66844
rect 1996 66716 2036 66725
rect 1996 66128 2036 66676
rect 1996 66079 2036 66088
rect 1900 63475 1940 63484
rect 1996 65960 2036 65969
rect 1900 63020 1940 63029
rect 1900 59576 1940 62980
rect 1996 61256 2036 65920
rect 2092 64112 2132 67264
rect 2092 64063 2132 64072
rect 1996 61207 2036 61216
rect 2092 63692 2132 63701
rect 1900 59527 1940 59536
rect 1996 60836 2036 60845
rect 1996 60332 2036 60796
rect 1804 59191 1844 59200
rect 1900 59324 1940 59333
rect 1804 57392 1844 57401
rect 1804 57056 1844 57352
rect 1804 57007 1844 57016
rect 1804 56888 1844 56897
rect 1804 54872 1844 56848
rect 1804 54823 1844 54832
rect 1708 54235 1748 54244
rect 1324 54151 1364 54160
rect 1708 54032 1748 54041
rect 556 53479 596 53488
rect 652 53864 692 53873
rect 556 53360 596 53369
rect 556 51848 596 53320
rect 652 52856 692 53824
rect 652 52807 692 52816
rect 1324 53192 1364 53201
rect 556 51799 596 51808
rect 652 52520 692 52529
rect 556 51596 596 51605
rect 556 51176 596 51556
rect 652 51260 692 52480
rect 652 51211 692 51220
rect 1324 51260 1364 53152
rect 1708 52604 1748 53992
rect 1900 53696 1940 59284
rect 1996 57056 2036 60292
rect 2092 59996 2132 63652
rect 2188 62012 2228 68356
rect 2284 64280 2324 68440
rect 2380 64364 2420 71968
rect 2476 71504 2516 72472
rect 2476 68816 2516 71464
rect 2572 71084 2612 72892
rect 2668 72260 2708 74236
rect 2668 72211 2708 72220
rect 2764 71420 2804 75748
rect 2860 74528 2900 74537
rect 2860 72512 2900 74488
rect 2956 73520 2996 76336
rect 3052 73688 3092 78268
rect 3148 78056 3188 78065
rect 3188 78016 3284 78056
rect 3148 78007 3188 78016
rect 3148 77720 3188 77729
rect 3148 77384 3188 77680
rect 3148 77335 3188 77344
rect 3052 73639 3092 73648
rect 3148 76628 3188 76637
rect 2956 73471 2996 73480
rect 2956 72932 2996 72941
rect 2956 72797 2996 72892
rect 2860 72463 2900 72472
rect 3052 72764 3092 72773
rect 2956 72260 2996 72269
rect 2956 72125 2996 72220
rect 2956 71756 2996 71765
rect 2764 71371 2804 71380
rect 2860 71504 2900 71513
rect 2860 71369 2900 71464
rect 2572 69908 2612 71044
rect 2764 70748 2804 70757
rect 2572 69859 2612 69868
rect 2668 70664 2708 70673
rect 2668 69152 2708 70624
rect 2764 70076 2804 70708
rect 2764 70027 2804 70036
rect 2860 69908 2900 69917
rect 2668 69103 2708 69112
rect 2764 69868 2860 69908
rect 2764 69236 2804 69868
rect 2860 69859 2900 69868
rect 2956 69908 2996 71716
rect 2956 69859 2996 69868
rect 2956 69740 2996 69749
rect 2764 69101 2804 69196
rect 2860 69152 2900 69247
rect 2860 69103 2900 69112
rect 2860 68984 2900 68993
rect 2476 68767 2516 68776
rect 2764 68944 2860 68984
rect 2476 68648 2516 68657
rect 2476 67724 2516 68608
rect 2476 67675 2516 67684
rect 2572 68228 2612 68237
rect 2476 67472 2516 67481
rect 2476 64532 2516 67432
rect 2572 66212 2612 68188
rect 2668 67724 2708 67733
rect 2764 67724 2804 68944
rect 2860 68916 2900 68944
rect 2956 68396 2996 69700
rect 3052 69236 3092 72724
rect 3052 69187 3092 69196
rect 2956 68347 2996 68356
rect 3052 69068 3092 69077
rect 2956 68144 2996 68153
rect 2860 67724 2900 67733
rect 2764 67684 2860 67724
rect 2668 66884 2708 67684
rect 2860 67656 2900 67684
rect 2956 67556 2996 68104
rect 2860 67516 2996 67556
rect 2708 66844 2804 66884
rect 2668 66835 2708 66844
rect 2572 66163 2612 66172
rect 2668 66716 2708 66725
rect 2476 64483 2516 64492
rect 2572 65792 2612 65801
rect 2572 64448 2612 65752
rect 2668 64700 2708 66676
rect 2764 65792 2804 66844
rect 2860 66296 2900 67516
rect 2860 66247 2900 66256
rect 2956 66884 2996 66893
rect 2860 66044 2900 66055
rect 2860 65960 2900 66004
rect 2860 65911 2900 65920
rect 2764 65743 2804 65752
rect 2956 65624 2996 66844
rect 3052 65876 3092 69028
rect 3052 65827 3092 65836
rect 2668 64651 2708 64660
rect 2764 65584 2956 65624
rect 2572 64408 2708 64448
rect 2380 64324 2612 64364
rect 2284 64240 2420 64280
rect 2284 64112 2324 64121
rect 2284 62348 2324 64072
rect 2380 63440 2420 64240
rect 2380 63391 2420 63400
rect 2476 64196 2516 64205
rect 2284 62308 2420 62348
rect 2188 61963 2228 61972
rect 2284 62180 2324 62189
rect 2092 59947 2132 59956
rect 2188 61508 2228 61517
rect 1996 55628 2036 57016
rect 1996 55579 2036 55588
rect 1900 53647 1940 53656
rect 1996 54788 2036 54797
rect 1708 52555 1748 52564
rect 1804 51848 1844 51857
rect 1804 51713 1844 51808
rect 1324 51211 1364 51220
rect 556 51127 596 51136
rect 1996 51008 2036 54748
rect 2188 54620 2228 61468
rect 2284 60248 2324 62140
rect 2284 60199 2324 60208
rect 2284 60080 2324 60089
rect 2284 59324 2324 60040
rect 2284 55796 2324 59284
rect 2380 58484 2420 62308
rect 2476 60500 2516 64156
rect 2572 61004 2612 64324
rect 2668 63188 2708 64408
rect 2764 63608 2804 65584
rect 2956 65575 2996 65584
rect 2860 65456 2900 65465
rect 2860 65321 2900 65416
rect 2956 65372 2996 65467
rect 2956 65323 2996 65332
rect 2956 65204 2996 65213
rect 2860 64616 2900 64625
rect 2860 63860 2900 64576
rect 2860 63776 2900 63820
rect 2860 63727 2900 63736
rect 2764 63568 2900 63608
rect 2668 61844 2708 63148
rect 2860 62852 2900 63568
rect 2668 61795 2708 61804
rect 2764 62812 2860 62852
rect 2764 62348 2804 62812
rect 2860 62803 2900 62812
rect 2860 62684 2900 62693
rect 2860 62516 2900 62644
rect 2860 62467 2900 62476
rect 2764 61676 2804 62308
rect 2956 62348 2996 65164
rect 3052 64700 3092 64795
rect 3052 64651 3092 64660
rect 3052 64448 3092 64457
rect 3052 63272 3092 64408
rect 3148 63524 3188 76588
rect 3244 73856 3284 78016
rect 3340 75956 3380 78772
rect 3436 78224 3476 81796
rect 3532 81332 3572 81341
rect 3532 80744 3572 81292
rect 3628 81248 3668 81257
rect 3628 81080 3668 81208
rect 3724 81164 3764 81880
rect 3820 81332 3860 81964
rect 4012 81953 4052 82048
rect 3820 81283 3860 81292
rect 4108 81416 4148 83560
rect 4204 82928 4244 90112
rect 4396 88976 4436 88985
rect 4396 88892 4436 88936
rect 4396 88841 4436 88852
rect 4396 88556 4436 88565
rect 4396 88136 4436 88516
rect 4396 88087 4436 88096
rect 4492 87800 4532 90532
rect 4492 86708 4532 87760
rect 4492 86659 4532 86668
rect 4396 86120 4436 86129
rect 4300 85532 4340 85541
rect 4300 84356 4340 85492
rect 4396 85448 4436 86080
rect 4396 85399 4436 85408
rect 4492 85700 4532 85709
rect 4396 85112 4436 85121
rect 4396 84977 4436 85072
rect 4492 84440 4532 85660
rect 4300 84307 4340 84316
rect 4396 84400 4532 84440
rect 4300 84188 4340 84197
rect 4300 83516 4340 84148
rect 4396 83768 4436 84400
rect 4396 83684 4436 83728
rect 4396 83635 4436 83644
rect 4492 84272 4532 84281
rect 4300 83467 4340 83476
rect 4396 83516 4436 83525
rect 4396 83348 4436 83476
rect 4396 83299 4436 83308
rect 4204 82879 4244 82888
rect 4300 83096 4340 83105
rect 4300 82844 4340 83056
rect 4108 81248 4148 81376
rect 4108 81199 4148 81208
rect 4204 82760 4244 82769
rect 3724 81115 3764 81124
rect 4204 81080 4244 82720
rect 4300 82760 4340 82804
rect 4300 82711 4340 82720
rect 4396 83096 4436 83105
rect 4300 82592 4340 82601
rect 4300 82004 4340 82552
rect 4396 82256 4436 83056
rect 4396 82207 4436 82216
rect 4396 82004 4436 82013
rect 4300 81964 4396 82004
rect 4396 81955 4436 81964
rect 3628 81031 3668 81040
rect 4108 81040 4244 81080
rect 4300 81332 4340 81341
rect 3688 80912 4056 80921
rect 3728 80872 3770 80912
rect 3810 80872 3852 80912
rect 3892 80872 3934 80912
rect 3974 80872 4016 80912
rect 3688 80863 4056 80872
rect 4012 80744 4052 80753
rect 3532 80704 3764 80744
rect 3628 80576 3668 80585
rect 3532 79736 3572 79745
rect 3532 78980 3572 79696
rect 3628 79568 3668 80536
rect 3724 79736 3764 80704
rect 3724 79687 3764 79696
rect 4012 79652 4052 80704
rect 4012 79603 4052 79612
rect 3628 79519 3668 79528
rect 3688 79400 4056 79409
rect 3728 79360 3770 79400
rect 3810 79360 3852 79400
rect 3892 79360 3934 79400
rect 3974 79360 4016 79400
rect 3688 79351 4056 79360
rect 3532 78560 3572 78940
rect 4108 78728 4148 81040
rect 4300 80492 4340 81292
rect 4108 78679 4148 78688
rect 4204 80324 4244 80333
rect 3532 78511 3572 78520
rect 3436 78175 3476 78184
rect 3532 78308 3572 78317
rect 3340 75907 3380 75916
rect 3436 77468 3476 77477
rect 3244 73807 3284 73816
rect 3340 75116 3380 75125
rect 3148 63475 3188 63484
rect 3244 73688 3284 73697
rect 3052 63223 3092 63232
rect 3148 63356 3188 63365
rect 3148 63104 3188 63316
rect 2956 62299 2996 62308
rect 3052 63064 3188 63104
rect 2572 60955 2612 60964
rect 2668 61004 2708 61013
rect 2668 60836 2708 60964
rect 2668 60787 2708 60796
rect 2668 60668 2708 60677
rect 2476 60460 2612 60500
rect 2380 58435 2420 58444
rect 2476 60332 2516 60341
rect 2476 60164 2516 60292
rect 2476 58652 2516 60124
rect 2476 57644 2516 58612
rect 2476 57595 2516 57604
rect 2572 56972 2612 60460
rect 2668 58736 2708 60628
rect 2764 60500 2804 61636
rect 2956 62180 2996 62189
rect 2956 61760 2996 62140
rect 2956 60668 2996 61720
rect 2956 60619 2996 60628
rect 3052 60500 3092 63064
rect 3148 62936 3188 62945
rect 3148 60836 3188 62896
rect 3148 60787 3188 60796
rect 2764 60460 2996 60500
rect 3052 60460 3188 60500
rect 2956 60416 2996 60460
rect 2956 60376 3092 60416
rect 2668 58687 2708 58696
rect 2764 60164 2804 60173
rect 2764 58988 2804 60124
rect 2764 58652 2804 58948
rect 2860 60080 2900 60089
rect 2860 58736 2900 60040
rect 3052 59324 3092 60376
rect 2860 58687 2900 58696
rect 2956 59284 3092 59324
rect 2764 58603 2804 58612
rect 2668 58568 2708 58577
rect 2668 57896 2708 58528
rect 2860 58484 2900 58493
rect 2668 57847 2708 57856
rect 2764 58444 2860 58484
rect 2668 57308 2708 57403
rect 2668 57259 2708 57268
rect 2572 56923 2612 56932
rect 2668 57140 2708 57149
rect 2668 56888 2708 57100
rect 2668 56839 2708 56848
rect 2284 54788 2324 55756
rect 2668 55712 2708 55721
rect 2284 54739 2324 54748
rect 2572 55628 2612 55637
rect 2572 54872 2612 55588
rect 2668 55124 2708 55672
rect 2764 55628 2804 58444
rect 2860 58416 2900 58444
rect 2956 56300 2996 59284
rect 3052 59156 3092 59165
rect 3052 57224 3092 59116
rect 3148 58400 3188 60460
rect 3148 58351 3188 58360
rect 3148 58232 3188 58241
rect 3148 57308 3188 58192
rect 3148 57259 3188 57268
rect 3052 57175 3092 57184
rect 2956 56251 2996 56260
rect 3148 56384 3188 56393
rect 3052 56132 3092 56141
rect 2764 55588 2996 55628
rect 2668 55075 2708 55084
rect 2764 55376 2804 55385
rect 2572 54788 2612 54832
rect 2572 54737 2612 54748
rect 2668 54956 2708 54965
rect 2188 54580 2420 54620
rect 2092 54116 2132 54125
rect 2092 53360 2132 54076
rect 2188 53528 2228 53537
rect 2188 53393 2228 53488
rect 2092 53311 2132 53320
rect 2380 51680 2420 54580
rect 2476 54116 2516 54125
rect 2476 52604 2516 54076
rect 2668 53192 2708 54916
rect 2764 54536 2804 55336
rect 2860 54956 2900 54965
rect 2860 54872 2900 54916
rect 2860 54821 2900 54832
rect 2764 54487 2804 54496
rect 2668 53143 2708 53152
rect 2860 53192 2900 53201
rect 2476 52555 2516 52564
rect 2860 51932 2900 53152
rect 2860 51883 2900 51892
rect 2380 51631 2420 51640
rect 2572 51848 2612 51857
rect 1996 50959 2036 50968
rect 2572 51008 2612 51808
rect 2860 51596 2900 51605
rect 2572 50873 2612 50968
rect 2764 51556 2860 51596
rect 2380 50840 2420 50849
rect 2380 50705 2420 50800
rect 2764 48824 2804 51556
rect 2860 51528 2900 51556
rect 2956 50672 2996 55588
rect 3052 54620 3092 56092
rect 3052 53444 3092 54580
rect 3052 53395 3092 53404
rect 2956 50623 2996 50632
rect 3052 53276 3092 53285
rect 1996 48152 2036 48161
rect 1996 47228 2036 48112
rect 2668 48068 2708 48077
rect 76 45800 116 45809
rect 76 45464 116 45760
rect 76 45415 116 45424
rect 76 44960 116 44969
rect 76 44792 116 44920
rect 1612 44960 1652 44969
rect 76 44743 116 44752
rect 1420 44792 1460 44801
rect 76 44288 116 44297
rect 76 44120 116 44248
rect 76 44071 116 44080
rect 1228 43784 1268 43793
rect 1036 42860 1076 42869
rect 172 41768 212 41777
rect 76 41096 116 41105
rect 76 40592 116 41056
rect 76 40543 116 40552
rect 172 40424 212 41728
rect 172 40375 212 40384
rect 460 41180 500 41189
rect 364 40088 404 40097
rect 364 38912 404 40048
rect 364 38863 404 38872
rect 460 38744 500 41140
rect 364 38704 500 38744
rect 940 39500 980 39509
rect 76 38240 116 38249
rect 76 33032 116 38200
rect 76 32983 116 32992
rect 172 35384 212 35393
rect 172 32864 212 35344
rect 172 32815 212 32824
rect 268 33368 308 33377
rect 76 32696 116 32705
rect 76 32561 116 32656
rect 172 31688 212 31697
rect 76 29672 116 29681
rect 76 25556 116 29632
rect 172 25640 212 31648
rect 268 27656 308 33328
rect 364 30596 404 38704
rect 748 38072 788 38081
rect 652 36728 692 36737
rect 652 35216 692 36688
rect 748 35888 788 38032
rect 844 37736 884 37745
rect 844 35972 884 37696
rect 844 35923 884 35932
rect 748 35839 788 35848
rect 652 35167 692 35176
rect 844 35720 884 35729
rect 844 34460 884 35680
rect 844 34411 884 34420
rect 364 30547 404 30556
rect 460 34376 500 34385
rect 460 29168 500 34336
rect 940 33140 980 39460
rect 460 29119 500 29128
rect 556 33100 980 33140
rect 1036 33140 1076 42820
rect 1228 41180 1268 43744
rect 1228 41131 1268 41140
rect 1420 41096 1460 44752
rect 1612 44456 1652 44920
rect 1612 44407 1652 44416
rect 1996 43112 2036 47188
rect 2188 47984 2228 47993
rect 2188 46724 2228 47944
rect 2668 47933 2708 48028
rect 2764 47984 2804 48784
rect 3052 48236 3092 53236
rect 2764 47935 2804 47944
rect 2956 48196 3092 48236
rect 2188 46675 2228 46684
rect 2860 47228 2900 47237
rect 2860 46556 2900 47188
rect 2284 46136 2324 46145
rect 2188 43364 2228 43373
rect 1996 43063 2036 43072
rect 2092 43280 2132 43289
rect 1804 42608 1844 42617
rect 1708 42524 1748 42533
rect 1612 41432 1652 41441
rect 1324 41056 1460 41096
rect 1516 41348 1556 41357
rect 1324 40928 1364 41056
rect 1132 40888 1364 40928
rect 1420 40928 1460 40937
rect 1132 33620 1172 40888
rect 1228 40760 1268 40769
rect 1228 39752 1268 40720
rect 1420 40508 1460 40888
rect 1516 40760 1556 41308
rect 1516 40711 1556 40720
rect 1228 39703 1268 39712
rect 1324 40468 1460 40508
rect 1516 40592 1556 40601
rect 1324 39584 1364 40468
rect 1420 40340 1460 40349
rect 1420 39752 1460 40300
rect 1420 39703 1460 39712
rect 1324 39544 1460 39584
rect 1228 39080 1268 39089
rect 1228 36728 1268 39040
rect 1324 38492 1364 38501
rect 1324 38156 1364 38452
rect 1324 38107 1364 38116
rect 1228 36679 1268 36688
rect 1420 36560 1460 39544
rect 1420 36511 1460 36520
rect 1420 36392 1460 36401
rect 1228 36056 1268 36065
rect 1228 34376 1268 36016
rect 1420 35216 1460 36352
rect 1420 35167 1460 35176
rect 1228 34327 1268 34336
rect 1324 35048 1364 35057
rect 1324 33788 1364 35008
rect 1324 33739 1364 33748
rect 1420 35048 1460 35057
rect 1132 33284 1172 33580
rect 1132 33235 1172 33244
rect 1420 33200 1460 35008
rect 1516 33704 1556 40552
rect 1612 40424 1652 41392
rect 1612 40375 1652 40384
rect 1708 40340 1748 42484
rect 1708 40291 1748 40300
rect 1804 40172 1844 42568
rect 1996 41936 2036 41945
rect 1900 41768 1940 41777
rect 1900 40676 1940 41728
rect 1900 40627 1940 40636
rect 1708 40132 1844 40172
rect 1900 40172 1940 40181
rect 1612 39668 1652 39677
rect 1612 38912 1652 39628
rect 1612 38863 1652 38872
rect 1708 39584 1748 40132
rect 1900 39920 1940 40132
rect 1900 39871 1940 39880
rect 1612 38744 1652 38753
rect 1612 36728 1652 38704
rect 1708 37484 1748 39544
rect 1708 37435 1748 37444
rect 1804 39668 1844 39677
rect 1612 36679 1652 36688
rect 1612 36560 1652 36569
rect 1612 35048 1652 36520
rect 1612 34999 1652 35008
rect 1708 36056 1748 36065
rect 1612 34712 1652 34723
rect 1612 34628 1652 34672
rect 1612 34579 1652 34588
rect 1516 33655 1556 33664
rect 1612 34040 1652 34049
rect 1420 33151 1460 33160
rect 1036 33100 1172 33140
rect 460 28328 500 28337
rect 460 28193 500 28288
rect 556 28076 596 33100
rect 940 32948 980 32957
rect 268 27607 308 27616
rect 364 28036 596 28076
rect 652 31352 692 31361
rect 172 25591 212 25600
rect 268 26648 308 26657
rect 76 25507 116 25516
rect 76 25304 116 25313
rect 76 18416 116 25264
rect 76 18367 116 18376
rect 172 22280 212 22289
rect 172 14048 212 22240
rect 268 20096 308 26608
rect 268 20047 308 20056
rect 268 19424 308 19433
rect 268 16400 308 19384
rect 364 18332 404 28036
rect 460 26984 500 26993
rect 460 20684 500 26944
rect 460 20635 500 20644
rect 556 25640 596 25649
rect 364 18283 404 18292
rect 460 19592 500 19601
rect 268 16360 404 16400
rect 172 13999 212 14008
rect 268 16232 308 16241
rect 76 13880 116 13889
rect 76 13376 116 13840
rect 76 13327 116 13336
rect 76 12872 116 12881
rect 116 12832 212 12872
rect 76 12823 116 12832
rect 172 12620 212 12832
rect 172 12571 212 12580
rect 268 10436 308 16192
rect 364 16064 404 16360
rect 364 15476 404 16024
rect 364 15427 404 15436
rect 268 10387 308 10396
rect 364 15224 404 15233
rect 172 10184 212 10193
rect 172 5564 212 10144
rect 364 9680 404 15184
rect 460 12452 500 19552
rect 556 18500 596 25600
rect 652 25220 692 31312
rect 652 25171 692 25180
rect 748 30680 788 30689
rect 556 18451 596 18460
rect 652 24632 692 24641
rect 460 12403 500 12412
rect 556 18248 596 18257
rect 556 11948 596 18208
rect 652 17744 692 24592
rect 748 23120 788 30640
rect 748 23071 788 23080
rect 844 30008 884 30017
rect 844 22280 884 29968
rect 844 22231 884 22240
rect 940 23876 980 32908
rect 1036 32108 1076 32117
rect 1036 29924 1076 32068
rect 1036 24548 1076 29884
rect 1132 28832 1172 33100
rect 1516 33116 1556 33125
rect 1420 32192 1460 32201
rect 1132 28783 1172 28792
rect 1228 32024 1268 32033
rect 1036 24499 1076 24508
rect 1132 28664 1172 28673
rect 940 21104 980 23836
rect 748 21064 980 21104
rect 1036 23960 1076 23969
rect 748 19424 788 21064
rect 940 20936 980 20945
rect 748 19375 788 19384
rect 844 19928 884 19937
rect 652 17695 692 17704
rect 748 19256 788 19265
rect 652 12956 692 12965
rect 652 12536 692 12916
rect 652 12487 692 12496
rect 748 12368 788 19216
rect 844 12536 884 19888
rect 940 13292 980 20896
rect 1036 16232 1076 23920
rect 1132 23060 1172 28624
rect 1228 25304 1268 31984
rect 1420 31436 1460 32152
rect 1420 31387 1460 31396
rect 1420 30596 1460 30605
rect 1324 29924 1364 29935
rect 1324 29840 1364 29884
rect 1324 29791 1364 29800
rect 1324 29336 1364 29345
rect 1324 28748 1364 29296
rect 1324 28699 1364 28708
rect 1324 28580 1364 28589
rect 1324 27236 1364 28540
rect 1324 27187 1364 27196
rect 1228 25255 1268 25264
rect 1324 25976 1364 25985
rect 1132 23020 1268 23060
rect 1132 22952 1172 22961
rect 1132 22448 1172 22912
rect 1132 22399 1172 22408
rect 1228 21608 1268 23020
rect 1228 21559 1268 21568
rect 1036 16183 1076 16192
rect 1132 21524 1172 21533
rect 1132 13964 1172 21484
rect 1228 20012 1268 20021
rect 1228 16988 1268 19972
rect 1324 18584 1364 25936
rect 1420 22028 1460 30556
rect 1420 21979 1460 21988
rect 1324 18535 1364 18544
rect 1420 21860 1460 21869
rect 1228 16939 1268 16948
rect 1324 15896 1364 15905
rect 1132 13915 1172 13924
rect 1228 14804 1268 14813
rect 1228 13880 1268 14764
rect 1228 13831 1268 13840
rect 940 13243 980 13252
rect 844 12487 884 12496
rect 748 12319 788 12328
rect 556 11899 596 11908
rect 748 12200 788 12209
rect 364 9631 404 9640
rect 460 11192 500 11201
rect 364 8168 404 8177
rect 172 5515 212 5524
rect 268 5816 308 5825
rect 268 5060 308 5776
rect 364 5732 404 8128
rect 460 6656 500 11152
rect 460 6607 500 6616
rect 652 10520 692 10529
rect 364 5683 404 5692
rect 556 6488 596 6497
rect 268 5011 308 5020
rect 364 4472 404 4481
rect 364 3632 404 4432
rect 556 4304 596 6448
rect 652 5648 692 10480
rect 748 7160 788 12160
rect 940 11864 980 11873
rect 748 7111 788 7120
rect 844 8504 884 8513
rect 652 5599 692 5608
rect 844 5228 884 8464
rect 940 6992 980 11824
rect 1324 11108 1364 15856
rect 1420 14048 1460 21820
rect 1516 17996 1556 33076
rect 1612 29168 1652 34000
rect 1708 33536 1748 36016
rect 1708 33487 1748 33496
rect 1804 33452 1844 39628
rect 1900 39584 1940 39593
rect 1900 39449 1940 39544
rect 1804 33403 1844 33412
rect 1900 38744 1940 38753
rect 1708 33200 1748 33209
rect 1708 33140 1748 33160
rect 1708 33100 1844 33140
rect 1708 32696 1748 32705
rect 1708 30932 1748 32656
rect 1708 30883 1748 30892
rect 1612 29119 1652 29128
rect 1708 30260 1748 30269
rect 1612 28412 1652 28507
rect 1612 28363 1652 28372
rect 1612 28160 1652 28169
rect 1612 25220 1652 28120
rect 1612 25171 1652 25180
rect 1612 24128 1652 24137
rect 1612 23372 1652 24088
rect 1612 23323 1652 23332
rect 1612 21608 1652 21703
rect 1612 21559 1652 21568
rect 1612 21356 1652 21365
rect 1612 20180 1652 21316
rect 1612 20131 1652 20140
rect 1516 17947 1556 17956
rect 1612 19340 1652 19349
rect 1612 17828 1652 19300
rect 1612 17779 1652 17788
rect 1612 16568 1652 16577
rect 1420 13999 1460 14008
rect 1516 14888 1556 14897
rect 1420 13880 1460 13889
rect 1420 13292 1460 13840
rect 1420 13040 1460 13252
rect 1420 12991 1460 13000
rect 1324 11059 1364 11068
rect 1420 12872 1460 12881
rect 1420 10100 1460 12832
rect 1516 10436 1556 14848
rect 1612 13460 1652 16528
rect 1708 16484 1748 30220
rect 1804 27824 1844 33100
rect 1900 32948 1940 38704
rect 1996 34208 2036 41896
rect 2092 37652 2132 43240
rect 2188 43280 2228 43324
rect 2188 43229 2228 43240
rect 2284 41936 2324 46096
rect 2860 45548 2900 46516
rect 2572 44876 2612 44885
rect 2284 41887 2324 41896
rect 2380 44792 2420 44801
rect 2284 41264 2324 41273
rect 2092 37603 2132 37612
rect 2188 40844 2228 40853
rect 2188 36140 2228 40804
rect 2284 40676 2324 41224
rect 2380 40844 2420 44752
rect 2476 44204 2516 44213
rect 2476 42524 2516 44164
rect 2476 42475 2516 42484
rect 2476 42020 2516 42029
rect 2476 41768 2516 41980
rect 2476 41180 2516 41728
rect 2476 41131 2516 41140
rect 2380 40795 2420 40804
rect 2572 40676 2612 44836
rect 2668 44120 2708 44129
rect 2668 41432 2708 44080
rect 2668 41383 2708 41392
rect 2764 43700 2804 43709
rect 2284 40627 2324 40636
rect 2380 40636 2612 40676
rect 2668 41180 2708 41189
rect 2284 40508 2324 40517
rect 2284 36812 2324 40468
rect 2380 36812 2420 40636
rect 2668 40592 2708 41140
rect 2668 40543 2708 40552
rect 2572 40508 2612 40517
rect 2476 40340 2516 40349
rect 2476 38996 2516 40300
rect 2476 38947 2516 38956
rect 2572 38408 2612 40468
rect 2668 40424 2708 40433
rect 2668 39752 2708 40384
rect 2668 39703 2708 39712
rect 2572 38359 2612 38368
rect 2668 39584 2708 39593
rect 2668 37316 2708 39544
rect 2764 38492 2804 43660
rect 2860 42020 2900 45508
rect 2956 42188 2996 48196
rect 3052 45632 3092 45641
rect 3052 44288 3092 45592
rect 3052 44239 3092 44248
rect 3148 43220 3188 56344
rect 3244 53444 3284 73648
rect 3340 73436 3380 75076
rect 3340 73184 3380 73396
rect 3340 73135 3380 73144
rect 3436 72932 3476 77428
rect 3532 76796 3572 78268
rect 4012 78308 4052 78317
rect 3724 78224 3764 78233
rect 3724 78089 3764 78184
rect 4012 78173 4052 78268
rect 4108 78224 4148 78233
rect 3688 77888 4056 77897
rect 3728 77848 3770 77888
rect 3810 77848 3852 77888
rect 3892 77848 3934 77888
rect 3974 77848 4016 77888
rect 3688 77839 4056 77848
rect 4108 77552 4148 78184
rect 4012 77512 4148 77552
rect 3820 77468 3860 77477
rect 3820 77333 3860 77428
rect 3532 76040 3572 76756
rect 4012 76712 4052 77512
rect 4012 76663 4052 76672
rect 3628 76628 3668 76637
rect 3628 76493 3668 76588
rect 3688 76376 4056 76385
rect 3728 76336 3770 76376
rect 3810 76336 3852 76376
rect 3892 76336 3934 76376
rect 3974 76336 4016 76376
rect 3688 76327 4056 76336
rect 3532 74528 3572 76000
rect 3628 75956 3668 75967
rect 3628 75872 3668 75916
rect 3628 75823 3668 75832
rect 4108 75032 4148 75041
rect 3688 74864 4056 74873
rect 3728 74824 3770 74864
rect 3810 74824 3852 74864
rect 3892 74824 3934 74864
rect 3974 74824 4016 74864
rect 3688 74815 4056 74824
rect 3532 74479 3572 74488
rect 3916 74528 3956 74537
rect 3532 74360 3572 74369
rect 3532 73856 3572 74320
rect 3916 74192 3956 74488
rect 3916 74143 3956 74152
rect 4012 74444 4052 74453
rect 3532 73721 3572 73816
rect 4012 73688 4052 74404
rect 4012 73639 4052 73648
rect 3688 73352 4056 73361
rect 3728 73312 3770 73352
rect 3810 73312 3852 73352
rect 3892 73312 3934 73352
rect 3974 73312 4016 73352
rect 3688 73303 4056 73312
rect 3340 72892 3476 72932
rect 3340 72428 3380 72892
rect 3340 72379 3380 72388
rect 3436 72764 3476 72773
rect 3340 72260 3380 72269
rect 3340 71504 3380 72220
rect 3340 69236 3380 71464
rect 3436 70748 3476 72724
rect 3436 70699 3476 70708
rect 3532 72344 3572 72353
rect 3340 69187 3380 69196
rect 3436 70496 3476 70505
rect 3340 69068 3380 69077
rect 3436 69068 3476 70456
rect 3380 69028 3476 69068
rect 3340 68144 3380 69028
rect 3340 68095 3380 68104
rect 3436 68816 3476 68825
rect 3340 67640 3380 67649
rect 3340 66296 3380 67600
rect 3340 66247 3380 66256
rect 3340 66128 3380 66137
rect 3340 65204 3380 66088
rect 3340 65155 3380 65164
rect 3340 64784 3380 64793
rect 3340 64700 3380 64744
rect 3340 64649 3380 64660
rect 3340 64028 3380 64037
rect 3340 61676 3380 63988
rect 3436 63440 3476 68776
rect 3532 65456 3572 72304
rect 3628 72176 3668 72187
rect 3628 72092 3668 72136
rect 3628 72043 3668 72052
rect 3688 71840 4056 71849
rect 3728 71800 3770 71840
rect 3810 71800 3852 71840
rect 3892 71800 3934 71840
rect 3974 71800 4016 71840
rect 3688 71791 4056 71800
rect 3628 71672 3668 71681
rect 3628 70496 3668 71632
rect 3820 71420 3860 71429
rect 3724 71336 3764 71345
rect 3724 70664 3764 71296
rect 3820 71252 3860 71380
rect 4108 71420 4148 74992
rect 4204 72344 4244 80284
rect 4300 79148 4340 80452
rect 4300 79099 4340 79108
rect 4396 81248 4436 81257
rect 4396 79904 4436 81208
rect 4300 78980 4340 78989
rect 4300 77468 4340 78940
rect 4396 78560 4436 79864
rect 4396 78511 4436 78520
rect 4300 77419 4340 77428
rect 4396 78308 4436 78317
rect 4396 76796 4436 78268
rect 4492 77048 4532 84232
rect 4588 78308 4628 93580
rect 4780 93260 4820 93269
rect 4684 90824 4724 90833
rect 4684 89564 4724 90784
rect 4684 88976 4724 89524
rect 4684 88927 4724 88936
rect 4780 88808 4820 93220
rect 4928 92252 5296 92261
rect 4968 92212 5010 92252
rect 5050 92212 5092 92252
rect 5132 92212 5174 92252
rect 5214 92212 5256 92252
rect 4928 92203 5296 92212
rect 5932 92084 5972 94816
rect 6028 94772 6068 96688
rect 6028 94723 6068 94732
rect 6220 94352 6260 96688
rect 6412 95024 6452 96688
rect 6412 94975 6452 94984
rect 6316 94856 6356 94865
rect 6316 94721 6356 94816
rect 6220 94303 6260 94312
rect 6604 94352 6644 96688
rect 6700 94856 6740 94865
rect 6700 94721 6740 94816
rect 6796 94772 6836 96688
rect 6796 94723 6836 94732
rect 6604 94303 6644 94312
rect 6988 94352 7028 96688
rect 7084 94856 7124 94865
rect 7084 94721 7124 94816
rect 7180 94688 7220 96688
rect 7180 94639 7220 94648
rect 6988 94303 7028 94312
rect 7372 94352 7412 96688
rect 7564 95024 7604 96688
rect 7564 94975 7604 94984
rect 7372 94303 7412 94312
rect 7564 94772 7604 94781
rect 6124 94184 6164 94193
rect 6124 94049 6164 94144
rect 6892 94184 6932 94193
rect 6028 93680 6068 93689
rect 6028 93620 6068 93640
rect 6028 93580 6164 93620
rect 5932 92035 5972 92044
rect 6028 90824 6068 90833
rect 4928 90740 5296 90749
rect 4968 90700 5010 90740
rect 5050 90700 5092 90740
rect 5132 90700 5174 90740
rect 5214 90700 5256 90740
rect 4928 90691 5296 90700
rect 5740 90152 5780 90161
rect 4928 89228 5296 89237
rect 4968 89188 5010 89228
rect 5050 89188 5092 89228
rect 5132 89188 5174 89228
rect 5214 89188 5256 89228
rect 4928 89179 5296 89188
rect 4684 88768 4820 88808
rect 5356 89060 5396 89069
rect 4684 84524 4724 88768
rect 4780 88640 4820 88649
rect 4780 87380 4820 88600
rect 5356 88052 5396 89020
rect 5356 88003 5396 88012
rect 5452 88136 5492 88145
rect 5356 87884 5396 87893
rect 4928 87716 5296 87725
rect 4968 87676 5010 87716
rect 5050 87676 5092 87716
rect 5132 87676 5174 87716
rect 5214 87676 5256 87716
rect 4928 87667 5296 87676
rect 4780 87331 4820 87340
rect 5164 87380 5204 87389
rect 5164 86624 5204 87340
rect 5164 86489 5204 86584
rect 5260 87212 5300 87221
rect 5260 86540 5300 87172
rect 5260 86491 5300 86500
rect 4780 86288 4820 86297
rect 4780 85868 4820 86248
rect 4928 86204 5296 86213
rect 4968 86164 5010 86204
rect 5050 86164 5092 86204
rect 5132 86164 5174 86204
rect 5214 86164 5256 86204
rect 4928 86155 5296 86164
rect 4780 85819 4820 85828
rect 4684 84475 4724 84484
rect 4780 85196 4820 85205
rect 4684 84356 4724 84365
rect 4684 83096 4724 84316
rect 4780 83516 4820 85156
rect 4928 84692 5296 84701
rect 4968 84652 5010 84692
rect 5050 84652 5092 84692
rect 5132 84652 5174 84692
rect 5214 84652 5256 84692
rect 4928 84643 5296 84652
rect 4780 83467 4820 83476
rect 5260 83768 5300 83777
rect 4684 83047 4724 83056
rect 4780 83348 4820 83357
rect 5260 83348 5300 83728
rect 5356 83516 5396 87844
rect 5452 87380 5492 88096
rect 5644 88052 5684 88061
rect 5548 87968 5588 87977
rect 5548 87464 5588 87928
rect 5548 87415 5588 87424
rect 5452 87331 5492 87340
rect 5644 87296 5684 88012
rect 5452 87128 5492 87137
rect 5452 86372 5492 87088
rect 5644 86960 5684 87256
rect 5740 87128 5780 90112
rect 5740 87079 5780 87088
rect 5836 88052 5876 88061
rect 5836 87380 5876 88012
rect 5644 86920 5780 86960
rect 5644 86792 5684 86801
rect 5452 85280 5492 86332
rect 5452 85231 5492 85240
rect 5548 86708 5588 86717
rect 5452 85112 5492 85121
rect 5452 83540 5492 85072
rect 5548 85028 5588 86668
rect 5644 86657 5684 86752
rect 5548 84979 5588 84988
rect 5644 86540 5684 86549
rect 5548 84524 5588 84533
rect 5548 84389 5588 84484
rect 5644 84440 5684 86500
rect 5644 84391 5684 84400
rect 5740 84524 5780 86920
rect 5836 86708 5876 87340
rect 5836 86659 5876 86668
rect 5932 87884 5972 87893
rect 5836 86540 5876 86549
rect 5836 86036 5876 86500
rect 5836 85987 5876 85996
rect 5740 84389 5780 84484
rect 5836 84356 5876 84365
rect 5644 84188 5684 84197
rect 5452 83500 5588 83540
rect 5356 83467 5396 83476
rect 5548 83432 5588 83500
rect 5452 83392 5588 83432
rect 5644 83432 5684 84148
rect 5836 83516 5876 84316
rect 5836 83467 5876 83476
rect 5644 83392 5780 83432
rect 5260 83308 5396 83348
rect 4684 82928 4724 82937
rect 4684 81500 4724 82888
rect 4684 80996 4724 81460
rect 4684 80947 4724 80956
rect 4780 82088 4820 83308
rect 4928 83180 5296 83189
rect 4968 83140 5010 83180
rect 5050 83140 5092 83180
rect 5132 83140 5174 83180
rect 5214 83140 5256 83180
rect 4928 83131 5296 83140
rect 4972 83012 5012 83021
rect 4972 82877 5012 82972
rect 4588 78259 4628 78268
rect 4684 80240 4724 80249
rect 4492 76999 4532 77008
rect 4588 77300 4628 77309
rect 4300 76628 4340 76637
rect 4300 76040 4340 76588
rect 4300 74780 4340 76000
rect 4300 74731 4340 74740
rect 4396 75956 4436 76756
rect 4396 74444 4436 75916
rect 4396 74395 4436 74404
rect 4492 76544 4532 76553
rect 4396 74024 4436 74033
rect 4300 73940 4340 73949
rect 4300 73772 4340 73900
rect 4396 73940 4436 73984
rect 4396 73889 4436 73900
rect 4300 73688 4340 73732
rect 4300 73639 4340 73648
rect 4204 72295 4244 72304
rect 4300 73520 4340 73529
rect 4300 72260 4340 73480
rect 4300 72211 4340 72220
rect 4396 72764 4436 72773
rect 4108 71371 4148 71380
rect 4204 72176 4244 72185
rect 4204 71252 4244 72136
rect 3820 71212 4244 71252
rect 3724 70615 3764 70624
rect 3916 70664 3956 70673
rect 3628 70447 3668 70456
rect 3916 70496 3956 70624
rect 3916 70447 3956 70456
rect 4108 70580 4148 70589
rect 3688 70328 4056 70337
rect 3728 70288 3770 70328
rect 3810 70288 3852 70328
rect 3892 70288 3934 70328
rect 3974 70288 4016 70328
rect 3688 70279 4056 70288
rect 4012 69824 4052 69833
rect 3628 69236 3668 69245
rect 3628 69101 3668 69196
rect 4012 69236 4052 69784
rect 4012 69187 4052 69196
rect 3688 68816 4056 68825
rect 3728 68776 3770 68816
rect 3810 68776 3852 68816
rect 3892 68776 3934 68816
rect 3974 68776 4016 68816
rect 3688 68767 4056 68776
rect 4012 68480 4052 68489
rect 3916 68396 3956 68407
rect 3916 68312 3956 68356
rect 3916 67808 3956 68272
rect 3916 67759 3956 67768
rect 4012 67472 4052 68440
rect 4108 67892 4148 70540
rect 4204 68312 4244 71212
rect 4396 70832 4436 72724
rect 4396 70783 4436 70792
rect 4300 70664 4340 70759
rect 4300 70615 4340 70624
rect 4300 70496 4340 70505
rect 4300 69236 4340 70456
rect 4492 70244 4532 76504
rect 4588 73772 4628 77260
rect 4684 76796 4724 80200
rect 4780 76964 4820 82048
rect 4876 82676 4916 82685
rect 4876 82004 4916 82636
rect 4876 81955 4916 81964
rect 5356 82004 5396 83308
rect 5356 81955 5396 81964
rect 4972 81836 5012 81931
rect 4972 81787 5012 81796
rect 4928 81668 5296 81677
rect 4968 81628 5010 81668
rect 5050 81628 5092 81668
rect 5132 81628 5174 81668
rect 5214 81628 5256 81668
rect 4928 81619 5296 81628
rect 5164 81500 5204 81509
rect 4972 81332 5012 81343
rect 4972 81248 5012 81292
rect 4972 81199 5012 81208
rect 5164 80324 5204 81460
rect 5356 81332 5396 81341
rect 5356 81197 5396 81292
rect 5452 80492 5492 83392
rect 5164 80275 5204 80284
rect 5356 80452 5492 80492
rect 5548 83264 5588 83273
rect 4928 80156 5296 80165
rect 4968 80116 5010 80156
rect 5050 80116 5092 80156
rect 5132 80116 5174 80156
rect 5214 80116 5256 80156
rect 4928 80107 5296 80116
rect 5260 79988 5300 79997
rect 5260 79568 5300 79948
rect 5260 79519 5300 79528
rect 4928 78644 5296 78653
rect 4968 78604 5010 78644
rect 5050 78604 5092 78644
rect 5132 78604 5174 78644
rect 5214 78604 5256 78644
rect 4928 78595 5296 78604
rect 5260 78224 5300 78233
rect 5260 77468 5300 78184
rect 5356 77552 5396 80452
rect 5452 79904 5492 79913
rect 5452 79148 5492 79864
rect 5452 79099 5492 79108
rect 5356 77503 5396 77512
rect 5452 78980 5492 78989
rect 5260 77419 5300 77428
rect 5356 77300 5396 77309
rect 4928 77132 5296 77141
rect 4968 77092 5010 77132
rect 5050 77092 5092 77132
rect 5132 77092 5174 77132
rect 5214 77092 5256 77132
rect 4928 77083 5296 77092
rect 4780 76915 4820 76924
rect 4684 76747 4724 76756
rect 5068 76796 5108 76805
rect 4684 76628 4724 76637
rect 4684 75788 4724 76588
rect 5068 75956 5108 76756
rect 5356 76796 5396 77260
rect 5356 76747 5396 76756
rect 5452 76376 5492 78940
rect 5452 76327 5492 76336
rect 5548 76208 5588 83224
rect 5356 76168 5588 76208
rect 5644 83180 5684 83189
rect 5068 75907 5108 75916
rect 5260 75956 5300 75965
rect 5260 75821 5300 75916
rect 4684 75739 4724 75748
rect 4588 73723 4628 73732
rect 4684 75620 4724 75629
rect 4684 75200 4724 75580
rect 4928 75620 5296 75629
rect 4968 75580 5010 75620
rect 5050 75580 5092 75620
rect 5132 75580 5174 75620
rect 5214 75580 5256 75620
rect 4928 75571 5296 75580
rect 4876 75284 4916 75379
rect 4876 75235 4916 75244
rect 4588 72176 4628 72185
rect 4588 72041 4628 72136
rect 4300 69187 4340 69196
rect 4396 70204 4532 70244
rect 4588 71504 4628 71513
rect 4300 68312 4340 68321
rect 4204 68272 4300 68312
rect 4108 67843 4148 67852
rect 4204 68144 4244 68153
rect 4012 67423 4052 67432
rect 4108 67724 4148 67733
rect 3688 67304 4056 67313
rect 3728 67264 3770 67304
rect 3810 67264 3852 67304
rect 3892 67264 3934 67304
rect 3974 67264 4016 67304
rect 3688 67255 4056 67264
rect 3628 67052 3668 67061
rect 3628 66212 3668 67012
rect 4108 66968 4148 67684
rect 3628 66128 3668 66172
rect 3628 66079 3668 66088
rect 3820 66800 3860 66809
rect 3820 66212 3860 66760
rect 3820 66077 3860 66172
rect 3688 65792 4056 65801
rect 3728 65752 3770 65792
rect 3810 65752 3852 65792
rect 3892 65752 3934 65792
rect 3974 65752 4016 65792
rect 3688 65743 4056 65752
rect 3532 65407 3572 65416
rect 4012 65624 4052 65633
rect 4012 65372 4052 65584
rect 4012 65323 4052 65332
rect 3436 63391 3476 63400
rect 3532 65204 3572 65213
rect 3340 61627 3380 61636
rect 3436 63272 3476 63281
rect 3436 61508 3476 63232
rect 3532 61676 3572 65164
rect 3628 65204 3668 65213
rect 3628 64616 3668 65164
rect 4012 65120 4052 65129
rect 3820 64952 3860 64961
rect 3820 64700 3860 64912
rect 3820 64651 3860 64660
rect 3628 64567 3668 64576
rect 4012 64448 4052 65080
rect 4012 64399 4052 64408
rect 3688 64280 4056 64289
rect 3728 64240 3770 64280
rect 3810 64240 3852 64280
rect 3892 64240 3934 64280
rect 3974 64240 4016 64280
rect 3688 64231 4056 64240
rect 4012 64028 4052 64037
rect 3916 63860 3956 63869
rect 3916 63188 3956 63820
rect 3916 63139 3956 63148
rect 4012 63020 4052 63988
rect 4012 62971 4052 62980
rect 3688 62768 4056 62777
rect 3728 62728 3770 62768
rect 3810 62728 3852 62768
rect 3892 62728 3934 62768
rect 3974 62728 4016 62768
rect 3688 62719 4056 62728
rect 3532 61627 3572 61636
rect 3628 62348 3668 62357
rect 3340 61468 3476 61508
rect 3340 60164 3380 61468
rect 3532 61424 3572 61433
rect 3340 58652 3380 60124
rect 3436 60920 3476 60929
rect 3436 59576 3476 60880
rect 3532 60164 3572 61384
rect 3628 61424 3668 62308
rect 4012 62348 4052 62357
rect 4012 62213 4052 62308
rect 4012 61592 4052 61601
rect 4012 61457 4052 61552
rect 3628 61375 3668 61384
rect 3688 61256 4056 61265
rect 3728 61216 3770 61256
rect 3810 61216 3852 61256
rect 3892 61216 3934 61256
rect 3974 61216 4016 61256
rect 3688 61207 4056 61216
rect 3532 60115 3572 60124
rect 3628 61088 3668 61097
rect 3628 59912 3668 61048
rect 3820 61088 3860 61097
rect 3724 61004 3764 61013
rect 3724 59996 3764 60964
rect 3820 60836 3860 61048
rect 4012 60920 4052 61015
rect 4012 60871 4052 60880
rect 3820 60500 3860 60796
rect 3916 60752 3956 60761
rect 3916 60617 3956 60712
rect 4012 60668 4052 60677
rect 3820 60460 3956 60500
rect 3724 59947 3764 59956
rect 3916 60332 3956 60460
rect 3916 59996 3956 60292
rect 3916 59947 3956 59956
rect 4012 60164 4052 60628
rect 4012 59996 4052 60124
rect 4012 59947 4052 59956
rect 3436 59527 3476 59536
rect 3532 59872 3668 59912
rect 3340 58603 3380 58612
rect 3436 59324 3476 59333
rect 3436 58736 3476 59284
rect 3244 53395 3284 53404
rect 3340 58400 3380 58409
rect 3244 51932 3284 51941
rect 3244 48152 3284 51892
rect 3340 49664 3380 58360
rect 3436 57896 3476 58696
rect 3532 58484 3572 59872
rect 3688 59744 4056 59753
rect 3728 59704 3770 59744
rect 3810 59704 3852 59744
rect 3892 59704 3934 59744
rect 3974 59704 4016 59744
rect 3688 59695 4056 59704
rect 3628 59576 3668 59585
rect 3628 59441 3668 59536
rect 3724 59492 3764 59501
rect 3724 58484 3764 59452
rect 3916 59408 3956 59417
rect 3820 59240 3860 59249
rect 3820 58652 3860 59200
rect 3916 58820 3956 59368
rect 3916 58771 3956 58780
rect 3820 58603 3860 58612
rect 3916 58568 3956 58577
rect 3916 58484 3956 58528
rect 3724 58444 3956 58484
rect 3532 58435 3572 58444
rect 3436 57140 3476 57856
rect 3436 57091 3476 57100
rect 3532 58316 3572 58325
rect 3436 56888 3476 56897
rect 3436 55796 3476 56848
rect 3436 55747 3476 55756
rect 3532 54788 3572 58276
rect 3688 58232 4056 58241
rect 3728 58192 3770 58232
rect 3810 58192 3852 58232
rect 3892 58192 3934 58232
rect 3974 58192 4016 58232
rect 3688 58183 4056 58192
rect 4012 57812 4052 57821
rect 4012 57677 4052 57772
rect 3628 57644 3668 57653
rect 3628 56888 3668 57604
rect 3628 56839 3668 56848
rect 3688 56720 4056 56729
rect 3728 56680 3770 56720
rect 3810 56680 3852 56720
rect 3892 56680 3934 56720
rect 3974 56680 4016 56720
rect 3688 56671 4056 56680
rect 3628 56552 3668 56561
rect 3628 56300 3668 56512
rect 3628 56251 3668 56260
rect 3688 55208 4056 55217
rect 3728 55168 3770 55208
rect 3810 55168 3852 55208
rect 3892 55168 3934 55208
rect 3974 55168 4016 55208
rect 3688 55159 4056 55168
rect 3436 54748 3572 54788
rect 3724 54872 3764 54881
rect 3436 53612 3476 54748
rect 3628 54704 3668 54713
rect 3532 54620 3572 54629
rect 3532 54368 3572 54580
rect 3532 54319 3572 54328
rect 3628 54116 3668 54664
rect 3724 54200 3764 54832
rect 3820 54704 3860 54713
rect 3820 54284 3860 54664
rect 3820 54235 3860 54244
rect 3916 54704 3956 54713
rect 3916 54536 3956 54664
rect 3724 54151 3764 54160
rect 3628 54067 3668 54076
rect 3916 54032 3956 54496
rect 3916 53983 3956 53992
rect 3724 53864 3764 53959
rect 3724 53815 3764 53824
rect 3688 53696 4056 53705
rect 3728 53656 3770 53696
rect 3810 53656 3852 53696
rect 3892 53656 3934 53696
rect 3974 53656 4016 53696
rect 3688 53647 4056 53656
rect 3436 53572 3572 53612
rect 3436 53444 3476 53453
rect 3436 51764 3476 53404
rect 3532 53360 3572 53572
rect 3532 53311 3572 53320
rect 4012 53276 4052 53285
rect 4108 53276 4148 66928
rect 4204 66884 4244 68104
rect 4204 66835 4244 66844
rect 4300 67556 4340 68272
rect 4396 67556 4436 70204
rect 4492 70076 4532 70085
rect 4492 67724 4532 70036
rect 4588 69908 4628 71464
rect 4684 70076 4724 75160
rect 4876 75116 4916 75125
rect 4684 70027 4724 70036
rect 4780 74444 4820 74453
rect 4588 69868 4724 69908
rect 4492 67675 4532 67684
rect 4588 69740 4628 69749
rect 4588 67724 4628 69700
rect 4684 68984 4724 69868
rect 4780 69068 4820 74404
rect 4876 74276 4916 75076
rect 5260 74696 5300 74705
rect 5068 74612 5108 74621
rect 5068 74444 5108 74572
rect 5260 74561 5300 74656
rect 5068 74395 5108 74404
rect 4876 74227 4916 74236
rect 5164 74360 5204 74371
rect 5164 74276 5204 74320
rect 5164 74227 5204 74236
rect 4928 74108 5296 74117
rect 4968 74068 5010 74108
rect 5050 74068 5092 74108
rect 5132 74068 5174 74108
rect 5214 74068 5256 74108
rect 4928 74059 5296 74068
rect 5356 73856 5396 76168
rect 5548 76040 5588 76049
rect 5356 73807 5396 73816
rect 5452 75788 5492 75797
rect 5164 73772 5204 73781
rect 4972 73688 5012 73697
rect 4972 72932 5012 73648
rect 5164 73460 5204 73732
rect 5164 73420 5396 73460
rect 4972 72883 5012 72892
rect 5260 73352 5300 73361
rect 5260 72764 5300 73312
rect 5260 72715 5300 72724
rect 4928 72596 5296 72605
rect 4968 72556 5010 72596
rect 5050 72556 5092 72596
rect 5132 72556 5174 72596
rect 5214 72556 5256 72596
rect 4928 72547 5296 72556
rect 5356 72344 5396 73420
rect 5068 72304 5396 72344
rect 5068 71504 5108 72304
rect 5164 72176 5204 72185
rect 5204 72136 5396 72176
rect 5164 72127 5204 72136
rect 5068 71455 5108 71464
rect 5260 71504 5300 71513
rect 5260 71369 5300 71464
rect 4928 71084 5296 71093
rect 4968 71044 5010 71084
rect 5050 71044 5092 71084
rect 5132 71044 5174 71084
rect 5214 71044 5256 71084
rect 4928 71035 5296 71044
rect 4972 70916 5012 70925
rect 4876 70748 4916 70757
rect 4876 70613 4916 70708
rect 4876 70412 4916 70421
rect 4876 69824 4916 70372
rect 4972 69908 5012 70876
rect 4972 69859 5012 69868
rect 5164 70916 5204 70925
rect 4876 69775 4916 69784
rect 5164 69740 5204 70876
rect 5164 69691 5204 69700
rect 4928 69572 5296 69581
rect 4968 69532 5010 69572
rect 5050 69532 5092 69572
rect 5132 69532 5174 69572
rect 5214 69532 5256 69572
rect 4928 69523 5296 69532
rect 5260 69404 5300 69413
rect 5260 69236 5300 69364
rect 5260 69187 5300 69196
rect 4780 69028 4916 69068
rect 4684 68944 4820 68984
rect 4588 67675 4628 67684
rect 4684 68816 4724 68825
rect 4396 67516 4628 67556
rect 4204 66716 4244 66725
rect 4204 66212 4244 66676
rect 4204 66163 4244 66172
rect 4300 65624 4340 67516
rect 4204 65584 4340 65624
rect 4396 67052 4436 67061
rect 4204 63944 4244 65584
rect 4300 65456 4340 65465
rect 4300 64868 4340 65416
rect 4300 64819 4340 64828
rect 4300 64616 4340 64625
rect 4300 64532 4340 64576
rect 4300 64481 4340 64492
rect 4204 63895 4244 63904
rect 4300 64364 4340 64373
rect 4300 63860 4340 64324
rect 4300 63811 4340 63820
rect 4204 63776 4244 63785
rect 4204 62768 4244 63736
rect 4204 62719 4244 62728
rect 4300 63608 4340 63617
rect 4204 62432 4244 62441
rect 4204 61676 4244 62392
rect 4204 57896 4244 61636
rect 4204 56384 4244 57856
rect 4204 56335 4244 56344
rect 4204 55880 4244 55889
rect 4204 54872 4244 55840
rect 4204 54823 4244 54832
rect 4204 54620 4244 54629
rect 4204 54116 4244 54580
rect 4204 54067 4244 54076
rect 4052 53236 4148 53276
rect 4012 53227 4052 53236
rect 4108 53108 4148 53236
rect 4204 53948 4244 53957
rect 4204 53276 4244 53908
rect 4204 53227 4244 53236
rect 4108 53068 4244 53108
rect 4108 52604 4148 52613
rect 3688 52184 4056 52193
rect 3728 52144 3770 52184
rect 3810 52144 3852 52184
rect 3892 52144 3934 52184
rect 3974 52144 4016 52184
rect 3688 52135 4056 52144
rect 3628 51764 3668 51773
rect 3436 51724 3628 51764
rect 3628 51715 3668 51724
rect 4108 51092 4148 52564
rect 4108 51043 4148 51052
rect 3688 50672 4056 50681
rect 3728 50632 3770 50672
rect 3810 50632 3852 50672
rect 3892 50632 3934 50672
rect 3974 50632 4016 50672
rect 3688 50623 4056 50632
rect 3340 49615 3380 49624
rect 3532 50084 3572 50093
rect 3244 47396 3284 48112
rect 3340 48068 3380 48077
rect 3340 47480 3380 48028
rect 3340 47431 3380 47440
rect 3244 47347 3284 47356
rect 3532 47312 3572 50044
rect 4108 49412 4148 49421
rect 3688 49160 4056 49169
rect 3728 49120 3770 49160
rect 3810 49120 3852 49160
rect 3892 49120 3934 49160
rect 3974 49120 4016 49160
rect 3688 49111 4056 49120
rect 4108 48068 4148 49372
rect 4204 48908 4244 53068
rect 4300 50252 4340 63568
rect 4396 63272 4436 67012
rect 4492 66296 4532 66305
rect 4492 64952 4532 66256
rect 4492 64903 4532 64912
rect 4492 64784 4532 64793
rect 4492 63440 4532 64744
rect 4492 63391 4532 63400
rect 4396 63232 4532 63272
rect 4396 63104 4436 63113
rect 4396 60332 4436 63064
rect 4492 62348 4532 63232
rect 4492 61676 4532 62308
rect 4492 61627 4532 61636
rect 4588 61592 4628 67516
rect 4684 64700 4724 68776
rect 4780 67892 4820 68944
rect 4876 68816 4916 69028
rect 4876 68767 4916 68776
rect 4972 68648 5012 68657
rect 4972 68228 5012 68608
rect 4972 68179 5012 68188
rect 4928 68060 5296 68069
rect 4968 68020 5010 68060
rect 5050 68020 5092 68060
rect 5132 68020 5174 68060
rect 5214 68020 5256 68060
rect 4928 68011 5296 68020
rect 4780 67852 5012 67892
rect 4876 67724 4916 67733
rect 4780 67640 4820 67649
rect 4780 66380 4820 67600
rect 4876 67556 4916 67684
rect 4876 67507 4916 67516
rect 4972 67052 5012 67852
rect 5356 67808 5396 72136
rect 5356 67759 5396 67768
rect 4972 67003 5012 67012
rect 4876 66968 4916 66977
rect 4876 66884 4916 66928
rect 4876 66833 4916 66844
rect 4928 66548 5296 66557
rect 4968 66508 5010 66548
rect 5050 66508 5092 66548
rect 5132 66508 5174 66548
rect 5214 66508 5256 66548
rect 4928 66499 5296 66508
rect 5356 66548 5396 66557
rect 4780 66331 4820 66340
rect 5356 66296 5396 66508
rect 5356 66247 5396 66256
rect 5356 65960 5396 65969
rect 5356 65792 5396 65920
rect 5356 65743 5396 65752
rect 5164 65372 5204 65381
rect 5164 65237 5204 65332
rect 4928 65036 5296 65045
rect 4968 64996 5010 65036
rect 5050 64996 5092 65036
rect 5132 64996 5174 65036
rect 5214 64996 5256 65036
rect 4928 64987 5296 64996
rect 4684 64651 4724 64660
rect 4876 64616 4916 64627
rect 4876 64532 4916 64576
rect 4876 64483 4916 64492
rect 5068 64280 5108 64289
rect 4780 64112 4820 64121
rect 4684 64072 4780 64112
rect 4684 63524 4724 64072
rect 4780 63977 4820 64072
rect 5068 63944 5108 64240
rect 5068 63895 5108 63904
rect 4684 63475 4724 63484
rect 4780 63692 4820 63701
rect 4588 61543 4628 61552
rect 4684 63188 4724 63197
rect 4588 61424 4628 61433
rect 4588 60836 4628 61384
rect 4396 59324 4436 60292
rect 4396 59275 4436 59284
rect 4492 60796 4588 60836
rect 4396 59156 4436 59165
rect 4396 53300 4436 59116
rect 4492 56300 4532 60796
rect 4588 60787 4628 60796
rect 4588 60668 4628 60677
rect 4588 57056 4628 60628
rect 4588 57007 4628 57016
rect 4492 55880 4532 56260
rect 4492 55831 4532 55840
rect 4492 54788 4532 54797
rect 4492 54116 4532 54748
rect 4492 54032 4532 54076
rect 4492 53952 4532 53992
rect 4396 53260 4532 53300
rect 4396 53108 4436 53117
rect 4396 51848 4436 53068
rect 4396 51799 4436 51808
rect 4492 51680 4532 53260
rect 4684 52520 4724 63148
rect 4780 63188 4820 63652
rect 5356 63692 5396 63701
rect 4928 63524 5296 63533
rect 4968 63484 5010 63524
rect 5050 63484 5092 63524
rect 5132 63484 5174 63524
rect 5214 63484 5256 63524
rect 4928 63475 5296 63484
rect 4780 63139 4820 63148
rect 5260 63356 5300 63365
rect 4972 63020 5012 63029
rect 4780 62936 4820 62945
rect 4780 61844 4820 62896
rect 4972 62852 5012 62980
rect 4972 62803 5012 62812
rect 4876 62768 4916 62777
rect 4876 62180 4916 62728
rect 5260 62180 5300 63316
rect 5356 62348 5396 63652
rect 5452 63188 5492 75748
rect 5548 73940 5588 76000
rect 5644 74360 5684 83140
rect 5740 75200 5780 83392
rect 5836 82760 5876 82769
rect 5836 82088 5876 82720
rect 5932 82256 5972 87844
rect 6028 87884 6068 90784
rect 6028 87835 6068 87844
rect 6124 86708 6164 93580
rect 6796 92420 6836 92429
rect 6316 89816 6356 89825
rect 6220 89480 6260 89489
rect 6220 89228 6260 89440
rect 6220 89179 6260 89188
rect 6220 88640 6260 88649
rect 6220 88052 6260 88600
rect 6220 88003 6260 88012
rect 6124 86659 6164 86668
rect 6220 87884 6260 87893
rect 6028 86624 6068 86633
rect 6028 84608 6068 86584
rect 6028 84559 6068 84568
rect 6124 86456 6164 86465
rect 5932 82207 5972 82216
rect 6028 84356 6068 84365
rect 6124 84356 6164 86416
rect 6068 84316 6164 84356
rect 5836 82048 5972 82088
rect 5836 81416 5876 81425
rect 5836 79904 5876 81376
rect 5932 81332 5972 82048
rect 5932 81283 5972 81292
rect 6028 81248 6068 84316
rect 6220 82844 6260 87844
rect 6220 82795 6260 82804
rect 6124 82592 6164 82601
rect 6124 81500 6164 82552
rect 6124 81451 6164 81460
rect 6220 82256 6260 82265
rect 6028 81199 6068 81208
rect 6124 81332 6164 81341
rect 5836 79855 5876 79864
rect 5932 81164 5972 81173
rect 5836 78980 5876 78989
rect 5836 78845 5876 78940
rect 5740 75151 5780 75160
rect 5836 76964 5876 76973
rect 5740 75032 5780 75041
rect 5740 74528 5780 74992
rect 5740 74479 5780 74488
rect 5836 74528 5876 76924
rect 5932 76208 5972 81124
rect 6028 80744 6068 80753
rect 6028 80660 6068 80704
rect 6028 80609 6068 80620
rect 6028 80408 6068 80417
rect 6028 80273 6068 80368
rect 6028 80156 6068 80165
rect 6028 79820 6068 80116
rect 6028 79652 6068 79780
rect 6028 79603 6068 79612
rect 6028 79232 6068 79241
rect 6028 76292 6068 79192
rect 6028 76243 6068 76252
rect 5932 76159 5972 76168
rect 5836 74479 5876 74488
rect 5932 76040 5972 76049
rect 5932 74444 5972 76000
rect 6124 75872 6164 81292
rect 6220 76292 6260 82216
rect 6316 77216 6356 89776
rect 6412 89396 6452 89405
rect 6412 87380 6452 89356
rect 6412 87331 6452 87340
rect 6604 87548 6644 87557
rect 6412 87128 6452 87137
rect 6412 86624 6452 87088
rect 6412 86575 6452 86584
rect 6412 86372 6452 86381
rect 6412 82256 6452 86332
rect 6508 85784 6548 85793
rect 6508 82508 6548 85744
rect 6508 82459 6548 82468
rect 6412 82207 6452 82216
rect 6508 82088 6548 82097
rect 6412 82048 6508 82088
rect 6412 81416 6452 82048
rect 6508 82039 6548 82048
rect 6412 81367 6452 81376
rect 6508 81668 6548 81677
rect 6508 81248 6548 81628
rect 6412 81208 6548 81248
rect 6412 79736 6452 81208
rect 6508 80996 6548 81005
rect 6508 80576 6548 80956
rect 6508 80527 6548 80536
rect 6508 80324 6548 80335
rect 6508 80240 6548 80284
rect 6508 80191 6548 80200
rect 6412 79696 6548 79736
rect 6412 79400 6452 79409
rect 6412 77972 6452 79360
rect 6412 77923 6452 77932
rect 6316 77167 6356 77176
rect 6220 76243 6260 76252
rect 6316 76964 6356 76973
rect 6316 76712 6356 76924
rect 6124 75823 6164 75832
rect 6220 76124 6260 76133
rect 6220 75620 6260 76084
rect 6220 75571 6260 75580
rect 5932 74395 5972 74404
rect 6124 75284 6164 75293
rect 5836 74360 5876 74369
rect 5644 74320 5780 74360
rect 5548 73891 5588 73900
rect 5740 73100 5780 74320
rect 5836 73940 5876 74320
rect 5836 73891 5876 73900
rect 5932 74108 5972 74117
rect 5932 73184 5972 74068
rect 6124 73772 6164 75244
rect 6220 74528 6260 74537
rect 6220 74393 6260 74488
rect 6316 74108 6356 76672
rect 6412 76544 6452 76553
rect 6412 75368 6452 76504
rect 6508 75956 6548 79696
rect 6604 78476 6644 87508
rect 6700 86372 6740 86381
rect 6700 85700 6740 86332
rect 6796 86288 6836 92380
rect 6892 91328 6932 94144
rect 7276 94184 7316 94193
rect 7180 94100 7220 94109
rect 7180 93596 7220 94060
rect 7180 93547 7220 93556
rect 6892 91279 6932 91288
rect 7276 91244 7316 94144
rect 7468 93932 7508 93941
rect 7468 93764 7508 93892
rect 7468 93715 7508 93724
rect 7276 91195 7316 91204
rect 7084 88640 7124 88649
rect 7084 87464 7124 88600
rect 7564 88640 7604 94732
rect 7756 94352 7796 96688
rect 7852 95024 7892 95033
rect 7948 95024 7988 96688
rect 7892 94984 7988 95024
rect 7852 94975 7892 94984
rect 8140 94772 8180 96688
rect 8332 95024 8372 96688
rect 8332 94975 8372 94984
rect 8140 94723 8180 94732
rect 7756 94303 7796 94312
rect 8428 94688 8468 94697
rect 8044 94184 8084 94193
rect 8044 94049 8084 94144
rect 8236 94184 8276 94193
rect 8140 94016 8180 94025
rect 7564 88591 7604 88600
rect 7660 93932 7700 93941
rect 7084 87415 7124 87424
rect 7372 87884 7412 87893
rect 7084 87296 7124 87305
rect 7084 86456 7124 87256
rect 7276 86708 7316 86717
rect 7084 86407 7124 86416
rect 7180 86624 7220 86633
rect 6796 86239 6836 86248
rect 7084 86288 7124 86297
rect 6740 85660 6836 85700
rect 6700 85651 6740 85660
rect 6700 84860 6740 84869
rect 6700 84440 6740 84820
rect 6700 84391 6740 84400
rect 6700 84272 6740 84281
rect 6700 82172 6740 84232
rect 6796 83516 6836 85660
rect 6892 84860 6932 84869
rect 6892 83768 6932 84820
rect 6988 84608 7028 84617
rect 6988 84356 7028 84568
rect 6988 84307 7028 84316
rect 7084 84272 7124 86248
rect 7180 86036 7220 86584
rect 7180 85868 7220 85996
rect 7180 85819 7220 85828
rect 7084 84223 7124 84232
rect 7180 85112 7220 85121
rect 6892 83719 6932 83728
rect 6796 82592 6836 83476
rect 6988 83600 7028 83609
rect 6988 83516 7028 83560
rect 7180 83540 7220 85072
rect 7276 83684 7316 86668
rect 7372 86540 7412 87844
rect 7372 86491 7412 86500
rect 7660 86372 7700 93892
rect 8044 91832 8084 91841
rect 8044 91697 8084 91792
rect 7948 91160 7988 91169
rect 7948 91025 7988 91120
rect 8044 88640 8084 88649
rect 7948 87380 7988 87389
rect 7852 87296 7892 87305
rect 7852 86624 7892 87256
rect 7852 86575 7892 86584
rect 7948 86792 7988 87340
rect 7948 86540 7988 86752
rect 7948 86405 7988 86500
rect 7372 86332 7700 86372
rect 7372 84104 7412 86332
rect 8044 86204 8084 88600
rect 8140 86372 8180 93976
rect 8236 93932 8276 94144
rect 8236 93883 8276 93892
rect 8332 91160 8372 91169
rect 8332 91025 8372 91120
rect 8140 86323 8180 86332
rect 8236 86540 8276 86549
rect 8044 86164 8180 86204
rect 7468 85112 7508 85121
rect 7468 84608 7508 85072
rect 7756 85112 7796 85121
rect 7468 84559 7508 84568
rect 7564 85028 7604 85037
rect 7372 84055 7412 84064
rect 7468 84356 7508 84365
rect 7468 83852 7508 84316
rect 7468 83803 7508 83812
rect 7564 83768 7604 84988
rect 7756 84977 7796 85072
rect 7852 85028 7892 85037
rect 7660 84944 7700 84953
rect 7660 84272 7700 84904
rect 7852 84524 7892 84988
rect 7852 84475 7892 84484
rect 8044 85028 8084 85037
rect 7852 84356 7892 84365
rect 7852 84272 7892 84316
rect 8044 84272 8084 84988
rect 8140 84860 8180 86164
rect 8140 84811 8180 84820
rect 7852 84232 8084 84272
rect 7660 84223 7700 84232
rect 7948 84104 7988 84113
rect 7564 83719 7604 83728
rect 7756 83852 7796 83861
rect 7276 83644 7508 83684
rect 7180 83500 7316 83540
rect 6988 83465 7028 83476
rect 7276 83432 7316 83500
rect 7468 83516 7508 83644
rect 7372 83432 7412 83441
rect 7276 83392 7372 83432
rect 6796 82543 6836 82552
rect 6988 83264 7028 83273
rect 6892 82424 6932 82433
rect 6700 82132 6836 82172
rect 6700 82004 6740 82013
rect 6700 81332 6740 81964
rect 6700 80744 6740 81292
rect 6700 80695 6740 80704
rect 6604 78427 6644 78436
rect 6700 80576 6740 80585
rect 6700 78308 6740 80536
rect 6796 78728 6836 82132
rect 6892 81668 6932 82384
rect 6892 81619 6932 81628
rect 6988 81920 7028 83224
rect 7372 82844 7412 83392
rect 7372 82795 7412 82804
rect 7468 82340 7508 83476
rect 7660 83432 7700 83441
rect 7660 83348 7700 83392
rect 7372 82300 7508 82340
rect 7564 83012 7604 83021
rect 7276 82004 7316 82013
rect 6892 81500 6932 81509
rect 6892 79400 6932 81460
rect 6988 79736 7028 81880
rect 7180 81920 7220 81929
rect 7084 81836 7124 81845
rect 7084 80576 7124 81796
rect 7180 81500 7220 81880
rect 7180 81451 7220 81460
rect 7084 80527 7124 80536
rect 7180 81332 7220 81341
rect 6988 79484 7028 79696
rect 6988 79444 7124 79484
rect 6892 79360 7028 79400
rect 6796 78679 6836 78688
rect 6700 78259 6740 78268
rect 6796 78476 6836 78485
rect 6700 77552 6740 77561
rect 6604 76796 6644 76805
rect 6604 76544 6644 76756
rect 6604 76495 6644 76504
rect 6508 75916 6644 75956
rect 6412 75319 6452 75328
rect 6508 75788 6548 75797
rect 6316 74059 6356 74068
rect 6220 73772 6260 73781
rect 6124 73732 6220 73772
rect 5932 73135 5972 73144
rect 5740 73051 5780 73060
rect 5548 72932 5588 72941
rect 5548 71420 5588 72892
rect 6220 72932 6260 73732
rect 6412 73520 6452 73529
rect 6412 73460 6452 73480
rect 6124 72764 6164 72773
rect 5548 70916 5588 71380
rect 5548 70867 5588 70876
rect 5644 72344 5684 72353
rect 5548 70580 5588 70589
rect 5548 69320 5588 70540
rect 5548 69271 5588 69280
rect 5548 69152 5588 69161
rect 5548 68228 5588 69112
rect 5548 68179 5588 68188
rect 5452 63139 5492 63148
rect 5548 67808 5588 67817
rect 5356 62299 5396 62308
rect 5452 63020 5492 63029
rect 5260 62140 5396 62180
rect 4876 62131 4916 62140
rect 4928 62012 5296 62021
rect 4968 61972 5010 62012
rect 5050 61972 5092 62012
rect 5132 61972 5174 62012
rect 5214 61972 5256 62012
rect 4928 61963 5296 61972
rect 4780 61795 4820 61804
rect 4780 61676 4820 61685
rect 4780 56300 4820 61636
rect 4928 60500 5296 60509
rect 4968 60460 5010 60500
rect 5050 60460 5092 60500
rect 5132 60460 5174 60500
rect 5214 60460 5256 60500
rect 4928 60451 5296 60460
rect 5356 60416 5396 62140
rect 5452 61676 5492 62980
rect 5548 62348 5588 67768
rect 5644 63692 5684 72304
rect 5932 72260 5972 72271
rect 5740 72176 5780 72185
rect 5740 71252 5780 72136
rect 5740 71203 5780 71212
rect 5836 72176 5876 72185
rect 5740 70496 5780 70505
rect 5740 69572 5780 70456
rect 5740 69523 5780 69532
rect 5740 69152 5780 69161
rect 5740 67724 5780 69112
rect 5740 63944 5780 67684
rect 5836 67136 5876 72136
rect 5932 72176 5972 72220
rect 6124 72260 6164 72724
rect 6124 72211 6164 72220
rect 5932 72127 5972 72136
rect 5836 67087 5876 67096
rect 5932 71336 5972 71345
rect 5932 68396 5972 71296
rect 6220 71336 6260 72892
rect 6220 71287 6260 71296
rect 6316 73420 6452 73460
rect 6028 71084 6068 71093
rect 6028 70748 6068 71044
rect 6028 70699 6068 70708
rect 6220 70580 6260 70589
rect 5836 66884 5876 66893
rect 5836 66128 5876 66844
rect 5836 66079 5876 66088
rect 5836 65960 5876 65969
rect 5836 64700 5876 65920
rect 5932 65624 5972 68356
rect 5932 65575 5972 65584
rect 6028 70496 6068 70505
rect 5836 64651 5876 64660
rect 5932 65204 5972 65213
rect 5740 63895 5780 63904
rect 5836 64280 5876 64289
rect 5644 63643 5684 63652
rect 5740 63776 5780 63785
rect 5740 63104 5780 63736
rect 5644 63064 5780 63104
rect 5644 62516 5684 63064
rect 5740 62936 5780 62945
rect 5740 62600 5780 62896
rect 5740 62551 5780 62560
rect 5644 62467 5684 62476
rect 5548 62308 5684 62348
rect 5452 61627 5492 61636
rect 5548 62180 5588 62189
rect 5548 61592 5588 62140
rect 5644 61760 5684 62308
rect 5644 61711 5684 61720
rect 5740 61844 5780 61853
rect 5548 61543 5588 61552
rect 5356 60367 5396 60376
rect 5452 61508 5492 61517
rect 4876 60332 4916 60341
rect 4876 59156 4916 60292
rect 4876 59107 4916 59116
rect 5356 60248 5396 60257
rect 4928 58988 5296 58997
rect 4968 58948 5010 58988
rect 5050 58948 5092 58988
rect 5132 58948 5174 58988
rect 5214 58948 5256 58988
rect 4928 58939 5296 58948
rect 4876 58820 4916 58829
rect 4876 58652 4916 58780
rect 4876 58603 4916 58612
rect 4876 57812 4916 57821
rect 4876 57677 4916 57772
rect 4928 57476 5296 57485
rect 4968 57436 5010 57476
rect 5050 57436 5092 57476
rect 5132 57436 5174 57476
rect 5214 57436 5256 57476
rect 4928 57427 5296 57436
rect 5356 57476 5396 60208
rect 5356 57427 5396 57436
rect 5452 57224 5492 61468
rect 5548 60836 5588 60845
rect 5548 60332 5588 60796
rect 5548 60283 5588 60292
rect 5644 60164 5684 60173
rect 5740 60164 5780 61804
rect 5684 60124 5780 60164
rect 5644 60115 5684 60124
rect 5644 59912 5684 59921
rect 5644 58820 5684 59872
rect 5740 59828 5780 60124
rect 5740 59408 5780 59788
rect 5740 59359 5780 59368
rect 5644 58771 5684 58780
rect 5836 58820 5876 64240
rect 5932 62432 5972 65164
rect 5932 62383 5972 62392
rect 5932 60164 5972 60173
rect 5932 60029 5972 60124
rect 5836 58771 5876 58780
rect 5932 59408 5972 59417
rect 5932 58988 5972 59368
rect 5644 58652 5684 58661
rect 5932 58652 5972 58948
rect 5548 58568 5588 58577
rect 5548 58064 5588 58528
rect 5548 58015 5588 58024
rect 5644 57812 5684 58612
rect 5644 57763 5684 57772
rect 5740 58612 5972 58652
rect 6028 58652 6068 70456
rect 6124 69824 6164 69833
rect 6124 68480 6164 69784
rect 6220 68648 6260 70540
rect 6220 68599 6260 68608
rect 6124 68431 6164 68440
rect 6220 66884 6260 66893
rect 6220 66212 6260 66844
rect 6220 66163 6260 66172
rect 6124 65876 6164 65885
rect 6124 64532 6164 65836
rect 6124 64483 6164 64492
rect 6220 65624 6260 65633
rect 6124 64196 6164 64205
rect 6124 63692 6164 64156
rect 6220 64028 6260 65584
rect 6316 65372 6356 73420
rect 6508 73016 6548 75748
rect 6604 73604 6644 75916
rect 6604 73555 6644 73564
rect 6700 74528 6740 77512
rect 6412 72976 6548 73016
rect 6412 66548 6452 72976
rect 6604 72932 6644 72941
rect 6412 66499 6452 66508
rect 6508 72848 6548 72857
rect 6316 65323 6356 65332
rect 6412 64784 6452 64793
rect 6220 63860 6260 63988
rect 6220 63811 6260 63820
rect 6316 64700 6356 64709
rect 6124 61676 6164 63652
rect 6124 61627 6164 61636
rect 6220 63692 6260 63701
rect 6124 60164 6164 60173
rect 6124 59828 6164 60124
rect 6124 59779 6164 59788
rect 4780 56251 4820 56260
rect 5260 57184 5492 57224
rect 5260 56132 5300 57184
rect 5548 57140 5588 57149
rect 5452 57100 5548 57140
rect 5260 56083 5300 56092
rect 5356 56300 5396 56309
rect 4928 55964 5296 55973
rect 4968 55924 5010 55964
rect 5050 55924 5092 55964
rect 5132 55924 5174 55964
rect 5214 55924 5256 55964
rect 4928 55915 5296 55924
rect 5356 55796 5396 56260
rect 5356 55747 5396 55756
rect 5452 56216 5492 57100
rect 5548 57091 5588 57100
rect 5452 55628 5492 56176
rect 5356 55588 5492 55628
rect 5548 56972 5588 56981
rect 4928 54452 5296 54461
rect 4968 54412 5010 54452
rect 5050 54412 5092 54452
rect 5132 54412 5174 54452
rect 5214 54412 5256 54452
rect 4928 54403 5296 54412
rect 5356 53024 5396 55588
rect 5548 55544 5588 56932
rect 4928 52940 5296 52949
rect 4968 52900 5010 52940
rect 5050 52900 5092 52940
rect 5132 52900 5174 52940
rect 5214 52900 5256 52940
rect 4928 52891 5296 52900
rect 4684 52471 4724 52480
rect 4492 51631 4532 51640
rect 5356 51596 5396 52984
rect 5356 51547 5396 51556
rect 5452 55504 5588 55544
rect 5644 56972 5684 56981
rect 5740 56972 5780 58612
rect 6028 58603 6068 58612
rect 6124 59492 6164 59501
rect 6124 59324 6164 59452
rect 6124 57476 6164 59284
rect 5684 56932 5780 56972
rect 5932 57436 6164 57476
rect 5932 57224 5972 57436
rect 6220 57392 6260 63652
rect 6316 62516 6356 64660
rect 6316 62467 6356 62476
rect 6316 62348 6356 62357
rect 6316 62264 6356 62308
rect 6316 61844 6356 62224
rect 6316 59492 6356 61804
rect 6316 59443 6356 59452
rect 6412 59240 6452 64744
rect 6412 57812 6452 59200
rect 6412 57763 6452 57772
rect 4928 51428 5296 51437
rect 4968 51388 5010 51428
rect 5050 51388 5092 51428
rect 5132 51388 5174 51428
rect 5214 51388 5256 51428
rect 4928 51379 5296 51388
rect 4492 51092 4532 51101
rect 4492 50672 4532 51052
rect 4492 50623 4532 50632
rect 4300 50203 4340 50212
rect 4928 49916 5296 49925
rect 4968 49876 5010 49916
rect 5050 49876 5092 49916
rect 5132 49876 5174 49916
rect 5214 49876 5256 49916
rect 4928 49867 5296 49876
rect 4204 48859 4244 48868
rect 4684 49328 4724 49337
rect 4396 48656 4436 48665
rect 4204 48572 4244 48581
rect 4204 48437 4244 48532
rect 4108 48019 4148 48028
rect 4204 47984 4244 47993
rect 3688 47648 4056 47657
rect 3728 47608 3770 47648
rect 3810 47608 3852 47648
rect 3892 47608 3934 47648
rect 3974 47608 4016 47648
rect 3688 47599 4056 47608
rect 4204 47540 4244 47944
rect 4204 47500 4340 47540
rect 3532 47263 3572 47272
rect 3436 47228 3476 47237
rect 3340 46724 3380 46733
rect 2956 42139 2996 42148
rect 3052 43180 3188 43220
rect 3244 46640 3284 46649
rect 3244 44120 3284 46600
rect 3340 46589 3380 46684
rect 3436 46472 3476 47188
rect 3916 47228 3956 47237
rect 3916 47093 3956 47188
rect 2860 41971 2900 41980
rect 3052 41348 3092 43180
rect 3052 41299 3092 41308
rect 3148 42692 3188 42701
rect 3148 41936 3188 42652
rect 3052 41180 3092 41189
rect 2956 40256 2996 40265
rect 2860 39836 2900 39845
rect 2956 39836 2996 40216
rect 2900 39796 2996 39836
rect 2860 39787 2900 39796
rect 2956 39668 2996 39677
rect 2764 38452 2900 38492
rect 2764 38324 2804 38333
rect 2764 37400 2804 38284
rect 2860 38072 2900 38452
rect 2860 38023 2900 38032
rect 2764 37351 2804 37360
rect 2860 37904 2900 37913
rect 2860 37484 2900 37864
rect 2668 37267 2708 37276
rect 2380 36772 2516 36812
rect 2284 36763 2324 36772
rect 2380 36644 2420 36653
rect 2092 36100 2228 36140
rect 2284 36604 2380 36644
rect 2092 35132 2132 36100
rect 2092 35083 2132 35092
rect 2188 35972 2228 35981
rect 1996 34159 2036 34168
rect 2092 34292 2132 34301
rect 2092 34157 2132 34252
rect 1900 32899 1940 32908
rect 1996 33704 2036 33713
rect 1900 32780 1940 32789
rect 1900 29840 1940 32740
rect 1900 29791 1940 29800
rect 1996 29168 2036 33664
rect 2092 33200 2132 33209
rect 2092 33116 2132 33160
rect 2092 33036 2132 33076
rect 2092 32948 2132 32957
rect 2092 29336 2132 32908
rect 2188 32276 2228 35932
rect 2188 32227 2228 32236
rect 2284 35888 2324 36604
rect 2380 36595 2420 36604
rect 2284 34460 2324 35848
rect 2380 35720 2420 35729
rect 2380 35300 2420 35680
rect 2380 35251 2420 35260
rect 2092 29287 2132 29296
rect 2188 31016 2228 31025
rect 1996 29119 2036 29128
rect 2092 29168 2132 29177
rect 1804 27775 1844 27784
rect 1996 27992 2036 28001
rect 1804 26900 1844 26911
rect 1804 26816 1844 26860
rect 1804 26767 1844 26776
rect 1900 26060 1940 26069
rect 1804 25388 1844 25397
rect 1804 20936 1844 25348
rect 1900 22532 1940 26020
rect 1996 23960 2036 27952
rect 2092 25472 2132 29128
rect 2188 26732 2228 30976
rect 2188 26683 2228 26692
rect 2092 25423 2132 25432
rect 2188 26396 2228 26405
rect 1996 23911 2036 23920
rect 2092 25136 2132 25145
rect 1900 22492 2036 22532
rect 1804 20012 1844 20896
rect 1900 22364 1940 22373
rect 1900 21440 1940 22324
rect 1900 20852 1940 21400
rect 1900 20803 1940 20812
rect 1804 19963 1844 19972
rect 1996 20012 2036 22492
rect 1900 19844 1940 19853
rect 1804 18752 1844 18761
rect 1804 18164 1844 18712
rect 1900 18416 1940 19804
rect 1996 19340 2036 19972
rect 1996 19291 2036 19300
rect 1900 18376 2036 18416
rect 1804 18115 1844 18124
rect 1708 16435 1748 16444
rect 1804 17912 1844 17921
rect 1804 16316 1844 17872
rect 1612 13411 1652 13420
rect 1708 16276 1844 16316
rect 1708 13292 1748 16276
rect 1996 14804 2036 18376
rect 1996 14755 2036 14764
rect 1996 14636 2036 14645
rect 1900 14300 1940 14309
rect 1900 14132 1940 14260
rect 1900 14083 1940 14092
rect 1612 13252 1748 13292
rect 1804 13544 1844 13553
rect 1612 11948 1652 13252
rect 1612 11899 1652 11908
rect 1708 13040 1748 13049
rect 1516 10387 1556 10396
rect 1612 10856 1652 10865
rect 1420 10060 1556 10100
rect 1228 9848 1268 9857
rect 1132 8840 1172 8849
rect 940 6943 980 6952
rect 1036 7496 1076 7505
rect 844 5179 884 5188
rect 556 4255 596 4264
rect 940 5144 980 5153
rect 940 3884 980 5104
rect 1036 4724 1076 7456
rect 1132 5144 1172 8800
rect 1228 6572 1268 9808
rect 1420 8756 1460 8765
rect 1420 7916 1460 8716
rect 1516 8000 1556 10060
rect 1516 7951 1556 7960
rect 1420 7867 1460 7876
rect 1228 6523 1268 6532
rect 1420 7160 1460 7169
rect 1132 5095 1172 5104
rect 1324 6152 1364 6161
rect 1036 4675 1076 4684
rect 1324 4304 1364 6112
rect 1420 5900 1460 7120
rect 1612 6656 1652 10816
rect 1708 10184 1748 13000
rect 1804 10772 1844 13504
rect 1900 13292 1940 13301
rect 1900 12980 1940 13252
rect 1900 12931 1940 12940
rect 1996 12872 2036 14596
rect 1900 12832 2036 12872
rect 1900 11276 1940 12832
rect 1900 11227 1940 11236
rect 1996 11528 2036 11537
rect 1804 10732 1940 10772
rect 1708 10135 1748 10144
rect 1804 10604 1844 10613
rect 1708 10016 1748 10025
rect 1708 9680 1748 9976
rect 1708 9631 1748 9640
rect 1612 6607 1652 6616
rect 1708 9428 1748 9437
rect 1612 6488 1652 6497
rect 1612 6152 1652 6448
rect 1612 6103 1652 6112
rect 1420 5851 1460 5860
rect 1708 5480 1748 9388
rect 1804 8756 1844 10564
rect 1900 8840 1940 10732
rect 1900 8791 1940 8800
rect 1804 8707 1844 8716
rect 1804 8588 1844 8597
rect 1804 7160 1844 8548
rect 1804 7111 1844 7120
rect 1996 7160 2036 11488
rect 2092 10520 2132 25096
rect 2188 17996 2228 26356
rect 2188 17947 2228 17956
rect 2188 15056 2228 15065
rect 2188 13964 2228 15016
rect 2284 14132 2324 34420
rect 2380 35048 2420 35057
rect 2380 29756 2420 35008
rect 2476 34376 2516 36772
rect 2476 34327 2516 34336
rect 2572 36728 2612 36737
rect 2572 33872 2612 36688
rect 2764 35972 2804 35981
rect 2764 34880 2804 35932
rect 2764 34831 2804 34840
rect 2668 34712 2708 34723
rect 2668 34628 2708 34672
rect 2668 34579 2708 34588
rect 2764 34544 2804 34553
rect 2572 33823 2612 33832
rect 2668 34460 2708 34469
rect 2572 33704 2612 33713
rect 2476 33620 2516 33629
rect 2476 32948 2516 33580
rect 2476 32108 2516 32908
rect 2476 32059 2516 32068
rect 2380 29707 2420 29716
rect 2476 30596 2516 30605
rect 2476 29336 2516 30556
rect 2572 29840 2612 33664
rect 2668 33536 2708 34420
rect 2764 33620 2804 34504
rect 2860 33788 2900 37444
rect 2956 35216 2996 39628
rect 3052 38240 3092 41140
rect 3148 40760 3188 41896
rect 3148 40711 3188 40720
rect 3148 40508 3188 40517
rect 3148 39752 3188 40468
rect 3148 39500 3188 39712
rect 3148 39451 3188 39460
rect 3244 38324 3284 44080
rect 3340 44204 3380 44213
rect 3340 43868 3380 44164
rect 3436 44036 3476 46432
rect 4300 46388 4340 47500
rect 4204 46304 4244 46313
rect 3688 46136 4056 46145
rect 3728 46096 3770 46136
rect 3810 46096 3852 46136
rect 3892 46096 3934 46136
rect 3974 46096 4016 46136
rect 3688 46087 4056 46096
rect 3916 45968 3956 45979
rect 3916 45884 3956 45928
rect 3916 45835 3956 45844
rect 4012 45800 4052 45809
rect 3916 45716 3956 45725
rect 3916 45128 3956 45676
rect 4012 45665 4052 45760
rect 4108 45716 4148 45725
rect 4108 45212 4148 45676
rect 4108 45163 4148 45172
rect 3916 45079 3956 45088
rect 4108 45044 4148 45053
rect 3688 44624 4056 44633
rect 3728 44584 3770 44624
rect 3810 44584 3852 44624
rect 3892 44584 3934 44624
rect 3974 44584 4016 44624
rect 3688 44575 4056 44584
rect 4012 44456 4052 44465
rect 3916 44372 3956 44381
rect 3436 43987 3476 43996
rect 3532 44204 3572 44213
rect 3340 43828 3476 43868
rect 3244 38275 3284 38284
rect 3340 40508 3380 40517
rect 3052 38191 3092 38200
rect 3340 38156 3380 40468
rect 3148 38116 3380 38156
rect 3052 38072 3092 38081
rect 3052 36812 3092 38032
rect 3052 36763 3092 36772
rect 2956 35167 2996 35176
rect 3052 36140 3092 36149
rect 2956 35048 2996 35057
rect 2956 34544 2996 35008
rect 2956 34495 2996 34504
rect 2860 33739 2900 33748
rect 2956 34376 2996 34385
rect 2764 33571 2804 33580
rect 2956 33536 2996 34336
rect 3052 33704 3092 36100
rect 3052 33655 3092 33664
rect 2668 30848 2708 33496
rect 2860 33496 2996 33536
rect 3052 33536 3092 33545
rect 2860 33140 2900 33496
rect 2764 33100 2900 33140
rect 2956 33368 2996 33377
rect 2764 31604 2804 33100
rect 2860 32108 2900 32117
rect 2956 32108 2996 33328
rect 2900 32068 2996 32108
rect 2860 32059 2900 32068
rect 3052 32024 3092 33496
rect 3148 33536 3188 38116
rect 3436 38072 3476 43828
rect 3532 42104 3572 44164
rect 3916 43952 3956 44332
rect 4012 44321 4052 44416
rect 3916 43903 3956 43912
rect 3628 43532 3668 43541
rect 3628 43397 3668 43492
rect 4108 43532 4148 45004
rect 4204 44288 4244 46264
rect 4204 44239 4244 44248
rect 4012 43448 4052 43457
rect 4012 43280 4052 43408
rect 4012 43231 4052 43240
rect 3688 43112 4056 43121
rect 3728 43072 3770 43112
rect 3810 43072 3852 43112
rect 3892 43072 3934 43112
rect 3974 43072 4016 43112
rect 3688 43063 4056 43072
rect 4108 42776 4148 43492
rect 3532 42055 3572 42064
rect 3628 42188 3668 42197
rect 3628 41768 3668 42148
rect 4108 41852 4148 42736
rect 4108 41803 4148 41812
rect 4204 43616 4244 43625
rect 3532 41728 3668 41768
rect 3532 40928 3572 41728
rect 3688 41600 4056 41609
rect 3728 41560 3770 41600
rect 3810 41560 3852 41600
rect 3892 41560 3934 41600
rect 3974 41560 4016 41600
rect 3688 41551 4056 41560
rect 4108 41432 4148 41441
rect 4108 41180 4148 41392
rect 4108 41131 4148 41140
rect 4012 41012 4052 41021
rect 3532 40888 3668 40928
rect 3532 40760 3572 40769
rect 3532 38492 3572 40720
rect 3628 40256 3668 40888
rect 4012 40508 4052 40972
rect 4108 40928 4148 41023
rect 4108 40879 4148 40888
rect 4012 40459 4052 40468
rect 3628 40207 3668 40216
rect 3688 40088 4056 40097
rect 3728 40048 3770 40088
rect 3810 40048 3852 40088
rect 3892 40048 3934 40088
rect 3974 40048 4016 40088
rect 3688 40039 4056 40048
rect 4204 39500 4244 43576
rect 4204 39451 4244 39460
rect 4300 39332 4340 46348
rect 4396 43220 4436 48616
rect 4492 48236 4532 48245
rect 4492 46472 4532 48196
rect 4492 46423 4532 46432
rect 4588 48068 4628 48077
rect 4492 45800 4532 45809
rect 4492 45632 4532 45760
rect 4492 45583 4532 45592
rect 4492 45464 4532 45475
rect 4492 45380 4532 45424
rect 4492 45331 4532 45340
rect 4492 44960 4532 44969
rect 4492 44372 4532 44920
rect 4492 44120 4532 44332
rect 4492 43784 4532 44080
rect 4492 43735 4532 43744
rect 4588 43700 4628 48028
rect 4684 47228 4724 49288
rect 4684 47179 4724 47188
rect 4780 48824 4820 48833
rect 4780 47060 4820 48784
rect 4928 48404 5296 48413
rect 4968 48364 5010 48404
rect 5050 48364 5092 48404
rect 5132 48364 5174 48404
rect 5214 48364 5256 48404
rect 4928 48355 5296 48364
rect 4876 47984 4916 47993
rect 4876 47849 4916 47944
rect 5356 47984 5396 47993
rect 4780 47011 4820 47020
rect 4928 46892 5296 46901
rect 4968 46852 5010 46892
rect 5050 46852 5092 46892
rect 5132 46852 5174 46892
rect 5214 46852 5256 46892
rect 4928 46843 5296 46852
rect 4684 46724 4724 46733
rect 4684 46589 4724 46684
rect 5164 46724 5204 46733
rect 4972 46388 5012 46397
rect 4780 45968 4820 45977
rect 4780 45884 4820 45928
rect 4780 45833 4820 45844
rect 4684 45800 4724 45811
rect 4684 45716 4724 45760
rect 4684 45667 4724 45676
rect 4972 45548 5012 46348
rect 5068 46052 5108 46061
rect 5068 45716 5108 46012
rect 5164 45884 5204 46684
rect 5356 46556 5396 47944
rect 5452 46724 5492 55504
rect 5548 54788 5588 54797
rect 5548 53276 5588 54748
rect 5548 53227 5588 53236
rect 5548 52604 5588 52613
rect 5548 51932 5588 52564
rect 5548 51883 5588 51892
rect 5644 48908 5684 56932
rect 5932 56552 5972 57184
rect 5932 56503 5972 56512
rect 6028 57352 6260 57392
rect 6412 57644 6452 57653
rect 5836 56300 5876 56309
rect 5740 54116 5780 54125
rect 5740 53696 5780 54076
rect 5740 53647 5780 53656
rect 5740 53276 5780 53285
rect 5740 52772 5780 53236
rect 5740 52723 5780 52732
rect 5836 53192 5876 56260
rect 6028 54788 6068 57352
rect 6412 57140 6452 57604
rect 6412 57091 6452 57100
rect 6028 54739 6068 54748
rect 6124 56972 6164 56981
rect 6028 54284 6068 54293
rect 5836 51092 5876 53152
rect 5932 53948 5972 53957
rect 5932 53612 5972 53908
rect 5932 52520 5972 53572
rect 5932 52471 5972 52480
rect 6028 53108 6068 54244
rect 6124 53948 6164 56932
rect 6412 56384 6452 56393
rect 6412 56249 6452 56344
rect 6316 55796 6356 55805
rect 6220 55376 6260 55385
rect 6220 55241 6260 55336
rect 6220 54284 6260 54379
rect 6220 54235 6260 54244
rect 6316 54116 6356 55756
rect 6124 53899 6164 53908
rect 6220 54076 6356 54116
rect 6412 55712 6452 55721
rect 6028 52604 6068 53068
rect 6028 52016 6068 52564
rect 6028 51967 6068 51976
rect 6124 53780 6164 53789
rect 5836 51043 5876 51052
rect 5452 46675 5492 46684
rect 5548 48868 5684 48908
rect 5740 50084 5780 50093
rect 5396 46516 5492 46556
rect 5356 46507 5396 46516
rect 5356 46388 5396 46397
rect 5164 45835 5204 45844
rect 5260 46052 5300 46061
rect 5260 45800 5300 46012
rect 5260 45751 5300 45760
rect 5068 45667 5108 45676
rect 4972 45499 5012 45508
rect 4780 45464 4820 45473
rect 4684 44960 4724 44969
rect 4684 44204 4724 44920
rect 4684 44155 4724 44164
rect 4588 43651 4628 43660
rect 4684 44036 4724 44045
rect 4396 43180 4532 43220
rect 4396 43112 4436 43121
rect 4396 39752 4436 43072
rect 4492 41264 4532 43180
rect 4684 42944 4724 43996
rect 4780 43280 4820 45424
rect 4928 45380 5296 45389
rect 4968 45340 5010 45380
rect 5050 45340 5092 45380
rect 5132 45340 5174 45380
rect 5214 45340 5256 45380
rect 4928 45331 5296 45340
rect 5356 45128 5396 46348
rect 5452 46136 5492 46516
rect 5452 46087 5492 46096
rect 5452 45968 5492 45979
rect 5452 45884 5492 45928
rect 5452 45835 5492 45844
rect 5452 45212 5492 45307
rect 5452 45163 5492 45172
rect 5356 45079 5396 45088
rect 5452 45044 5492 45053
rect 5164 44876 5204 44885
rect 5068 44372 5108 44381
rect 4876 44288 4916 44297
rect 4876 44036 4916 44248
rect 5068 44237 5108 44332
rect 4876 43987 4916 43996
rect 5164 44036 5204 44836
rect 5260 44624 5300 44633
rect 5260 44456 5300 44584
rect 5452 44540 5492 45004
rect 5452 44491 5492 44500
rect 5260 44407 5300 44416
rect 5260 44288 5300 44297
rect 5300 44248 5396 44288
rect 5260 44153 5300 44248
rect 5164 43987 5204 43996
rect 4928 43868 5296 43877
rect 4968 43828 5010 43868
rect 5050 43828 5092 43868
rect 5132 43828 5174 43868
rect 5214 43828 5256 43868
rect 4928 43819 5296 43828
rect 5356 43868 5396 44248
rect 5452 44120 5492 44129
rect 5452 43985 5492 44080
rect 5356 43819 5396 43828
rect 5452 43868 5492 43877
rect 5260 43700 5300 43709
rect 5260 43616 5300 43660
rect 5260 43565 5300 43576
rect 5356 43616 5396 43625
rect 4972 43364 5012 43373
rect 4780 43231 4820 43240
rect 4876 43280 4916 43289
rect 4684 42895 4724 42904
rect 4588 42860 4628 42869
rect 4588 42524 4628 42820
rect 4684 42692 4724 42787
rect 4684 42643 4724 42652
rect 4684 42524 4724 42533
rect 4876 42524 4916 43240
rect 4972 42944 5012 43324
rect 4972 42895 5012 42904
rect 5260 43364 5300 43373
rect 5164 42860 5204 42869
rect 5164 42725 5204 42820
rect 4588 42484 4684 42524
rect 4588 42020 4628 42029
rect 4588 41600 4628 41980
rect 4588 41551 4628 41560
rect 4588 41432 4628 41441
rect 4588 41297 4628 41392
rect 4492 40676 4532 41224
rect 4684 41180 4724 42484
rect 4780 42484 4916 42524
rect 5260 42608 5300 43324
rect 5356 42692 5396 43576
rect 5356 42643 5396 42652
rect 5260 42524 5300 42568
rect 5260 42484 5396 42524
rect 4780 42356 4820 42484
rect 4780 42307 4820 42316
rect 4928 42356 5296 42365
rect 4968 42316 5010 42356
rect 5050 42316 5092 42356
rect 5132 42316 5174 42356
rect 5214 42316 5256 42356
rect 4928 42307 5296 42316
rect 5356 42104 5396 42484
rect 5260 42064 5396 42104
rect 4492 40627 4532 40636
rect 4588 41140 4724 41180
rect 4780 41852 4820 41861
rect 4396 39703 4436 39712
rect 4492 39752 4532 39763
rect 4492 39668 4532 39712
rect 4492 39619 4532 39628
rect 4300 39283 4340 39292
rect 4396 39584 4436 39593
rect 3724 39248 3764 39259
rect 3724 39164 3764 39208
rect 3724 39115 3764 39124
rect 4012 38996 4052 39005
rect 4300 38996 4340 39005
rect 4052 38956 4148 38996
rect 4012 38947 4052 38956
rect 4108 38912 4148 38956
rect 3688 38576 4056 38585
rect 3728 38536 3770 38576
rect 3810 38536 3852 38576
rect 3892 38536 3934 38576
rect 3974 38536 4016 38576
rect 3688 38527 4056 38536
rect 3532 38443 3572 38452
rect 3148 33487 3188 33496
rect 3244 38032 3476 38072
rect 3532 38324 3572 38333
rect 3148 33368 3188 33377
rect 3148 32192 3188 33328
rect 3148 32143 3188 32152
rect 2956 31940 2996 31949
rect 2764 31564 2900 31604
rect 2860 31184 2900 31564
rect 2860 31135 2900 31144
rect 2668 30799 2708 30808
rect 2668 30512 2708 30521
rect 2668 30344 2708 30472
rect 2668 30295 2708 30304
rect 2860 30176 2900 30185
rect 2668 30136 2860 30176
rect 2668 30092 2708 30136
rect 2860 30127 2900 30136
rect 2668 30043 2708 30052
rect 2572 29791 2612 29800
rect 2860 29672 2900 29681
rect 2380 29296 2516 29336
rect 2764 29632 2860 29672
rect 2380 26060 2420 29296
rect 2476 29168 2516 29177
rect 2476 28244 2516 29128
rect 2668 29084 2708 29093
rect 2476 27740 2516 28204
rect 2476 27691 2516 27700
rect 2572 28916 2612 28925
rect 2380 26011 2420 26020
rect 2476 27572 2516 27581
rect 2476 25388 2516 27532
rect 2572 26984 2612 28876
rect 2668 27824 2708 29044
rect 2764 28580 2804 29632
rect 2860 29604 2900 29632
rect 2860 29084 2900 29179
rect 2860 29035 2900 29044
rect 2860 28832 2900 28927
rect 2860 28783 2900 28792
rect 2860 28580 2900 28589
rect 2764 28540 2860 28580
rect 2860 28512 2900 28540
rect 2668 27775 2708 27784
rect 2764 28412 2804 28421
rect 2572 26935 2612 26944
rect 2668 27656 2708 27665
rect 2668 26060 2708 27616
rect 2764 27572 2804 28372
rect 2764 26900 2804 27532
rect 2956 27404 2996 31900
rect 3052 31520 3092 31984
rect 3052 31471 3092 31480
rect 3148 31772 3188 31781
rect 3052 31352 3092 31361
rect 3052 30764 3092 31312
rect 3052 30680 3092 30724
rect 3052 30600 3092 30640
rect 3148 30260 3188 31732
rect 3052 30220 3188 30260
rect 3052 29336 3092 30220
rect 3052 28412 3092 29296
rect 3148 30092 3188 30101
rect 3148 29168 3188 30052
rect 3148 29119 3188 29128
rect 3052 28363 3092 28372
rect 3148 28496 3188 28505
rect 3148 28361 3188 28456
rect 2764 26851 2804 26860
rect 2860 27364 2956 27404
rect 2764 26060 2804 26069
rect 2668 26020 2764 26060
rect 2764 26011 2804 26020
rect 2764 25892 2804 25901
rect 2476 25348 2708 25388
rect 2476 25220 2516 25229
rect 2380 23288 2420 23297
rect 2380 23036 2420 23248
rect 2380 22901 2420 22996
rect 2380 22196 2420 22205
rect 2380 21608 2420 22156
rect 2380 21559 2420 21568
rect 2380 21356 2420 21365
rect 2380 21221 2420 21316
rect 2380 20852 2420 20861
rect 2380 20717 2420 20812
rect 2380 18500 2420 18509
rect 2380 17156 2420 18460
rect 2380 17107 2420 17116
rect 2380 16400 2420 16411
rect 2380 16316 2420 16360
rect 2380 16267 2420 16276
rect 2284 14083 2324 14092
rect 2380 14048 2420 14057
rect 2188 13924 2324 13964
rect 2092 10471 2132 10480
rect 1996 7111 2036 7120
rect 2092 10352 2132 10361
rect 2092 5816 2132 10312
rect 2284 10352 2324 13924
rect 2380 12536 2420 14008
rect 2476 13880 2516 25180
rect 2572 24548 2612 24557
rect 2572 23876 2612 24508
rect 2572 20012 2612 23836
rect 2668 20768 2708 25348
rect 2764 24548 2804 25852
rect 2860 24884 2900 27364
rect 2956 27355 2996 27364
rect 3052 28076 3092 28085
rect 3052 26144 3092 28036
rect 2860 24835 2900 24844
rect 2956 25472 2996 25481
rect 2860 24548 2900 24557
rect 2764 24508 2860 24548
rect 2860 24480 2900 24508
rect 2860 24380 2900 24389
rect 2860 21776 2900 24340
rect 2956 23372 2996 25432
rect 3052 24800 3092 26104
rect 3052 24751 3092 24760
rect 3148 26312 3188 26321
rect 3148 24716 3188 26272
rect 3148 24667 3188 24676
rect 2956 23323 2996 23332
rect 3052 24464 3092 24473
rect 3052 23792 3092 24424
rect 3052 23204 3092 23752
rect 3244 23540 3284 38032
rect 3436 37568 3476 37577
rect 3340 37232 3380 37241
rect 3340 36140 3380 37192
rect 3436 36560 3476 37528
rect 3532 36896 3572 38284
rect 4108 38156 4148 38872
rect 4108 38107 4148 38116
rect 4204 38912 4244 38921
rect 3820 37736 3860 37745
rect 3820 37484 3860 37696
rect 3820 37435 3860 37444
rect 4108 37232 4148 37241
rect 3688 37064 4056 37073
rect 3728 37024 3770 37064
rect 3810 37024 3852 37064
rect 3892 37024 3934 37064
rect 3974 37024 4016 37064
rect 3688 37015 4056 37024
rect 3532 36856 3764 36896
rect 3628 36728 3668 36737
rect 3436 36511 3476 36520
rect 3532 36644 3572 36653
rect 3340 36091 3380 36100
rect 3436 35972 3476 35981
rect 3340 35804 3380 35813
rect 3340 34376 3380 35764
rect 3340 34327 3380 34336
rect 3340 34208 3380 34217
rect 3340 33536 3380 34168
rect 3340 33487 3380 33496
rect 3340 33368 3380 33377
rect 3340 32108 3380 33328
rect 3436 33116 3476 35932
rect 3532 35384 3572 36604
rect 3628 35888 3668 36688
rect 3628 35839 3668 35848
rect 3724 35888 3764 36856
rect 3724 35839 3764 35848
rect 3820 36560 3860 36569
rect 3820 35804 3860 36520
rect 4012 36140 4052 36235
rect 4012 36091 4052 36100
rect 4108 36056 4148 37192
rect 4108 36007 4148 36016
rect 3820 35755 3860 35764
rect 4108 35888 4148 35897
rect 3688 35552 4056 35561
rect 3728 35512 3770 35552
rect 3810 35512 3852 35552
rect 3892 35512 3934 35552
rect 3974 35512 4016 35552
rect 3688 35503 4056 35512
rect 3532 35335 3572 35344
rect 4012 35132 4052 35141
rect 3436 33067 3476 33076
rect 3532 34460 3572 34469
rect 3532 33704 3572 34420
rect 4012 34208 4052 35092
rect 4012 34159 4052 34168
rect 3688 34040 4056 34049
rect 3728 34000 3770 34040
rect 3810 34000 3852 34040
rect 3892 34000 3934 34040
rect 3974 34000 4016 34040
rect 3688 33991 4056 34000
rect 4108 33872 4148 35848
rect 4204 35384 4244 38872
rect 4300 38861 4340 38956
rect 4300 38408 4340 38503
rect 4300 38359 4340 38368
rect 4300 38240 4340 38249
rect 4300 38105 4340 38200
rect 4204 35335 4244 35344
rect 4396 35300 4436 39544
rect 4492 39500 4532 39509
rect 4492 36224 4532 39460
rect 4492 36175 4532 36184
rect 4588 36056 4628 41140
rect 4684 41012 4724 41021
rect 4684 39164 4724 40972
rect 4780 39920 4820 41812
rect 5164 41180 5204 41191
rect 5164 41096 5204 41140
rect 5164 41047 5204 41056
rect 5260 41096 5300 42064
rect 5356 41936 5396 41947
rect 5356 41852 5396 41896
rect 5356 41803 5396 41812
rect 5356 41348 5396 41357
rect 5356 41264 5396 41308
rect 5356 41213 5396 41224
rect 5260 41047 5300 41056
rect 5356 41012 5396 41021
rect 4928 40844 5296 40853
rect 4968 40804 5010 40844
rect 5050 40804 5092 40844
rect 5132 40804 5174 40844
rect 5214 40804 5256 40844
rect 4928 40795 5296 40804
rect 4972 40676 5012 40685
rect 4876 40340 4916 40349
rect 4876 40088 4916 40300
rect 4876 40039 4916 40048
rect 4780 39880 4916 39920
rect 4684 39115 4724 39124
rect 4780 39752 4820 39761
rect 4684 38996 4724 39005
rect 4684 37484 4724 38956
rect 4780 38912 4820 39712
rect 4876 39500 4916 39880
rect 4972 39584 5012 40636
rect 5068 40676 5108 40685
rect 5068 39668 5108 40636
rect 5164 40508 5204 40517
rect 5164 40373 5204 40468
rect 5260 40424 5300 40519
rect 5260 40375 5300 40384
rect 5164 39836 5204 39845
rect 5164 39701 5204 39796
rect 5356 39752 5396 40972
rect 5356 39703 5396 39712
rect 5068 39619 5108 39628
rect 4972 39535 5012 39544
rect 4876 39451 4916 39460
rect 5164 39500 5204 39595
rect 5164 39451 5204 39460
rect 4928 39332 5296 39341
rect 4968 39292 5010 39332
rect 5050 39292 5092 39332
rect 5132 39292 5174 39332
rect 5214 39292 5256 39332
rect 4928 39283 5296 39292
rect 5356 39332 5396 39341
rect 4780 38863 4820 38872
rect 4876 39164 4916 39173
rect 4876 38660 4916 39124
rect 4684 37435 4724 37444
rect 4780 38620 4916 38660
rect 4780 37484 4820 38620
rect 4928 37820 5296 37829
rect 4968 37780 5010 37820
rect 5050 37780 5092 37820
rect 5132 37780 5174 37820
rect 5214 37780 5256 37820
rect 4928 37771 5296 37780
rect 4588 36007 4628 36016
rect 4684 37316 4724 37325
rect 4684 36560 4724 37276
rect 4396 35251 4436 35260
rect 4492 35972 4532 35981
rect 4492 35468 4532 35932
rect 3532 32948 3572 33664
rect 3340 32059 3380 32068
rect 3436 32908 3572 32948
rect 3628 33832 4148 33872
rect 4204 35216 4244 35225
rect 3340 31940 3380 31949
rect 3340 31772 3380 31900
rect 3340 31723 3380 31732
rect 3340 30764 3380 30773
rect 3340 28328 3380 30724
rect 3340 28279 3380 28288
rect 3340 27740 3380 27749
rect 3340 24632 3380 27700
rect 3340 23708 3380 24592
rect 3340 23659 3380 23668
rect 3244 23500 3380 23540
rect 3340 23288 3380 23500
rect 3244 23248 3380 23288
rect 3436 23288 3476 32908
rect 3628 32780 3668 33832
rect 4204 33788 4244 35176
rect 4396 34460 4436 34469
rect 3916 33748 4244 33788
rect 4300 34124 4340 34133
rect 3724 33704 3764 33713
rect 3724 33452 3764 33664
rect 3724 33403 3764 33412
rect 3820 33620 3860 33629
rect 3820 32948 3860 33580
rect 3916 33032 3956 33748
rect 4204 33620 4244 33629
rect 4204 33140 4244 33580
rect 3916 32983 3956 32992
rect 4108 33100 4244 33140
rect 3820 32899 3860 32908
rect 3628 32731 3668 32740
rect 3688 32528 4056 32537
rect 3728 32488 3770 32528
rect 3810 32488 3852 32528
rect 3892 32488 3934 32528
rect 3974 32488 4016 32528
rect 3688 32479 4056 32488
rect 3532 32444 3572 32453
rect 3532 32360 3572 32404
rect 3532 32309 3572 32320
rect 3532 31184 3572 31193
rect 3532 29168 3572 31144
rect 3688 31016 4056 31025
rect 3728 30976 3770 31016
rect 3810 30976 3852 31016
rect 3892 30976 3934 31016
rect 3974 30976 4016 31016
rect 3688 30967 4056 30976
rect 3916 30596 3956 30605
rect 3916 30344 3956 30556
rect 3916 30295 3956 30304
rect 4012 29672 4052 29767
rect 4012 29623 4052 29632
rect 3688 29504 4056 29513
rect 3728 29464 3770 29504
rect 3810 29464 3852 29504
rect 3892 29464 3934 29504
rect 3974 29464 4016 29504
rect 3688 29455 4056 29464
rect 4012 29336 4052 29345
rect 3532 29128 3668 29168
rect 3532 29000 3572 29009
rect 3532 27740 3572 28960
rect 3628 28160 3668 29128
rect 3724 29084 3764 29093
rect 3724 28328 3764 29044
rect 3916 28916 3956 28925
rect 3916 28496 3956 28876
rect 4012 28832 4052 29296
rect 4012 28783 4052 28792
rect 4012 28664 4052 28673
rect 4012 28529 4052 28624
rect 3916 28447 3956 28456
rect 3724 28279 3764 28288
rect 3628 28111 3668 28120
rect 3688 27992 4056 28001
rect 3728 27952 3770 27992
rect 3810 27952 3852 27992
rect 3892 27952 3934 27992
rect 3974 27952 4016 27992
rect 3688 27943 4056 27952
rect 3532 27691 3572 27700
rect 3916 27740 3956 27749
rect 3532 27572 3572 27581
rect 3532 26900 3572 27532
rect 3916 27572 3956 27700
rect 3916 27523 3956 27532
rect 4012 27488 4052 27499
rect 4012 27404 4052 27448
rect 4012 27355 4052 27364
rect 3532 26851 3572 26860
rect 3628 27068 3668 27077
rect 3628 26648 3668 27028
rect 3820 26900 3860 26909
rect 3820 26765 3860 26860
rect 3532 26608 3668 26648
rect 3532 26144 3572 26608
rect 3688 26480 4056 26489
rect 3728 26440 3770 26480
rect 3810 26440 3852 26480
rect 3892 26440 3934 26480
rect 3974 26440 4016 26480
rect 3688 26431 4056 26440
rect 3916 26312 3956 26321
rect 3628 26144 3668 26153
rect 3532 26104 3628 26144
rect 3628 26095 3668 26104
rect 2956 23164 3092 23204
rect 3148 23204 3188 23213
rect 2956 22196 2996 23164
rect 3052 23060 3092 23069
rect 3052 22448 3092 23020
rect 3148 22532 3188 23164
rect 3244 22952 3284 23248
rect 3436 23239 3476 23248
rect 3532 25976 3572 25985
rect 3244 22903 3284 22912
rect 3340 23120 3380 23129
rect 3148 22492 3284 22532
rect 3052 22408 3188 22448
rect 3052 22196 3092 22205
rect 2956 22156 3052 22196
rect 2860 21727 2900 21736
rect 2956 21608 2996 21617
rect 2668 20719 2708 20728
rect 2764 20852 2804 20861
rect 2572 19340 2612 19972
rect 2572 15980 2612 19300
rect 2668 18668 2708 18677
rect 2668 18416 2708 18628
rect 2668 18367 2708 18376
rect 2572 15931 2612 15940
rect 2668 17996 2708 18005
rect 2476 13831 2516 13840
rect 2572 14552 2612 14561
rect 2572 12980 2612 14512
rect 2668 14048 2708 17956
rect 2764 17828 2804 20812
rect 2860 20600 2900 20609
rect 2860 20465 2900 20560
rect 2860 19424 2900 19433
rect 2860 18500 2900 19384
rect 2956 19256 2996 21568
rect 3052 21440 3092 22156
rect 3052 19424 3092 21400
rect 3052 19375 3092 19384
rect 2956 19216 3092 19256
rect 3052 19172 3092 19216
rect 2860 18451 2900 18460
rect 2956 18584 2996 18593
rect 3052 18584 3092 19132
rect 2996 18544 3092 18584
rect 2860 17828 2900 17837
rect 2764 17788 2860 17828
rect 2764 17156 2804 17788
rect 2860 17760 2900 17788
rect 2956 17828 2996 18544
rect 2956 17779 2996 17788
rect 3052 18416 3092 18425
rect 3052 17576 3092 18376
rect 3052 17527 3092 17536
rect 2860 17156 2900 17184
rect 2764 17116 2860 17156
rect 2860 17107 2900 17116
rect 2860 16988 2900 16997
rect 2764 16948 2860 16988
rect 2764 15728 2804 16948
rect 2860 16920 2900 16948
rect 2764 15679 2804 15688
rect 2956 16316 2996 16325
rect 2956 15560 2996 16276
rect 2668 13999 2708 14008
rect 2764 15520 2996 15560
rect 2764 15476 2804 15520
rect 2380 11696 2420 12496
rect 2380 11647 2420 11656
rect 2476 12940 2612 12980
rect 2668 13880 2708 13889
rect 2284 10303 2324 10312
rect 2380 11444 2420 11453
rect 2284 10184 2324 10193
rect 1708 5431 1748 5440
rect 1804 5776 2132 5816
rect 2188 10100 2228 10109
rect 1804 5312 1844 5776
rect 1708 5272 1844 5312
rect 1996 5648 2036 5657
rect 1420 4976 1460 4985
rect 1420 4640 1460 4936
rect 1420 4591 1460 4600
rect 1324 4255 1364 4264
rect 940 3835 980 3844
rect 1516 4052 1556 4061
rect 364 3583 404 3592
rect 1516 3632 1556 4012
rect 1516 3583 1556 3592
rect 76 3128 116 3137
rect 76 2960 116 3088
rect 76 2911 116 2920
rect 1420 2960 1460 2969
rect 1420 2624 1460 2920
rect 1420 2575 1460 2584
rect 1708 2624 1748 5272
rect 1996 5144 2036 5608
rect 1996 5095 2036 5104
rect 2092 5564 2132 5573
rect 2092 4724 2132 5524
rect 2092 4675 2132 4684
rect 2188 4136 2228 10060
rect 2284 10049 2324 10144
rect 2284 9596 2324 9605
rect 2284 9428 2324 9556
rect 2284 8084 2324 9388
rect 2284 7244 2324 8044
rect 2284 6488 2324 7204
rect 2284 6439 2324 6448
rect 2380 5648 2420 11404
rect 2476 10772 2516 12940
rect 2476 10723 2516 10732
rect 2572 12368 2612 12377
rect 2476 10520 2516 10529
rect 2476 9596 2516 10480
rect 2476 9547 2516 9556
rect 2476 9428 2516 9437
rect 2476 8756 2516 9388
rect 2572 8924 2612 12328
rect 2668 11192 2708 13840
rect 2764 13712 2804 15436
rect 3148 15476 3188 22408
rect 3244 18584 3284 22492
rect 3340 20096 3380 23080
rect 3436 23120 3476 23129
rect 3436 22532 3476 23080
rect 3532 23036 3572 25936
rect 3628 25640 3668 25649
rect 3628 25304 3668 25600
rect 3820 25640 3860 25649
rect 3820 25472 3860 25600
rect 3820 25423 3860 25432
rect 3916 25472 3956 26272
rect 4012 25892 4052 25901
rect 4012 25724 4052 25852
rect 4012 25675 4052 25684
rect 3916 25423 3956 25432
rect 3628 25255 3668 25264
rect 3688 24968 4056 24977
rect 3728 24928 3770 24968
rect 3810 24928 3852 24968
rect 3892 24928 3934 24968
rect 3974 24928 4016 24968
rect 3688 24919 4056 24928
rect 3628 24800 3668 24809
rect 3628 24548 3668 24760
rect 3628 23792 3668 24508
rect 3724 24716 3764 24725
rect 3724 23960 3764 24676
rect 3724 23911 3764 23920
rect 3916 24044 3956 24053
rect 3628 23657 3668 23752
rect 3724 23624 3764 23719
rect 3724 23575 3764 23584
rect 3916 23624 3956 24004
rect 4108 23960 4148 33100
rect 4204 33032 4244 33041
rect 4204 31772 4244 32992
rect 4300 33032 4340 34084
rect 4396 33116 4436 34420
rect 4492 33200 4532 35428
rect 4492 33151 4532 33160
rect 4588 35888 4628 35897
rect 4396 33067 4436 33076
rect 4300 32983 4340 32992
rect 4396 32948 4436 32957
rect 4204 31723 4244 31732
rect 4300 32780 4340 32789
rect 4300 31604 4340 32740
rect 4204 31436 4244 31445
rect 4204 31100 4244 31396
rect 4204 31051 4244 31060
rect 4300 30764 4340 31564
rect 4300 30715 4340 30724
rect 4204 30512 4244 30521
rect 4204 30092 4244 30472
rect 4204 30043 4244 30052
rect 4300 30344 4340 30353
rect 4300 29924 4340 30304
rect 4204 29884 4340 29924
rect 4204 28580 4244 29884
rect 4300 29756 4340 29765
rect 4300 29168 4340 29716
rect 4300 29119 4340 29128
rect 4204 28531 4244 28540
rect 4300 29000 4340 29009
rect 4300 28496 4340 28960
rect 4300 28447 4340 28456
rect 4396 28076 4436 32908
rect 4492 32948 4532 32957
rect 4492 31688 4532 32908
rect 4588 32864 4628 35848
rect 4588 32815 4628 32824
rect 4492 31639 4532 31648
rect 4588 32696 4628 32705
rect 4492 31016 4532 31025
rect 4492 30848 4532 30976
rect 4492 30799 4532 30808
rect 4492 30680 4532 30689
rect 4492 30596 4532 30640
rect 4492 30545 4532 30556
rect 4588 30260 4628 32656
rect 4492 30220 4628 30260
rect 4492 29756 4532 30220
rect 4492 28412 4532 29716
rect 4492 28363 4532 28372
rect 4588 29672 4628 29681
rect 4588 28412 4628 29632
rect 4588 28363 4628 28372
rect 4588 28160 4628 28169
rect 4396 28036 4532 28076
rect 4204 27404 4244 27413
rect 4204 25724 4244 27364
rect 4300 26312 4340 26321
rect 4300 25724 4340 26272
rect 4492 26144 4532 28036
rect 4588 28025 4628 28120
rect 4588 27656 4628 27665
rect 4588 27152 4628 27616
rect 4684 27572 4724 36520
rect 4780 35720 4820 37444
rect 4928 36308 5296 36317
rect 4968 36268 5010 36308
rect 5050 36268 5092 36308
rect 5132 36268 5174 36308
rect 5214 36268 5256 36308
rect 4928 36259 5296 36268
rect 5356 35888 5396 39292
rect 5452 38996 5492 43828
rect 5548 43364 5588 48868
rect 5644 48740 5684 48749
rect 5644 48605 5684 48700
rect 5740 48068 5780 50044
rect 6124 49580 6164 53740
rect 6124 49531 6164 49540
rect 6220 49412 6260 54076
rect 6316 53948 6356 53957
rect 6316 52604 6356 53908
rect 6316 51680 6356 52564
rect 6316 51631 6356 51640
rect 6220 49363 6260 49372
rect 6124 48908 6164 48917
rect 6124 48740 6164 48868
rect 6124 48691 6164 48700
rect 5740 48019 5780 48028
rect 5836 48488 5876 48497
rect 5644 47060 5684 47069
rect 5644 45968 5684 47020
rect 5644 45128 5684 45928
rect 5740 46052 5780 46061
rect 5740 45212 5780 46012
rect 5740 45163 5780 45172
rect 5644 45079 5684 45088
rect 5548 43315 5588 43324
rect 5644 44540 5684 44549
rect 5548 43112 5588 43121
rect 5548 39752 5588 43072
rect 5644 42692 5684 44500
rect 5740 44372 5780 44381
rect 5740 43532 5780 44332
rect 5836 43868 5876 48448
rect 6412 48236 6452 55672
rect 6508 55544 6548 72808
rect 6604 72008 6644 72892
rect 6700 72260 6740 74488
rect 6796 73520 6836 78436
rect 6892 78308 6932 78317
rect 6892 77468 6932 78268
rect 6892 76544 6932 77428
rect 6892 76495 6932 76504
rect 6988 75956 7028 79360
rect 6988 75907 7028 75916
rect 6796 73471 6836 73480
rect 6892 75872 6932 75881
rect 6796 73268 6836 73277
rect 6796 72428 6836 73228
rect 6796 72379 6836 72388
rect 6740 72220 6836 72260
rect 6700 72211 6740 72220
rect 6604 71420 6644 71968
rect 6604 70916 6644 71380
rect 6604 70867 6644 70876
rect 6700 72008 6740 72017
rect 6604 70580 6644 70589
rect 6604 66716 6644 70540
rect 6700 68984 6740 71968
rect 6796 70832 6836 72220
rect 6892 72176 6932 75832
rect 6988 75788 7028 75797
rect 6988 75284 7028 75748
rect 6988 75235 7028 75244
rect 6988 75116 7028 75125
rect 6988 74024 7028 75076
rect 7084 74612 7124 79444
rect 7180 78476 7220 81292
rect 7276 80912 7316 81964
rect 7372 81332 7412 82300
rect 7468 82172 7508 82181
rect 7468 81836 7508 82132
rect 7564 82004 7604 82972
rect 7564 81955 7604 81964
rect 7468 81796 7604 81836
rect 7372 81283 7412 81292
rect 7468 81668 7508 81677
rect 7276 80863 7316 80872
rect 7468 80324 7508 81628
rect 7564 81080 7604 81796
rect 7660 81416 7700 83308
rect 7660 81367 7700 81376
rect 7564 81031 7604 81040
rect 7660 81248 7700 81257
rect 7372 80240 7412 80249
rect 7276 79988 7316 79997
rect 7276 79568 7316 79948
rect 7372 79820 7412 80200
rect 7468 79988 7508 80284
rect 7468 79939 7508 79948
rect 7564 80240 7604 80249
rect 7372 79771 7412 79780
rect 7468 79736 7508 79745
rect 7468 79601 7508 79696
rect 7276 79519 7316 79528
rect 7468 79064 7508 79073
rect 7180 77552 7220 78436
rect 7372 78560 7412 78569
rect 7180 77503 7220 77512
rect 7276 77888 7316 77897
rect 7084 74563 7124 74572
rect 7180 77300 7220 77309
rect 6988 73975 7028 73984
rect 7084 74444 7124 74453
rect 7084 73856 7124 74404
rect 6892 72092 6932 72136
rect 6892 72012 6932 72052
rect 6988 73816 7084 73856
rect 6988 72428 7028 73816
rect 7084 73807 7124 73816
rect 7180 73772 7220 77260
rect 7180 73723 7220 73732
rect 7084 73604 7124 73613
rect 7084 73184 7124 73564
rect 7084 73135 7124 73144
rect 7180 73436 7220 73445
rect 7180 73016 7220 73396
rect 6796 70783 6836 70792
rect 6988 70076 7028 72388
rect 6700 68935 6740 68944
rect 6796 70036 7028 70076
rect 7084 72976 7220 73016
rect 6604 66667 6644 66676
rect 6604 66128 6644 66137
rect 6644 66088 6740 66128
rect 6604 66079 6644 66088
rect 6604 65960 6644 65969
rect 6604 63188 6644 65920
rect 6700 65288 6740 66088
rect 6700 65239 6740 65248
rect 6700 63944 6740 63953
rect 6700 63524 6740 63904
rect 6700 63475 6740 63484
rect 6700 63356 6740 63365
rect 6700 63221 6740 63316
rect 6604 62768 6644 63148
rect 6604 62719 6644 62728
rect 6700 63020 6740 63029
rect 6700 62600 6740 62980
rect 6700 62551 6740 62560
rect 6604 62180 6644 62189
rect 6604 59324 6644 62140
rect 6700 61844 6740 61853
rect 6700 61676 6740 61804
rect 6700 61627 6740 61636
rect 6604 59275 6644 59284
rect 6700 61508 6740 61517
rect 6700 59660 6740 61468
rect 6700 59156 6740 59620
rect 6604 59116 6740 59156
rect 6604 56384 6644 59116
rect 6604 56335 6644 56344
rect 6700 57980 6740 57989
rect 6508 52604 6548 55504
rect 6700 55628 6740 57940
rect 6604 53864 6644 53873
rect 6604 53276 6644 53824
rect 6700 53780 6740 55588
rect 6700 53731 6740 53740
rect 6604 53227 6644 53236
rect 6604 53108 6644 53117
rect 6604 52772 6644 53068
rect 6604 52723 6644 52732
rect 6508 52555 6548 52564
rect 6508 52436 6548 52445
rect 6508 51764 6548 52396
rect 6508 51715 6548 51724
rect 6508 51092 6548 51101
rect 6508 49496 6548 51052
rect 6508 49447 6548 49456
rect 6604 49328 6644 49337
rect 6604 48740 6644 49288
rect 6604 48691 6644 48700
rect 6796 48572 6836 70036
rect 6892 69908 6932 69917
rect 6892 69236 6932 69868
rect 6892 69187 6932 69196
rect 6988 69320 7028 69329
rect 6892 67724 6932 67733
rect 6892 66464 6932 67684
rect 6988 67472 7028 69280
rect 7084 67976 7124 72976
rect 7276 72764 7316 77848
rect 7372 75788 7412 78520
rect 7468 78308 7508 79024
rect 7468 78259 7508 78268
rect 7372 75739 7412 75748
rect 7468 76040 7508 76049
rect 7372 74360 7412 74369
rect 7372 73772 7412 74320
rect 7468 74276 7508 76000
rect 7468 74227 7508 74236
rect 7372 73723 7412 73732
rect 7564 73688 7604 80200
rect 7660 78896 7700 81208
rect 7660 74696 7700 78856
rect 7756 77468 7796 83812
rect 7852 81752 7892 81761
rect 7852 81500 7892 81712
rect 7852 81451 7892 81460
rect 7852 81332 7892 81341
rect 7852 80408 7892 81292
rect 7852 80359 7892 80368
rect 7852 79820 7892 79829
rect 7852 78980 7892 79780
rect 7852 78931 7892 78940
rect 7948 78224 7988 84064
rect 8044 83684 8084 84232
rect 8044 83635 8084 83644
rect 8140 84188 8180 84197
rect 7948 78175 7988 78184
rect 8044 83180 8084 83189
rect 7756 76796 7796 77428
rect 7756 76747 7796 76756
rect 7852 77552 7892 77561
rect 7852 76124 7892 77512
rect 8044 77468 8084 83140
rect 8140 82256 8180 84148
rect 8140 82207 8180 82216
rect 8140 81332 8180 81341
rect 8140 79820 8180 81292
rect 8236 80156 8276 86500
rect 8428 85952 8468 94648
rect 8524 94352 8564 96688
rect 8716 94940 8756 96688
rect 8716 94891 8756 94900
rect 8812 94688 8852 94697
rect 8812 94553 8852 94648
rect 8524 94303 8564 94312
rect 8908 94268 8948 96688
rect 9100 94940 9140 96688
rect 9100 94891 9140 94900
rect 8908 94219 8948 94228
rect 9292 94184 9332 96688
rect 9484 94940 9524 96688
rect 9484 94891 9524 94900
rect 9388 94688 9428 94697
rect 9388 94553 9428 94648
rect 9676 94268 9716 96688
rect 9868 94940 9908 96688
rect 9868 94891 9908 94900
rect 9772 94688 9812 94697
rect 9772 94553 9812 94648
rect 9676 94219 9716 94228
rect 9292 94135 9332 94144
rect 10060 94184 10100 96688
rect 10252 94940 10292 96688
rect 10252 94891 10292 94900
rect 10444 94268 10484 96688
rect 10636 94940 10676 96688
rect 10636 94891 10676 94900
rect 10732 94772 10772 94781
rect 10540 94688 10580 94697
rect 10540 94553 10580 94648
rect 10732 94637 10772 94732
rect 10444 94219 10484 94228
rect 10060 94135 10100 94144
rect 10828 94184 10868 96688
rect 11020 94940 11060 96688
rect 11020 94891 11060 94900
rect 11212 94940 11252 96688
rect 11212 94891 11252 94900
rect 11308 95024 11348 95033
rect 11212 94688 11252 94697
rect 11212 94553 11252 94648
rect 10828 94135 10868 94144
rect 9484 94100 9524 94109
rect 8620 93848 8660 93857
rect 8428 85903 8468 85912
rect 8524 88556 8564 88565
rect 8524 85784 8564 88516
rect 8620 88304 8660 93808
rect 8620 88255 8660 88264
rect 8716 92924 8756 92933
rect 8716 88892 8756 92884
rect 8716 88052 8756 88852
rect 9292 89564 9332 89573
rect 9292 88808 9332 89524
rect 8716 88003 8756 88012
rect 8908 88136 8948 88145
rect 8620 87968 8660 87977
rect 8620 86708 8660 87928
rect 8716 87548 8756 87557
rect 8716 87413 8756 87508
rect 8812 87212 8852 87221
rect 8620 86668 8756 86708
rect 8620 86540 8660 86549
rect 8620 86036 8660 86500
rect 8620 85987 8660 85996
rect 8716 86456 8756 86668
rect 8428 85744 8564 85784
rect 8620 85868 8660 85877
rect 8332 84944 8372 84953
rect 8332 84440 8372 84904
rect 8332 84391 8372 84400
rect 8332 84188 8372 84197
rect 8332 84053 8372 84148
rect 8332 83852 8372 83861
rect 8332 83516 8372 83812
rect 8332 83012 8372 83476
rect 8428 83180 8468 85744
rect 8524 85196 8564 85205
rect 8524 84944 8564 85156
rect 8524 84895 8564 84904
rect 8524 84776 8564 84785
rect 8524 84356 8564 84736
rect 8524 84307 8564 84316
rect 8524 84104 8564 84113
rect 8524 83600 8564 84064
rect 8524 83551 8564 83560
rect 8524 83432 8564 83441
rect 8524 83264 8564 83392
rect 8524 83215 8564 83224
rect 8428 83131 8468 83140
rect 8332 82963 8372 82972
rect 8524 82760 8564 82769
rect 8428 82676 8468 82685
rect 8428 82088 8468 82636
rect 8428 82039 8468 82048
rect 8428 81920 8468 81929
rect 8332 81836 8372 81845
rect 8332 81164 8372 81796
rect 8428 81332 8468 81880
rect 8428 81283 8468 81292
rect 8332 81124 8468 81164
rect 8428 80660 8468 81124
rect 8236 80107 8276 80116
rect 8332 80620 8468 80660
rect 8332 80492 8372 80620
rect 8236 79820 8276 79829
rect 8140 79780 8236 79820
rect 7756 76084 7892 76124
rect 7948 77428 8084 77468
rect 8140 79064 8180 79073
rect 7948 76124 7988 77428
rect 7756 75284 7796 76084
rect 7948 75989 7988 76084
rect 8044 77300 8084 77309
rect 8044 76880 8084 77260
rect 8140 76964 8180 79024
rect 8140 76915 8180 76924
rect 7756 75235 7796 75244
rect 7852 75956 7892 75965
rect 7660 74647 7700 74656
rect 7756 75032 7796 75041
rect 7660 74276 7700 74285
rect 7660 74141 7700 74236
rect 7756 73856 7796 74992
rect 7756 73807 7796 73816
rect 7852 73688 7892 75916
rect 7948 75452 7988 75461
rect 7948 75368 7988 75412
rect 7948 75317 7988 75328
rect 8044 75200 8084 76840
rect 8236 76796 8276 79780
rect 8332 77384 8372 80452
rect 8524 79652 8564 82720
rect 8332 77335 8372 77344
rect 8428 79612 8564 79652
rect 8428 78308 8468 79612
rect 8044 75151 8084 75160
rect 8140 76756 8276 76796
rect 7948 75032 7988 75041
rect 8140 75032 8180 76756
rect 8332 76712 8372 76721
rect 8236 76628 8276 76637
rect 8236 75284 8276 76588
rect 8332 76208 8372 76672
rect 8428 76712 8468 78268
rect 8524 79484 8564 79493
rect 8524 77972 8564 79444
rect 8524 77923 8564 77932
rect 8524 77468 8564 77477
rect 8524 77333 8564 77428
rect 8428 76663 8468 76672
rect 8332 76159 8372 76168
rect 8620 75620 8660 85828
rect 8716 85280 8756 86416
rect 8812 86036 8852 87172
rect 8908 86792 8948 88096
rect 9292 88052 9332 88768
rect 9292 88003 9332 88012
rect 9292 87884 9332 87893
rect 9196 87800 9236 87809
rect 8908 86743 8948 86752
rect 9100 87044 9140 87053
rect 8812 85868 8852 85996
rect 8812 85819 8852 85828
rect 9004 85784 9044 85793
rect 8716 85231 8756 85240
rect 8812 85700 8852 85709
rect 8716 83936 8756 83945
rect 8716 81584 8756 83896
rect 8812 82256 8852 85660
rect 8908 85616 8948 85625
rect 8908 84776 8948 85576
rect 8908 84356 8948 84736
rect 8908 84307 8948 84316
rect 9004 85112 9044 85744
rect 8812 82207 8852 82216
rect 8908 84188 8948 84197
rect 8908 82592 8948 84148
rect 8908 82088 8948 82552
rect 8908 82039 8948 82048
rect 8716 81535 8756 81544
rect 8812 82004 8852 82013
rect 8524 75580 8660 75620
rect 8716 81416 8756 81425
rect 8428 75452 8468 75463
rect 8428 75368 8468 75412
rect 8428 75319 8468 75328
rect 8236 75235 8276 75244
rect 8428 75116 8468 75125
rect 8140 74992 8372 75032
rect 7948 74897 7988 74992
rect 7564 73639 7604 73648
rect 7756 73648 7892 73688
rect 7948 74612 7988 74621
rect 7948 74528 7988 74572
rect 7276 72715 7316 72724
rect 7276 72596 7316 72605
rect 7276 71336 7316 72556
rect 7372 72260 7412 72269
rect 7372 71504 7412 72220
rect 7372 71455 7412 71464
rect 7660 71672 7700 71681
rect 7276 71287 7316 71296
rect 7660 71168 7700 71632
rect 7660 71119 7700 71128
rect 7468 70916 7508 70925
rect 7180 70832 7220 70841
rect 7180 70697 7220 70792
rect 7372 70748 7412 70843
rect 7372 70699 7412 70708
rect 7276 70664 7316 70673
rect 7180 70496 7220 70505
rect 7180 69908 7220 70456
rect 7180 69859 7220 69868
rect 7180 69740 7220 69749
rect 7180 68480 7220 69700
rect 7276 69068 7316 70624
rect 7372 70580 7412 70589
rect 7372 69908 7412 70540
rect 7372 69859 7412 69868
rect 7468 69656 7508 70876
rect 7660 70916 7700 70925
rect 7564 70748 7604 70757
rect 7564 70076 7604 70708
rect 7660 70244 7700 70876
rect 7660 70195 7700 70204
rect 7604 70036 7700 70076
rect 7564 70027 7604 70036
rect 7372 69616 7508 69656
rect 7372 69488 7412 69616
rect 7372 69439 7412 69448
rect 7564 69404 7604 69413
rect 7564 69269 7604 69364
rect 7276 69019 7316 69028
rect 7372 69236 7412 69245
rect 7372 68816 7412 69196
rect 7372 68767 7412 68776
rect 7564 68984 7604 68993
rect 7180 68345 7220 68440
rect 7276 68564 7316 68573
rect 7084 67927 7124 67936
rect 7180 68228 7220 68237
rect 6988 67423 7028 67432
rect 7180 67808 7220 68188
rect 6892 66415 6932 66424
rect 6988 66380 7028 66389
rect 6892 66212 6932 66221
rect 6892 66128 6932 66172
rect 6892 66077 6932 66088
rect 6988 63524 7028 66340
rect 7180 66044 7220 67768
rect 7276 66380 7316 68524
rect 7468 68564 7508 68573
rect 7468 68480 7508 68524
rect 7468 68429 7508 68440
rect 7564 68480 7604 68944
rect 7564 68431 7604 68440
rect 7372 68396 7412 68405
rect 7372 66800 7412 68356
rect 7372 66751 7412 66760
rect 7468 68312 7508 68321
rect 7276 66331 7316 66340
rect 7372 66632 7412 66641
rect 7180 64700 7220 66004
rect 7180 64651 7220 64660
rect 7276 66212 7316 66221
rect 7276 64532 7316 66172
rect 6892 63484 7028 63524
rect 7180 64492 7316 64532
rect 6892 57812 6932 63484
rect 7180 63380 7220 64492
rect 6988 63340 7220 63380
rect 7276 63860 7316 63869
rect 6988 63272 7028 63340
rect 6988 63232 7124 63272
rect 6892 55796 6932 57772
rect 6988 63104 7028 63113
rect 6988 56804 7028 63064
rect 7084 62852 7124 63232
rect 7084 62803 7124 62812
rect 7084 62600 7124 62609
rect 7084 61676 7124 62560
rect 7084 61627 7124 61636
rect 7180 62516 7220 62525
rect 7084 61508 7124 61517
rect 7084 58064 7124 61468
rect 7180 58904 7220 62476
rect 7276 60836 7316 63820
rect 7372 62516 7412 66592
rect 7372 62467 7412 62476
rect 7372 62348 7412 62357
rect 7372 61844 7412 62308
rect 7468 62012 7508 68272
rect 7564 68060 7604 68069
rect 7564 63104 7604 68020
rect 7660 66968 7700 70036
rect 7660 66919 7700 66928
rect 7564 63055 7604 63064
rect 7660 66800 7700 66809
rect 7468 61963 7508 61972
rect 7564 62516 7604 62525
rect 7372 61795 7412 61804
rect 7564 61928 7604 62476
rect 7276 60500 7316 60796
rect 7276 60451 7316 60460
rect 7372 61676 7412 61685
rect 7372 60920 7412 61636
rect 7564 61004 7604 61888
rect 7564 60955 7604 60964
rect 7276 59912 7316 59921
rect 7276 59324 7316 59872
rect 7276 59275 7316 59284
rect 7180 58855 7220 58864
rect 7084 58024 7220 58064
rect 6988 56755 7028 56764
rect 7084 57896 7124 57905
rect 6892 55747 6932 55756
rect 6892 54788 6932 54797
rect 6892 53444 6932 54748
rect 6892 53192 6932 53404
rect 6988 53696 7028 53705
rect 6988 53300 7028 53656
rect 6988 53251 7028 53260
rect 6892 53152 7028 53192
rect 6892 52772 6932 52781
rect 6892 52604 6932 52732
rect 6892 52555 6932 52564
rect 6796 48523 6836 48532
rect 6892 52436 6932 52445
rect 6412 48187 6452 48196
rect 6316 47732 6356 47741
rect 6220 46052 6260 46061
rect 5932 45716 5972 45725
rect 5932 45581 5972 45676
rect 6124 45716 6164 45725
rect 6028 45212 6068 45221
rect 5932 45172 6028 45212
rect 5932 44792 5972 45172
rect 6028 45163 6068 45172
rect 5932 44743 5972 44752
rect 6028 45044 6068 45053
rect 6028 44540 6068 45004
rect 6028 44491 6068 44500
rect 5932 44288 5972 44383
rect 5932 44239 5972 44248
rect 5836 43819 5876 43828
rect 5932 44120 5972 44129
rect 5740 43483 5780 43492
rect 5836 43616 5876 43625
rect 5644 42643 5684 42652
rect 5740 43364 5780 43373
rect 5644 41936 5684 41945
rect 5644 40508 5684 41896
rect 5644 40459 5684 40468
rect 5644 40340 5684 40349
rect 5644 40256 5684 40300
rect 5644 40205 5684 40216
rect 5548 39712 5684 39752
rect 5644 39332 5684 39712
rect 5644 39283 5684 39292
rect 5452 38947 5492 38956
rect 5548 39164 5588 39173
rect 5740 39164 5780 43324
rect 5836 42860 5876 43576
rect 5932 42944 5972 44080
rect 5932 42895 5972 42904
rect 6028 43532 6068 43541
rect 5836 42811 5876 42820
rect 6028 42860 6068 43492
rect 6124 43364 6164 45676
rect 6220 45296 6260 46012
rect 6220 45247 6260 45256
rect 6316 45128 6356 47692
rect 6700 46556 6740 46565
rect 6604 46304 6644 46313
rect 6412 45968 6452 45977
rect 6412 45716 6452 45928
rect 6412 45667 6452 45676
rect 6604 45716 6644 46264
rect 6700 46136 6740 46516
rect 6700 46087 6740 46096
rect 6604 45667 6644 45676
rect 6796 45800 6836 45811
rect 6796 45716 6836 45760
rect 6796 45667 6836 45676
rect 6700 45632 6740 45641
rect 6700 45497 6740 45592
rect 6604 45464 6644 45473
rect 6316 45079 6356 45088
rect 6412 45380 6452 45389
rect 6316 44792 6356 44801
rect 6124 43315 6164 43324
rect 6220 44624 6260 44633
rect 6028 42776 6068 42820
rect 5932 42736 6068 42776
rect 5932 41936 5972 42736
rect 6028 42725 6068 42736
rect 6124 42944 6164 42953
rect 6124 42692 6164 42904
rect 5932 41887 5972 41896
rect 6028 42608 6068 42617
rect 5836 41852 5876 41861
rect 5836 39836 5876 41812
rect 6028 41180 6068 42568
rect 6124 41348 6164 42652
rect 6220 42020 6260 44584
rect 6316 44204 6356 44752
rect 6412 44708 6452 45340
rect 6412 44659 6452 44668
rect 6412 44540 6452 44549
rect 6412 44288 6452 44500
rect 6412 44239 6452 44248
rect 6508 44372 6548 44381
rect 6508 44237 6548 44332
rect 6316 44155 6356 44164
rect 6508 43616 6548 43625
rect 6412 43448 6452 43457
rect 6316 43028 6356 43039
rect 6316 42944 6356 42988
rect 6316 42895 6356 42904
rect 6412 42692 6452 43408
rect 6412 42643 6452 42652
rect 6508 43448 6548 43576
rect 6508 42776 6548 43408
rect 6220 41971 6260 41980
rect 6508 41432 6548 42736
rect 6508 41383 6548 41392
rect 6124 41299 6164 41308
rect 6508 41264 6548 41273
rect 6508 41180 6548 41224
rect 6028 41045 6068 41140
rect 6412 41140 6548 41180
rect 6124 41096 6164 41105
rect 5836 39787 5876 39796
rect 5932 41012 5972 41021
rect 5932 39668 5972 40972
rect 6028 40844 6068 40853
rect 6028 40760 6068 40804
rect 6028 40709 6068 40720
rect 6028 40508 6068 40603
rect 6028 40459 6068 40468
rect 6124 40592 6164 41056
rect 6316 41096 6356 41105
rect 6220 41012 6260 41021
rect 6220 40676 6260 40972
rect 6220 40627 6260 40636
rect 6124 40340 6164 40552
rect 5932 39619 5972 39628
rect 6028 40300 6164 40340
rect 6220 40508 6260 40517
rect 6028 39584 6068 40300
rect 6124 40004 6164 40015
rect 6124 39920 6164 39964
rect 6124 39871 6164 39880
rect 5452 38576 5492 38585
rect 5452 38492 5492 38536
rect 5452 38441 5492 38452
rect 5548 38240 5588 39124
rect 5548 38191 5588 38200
rect 5644 39124 5780 39164
rect 5836 39500 5876 39509
rect 5644 38072 5684 39124
rect 5548 38032 5684 38072
rect 5740 38996 5780 39005
rect 5452 37988 5492 37997
rect 5452 37652 5492 37948
rect 5452 37603 5492 37612
rect 5452 36980 5492 36989
rect 5452 36845 5492 36940
rect 5356 35839 5396 35848
rect 4780 35671 4820 35680
rect 5356 35720 5396 35729
rect 5164 35552 5204 35561
rect 4780 35300 4820 35309
rect 4780 34292 4820 35260
rect 5164 35132 5204 35512
rect 5164 35083 5204 35092
rect 5356 35048 5396 35680
rect 4928 34796 5296 34805
rect 4968 34756 5010 34796
rect 5050 34756 5092 34796
rect 5132 34756 5174 34796
rect 5214 34756 5256 34796
rect 4928 34747 5296 34756
rect 4972 34628 5012 34637
rect 4780 34040 4820 34252
rect 4780 33991 4820 34000
rect 4876 34460 4916 34469
rect 4876 33788 4916 34420
rect 4972 34376 5012 34588
rect 5260 34628 5300 34637
rect 5260 34460 5300 34588
rect 5260 34411 5300 34420
rect 4972 34327 5012 34336
rect 4780 33748 4916 33788
rect 4780 32108 4820 33748
rect 4928 33284 5296 33293
rect 4968 33244 5010 33284
rect 5050 33244 5092 33284
rect 5132 33244 5174 33284
rect 5214 33244 5256 33284
rect 4928 33235 5296 33244
rect 5164 32948 5204 32957
rect 5164 32360 5204 32908
rect 5164 32311 5204 32320
rect 5260 32864 5300 32873
rect 4780 30092 4820 32068
rect 5260 31940 5300 32824
rect 5260 31891 5300 31900
rect 4928 31772 5296 31781
rect 4968 31732 5010 31772
rect 5050 31732 5092 31772
rect 5132 31732 5174 31772
rect 5214 31732 5256 31772
rect 4928 31723 5296 31732
rect 5164 31604 5204 31613
rect 5164 31436 5204 31564
rect 4876 31100 4916 31109
rect 4876 31016 4916 31060
rect 4876 30965 4916 30976
rect 5068 30932 5108 30941
rect 5068 30596 5108 30892
rect 5164 30848 5204 31396
rect 5260 31520 5300 31529
rect 5260 31385 5300 31480
rect 5164 30799 5204 30808
rect 5068 30461 5108 30556
rect 4928 30260 5296 30269
rect 4968 30220 5010 30260
rect 5050 30220 5092 30260
rect 5132 30220 5174 30260
rect 5214 30220 5256 30260
rect 4928 30211 5296 30220
rect 4780 30052 4916 30092
rect 4876 30008 4916 30052
rect 4780 29924 4820 29933
rect 4780 28664 4820 29884
rect 4876 29336 4916 29968
rect 4876 29287 4916 29296
rect 5260 30008 5300 30017
rect 4876 28916 4916 29011
rect 4876 28867 4916 28876
rect 5260 28916 5300 29968
rect 5260 28867 5300 28876
rect 4928 28748 5296 28757
rect 4968 28708 5010 28748
rect 5050 28708 5092 28748
rect 5132 28708 5174 28748
rect 5214 28708 5256 28748
rect 4928 28699 5296 28708
rect 4780 28615 4820 28624
rect 4876 28580 4916 28589
rect 4780 28412 4820 28421
rect 4780 28277 4820 28372
rect 4876 27656 4916 28540
rect 5068 28580 5108 28589
rect 5068 28412 5108 28540
rect 5260 28580 5300 28589
rect 5260 28445 5300 28540
rect 5068 28363 5108 28372
rect 4876 27607 4916 27616
rect 5260 27740 5300 27749
rect 4684 27532 4820 27572
rect 4588 27103 4628 27112
rect 4684 27404 4724 27413
rect 4492 26095 4532 26104
rect 4588 26984 4628 26993
rect 4588 26060 4628 26944
rect 4300 25684 4532 25724
rect 4204 25675 4244 25684
rect 4300 25556 4340 25565
rect 4300 24548 4340 25516
rect 4300 24499 4340 24508
rect 4300 24380 4340 24389
rect 4108 23920 4244 23960
rect 4012 23876 4052 23885
rect 4052 23836 4148 23876
rect 4012 23827 4052 23836
rect 3916 23575 3956 23584
rect 3688 23456 4056 23465
rect 3728 23416 3770 23456
rect 3810 23416 3852 23456
rect 3892 23416 3934 23456
rect 3974 23416 4016 23456
rect 3688 23407 4056 23416
rect 3532 22987 3572 22996
rect 3628 23288 3668 23297
rect 3436 22483 3476 22492
rect 3532 22868 3572 22877
rect 3436 22364 3476 22373
rect 3436 22229 3476 22324
rect 3532 22280 3572 22828
rect 3532 22231 3572 22240
rect 3340 20047 3380 20056
rect 3436 22112 3476 22121
rect 3628 22112 3668 23248
rect 3820 23288 3860 23297
rect 3436 19928 3476 22072
rect 3532 22072 3668 22112
rect 3724 23204 3764 23213
rect 3724 22112 3764 23164
rect 3820 22196 3860 23248
rect 4012 23288 4052 23297
rect 3820 22147 3860 22156
rect 3916 23120 3956 23129
rect 3916 22196 3956 23080
rect 4012 22952 4052 23248
rect 4012 22903 4052 22912
rect 3916 22147 3956 22156
rect 4108 22364 4148 23836
rect 4204 23288 4244 23920
rect 4204 23239 4244 23248
rect 4300 23120 4340 24340
rect 4300 23071 4340 23080
rect 4396 23540 4436 23549
rect 4300 22952 4340 22961
rect 3532 21524 3572 22072
rect 3724 22063 3764 22072
rect 3688 21944 4056 21953
rect 3728 21904 3770 21944
rect 3810 21904 3852 21944
rect 3892 21904 3934 21944
rect 3974 21904 4016 21944
rect 3688 21895 4056 21904
rect 3820 21776 3860 21785
rect 3820 21692 3860 21736
rect 3628 21524 3668 21533
rect 3532 21484 3628 21524
rect 3628 21475 3668 21484
rect 3436 19879 3476 19888
rect 3532 21356 3572 21365
rect 3532 20264 3572 21316
rect 3820 20852 3860 21652
rect 3820 20803 3860 20812
rect 3916 21608 3956 21617
rect 3628 20684 3668 20779
rect 3916 20768 3956 21568
rect 4012 21608 4052 21617
rect 4012 21020 4052 21568
rect 4012 20971 4052 20980
rect 3916 20719 3956 20728
rect 3628 20635 3668 20644
rect 3688 20432 4056 20441
rect 3728 20392 3770 20432
rect 3810 20392 3852 20432
rect 3892 20392 3934 20432
rect 3974 20392 4016 20432
rect 3688 20383 4056 20392
rect 3532 19592 3572 20224
rect 3244 18535 3284 18544
rect 3340 19552 3572 19592
rect 3628 19928 3668 19937
rect 3340 18500 3380 19552
rect 3532 19340 3572 19349
rect 3436 19088 3476 19097
rect 3436 18752 3476 19048
rect 3532 18920 3572 19300
rect 3628 19256 3668 19888
rect 3628 19121 3668 19216
rect 3532 18871 3572 18880
rect 3688 18920 4056 18929
rect 3728 18880 3770 18920
rect 3810 18880 3852 18920
rect 3892 18880 3934 18920
rect 3974 18880 4016 18920
rect 3688 18871 4056 18880
rect 3532 18752 3572 18761
rect 3436 18712 3532 18752
rect 3244 18416 3284 18427
rect 3244 18332 3284 18376
rect 3244 18283 3284 18292
rect 3148 15427 3188 15436
rect 3244 17828 3284 17837
rect 2956 15392 2996 15401
rect 2860 13964 2900 13973
rect 2860 13829 2900 13924
rect 2764 13672 2900 13712
rect 2764 13544 2804 13553
rect 2764 12284 2804 13504
rect 2764 12235 2804 12244
rect 2860 13040 2900 13672
rect 2860 11780 2900 13000
rect 2668 11143 2708 11152
rect 2764 11740 2860 11780
rect 2764 10940 2804 11740
rect 2860 11712 2900 11740
rect 2860 11612 2900 11621
rect 2860 11477 2900 11572
rect 2956 11024 2996 15352
rect 3148 15308 3188 15317
rect 3148 13544 3188 15268
rect 3148 13495 3188 13504
rect 3244 13460 3284 17788
rect 3340 17492 3380 18460
rect 3532 17828 3572 18712
rect 4012 18500 4052 18509
rect 3628 18416 3668 18425
rect 3628 18281 3668 18376
rect 4012 17996 4052 18460
rect 4012 17947 4052 17956
rect 3340 17443 3380 17452
rect 3436 17788 3532 17828
rect 3340 17324 3380 17333
rect 3340 16484 3380 17284
rect 3436 17156 3476 17788
rect 3532 17779 3572 17788
rect 3916 17828 3956 17837
rect 3916 17693 3956 17788
rect 4012 17744 4052 17753
rect 4012 17609 4052 17704
rect 3436 17107 3476 17116
rect 3532 17492 3572 17501
rect 3340 16435 3380 16444
rect 3436 16988 3476 16997
rect 3340 16316 3380 16325
rect 3340 14972 3380 16276
rect 3340 14923 3380 14932
rect 3244 13411 3284 13420
rect 3340 14300 3380 14309
rect 3340 14048 3380 14260
rect 3148 13376 3188 13385
rect 3052 13040 3092 13049
rect 3052 12536 3092 13000
rect 3052 12487 3092 12496
rect 2956 10975 2996 10984
rect 3052 12368 3092 12377
rect 2764 10891 2804 10900
rect 2572 8875 2612 8884
rect 2668 10688 2708 10697
rect 2476 8707 2516 8716
rect 2380 5599 2420 5608
rect 2380 4976 2420 4985
rect 2380 4472 2420 4936
rect 2380 4423 2420 4432
rect 2188 4087 2228 4096
rect 1996 4052 2036 4061
rect 1804 3212 1844 3221
rect 1804 2792 1844 3172
rect 1804 2743 1844 2752
rect 1900 3128 1940 3137
rect 1708 2575 1748 2584
rect 1900 1784 1940 3088
rect 1804 1744 1940 1784
rect 1804 80 1844 1744
rect 1996 80 2036 4012
rect 2188 3632 2228 3641
rect 2092 2624 2132 2633
rect 2092 2489 2132 2584
rect 2188 80 2228 3592
rect 2668 3548 2708 10648
rect 2860 10520 2900 10529
rect 2764 10268 2804 10277
rect 2764 8168 2804 10228
rect 2860 10184 2900 10480
rect 2860 10135 2900 10144
rect 2956 10436 2996 10445
rect 2956 10016 2996 10396
rect 2956 9965 2996 9976
rect 2956 8504 2996 8513
rect 2860 8168 2900 8177
rect 2764 8128 2860 8168
rect 2860 8100 2900 8128
rect 2764 7916 2804 7925
rect 2764 7244 2804 7876
rect 2764 6656 2804 7204
rect 2860 7160 2900 7169
rect 2860 6908 2900 7120
rect 2860 6859 2900 6868
rect 2764 6607 2804 6616
rect 2860 6320 2900 6329
rect 2860 6185 2900 6280
rect 2668 3499 2708 3508
rect 2380 3464 2420 3473
rect 2380 3329 2420 3424
rect 2956 2900 2996 8464
rect 3052 4388 3092 12328
rect 3148 9680 3188 13336
rect 3340 13376 3380 14008
rect 3340 13327 3380 13336
rect 3436 13292 3476 16948
rect 3532 13460 3572 17452
rect 3688 17408 4056 17417
rect 3728 17368 3770 17408
rect 3810 17368 3852 17408
rect 3892 17368 3934 17408
rect 3974 17368 4016 17408
rect 3688 17359 4056 17368
rect 3820 17156 3860 17165
rect 3628 16988 3668 16997
rect 3628 16232 3668 16948
rect 3820 16904 3860 17116
rect 4012 17072 4052 17081
rect 4108 17072 4148 22324
rect 4204 22784 4244 22793
rect 4204 21440 4244 22744
rect 4300 21608 4340 22912
rect 4396 22280 4436 23500
rect 4396 22231 4436 22240
rect 4300 21559 4340 21568
rect 4396 21776 4436 21785
rect 4204 19508 4244 21400
rect 4204 19459 4244 19468
rect 4300 21440 4340 21449
rect 4204 19340 4244 19349
rect 4300 19340 4340 21400
rect 4396 20012 4436 21736
rect 4396 19963 4436 19972
rect 4244 19300 4340 19340
rect 4396 19844 4436 19853
rect 4204 19088 4244 19300
rect 4396 19172 4436 19804
rect 4396 19123 4436 19132
rect 4204 18332 4244 19048
rect 4300 18920 4340 18929
rect 4300 18584 4340 18880
rect 4492 18584 4532 25684
rect 4588 24800 4628 26020
rect 4684 26060 4724 27364
rect 4684 26011 4724 26020
rect 4588 24751 4628 24760
rect 4684 25892 4724 25901
rect 4588 24548 4628 24557
rect 4588 23060 4628 24508
rect 4684 23876 4724 25852
rect 4684 23827 4724 23836
rect 4684 23624 4724 23633
rect 4684 23372 4724 23584
rect 4684 23323 4724 23332
rect 4588 23020 4724 23060
rect 4588 22364 4628 22373
rect 4588 22196 4628 22324
rect 4588 21440 4628 22156
rect 4588 21391 4628 21400
rect 4300 18535 4340 18544
rect 4396 18544 4532 18584
rect 4588 20768 4628 20777
rect 4588 18584 4628 20728
rect 4204 18283 4244 18292
rect 4052 17032 4148 17072
rect 4012 17023 4052 17032
rect 3628 16183 3668 16192
rect 3724 16568 3764 16577
rect 3724 16148 3764 16528
rect 3820 16316 3860 16864
rect 3820 16267 3860 16276
rect 4108 16316 4148 17032
rect 4204 17156 4244 17165
rect 4204 16652 4244 17116
rect 4300 16988 4340 17083
rect 4300 16939 4340 16948
rect 4204 16603 4244 16612
rect 4300 16820 4340 16829
rect 3724 16099 3764 16108
rect 3688 15896 4056 15905
rect 3728 15856 3770 15896
rect 3810 15856 3852 15896
rect 3892 15856 3934 15896
rect 3974 15856 4016 15896
rect 3688 15847 4056 15856
rect 3628 15644 3668 15653
rect 3628 15476 3668 15604
rect 3628 15427 3668 15436
rect 3628 15056 3668 15065
rect 3628 14804 3668 15016
rect 3628 14755 3668 14764
rect 3688 14384 4056 14393
rect 3728 14344 3770 14384
rect 3810 14344 3852 14384
rect 3892 14344 3934 14384
rect 3974 14344 4016 14384
rect 3688 14335 4056 14344
rect 4108 14216 4148 16276
rect 4300 15896 4340 16780
rect 4300 15847 4340 15856
rect 4012 14176 4148 14216
rect 4204 15644 4244 15653
rect 3532 13411 3572 13420
rect 3628 13964 3668 13973
rect 3628 13292 3668 13924
rect 3436 13243 3476 13252
rect 3532 13252 3668 13292
rect 3340 13208 3380 13217
rect 3340 12872 3380 13168
rect 3340 12823 3380 12832
rect 3532 12620 3572 13252
rect 4012 13040 4052 14176
rect 4012 12991 4052 13000
rect 4108 13964 4148 13973
rect 3688 12872 4056 12881
rect 3728 12832 3770 12872
rect 3810 12832 3852 12872
rect 3892 12832 3934 12872
rect 3974 12832 4016 12872
rect 3688 12823 4056 12832
rect 3916 12704 3956 12713
rect 3532 12571 3572 12580
rect 3724 12620 3764 12629
rect 3340 12536 3380 12545
rect 3244 12452 3284 12461
rect 3244 10352 3284 12412
rect 3244 10303 3284 10312
rect 3148 9631 3188 9640
rect 3340 9008 3380 12496
rect 3724 12536 3764 12580
rect 3724 12485 3764 12496
rect 3628 12452 3668 12461
rect 3532 12412 3628 12452
rect 3436 11192 3476 11201
rect 3436 11057 3476 11152
rect 3436 10268 3476 10277
rect 3436 10184 3476 10228
rect 3436 10133 3476 10144
rect 3244 8968 3380 9008
rect 3436 9764 3476 9773
rect 3148 7748 3188 7757
rect 3148 6656 3188 7708
rect 3148 6607 3188 6616
rect 3148 5564 3188 5573
rect 3148 5429 3188 5524
rect 3148 5144 3188 5153
rect 3148 4808 3188 5104
rect 3148 4759 3188 4768
rect 3052 4339 3092 4348
rect 3052 3548 3092 3557
rect 3244 3548 3284 8968
rect 3340 8840 3380 8849
rect 3340 6572 3380 8800
rect 3436 8756 3476 9724
rect 3532 9596 3572 12412
rect 3628 12403 3668 12412
rect 3916 11612 3956 12664
rect 4108 11948 4148 13924
rect 4108 11899 4148 11908
rect 4012 11864 4052 11873
rect 4012 11780 4052 11824
rect 4204 11780 4244 15604
rect 4300 15476 4340 15485
rect 4300 14972 4340 15436
rect 4300 14636 4340 14932
rect 4300 13460 4340 14596
rect 4396 14048 4436 18544
rect 4588 18535 4628 18544
rect 4684 17996 4724 23020
rect 4780 23036 4820 27532
rect 5260 27488 5300 27700
rect 5260 27439 5300 27448
rect 4928 27236 5296 27245
rect 4968 27196 5010 27236
rect 5050 27196 5092 27236
rect 5132 27196 5174 27236
rect 5214 27196 5256 27236
rect 4928 27187 5296 27196
rect 5356 26312 5396 35008
rect 5452 34040 5492 34049
rect 5452 32108 5492 34000
rect 5548 33140 5588 38032
rect 5644 36224 5684 36233
rect 5644 34040 5684 36184
rect 5740 35804 5780 38956
rect 5836 38324 5876 39460
rect 6028 39416 6068 39544
rect 6220 39584 6260 40468
rect 6316 40424 6356 41056
rect 6316 40375 6356 40384
rect 6316 40256 6356 40265
rect 6316 39668 6356 40216
rect 6412 39920 6452 41140
rect 6604 41096 6644 45424
rect 6892 45380 6932 52396
rect 6988 51848 7028 53152
rect 7084 52856 7124 57856
rect 7180 54704 7220 58024
rect 7372 56552 7412 60880
rect 7180 54655 7220 54664
rect 7276 56512 7412 56552
rect 7468 60500 7508 60509
rect 7276 55376 7316 56512
rect 7276 54284 7316 55336
rect 7276 54235 7316 54244
rect 7372 56384 7412 56393
rect 7180 54116 7220 54125
rect 7220 54076 7316 54116
rect 7180 54067 7220 54076
rect 7180 53948 7220 53957
rect 7180 53360 7220 53908
rect 7180 53311 7220 53320
rect 7276 53444 7316 54076
rect 7276 53276 7316 53404
rect 7276 53227 7316 53236
rect 7084 52807 7124 52816
rect 7180 53192 7220 53201
rect 7084 51848 7124 51857
rect 6988 51808 7084 51848
rect 7084 51799 7124 51808
rect 6988 51680 7028 51689
rect 6988 51545 7028 51640
rect 7180 51008 7220 53152
rect 7372 52688 7412 56344
rect 7372 52639 7412 52648
rect 7180 50959 7220 50968
rect 7180 49580 7220 49589
rect 7180 48740 7220 49540
rect 7180 48691 7220 48700
rect 7468 48152 7508 60460
rect 7564 59072 7604 59081
rect 7564 50756 7604 59032
rect 7660 55712 7700 66760
rect 7756 65288 7796 73648
rect 7852 72260 7892 72269
rect 7852 71672 7892 72220
rect 7852 71623 7892 71632
rect 7852 71504 7892 71513
rect 7852 68564 7892 71464
rect 7852 68515 7892 68524
rect 7948 68396 7988 74488
rect 8044 74360 8084 74369
rect 8044 74024 8084 74320
rect 8236 74192 8276 74201
rect 8236 74108 8276 74152
rect 8236 74057 8276 74068
rect 8140 74024 8180 74052
rect 8044 73984 8140 74024
rect 8044 72428 8084 73984
rect 8140 73975 8180 73984
rect 8332 73940 8372 74992
rect 8428 74696 8468 75076
rect 8428 74647 8468 74656
rect 8236 73900 8372 73940
rect 8140 73688 8180 73697
rect 8140 73184 8180 73648
rect 8140 73135 8180 73144
rect 8140 73016 8180 73025
rect 8140 72881 8180 72976
rect 8044 72388 8180 72428
rect 8044 71420 8084 71429
rect 8044 69404 8084 71380
rect 8140 70160 8180 72388
rect 8140 70111 8180 70120
rect 8236 69992 8276 73900
rect 8428 73520 8468 73529
rect 8332 73480 8428 73520
rect 8332 72932 8372 73480
rect 8428 73471 8468 73480
rect 8332 72883 8372 72892
rect 8428 73352 8468 73361
rect 8236 69943 8276 69952
rect 8332 72764 8372 72773
rect 8044 69355 8084 69364
rect 8140 69824 8180 69833
rect 7756 64700 7796 65248
rect 7756 64651 7796 64660
rect 7852 68356 7988 68396
rect 8044 69236 8084 69245
rect 7756 64280 7796 64289
rect 7756 63944 7796 64240
rect 7756 63895 7796 63904
rect 7756 63692 7796 63701
rect 7756 63557 7796 63652
rect 7756 63188 7796 63197
rect 7756 62684 7796 63148
rect 7756 62635 7796 62644
rect 7756 62180 7796 62189
rect 7756 61592 7796 62140
rect 7756 61543 7796 61552
rect 7756 61004 7796 61013
rect 7756 57140 7796 60964
rect 7852 59576 7892 68356
rect 8044 67556 8084 69196
rect 8044 67507 8084 67516
rect 8140 66884 8180 69784
rect 8236 69740 8276 69749
rect 8236 69320 8276 69700
rect 8236 69185 8276 69280
rect 8236 69068 8276 69077
rect 8236 68480 8276 69028
rect 8236 68431 8276 68440
rect 8236 68228 8276 68237
rect 8236 68093 8276 68188
rect 8140 66835 8180 66844
rect 8236 67724 8276 67733
rect 7948 66212 7988 66221
rect 7948 65540 7988 66172
rect 7948 65491 7988 65500
rect 8140 64700 8180 64709
rect 7948 64364 7988 64373
rect 7948 63608 7988 64324
rect 7948 63559 7988 63568
rect 8044 63944 8084 63953
rect 7948 63440 7988 63449
rect 7948 60164 7988 63400
rect 8044 63188 8084 63904
rect 8140 63944 8180 64660
rect 8140 63895 8180 63904
rect 8236 63524 8276 67684
rect 8332 66716 8372 72724
rect 8428 67724 8468 73312
rect 8428 67675 8468 67684
rect 8332 63776 8372 66676
rect 8524 66632 8564 75580
rect 8620 75284 8660 75293
rect 8620 75149 8660 75244
rect 8716 74612 8756 81376
rect 8812 81332 8852 81964
rect 8812 81283 8852 81292
rect 8908 81920 8948 81929
rect 8908 81164 8948 81880
rect 8908 81115 8948 81124
rect 8908 80912 8948 80921
rect 8812 80156 8852 80165
rect 8812 79820 8852 80116
rect 8812 79568 8852 79780
rect 8812 79519 8852 79528
rect 8812 79148 8852 79157
rect 8812 76796 8852 79108
rect 8908 78980 8948 80872
rect 8908 76880 8948 78940
rect 8908 76831 8948 76840
rect 8812 75284 8852 76756
rect 8908 76124 8948 76133
rect 8908 75536 8948 76084
rect 8908 75487 8948 75496
rect 8908 75284 8948 75293
rect 8812 75244 8908 75284
rect 8908 75235 8948 75244
rect 8908 74780 8948 74789
rect 8908 74645 8948 74740
rect 8716 74572 8852 74612
rect 8716 74444 8756 74453
rect 8620 72932 8660 72941
rect 8620 72344 8660 72892
rect 8620 72295 8660 72304
rect 8620 72092 8660 72101
rect 8620 69908 8660 72052
rect 8716 71420 8756 74404
rect 8716 69992 8756 71380
rect 8716 69943 8756 69952
rect 8812 73016 8852 74572
rect 8620 69488 8660 69868
rect 8620 67052 8660 69448
rect 8716 68564 8756 68575
rect 8716 68480 8756 68524
rect 8716 68431 8756 68440
rect 8620 67003 8660 67012
rect 8524 66583 8564 66592
rect 8812 65708 8852 72976
rect 8908 73520 8948 73529
rect 8908 72932 8948 73480
rect 8908 72883 8948 72892
rect 8908 72092 8948 72101
rect 8908 70580 8948 72052
rect 9004 71924 9044 85072
rect 9100 82088 9140 87004
rect 9196 83936 9236 87760
rect 9292 86624 9332 87844
rect 9292 85028 9332 86584
rect 9292 84979 9332 84988
rect 9388 87128 9428 87137
rect 9196 83887 9236 83896
rect 9292 84860 9332 84869
rect 9292 83936 9332 84820
rect 9292 83887 9332 83896
rect 9292 83768 9332 83777
rect 9100 82039 9140 82048
rect 9196 83684 9236 83693
rect 9100 81584 9140 81593
rect 9100 78980 9140 81544
rect 9100 78308 9140 78940
rect 9100 78259 9140 78268
rect 9100 78140 9140 78151
rect 9100 78056 9140 78100
rect 9100 78007 9140 78016
rect 9100 77720 9140 77729
rect 9100 76712 9140 77680
rect 9100 76663 9140 76672
rect 9196 75956 9236 83644
rect 9292 80576 9332 83728
rect 9292 80527 9332 80536
rect 9292 80240 9332 80251
rect 9292 80156 9332 80200
rect 9292 80107 9332 80116
rect 9292 79652 9332 79661
rect 9292 79400 9332 79612
rect 9292 79351 9332 79360
rect 9100 75916 9236 75956
rect 9292 78896 9332 78905
rect 9100 74444 9140 75916
rect 9100 74395 9140 74404
rect 9196 75200 9236 75209
rect 9100 73520 9140 73615
rect 9100 73471 9140 73480
rect 9100 73016 9140 73025
rect 9100 72092 9140 72976
rect 9196 72428 9236 75160
rect 9292 73688 9332 78856
rect 9388 76880 9428 87088
rect 9484 81500 9524 94060
rect 9484 81451 9524 81460
rect 9580 94016 9620 94025
rect 9580 81248 9620 93976
rect 9964 94016 10004 94025
rect 9964 93881 10004 93976
rect 11020 94016 11060 94025
rect 10156 93932 10196 93941
rect 10156 93797 10196 93892
rect 10828 93932 10868 93941
rect 10828 93797 10868 93892
rect 11020 93881 11060 93976
rect 9676 91664 9716 91673
rect 9676 83768 9716 91624
rect 10828 91412 10868 91421
rect 9964 90992 10004 91001
rect 9676 83719 9716 83728
rect 9772 89396 9812 89405
rect 9772 84356 9812 89356
rect 9868 88640 9908 88649
rect 9868 87632 9908 88600
rect 9868 87583 9908 87592
rect 9772 81500 9812 84316
rect 9772 81451 9812 81460
rect 9868 85280 9908 85289
rect 9580 81208 9812 81248
rect 9484 81164 9524 81173
rect 9484 78980 9524 81124
rect 9484 78931 9524 78940
rect 9580 79988 9620 79997
rect 9484 78728 9524 78823
rect 9484 78679 9524 78688
rect 9388 76831 9428 76840
rect 9292 73639 9332 73648
rect 9388 76712 9428 76721
rect 9388 73460 9428 76672
rect 9484 75956 9524 75965
rect 9484 74696 9524 75916
rect 9484 74647 9524 74656
rect 9196 72379 9236 72388
rect 9292 73420 9428 73460
rect 9484 73856 9524 73865
rect 9100 72043 9140 72052
rect 9196 72176 9236 72185
rect 9004 71884 9140 71924
rect 8908 70531 8948 70540
rect 9004 70412 9044 70421
rect 9004 67640 9044 70372
rect 8908 67136 8948 67145
rect 8908 67001 8948 67096
rect 9004 66884 9044 67600
rect 8716 65668 8812 65708
rect 8524 65204 8564 65213
rect 8524 64700 8564 65164
rect 8620 65036 8660 65045
rect 8620 64901 8660 64996
rect 8428 64660 8524 64700
rect 8428 63944 8468 64660
rect 8524 64651 8564 64660
rect 8620 64532 8660 64541
rect 8620 64028 8660 64492
rect 8620 63979 8660 63988
rect 8428 63895 8468 63904
rect 8524 63860 8564 63869
rect 8332 63736 8468 63776
rect 8140 63484 8276 63524
rect 8140 63440 8180 63484
rect 8140 63391 8180 63400
rect 8332 63272 8372 63281
rect 8044 62432 8084 63148
rect 8236 63188 8276 63197
rect 8044 62383 8084 62392
rect 8140 63104 8180 63113
rect 7948 60115 7988 60124
rect 8044 60584 8084 60593
rect 8044 59576 8084 60544
rect 7852 59527 7892 59536
rect 7948 59536 8084 59576
rect 8140 59576 8180 63064
rect 8236 60332 8276 63148
rect 8332 60920 8372 63232
rect 8332 60871 8372 60880
rect 8236 60283 8276 60292
rect 8332 60752 8372 60761
rect 7852 59240 7892 59249
rect 7852 57812 7892 59200
rect 7852 57763 7892 57772
rect 7852 57140 7892 57149
rect 7756 57100 7852 57140
rect 7756 56384 7796 57100
rect 7852 57091 7892 57100
rect 7852 56972 7892 56981
rect 7852 56552 7892 56932
rect 7852 56503 7892 56512
rect 7756 56335 7796 56344
rect 7660 55663 7700 55672
rect 7948 55544 7988 59536
rect 8140 59527 8180 59536
rect 7564 50707 7604 50716
rect 7660 55504 7988 55544
rect 8044 59408 8084 59417
rect 8044 57644 8084 59368
rect 8044 55544 8084 57604
rect 8140 57812 8180 57821
rect 8140 56300 8180 57772
rect 8332 56804 8372 60712
rect 8332 56755 8372 56764
rect 8428 57056 8468 63736
rect 8524 63020 8564 63820
rect 8620 63524 8660 63533
rect 8620 63272 8660 63484
rect 8620 63223 8660 63232
rect 8524 62971 8564 62980
rect 8620 63104 8660 63113
rect 8524 62432 8564 62441
rect 8524 62297 8564 62392
rect 8524 60920 8564 60929
rect 8524 58736 8564 60880
rect 8620 59912 8660 63064
rect 8716 62348 8756 65668
rect 8812 65659 8852 65668
rect 8908 66844 9044 66884
rect 8812 65204 8852 65213
rect 8812 65036 8852 65164
rect 8812 64987 8852 64996
rect 8812 64700 8852 64795
rect 8812 64651 8852 64660
rect 8812 64448 8852 64457
rect 8812 63272 8852 64408
rect 8908 64028 8948 66844
rect 8908 63979 8948 63988
rect 9004 64616 9044 64625
rect 9004 63944 9044 64576
rect 9004 63860 9044 63904
rect 8908 63820 9044 63860
rect 8908 63524 8948 63820
rect 8908 63475 8948 63484
rect 9004 63692 9044 63701
rect 8812 63223 8852 63232
rect 8908 63380 8948 63389
rect 8908 62936 8948 63340
rect 9004 63104 9044 63652
rect 9004 63055 9044 63064
rect 9100 63020 9140 71884
rect 9196 70244 9236 72136
rect 9292 72092 9332 73420
rect 9388 72680 9428 72689
rect 9388 72176 9428 72640
rect 9388 72127 9428 72136
rect 9292 72043 9332 72052
rect 9484 72008 9524 73816
rect 9388 71968 9524 72008
rect 9292 71924 9332 71933
rect 9292 70748 9332 71884
rect 9292 70699 9332 70708
rect 9196 70195 9236 70204
rect 9292 69404 9332 69413
rect 9292 67724 9332 69364
rect 9292 67675 9332 67684
rect 9292 65624 9332 65633
rect 9292 65540 9332 65584
rect 9292 64952 9332 65500
rect 9292 64868 9332 64912
rect 9292 64819 9332 64828
rect 9292 64700 9332 64709
rect 9196 64112 9236 64121
rect 9196 63977 9236 64072
rect 9292 63860 9332 64660
rect 9292 63811 9332 63820
rect 9196 63776 9236 63785
rect 9196 63356 9236 63736
rect 9388 63692 9428 71968
rect 9484 71840 9524 71849
rect 9484 68648 9524 71800
rect 9484 68599 9524 68608
rect 9484 68480 9524 68489
rect 9484 67808 9524 68440
rect 9484 66884 9524 67768
rect 9484 66212 9524 66844
rect 9484 66163 9524 66172
rect 9484 65960 9524 65969
rect 9484 65456 9524 65920
rect 9484 65407 9524 65416
rect 9484 65204 9524 65213
rect 9484 64700 9524 65164
rect 9484 64651 9524 64660
rect 9196 63307 9236 63316
rect 9292 63652 9428 63692
rect 9484 63860 9524 63869
rect 9100 62980 9236 63020
rect 8908 62896 9140 62936
rect 8716 60836 8756 62308
rect 8908 62600 8948 62609
rect 8716 60787 8756 60796
rect 8812 61256 8852 61265
rect 8812 59996 8852 61216
rect 8812 59947 8852 59956
rect 8620 59324 8660 59872
rect 8620 59275 8660 59284
rect 8524 57140 8564 58696
rect 8620 59156 8660 59165
rect 8620 58652 8660 59116
rect 8620 58603 8660 58612
rect 8812 58904 8852 58913
rect 8524 57091 8564 57100
rect 8620 57812 8660 57821
rect 8332 56636 8372 56645
rect 8332 56300 8372 56596
rect 8140 56260 8276 56300
rect 7468 48103 7508 48112
rect 7564 48656 7604 48665
rect 6892 45331 6932 45340
rect 6988 46556 7028 46565
rect 6988 45632 7028 46516
rect 7180 46556 7220 46565
rect 7180 45884 7220 46516
rect 7180 45835 7220 45844
rect 7468 46556 7508 46565
rect 7564 46556 7604 48616
rect 7660 47396 7700 55504
rect 7756 54620 7796 54629
rect 7756 54116 7796 54580
rect 7948 54284 7988 54293
rect 7756 54067 7796 54076
rect 7852 54200 7892 54209
rect 7756 53948 7796 53957
rect 7756 51008 7796 53908
rect 7852 53276 7892 54160
rect 7948 54149 7988 54244
rect 7852 53227 7892 53236
rect 7948 51764 7988 51773
rect 7948 51092 7988 51724
rect 7948 51043 7988 51052
rect 7756 50672 7796 50968
rect 7756 50623 7796 50632
rect 7948 49580 7988 49589
rect 7948 48740 7988 49540
rect 7948 48691 7988 48700
rect 7660 47347 7700 47356
rect 8044 47984 8084 55504
rect 8140 56132 8180 56141
rect 8140 50420 8180 56092
rect 8236 53948 8276 56260
rect 8236 53899 8276 53908
rect 8236 53276 8276 53285
rect 8236 52016 8276 53236
rect 8236 51967 8276 51976
rect 8332 50504 8372 56260
rect 8428 53444 8468 57016
rect 8620 56132 8660 57772
rect 8428 52520 8468 53404
rect 8428 52471 8468 52480
rect 8524 54284 8564 54293
rect 8428 51680 8468 51689
rect 8428 51545 8468 51640
rect 8332 50455 8372 50464
rect 8140 50380 8276 50420
rect 7508 46516 7604 46556
rect 6700 45296 6740 45305
rect 6700 45044 6740 45256
rect 6892 45212 6932 45221
rect 6700 44995 6740 45004
rect 6796 45128 6836 45137
rect 6700 44876 6740 44885
rect 6700 44540 6740 44836
rect 6700 44120 6740 44500
rect 6700 43616 6740 44080
rect 6796 44120 6836 45088
rect 6796 44071 6836 44080
rect 6892 44960 6932 45172
rect 6988 45128 7028 45592
rect 7180 45632 7220 45641
rect 6988 45079 7028 45088
rect 7084 45296 7124 45305
rect 6796 43952 6836 43961
rect 6796 43868 6836 43912
rect 6796 43817 6836 43828
rect 6700 43567 6740 43576
rect 6796 43700 6836 43709
rect 6604 41047 6644 41056
rect 6700 43364 6740 43373
rect 6412 39871 6452 39880
rect 6508 41012 6548 41021
rect 6316 39619 6356 39628
rect 6220 39500 6260 39544
rect 6220 39420 6260 39460
rect 6412 39584 6452 39593
rect 6028 39367 6068 39376
rect 6028 39164 6068 39173
rect 5836 38275 5876 38284
rect 5932 39080 5972 39089
rect 5932 38240 5972 39040
rect 5836 38072 5876 38081
rect 5836 37937 5876 38032
rect 5932 37820 5972 38200
rect 5740 35755 5780 35764
rect 5836 37780 5972 37820
rect 5836 37652 5876 37780
rect 5836 35636 5876 37612
rect 5740 35596 5876 35636
rect 5932 37484 5972 37493
rect 5740 34544 5780 35596
rect 5740 34495 5780 34504
rect 5836 35132 5876 35141
rect 5836 34712 5876 35092
rect 5644 33991 5684 34000
rect 5740 34292 5780 34301
rect 5548 33100 5684 33140
rect 5548 33032 5588 33041
rect 5548 32948 5588 32992
rect 5548 32897 5588 32908
rect 5452 32059 5492 32068
rect 5548 32528 5588 32537
rect 5548 31940 5588 32488
rect 5356 26263 5396 26272
rect 5452 31900 5588 31940
rect 4928 25724 5296 25733
rect 4968 25684 5010 25724
rect 5050 25684 5092 25724
rect 5132 25684 5174 25724
rect 5214 25684 5256 25724
rect 4928 25675 5296 25684
rect 4972 25556 5012 25565
rect 4876 25388 4916 25397
rect 4876 25304 4916 25348
rect 4876 25253 4916 25264
rect 4972 24632 5012 25516
rect 4972 24583 5012 24592
rect 5260 25052 5300 25061
rect 5260 24632 5300 25012
rect 5452 24716 5492 31900
rect 5548 31772 5588 31781
rect 5548 30680 5588 31732
rect 5644 31436 5684 33100
rect 5740 32360 5780 34252
rect 5836 33140 5876 34672
rect 5932 34880 5972 37444
rect 5932 34376 5972 34840
rect 5932 34327 5972 34336
rect 5932 34124 5972 34133
rect 5932 33284 5972 34084
rect 5932 33235 5972 33244
rect 5836 33100 5972 33140
rect 5740 32311 5780 32320
rect 5836 32864 5876 32873
rect 5836 31940 5876 32824
rect 5836 31891 5876 31900
rect 5644 31387 5684 31396
rect 5836 31520 5876 31529
rect 5740 31184 5780 31193
rect 5548 29168 5588 30640
rect 5548 29119 5588 29128
rect 5644 31144 5740 31184
rect 5260 24583 5300 24592
rect 5356 24676 5452 24716
rect 4876 24464 4916 24559
rect 4876 24415 4916 24424
rect 4928 24212 5296 24221
rect 4968 24172 5010 24212
rect 5050 24172 5092 24212
rect 5132 24172 5174 24212
rect 5214 24172 5256 24212
rect 4928 24163 5296 24172
rect 4972 23960 5012 23969
rect 4972 23792 5012 23920
rect 4972 23743 5012 23752
rect 4780 22987 4820 22996
rect 4928 22700 5296 22709
rect 4968 22660 5010 22700
rect 5050 22660 5092 22700
rect 5132 22660 5174 22700
rect 5214 22660 5256 22700
rect 4928 22651 5296 22660
rect 5356 22532 5396 24676
rect 5452 24667 5492 24676
rect 5548 28832 5588 28841
rect 5452 23792 5492 23801
rect 5452 22700 5492 23752
rect 5548 22868 5588 28792
rect 5644 28328 5684 31144
rect 5740 31135 5780 31144
rect 5740 30848 5780 30857
rect 5740 30008 5780 30808
rect 5740 29959 5780 29968
rect 5644 28279 5684 28288
rect 5740 29840 5780 29849
rect 5644 27572 5684 27581
rect 5740 27572 5780 29800
rect 5836 28160 5876 31480
rect 5836 28111 5876 28120
rect 5740 27532 5876 27572
rect 5644 27068 5684 27532
rect 5644 27019 5684 27028
rect 5740 27404 5780 27413
rect 5548 22819 5588 22828
rect 5644 25808 5684 25817
rect 5452 22660 5588 22700
rect 5260 22492 5396 22532
rect 5452 22532 5492 22541
rect 5260 21356 5300 22492
rect 5260 21307 5300 21316
rect 5356 22364 5396 22373
rect 4928 21188 5296 21197
rect 4968 21148 5010 21188
rect 5050 21148 5092 21188
rect 5132 21148 5174 21188
rect 5214 21148 5256 21188
rect 4928 21139 5296 21148
rect 4780 21020 4820 21029
rect 4780 19424 4820 20980
rect 5356 21020 5396 22324
rect 5356 20971 5396 20980
rect 5260 20936 5300 20945
rect 5164 20852 5204 20861
rect 5164 20348 5204 20812
rect 5260 20768 5300 20896
rect 5260 20719 5300 20728
rect 5356 20852 5396 20861
rect 5164 20299 5204 20308
rect 5356 20012 5396 20812
rect 4928 19676 5296 19685
rect 4968 19636 5010 19676
rect 5050 19636 5092 19676
rect 5132 19636 5174 19676
rect 5214 19636 5256 19676
rect 4928 19627 5296 19636
rect 5356 19676 5396 19972
rect 5452 19844 5492 22492
rect 5548 22448 5588 22660
rect 5548 22399 5588 22408
rect 5548 21356 5588 21365
rect 5548 20432 5588 21316
rect 5548 20383 5588 20392
rect 5452 19795 5492 19804
rect 5548 20264 5588 20273
rect 5356 19627 5396 19636
rect 5452 19592 5492 19601
rect 4780 19375 4820 19384
rect 5164 19508 5204 19517
rect 4780 18584 4820 18593
rect 4780 18248 4820 18544
rect 5068 18584 5108 18593
rect 4972 18416 5012 18511
rect 5068 18449 5108 18544
rect 4972 18367 5012 18376
rect 5164 18416 5204 19468
rect 5260 19508 5300 19517
rect 5300 19468 5396 19508
rect 5260 19459 5300 19468
rect 5164 18367 5204 18376
rect 4780 18199 4820 18208
rect 4928 18164 5296 18173
rect 4968 18124 5010 18164
rect 5050 18124 5092 18164
rect 5132 18124 5174 18164
rect 5214 18124 5256 18164
rect 4928 18115 5296 18124
rect 4684 17956 4820 17996
rect 4492 17828 4532 17837
rect 4492 16232 4532 17788
rect 4684 17828 4724 17837
rect 4492 15224 4532 16192
rect 4492 15175 4532 15184
rect 4588 17240 4628 17249
rect 4396 13999 4436 14008
rect 4492 14552 4532 14561
rect 4492 13964 4532 14512
rect 4492 13915 4532 13924
rect 4300 13411 4340 13420
rect 4396 13880 4436 13889
rect 4300 13040 4340 13049
rect 4300 12536 4340 13000
rect 4300 12487 4340 12496
rect 4300 12284 4340 12293
rect 4300 11948 4340 12244
rect 4300 11899 4340 11908
rect 4396 11780 4436 13840
rect 4588 13880 4628 17200
rect 4684 15728 4724 17788
rect 4684 15679 4724 15688
rect 4588 13831 4628 13840
rect 4684 14804 4724 14813
rect 4012 11740 4244 11780
rect 4300 11740 4436 11780
rect 4492 13796 4532 13805
rect 3916 11572 4148 11612
rect 3688 11360 4056 11369
rect 3728 11320 3770 11360
rect 3810 11320 3852 11360
rect 3892 11320 3934 11360
rect 3974 11320 4016 11360
rect 3688 11311 4056 11320
rect 3724 11192 3764 11201
rect 3628 10352 3668 10363
rect 3628 10268 3668 10312
rect 3628 10219 3668 10228
rect 3724 10016 3764 11152
rect 3724 9967 3764 9976
rect 3688 9848 4056 9857
rect 3728 9808 3770 9848
rect 3810 9808 3852 9848
rect 3892 9808 3934 9848
rect 3974 9808 4016 9848
rect 3688 9799 4056 9808
rect 3532 9547 3572 9556
rect 4012 9512 4052 9521
rect 3436 8707 3476 8716
rect 3532 9176 3572 9185
rect 3340 6523 3380 6532
rect 3436 8000 3476 8009
rect 3340 5816 3380 5825
rect 3340 5144 3380 5776
rect 3340 5095 3380 5104
rect 3092 3508 3284 3548
rect 3052 3499 3092 3508
rect 3436 2900 3476 7960
rect 3532 6992 3572 9136
rect 3916 9008 3956 9017
rect 3820 8672 3860 8681
rect 3820 8537 3860 8632
rect 3916 8588 3956 8968
rect 4012 8924 4052 9472
rect 4108 9260 4148 11572
rect 4300 10940 4340 11740
rect 4492 11696 4532 13756
rect 4588 13712 4628 13721
rect 4588 12116 4628 13672
rect 4588 12067 4628 12076
rect 4684 12032 4724 14764
rect 4684 11983 4724 11992
rect 4492 11647 4532 11656
rect 4684 11864 4724 11873
rect 4204 10900 4340 10940
rect 4396 11612 4436 11621
rect 4204 10520 4244 10900
rect 4300 10772 4340 10781
rect 4300 10637 4340 10732
rect 4204 10480 4340 10520
rect 4108 9211 4148 9220
rect 4204 10268 4244 10277
rect 4012 8875 4052 8884
rect 3916 8539 3956 8548
rect 4108 8756 4148 8765
rect 3688 8336 4056 8345
rect 3728 8296 3770 8336
rect 3810 8296 3852 8336
rect 3892 8296 3934 8336
rect 3974 8296 4016 8336
rect 3688 8287 4056 8296
rect 3532 6943 3572 6952
rect 3688 6824 4056 6833
rect 3728 6784 3770 6824
rect 3810 6784 3852 6824
rect 3892 6784 3934 6824
rect 3974 6784 4016 6824
rect 3688 6775 4056 6784
rect 4108 6656 4148 8716
rect 4204 7412 4244 10228
rect 4300 8168 4340 10480
rect 4300 8119 4340 8128
rect 4396 8000 4436 11572
rect 4588 10436 4628 10445
rect 4492 9344 4532 9353
rect 4492 8168 4532 9304
rect 4588 8672 4628 10396
rect 4684 10268 4724 11824
rect 4684 9512 4724 10228
rect 4684 9463 4724 9472
rect 4684 9344 4724 9353
rect 4684 8840 4724 9304
rect 4684 8791 4724 8800
rect 4588 8623 4628 8632
rect 4492 8119 4532 8128
rect 4588 8168 4628 8177
rect 4204 7363 4244 7372
rect 4300 7960 4436 8000
rect 4108 6607 4148 6616
rect 4204 7244 4244 7253
rect 4204 6404 4244 7204
rect 4204 6355 4244 6364
rect 4108 5732 4148 5741
rect 3688 5312 4056 5321
rect 3728 5272 3770 5312
rect 3810 5272 3852 5312
rect 3892 5272 3934 5312
rect 3974 5272 4016 5312
rect 3688 5263 4056 5272
rect 3688 3800 4056 3809
rect 3728 3760 3770 3800
rect 3810 3760 3852 3800
rect 3892 3760 3934 3800
rect 3974 3760 4016 3800
rect 3688 3751 4056 3760
rect 3532 3464 3572 3473
rect 3532 3128 3572 3424
rect 3532 3079 3572 3088
rect 2956 2860 3092 2900
rect 2764 2624 2804 2633
rect 2476 2540 2516 2549
rect 2476 2372 2516 2500
rect 2764 2489 2804 2584
rect 2476 2323 2516 2332
rect 3052 2204 3092 2860
rect 3244 2860 3476 2900
rect 4108 2876 4148 5692
rect 4300 5732 4340 7960
rect 4588 7328 4628 8128
rect 4780 7916 4820 17956
rect 5356 17744 5396 19468
rect 5356 17695 5396 17704
rect 4876 17660 4916 17669
rect 4876 17324 4916 17620
rect 5452 17408 5492 19552
rect 5548 19424 5588 20224
rect 5548 19375 5588 19384
rect 5548 17912 5588 17921
rect 5548 17777 5588 17872
rect 4876 17275 4916 17284
rect 5356 17368 5492 17408
rect 5068 16988 5108 16999
rect 5068 16904 5108 16948
rect 5068 16855 5108 16864
rect 4928 16652 5296 16661
rect 4968 16612 5010 16652
rect 5050 16612 5092 16652
rect 5132 16612 5174 16652
rect 5214 16612 5256 16652
rect 4928 16603 5296 16612
rect 4972 16316 5012 16325
rect 4972 16181 5012 16276
rect 5260 16316 5300 16325
rect 5260 15644 5300 16276
rect 5260 15595 5300 15604
rect 4928 15140 5296 15149
rect 4968 15100 5010 15140
rect 5050 15100 5092 15140
rect 5132 15100 5174 15140
rect 5214 15100 5256 15140
rect 4928 15091 5296 15100
rect 5356 13880 5396 17368
rect 5644 17324 5684 25768
rect 5740 23288 5780 27364
rect 5836 26060 5876 27532
rect 5836 25052 5876 26020
rect 5932 26984 5972 33100
rect 6028 29504 6068 39124
rect 6220 39164 6260 39173
rect 6220 39080 6260 39124
rect 6220 39029 6260 39040
rect 6124 38996 6164 39005
rect 6124 38324 6164 38956
rect 6124 38275 6164 38284
rect 6220 38240 6260 38249
rect 6124 38072 6164 38081
rect 6124 37820 6164 38032
rect 6124 37771 6164 37780
rect 6124 37484 6164 37493
rect 6124 36644 6164 37444
rect 6124 36595 6164 36604
rect 6124 36476 6164 36485
rect 6220 36476 6260 38200
rect 6316 38072 6356 38083
rect 6316 37988 6356 38032
rect 6316 37939 6356 37948
rect 6412 37820 6452 39544
rect 6508 39164 6548 40972
rect 6604 40928 6644 40937
rect 6604 39752 6644 40888
rect 6604 39703 6644 39712
rect 6700 39584 6740 43324
rect 6796 41852 6836 43660
rect 6892 42776 6932 44920
rect 7084 43700 7124 45256
rect 7180 44876 7220 45592
rect 7468 45464 7508 46516
rect 7852 45968 7892 45977
rect 7468 45415 7508 45424
rect 7660 45464 7700 45473
rect 7564 45380 7604 45389
rect 7564 45245 7604 45340
rect 7660 45128 7700 45424
rect 7660 45079 7700 45088
rect 7468 45044 7508 45053
rect 7180 44827 7220 44836
rect 7276 44960 7316 44969
rect 7276 44456 7316 44920
rect 7276 44407 7316 44416
rect 7084 43651 7124 43660
rect 7180 44036 7220 44045
rect 6892 42727 6932 42736
rect 6988 43532 7028 43541
rect 6796 41803 6836 41812
rect 6892 42608 6932 42617
rect 6892 42440 6932 42568
rect 6508 39115 6548 39124
rect 6604 39544 6740 39584
rect 6796 41180 6836 41189
rect 6796 40760 6836 41140
rect 6796 39836 6836 40720
rect 6604 39080 6644 39544
rect 6604 39031 6644 39040
rect 6700 39416 6740 39425
rect 6700 38912 6740 39376
rect 6796 39080 6836 39796
rect 6796 39031 6836 39040
rect 6892 40256 6932 42400
rect 6892 39080 6932 40216
rect 6988 42524 7028 43492
rect 6988 39500 7028 42484
rect 7084 43448 7124 43457
rect 7180 43448 7220 43996
rect 7468 44036 7508 45004
rect 7852 45044 7892 45928
rect 7468 43987 7508 43996
rect 7564 44204 7604 44213
rect 7124 43408 7220 43448
rect 7084 40844 7124 43408
rect 7180 42776 7220 42785
rect 7180 42020 7220 42736
rect 7372 42272 7412 42281
rect 7180 41980 7316 42020
rect 7180 41852 7220 41861
rect 7180 41600 7220 41812
rect 7180 41180 7220 41560
rect 7180 41012 7220 41140
rect 7180 40963 7220 40972
rect 7084 40795 7124 40804
rect 7180 40676 7220 40685
rect 6988 39365 7028 39460
rect 7084 40592 7124 40601
rect 7084 39752 7124 40552
rect 7180 40592 7220 40636
rect 7180 40541 7220 40552
rect 7084 39668 7124 39712
rect 6988 39248 7028 39257
rect 6988 39113 7028 39208
rect 6892 39031 6932 39040
rect 6988 38996 7028 39005
rect 6604 38872 6700 38912
rect 6508 38324 6548 38333
rect 6508 38072 6548 38284
rect 6508 38023 6548 38032
rect 6164 36436 6260 36476
rect 6124 36427 6164 36436
rect 6124 35888 6164 35897
rect 6124 34964 6164 35848
rect 6124 32192 6164 34924
rect 6220 33956 6260 36436
rect 6316 37232 6356 37241
rect 6316 35972 6356 37192
rect 6316 35923 6356 35932
rect 6220 33907 6260 33916
rect 6316 34880 6356 34889
rect 6220 33788 6260 33797
rect 6220 32528 6260 33748
rect 6316 32948 6356 34840
rect 6412 33872 6452 37780
rect 6412 33823 6452 33832
rect 6508 37904 6548 37913
rect 6316 32899 6356 32908
rect 6220 32479 6260 32488
rect 6412 32192 6452 32201
rect 6124 32152 6412 32192
rect 6028 29455 6068 29464
rect 6124 31940 6164 31949
rect 6124 31352 6164 31900
rect 6220 31352 6260 31361
rect 6124 31312 6220 31352
rect 6124 31268 6164 31312
rect 6220 31303 6260 31312
rect 6124 29420 6164 31228
rect 6220 30764 6260 30773
rect 6220 29924 6260 30724
rect 6316 30092 6356 32152
rect 6412 32143 6452 32152
rect 6316 30043 6356 30052
rect 6412 31604 6452 31613
rect 6220 29875 6260 29884
rect 6412 29588 6452 31564
rect 6412 29539 6452 29548
rect 6124 29371 6164 29380
rect 6316 29504 6356 29513
rect 6028 29336 6068 29345
rect 6028 27908 6068 29296
rect 6028 27859 6068 27868
rect 6124 28916 6164 28925
rect 5932 25220 5972 26944
rect 6028 27404 6068 27413
rect 6028 26312 6068 27364
rect 6124 26396 6164 28876
rect 6124 26347 6164 26356
rect 6220 28244 6260 28253
rect 6028 26263 6068 26272
rect 5932 25171 5972 25180
rect 6028 26144 6068 26153
rect 6028 25808 6068 26104
rect 5836 23876 5876 25012
rect 5932 25052 5972 25061
rect 5932 24800 5972 25012
rect 5932 24751 5972 24760
rect 5836 23827 5876 23836
rect 5932 24632 5972 24641
rect 5932 23792 5972 24592
rect 5932 23743 5972 23752
rect 5740 23239 5780 23248
rect 5932 23204 5972 23213
rect 5740 23120 5780 23129
rect 5740 18584 5780 23080
rect 5740 18535 5780 18544
rect 5836 22616 5876 22625
rect 5836 18416 5876 22576
rect 5932 22196 5972 23164
rect 6028 23060 6068 25768
rect 6124 24800 6164 24809
rect 6124 23204 6164 24760
rect 6124 23155 6164 23164
rect 6028 23036 6164 23060
rect 6068 23020 6164 23036
rect 6028 22987 6068 22996
rect 5932 20096 5972 22156
rect 6028 22280 6068 22289
rect 6028 21608 6068 22240
rect 6028 20264 6068 21568
rect 6124 20852 6164 23020
rect 6124 20803 6164 20812
rect 6028 20215 6068 20224
rect 6124 20684 6164 20693
rect 5932 20056 6068 20096
rect 5932 19760 5972 19855
rect 5932 19711 5972 19720
rect 5740 18376 5876 18416
rect 5932 19592 5972 19601
rect 5740 17744 5780 18376
rect 5740 17695 5780 17704
rect 5836 17996 5876 18005
rect 5356 13831 5396 13840
rect 5452 17284 5684 17324
rect 5740 17408 5780 17417
rect 4928 13628 5296 13637
rect 4968 13588 5010 13628
rect 5050 13588 5092 13628
rect 5132 13588 5174 13628
rect 5214 13588 5256 13628
rect 4928 13579 5296 13588
rect 5356 13544 5396 13553
rect 5164 13460 5204 13469
rect 4876 12704 4916 12713
rect 4876 12536 4916 12664
rect 4876 12487 4916 12496
rect 5164 12536 5204 13420
rect 5260 13208 5300 13217
rect 5260 12704 5300 13168
rect 5260 12655 5300 12664
rect 5164 12284 5204 12496
rect 5164 12235 5204 12244
rect 4928 12116 5296 12125
rect 4968 12076 5010 12116
rect 5050 12076 5092 12116
rect 5132 12076 5174 12116
rect 5214 12076 5256 12116
rect 4928 12067 5296 12076
rect 5260 11948 5300 11957
rect 4972 11864 5012 11873
rect 4972 11612 5012 11824
rect 4972 11563 5012 11572
rect 5260 10772 5300 11908
rect 5356 10940 5396 13504
rect 5356 10891 5396 10900
rect 5260 10732 5396 10772
rect 4928 10604 5296 10613
rect 4968 10564 5010 10604
rect 5050 10564 5092 10604
rect 5132 10564 5174 10604
rect 5214 10564 5256 10604
rect 4928 10555 5296 10564
rect 5164 10436 5204 10445
rect 5164 9428 5204 10396
rect 5164 9379 5204 9388
rect 4928 9092 5296 9101
rect 4968 9052 5010 9092
rect 5050 9052 5092 9092
rect 5132 9052 5174 9092
rect 5214 9052 5256 9092
rect 4928 9043 5296 9052
rect 5356 9008 5396 10732
rect 5356 8959 5396 8968
rect 5068 8924 5108 8933
rect 5068 8789 5108 8884
rect 5356 8840 5396 8849
rect 4492 7288 4628 7328
rect 4684 7876 4820 7916
rect 4396 7160 4436 7169
rect 4396 6824 4436 7120
rect 4396 6775 4436 6784
rect 4300 5683 4340 5692
rect 4492 4724 4532 7288
rect 4588 7160 4628 7169
rect 4588 5900 4628 7120
rect 4588 5851 4628 5860
rect 4492 4675 4532 4684
rect 4684 4556 4724 7876
rect 4928 7580 5296 7589
rect 4968 7540 5010 7580
rect 5050 7540 5092 7580
rect 5132 7540 5174 7580
rect 5214 7540 5256 7580
rect 4928 7531 5296 7540
rect 5356 7160 5396 8800
rect 5452 7916 5492 17284
rect 5740 16232 5780 17368
rect 5548 16192 5780 16232
rect 5836 16232 5876 17956
rect 5548 13712 5588 16192
rect 5836 16183 5876 16192
rect 5548 13663 5588 13672
rect 5644 16064 5684 16073
rect 5548 13544 5588 13553
rect 5548 13292 5588 13504
rect 5548 13243 5588 13252
rect 5548 13040 5588 13049
rect 5548 12536 5588 13000
rect 5548 12487 5588 12496
rect 5548 12284 5588 12293
rect 5548 9680 5588 12244
rect 5644 11948 5684 16024
rect 5836 15896 5876 15905
rect 5740 15476 5780 15485
rect 5740 14888 5780 15436
rect 5740 14839 5780 14848
rect 5836 14720 5876 15856
rect 5644 11899 5684 11908
rect 5740 14680 5876 14720
rect 5740 11780 5780 14680
rect 5836 14048 5876 14057
rect 5932 14048 5972 19552
rect 6028 17828 6068 20056
rect 6124 19424 6164 20644
rect 6220 19676 6260 28204
rect 6316 24632 6356 29464
rect 6412 29420 6452 29429
rect 6412 28580 6452 29380
rect 6508 29336 6548 37864
rect 6604 35384 6644 38872
rect 6700 38863 6740 38872
rect 6892 38912 6932 38921
rect 6700 38492 6740 38501
rect 6700 37484 6740 38452
rect 6796 38072 6836 38081
rect 6796 37988 6836 38032
rect 6796 37937 6836 37948
rect 6892 38072 6932 38872
rect 6988 38408 7028 38956
rect 6988 38359 7028 38368
rect 6892 37820 6932 38032
rect 6892 37771 6932 37780
rect 6988 38156 7028 38165
rect 6700 37435 6740 37444
rect 6988 37148 7028 38116
rect 7084 38072 7124 39628
rect 7276 39164 7316 41980
rect 7372 40676 7412 42232
rect 7372 40627 7412 40636
rect 7468 41180 7508 41189
rect 7468 40928 7508 41140
rect 7372 40508 7412 40517
rect 7372 40424 7412 40468
rect 7372 40373 7412 40384
rect 7276 39124 7412 39164
rect 7276 38996 7316 39005
rect 7084 37988 7124 38032
rect 7084 37908 7124 37948
rect 7180 38912 7220 38921
rect 6988 37108 7124 37148
rect 6796 36812 6836 36821
rect 6700 36644 6740 36653
rect 6700 36140 6740 36604
rect 6700 36091 6740 36100
rect 6604 35335 6644 35344
rect 6796 35888 6836 36772
rect 6796 35468 6836 35848
rect 6700 34796 6740 34805
rect 6508 29287 6548 29296
rect 6604 34040 6644 34049
rect 6412 28531 6452 28540
rect 6604 28244 6644 34000
rect 6604 28195 6644 28204
rect 6700 28076 6740 34756
rect 6796 33620 6836 35428
rect 6796 33571 6836 33580
rect 6988 36392 7028 36401
rect 6796 32948 6836 32957
rect 6796 32360 6836 32908
rect 6796 32311 6836 32320
rect 6892 32864 6932 32873
rect 6892 32108 6932 32824
rect 6988 32276 7028 36352
rect 7084 34964 7124 37108
rect 7180 35132 7220 38872
rect 7276 38156 7316 38956
rect 7276 38107 7316 38116
rect 7372 38240 7412 39124
rect 7372 38156 7412 38200
rect 7372 38107 7412 38116
rect 7372 37988 7412 37997
rect 7276 37316 7316 37325
rect 7276 37181 7316 37276
rect 7276 36392 7316 36401
rect 7276 36056 7316 36352
rect 7276 36007 7316 36016
rect 7180 35083 7220 35092
rect 7276 35552 7316 35561
rect 7084 34924 7220 34964
rect 7084 32696 7124 32705
rect 7084 32444 7124 32656
rect 7084 32395 7124 32404
rect 7084 32276 7124 32285
rect 6988 32236 7084 32276
rect 7084 32227 7124 32236
rect 6796 32068 6932 32108
rect 7084 32108 7124 32117
rect 6796 31436 6836 32068
rect 6988 31940 7028 31949
rect 6892 31856 6932 31865
rect 6892 31721 6932 31816
rect 6796 31387 6836 31396
rect 6892 31520 6932 31529
rect 6796 31100 6836 31109
rect 6796 30965 6836 31060
rect 6892 30680 6932 31480
rect 6892 29924 6932 30640
rect 6892 29084 6932 29884
rect 6892 29035 6932 29044
rect 6796 29000 6836 29009
rect 6796 28580 6836 28960
rect 6796 28531 6836 28540
rect 6316 24583 6356 24592
rect 6412 28036 6740 28076
rect 6796 28412 6836 28421
rect 6316 24464 6356 24473
rect 6316 20180 6356 24424
rect 6412 22532 6452 28036
rect 6508 27320 6548 27329
rect 6508 26984 6548 27280
rect 6508 26935 6548 26944
rect 6604 27236 6644 27245
rect 6508 25136 6548 25145
rect 6508 24884 6548 25096
rect 6508 24835 6548 24844
rect 6412 22483 6452 22492
rect 6412 22364 6452 22373
rect 6412 21776 6452 22324
rect 6412 21727 6452 21736
rect 6412 21524 6452 21533
rect 6412 21188 6452 21484
rect 6412 21020 6452 21148
rect 6412 20971 6452 20980
rect 6508 21440 6548 21449
rect 6316 20140 6452 20180
rect 6220 19627 6260 19636
rect 6316 20012 6356 20021
rect 6124 19384 6260 19424
rect 6124 19256 6164 19265
rect 6124 19121 6164 19216
rect 6220 19172 6260 19384
rect 6028 17779 6068 17788
rect 6124 18836 6164 18845
rect 6124 16988 6164 18796
rect 6220 17744 6260 19132
rect 6220 17695 6260 17704
rect 6316 19088 6356 19972
rect 6124 16939 6164 16948
rect 6220 17324 6260 17333
rect 6028 16568 6068 16577
rect 6028 16232 6068 16528
rect 6124 16484 6164 16493
rect 6124 16349 6164 16444
rect 6028 16183 6068 16192
rect 5876 14008 5972 14048
rect 6028 16064 6068 16073
rect 5836 13999 5876 14008
rect 5836 13880 5876 13920
rect 5836 13796 5876 13840
rect 5836 12704 5876 13756
rect 5932 13880 5972 13889
rect 5932 13628 5972 13840
rect 5932 13579 5972 13588
rect 5932 13376 5972 13385
rect 5932 12872 5972 13336
rect 5932 12823 5972 12832
rect 5836 12664 5972 12704
rect 5548 9631 5588 9640
rect 5644 11740 5740 11780
rect 5644 8000 5684 11740
rect 5740 11731 5780 11740
rect 5836 12536 5876 12545
rect 5836 10436 5876 12496
rect 5932 12284 5972 12664
rect 5932 12235 5972 12244
rect 5836 10387 5876 10396
rect 5932 10268 5972 10277
rect 5836 9680 5876 9689
rect 5836 9545 5876 9640
rect 5836 8756 5876 8765
rect 5836 8168 5876 8716
rect 5836 8119 5876 8128
rect 5644 7960 5780 8000
rect 5452 7876 5684 7916
rect 5356 7111 5396 7120
rect 4928 6068 5296 6077
rect 4968 6028 5010 6068
rect 5050 6028 5092 6068
rect 5132 6028 5174 6068
rect 5214 6028 5256 6068
rect 4928 6019 5296 6028
rect 4876 5648 4916 5657
rect 4876 5513 4916 5608
rect 4780 5480 4820 5489
rect 4780 5345 4820 5440
rect 3052 2155 3092 2164
rect 3148 2624 3188 2633
rect 2284 2120 2324 2129
rect 2284 1985 2324 2080
rect 2572 2120 2612 2129
rect 2380 2036 2420 2045
rect 2380 80 2420 1996
rect 2572 1985 2612 2080
rect 2764 1868 2804 1877
rect 2476 1784 2516 1793
rect 2476 1700 2516 1744
rect 2476 1649 2516 1660
rect 2572 1784 2612 1793
rect 2572 80 2612 1744
rect 2764 80 2804 1828
rect 2956 1868 2996 1877
rect 2956 80 2996 1828
rect 3148 80 3188 2584
rect 3244 1784 3284 2860
rect 4108 2827 4148 2836
rect 4396 4516 4724 4556
rect 4928 4556 5296 4565
rect 4968 4516 5010 4556
rect 5050 4516 5092 4556
rect 5132 4516 5174 4556
rect 5214 4516 5256 4556
rect 3532 2792 3572 2801
rect 3532 2657 3572 2752
rect 3628 2624 3668 2633
rect 3628 2456 3668 2584
rect 3532 2416 3668 2456
rect 4108 2624 4148 2633
rect 3340 2120 3380 2215
rect 3340 2071 3380 2080
rect 3244 1735 3284 1744
rect 3340 1868 3380 1877
rect 3340 80 3380 1828
rect 3532 80 3572 2416
rect 3688 2288 4056 2297
rect 3728 2248 3770 2288
rect 3810 2248 3852 2288
rect 3892 2248 3934 2288
rect 3974 2248 4016 2288
rect 3688 2239 4056 2248
rect 3724 2036 3764 2045
rect 3724 80 3764 1996
rect 4108 1364 4148 2584
rect 4300 2624 4340 2633
rect 4204 2204 4244 2213
rect 4204 2120 4244 2164
rect 4204 2069 4244 2080
rect 3916 1324 4148 1364
rect 4204 1868 4244 1877
rect 3916 80 3956 1324
rect 4204 1028 4244 1828
rect 4108 988 4244 1028
rect 4108 80 4148 988
rect 4300 80 4340 2584
rect 4396 1616 4436 4516
rect 4928 4507 5296 4516
rect 5356 4304 5396 4313
rect 4684 3800 4724 3809
rect 4684 2876 4724 3760
rect 4928 3044 5296 3053
rect 4968 3004 5010 3044
rect 5050 3004 5092 3044
rect 5132 3004 5174 3044
rect 5214 3004 5256 3044
rect 4928 2995 5296 3004
rect 5356 2900 5396 4264
rect 4684 2827 4724 2836
rect 4876 2876 4916 2885
rect 4876 2792 4916 2836
rect 4876 2741 4916 2752
rect 5260 2860 5396 2900
rect 5548 3548 5588 3557
rect 4684 2624 4724 2633
rect 4396 1567 4436 1576
rect 4492 1868 4532 1877
rect 4492 80 4532 1828
rect 4684 80 4724 2584
rect 5260 2456 5300 2860
rect 5260 2407 5300 2416
rect 5356 2624 5396 2633
rect 4780 1868 4820 1877
rect 4780 860 4820 1828
rect 4928 1532 5296 1541
rect 4968 1492 5010 1532
rect 5050 1492 5092 1532
rect 5132 1492 5174 1532
rect 5214 1492 5256 1532
rect 4928 1483 5296 1492
rect 5356 1364 5396 2584
rect 5068 1324 5396 1364
rect 5452 2540 5492 2549
rect 4780 820 4916 860
rect 4876 80 4916 820
rect 5068 80 5108 1324
rect 5260 1028 5300 1037
rect 5260 80 5300 988
rect 5452 80 5492 2500
rect 5548 2120 5588 3508
rect 5644 2456 5684 7876
rect 5740 7244 5780 7960
rect 5740 6404 5780 7204
rect 5740 6355 5780 6364
rect 5932 6236 5972 10228
rect 6028 6824 6068 16024
rect 6124 15812 6164 15821
rect 6124 13796 6164 15772
rect 6220 15140 6260 17284
rect 6220 15091 6260 15100
rect 6220 14300 6260 14309
rect 6220 14048 6260 14260
rect 6220 13913 6260 14008
rect 6124 13756 6260 13796
rect 6124 13628 6164 13637
rect 6124 12452 6164 13588
rect 6124 12403 6164 12412
rect 6124 12284 6164 12293
rect 6124 10856 6164 12244
rect 6124 8840 6164 10816
rect 6220 10268 6260 13756
rect 6220 10219 6260 10228
rect 6316 13208 6356 19048
rect 6316 11780 6356 13168
rect 6412 12200 6452 20140
rect 6508 18836 6548 21400
rect 6508 18787 6548 18796
rect 6508 18584 6548 18679
rect 6508 18535 6548 18544
rect 6508 18416 6548 18425
rect 6508 17912 6548 18376
rect 6508 17863 6548 17872
rect 6508 17744 6548 17753
rect 6508 17324 6548 17704
rect 6508 17275 6548 17284
rect 6508 16988 6548 16997
rect 6508 16652 6548 16948
rect 6604 16820 6644 27196
rect 6796 26816 6836 28372
rect 6892 27992 6932 28001
rect 6892 27572 6932 27952
rect 6892 27523 6932 27532
rect 6988 26900 7028 31900
rect 6988 26851 7028 26860
rect 6796 26767 6836 26776
rect 6796 26648 6836 26657
rect 6700 26564 6740 26573
rect 6700 25388 6740 26524
rect 6796 26228 6836 26608
rect 6796 26179 6836 26188
rect 6700 25339 6740 25348
rect 6796 25640 6836 25649
rect 6604 16771 6644 16780
rect 6700 25220 6740 25229
rect 6508 16612 6644 16652
rect 6508 16484 6548 16493
rect 6508 15560 6548 16444
rect 6604 16400 6644 16612
rect 6604 16351 6644 16360
rect 6604 16232 6644 16241
rect 6604 15980 6644 16192
rect 6604 15931 6644 15940
rect 6508 15511 6548 15520
rect 6604 15644 6644 15653
rect 6604 15509 6644 15604
rect 6700 15392 6740 25180
rect 6796 23960 6836 25600
rect 7084 25640 7124 32068
rect 7084 25591 7124 25600
rect 7180 25472 7220 34924
rect 7276 34460 7316 35512
rect 7276 33620 7316 34420
rect 7276 33571 7316 33580
rect 7372 33140 7412 37948
rect 7468 36308 7508 40888
rect 7468 36259 7508 36268
rect 7372 33091 7412 33100
rect 7468 35132 7508 35141
rect 7468 34208 7508 35092
rect 7372 33032 7412 33041
rect 7276 32696 7316 32705
rect 7276 32108 7316 32656
rect 7372 32528 7412 32992
rect 7468 32948 7508 34168
rect 7468 32899 7508 32908
rect 7564 34460 7604 44164
rect 7660 43532 7700 43541
rect 7660 40928 7700 43492
rect 7756 43532 7796 43541
rect 7756 42608 7796 43492
rect 7756 41684 7796 42568
rect 7852 41852 7892 45004
rect 7948 45296 7988 45305
rect 7948 45128 7988 45256
rect 7948 44120 7988 45088
rect 7948 43532 7988 44080
rect 7948 42692 7988 43492
rect 8044 43220 8084 47944
rect 8140 50252 8180 50261
rect 8140 47816 8180 50212
rect 8236 48488 8276 50380
rect 8524 50252 8564 54244
rect 8524 50203 8564 50212
rect 8620 48908 8660 56092
rect 8812 55544 8852 58864
rect 8908 57308 8948 62560
rect 9004 59324 9044 59333
rect 9004 58568 9044 59284
rect 9004 57896 9044 58528
rect 9004 57847 9044 57856
rect 8908 57259 8948 57268
rect 9004 55796 9044 55805
rect 8812 54536 8852 55504
rect 8812 54487 8852 54496
rect 8908 55712 8948 55721
rect 8908 54032 8948 55672
rect 9004 55628 9044 55756
rect 9004 55579 9044 55588
rect 9004 54872 9044 54881
rect 9004 54788 9044 54832
rect 9004 54284 9044 54748
rect 9004 54235 9044 54244
rect 8812 53948 8852 53957
rect 8716 52016 8756 52025
rect 8716 50840 8756 51976
rect 8716 50791 8756 50800
rect 8620 48859 8660 48868
rect 8812 48740 8852 53908
rect 8908 50504 8948 53992
rect 9100 51680 9140 62896
rect 9196 57812 9236 62980
rect 9292 61760 9332 63652
rect 9388 63524 9428 63533
rect 9388 63188 9428 63484
rect 9388 63139 9428 63148
rect 9388 63020 9428 63029
rect 9388 62600 9428 62980
rect 9388 62551 9428 62560
rect 9484 62348 9524 63820
rect 9484 62299 9524 62308
rect 9484 62012 9524 62021
rect 9292 61720 9428 61760
rect 9292 59576 9332 59585
rect 9292 58904 9332 59536
rect 9292 58652 9332 58864
rect 9292 58603 9332 58612
rect 9196 57763 9236 57772
rect 9292 57644 9332 57653
rect 9292 57140 9332 57604
rect 9292 57091 9332 57100
rect 9292 56300 9332 56309
rect 9292 55880 9332 56260
rect 9292 54872 9332 55840
rect 9292 54823 9332 54832
rect 9100 51631 9140 51640
rect 9196 54788 9236 54797
rect 8908 50464 9140 50504
rect 9004 50336 9044 50345
rect 8812 48691 8852 48700
rect 8908 48824 8948 48833
rect 8236 48439 8276 48448
rect 8908 47900 8948 48784
rect 8140 46640 8180 47776
rect 8812 47816 8852 47825
rect 8620 47228 8660 47237
rect 8620 47093 8660 47188
rect 8140 46591 8180 46600
rect 8524 46976 8564 46985
rect 8236 46052 8276 46061
rect 8140 45884 8180 45893
rect 8140 45044 8180 45844
rect 8140 44995 8180 45004
rect 8236 45716 8276 46012
rect 8236 44204 8276 45676
rect 8428 45800 8468 45809
rect 8236 44155 8276 44164
rect 8332 45632 8372 45641
rect 8332 44036 8372 45592
rect 8236 43700 8276 43709
rect 8044 43180 8180 43220
rect 7948 42188 7988 42652
rect 7948 42139 7988 42148
rect 7852 41803 7892 41812
rect 7948 41936 7988 41945
rect 7852 41684 7892 41693
rect 7756 41644 7852 41684
rect 7756 41096 7796 41644
rect 7852 41635 7892 41644
rect 7756 41047 7796 41056
rect 7660 40888 7892 40928
rect 7756 40592 7796 40601
rect 7660 40484 7700 40493
rect 7660 40004 7700 40444
rect 7660 39955 7700 39964
rect 7756 38240 7796 40552
rect 7852 39668 7892 40888
rect 7852 39619 7892 39628
rect 7756 38191 7796 38200
rect 7660 37484 7700 37493
rect 7660 36476 7700 37444
rect 7660 36427 7700 36436
rect 7756 37400 7796 37409
rect 7756 36644 7796 37360
rect 7948 36896 7988 41896
rect 8044 41600 8084 41609
rect 8044 41264 8084 41560
rect 8044 41215 8084 41224
rect 8044 40424 8084 40433
rect 8044 40088 8084 40384
rect 8044 40039 8084 40048
rect 7948 36847 7988 36856
rect 8044 37568 8084 37577
rect 7468 32696 7508 32791
rect 7468 32647 7508 32656
rect 7372 32488 7508 32528
rect 7276 32059 7316 32068
rect 7372 32360 7412 32369
rect 7372 31856 7412 32320
rect 7372 31807 7412 31816
rect 7276 31436 7316 31445
rect 7276 30764 7316 31396
rect 7276 30715 7316 30724
rect 7468 30596 7508 32488
rect 7564 32192 7604 34420
rect 7660 36308 7700 36317
rect 7660 32360 7700 36268
rect 7756 36056 7796 36604
rect 7756 36007 7796 36016
rect 8044 35804 8084 37528
rect 8044 35755 8084 35764
rect 7756 35216 7796 35225
rect 7756 33872 7796 35176
rect 8044 35132 8084 35141
rect 7948 35048 7988 35057
rect 7756 33032 7796 33832
rect 7756 32983 7796 32992
rect 7852 34964 7892 34973
rect 7660 32311 7700 32320
rect 7756 32864 7796 32873
rect 7564 32143 7604 32152
rect 7660 31940 7700 31949
rect 7372 30512 7412 30521
rect 7276 30428 7316 30437
rect 7276 30260 7316 30388
rect 7276 30211 7316 30220
rect 7372 29756 7412 30472
rect 7372 29091 7412 29716
rect 7276 29000 7316 29009
rect 7276 28412 7316 28960
rect 7372 29000 7416 29091
rect 7468 29084 7508 30556
rect 7468 29035 7508 29044
rect 7564 30680 7604 30689
rect 7564 29924 7604 30640
rect 7564 29168 7604 29884
rect 7372 28951 7416 28960
rect 7564 28412 7604 29128
rect 7316 28372 7412 28412
rect 7276 28363 7316 28372
rect 7276 28244 7316 28253
rect 7276 26648 7316 28204
rect 7276 26599 7316 26608
rect 7276 26480 7316 26489
rect 7276 26312 7316 26440
rect 7276 26263 7316 26272
rect 7276 26060 7316 26069
rect 7276 25556 7316 26020
rect 7276 25507 7316 25516
rect 7084 25432 7220 25472
rect 6988 24968 7028 24977
rect 6988 24833 7028 24928
rect 6988 24632 7028 24641
rect 6796 23911 6836 23920
rect 6892 24548 6932 24557
rect 6796 23456 6836 23465
rect 6796 21860 6836 23416
rect 6796 21811 6836 21820
rect 6796 21692 6836 21701
rect 6796 19088 6836 21652
rect 6892 21356 6932 24508
rect 6988 24497 7028 24592
rect 7084 24548 7124 25432
rect 7276 25388 7316 25397
rect 7084 24499 7124 24508
rect 7180 25304 7220 25313
rect 7180 24044 7220 25264
rect 7180 23995 7220 24004
rect 6988 23876 7028 23885
rect 7276 23876 7316 25348
rect 6988 21692 7028 23836
rect 7180 23836 7276 23876
rect 6988 21643 7028 21652
rect 7084 23624 7124 23633
rect 7084 22616 7124 23584
rect 6892 21307 6932 21316
rect 6988 21524 7028 21533
rect 6892 20684 6932 20693
rect 6892 20264 6932 20644
rect 6892 20215 6932 20224
rect 6796 19048 6932 19088
rect 6412 12151 6452 12160
rect 6508 15352 6740 15392
rect 6796 18920 6836 18929
rect 6508 12032 6548 15352
rect 6700 15224 6740 15233
rect 6604 15140 6644 15149
rect 6604 13796 6644 15100
rect 6604 13747 6644 13756
rect 6604 12620 6644 12631
rect 6604 12536 6644 12580
rect 6604 12487 6644 12496
rect 6316 10184 6356 11740
rect 6412 11992 6548 12032
rect 6604 12368 6644 12377
rect 6412 11192 6452 11992
rect 6604 11948 6644 12328
rect 6604 11899 6644 11908
rect 6412 11143 6452 11152
rect 6508 11780 6548 11789
rect 6220 10016 6260 10025
rect 6220 9428 6260 9976
rect 6220 9379 6260 9388
rect 6124 8791 6164 8800
rect 6220 9176 6260 9185
rect 6220 8672 6260 9136
rect 6220 8623 6260 8632
rect 6316 8084 6356 10144
rect 6412 11024 6452 11033
rect 6412 10352 6452 10984
rect 6412 8588 6452 10312
rect 6508 10268 6548 11740
rect 6508 10219 6548 10228
rect 6604 11192 6644 11201
rect 6604 9428 6644 11152
rect 6700 10940 6740 15184
rect 6796 11024 6836 18880
rect 6892 13460 6932 19048
rect 6988 18500 7028 21484
rect 7084 20180 7124 22576
rect 7180 21608 7220 23836
rect 7276 23827 7316 23836
rect 7372 23708 7412 28372
rect 7468 28328 7508 28337
rect 7468 27068 7508 28288
rect 7468 27019 7508 27028
rect 7468 26900 7508 26909
rect 7468 26144 7508 26860
rect 7468 26095 7508 26104
rect 7468 25976 7508 25985
rect 7468 25841 7508 25936
rect 7468 24968 7508 24977
rect 7468 24800 7508 24928
rect 7468 24751 7508 24760
rect 7468 24548 7508 24557
rect 7468 24413 7508 24508
rect 7564 24380 7604 28372
rect 7660 25220 7700 31900
rect 7756 30176 7796 32824
rect 7756 30127 7796 30136
rect 7756 30008 7796 30017
rect 7852 30008 7892 34924
rect 7948 33116 7988 35008
rect 7948 33067 7988 33076
rect 7948 32948 7988 32957
rect 7948 32696 7988 32908
rect 8044 32780 8084 35092
rect 8044 32731 8084 32740
rect 7948 32647 7988 32656
rect 7948 32528 7988 32537
rect 7948 31856 7988 32488
rect 8044 32444 8084 32453
rect 8044 32309 8084 32404
rect 8140 32024 8180 43180
rect 8236 42776 8276 43660
rect 8236 42727 8276 42736
rect 8332 42692 8372 43996
rect 8428 45044 8468 45760
rect 8428 43616 8468 45004
rect 8428 43567 8468 43576
rect 8332 42643 8372 42652
rect 8428 42020 8468 42029
rect 8428 39920 8468 41980
rect 8236 39668 8276 39677
rect 8236 38912 8276 39628
rect 8236 38863 8276 38872
rect 8332 39080 8372 39089
rect 8236 37232 8276 37241
rect 8236 36728 8276 37192
rect 8236 36679 8276 36688
rect 8236 35972 8276 35981
rect 8236 35837 8276 35932
rect 8236 35048 8276 35057
rect 8236 33200 8276 35008
rect 8236 33151 8276 33160
rect 8332 32864 8372 39040
rect 8428 38996 8468 39880
rect 8524 39332 8564 46936
rect 8620 45632 8660 45641
rect 8620 45128 8660 45592
rect 8620 45079 8660 45088
rect 8716 44624 8756 44633
rect 8716 44456 8756 44584
rect 8716 44407 8756 44416
rect 8716 43616 8756 43625
rect 8716 42020 8756 43576
rect 8716 41180 8756 41980
rect 8716 41131 8756 41140
rect 8716 40760 8756 40769
rect 8620 40424 8660 40433
rect 8620 40088 8660 40384
rect 8620 40039 8660 40048
rect 8524 39283 8564 39292
rect 8428 38947 8468 38956
rect 8620 39248 8660 39257
rect 8428 38828 8468 38837
rect 8428 38240 8468 38788
rect 8620 38324 8660 39208
rect 8620 38275 8660 38284
rect 8428 38191 8468 38200
rect 8620 37988 8660 37997
rect 8620 37400 8660 37948
rect 8620 37351 8660 37360
rect 8428 36476 8468 36485
rect 8428 34628 8468 36436
rect 8428 34579 8468 34588
rect 8524 36056 8564 36065
rect 8428 33956 8468 33965
rect 8428 33200 8468 33916
rect 8428 33151 8468 33160
rect 7948 31807 7988 31816
rect 8044 31984 8180 32024
rect 8236 32824 8372 32864
rect 8428 32948 8468 32957
rect 7948 31352 7988 31361
rect 7948 30092 7988 31312
rect 7948 30043 7988 30052
rect 7796 29968 7892 30008
rect 7756 28328 7796 29968
rect 7948 29924 7988 29933
rect 7756 28279 7796 28288
rect 7852 28412 7892 28421
rect 7852 27572 7892 28372
rect 7948 28412 7988 29884
rect 7948 28363 7988 28372
rect 7852 27523 7892 27532
rect 7756 27488 7796 27497
rect 7756 26900 7796 27448
rect 7948 27488 7988 27497
rect 7948 27068 7988 27448
rect 7948 27019 7988 27028
rect 7756 26851 7796 26860
rect 7948 26900 7988 26909
rect 7852 26816 7892 26825
rect 7660 25171 7700 25180
rect 7756 26732 7796 26741
rect 7564 24331 7604 24340
rect 7180 21559 7220 21568
rect 7276 23668 7412 23708
rect 7084 20131 7124 20140
rect 7180 20852 7220 20861
rect 7180 20096 7220 20812
rect 7180 20047 7220 20056
rect 7084 20012 7124 20021
rect 7084 19877 7124 19972
rect 6988 18451 7028 18460
rect 7180 19256 7220 19265
rect 7180 18416 7220 19216
rect 7276 18668 7316 23668
rect 7372 23120 7412 23129
rect 7372 23036 7412 23080
rect 7372 22985 7412 22996
rect 7564 22868 7604 22877
rect 7468 22364 7508 22373
rect 7372 21608 7412 21617
rect 7372 18836 7412 21568
rect 7372 18787 7412 18796
rect 7276 18619 7316 18628
rect 7180 18367 7220 18376
rect 7276 18500 7316 18509
rect 7180 17576 7220 17585
rect 7084 17492 7124 17501
rect 6988 16232 7028 16327
rect 6988 16183 7028 16192
rect 6988 15980 7028 15989
rect 6988 15728 7028 15940
rect 6988 14888 7028 15688
rect 6988 14839 7028 14848
rect 7084 14804 7124 17452
rect 7180 17441 7220 17536
rect 7276 17240 7316 18460
rect 7276 17191 7316 17200
rect 7372 17828 7412 17837
rect 7180 16484 7220 16493
rect 7180 16349 7220 16444
rect 7180 15476 7220 15485
rect 7180 14972 7220 15436
rect 7180 14923 7220 14932
rect 7276 15224 7316 15233
rect 7084 14764 7220 14804
rect 6892 11192 6932 13420
rect 6988 14720 7028 14729
rect 6988 11780 7028 14680
rect 7084 14552 7124 14561
rect 7084 13964 7124 14512
rect 7084 13915 7124 13924
rect 6988 11731 7028 11740
rect 7084 13796 7124 13805
rect 6892 11143 6932 11152
rect 6796 10984 7028 11024
rect 6740 10900 6836 10940
rect 6700 10891 6740 10900
rect 6412 8539 6452 8548
rect 6508 9388 6644 9428
rect 6220 7916 6260 7925
rect 6220 7328 6260 7876
rect 6220 6992 6260 7288
rect 6220 6943 6260 6952
rect 6028 6775 6068 6784
rect 6124 6908 6164 6917
rect 6124 6773 6164 6868
rect 5740 6196 5972 6236
rect 6316 6320 6356 8044
rect 5740 2792 5780 6196
rect 5836 5984 5876 5993
rect 5836 2876 5876 5944
rect 6316 5732 6356 6280
rect 6316 5683 6356 5692
rect 6412 8252 6452 8261
rect 6412 2900 6452 8212
rect 6508 5816 6548 9388
rect 6796 9344 6836 10900
rect 6892 10856 6932 10865
rect 6892 10688 6932 10816
rect 6892 10639 6932 10648
rect 6604 9260 6644 9269
rect 6604 5984 6644 9220
rect 6700 8840 6740 8935
rect 6700 8791 6740 8800
rect 6700 8672 6740 8681
rect 6796 8672 6836 9304
rect 6892 8672 6932 8681
rect 6796 8632 6892 8672
rect 6700 7412 6740 8632
rect 6892 8623 6932 8632
rect 6700 7363 6740 7372
rect 6988 6572 7028 10984
rect 7084 10352 7124 13756
rect 7180 13292 7220 14764
rect 7276 14720 7316 15184
rect 7372 14972 7412 17788
rect 7468 16988 7508 22324
rect 7564 20852 7604 22828
rect 7564 20180 7604 20812
rect 7564 20140 7700 20180
rect 7660 18500 7700 20140
rect 7660 18451 7700 18460
rect 7564 18332 7604 18341
rect 7564 17660 7604 18292
rect 7564 17611 7604 17620
rect 7660 18248 7700 18257
rect 7468 16939 7508 16948
rect 7564 16988 7604 16997
rect 7372 14923 7412 14932
rect 7468 16232 7508 16241
rect 7276 14671 7316 14680
rect 7468 14384 7508 16192
rect 7276 14344 7508 14384
rect 7276 13544 7316 14344
rect 7468 14216 7508 14225
rect 7372 14048 7412 14057
rect 7372 13880 7412 14008
rect 7372 13831 7412 13840
rect 7276 13495 7316 13504
rect 7372 13460 7412 13555
rect 7372 13411 7412 13420
rect 7372 13292 7412 13301
rect 7180 13252 7372 13292
rect 7372 13243 7412 13252
rect 7084 10303 7124 10312
rect 7180 12872 7220 12881
rect 7180 9176 7220 12832
rect 6988 6523 7028 6532
rect 7084 8756 7124 8765
rect 6604 5935 6644 5944
rect 6892 6404 6932 6413
rect 6508 5312 6548 5776
rect 6892 5732 6932 6364
rect 6508 4892 6548 5272
rect 6508 4843 6548 4852
rect 6700 5480 6740 5489
rect 6700 4472 6740 5440
rect 6892 4556 6932 5692
rect 7084 5480 7124 8716
rect 7180 7916 7220 9136
rect 7180 7867 7220 7876
rect 7276 12032 7316 12041
rect 7084 5431 7124 5440
rect 7276 4808 7316 11992
rect 7372 11024 7412 11033
rect 7372 8924 7412 10984
rect 7372 8756 7412 8884
rect 7372 8707 7412 8716
rect 7276 4759 7316 4768
rect 7372 5396 7412 5405
rect 6892 4507 6932 4516
rect 6700 4423 6740 4432
rect 5836 2827 5876 2836
rect 6316 2860 6452 2900
rect 6700 3128 6740 3137
rect 5740 2743 5780 2752
rect 5644 2407 5684 2416
rect 5836 2624 5876 2633
rect 5548 2071 5588 2080
rect 5644 2036 5684 2045
rect 5548 1868 5588 1877
rect 5548 1028 5588 1828
rect 5548 979 5588 988
rect 5644 80 5684 1996
rect 5836 80 5876 2584
rect 6028 2372 6068 2381
rect 6028 2237 6068 2332
rect 6316 2120 6356 2860
rect 6316 2071 6356 2080
rect 6700 2120 6740 3088
rect 7276 2456 7316 2465
rect 6700 2071 6740 2080
rect 6892 2120 6932 2129
rect 6892 1985 6932 2080
rect 7084 2036 7124 2045
rect 6412 1952 6452 1961
rect 6028 1868 6068 1877
rect 6028 80 6068 1828
rect 6220 1868 6260 1877
rect 6220 80 6260 1828
rect 6412 80 6452 1912
rect 6604 1952 6644 1961
rect 6604 80 6644 1912
rect 6988 1952 7028 1961
rect 6796 1868 6836 1877
rect 6796 80 6836 1828
rect 6988 80 7028 1912
rect 7084 1901 7124 1996
rect 7276 2036 7316 2416
rect 7276 1987 7316 1996
rect 7180 1196 7220 1205
rect 7180 80 7220 1156
rect 7372 80 7412 5356
rect 7468 5144 7508 14176
rect 7564 11864 7604 16948
rect 7660 15476 7700 18208
rect 7756 17996 7796 26692
rect 7852 26564 7892 26776
rect 7948 26648 7988 26860
rect 7948 26599 7988 26608
rect 7852 26515 7892 26524
rect 7948 26144 7988 26155
rect 7948 26060 7988 26104
rect 7948 26011 7988 26020
rect 7852 25556 7892 25565
rect 7852 25388 7892 25516
rect 7852 24884 7892 25348
rect 7852 24835 7892 24844
rect 8044 24716 8084 31984
rect 8140 31856 8180 31865
rect 8140 27320 8180 31816
rect 8236 31352 8276 32824
rect 8236 31303 8276 31312
rect 8332 32696 8372 32705
rect 8236 31184 8276 31193
rect 8236 29924 8276 31144
rect 8236 29875 8276 29884
rect 8332 28580 8372 32656
rect 8332 28531 8372 28540
rect 8332 28412 8372 28421
rect 8332 27824 8372 28372
rect 8332 27775 8372 27784
rect 8332 27572 8372 27581
rect 8140 27280 8276 27320
rect 8140 26816 8180 26825
rect 8140 26144 8180 26776
rect 8140 25976 8180 26104
rect 8140 25927 8180 25936
rect 8044 24667 8084 24676
rect 7948 24632 7988 24641
rect 7852 24548 7892 24557
rect 7852 24044 7892 24508
rect 7852 23995 7892 24004
rect 7948 23624 7988 24592
rect 7852 23204 7892 23213
rect 7852 23120 7892 23164
rect 7852 23069 7892 23080
rect 7852 22952 7892 22961
rect 7852 19928 7892 22912
rect 7948 22448 7988 23584
rect 7948 22399 7988 22408
rect 8044 24128 8084 24137
rect 8044 22364 8084 24088
rect 8044 22315 8084 22324
rect 8140 23120 8180 23129
rect 8044 21860 8084 21869
rect 7852 19879 7892 19888
rect 7948 21608 7988 21617
rect 7852 19760 7892 19769
rect 7852 19256 7892 19720
rect 7852 18584 7892 19216
rect 7852 18535 7892 18544
rect 7756 17947 7796 17956
rect 7852 17828 7892 17837
rect 7948 17828 7988 21568
rect 8044 20600 8084 21820
rect 8044 20551 8084 20560
rect 8140 20768 8180 23080
rect 8044 19172 8084 19181
rect 8044 18164 8084 19132
rect 8140 18500 8180 20728
rect 8140 18365 8180 18460
rect 8044 18115 8084 18124
rect 7892 17788 7988 17828
rect 8044 17996 8084 18005
rect 7852 17072 7892 17788
rect 7852 17023 7892 17032
rect 7948 16988 7988 16997
rect 7660 15427 7700 15436
rect 7852 16904 7892 16913
rect 7756 14300 7796 14309
rect 7660 13880 7700 13889
rect 7660 13208 7700 13840
rect 7660 13159 7700 13168
rect 7564 11815 7604 11824
rect 7660 13040 7700 13049
rect 7564 10772 7604 10781
rect 7564 10268 7604 10732
rect 7564 10219 7604 10228
rect 7564 9428 7604 9437
rect 7564 8588 7604 9388
rect 7660 9008 7700 13000
rect 7660 8959 7700 8968
rect 7564 7244 7604 8548
rect 7564 7195 7604 7204
rect 7468 5095 7508 5104
rect 7756 4388 7796 14260
rect 7852 13964 7892 16864
rect 7948 16400 7988 16948
rect 7948 16351 7988 16360
rect 7892 13924 7988 13964
rect 7852 13915 7892 13924
rect 7852 13796 7892 13805
rect 7852 13208 7892 13756
rect 7852 13159 7892 13168
rect 7852 12704 7892 12713
rect 7852 12536 7892 12664
rect 7852 12487 7892 12496
rect 7948 11024 7988 13924
rect 8044 12620 8084 17956
rect 8140 17828 8180 17837
rect 8140 17240 8180 17788
rect 8140 17191 8180 17200
rect 8140 14384 8180 14393
rect 8140 13964 8180 14344
rect 8140 13915 8180 13924
rect 8044 12571 8084 12580
rect 8140 12788 8180 12797
rect 8140 12452 8180 12748
rect 8044 12412 8180 12452
rect 8044 11864 8084 12412
rect 8044 11815 8084 11824
rect 8140 12284 8180 12293
rect 7948 10975 7988 10984
rect 8140 11780 8180 12244
rect 8044 10940 8084 10949
rect 7852 10772 7892 10781
rect 7852 10184 7892 10732
rect 8044 10436 8084 10900
rect 8044 10387 8084 10396
rect 7852 10135 7892 10144
rect 7948 10016 7988 10025
rect 7852 8756 7892 8765
rect 7852 8168 7892 8716
rect 7852 8119 7892 8128
rect 7948 6656 7988 9976
rect 7948 6607 7988 6616
rect 8140 7916 8180 11740
rect 8140 7244 8180 7876
rect 8044 6404 8084 6413
rect 7756 4339 7796 4348
rect 7948 5564 7988 5573
rect 7756 3380 7796 3389
rect 7756 2120 7796 3340
rect 7756 2071 7796 2080
rect 7756 1448 7796 1457
rect 7564 356 7604 365
rect 7564 80 7604 316
rect 7756 80 7796 1408
rect 7948 80 7988 5524
rect 8044 5144 8084 6364
rect 8044 5095 8084 5104
rect 8140 5732 8180 7204
rect 8140 4892 8180 5692
rect 8140 4843 8180 4852
rect 8236 1952 8276 27280
rect 8332 27068 8372 27532
rect 8332 27019 8372 27028
rect 8332 23792 8372 23801
rect 8332 22868 8372 23752
rect 8428 23120 8468 32908
rect 8524 28916 8564 36016
rect 8524 28867 8564 28876
rect 8620 33200 8660 33209
rect 8524 26900 8564 26909
rect 8524 26060 8564 26860
rect 8524 26011 8564 26020
rect 8428 23071 8468 23080
rect 8524 24632 8564 24641
rect 8332 22819 8372 22828
rect 8332 22616 8372 22711
rect 8332 22567 8372 22576
rect 8332 22364 8372 22373
rect 8332 21860 8372 22324
rect 8428 22280 8468 22289
rect 8428 22145 8468 22240
rect 8332 21811 8372 21820
rect 8332 21440 8372 21449
rect 8332 20936 8372 21400
rect 8332 20887 8372 20896
rect 8332 19340 8372 19349
rect 8332 19205 8372 19300
rect 8428 19256 8468 19265
rect 8428 18920 8468 19216
rect 8428 18871 8468 18880
rect 8524 18668 8564 24592
rect 8620 23960 8660 33160
rect 8716 31520 8756 40720
rect 8812 40256 8852 47776
rect 8908 47060 8948 47860
rect 8908 46556 8948 47020
rect 8908 46507 8948 46516
rect 8908 45800 8948 45809
rect 8908 44960 8948 45760
rect 8908 44911 8948 44920
rect 8908 44204 8948 44213
rect 8908 43616 8948 44164
rect 8908 43567 8948 43576
rect 9004 40424 9044 50296
rect 8812 40207 8852 40216
rect 8908 40340 8948 40349
rect 8908 40256 8948 40300
rect 8908 40205 8948 40216
rect 8812 40088 8852 40097
rect 8812 39248 8852 40048
rect 8812 38996 8852 39208
rect 8908 39164 8948 39173
rect 9004 39164 9044 40384
rect 8948 39124 9044 39164
rect 8908 39115 8948 39124
rect 8812 37316 8852 38956
rect 8812 37267 8852 37276
rect 9100 36560 9140 50464
rect 9196 50420 9236 54748
rect 9292 54620 9332 54629
rect 9292 54116 9332 54580
rect 9292 54067 9332 54076
rect 9292 53024 9332 53033
rect 9292 52604 9332 52984
rect 9292 52555 9332 52564
rect 9196 50371 9236 50380
rect 9292 51680 9332 51689
rect 9292 50084 9332 51640
rect 9292 50035 9332 50044
rect 9196 48824 9236 48835
rect 9196 48740 9236 48784
rect 9196 48691 9236 48700
rect 9388 47480 9428 61720
rect 9484 61004 9524 61972
rect 9580 61172 9620 79948
rect 9676 79904 9716 79999
rect 9676 79855 9716 79864
rect 9676 79736 9716 79747
rect 9676 79652 9716 79696
rect 9676 79603 9716 79612
rect 9676 79148 9716 79157
rect 9676 70580 9716 79108
rect 9772 72764 9812 81208
rect 9868 78056 9908 85240
rect 9964 83684 10004 90952
rect 10636 89732 10676 89741
rect 10060 89480 10100 89489
rect 10060 89345 10100 89440
rect 10636 88808 10676 89692
rect 10540 88640 10580 88649
rect 10348 88472 10388 88481
rect 9964 83635 10004 83644
rect 10060 87716 10100 87725
rect 10060 86792 10100 87676
rect 9964 83516 10004 83525
rect 9964 83381 10004 83476
rect 9964 82004 10004 82013
rect 9964 78224 10004 81964
rect 10060 80576 10100 86752
rect 10252 85868 10292 85877
rect 10156 85028 10196 85037
rect 10156 80744 10196 84988
rect 10252 85028 10292 85828
rect 10252 84356 10292 84988
rect 10252 84307 10292 84316
rect 10252 82844 10292 82853
rect 10252 82004 10292 82804
rect 10252 81955 10292 81964
rect 10156 80695 10196 80704
rect 10060 80536 10292 80576
rect 10060 80408 10100 80417
rect 10060 78308 10100 80368
rect 10060 78259 10100 78268
rect 10156 78728 10196 78737
rect 9964 78175 10004 78184
rect 9868 77552 9908 78016
rect 9868 77503 9908 77512
rect 9868 77384 9908 77393
rect 9868 77249 9908 77344
rect 9868 76796 9908 76805
rect 9868 76208 9908 76756
rect 9868 76159 9908 76168
rect 9964 76628 10004 76637
rect 9964 75956 10004 76588
rect 10060 76460 10100 76469
rect 10060 76325 10100 76420
rect 9772 72715 9812 72724
rect 9868 75916 10004 75956
rect 9772 72260 9812 72269
rect 9772 71000 9812 72220
rect 9772 70951 9812 70960
rect 9676 70531 9716 70540
rect 9772 70748 9812 70757
rect 9772 69908 9812 70708
rect 9772 69859 9812 69868
rect 9868 69152 9908 75916
rect 10060 75452 10100 75461
rect 10060 75317 10100 75412
rect 10060 73352 10100 73361
rect 10060 73217 10100 73312
rect 9964 72176 10004 72185
rect 9964 72041 10004 72136
rect 10060 70664 10100 70673
rect 10060 70496 10100 70624
rect 10060 70447 10100 70456
rect 9868 69112 10004 69152
rect 9772 69068 9812 69077
rect 9676 68648 9716 68657
rect 9676 67640 9716 68608
rect 9676 66800 9716 67600
rect 9676 66751 9716 66760
rect 9676 65288 9716 65297
rect 9676 64868 9716 65248
rect 9676 64819 9716 64828
rect 9676 63944 9716 63953
rect 9676 63356 9716 63904
rect 9676 63307 9716 63316
rect 9676 63188 9716 63197
rect 9676 62600 9716 63148
rect 9676 62551 9716 62560
rect 9580 61123 9620 61132
rect 9484 60964 9620 61004
rect 9484 60836 9524 60845
rect 9484 58904 9524 60796
rect 9484 57224 9524 58864
rect 9484 57175 9524 57184
rect 9580 58568 9620 60964
rect 9772 60836 9812 69028
rect 9868 68984 9908 68993
rect 9868 68396 9908 68944
rect 9868 68347 9908 68356
rect 9868 68228 9908 68237
rect 9868 64280 9908 68188
rect 9964 65960 10004 69112
rect 10060 68648 10100 68657
rect 10060 68513 10100 68608
rect 10060 68144 10100 68153
rect 10060 68009 10100 68104
rect 9964 65911 10004 65920
rect 10156 66884 10196 78688
rect 10252 78392 10292 80536
rect 10348 78476 10388 88432
rect 10540 88052 10580 88600
rect 10540 88003 10580 88012
rect 10636 88136 10676 88768
rect 10444 87716 10484 87725
rect 10444 86792 10484 87676
rect 10444 86743 10484 86752
rect 10636 86540 10676 88096
rect 10732 88892 10772 88901
rect 10732 87296 10772 88852
rect 10732 86876 10772 87256
rect 10732 86827 10772 86836
rect 10828 86540 10868 91372
rect 11020 90236 11060 90245
rect 10636 86491 10676 86500
rect 10732 86500 10868 86540
rect 10924 88724 10964 88733
rect 10924 88136 10964 88684
rect 10444 85616 10484 85625
rect 10444 85481 10484 85576
rect 10636 85448 10676 85457
rect 10540 85280 10580 85289
rect 10444 84860 10484 84869
rect 10444 82844 10484 84820
rect 10444 82795 10484 82804
rect 10348 78427 10388 78436
rect 10444 82088 10484 82097
rect 10444 81248 10484 82048
rect 10444 80576 10484 81208
rect 10252 77132 10292 78352
rect 10252 77083 10292 77092
rect 10348 78308 10388 78317
rect 10348 77468 10388 78268
rect 10444 78140 10484 80536
rect 10540 79064 10580 85240
rect 10636 85028 10676 85408
rect 10636 84979 10676 84988
rect 10636 84356 10676 84365
rect 10636 84188 10676 84316
rect 10636 84139 10676 84148
rect 10636 83684 10676 83693
rect 10636 82088 10676 83644
rect 10636 82039 10676 82048
rect 10732 81920 10772 86500
rect 10636 81880 10772 81920
rect 10828 84272 10868 84281
rect 10828 83516 10868 84232
rect 10636 80408 10676 81880
rect 10732 81752 10772 81761
rect 10732 80660 10772 81712
rect 10828 81500 10868 83476
rect 10828 81451 10868 81460
rect 10732 80620 10868 80660
rect 10636 80359 10676 80368
rect 10732 80492 10772 80501
rect 10636 80156 10676 80165
rect 10636 79820 10676 80116
rect 10636 79771 10676 79780
rect 10732 79820 10772 80452
rect 10540 79015 10580 79024
rect 10636 79316 10676 79325
rect 10540 78896 10580 78905
rect 10636 78896 10676 79276
rect 10732 79064 10772 79780
rect 10732 79015 10772 79024
rect 10636 78856 10772 78896
rect 10540 78761 10580 78856
rect 10636 78644 10676 78653
rect 10540 78560 10580 78569
rect 10540 78308 10580 78520
rect 10540 78259 10580 78268
rect 10444 78091 10484 78100
rect 10252 76964 10292 76973
rect 10252 76829 10292 76924
rect 10252 76712 10292 76721
rect 10252 75284 10292 76672
rect 10252 75235 10292 75244
rect 10252 75116 10292 75125
rect 10252 74528 10292 75076
rect 10252 74479 10292 74488
rect 10252 73772 10292 73781
rect 10252 71420 10292 73732
rect 10252 71371 10292 71380
rect 10348 71504 10388 77428
rect 10540 77468 10580 77477
rect 10540 77333 10580 77428
rect 10444 77300 10484 77309
rect 10444 77216 10484 77260
rect 10444 77176 10580 77216
rect 10444 76628 10484 76723
rect 10444 76579 10484 76588
rect 10348 70748 10388 71464
rect 10348 70699 10388 70708
rect 10444 76460 10484 76469
rect 10540 76460 10580 77176
rect 10636 76796 10676 78604
rect 10732 77300 10772 78856
rect 10732 77251 10772 77260
rect 10732 77132 10772 77141
rect 10732 76880 10772 77092
rect 10732 76831 10772 76840
rect 10636 76747 10676 76756
rect 10540 76420 10676 76460
rect 10252 70496 10292 70505
rect 10252 69320 10292 70456
rect 10252 69271 10292 69280
rect 10348 69992 10388 70001
rect 10252 69152 10292 69161
rect 10252 68312 10292 69112
rect 10252 68263 10292 68272
rect 10348 69068 10388 69952
rect 10060 65372 10100 65381
rect 9868 64231 9908 64240
rect 9964 65204 10004 65213
rect 9964 63944 10004 65164
rect 10060 64616 10100 65332
rect 10156 65288 10196 66844
rect 10252 68144 10292 68153
rect 10252 65540 10292 68104
rect 10348 67724 10388 69028
rect 10348 67675 10388 67684
rect 10252 65491 10292 65500
rect 10348 67556 10388 67565
rect 10156 64952 10196 65248
rect 10156 64903 10196 64912
rect 10252 65372 10292 65381
rect 10252 64868 10292 65332
rect 10156 64784 10196 64793
rect 10156 64649 10196 64744
rect 10060 64567 10100 64576
rect 10252 64532 10292 64828
rect 9964 63895 10004 63904
rect 10156 64492 10292 64532
rect 10060 63692 10100 63701
rect 9964 63440 10004 63449
rect 9964 62768 10004 63400
rect 9964 62719 10004 62728
rect 9964 62432 10004 62441
rect 9964 62264 10004 62392
rect 10060 62432 10100 63652
rect 10060 62383 10100 62392
rect 10156 62516 10196 64492
rect 10348 63692 10388 67516
rect 10348 63643 10388 63652
rect 10444 63524 10484 76420
rect 10540 76292 10580 76301
rect 10540 70076 10580 76252
rect 10636 73460 10676 76420
rect 10732 76124 10772 76133
rect 10732 75956 10772 76084
rect 10732 75907 10772 75916
rect 10636 73420 10772 73460
rect 10636 72596 10676 72605
rect 10636 72176 10676 72556
rect 10636 72127 10676 72136
rect 10540 70027 10580 70036
rect 10636 71420 10676 71429
rect 10636 70832 10676 71380
rect 10540 69908 10580 69917
rect 10540 69152 10580 69868
rect 10540 67892 10580 69112
rect 10636 67976 10676 70792
rect 10636 67927 10676 67936
rect 10540 67843 10580 67852
rect 10636 65960 10676 65969
rect 10540 65372 10580 65381
rect 10540 64700 10580 65332
rect 10540 64651 10580 64660
rect 10636 64532 10676 65920
rect 9868 62224 9964 62264
rect 9868 61676 9908 62224
rect 9964 62215 10004 62224
rect 9868 61627 9908 61636
rect 9964 62096 10004 62105
rect 9580 55796 9620 58528
rect 9580 54872 9620 55756
rect 9676 60796 9812 60836
rect 9868 61172 9908 61181
rect 9676 58736 9716 60796
rect 9676 55628 9716 58696
rect 9676 54956 9716 55588
rect 9676 54907 9716 54916
rect 9772 60668 9812 60677
rect 9580 54200 9620 54832
rect 9580 54065 9620 54160
rect 9676 54788 9716 54797
rect 9676 54116 9716 54748
rect 9676 54067 9716 54076
rect 9772 53300 9812 60628
rect 9484 53276 9524 53285
rect 9484 52856 9524 53236
rect 9484 52688 9524 52816
rect 9484 51764 9524 52648
rect 9484 51715 9524 51724
rect 9580 53260 9812 53300
rect 9388 47431 9428 47440
rect 9484 49580 9524 49589
rect 9388 47228 9428 47237
rect 9388 46724 9428 47188
rect 9388 46675 9428 46684
rect 9388 45716 9428 45725
rect 9388 45548 9428 45676
rect 9388 45499 9428 45508
rect 9196 45212 9236 45221
rect 9196 44204 9236 45172
rect 9196 44155 9236 44164
rect 9292 44960 9332 44969
rect 9292 43532 9332 44920
rect 9388 44540 9428 44549
rect 9388 44120 9428 44500
rect 9388 44071 9428 44080
rect 9292 43220 9332 43492
rect 9292 43180 9428 43220
rect 9100 36511 9140 36520
rect 9196 40256 9236 40265
rect 9196 38240 9236 40216
rect 9292 39500 9332 39509
rect 9292 39164 9332 39460
rect 9292 39115 9332 39124
rect 8812 36308 8852 36317
rect 8812 34712 8852 36268
rect 9004 35636 9044 35645
rect 8908 34880 8948 34889
rect 8908 34745 8948 34840
rect 8812 34663 8852 34672
rect 8812 34544 8852 34553
rect 8812 33620 8852 34504
rect 8812 33571 8852 33580
rect 8908 34460 8948 34469
rect 8908 33452 8948 34420
rect 8812 33412 8908 33452
rect 8812 32864 8852 33412
rect 8908 33403 8948 33412
rect 8812 32815 8852 32824
rect 8908 33284 8948 33293
rect 8812 32612 8852 32621
rect 8812 32360 8852 32572
rect 8812 32311 8852 32320
rect 8908 32192 8948 33244
rect 9004 33284 9044 35596
rect 9004 32444 9044 33244
rect 9004 32395 9044 32404
rect 9100 34964 9140 34973
rect 9100 32444 9140 34924
rect 9196 34628 9236 38200
rect 9292 36644 9332 36653
rect 9292 35384 9332 36604
rect 9292 35335 9332 35344
rect 9196 34579 9236 34588
rect 8716 31471 8756 31480
rect 8812 32152 8908 32192
rect 8716 30428 8756 30437
rect 8716 29924 8756 30388
rect 8716 29875 8756 29884
rect 8716 29756 8756 29765
rect 8716 29420 8756 29716
rect 8716 29371 8756 29380
rect 8812 29084 8852 32152
rect 8908 32143 8948 32152
rect 9004 30932 9044 30941
rect 8908 30512 8948 30523
rect 8908 30428 8948 30472
rect 8908 30379 8948 30388
rect 8908 29924 8948 29933
rect 8908 29504 8948 29884
rect 8908 29455 8948 29464
rect 9004 29168 9044 30892
rect 9100 30848 9140 32404
rect 9100 30799 9140 30808
rect 9196 34460 9236 34469
rect 9196 30008 9236 34420
rect 9388 32948 9428 43180
rect 9484 41432 9524 49540
rect 9580 48236 9620 53260
rect 9676 53192 9716 53201
rect 9676 52604 9716 53152
rect 9676 51848 9716 52564
rect 9676 51799 9716 51808
rect 9772 53108 9812 53117
rect 9772 50420 9812 53068
rect 9676 50380 9812 50420
rect 9676 48992 9716 50380
rect 9772 50252 9812 50261
rect 9772 49580 9812 50212
rect 9772 49445 9812 49540
rect 9868 48992 9908 61132
rect 9964 58736 10004 62056
rect 10156 61676 10196 62476
rect 10156 61627 10196 61636
rect 10252 63484 10484 63524
rect 10540 64492 10676 64532
rect 10060 60836 10100 60845
rect 10060 60164 10100 60796
rect 10060 60115 10100 60124
rect 9964 58687 10004 58696
rect 10156 59156 10196 59165
rect 10156 58568 10196 59116
rect 10156 57644 10196 58528
rect 9964 56888 10004 56897
rect 9964 56384 10004 56848
rect 10060 56552 10100 56561
rect 10060 56417 10100 56512
rect 9964 56335 10004 56344
rect 9964 56132 10004 56141
rect 9964 55628 10004 56092
rect 10156 55712 10196 57604
rect 10156 55663 10196 55672
rect 9964 55579 10004 55588
rect 9964 54536 10004 54545
rect 9964 54032 10004 54496
rect 9964 53983 10004 53992
rect 10060 53864 10100 53873
rect 9964 53612 10004 53621
rect 10060 53612 10100 53824
rect 10004 53572 10100 53612
rect 9964 53563 10004 53572
rect 10060 53444 10100 53453
rect 9964 53108 10004 53117
rect 9964 52604 10004 53068
rect 9964 52555 10004 52564
rect 9964 52436 10004 52445
rect 9964 51932 10004 52396
rect 9964 51883 10004 51892
rect 10060 51764 10100 53404
rect 10060 51715 10100 51724
rect 10156 53360 10196 53369
rect 10156 51680 10196 53320
rect 10156 51631 10196 51640
rect 10060 50336 10100 50345
rect 10060 50201 10100 50296
rect 10156 50252 10196 50261
rect 10156 50117 10196 50212
rect 10156 49580 10196 49589
rect 10156 49445 10196 49540
rect 10252 49496 10292 63484
rect 10540 63380 10580 64492
rect 10444 63340 10580 63380
rect 10636 64364 10676 64373
rect 10348 63188 10388 63197
rect 10348 60836 10388 63148
rect 10444 62600 10484 63340
rect 10636 62936 10676 64324
rect 10444 62551 10484 62560
rect 10540 62896 10676 62936
rect 10732 63860 10772 73420
rect 10828 73184 10868 80620
rect 10924 78728 10964 88096
rect 10924 78679 10964 78688
rect 11020 78560 11060 90196
rect 11308 88724 11348 94984
rect 11404 94856 11444 96688
rect 11404 94807 11444 94816
rect 11596 94856 11636 96688
rect 11596 94807 11636 94816
rect 11500 94772 11540 94781
rect 11500 94184 11540 94732
rect 11788 94772 11828 96688
rect 11980 94940 12020 96688
rect 11980 94891 12020 94900
rect 12172 94940 12212 96688
rect 12364 95696 12404 96688
rect 12364 95656 12500 95696
rect 12172 94891 12212 94900
rect 11788 94723 11828 94732
rect 12364 94772 12404 94781
rect 11596 94688 11636 94697
rect 11596 94553 11636 94648
rect 12172 94688 12212 94697
rect 11788 94604 11828 94613
rect 11500 94135 11540 94144
rect 11692 94100 11732 94109
rect 11404 90404 11444 90413
rect 11404 89564 11444 90364
rect 11596 89900 11636 89909
rect 11404 89515 11444 89524
rect 11500 89816 11540 89825
rect 11308 88684 11444 88724
rect 11212 88052 11252 88061
rect 11020 78511 11060 78520
rect 11116 87968 11156 87977
rect 10924 78476 10964 78485
rect 10924 78392 10964 78436
rect 10924 78352 11060 78392
rect 10924 76628 10964 76637
rect 10924 76493 10964 76588
rect 10924 76040 10964 76049
rect 10924 75116 10964 76000
rect 10924 75067 10964 75076
rect 10828 73135 10868 73144
rect 10924 73604 10964 73613
rect 10828 72932 10868 72941
rect 10828 72260 10868 72892
rect 10828 69992 10868 72220
rect 10828 69943 10868 69952
rect 10924 68732 10964 73564
rect 11020 73100 11060 78352
rect 11116 73856 11156 87928
rect 11212 86792 11252 88012
rect 11212 86743 11252 86752
rect 11308 87884 11348 87893
rect 11308 87128 11348 87844
rect 11212 84104 11252 84113
rect 11212 83600 11252 84064
rect 11212 83551 11252 83560
rect 11212 80660 11252 80669
rect 11212 80408 11252 80620
rect 11212 80359 11252 80368
rect 11212 79988 11252 79997
rect 11212 79736 11252 79948
rect 11212 79687 11252 79696
rect 11212 79568 11252 79577
rect 11212 79316 11252 79528
rect 11212 79267 11252 79276
rect 11212 79148 11252 79157
rect 11212 78980 11252 79108
rect 11212 78931 11252 78940
rect 11116 73807 11156 73816
rect 11212 78476 11252 78485
rect 11020 73051 11060 73060
rect 11116 73688 11156 73697
rect 11020 72932 11060 72941
rect 11020 72680 11060 72892
rect 11020 70412 11060 72640
rect 11020 69320 11060 70372
rect 11020 69271 11060 69280
rect 10924 68683 10964 68692
rect 11116 68396 11156 73648
rect 11212 72344 11252 78436
rect 11308 72848 11348 87088
rect 11404 83852 11444 88684
rect 11500 84692 11540 89776
rect 11500 84643 11540 84652
rect 11404 83803 11444 83812
rect 11500 84356 11540 84365
rect 11308 72799 11348 72808
rect 11404 83516 11444 83525
rect 11404 82760 11444 83476
rect 11404 82004 11444 82720
rect 11404 81332 11444 81964
rect 11404 79652 11444 81292
rect 11212 72304 11348 72344
rect 10540 62348 10580 62896
rect 10348 60787 10388 60796
rect 10444 62308 10580 62348
rect 10636 62768 10676 62777
rect 10348 59408 10388 59417
rect 10348 59324 10388 59368
rect 10348 59273 10388 59284
rect 10444 58652 10484 62308
rect 10348 58612 10484 58652
rect 10540 58652 10580 58661
rect 10348 53864 10388 58612
rect 10444 58484 10484 58493
rect 10444 58400 10484 58444
rect 10444 58349 10484 58360
rect 10540 58064 10580 58612
rect 10540 58015 10580 58024
rect 10540 57812 10580 57821
rect 10540 57677 10580 57772
rect 10636 56972 10676 62728
rect 10732 61844 10772 63820
rect 10828 68356 11156 68396
rect 11212 72176 11252 72185
rect 11212 70664 11252 72136
rect 10828 63188 10868 68356
rect 11212 68312 11252 70624
rect 11308 69908 11348 72304
rect 11308 69859 11348 69868
rect 10828 63139 10868 63148
rect 10924 68272 11252 68312
rect 11308 69740 11348 69749
rect 10732 60164 10772 61804
rect 10732 60115 10772 60124
rect 10828 62348 10868 62357
rect 10828 62180 10868 62308
rect 10828 61676 10868 62140
rect 10828 59996 10868 61636
rect 10924 60080 10964 68272
rect 11116 67976 11156 67985
rect 11116 67724 11156 67936
rect 11116 67675 11156 67684
rect 11116 66716 11156 66725
rect 11020 65960 11060 65969
rect 11020 65372 11060 65920
rect 11020 65323 11060 65332
rect 11116 64700 11156 66676
rect 11212 66128 11252 66137
rect 11212 65876 11252 66088
rect 11212 65827 11252 65836
rect 11212 65204 11252 65213
rect 11212 65069 11252 65164
rect 11116 64651 11156 64660
rect 11212 64952 11252 64961
rect 10924 60031 10964 60040
rect 11020 64616 11060 64625
rect 11020 62936 11060 64576
rect 11116 64448 11156 64457
rect 11116 63524 11156 64408
rect 11116 63475 11156 63484
rect 10540 56932 10676 56972
rect 10732 59956 10868 59996
rect 10444 54788 10484 54797
rect 10444 54116 10484 54748
rect 10444 54067 10484 54076
rect 10348 53815 10388 53824
rect 10444 53864 10484 53873
rect 10444 53444 10484 53824
rect 10444 53395 10484 53404
rect 10348 53360 10388 53369
rect 10348 52772 10388 53320
rect 10540 53108 10580 56932
rect 10732 54872 10772 59956
rect 10828 59828 10868 59837
rect 10828 59492 10868 59788
rect 10828 59443 10868 59452
rect 10828 59324 10868 59333
rect 10828 59156 10868 59284
rect 10828 59107 10868 59116
rect 10828 58568 10868 58577
rect 10828 57644 10868 58528
rect 10924 58484 10964 58493
rect 10924 58148 10964 58444
rect 11020 58400 11060 62896
rect 11116 61844 11156 61853
rect 11116 61709 11156 61804
rect 11116 61592 11156 61601
rect 11116 61088 11156 61552
rect 11116 61039 11156 61048
rect 11212 59996 11252 64912
rect 11308 64196 11348 69700
rect 11308 64147 11348 64156
rect 11404 66884 11444 79612
rect 11500 77384 11540 84316
rect 11500 75956 11540 77344
rect 11500 75907 11540 75916
rect 11500 75284 11540 75293
rect 11500 74444 11540 75244
rect 11500 73940 11540 74404
rect 11500 73891 11540 73900
rect 11500 73772 11540 73781
rect 11500 73016 11540 73732
rect 11596 73436 11636 89860
rect 11692 89060 11732 94060
rect 11692 89011 11732 89020
rect 11692 86708 11732 86717
rect 11692 84776 11732 86668
rect 11692 84727 11732 84736
rect 11788 83540 11828 94564
rect 12172 94553 12212 94648
rect 12364 94637 12404 94732
rect 12460 94604 12500 95656
rect 12460 94555 12500 94564
rect 12556 94184 12596 96688
rect 12748 95024 12788 96688
rect 12940 96368 12980 96688
rect 12748 94975 12788 94984
rect 12844 96328 12980 96368
rect 12844 94268 12884 96328
rect 13132 94940 13172 96688
rect 13132 94891 13172 94900
rect 13228 94772 13268 94781
rect 13036 94688 13076 94697
rect 12940 94268 12980 94277
rect 12844 94228 12940 94268
rect 12940 94219 12980 94228
rect 12556 94135 12596 94144
rect 12076 94016 12116 94025
rect 11980 88892 12020 88901
rect 11980 88052 12020 88852
rect 11980 88003 12020 88012
rect 11884 85868 11924 85877
rect 11884 85028 11924 85828
rect 11884 84356 11924 84988
rect 11980 84524 12020 84533
rect 11980 84389 12020 84484
rect 11884 84307 11924 84316
rect 11596 73387 11636 73396
rect 11692 83516 11828 83540
rect 11732 83500 11828 83516
rect 11980 83600 12020 83609
rect 11692 82760 11732 83476
rect 11692 82004 11732 82720
rect 11692 81248 11732 81964
rect 11692 79820 11732 81208
rect 11788 82844 11828 82853
rect 11788 82088 11828 82804
rect 11980 82844 12020 83560
rect 12076 83516 12116 93976
rect 12652 93932 12692 93941
rect 12268 93764 12308 93773
rect 12172 88892 12212 88901
rect 12172 88304 12212 88852
rect 12172 88255 12212 88264
rect 12076 83467 12116 83476
rect 12172 87380 12212 87389
rect 12172 86540 12212 87340
rect 11980 82795 12020 82804
rect 12076 83348 12116 83357
rect 11788 81332 11828 82048
rect 11788 80660 11828 81292
rect 11788 80611 11828 80620
rect 11884 81836 11924 81845
rect 11788 80408 11828 80417
rect 11788 79988 11828 80368
rect 11788 79939 11828 79948
rect 11500 72428 11540 72976
rect 11500 72379 11540 72388
rect 11500 72260 11540 72269
rect 11500 71420 11540 72220
rect 11500 71371 11540 71380
rect 11596 72008 11636 72017
rect 11500 70412 11540 70421
rect 11500 69236 11540 70372
rect 11500 69187 11540 69196
rect 11212 59947 11252 59956
rect 11308 63608 11348 63617
rect 11116 59660 11156 59669
rect 11116 59324 11156 59620
rect 11116 59275 11156 59284
rect 11212 59408 11252 59417
rect 11212 58988 11252 59368
rect 11212 58939 11252 58948
rect 11020 58351 11060 58360
rect 11116 58652 11156 58661
rect 10924 58099 10964 58108
rect 11116 58148 11156 58612
rect 11212 58568 11252 58579
rect 11212 58484 11252 58528
rect 11212 58435 11252 58444
rect 11308 58316 11348 63568
rect 11116 58099 11156 58108
rect 11212 58276 11348 58316
rect 10924 57980 10964 57989
rect 10924 57845 10964 57940
rect 11020 57896 11060 57905
rect 10828 57308 10868 57604
rect 10924 57728 10964 57737
rect 10924 57593 10964 57688
rect 10828 57259 10868 57268
rect 10636 53864 10676 53873
rect 10636 53729 10676 53824
rect 10636 53444 10676 53453
rect 10636 53309 10676 53404
rect 10540 53059 10580 53068
rect 10732 53024 10772 54832
rect 10732 52975 10772 52984
rect 10828 56300 10868 56309
rect 10348 52723 10388 52732
rect 10732 52772 10772 52781
rect 10540 52688 10580 52697
rect 10444 52604 10484 52613
rect 10348 52520 10388 52529
rect 10348 51764 10388 52480
rect 10444 52100 10484 52564
rect 10444 52051 10484 52060
rect 10540 51848 10580 52648
rect 10732 52637 10772 52732
rect 10636 52520 10676 52529
rect 10636 52016 10676 52480
rect 10636 51967 10676 51976
rect 10540 51799 10580 51808
rect 10348 51715 10388 51724
rect 10828 51092 10868 56260
rect 10924 55376 10964 55385
rect 10924 54116 10964 55336
rect 10924 54067 10964 54076
rect 10924 53444 10964 53539
rect 10924 53395 10964 53404
rect 10924 52436 10964 52445
rect 10924 52016 10964 52396
rect 10924 51967 10964 51976
rect 10828 51043 10868 51052
rect 10444 51008 10484 51017
rect 10348 50840 10388 50849
rect 10348 50252 10388 50800
rect 10348 50203 10388 50212
rect 10444 49664 10484 50968
rect 11020 51008 11060 57856
rect 11020 50504 11060 50968
rect 11020 50455 11060 50464
rect 11116 57812 11156 57821
rect 11116 57140 11156 57772
rect 11116 50504 11156 57100
rect 10444 49615 10484 49624
rect 10924 49748 10964 49757
rect 10252 49447 10292 49456
rect 10732 49580 10772 49589
rect 10732 49445 10772 49540
rect 9676 48952 9812 48992
rect 9868 48980 10100 48992
rect 9868 48952 10292 48980
rect 9676 48824 9716 48833
rect 9676 48689 9716 48784
rect 9580 48196 9716 48236
rect 9484 41383 9524 41392
rect 9580 46556 9620 46565
rect 9484 40676 9524 40685
rect 9484 40424 9524 40636
rect 9484 39668 9524 40384
rect 9484 39619 9524 39628
rect 9484 39416 9524 39425
rect 9484 39281 9524 39376
rect 9484 38240 9524 38249
rect 9484 37820 9524 38200
rect 9484 37736 9524 37780
rect 9484 37685 9524 37696
rect 9484 36728 9524 36737
rect 9484 35300 9524 36688
rect 9484 33284 9524 35260
rect 9580 34460 9620 46516
rect 9580 33620 9620 34420
rect 9580 33571 9620 33580
rect 9484 33235 9524 33244
rect 9580 33452 9620 33461
rect 9580 33032 9620 33412
rect 9580 32983 9620 32992
rect 9100 29840 9140 29851
rect 9100 29756 9140 29800
rect 9100 29707 9140 29716
rect 9004 29119 9044 29128
rect 8716 28664 8756 28673
rect 8716 28244 8756 28624
rect 8716 28195 8756 28204
rect 8812 26816 8852 29044
rect 8908 29084 8948 29093
rect 8908 27488 8948 29044
rect 9100 28916 9140 28925
rect 9004 28832 9044 28841
rect 9004 28580 9044 28792
rect 9004 28531 9044 28540
rect 8908 27439 8948 27448
rect 9004 28328 9044 28337
rect 8812 26144 8852 26776
rect 8812 26095 8852 26104
rect 8908 26900 8948 26909
rect 8908 26060 8948 26860
rect 8620 23911 8660 23920
rect 8812 24884 8852 24893
rect 8812 24464 8852 24844
rect 8620 22448 8660 22457
rect 8620 21776 8660 22408
rect 8716 22280 8756 22289
rect 8716 22112 8756 22240
rect 8716 22063 8756 22072
rect 8620 21727 8660 21736
rect 8812 21188 8852 24424
rect 8812 21139 8852 21148
rect 8908 21188 8948 26020
rect 9004 25808 9044 28288
rect 9004 24716 9044 25768
rect 9100 26396 9140 28876
rect 9196 27572 9236 29968
rect 9292 32276 9332 32285
rect 9292 31268 9332 32236
rect 9388 32192 9428 32908
rect 9580 32864 9620 32873
rect 9388 32143 9428 32152
rect 9484 32276 9524 32285
rect 9580 32276 9620 32824
rect 9676 32696 9716 48196
rect 9772 46640 9812 48952
rect 10060 48940 10292 48952
rect 9964 48740 10004 48749
rect 9772 46600 9908 46640
rect 9772 46472 9812 46481
rect 9772 45968 9812 46432
rect 9772 45919 9812 45928
rect 9868 44540 9908 46600
rect 9868 44491 9908 44500
rect 9772 44288 9812 44297
rect 9772 42944 9812 44248
rect 9868 44204 9908 44213
rect 9868 44069 9908 44164
rect 9772 42895 9812 42904
rect 9868 43868 9908 43877
rect 9868 43280 9908 43828
rect 9868 42692 9908 43240
rect 9868 42643 9908 42652
rect 9868 42020 9908 42029
rect 9772 41936 9812 41945
rect 9772 40676 9812 41896
rect 9772 40627 9812 40636
rect 9772 40508 9812 40548
rect 9772 40424 9812 40468
rect 9772 39836 9812 40384
rect 9772 39787 9812 39796
rect 9772 35972 9812 35981
rect 9772 35132 9812 35932
rect 9772 35083 9812 35092
rect 9868 34460 9908 41980
rect 9964 40760 10004 48700
rect 10252 46556 10292 48940
rect 10636 48740 10676 48749
rect 10636 47900 10676 48700
rect 10540 47816 10580 47825
rect 10444 47228 10484 47237
rect 10156 46472 10196 46481
rect 10156 45968 10196 46432
rect 10252 46421 10292 46516
rect 10348 46724 10388 46733
rect 10156 45919 10196 45928
rect 10156 45800 10196 45809
rect 10156 45044 10196 45760
rect 10348 45128 10388 46684
rect 10444 46640 10484 47188
rect 10444 46591 10484 46600
rect 10444 46472 10484 46481
rect 10444 45212 10484 46432
rect 10444 45163 10484 45172
rect 10348 45079 10388 45088
rect 10156 44995 10196 45004
rect 10348 44288 10388 44297
rect 10252 44036 10292 44045
rect 10252 41768 10292 43996
rect 10156 41180 10196 41189
rect 10156 41045 10196 41140
rect 9964 40711 10004 40720
rect 9964 40592 10004 40601
rect 9964 40340 10004 40552
rect 10252 40508 10292 41728
rect 10348 40844 10388 44248
rect 10540 44288 10580 47776
rect 10636 47765 10676 47860
rect 10732 47816 10772 47825
rect 10732 47648 10772 47776
rect 10636 46472 10676 46481
rect 10636 45968 10676 46432
rect 10636 45919 10676 45928
rect 10540 44239 10580 44248
rect 10636 44960 10676 44969
rect 10540 44120 10580 44129
rect 10444 42776 10484 42785
rect 10444 42188 10484 42736
rect 10444 42139 10484 42148
rect 10348 40795 10388 40804
rect 10252 40459 10292 40468
rect 10060 40340 10100 40349
rect 9964 40300 10060 40340
rect 10060 40272 10100 40300
rect 9964 40172 10004 40181
rect 9964 39080 10004 40132
rect 10060 39836 10100 39847
rect 10060 39752 10100 39796
rect 10060 39703 10100 39712
rect 10252 39836 10292 39845
rect 10156 39584 10196 39593
rect 10060 39416 10100 39425
rect 10060 39281 10100 39376
rect 9964 39031 10004 39040
rect 9964 38324 10004 38333
rect 9964 37484 10004 38284
rect 9964 37435 10004 37444
rect 10060 37568 10100 37577
rect 10060 37433 10100 37528
rect 9868 34411 9908 34420
rect 9964 36644 10004 36653
rect 9868 33536 9908 33545
rect 9868 33140 9908 33496
rect 9676 32647 9716 32656
rect 9772 33100 9908 33140
rect 9580 32236 9716 32276
rect 9388 32024 9428 32033
rect 9388 31940 9428 31984
rect 9388 31889 9428 31900
rect 9292 29840 9332 31228
rect 9292 29791 9332 29800
rect 9388 29756 9428 29765
rect 9292 29672 9332 29681
rect 9292 29537 9332 29632
rect 9388 29621 9428 29716
rect 9292 29420 9332 29429
rect 9292 29285 9332 29380
rect 9484 29252 9524 32236
rect 9580 32024 9620 32033
rect 9580 30764 9620 31984
rect 9676 31436 9716 32236
rect 9676 31387 9716 31396
rect 9772 32192 9812 33100
rect 9580 30715 9620 30724
rect 9676 29924 9716 29933
rect 9388 29212 9524 29252
rect 9580 29840 9620 29849
rect 9292 29168 9332 29177
rect 9292 27656 9332 29128
rect 9292 27607 9332 27616
rect 9196 27523 9236 27532
rect 9292 27236 9332 27245
rect 9292 27068 9332 27196
rect 9292 27019 9332 27028
rect 9100 25640 9140 26356
rect 9196 26648 9236 26657
rect 9196 26144 9236 26608
rect 9292 26312 9332 26321
rect 9292 26177 9332 26272
rect 9196 26095 9236 26104
rect 9100 25591 9140 25600
rect 9196 25892 9236 25901
rect 9004 24667 9044 24676
rect 9100 25472 9140 25512
rect 9100 25388 9140 25432
rect 9100 25136 9140 25348
rect 9100 23876 9140 25096
rect 9196 23876 9236 25852
rect 9292 25388 9332 25397
rect 9292 24044 9332 25348
rect 9388 24800 9428 29212
rect 9388 24751 9428 24760
rect 9484 29084 9524 29093
rect 9292 23995 9332 24004
rect 9388 24380 9428 24389
rect 9196 23836 9332 23876
rect 9100 23827 9140 23836
rect 9100 23708 9140 23717
rect 9004 23120 9044 23215
rect 9004 23071 9044 23080
rect 9004 22952 9044 22961
rect 9004 21776 9044 22912
rect 9004 21727 9044 21736
rect 9100 22364 9140 23668
rect 9100 21692 9140 22324
rect 9100 21643 9140 21652
rect 8908 21139 8948 21148
rect 9100 21440 9140 21449
rect 8716 21020 8756 21029
rect 8332 18628 8564 18668
rect 8620 20852 8660 20861
rect 8332 17492 8372 18628
rect 8524 18500 8564 18509
rect 8332 17443 8372 17452
rect 8428 18416 8468 18425
rect 8428 17912 8468 18376
rect 8332 17072 8372 17081
rect 8332 4388 8372 17032
rect 8332 4339 8372 4348
rect 8428 3632 8468 17872
rect 8524 17744 8564 18460
rect 8620 17912 8660 20812
rect 8716 19256 8756 20980
rect 9100 20936 9140 21400
rect 9292 21188 9332 23836
rect 9388 23792 9428 24340
rect 9388 23743 9428 23752
rect 9292 21139 9332 21148
rect 9388 23120 9428 23129
rect 9292 21020 9332 21029
rect 9100 20887 9140 20896
rect 9196 20936 9236 20945
rect 9004 20852 9044 20861
rect 8716 19207 8756 19216
rect 8812 20684 8852 20693
rect 8620 17863 8660 17872
rect 8716 18584 8756 18593
rect 8524 17695 8564 17704
rect 8524 17492 8564 17501
rect 8524 15056 8564 17452
rect 8716 17492 8756 18544
rect 8812 17828 8852 20644
rect 8908 20012 8948 20021
rect 8908 19676 8948 19972
rect 9004 19928 9044 20812
rect 9004 19879 9044 19888
rect 9100 20600 9140 20609
rect 8908 19627 8948 19636
rect 9100 19256 9140 20560
rect 9100 19207 9140 19216
rect 8812 17779 8852 17788
rect 8908 18920 8948 18929
rect 8756 17452 8852 17492
rect 8716 17443 8756 17452
rect 8716 16316 8756 16325
rect 8620 16232 8660 16241
rect 8620 16097 8660 16192
rect 8716 16064 8756 16276
rect 8620 15308 8660 15317
rect 8620 15173 8660 15268
rect 8524 15016 8660 15056
rect 8524 14048 8564 14057
rect 8524 13913 8564 14008
rect 8620 13544 8660 15016
rect 8620 13495 8660 13504
rect 8524 12872 8564 12881
rect 8524 12620 8564 12832
rect 8524 12571 8564 12580
rect 8524 11780 8564 11789
rect 8524 11192 8564 11740
rect 8716 11612 8756 16024
rect 8812 14888 8852 17452
rect 8908 17408 8948 18880
rect 8908 17359 8948 17368
rect 9004 18752 9044 18761
rect 9004 18416 9044 18712
rect 8812 14753 8852 14848
rect 8908 15476 8948 15485
rect 8812 14048 8852 14057
rect 8812 12452 8852 14008
rect 8908 12704 8948 15436
rect 9004 14636 9044 18376
rect 9100 18500 9140 18509
rect 9100 17996 9140 18460
rect 9100 17947 9140 17956
rect 9100 17828 9140 17837
rect 9100 16988 9140 17788
rect 9100 16939 9140 16948
rect 9196 16400 9236 20896
rect 9292 19256 9332 20980
rect 9388 20684 9428 23080
rect 9484 20852 9524 29044
rect 9580 28832 9620 29800
rect 9580 22952 9620 28792
rect 9676 25892 9716 29884
rect 9772 29168 9812 32152
rect 9772 29119 9812 29128
rect 9868 33032 9908 33041
rect 9772 28412 9812 28421
rect 9772 27656 9812 28372
rect 9772 27607 9812 27616
rect 9676 25843 9716 25852
rect 9772 26900 9812 26909
rect 9676 25640 9716 25649
rect 9676 23708 9716 25600
rect 9772 25556 9812 26860
rect 9772 25507 9812 25516
rect 9772 25388 9812 25397
rect 9772 25253 9812 25348
rect 9676 23659 9716 23668
rect 9676 23204 9716 23213
rect 9676 23120 9716 23164
rect 9676 23069 9716 23080
rect 9580 22912 9812 22952
rect 9580 20852 9620 20861
rect 9484 20812 9580 20852
rect 9388 20635 9428 20644
rect 9292 19207 9332 19216
rect 9484 17828 9524 17837
rect 9484 17072 9524 17788
rect 9484 17023 9524 17032
rect 9196 16316 9236 16360
rect 9196 16265 9236 16276
rect 9292 15644 9332 15653
rect 9292 15308 9332 15604
rect 9292 15259 9332 15268
rect 9196 15140 9236 15149
rect 9196 14804 9236 15100
rect 9484 15056 9524 15065
rect 9484 14804 9524 15016
rect 9236 14764 9428 14804
rect 9196 14755 9236 14764
rect 9004 14587 9044 14596
rect 9292 14636 9332 14645
rect 8908 12620 8948 12664
rect 8908 12569 8948 12580
rect 9100 13964 9140 13973
rect 9004 12452 9044 12461
rect 8812 12412 8948 12452
rect 8812 12284 8852 12293
rect 8812 11780 8852 12244
rect 8812 11731 8852 11740
rect 8716 11572 8852 11612
rect 8524 11143 8564 11152
rect 8524 10772 8564 10781
rect 8524 10520 8564 10732
rect 8524 10471 8564 10480
rect 8812 9428 8852 11572
rect 8908 9848 8948 12412
rect 8908 9799 8948 9808
rect 9004 10604 9044 12412
rect 9100 11948 9140 13924
rect 9196 12536 9236 12545
rect 9196 12200 9236 12496
rect 9196 12151 9236 12160
rect 9100 11899 9140 11908
rect 9292 11864 9332 14596
rect 9292 11815 9332 11824
rect 9388 11780 9428 14764
rect 9484 14755 9524 14764
rect 9388 11731 9428 11740
rect 9484 14636 9524 14645
rect 9004 9764 9044 10564
rect 9292 11696 9332 11705
rect 9292 10184 9332 11656
rect 9292 10135 9332 10144
rect 9004 9715 9044 9724
rect 9196 9512 9236 9521
rect 8908 9428 8948 9437
rect 8812 9388 8908 9428
rect 8620 8756 8660 8765
rect 8620 7916 8660 8716
rect 8620 7867 8660 7876
rect 8908 8756 8948 9388
rect 8716 7328 8756 7337
rect 8620 6572 8660 6581
rect 8620 5228 8660 6532
rect 8716 6404 8756 7288
rect 8716 6355 8756 6364
rect 8812 7160 8852 7169
rect 8620 5179 8660 5188
rect 8428 3583 8468 3592
rect 8620 3632 8660 3641
rect 8428 2876 8468 2885
rect 8428 2741 8468 2836
rect 8236 1903 8276 1912
rect 8620 1952 8660 3592
rect 8620 1903 8660 1912
rect 8812 1868 8852 7120
rect 8908 6320 8948 8716
rect 8908 6271 8948 6280
rect 9100 7916 9140 7925
rect 9004 5312 9044 5321
rect 9004 4892 9044 5272
rect 9004 4843 9044 4852
rect 8812 1819 8852 1828
rect 8908 2456 8948 2465
rect 8716 1700 8756 1709
rect 8140 1448 8180 1457
rect 8140 80 8180 1408
rect 8332 1448 8372 1457
rect 8332 80 8372 1408
rect 8524 1448 8564 1457
rect 8524 80 8564 1408
rect 8716 80 8756 1660
rect 8908 80 8948 2416
rect 9004 1952 9044 1961
rect 9004 1817 9044 1912
rect 9100 1868 9140 7876
rect 9196 7244 9236 9472
rect 9196 6488 9236 7204
rect 9196 6439 9236 6448
rect 9388 6068 9428 6077
rect 9388 5564 9428 6028
rect 9388 5515 9428 5524
rect 9484 5564 9524 14596
rect 9580 6236 9620 20812
rect 9676 20348 9716 20357
rect 9676 19256 9716 20308
rect 9676 19207 9716 19216
rect 9676 19088 9716 19097
rect 9676 18668 9716 19048
rect 9676 18619 9716 18628
rect 9772 12980 9812 22912
rect 9868 16988 9908 32992
rect 9964 32276 10004 36604
rect 9964 32227 10004 32236
rect 10060 34460 10100 34469
rect 10060 33704 10100 34420
rect 10060 32192 10100 33664
rect 10156 33452 10196 39544
rect 10252 34376 10292 39796
rect 10348 39752 10388 39761
rect 10348 37652 10388 39712
rect 10348 37603 10388 37612
rect 10444 38744 10484 38753
rect 10348 37316 10388 37325
rect 10348 35132 10388 37276
rect 10444 36644 10484 38704
rect 10540 38156 10580 44080
rect 10636 42020 10676 44920
rect 10732 44120 10772 47608
rect 10828 47396 10868 47405
rect 10828 46472 10868 47356
rect 10828 46423 10868 46432
rect 10828 46304 10868 46313
rect 10828 45044 10868 46264
rect 10828 44995 10868 45004
rect 10732 44071 10772 44080
rect 10828 44708 10868 44717
rect 10732 43532 10772 43541
rect 10732 42188 10772 43492
rect 10732 42139 10772 42148
rect 10636 41971 10676 41980
rect 10828 41516 10868 44668
rect 10828 41467 10868 41476
rect 10924 41432 10964 49708
rect 11116 49664 11156 50464
rect 11212 49748 11252 58276
rect 11308 57812 11348 57821
rect 11308 57560 11348 57772
rect 11308 57511 11348 57520
rect 11308 54788 11348 54797
rect 11308 54284 11348 54748
rect 11308 54235 11348 54244
rect 11404 53300 11444 66844
rect 11500 66968 11540 66977
rect 11500 66833 11540 66928
rect 11500 65960 11540 65969
rect 11500 64364 11540 65920
rect 11500 64315 11540 64324
rect 11500 63860 11540 63869
rect 11500 63188 11540 63820
rect 11500 63139 11540 63148
rect 11500 62180 11540 62189
rect 11500 61508 11540 62140
rect 11500 58652 11540 61468
rect 11596 61088 11636 71968
rect 11692 66884 11732 79780
rect 11788 79736 11828 79745
rect 11788 79601 11828 79696
rect 11788 79232 11828 79241
rect 11788 78980 11828 79192
rect 11788 77468 11828 78940
rect 11788 77419 11828 77428
rect 11884 78308 11924 81796
rect 11980 80492 12020 80501
rect 11980 79988 12020 80452
rect 11980 79939 12020 79948
rect 11980 79820 12020 79829
rect 11980 79736 12020 79780
rect 11980 78476 12020 79696
rect 11980 78427 12020 78436
rect 11884 75200 11924 78268
rect 11884 73940 11924 75160
rect 11884 73891 11924 73900
rect 11980 78308 12020 78317
rect 11884 73436 11924 73445
rect 11788 71336 11828 71345
rect 11788 69404 11828 71296
rect 11788 69355 11828 69364
rect 11692 66835 11732 66844
rect 11788 69236 11828 69245
rect 11788 68396 11828 69196
rect 11788 66716 11828 68356
rect 11884 67976 11924 73396
rect 11980 73184 12020 78268
rect 12076 73604 12116 83308
rect 12172 80324 12212 86500
rect 12268 83684 12308 93724
rect 12556 89312 12596 89321
rect 12556 89228 12596 89272
rect 12556 89177 12596 89188
rect 12556 88052 12596 88061
rect 12364 87548 12404 87557
rect 12364 86792 12404 87508
rect 12364 86743 12404 86752
rect 12556 86372 12596 88012
rect 12556 86323 12596 86332
rect 12460 86204 12500 86213
rect 12460 86069 12500 86164
rect 12556 86120 12596 86129
rect 12556 86036 12596 86080
rect 12556 85985 12596 85996
rect 12364 85868 12404 85963
rect 12364 85819 12404 85828
rect 12556 85616 12596 85625
rect 12364 85448 12404 85457
rect 12364 85112 12404 85408
rect 12364 84524 12404 85072
rect 12460 85028 12500 85039
rect 12460 84944 12500 84988
rect 12460 84895 12500 84904
rect 12364 84475 12404 84484
rect 12460 84776 12500 84785
rect 12268 83635 12308 83644
rect 12268 83432 12308 83441
rect 12268 82844 12308 83392
rect 12268 82004 12308 82804
rect 12364 82004 12404 82013
rect 12268 81964 12364 82004
rect 12364 81332 12404 81964
rect 12268 80492 12308 80501
rect 12268 80408 12308 80452
rect 12268 80357 12308 80368
rect 12172 79232 12212 80284
rect 12364 80324 12404 81292
rect 12364 80275 12404 80284
rect 12460 80156 12500 84736
rect 12556 84356 12596 85576
rect 12556 84221 12596 84316
rect 12556 83936 12596 83945
rect 12556 83600 12596 83896
rect 12556 83551 12596 83560
rect 12556 82592 12596 82601
rect 12556 82004 12596 82552
rect 12556 81955 12596 81964
rect 12172 79183 12212 79192
rect 12268 80116 12500 80156
rect 12172 78812 12212 78907
rect 12172 78763 12212 78772
rect 12172 77468 12212 77563
rect 12172 77419 12212 77428
rect 12172 77300 12212 77309
rect 12172 75956 12212 77260
rect 12172 75907 12212 75916
rect 12076 73555 12116 73564
rect 12172 75032 12212 75041
rect 11980 73135 12020 73144
rect 12076 73436 12116 73445
rect 11980 72932 12020 72941
rect 11980 72344 12020 72892
rect 11980 71336 12020 72304
rect 12076 72008 12116 73396
rect 12172 72932 12212 74992
rect 12172 72883 12212 72892
rect 12076 71959 12116 71968
rect 11980 71287 12020 71296
rect 12076 71840 12116 71849
rect 12076 71420 12116 71800
rect 11884 67927 11924 67936
rect 11980 70916 12020 70925
rect 11692 66676 11828 66716
rect 11692 65456 11732 66676
rect 11884 66632 11924 66641
rect 11692 65120 11732 65416
rect 11692 65071 11732 65080
rect 11788 66212 11828 66221
rect 11692 64028 11732 64037
rect 11692 63188 11732 63988
rect 11788 63776 11828 66172
rect 11788 63727 11828 63736
rect 11692 63139 11732 63148
rect 11788 63608 11828 63617
rect 11692 62936 11732 62945
rect 11692 62348 11732 62896
rect 11692 62299 11732 62308
rect 11596 61048 11732 61088
rect 11500 58603 11540 58612
rect 11596 60920 11636 60929
rect 11500 58400 11540 58409
rect 11500 53864 11540 58360
rect 11500 53815 11540 53824
rect 11404 53260 11540 53300
rect 11308 51848 11348 51857
rect 11308 50084 11348 51808
rect 11404 50336 11444 50345
rect 11404 50201 11444 50296
rect 11308 49949 11348 50044
rect 11212 49708 11444 49748
rect 11116 49615 11156 49624
rect 11212 49580 11252 49589
rect 11212 48992 11252 49540
rect 11212 48943 11252 48952
rect 11308 49496 11348 49505
rect 11308 47984 11348 49456
rect 11308 47935 11348 47944
rect 11212 46976 11252 46985
rect 11116 46556 11156 46565
rect 11020 43532 11060 43541
rect 11020 43397 11060 43492
rect 11116 43196 11156 46516
rect 11212 45212 11252 46936
rect 11212 45163 11252 45172
rect 11308 46556 11348 46565
rect 11308 45044 11348 46516
rect 11212 45004 11348 45044
rect 11212 44792 11252 45004
rect 11212 44743 11252 44752
rect 11308 44624 11348 44633
rect 11308 44288 11348 44584
rect 11308 43220 11348 44248
rect 11404 43532 11444 49708
rect 11500 47648 11540 53260
rect 11596 50420 11636 60880
rect 11692 58904 11732 61048
rect 11788 59660 11828 63568
rect 11788 59611 11828 59620
rect 11692 51092 11732 58864
rect 11788 59492 11828 59501
rect 11788 58064 11828 59452
rect 11788 58015 11828 58024
rect 11884 57896 11924 66592
rect 11980 65456 12020 70876
rect 12076 70832 12116 71380
rect 12076 70783 12116 70792
rect 12172 71588 12212 71597
rect 12172 70748 12212 71548
rect 12172 70699 12212 70708
rect 12076 69992 12116 70001
rect 12076 66212 12116 69952
rect 12172 67724 12212 67733
rect 12172 66380 12212 67684
rect 12172 66331 12212 66340
rect 12076 66163 12116 66172
rect 12172 66212 12212 66221
rect 11980 65416 12116 65456
rect 11980 65204 12020 65213
rect 11980 63860 12020 65164
rect 12076 64784 12116 65416
rect 12076 64735 12116 64744
rect 12076 64616 12116 64625
rect 12076 64028 12116 64576
rect 12076 63979 12116 63988
rect 11980 63811 12020 63820
rect 12076 63692 12116 63701
rect 12076 63557 12116 63652
rect 12172 63380 12212 66172
rect 11788 57856 11924 57896
rect 11980 63340 12212 63380
rect 12268 63944 12308 80116
rect 12364 79904 12404 79913
rect 12364 78308 12404 79864
rect 12556 79736 12596 79745
rect 12556 79064 12596 79696
rect 12556 79015 12596 79024
rect 12364 78259 12404 78268
rect 12460 78812 12500 78821
rect 12364 78140 12404 78149
rect 12364 78005 12404 78100
rect 12364 77216 12404 77225
rect 12364 76376 12404 77176
rect 12364 76327 12404 76336
rect 11788 57812 11828 57856
rect 11788 57140 11828 57772
rect 11788 55040 11828 57100
rect 11788 54788 11828 55000
rect 11788 54200 11828 54748
rect 11788 54151 11828 54160
rect 11884 57728 11924 57737
rect 11692 51043 11732 51052
rect 11788 53444 11828 53453
rect 11596 50371 11636 50380
rect 11692 50504 11732 50515
rect 11692 50420 11732 50464
rect 11692 50371 11732 50380
rect 11788 48236 11828 53404
rect 11884 51764 11924 57688
rect 11980 53300 12020 63340
rect 12268 63272 12308 63904
rect 12076 63232 12308 63272
rect 12364 76208 12404 76217
rect 12076 59072 12116 63232
rect 12172 63104 12212 63115
rect 12172 63020 12212 63064
rect 12172 62348 12212 62980
rect 12172 61676 12212 62308
rect 12268 62516 12308 62525
rect 12268 61844 12308 62476
rect 12268 61795 12308 61804
rect 12172 61627 12212 61636
rect 12172 61424 12212 61433
rect 12172 60836 12212 61384
rect 12172 60080 12212 60796
rect 12268 60248 12308 60257
rect 12268 60113 12308 60208
rect 12172 60031 12212 60040
rect 12172 59912 12212 59921
rect 12172 59408 12212 59872
rect 12172 59359 12212 59368
rect 12268 59240 12308 59335
rect 12268 59191 12308 59200
rect 12076 59032 12308 59072
rect 12076 58904 12116 58913
rect 12076 58232 12116 58864
rect 12172 58736 12212 58745
rect 12172 58601 12212 58696
rect 12172 58484 12212 58493
rect 12172 58349 12212 58444
rect 12076 58183 12116 58192
rect 12172 58232 12212 58241
rect 12076 57980 12116 57989
rect 12076 57728 12116 57940
rect 12076 57679 12116 57688
rect 12076 57560 12116 57569
rect 12076 57425 12116 57520
rect 12172 56636 12212 58192
rect 12172 56587 12212 56596
rect 12076 56300 12116 56309
rect 12076 55628 12116 56260
rect 12076 55579 12116 55588
rect 12268 56216 12308 59032
rect 12268 55544 12308 56176
rect 12268 55495 12308 55504
rect 12172 54956 12212 54965
rect 11980 53260 12116 53300
rect 11884 51715 11924 51724
rect 11788 48187 11828 48196
rect 11884 51008 11924 51017
rect 11884 50084 11924 50968
rect 11500 47608 11636 47648
rect 11596 47396 11636 47608
rect 11596 47356 11732 47396
rect 11500 47312 11540 47321
rect 11500 46556 11540 47272
rect 11500 46507 11540 46516
rect 11596 47228 11636 47237
rect 11500 46388 11540 46397
rect 11500 46136 11540 46348
rect 11500 46087 11540 46096
rect 11596 45716 11636 47188
rect 11692 46808 11732 47356
rect 11692 46759 11732 46768
rect 11500 45632 11540 45641
rect 11500 44960 11540 45592
rect 11500 44624 11540 44920
rect 11500 44575 11540 44584
rect 11404 43483 11444 43492
rect 11500 43448 11540 43457
rect 11116 42104 11156 43156
rect 11212 43180 11348 43220
rect 11404 43364 11444 43373
rect 11212 42692 11252 43180
rect 11212 42643 11252 42652
rect 11116 42055 11156 42064
rect 11212 42440 11252 42449
rect 10924 41392 11156 41432
rect 10636 41180 10676 41189
rect 10636 39500 10676 41140
rect 11020 41180 11060 41189
rect 10636 39451 10676 39460
rect 10732 41096 10772 41105
rect 10732 41012 10772 41056
rect 10540 38107 10580 38116
rect 10636 38912 10676 38921
rect 10540 37988 10580 37997
rect 10540 37820 10580 37948
rect 10540 37484 10580 37780
rect 10540 37435 10580 37444
rect 10444 36595 10484 36604
rect 10348 34544 10388 35092
rect 10540 36224 10580 36233
rect 10540 35048 10580 36184
rect 10540 34999 10580 35008
rect 10348 34495 10388 34504
rect 10252 33620 10292 34336
rect 10444 34460 10484 34469
rect 10444 33788 10484 34420
rect 10444 33739 10484 33748
rect 10292 33580 10484 33620
rect 10252 33571 10292 33580
rect 10156 33412 10292 33452
rect 9964 32024 10004 32033
rect 9964 31604 10004 31984
rect 9964 31555 10004 31564
rect 9964 31436 10004 31445
rect 9964 28412 10004 31396
rect 10060 29840 10100 32152
rect 10060 29791 10100 29800
rect 10156 33284 10196 33293
rect 10060 28916 10100 28925
rect 10060 28781 10100 28876
rect 10156 28580 10196 33244
rect 10252 31184 10292 33412
rect 10252 31135 10292 31144
rect 10348 32696 10388 32705
rect 10156 28531 10196 28540
rect 10252 30092 10292 30101
rect 9964 28363 10004 28372
rect 10060 28328 10100 28337
rect 10060 28193 10100 28288
rect 10156 28160 10196 28169
rect 9964 28076 10004 28085
rect 9964 27404 10004 28036
rect 10060 27992 10100 28001
rect 10060 27857 10100 27952
rect 9964 27355 10004 27364
rect 10060 27236 10100 27245
rect 9964 26900 10004 26909
rect 9964 26228 10004 26860
rect 10060 26900 10100 27196
rect 10060 26851 10100 26860
rect 10060 26564 10100 26573
rect 10060 26429 10100 26524
rect 9964 26179 10004 26188
rect 10060 26144 10100 26153
rect 9964 26060 10004 26069
rect 9964 25556 10004 26020
rect 10060 26009 10100 26104
rect 10060 25808 10100 25817
rect 10060 25673 10100 25768
rect 9964 25507 10004 25516
rect 9964 25304 10004 25313
rect 9964 23624 10004 25264
rect 9964 23575 10004 23584
rect 10156 23372 10196 28120
rect 10252 23792 10292 30052
rect 10348 30008 10388 32656
rect 10444 32108 10484 33580
rect 10540 32528 10580 32537
rect 10540 32276 10580 32488
rect 10540 32227 10580 32236
rect 10444 32024 10484 32068
rect 10444 31944 10484 31984
rect 10444 31772 10484 31781
rect 10444 30092 10484 31732
rect 10444 30043 10484 30052
rect 10540 31520 10580 31529
rect 10348 29959 10388 29968
rect 10444 29924 10484 29933
rect 10444 29789 10484 29884
rect 10348 29168 10388 29177
rect 10348 28832 10388 29128
rect 10444 29084 10484 29093
rect 10444 28916 10484 29044
rect 10444 28867 10484 28876
rect 10348 28783 10388 28792
rect 10252 23743 10292 23752
rect 10348 28664 10388 28673
rect 10348 26060 10388 28624
rect 10348 25388 10388 26020
rect 10156 23323 10196 23332
rect 10252 23624 10292 23633
rect 10060 23288 10100 23297
rect 9964 22868 10004 22877
rect 9964 22448 10004 22828
rect 9964 22399 10004 22408
rect 9964 20180 10004 20189
rect 9964 17660 10004 20140
rect 10060 19340 10100 23248
rect 10156 22196 10196 22205
rect 10156 21524 10196 22156
rect 10156 21475 10196 21484
rect 10060 19291 10100 19300
rect 10156 20852 10196 20861
rect 10156 19844 10196 20812
rect 10156 18500 10196 19804
rect 10252 19508 10292 23584
rect 10348 23288 10388 25348
rect 10348 23239 10388 23248
rect 10444 27488 10484 27497
rect 10444 23876 10484 27448
rect 10540 25556 10580 31480
rect 10636 30680 10676 38872
rect 10636 30092 10676 30640
rect 10636 30043 10676 30052
rect 10636 29924 10676 29935
rect 10636 29840 10676 29884
rect 10636 29791 10676 29800
rect 10636 29168 10676 29177
rect 10636 28748 10676 29128
rect 10636 28699 10676 28708
rect 10636 28496 10676 28505
rect 10636 27824 10676 28456
rect 10636 26816 10676 27784
rect 10636 26767 10676 26776
rect 10540 25507 10580 25516
rect 10636 25892 10676 25901
rect 10348 23036 10388 23045
rect 10348 22532 10388 22996
rect 10348 22483 10388 22492
rect 10348 21524 10388 21533
rect 10348 21389 10388 21484
rect 10348 21272 10388 21281
rect 10348 20180 10388 21232
rect 10348 20131 10388 20140
rect 10444 19676 10484 23836
rect 10636 24548 10676 25852
rect 10444 19627 10484 19636
rect 10540 20852 10580 20861
rect 10252 19459 10292 19468
rect 9964 17611 10004 17620
rect 10060 18460 10196 18500
rect 10444 19424 10484 19433
rect 9868 16853 9908 16948
rect 9964 16904 10004 16913
rect 9868 15224 9908 15233
rect 9868 14804 9908 15184
rect 9868 14755 9908 14764
rect 9676 12940 9812 12980
rect 9676 8252 9716 12940
rect 9772 12620 9812 12629
rect 9772 12536 9812 12580
rect 9772 12485 9812 12496
rect 9868 12452 9908 12461
rect 9676 8203 9716 8212
rect 9772 11780 9812 11789
rect 9772 7244 9812 11740
rect 9868 11276 9908 12412
rect 9868 10856 9908 11236
rect 9868 10807 9908 10816
rect 9868 9680 9908 9689
rect 9868 9512 9908 9640
rect 9868 9463 9908 9472
rect 9772 6404 9812 7204
rect 9868 9344 9908 9353
rect 9868 7076 9908 9304
rect 9964 7916 10004 16864
rect 10060 12980 10100 18460
rect 10156 18164 10196 18173
rect 10156 17744 10196 18124
rect 10156 17695 10196 17704
rect 10348 17576 10388 17585
rect 10252 16820 10292 16829
rect 10156 14636 10196 14645
rect 10156 14048 10196 14596
rect 10156 13999 10196 14008
rect 10060 12940 10196 12980
rect 10060 12284 10100 12293
rect 10060 11864 10100 12244
rect 10060 11815 10100 11824
rect 10060 10184 10100 10193
rect 10060 9428 10100 10144
rect 10060 9293 10100 9388
rect 10156 9344 10196 12940
rect 10252 10772 10292 16780
rect 10348 15728 10388 17536
rect 10348 14720 10388 15688
rect 10444 15476 10484 19384
rect 10540 15560 10580 20812
rect 10636 18500 10676 24508
rect 10732 23060 10772 40972
rect 10924 41096 10964 41105
rect 10924 40961 10964 41056
rect 10828 40508 10868 40517
rect 10828 39668 10868 40468
rect 11020 39836 11060 41140
rect 10828 38912 10868 39628
rect 10924 39752 10964 39761
rect 10924 39617 10964 39712
rect 11020 39584 11060 39796
rect 11020 39535 11060 39544
rect 10924 39332 10964 39341
rect 10924 38996 10964 39292
rect 11116 39080 11156 41392
rect 11116 39031 11156 39040
rect 10924 38947 10964 38956
rect 10828 38863 10868 38872
rect 11116 38912 11156 38921
rect 11020 38828 11060 38837
rect 11020 38660 11060 38788
rect 11116 38777 11156 38872
rect 11020 38620 11156 38660
rect 11020 38156 11060 38165
rect 10828 38072 10868 38081
rect 10828 33872 10868 38032
rect 10924 36644 10964 36653
rect 10924 36224 10964 36604
rect 10924 36175 10964 36184
rect 10924 35720 10964 35729
rect 10924 34460 10964 35680
rect 10924 34411 10964 34420
rect 10828 33832 10964 33872
rect 10924 33788 10964 33832
rect 10924 33739 10964 33748
rect 10828 33704 10868 33713
rect 10828 32108 10868 33664
rect 10924 33620 10964 33629
rect 10924 33116 10964 33580
rect 10924 33067 10964 33076
rect 10828 31973 10868 32068
rect 10924 32948 10964 32957
rect 10828 30848 10868 30857
rect 10828 30713 10868 30808
rect 10924 30092 10964 32908
rect 10828 30052 10964 30092
rect 10828 29168 10868 30052
rect 10828 29119 10868 29128
rect 10924 29924 10964 29933
rect 10924 29084 10964 29884
rect 10924 29035 10964 29044
rect 10828 29000 10868 29009
rect 10828 27740 10868 28960
rect 10828 27691 10868 27700
rect 10924 28916 10964 28925
rect 10828 27572 10868 27581
rect 10828 27068 10868 27532
rect 10828 26480 10868 27028
rect 10828 26431 10868 26440
rect 10828 23624 10868 23633
rect 10828 23288 10868 23584
rect 10828 23239 10868 23248
rect 10732 23020 10868 23060
rect 10732 21188 10772 21197
rect 10732 20516 10772 21148
rect 10732 20467 10772 20476
rect 10636 18451 10676 18460
rect 10732 20264 10772 20273
rect 10636 17828 10676 17837
rect 10636 16484 10676 17788
rect 10732 17156 10772 20224
rect 10732 17107 10772 17116
rect 10636 16435 10676 16444
rect 10732 16988 10772 16997
rect 10636 16316 10676 16325
rect 10636 16148 10676 16276
rect 10636 15980 10676 16108
rect 10636 15931 10676 15940
rect 10732 15728 10772 16948
rect 10732 15679 10772 15688
rect 10540 15520 10772 15560
rect 10444 15436 10580 15476
rect 10348 14132 10388 14680
rect 10348 14083 10388 14092
rect 10444 14552 10484 14561
rect 10444 13964 10484 14512
rect 10348 13924 10484 13964
rect 10348 11696 10388 13924
rect 10348 11647 10388 11656
rect 10444 13208 10484 13217
rect 10252 10723 10292 10732
rect 10348 11528 10388 11537
rect 10252 9764 10292 9773
rect 10252 9512 10292 9724
rect 10252 9463 10292 9472
rect 10156 9260 10196 9304
rect 10156 9211 10196 9220
rect 10252 9260 10292 9269
rect 10060 8924 10100 8933
rect 10060 8789 10100 8884
rect 10252 8504 10292 9220
rect 10252 8455 10292 8464
rect 9964 7867 10004 7876
rect 9868 6488 9908 7036
rect 9868 6439 9908 6448
rect 9772 6355 9812 6364
rect 9964 6404 10004 6413
rect 9868 6236 9908 6245
rect 9580 6196 9812 6236
rect 9484 5515 9524 5524
rect 9676 6068 9716 6077
rect 9196 2708 9236 2719
rect 9196 2624 9236 2668
rect 9196 2575 9236 2584
rect 9676 2624 9716 6028
rect 9772 2900 9812 6196
rect 9868 4724 9908 6196
rect 9964 6068 10004 6364
rect 10156 6236 10196 6245
rect 9964 6019 10004 6028
rect 10060 6152 10100 6161
rect 10060 6017 10100 6112
rect 10156 5648 10196 6196
rect 10156 5599 10196 5608
rect 10156 5480 10196 5489
rect 10060 5228 10100 5237
rect 10060 5093 10100 5188
rect 10156 5060 10196 5440
rect 10156 5011 10196 5020
rect 10252 4808 10292 4817
rect 10348 4808 10388 11488
rect 10444 6068 10484 13168
rect 10444 6019 10484 6028
rect 10540 8756 10580 15436
rect 10636 15392 10676 15401
rect 10636 14636 10676 15352
rect 10636 14587 10676 14596
rect 10540 6404 10580 8716
rect 10540 5816 10580 6364
rect 10540 5767 10580 5776
rect 10636 13376 10676 13385
rect 10292 4768 10388 4808
rect 10252 4759 10292 4768
rect 9868 4675 9908 4684
rect 10636 4556 10676 13336
rect 10732 12980 10772 15520
rect 10828 13292 10868 23020
rect 10924 20684 10964 28876
rect 11020 27656 11060 38116
rect 11116 35972 11156 38620
rect 11116 35923 11156 35932
rect 11020 27607 11060 27616
rect 11116 34544 11156 34553
rect 11020 27404 11060 27413
rect 11020 25136 11060 27364
rect 11020 24548 11060 25096
rect 11020 24499 11060 24508
rect 11020 21356 11060 21365
rect 11020 20852 11060 21316
rect 11020 20803 11060 20812
rect 10924 20635 10964 20644
rect 11020 20348 11060 20357
rect 10924 20096 10964 20105
rect 10924 19961 10964 20056
rect 10828 13243 10868 13252
rect 10924 18500 10964 18509
rect 10732 12940 10868 12980
rect 10732 11528 10772 11537
rect 10732 10268 10772 11488
rect 10828 11024 10868 12940
rect 10828 10975 10868 10984
rect 10732 10219 10772 10228
rect 10828 10856 10868 10865
rect 10732 10100 10772 10109
rect 10732 9764 10772 10060
rect 10732 9715 10772 9724
rect 10732 7076 10772 7085
rect 10732 6488 10772 7036
rect 10732 6439 10772 6448
rect 10732 5732 10772 5741
rect 10732 5144 10772 5692
rect 10732 5095 10772 5104
rect 10636 4220 10676 4516
rect 10636 4171 10676 4180
rect 10828 4136 10868 10816
rect 10924 8840 10964 18460
rect 11020 17744 11060 20308
rect 11116 20264 11156 34504
rect 11212 33452 11252 42400
rect 11212 33403 11252 33412
rect 11308 41264 11348 41273
rect 11212 33284 11252 33293
rect 11212 32948 11252 33244
rect 11212 30512 11252 32908
rect 11308 31772 11348 41224
rect 11404 35384 11444 43324
rect 11500 43112 11540 43408
rect 11500 43063 11540 43072
rect 11596 42692 11636 45676
rect 11596 42643 11636 42652
rect 11692 46304 11732 46313
rect 11596 41936 11636 41945
rect 11500 41852 11540 41861
rect 11500 41180 11540 41812
rect 11500 41131 11540 41140
rect 11596 41096 11636 41896
rect 11596 41047 11636 41056
rect 11596 40172 11636 40181
rect 11500 39836 11540 39845
rect 11500 39416 11540 39796
rect 11500 39367 11540 39376
rect 11596 38492 11636 40132
rect 11596 38072 11636 38452
rect 11596 38023 11636 38032
rect 11500 37904 11540 37913
rect 11500 37769 11540 37864
rect 11692 37904 11732 46264
rect 11788 45800 11828 45809
rect 11788 44288 11828 45760
rect 11788 43280 11828 44248
rect 11788 43231 11828 43240
rect 11692 37855 11732 37864
rect 11788 42104 11828 42113
rect 11596 37820 11636 37829
rect 11500 37484 11540 37493
rect 11500 36476 11540 37444
rect 11500 36427 11540 36436
rect 11404 35335 11444 35344
rect 11500 36056 11540 36065
rect 11500 35216 11540 36016
rect 11404 35176 11540 35216
rect 11404 32528 11444 35176
rect 11404 32479 11444 32488
rect 11500 35048 11540 35057
rect 11500 32276 11540 35008
rect 11596 34544 11636 37780
rect 11692 37484 11732 37493
rect 11692 36644 11732 37444
rect 11788 36896 11828 42064
rect 11884 39164 11924 50044
rect 11980 50840 12020 50849
rect 11980 48824 12020 50800
rect 11980 48775 12020 48784
rect 12076 46976 12116 53260
rect 12172 51680 12212 54916
rect 12172 51631 12212 51640
rect 12268 50336 12308 50345
rect 12268 50201 12308 50296
rect 11980 46936 12116 46976
rect 12172 48824 12212 48833
rect 11980 42944 12020 46936
rect 11980 42895 12020 42904
rect 12076 46808 12116 46817
rect 11980 40928 12020 40937
rect 11980 40256 12020 40888
rect 11980 40207 12020 40216
rect 11980 40004 12020 40013
rect 11980 39869 12020 39964
rect 11884 39124 12020 39164
rect 11884 38996 11924 39005
rect 11884 38156 11924 38956
rect 11884 37568 11924 38116
rect 11884 37519 11924 37528
rect 11788 36847 11828 36856
rect 11692 36595 11732 36604
rect 11788 36728 11828 36737
rect 11788 36593 11828 36688
rect 11884 36644 11924 36653
rect 11596 34495 11636 34504
rect 11692 36476 11732 36485
rect 11692 34376 11732 36436
rect 11308 31723 11348 31732
rect 11404 32236 11540 32276
rect 11596 34336 11732 34376
rect 11788 35972 11828 35981
rect 11404 31436 11444 32236
rect 11500 32108 11540 32117
rect 11500 31604 11540 32068
rect 11500 31555 11540 31564
rect 11404 31396 11540 31436
rect 11212 30472 11444 30512
rect 11212 29924 11252 29933
rect 11212 27824 11252 29884
rect 11308 29420 11348 29431
rect 11308 29336 11348 29380
rect 11308 29287 11348 29296
rect 11308 29084 11348 29093
rect 11308 28580 11348 29044
rect 11308 28531 11348 28540
rect 11212 27775 11252 27784
rect 11308 28328 11348 28337
rect 11404 28328 11444 30472
rect 11348 28288 11444 28328
rect 11212 27656 11252 27665
rect 11212 22196 11252 27616
rect 11308 27572 11348 28288
rect 11500 27572 11540 31396
rect 11308 27523 11348 27532
rect 11404 27532 11540 27572
rect 11596 28412 11636 34336
rect 11692 33368 11732 33377
rect 11692 32948 11732 33328
rect 11692 32780 11732 32908
rect 11692 32731 11732 32740
rect 11692 32360 11732 32369
rect 11692 29336 11732 32320
rect 11788 30344 11828 35932
rect 11788 30295 11828 30304
rect 11884 32192 11924 36604
rect 11980 36140 12020 39124
rect 12076 36476 12116 46768
rect 12172 43616 12212 48784
rect 12268 48740 12308 48751
rect 12268 48656 12308 48700
rect 12268 48607 12308 48616
rect 12268 47228 12308 47237
rect 12268 46304 12308 47188
rect 12268 46255 12308 46264
rect 12172 43567 12212 43576
rect 12268 46136 12308 46145
rect 12268 43220 12308 46096
rect 12364 46052 12404 76168
rect 12460 75872 12500 78772
rect 12460 75823 12500 75832
rect 12556 78308 12596 78317
rect 12460 74864 12500 74873
rect 12460 73688 12500 74824
rect 12556 73940 12596 78268
rect 12556 73891 12596 73900
rect 12460 73639 12500 73648
rect 12652 73460 12692 93892
rect 12940 93932 12980 93941
rect 12940 93797 12980 93892
rect 13036 93764 13076 94648
rect 13228 94637 13268 94732
rect 13324 94184 13364 96688
rect 13516 95108 13556 96688
rect 13516 95059 13556 95068
rect 13324 94135 13364 94144
rect 13420 94520 13460 94529
rect 13420 94016 13460 94480
rect 13708 94268 13748 96688
rect 13900 94604 13940 96688
rect 13900 94555 13940 94564
rect 13708 94219 13748 94228
rect 14092 94184 14132 96688
rect 14284 95948 14324 96688
rect 14284 95899 14324 95908
rect 14380 94772 14420 94781
rect 14380 94637 14420 94732
rect 14476 94268 14516 96688
rect 14668 96620 14708 96688
rect 14668 96571 14708 96580
rect 14476 94219 14516 94228
rect 14572 94688 14612 94697
rect 14092 94135 14132 94144
rect 13420 93967 13460 93976
rect 13900 93932 13940 93941
rect 13900 93797 13940 93892
rect 14284 93932 14324 93941
rect 14284 93797 14324 93892
rect 14476 93848 14516 93857
rect 13036 93715 13076 93724
rect 13612 92756 13652 92765
rect 13132 90404 13172 90413
rect 13036 90152 13076 90161
rect 13036 89648 13076 90112
rect 13036 89599 13076 89608
rect 12748 89564 12788 89573
rect 12748 88304 12788 89524
rect 12748 87884 12788 88264
rect 12844 89480 12884 89489
rect 12844 89144 12884 89440
rect 12844 88892 12884 89104
rect 13132 89312 13172 90364
rect 13132 89060 13172 89272
rect 13228 89732 13268 89741
rect 13228 89228 13268 89692
rect 13228 89179 13268 89188
rect 13516 89648 13556 89657
rect 13132 89011 13172 89020
rect 12844 87968 12884 88852
rect 13516 88892 13556 89608
rect 13132 88808 13172 88817
rect 13132 88556 13172 88768
rect 13132 88220 13172 88516
rect 13132 88171 13172 88180
rect 13516 88556 13556 88852
rect 13516 88136 13556 88516
rect 12844 87919 12884 87928
rect 13132 88052 13172 88063
rect 13132 87968 13172 88012
rect 13132 87919 13172 87928
rect 12748 87835 12788 87844
rect 12844 87800 12884 87809
rect 12844 87632 12884 87760
rect 12940 87632 12980 87641
rect 12844 87592 12940 87632
rect 12940 87583 12980 87592
rect 13036 87548 13076 87557
rect 12940 87380 12980 87389
rect 12940 86624 12980 87340
rect 13036 86708 13076 87508
rect 13324 87548 13364 87557
rect 13036 86659 13076 86668
rect 13132 87464 13172 87473
rect 12940 86575 12980 86584
rect 13036 86456 13076 86465
rect 13036 86321 13076 86416
rect 12844 86204 12884 86215
rect 12844 86120 12884 86164
rect 12844 86071 12884 86080
rect 12748 85952 12788 85961
rect 12748 85448 12788 85912
rect 13036 85784 13076 85793
rect 12748 85399 12788 85408
rect 12844 85616 12884 85625
rect 12748 85280 12788 85289
rect 12748 85112 12788 85240
rect 12748 83768 12788 85072
rect 12748 83540 12788 83728
rect 12844 83684 12884 85576
rect 12940 85028 12980 85123
rect 12940 84979 12980 84988
rect 12940 84860 12980 84869
rect 12940 84440 12980 84820
rect 12940 84391 12980 84400
rect 13036 84272 13076 85744
rect 13132 85364 13172 87424
rect 13324 87380 13364 87508
rect 13324 87331 13364 87340
rect 13324 87212 13364 87221
rect 13228 87128 13268 87137
rect 13228 86624 13268 87088
rect 13228 86575 13268 86584
rect 13228 86456 13268 86465
rect 13228 86120 13268 86416
rect 13228 86071 13268 86080
rect 13132 85324 13268 85364
rect 13132 85196 13172 85205
rect 13132 84356 13172 85156
rect 13132 84307 13172 84316
rect 13036 84223 13076 84232
rect 13228 84020 13268 85324
rect 13228 83971 13268 83980
rect 12844 83635 12884 83644
rect 13228 83600 13268 83609
rect 12748 83500 12884 83540
rect 12748 82844 12788 82853
rect 12844 82844 12884 83500
rect 12844 82804 13172 82844
rect 12748 82709 12788 82804
rect 13036 82676 13076 82685
rect 13036 82256 13076 82636
rect 13036 82207 13076 82216
rect 13036 82004 13076 82013
rect 12748 80576 12788 80585
rect 12748 80441 12788 80536
rect 13036 80492 13076 81964
rect 13036 80443 13076 80452
rect 12748 80324 12788 80333
rect 12748 79904 12788 80284
rect 12748 79855 12788 79864
rect 12844 79904 12884 79913
rect 12748 79652 12788 79661
rect 12748 79064 12788 79612
rect 12844 79232 12884 79864
rect 12940 79736 12980 79745
rect 12940 79601 12980 79696
rect 12844 79183 12884 79192
rect 13036 79316 13076 79325
rect 12748 79015 12788 79024
rect 12940 79064 12980 79073
rect 12748 78812 12788 78821
rect 12748 78308 12788 78772
rect 12940 78476 12980 79024
rect 13036 78728 13076 79276
rect 13036 78679 13076 78688
rect 12940 78427 12980 78436
rect 13036 78560 13076 78569
rect 12748 78268 12884 78308
rect 12844 77888 12884 78268
rect 12748 77552 12788 77561
rect 12748 75200 12788 77512
rect 12844 76460 12884 77848
rect 12940 77384 12980 77393
rect 12940 76796 12980 77344
rect 12940 76747 12980 76756
rect 12844 76411 12884 76420
rect 12844 76124 12884 76133
rect 13036 76124 13076 78520
rect 13132 76292 13172 82804
rect 13228 80156 13268 83560
rect 13324 81752 13364 87172
rect 13516 85868 13556 88096
rect 13612 86540 13652 92716
rect 14476 90740 14516 93808
rect 14572 93680 14612 94648
rect 14764 94688 14804 94697
rect 14668 93932 14708 93941
rect 14668 93797 14708 93892
rect 14572 93631 14612 93640
rect 14476 90691 14516 90700
rect 14188 90488 14228 90497
rect 13612 85952 13652 86500
rect 13612 85903 13652 85912
rect 13708 89564 13748 89573
rect 13708 88724 13748 89524
rect 13420 85828 13556 85868
rect 13420 84860 13460 85828
rect 13612 85784 13652 85793
rect 13612 84860 13652 85744
rect 13708 85280 13748 88684
rect 13708 85231 13748 85240
rect 13804 89480 13844 89489
rect 13804 88640 13844 89440
rect 13420 84820 13556 84860
rect 13324 81703 13364 81712
rect 13420 83852 13460 83861
rect 13228 80107 13268 80116
rect 13324 80576 13364 80585
rect 13324 80492 13364 80536
rect 13324 79820 13364 80452
rect 13324 79771 13364 79780
rect 13228 79736 13268 79745
rect 13228 78980 13268 79696
rect 13228 78931 13268 78940
rect 13324 79400 13364 79409
rect 13132 76243 13172 76252
rect 13228 78812 13268 78821
rect 12844 75989 12884 76084
rect 12940 76084 13076 76124
rect 12748 75151 12788 75160
rect 12844 75872 12884 75881
rect 12748 74696 12788 74705
rect 12748 74561 12788 74656
rect 12748 74444 12788 74453
rect 12748 73688 12788 74404
rect 12748 73639 12788 73648
rect 12844 73460 12884 75832
rect 12940 75788 12980 76084
rect 13036 75956 13076 75965
rect 13228 75956 13268 78772
rect 13324 78056 13364 79360
rect 13324 78007 13364 78016
rect 13076 75916 13268 75956
rect 13324 76292 13364 76301
rect 13324 75956 13364 76252
rect 13036 75907 13076 75916
rect 13324 75872 13364 75916
rect 13228 75832 13364 75872
rect 13132 75788 13172 75797
rect 12940 75748 13076 75788
rect 13036 75452 13076 75748
rect 13036 75403 13076 75412
rect 13036 74276 13076 74285
rect 13036 73772 13076 74236
rect 13132 73856 13172 75748
rect 13132 73807 13172 73816
rect 12556 73420 12692 73460
rect 12748 73420 12884 73460
rect 12940 73732 13076 73772
rect 12460 70832 12500 70841
rect 12460 70697 12500 70792
rect 12556 69992 12596 73420
rect 12460 69952 12596 69992
rect 12652 73184 12692 73193
rect 12652 69992 12692 73144
rect 12460 68984 12500 69952
rect 12652 69943 12692 69952
rect 12748 69908 12788 73420
rect 12844 73352 12884 73361
rect 12844 72260 12884 73312
rect 12940 73184 12980 73732
rect 13132 73688 13172 73697
rect 12940 73135 12980 73144
rect 13036 73604 13076 73613
rect 12844 72125 12884 72220
rect 12844 71420 12884 71515
rect 12844 71371 12884 71380
rect 13036 71420 13076 73564
rect 13132 72932 13172 73648
rect 13132 72883 13172 72892
rect 13036 71371 13076 71380
rect 13132 72512 13172 72521
rect 12844 71252 12884 71261
rect 12844 70664 12884 71212
rect 13036 71000 13076 71009
rect 13036 70832 13076 70960
rect 13132 70916 13172 72472
rect 13132 70867 13172 70876
rect 13036 70783 13076 70792
rect 12844 70615 12884 70624
rect 13132 70748 13172 70757
rect 12748 69859 12788 69868
rect 13036 70580 13076 70589
rect 12460 68935 12500 68944
rect 12556 69824 12596 69833
rect 12460 68732 12500 68741
rect 12460 68396 12500 68692
rect 12460 68347 12500 68356
rect 12460 66212 12500 66221
rect 12460 64616 12500 66172
rect 12460 64567 12500 64576
rect 12460 64448 12500 64457
rect 12556 64448 12596 69784
rect 13036 68900 13076 70540
rect 13132 69068 13172 70708
rect 13228 70496 13268 75832
rect 13420 75452 13460 83812
rect 13516 83684 13556 84820
rect 13612 84811 13652 84820
rect 13708 84440 13748 84449
rect 13804 84440 13844 88600
rect 13748 84400 13844 84440
rect 13900 89228 13940 89237
rect 13708 84104 13748 84400
rect 13900 84356 13940 89188
rect 13708 84055 13748 84064
rect 13804 84316 13940 84356
rect 13996 88892 14036 88901
rect 13996 88052 14036 88852
rect 14092 88052 14132 88061
rect 13996 88012 14092 88052
rect 13996 85112 14036 88012
rect 14092 88003 14132 88012
rect 13516 83635 13556 83644
rect 13612 84020 13652 84029
rect 13516 82088 13556 82097
rect 13516 81752 13556 82048
rect 13516 81703 13556 81712
rect 13516 81584 13556 81593
rect 13516 78812 13556 81544
rect 13516 78763 13556 78772
rect 13612 78644 13652 83980
rect 13708 83936 13748 83945
rect 13708 81332 13748 83896
rect 13804 83096 13844 84316
rect 13996 83768 14036 85072
rect 14092 85868 14132 85877
rect 14092 83936 14132 85828
rect 14188 85196 14228 90448
rect 14380 89396 14420 89405
rect 14284 89060 14324 89069
rect 14284 88925 14324 89020
rect 14380 88892 14420 89356
rect 14380 88843 14420 88852
rect 14284 88808 14324 88817
rect 14284 88556 14324 88768
rect 14284 88507 14324 88516
rect 14188 85147 14228 85156
rect 14284 86036 14324 86045
rect 14188 85028 14228 85037
rect 14188 84944 14228 84988
rect 14188 84893 14228 84904
rect 14188 84692 14228 84701
rect 14188 84272 14228 84652
rect 14284 84440 14324 85996
rect 14380 85616 14420 85625
rect 14380 84524 14420 85576
rect 14380 84475 14420 84484
rect 14668 84860 14708 84869
rect 14284 84391 14324 84400
rect 14668 84440 14708 84820
rect 14668 84391 14708 84400
rect 14380 84356 14420 84365
rect 14188 84232 14324 84272
rect 14092 83887 14132 83896
rect 14188 84104 14228 84113
rect 13804 83047 13844 83056
rect 13900 83600 13940 83609
rect 13804 82844 13844 82853
rect 13804 82172 13844 82804
rect 13804 82004 13844 82132
rect 13804 81955 13844 81964
rect 13708 80576 13748 81292
rect 13708 80527 13748 80536
rect 13804 81836 13844 81845
rect 13804 78896 13844 81796
rect 13900 79316 13940 83560
rect 13996 81920 14036 83728
rect 14092 83768 14132 83777
rect 14092 82928 14132 83728
rect 14188 83012 14228 84064
rect 14284 83684 14324 84232
rect 14284 83549 14324 83644
rect 14380 83180 14420 84316
rect 14380 83131 14420 83140
rect 14476 84272 14516 84281
rect 14284 83012 14324 83021
rect 14188 82972 14284 83012
rect 14324 82972 14420 83012
rect 14092 82888 14228 82928
rect 14092 82760 14132 82769
rect 14092 82625 14132 82720
rect 13996 81871 14036 81880
rect 14092 82508 14132 82517
rect 14092 82004 14132 82468
rect 14092 81836 14132 81964
rect 14092 81787 14132 81796
rect 13900 79267 13940 79276
rect 13996 81752 14036 81761
rect 13420 75403 13460 75412
rect 13516 78604 13652 78644
rect 13708 78856 13804 78896
rect 13516 77636 13556 78604
rect 13612 78140 13652 78149
rect 13612 78005 13652 78100
rect 13708 77888 13748 78856
rect 13804 78847 13844 78856
rect 13900 78896 13940 78907
rect 13900 78812 13940 78856
rect 13900 78763 13940 78772
rect 13420 75284 13460 75293
rect 13324 75116 13364 75125
rect 13324 74981 13364 75076
rect 13324 74528 13364 74537
rect 13324 74393 13364 74488
rect 13420 73688 13460 75244
rect 13516 73772 13556 77596
rect 13612 77848 13748 77888
rect 13804 78308 13844 78317
rect 13612 75956 13652 77848
rect 13804 76796 13844 78268
rect 13708 76124 13748 76133
rect 13708 76040 13748 76084
rect 13708 75989 13748 76000
rect 13612 75536 13652 75916
rect 13612 75487 13652 75496
rect 13708 75788 13748 75797
rect 13708 75284 13748 75748
rect 13708 75235 13748 75244
rect 13804 74948 13844 76756
rect 13804 74444 13844 74908
rect 13708 74404 13804 74444
rect 13708 73856 13748 74404
rect 13804 74395 13844 74404
rect 13900 78056 13940 78065
rect 13804 74276 13844 74285
rect 13804 74141 13844 74236
rect 13900 74108 13940 78016
rect 13996 75788 14036 81712
rect 14188 79904 14228 82888
rect 14284 82877 14324 82972
rect 14284 82676 14324 82685
rect 14284 80828 14324 82636
rect 14380 82256 14420 82972
rect 14380 82207 14420 82216
rect 14380 82088 14420 82097
rect 14380 81836 14420 82048
rect 14476 82004 14516 84232
rect 14476 81955 14516 81964
rect 14572 84188 14612 84197
rect 14380 81796 14516 81836
rect 14284 80779 14324 80788
rect 14380 81164 14420 81173
rect 14188 79855 14228 79864
rect 14284 80324 14324 80333
rect 14092 79820 14132 79829
rect 14092 78224 14132 79780
rect 14092 78175 14132 78184
rect 14188 79652 14228 79661
rect 14092 78056 14132 78065
rect 14092 76964 14132 78016
rect 14092 76915 14132 76924
rect 14092 76712 14132 76807
rect 14092 76663 14132 76672
rect 13996 75739 14036 75748
rect 14092 76292 14132 76301
rect 13900 74059 13940 74068
rect 13996 75200 14036 75209
rect 13708 73807 13748 73816
rect 13516 73723 13556 73732
rect 13804 73772 13844 73781
rect 13420 73604 13460 73648
rect 13324 73564 13460 73604
rect 13324 73016 13364 73564
rect 13804 73352 13844 73732
rect 13324 72967 13364 72976
rect 13708 73184 13748 73193
rect 13420 72008 13460 72017
rect 13420 71420 13460 71968
rect 13420 71371 13460 71380
rect 13228 70447 13268 70456
rect 13324 71336 13364 71345
rect 13324 69152 13364 71296
rect 13420 71252 13460 71261
rect 13420 71084 13460 71212
rect 13420 71035 13460 71044
rect 13708 70916 13748 73144
rect 13804 72932 13844 73312
rect 13804 72883 13844 72892
rect 13900 73772 13940 73781
rect 13228 69068 13268 69077
rect 13132 69028 13228 69068
rect 12652 68860 13076 68900
rect 12652 68564 12692 68860
rect 12652 68515 12692 68524
rect 12940 68564 12980 68573
rect 12980 68524 13076 68564
rect 12940 68496 12980 68524
rect 12940 68312 12980 68321
rect 12940 68177 12980 68272
rect 12748 67892 12788 67901
rect 12748 67724 12788 67852
rect 13036 67892 13076 68524
rect 13036 67843 13076 67852
rect 13228 68396 13268 69028
rect 13324 69017 13364 69112
rect 13420 70876 13748 70916
rect 13804 71168 13844 71177
rect 12748 67675 12788 67684
rect 13132 67136 13172 67145
rect 12844 67052 12884 67061
rect 12748 66800 12788 66809
rect 12652 66296 12692 66305
rect 12652 65624 12692 66256
rect 12652 65575 12692 65584
rect 12748 65372 12788 66760
rect 12748 65237 12788 65332
rect 12844 65456 12884 67012
rect 13132 67001 13172 67096
rect 13036 66716 13076 66725
rect 13036 66128 13076 66676
rect 13036 66079 13076 66088
rect 13228 66128 13268 68356
rect 13420 68396 13460 70876
rect 13612 70748 13652 70757
rect 13612 70412 13652 70708
rect 13420 68347 13460 68356
rect 13516 69740 13556 69749
rect 13420 67808 13460 67817
rect 13420 66464 13460 67768
rect 13516 66884 13556 69700
rect 13612 67052 13652 70372
rect 13708 70076 13748 70085
rect 13708 67220 13748 70036
rect 13804 69152 13844 71128
rect 13804 69103 13844 69112
rect 13804 68900 13844 68909
rect 13804 68396 13844 68860
rect 13804 68347 13844 68356
rect 13708 67171 13748 67180
rect 13612 67012 13748 67052
rect 13516 66632 13556 66844
rect 13516 66583 13556 66592
rect 13420 66424 13652 66464
rect 13228 66079 13268 66088
rect 13516 66128 13556 66137
rect 12500 64408 12596 64448
rect 12652 64784 12692 64793
rect 12460 60248 12500 64408
rect 12556 64280 12596 64289
rect 12556 64112 12596 64240
rect 12556 63356 12596 64072
rect 12652 63944 12692 64744
rect 12652 63608 12692 63904
rect 12652 63559 12692 63568
rect 12748 64616 12788 64625
rect 12748 63608 12788 64576
rect 12748 63559 12788 63568
rect 12556 61172 12596 63316
rect 12652 63440 12692 63449
rect 12652 62348 12692 63400
rect 12748 63188 12788 63197
rect 12748 62516 12788 63148
rect 12748 62467 12788 62476
rect 12844 62516 12884 65416
rect 13132 65456 13172 65465
rect 12940 65036 12980 65045
rect 12940 64901 12980 64996
rect 13132 65036 13172 65416
rect 13516 65456 13556 66088
rect 13516 65407 13556 65416
rect 13132 64987 13172 64996
rect 13420 65372 13460 65381
rect 12940 64280 12980 64289
rect 12940 63608 12980 64240
rect 13132 63860 13172 63869
rect 12940 63568 13076 63608
rect 12844 62467 12884 62476
rect 12940 63440 12980 63449
rect 12652 62308 12788 62348
rect 12556 61123 12596 61132
rect 12652 60752 12692 60761
rect 12652 60500 12692 60712
rect 12652 60451 12692 60460
rect 12652 60332 12692 60341
rect 12460 60208 12596 60248
rect 12460 60080 12500 60089
rect 12460 53360 12500 60040
rect 12556 57812 12596 60208
rect 12652 60197 12692 60292
rect 12556 57224 12596 57772
rect 12556 56300 12596 57184
rect 12556 56251 12596 56260
rect 12652 60080 12692 60089
rect 12652 59912 12692 60040
rect 12652 57140 12692 59872
rect 12748 57560 12788 62308
rect 12748 57511 12788 57520
rect 12844 61760 12884 61769
rect 12844 61592 12884 61720
rect 12652 56216 12692 57100
rect 12652 53696 12692 56176
rect 12748 55628 12788 55637
rect 12748 54788 12788 55588
rect 12844 54956 12884 61552
rect 12940 61508 12980 63400
rect 12940 61459 12980 61468
rect 12940 59576 12980 59585
rect 12940 59324 12980 59536
rect 12940 59275 12980 59284
rect 12940 58988 12980 58997
rect 12940 57896 12980 58948
rect 13036 58820 13076 63568
rect 13132 62684 13172 63820
rect 13228 63776 13268 63785
rect 13268 63736 13364 63776
rect 13228 63727 13268 63736
rect 13324 63272 13364 63736
rect 13420 63524 13460 65332
rect 13420 63475 13460 63484
rect 13516 65288 13556 65297
rect 13324 63223 13364 63232
rect 13132 62635 13172 62644
rect 13228 63188 13268 63197
rect 13036 58771 13076 58780
rect 13132 60080 13172 60089
rect 12940 57847 12980 57856
rect 13036 58652 13076 58661
rect 12844 54907 12884 54916
rect 13036 57476 13076 58612
rect 13132 58568 13172 60040
rect 13132 58433 13172 58528
rect 12748 54748 12884 54788
rect 12652 53647 12692 53656
rect 12460 51260 12500 53320
rect 12748 53528 12788 53537
rect 12748 52604 12788 53488
rect 12844 53276 12884 54748
rect 12940 54284 12980 54293
rect 13036 54284 13076 57436
rect 12980 54244 13076 54284
rect 13132 58316 13172 58325
rect 12940 54216 12980 54244
rect 12844 53227 12884 53236
rect 12460 51211 12500 51220
rect 12556 51764 12596 51773
rect 12556 50252 12596 51724
rect 12748 51764 12788 52564
rect 12844 52772 12884 52781
rect 12844 51932 12884 52732
rect 12844 51883 12884 51892
rect 12748 51596 12788 51724
rect 12748 51092 12788 51556
rect 13132 51512 13172 58276
rect 13228 57392 13268 63148
rect 13324 63104 13364 63113
rect 13324 58316 13364 63064
rect 13420 62684 13460 62693
rect 13420 61676 13460 62644
rect 13516 62600 13556 65248
rect 13612 64868 13652 66424
rect 13612 64819 13652 64828
rect 13612 63524 13652 63533
rect 13708 63524 13748 67012
rect 13804 66380 13844 66389
rect 13804 65876 13844 66340
rect 13804 65827 13844 65836
rect 13804 64700 13844 64709
rect 13804 63608 13844 64660
rect 13900 63776 13940 73732
rect 13996 68984 14036 75160
rect 14092 74528 14132 76252
rect 14188 75956 14228 79612
rect 14188 75907 14228 75916
rect 14284 75284 14324 80284
rect 14380 79820 14420 81124
rect 14380 78308 14420 79780
rect 14380 75956 14420 78268
rect 14476 79064 14516 81796
rect 14572 79736 14612 84148
rect 14668 84188 14708 84197
rect 14668 82760 14708 84148
rect 14764 83540 14804 94648
rect 14860 94100 14900 96688
rect 15052 94268 15092 96688
rect 15052 94219 15092 94228
rect 15244 94184 15284 96688
rect 15436 95696 15476 96688
rect 15436 95647 15476 95656
rect 15628 95024 15668 96688
rect 15820 95024 15860 96688
rect 15916 95024 15956 95033
rect 15820 94984 15916 95024
rect 15628 94975 15668 94984
rect 15916 94975 15956 94984
rect 16012 94688 16052 96688
rect 16204 95024 16244 96688
rect 16204 94975 16244 94984
rect 16396 94940 16436 96688
rect 16396 94891 16436 94900
rect 16012 94639 16052 94648
rect 16300 94856 16340 94865
rect 15244 94135 15284 94144
rect 15340 94604 15380 94613
rect 14860 94051 14900 94060
rect 15148 93932 15188 93941
rect 15148 93797 15188 93892
rect 14956 93764 14996 93773
rect 14860 89396 14900 89405
rect 14860 89261 14900 89356
rect 14860 85532 14900 85541
rect 14860 84524 14900 85492
rect 14860 84475 14900 84484
rect 14860 84356 14900 84365
rect 14860 84221 14900 84316
rect 14764 83500 14900 83540
rect 14764 83096 14804 83191
rect 14764 83047 14804 83056
rect 14668 81416 14708 82720
rect 14764 82928 14804 82937
rect 14764 81836 14804 82888
rect 14860 82172 14900 83500
rect 14956 82424 14996 93724
rect 15340 93620 15380 94564
rect 16204 94184 16244 94193
rect 16204 94049 16244 94144
rect 15244 93580 15380 93620
rect 15436 93680 15476 93689
rect 15244 86204 15284 93580
rect 15340 90404 15380 90413
rect 15340 89648 15380 90364
rect 15340 89599 15380 89608
rect 15340 87884 15380 87893
rect 15340 87749 15380 87844
rect 15244 86155 15284 86164
rect 15340 86456 15380 86465
rect 15052 85868 15092 85877
rect 15052 84524 15092 85828
rect 15052 84475 15092 84484
rect 15244 85028 15284 85037
rect 15244 84944 15284 84988
rect 15244 84356 15284 84904
rect 15340 84440 15380 86416
rect 15340 84391 15380 84400
rect 15052 83600 15092 83695
rect 15052 83551 15092 83560
rect 14956 82375 14996 82384
rect 15052 83432 15092 83441
rect 14860 82123 14900 82132
rect 15052 82088 15092 83392
rect 15052 82039 15092 82048
rect 15148 82760 15188 82769
rect 15148 82256 15188 82720
rect 15244 82508 15284 84316
rect 15244 82459 15284 82468
rect 15340 83348 15380 83357
rect 15340 83180 15380 83308
rect 15340 82760 15380 83140
rect 14764 81787 14804 81796
rect 14860 82004 14900 82013
rect 14668 79820 14708 81376
rect 14860 81500 14900 81964
rect 14764 81332 14804 81341
rect 14764 80492 14804 81292
rect 14764 80443 14804 80452
rect 14668 79780 14804 79820
rect 14572 79696 14708 79736
rect 14476 77804 14516 79024
rect 14476 77755 14516 77764
rect 14572 79568 14612 79577
rect 14476 77636 14516 77645
rect 14476 77048 14516 77596
rect 14476 76999 14516 77008
rect 14380 75907 14420 75916
rect 14284 75235 14324 75244
rect 14188 75200 14228 75209
rect 14188 74612 14228 75160
rect 14188 74563 14228 74572
rect 14284 75116 14324 75125
rect 14092 74479 14132 74488
rect 14188 74276 14228 74285
rect 14092 74108 14132 74117
rect 14092 69908 14132 74068
rect 14188 73772 14228 74236
rect 14188 73723 14228 73732
rect 14092 69859 14132 69868
rect 14188 73268 14228 73277
rect 14188 69152 14228 73228
rect 14188 69103 14228 69112
rect 13996 68935 14036 68944
rect 14188 68984 14228 68993
rect 13996 68312 14036 68407
rect 13996 68263 14036 68272
rect 13996 68060 14036 68069
rect 13996 67556 14036 68020
rect 13996 67507 14036 67516
rect 14092 67724 14132 67733
rect 13996 66968 14036 66977
rect 13996 63860 14036 66928
rect 14092 66884 14132 67684
rect 14092 66835 14132 66844
rect 14092 65372 14132 65381
rect 14092 64868 14132 65332
rect 14092 64819 14132 64828
rect 13996 63811 14036 63820
rect 14092 63944 14132 63953
rect 13900 63727 13940 63736
rect 14092 63776 14132 63904
rect 14092 63727 14132 63736
rect 13996 63692 14036 63701
rect 13804 63568 13940 63608
rect 13708 63484 13844 63524
rect 13612 63356 13652 63484
rect 13612 63307 13652 63316
rect 13708 63272 13748 63281
rect 13516 62551 13556 62560
rect 13612 63188 13652 63197
rect 13420 58484 13460 61636
rect 13420 58435 13460 58444
rect 13516 62264 13556 62273
rect 13516 58484 13556 62224
rect 13612 61844 13652 63148
rect 13612 61795 13652 61804
rect 13708 61676 13748 63232
rect 13516 58435 13556 58444
rect 13612 61172 13652 61181
rect 13324 58276 13556 58316
rect 13228 57343 13268 57352
rect 13324 57812 13364 57821
rect 13324 55124 13364 57772
rect 13420 57140 13460 57149
rect 13420 56384 13460 57100
rect 13420 56335 13460 56344
rect 13324 54788 13364 55084
rect 13420 56216 13460 56225
rect 13420 55040 13460 56176
rect 13420 54991 13460 55000
rect 13324 54739 13364 54748
rect 13324 54032 13364 54041
rect 13324 53360 13364 53992
rect 13324 53311 13364 53320
rect 13132 51463 13172 51472
rect 13228 51680 13268 51689
rect 12748 51043 12788 51052
rect 12556 50203 12596 50212
rect 13228 51008 13268 51640
rect 13228 49580 13268 50968
rect 13228 49531 13268 49540
rect 12844 49412 12884 49421
rect 12748 48740 12788 48749
rect 12364 46003 12404 46012
rect 12460 48656 12500 48665
rect 12460 43868 12500 48616
rect 12652 48656 12692 48665
rect 12556 47060 12596 47069
rect 12556 46556 12596 47020
rect 12556 46507 12596 46516
rect 12556 46304 12596 46313
rect 12556 46169 12596 46264
rect 12364 43828 12500 43868
rect 12556 46052 12596 46061
rect 12364 43532 12404 43828
rect 12364 43483 12404 43492
rect 12460 43700 12500 43709
rect 12172 43180 12308 43220
rect 12172 38324 12212 43180
rect 12460 42020 12500 43660
rect 12268 41852 12308 41861
rect 12268 39752 12308 41812
rect 12460 41432 12500 41980
rect 12460 41264 12500 41392
rect 12460 41215 12500 41224
rect 12364 41180 12404 41189
rect 12364 40676 12404 41140
rect 12364 40627 12404 40636
rect 12364 40508 12404 40517
rect 12556 40508 12596 46012
rect 12652 42776 12692 48616
rect 12748 48605 12788 48700
rect 12652 41012 12692 42736
rect 12748 48236 12788 48245
rect 12748 41936 12788 48196
rect 12844 47228 12884 49372
rect 13420 49328 13460 49337
rect 13420 48740 13460 49288
rect 13420 48691 13460 48700
rect 13516 48572 13556 58276
rect 13612 54452 13652 61132
rect 13708 58988 13748 61636
rect 13708 58939 13748 58948
rect 13804 57140 13844 63484
rect 13900 63440 13940 63568
rect 13900 63391 13940 63400
rect 13900 63188 13940 63197
rect 13900 57812 13940 63148
rect 13996 62600 14036 63652
rect 14092 63440 14132 63449
rect 14092 63104 14132 63400
rect 14092 63055 14132 63064
rect 13996 62551 14036 62560
rect 14092 62936 14132 62945
rect 13996 62432 14036 62441
rect 13996 60836 14036 62392
rect 13996 60787 14036 60796
rect 13900 57763 13940 57772
rect 13996 58652 14036 58661
rect 13612 54403 13652 54412
rect 13708 57100 13844 57140
rect 13708 55628 13748 57100
rect 13900 57056 13940 57065
rect 13804 56972 13844 56981
rect 13804 56384 13844 56932
rect 13804 56300 13844 56344
rect 13804 56220 13844 56260
rect 13900 56804 13940 57016
rect 13900 56300 13940 56764
rect 13900 56251 13940 56260
rect 13708 54788 13748 55588
rect 13708 52688 13748 54748
rect 13708 52639 13748 52648
rect 13996 50252 14036 58612
rect 14092 55460 14132 62896
rect 14188 61088 14228 68944
rect 14284 63692 14324 75076
rect 14572 74528 14612 79528
rect 14668 77468 14708 79696
rect 14668 77419 14708 77428
rect 14764 78980 14804 79780
rect 14572 74479 14612 74488
rect 14668 76796 14708 76805
rect 14476 74444 14516 74453
rect 14380 73772 14420 73781
rect 14380 68648 14420 73732
rect 14380 68599 14420 68608
rect 14380 68396 14420 68405
rect 14380 67556 14420 68356
rect 14380 67507 14420 67516
rect 14380 66548 14420 66557
rect 14380 66212 14420 66508
rect 14380 66163 14420 66172
rect 14284 63643 14324 63652
rect 14380 63692 14420 63701
rect 14188 61039 14228 61048
rect 14284 63524 14324 63533
rect 14092 54116 14132 55420
rect 14092 53360 14132 54076
rect 14092 53311 14132 53320
rect 14188 58400 14228 58409
rect 14188 57392 14228 58360
rect 14284 58064 14324 63484
rect 14380 63356 14420 63652
rect 14380 63307 14420 63316
rect 14380 63188 14420 63197
rect 14380 63053 14420 63148
rect 14380 62936 14420 62945
rect 14380 62432 14420 62896
rect 14380 62383 14420 62392
rect 14380 62180 14420 62189
rect 14380 61760 14420 62140
rect 14380 61711 14420 61720
rect 14380 61424 14420 61433
rect 14380 60248 14420 61384
rect 14380 60199 14420 60208
rect 14380 60080 14420 60089
rect 14380 59945 14420 60040
rect 14284 58015 14324 58024
rect 14380 59324 14420 59333
rect 14380 58652 14420 59284
rect 14188 55628 14228 57352
rect 14284 57812 14324 57821
rect 14284 57140 14324 57772
rect 14284 56300 14324 57100
rect 14284 56251 14324 56260
rect 14188 52772 14228 55588
rect 14284 53528 14324 53537
rect 14284 52856 14324 53488
rect 14380 53528 14420 58612
rect 14476 58484 14516 74404
rect 14572 74360 14612 74369
rect 14572 71588 14612 74320
rect 14668 74024 14708 76756
rect 14764 76292 14804 78940
rect 14860 78812 14900 81460
rect 14860 78763 14900 78772
rect 14956 82004 14996 82013
rect 14860 78224 14900 78233
rect 14860 77132 14900 78184
rect 14860 76460 14900 77092
rect 14860 76411 14900 76420
rect 14764 76243 14804 76252
rect 14860 76208 14900 76217
rect 14668 73975 14708 73984
rect 14764 76040 14804 76049
rect 14668 73688 14708 73697
rect 14668 72764 14708 73648
rect 14764 73460 14804 76000
rect 14860 75200 14900 76168
rect 14860 75151 14900 75160
rect 14764 73420 14900 73460
rect 14668 72715 14708 72724
rect 14668 72596 14708 72605
rect 14668 72428 14708 72556
rect 14668 72379 14708 72388
rect 14572 71420 14612 71548
rect 14572 71371 14612 71380
rect 14668 72260 14708 72269
rect 14668 72008 14708 72220
rect 14572 71252 14612 71261
rect 14572 71117 14612 71212
rect 14572 70748 14612 70757
rect 14572 69992 14612 70708
rect 14572 69943 14612 69952
rect 14572 69236 14612 69245
rect 14572 68816 14612 69196
rect 14572 68312 14612 68776
rect 14572 65960 14612 68272
rect 14668 67472 14708 71968
rect 14860 71588 14900 73420
rect 14956 72428 14996 81964
rect 15148 81668 15188 82216
rect 15340 82172 15380 82720
rect 15340 82123 15380 82132
rect 15340 82004 15380 82013
rect 15148 81628 15284 81668
rect 15148 81080 15188 81089
rect 15052 79148 15092 79157
rect 15052 77552 15092 79108
rect 15148 78980 15188 81040
rect 15148 78931 15188 78940
rect 15052 77503 15092 77512
rect 15148 78812 15188 78821
rect 15148 77384 15188 78772
rect 15052 77344 15188 77384
rect 15052 76376 15092 77344
rect 15052 76327 15092 76336
rect 15148 76964 15188 76973
rect 15052 76208 15092 76217
rect 15052 75620 15092 76168
rect 15052 73688 15092 75580
rect 15052 73639 15092 73648
rect 14956 72379 14996 72388
rect 15052 73520 15092 73529
rect 14956 72260 14996 72269
rect 14956 72008 14996 72220
rect 14956 71959 14996 71968
rect 14764 71548 14900 71588
rect 14764 70412 14804 71548
rect 14956 71420 14996 71429
rect 14764 70363 14804 70372
rect 14860 71336 14900 71345
rect 14668 67423 14708 67432
rect 14764 69488 14804 69497
rect 14764 69152 14804 69448
rect 14572 65911 14612 65920
rect 14668 66296 14708 66305
rect 14668 65372 14708 66256
rect 14764 66128 14804 69112
rect 14860 68144 14900 71296
rect 14956 69320 14996 71380
rect 15052 69488 15092 73480
rect 15052 69439 15092 69448
rect 14956 69280 15092 69320
rect 14860 68095 14900 68104
rect 14956 68984 14996 68993
rect 14764 66079 14804 66088
rect 14860 67640 14900 67649
rect 14860 66884 14900 67600
rect 14668 65288 14708 65332
rect 14476 57308 14516 58444
rect 14572 65204 14612 65213
rect 14572 57980 14612 65164
rect 14668 63356 14708 65248
rect 14764 65960 14804 65969
rect 14764 64532 14804 65920
rect 14860 64700 14900 66844
rect 14860 64651 14900 64660
rect 14764 64492 14900 64532
rect 14668 62180 14708 63316
rect 14668 62131 14708 62140
rect 14764 64364 14804 64373
rect 14668 60164 14708 60175
rect 14668 60080 14708 60124
rect 14668 60031 14708 60040
rect 14572 57931 14612 57940
rect 14668 59828 14708 59837
rect 14668 59408 14708 59788
rect 14668 57896 14708 59368
rect 14764 58904 14804 64324
rect 14764 58855 14804 58864
rect 14668 57847 14708 57856
rect 14764 58148 14804 58157
rect 14476 57259 14516 57268
rect 14668 56216 14708 56225
rect 14380 53479 14420 53488
rect 14476 54200 14516 54209
rect 14380 53360 14420 53371
rect 14380 53276 14420 53320
rect 14380 53196 14420 53236
rect 14284 52816 14420 52856
rect 14188 52732 14324 52772
rect 14188 52604 14228 52613
rect 13996 50203 14036 50212
rect 14092 52100 14132 52109
rect 13516 48523 13556 48532
rect 12940 48068 12980 48077
rect 13228 48068 13268 48077
rect 12980 48028 13076 48068
rect 12940 48000 12980 48028
rect 12844 47179 12884 47188
rect 12940 45800 12980 45809
rect 13036 45800 13076 48028
rect 12980 45760 13076 45800
rect 12940 45732 12980 45760
rect 13228 45716 13268 48028
rect 13996 47228 14036 47237
rect 13996 46640 14036 47188
rect 13996 46591 14036 46600
rect 13612 46556 13652 46565
rect 13420 46472 13460 46481
rect 13420 45968 13460 46432
rect 13420 45919 13460 45928
rect 13228 45667 13268 45676
rect 13516 45716 13556 45725
rect 13420 45044 13460 45053
rect 12844 44792 12884 44801
rect 12844 43784 12884 44752
rect 13420 44456 13460 45004
rect 13420 44407 13460 44416
rect 12844 43448 12884 43744
rect 12844 43399 12884 43408
rect 13228 43784 13268 43793
rect 13036 43364 13076 43373
rect 13036 43280 13076 43324
rect 13036 43229 13076 43240
rect 12748 41887 12788 41896
rect 12844 43196 12884 43205
rect 12652 40963 12692 40972
rect 12364 39920 12404 40468
rect 12364 39871 12404 39880
rect 12460 40468 12596 40508
rect 12652 40844 12692 40853
rect 12268 39703 12308 39712
rect 12268 39650 12308 39659
rect 12268 38492 12308 39610
rect 12268 38443 12308 38452
rect 12364 39584 12404 39593
rect 12212 38284 12308 38324
rect 12172 38275 12212 38284
rect 12172 38156 12212 38165
rect 12172 37652 12212 38116
rect 12172 37603 12212 37612
rect 12268 37904 12308 38284
rect 12268 36812 12308 37864
rect 12364 37148 12404 39544
rect 12460 39164 12500 40468
rect 12556 40256 12596 40265
rect 12556 40004 12596 40216
rect 12556 39668 12596 39964
rect 12652 39752 12692 40804
rect 12844 40508 12884 43156
rect 13036 43112 13076 43121
rect 12940 42440 12980 42449
rect 13036 42440 13076 43072
rect 12980 42400 13076 42440
rect 12940 42372 12980 42400
rect 13036 42272 13076 42281
rect 13036 42104 13076 42232
rect 13036 42055 13076 42064
rect 12940 41936 12980 41945
rect 12980 41896 13076 41936
rect 12940 41868 12980 41896
rect 12940 40844 12980 40853
rect 12940 40709 12980 40804
rect 12748 40468 12884 40508
rect 12748 39836 12788 40468
rect 12844 40340 12884 40349
rect 12844 40205 12884 40300
rect 12940 40172 12980 40181
rect 13036 40172 13076 41896
rect 13228 40592 13268 43744
rect 13420 43448 13460 43457
rect 13324 43112 13364 43121
rect 13324 42977 13364 43072
rect 13324 42692 13364 42701
rect 13324 41348 13364 42652
rect 13420 42188 13460 43408
rect 13420 42139 13460 42148
rect 13516 41432 13556 45676
rect 13612 44960 13652 46516
rect 13612 44204 13652 44920
rect 13612 42356 13652 44164
rect 13900 46556 13940 46565
rect 13900 45632 13940 46516
rect 13900 45044 13940 45592
rect 13612 42307 13652 42316
rect 13708 43364 13748 43373
rect 13708 42188 13748 43324
rect 13804 42776 13844 42871
rect 13804 42727 13844 42736
rect 13324 41299 13364 41308
rect 13420 41392 13556 41432
rect 13612 42148 13748 42188
rect 13804 42608 13844 42617
rect 13420 40760 13460 41392
rect 13612 41348 13652 42148
rect 13420 40711 13460 40720
rect 13516 41308 13652 41348
rect 13708 42020 13748 42029
rect 13708 41348 13748 41980
rect 13804 41852 13844 42568
rect 13804 41803 13844 41812
rect 13804 41684 13844 41693
rect 13804 41549 13844 41644
rect 13708 41308 13844 41348
rect 13228 40543 13268 40552
rect 13324 40508 13364 40517
rect 12980 40132 13076 40172
rect 13132 40424 13172 40433
rect 12940 40104 12980 40132
rect 12748 39796 12884 39836
rect 12652 39712 12788 39752
rect 12556 39619 12596 39628
rect 12652 39584 12692 39593
rect 12652 39449 12692 39544
rect 12652 39248 12692 39257
rect 12652 39164 12692 39208
rect 12460 39124 12596 39164
rect 12460 38912 12500 38921
rect 12460 38408 12500 38872
rect 12460 38359 12500 38368
rect 12556 37988 12596 39124
rect 12652 39113 12692 39124
rect 12748 38912 12788 39712
rect 12748 38863 12788 38872
rect 12460 37948 12596 37988
rect 12652 38660 12692 38669
rect 12460 37316 12500 37948
rect 12460 37267 12500 37276
rect 12556 37736 12596 37745
rect 12364 37108 12500 37148
rect 12076 36427 12116 36436
rect 12172 36772 12308 36812
rect 11980 36091 12020 36100
rect 11980 35972 12020 35983
rect 11980 35888 12020 35932
rect 11980 35839 12020 35848
rect 12172 35552 12212 36772
rect 12268 36644 12308 36653
rect 12268 36140 12308 36604
rect 12268 36091 12308 36100
rect 12364 36140 12404 36149
rect 12076 35512 12212 35552
rect 12268 35888 12308 35897
rect 12076 34628 12116 35512
rect 12076 34579 12116 34588
rect 12172 35300 12212 35309
rect 11692 29287 11732 29296
rect 11788 29672 11828 29681
rect 11692 28580 11732 28591
rect 11692 28496 11732 28540
rect 11692 28447 11732 28456
rect 11308 27152 11348 27161
rect 11308 27068 11348 27112
rect 11308 27017 11348 27028
rect 11404 26900 11444 27532
rect 11404 26851 11444 26860
rect 11500 27404 11540 27413
rect 11308 26732 11348 26741
rect 11348 26692 11444 26732
rect 11308 26683 11348 26692
rect 11308 26480 11348 26489
rect 11308 25976 11348 26440
rect 11308 25927 11348 25936
rect 11308 25808 11348 25817
rect 11308 25556 11348 25768
rect 11308 25507 11348 25516
rect 11308 25388 11348 25397
rect 11308 24800 11348 25348
rect 11308 24751 11348 24760
rect 11308 22196 11348 22205
rect 11212 22156 11308 22196
rect 11212 21944 11252 21953
rect 11212 21809 11252 21904
rect 11308 21860 11348 22156
rect 11308 21811 11348 21820
rect 11212 21356 11252 21365
rect 11212 20432 11252 21316
rect 11212 20383 11252 20392
rect 11308 20600 11348 20609
rect 11116 20215 11156 20224
rect 11212 20012 11252 20021
rect 11020 17695 11060 17704
rect 11116 19972 11212 20012
rect 11116 19508 11156 19972
rect 11212 19963 11252 19972
rect 11020 17324 11060 17333
rect 11020 14552 11060 17284
rect 11020 14503 11060 14512
rect 10924 8252 10964 8800
rect 11020 14384 11060 14393
rect 11020 8420 11060 14344
rect 11116 10352 11156 19468
rect 11212 19676 11252 19685
rect 11212 14384 11252 19636
rect 11212 14335 11252 14344
rect 11116 10303 11156 10312
rect 11212 13544 11252 13553
rect 11020 8371 11060 8380
rect 11116 10016 11156 10025
rect 10924 8203 10964 8212
rect 11116 6488 11156 9976
rect 11020 6448 11156 6488
rect 10924 5816 10964 5825
rect 10924 4892 10964 5776
rect 10924 4843 10964 4852
rect 10828 4087 10868 4096
rect 10924 4220 10964 4229
rect 10060 2960 10100 2969
rect 9772 2860 10004 2900
rect 9676 2575 9716 2584
rect 9292 2456 9332 2465
rect 9100 1828 9236 1868
rect 9196 1784 9236 1828
rect 9196 1735 9236 1744
rect 9100 1700 9140 1709
rect 9100 80 9140 1660
rect 9292 80 9332 2416
rect 9676 2456 9716 2465
rect 9388 2372 9428 2381
rect 9388 1952 9428 2332
rect 9388 1903 9428 1912
rect 9484 1700 9524 1709
rect 9484 80 9524 1660
rect 9676 80 9716 2416
rect 9772 2456 9812 2465
rect 9772 1952 9812 2416
rect 9772 1903 9812 1912
rect 9868 1700 9908 1709
rect 9868 80 9908 1660
rect 9964 1532 10004 2860
rect 10060 2825 10100 2920
rect 10156 2708 10196 2717
rect 9964 1483 10004 1492
rect 10060 2456 10100 2465
rect 10060 80 10100 2416
rect 10156 1952 10196 2668
rect 10348 2624 10388 2633
rect 10348 2489 10388 2584
rect 10732 2624 10772 2633
rect 10156 1903 10196 1912
rect 10444 2456 10484 2465
rect 10252 1700 10292 1709
rect 10252 80 10292 1660
rect 10444 80 10484 2416
rect 10636 1700 10676 1709
rect 10636 80 10676 1660
rect 10732 1532 10772 2584
rect 10732 1483 10772 1492
rect 10828 2456 10868 2465
rect 10828 80 10868 2416
rect 10924 1952 10964 4180
rect 11020 2708 11060 6448
rect 11212 2900 11252 13504
rect 11308 10856 11348 20560
rect 11404 18836 11444 26692
rect 11500 26144 11540 27364
rect 11596 26228 11636 28372
rect 11788 28160 11828 29632
rect 11788 28111 11828 28120
rect 11788 27656 11828 27665
rect 11596 26179 11636 26188
rect 11692 27320 11732 27329
rect 11692 26312 11732 27280
rect 11500 26095 11540 26104
rect 11692 26144 11732 26272
rect 11692 26095 11732 26104
rect 11596 26060 11636 26069
rect 11500 25976 11540 25985
rect 11500 22784 11540 25936
rect 11500 22735 11540 22744
rect 11596 24548 11636 26020
rect 11788 25388 11828 27616
rect 11500 22364 11540 22459
rect 11500 22315 11540 22324
rect 11500 22112 11540 22121
rect 11500 21977 11540 22072
rect 11404 18787 11444 18796
rect 11500 21860 11540 21869
rect 11404 17156 11444 17165
rect 11404 14384 11444 17116
rect 11500 17072 11540 21820
rect 11596 19424 11636 24508
rect 11692 25348 11828 25388
rect 11692 20264 11732 25348
rect 11884 24548 11924 32152
rect 11980 34460 12020 34469
rect 11980 33200 12020 34420
rect 11980 32948 12020 33160
rect 11980 29756 12020 32908
rect 12076 34376 12116 34385
rect 12076 32192 12116 34336
rect 12076 31436 12116 32152
rect 12076 31387 12116 31396
rect 12076 31184 12116 31195
rect 12076 31100 12116 31144
rect 12076 31051 12116 31060
rect 11980 29716 12116 29756
rect 11980 29588 12020 29597
rect 11980 29084 12020 29548
rect 11980 27572 12020 29044
rect 11980 27523 12020 27532
rect 11980 27404 12020 27413
rect 11980 26144 12020 27364
rect 11980 25892 12020 26104
rect 11980 25843 12020 25852
rect 11884 23876 11924 24508
rect 11884 23827 11924 23836
rect 11980 23792 12020 23801
rect 11884 23288 11924 23297
rect 11788 23036 11828 23045
rect 11788 21608 11828 22996
rect 11788 21559 11828 21568
rect 11692 20215 11732 20224
rect 11788 20852 11828 20861
rect 11596 19375 11636 19384
rect 11692 20012 11732 20021
rect 11692 18668 11732 19972
rect 11500 17023 11540 17032
rect 11596 18628 11732 18668
rect 11596 14972 11636 18628
rect 11596 14923 11636 14932
rect 11692 18500 11732 18509
rect 11692 17744 11732 18460
rect 11404 14335 11444 14344
rect 11404 13964 11444 13973
rect 11404 13829 11444 13924
rect 11596 13964 11636 13973
rect 11500 13124 11540 13133
rect 11500 12980 11540 13084
rect 11308 10807 11348 10816
rect 11404 12940 11540 12980
rect 11308 10688 11348 10697
rect 11308 7160 11348 10648
rect 11404 10268 11444 12940
rect 11404 10219 11444 10228
rect 11500 11192 11540 11201
rect 11308 5816 11348 7120
rect 11308 5767 11348 5776
rect 11404 10100 11444 10109
rect 11404 8924 11444 10060
rect 11500 9764 11540 11152
rect 11500 9715 11540 9724
rect 11404 5312 11444 8884
rect 11596 8756 11636 13924
rect 11692 11948 11732 17704
rect 11788 13292 11828 20812
rect 11788 13243 11828 13252
rect 11788 13040 11828 13049
rect 11788 12536 11828 13000
rect 11788 12487 11828 12496
rect 11692 11908 11828 11948
rect 11692 11780 11732 11789
rect 11692 11444 11732 11740
rect 11692 11395 11732 11404
rect 11788 11276 11828 11908
rect 11788 10268 11828 11236
rect 11884 11192 11924 23248
rect 11980 20264 12020 23752
rect 12076 22280 12116 29716
rect 12172 28916 12212 35260
rect 12268 31856 12308 35848
rect 12268 31807 12308 31816
rect 12268 31100 12308 31109
rect 12268 29252 12308 31060
rect 12268 29203 12308 29212
rect 12364 30596 12404 36100
rect 12460 35888 12500 37108
rect 12556 36728 12596 37696
rect 12652 37484 12692 38620
rect 12748 38492 12788 38501
rect 12748 38156 12788 38452
rect 12748 38107 12788 38116
rect 12844 38240 12884 39796
rect 12940 39752 12980 39761
rect 12940 39617 12980 39712
rect 13036 39584 13076 39593
rect 13036 39449 13076 39544
rect 13132 39500 13172 40384
rect 13132 39451 13172 39460
rect 13228 40340 13268 40349
rect 13228 39416 13268 40300
rect 13228 39332 13268 39376
rect 13228 39281 13268 39292
rect 13036 39248 13076 39257
rect 13036 38912 13076 39208
rect 13036 38863 13076 38872
rect 13132 39248 13172 39257
rect 12652 37435 12692 37444
rect 12748 37988 12788 37997
rect 12748 37400 12788 37948
rect 12844 37820 12884 38200
rect 12844 37771 12884 37780
rect 13036 38240 13076 38249
rect 12748 37351 12788 37360
rect 12844 37568 12884 37577
rect 12556 36679 12596 36688
rect 12652 37316 12692 37325
rect 12460 35839 12500 35848
rect 12460 35720 12500 35729
rect 12460 34712 12500 35680
rect 12556 35720 12596 35729
rect 12556 35300 12596 35680
rect 12556 35251 12596 35260
rect 12556 34880 12596 34889
rect 12652 34880 12692 37276
rect 12748 36896 12788 36905
rect 12748 36392 12788 36856
rect 12844 36728 12884 37528
rect 13036 37484 13076 38200
rect 13132 37652 13172 39208
rect 13228 38996 13268 39005
rect 13228 38324 13268 38956
rect 13228 38275 13268 38284
rect 13132 37603 13172 37612
rect 13324 37568 13364 40468
rect 13516 39752 13556 41308
rect 13708 41180 13748 41189
rect 13420 39668 13460 39677
rect 13420 39248 13460 39628
rect 13516 39617 13556 39712
rect 13612 40676 13652 40685
rect 13420 39199 13460 39208
rect 13516 39416 13556 39425
rect 13516 38996 13556 39376
rect 13516 38240 13556 38956
rect 13516 38191 13556 38200
rect 13516 38072 13556 38081
rect 13324 37519 13364 37528
rect 13420 37652 13460 37661
rect 13036 37444 13268 37484
rect 12844 36688 13172 36728
rect 12940 36476 12980 36485
rect 12844 36392 12884 36401
rect 12748 36352 12844 36392
rect 12748 35972 12788 35981
rect 12748 35837 12788 35932
rect 12596 34840 12692 34880
rect 12556 34831 12596 34840
rect 12844 34796 12884 36352
rect 12940 35888 12980 36436
rect 12940 35839 12980 35848
rect 13036 35972 13076 35981
rect 13036 35132 13076 35932
rect 13036 35083 13076 35092
rect 12652 34756 12884 34796
rect 12460 34672 12596 34712
rect 12460 34544 12500 34553
rect 12460 34409 12500 34504
rect 12556 34376 12596 34672
rect 12556 34327 12596 34336
rect 12460 32528 12500 32537
rect 12460 32360 12500 32488
rect 12460 32311 12500 32320
rect 12556 32444 12596 32453
rect 12556 31940 12596 32404
rect 12364 29840 12404 30556
rect 12172 28867 12212 28876
rect 12172 27572 12212 27581
rect 12172 26816 12212 27532
rect 12268 27572 12308 27581
rect 12268 26900 12308 27532
rect 12268 26851 12308 26860
rect 12172 26767 12212 26776
rect 12076 21524 12116 22240
rect 12076 21475 12116 21484
rect 12172 26648 12212 26657
rect 12172 23708 12212 26608
rect 12268 26648 12308 26657
rect 12268 26060 12308 26608
rect 12268 25388 12308 26020
rect 12268 25339 12308 25348
rect 12364 25220 12404 29800
rect 11980 20215 12020 20224
rect 12076 20264 12116 20273
rect 11980 20012 12020 20021
rect 11980 19508 12020 19972
rect 11980 19459 12020 19468
rect 12076 18332 12116 20224
rect 12076 18283 12116 18292
rect 12172 18164 12212 23668
rect 12268 25180 12404 25220
rect 12460 31856 12500 31865
rect 12268 23120 12308 25180
rect 12268 23071 12308 23080
rect 12364 25052 12404 25061
rect 12268 22952 12308 22961
rect 12364 22952 12404 25012
rect 12460 23624 12500 31816
rect 12556 29084 12596 31900
rect 12652 30008 12692 34756
rect 13132 34712 13172 36688
rect 12652 29959 12692 29968
rect 12748 34672 13172 34712
rect 12748 31436 12788 34672
rect 12940 34544 12980 34553
rect 12980 34504 13076 34544
rect 12940 34476 12980 34504
rect 13036 33536 13076 34504
rect 12844 33496 13076 33536
rect 12844 32948 12884 33496
rect 13228 33200 13268 37444
rect 13420 36224 13460 37612
rect 13516 37484 13556 38032
rect 13516 37435 13556 37444
rect 13612 37400 13652 40636
rect 13708 38996 13748 41140
rect 13804 41012 13844 41308
rect 13804 40963 13844 40972
rect 13804 40508 13844 40517
rect 13804 39248 13844 40468
rect 13804 39199 13844 39208
rect 13900 39920 13940 45004
rect 13996 42020 14036 42029
rect 13996 41600 14036 41980
rect 13996 41551 14036 41560
rect 13708 38947 13748 38956
rect 13804 38996 13844 39005
rect 13804 38324 13844 38956
rect 13612 37351 13652 37360
rect 13708 38284 13844 38324
rect 13708 37232 13748 38284
rect 13804 38156 13844 38165
rect 13804 37484 13844 38116
rect 13804 37435 13844 37444
rect 13420 36175 13460 36184
rect 13516 37192 13748 37232
rect 13420 36056 13460 36065
rect 13324 35972 13364 35981
rect 13324 35384 13364 35932
rect 13324 35335 13364 35344
rect 13228 33151 13268 33160
rect 13324 35048 13364 35057
rect 13324 34880 13364 35008
rect 13420 34964 13460 36016
rect 13420 34915 13460 34924
rect 13228 33032 13268 33041
rect 12844 32908 13076 32948
rect 12748 29672 12788 31396
rect 12844 31016 12884 31025
rect 12844 30344 12884 30976
rect 12940 30764 12980 30773
rect 12940 30629 12980 30724
rect 12844 30295 12884 30304
rect 12940 30176 12980 30185
rect 12844 30008 12884 30017
rect 12844 29873 12884 29968
rect 12940 29840 12980 30136
rect 12940 29791 12980 29800
rect 12556 29035 12596 29044
rect 12652 29252 12692 29261
rect 12556 28916 12596 28925
rect 12556 23708 12596 28876
rect 12652 27488 12692 29212
rect 12748 28580 12788 29632
rect 12844 29672 12884 29681
rect 12844 29000 12884 29632
rect 12844 28951 12884 28960
rect 12940 29336 12980 29345
rect 12748 28531 12788 28540
rect 12844 28160 12884 28169
rect 12652 27439 12692 27448
rect 12748 27740 12788 27749
rect 12652 26984 12692 26993
rect 12652 23876 12692 26944
rect 12748 25388 12788 27700
rect 12844 25976 12884 28120
rect 12940 26144 12980 29296
rect 13036 26984 13076 32908
rect 13132 31520 13172 31529
rect 13132 31268 13172 31480
rect 13132 31219 13172 31228
rect 13132 30932 13172 30941
rect 13132 30797 13172 30892
rect 13132 30512 13172 30607
rect 13132 30463 13172 30472
rect 13132 30344 13172 30353
rect 13132 29252 13172 30304
rect 13132 29203 13172 29212
rect 13036 26935 13076 26944
rect 13132 27572 13172 27581
rect 12940 26095 12980 26104
rect 13036 26564 13076 26573
rect 12844 25936 12980 25976
rect 12748 25348 12884 25388
rect 12652 23827 12692 23836
rect 12748 25220 12788 25229
rect 12748 24884 12788 25180
rect 12556 23668 12692 23708
rect 12460 23584 12596 23624
rect 12308 22912 12404 22952
rect 12460 23456 12500 23465
rect 12268 18752 12308 22912
rect 12364 21440 12404 21449
rect 12364 21305 12404 21400
rect 12460 20012 12500 23416
rect 12364 19844 12404 19853
rect 12364 18920 12404 19804
rect 12460 19340 12500 19972
rect 12460 19291 12500 19300
rect 12364 18871 12404 18880
rect 12268 18712 12500 18752
rect 11980 18124 12212 18164
rect 12268 18332 12308 18341
rect 11980 17828 12020 18124
rect 11980 17779 12020 17788
rect 12076 17996 12116 18005
rect 12076 12620 12116 17956
rect 12268 17912 12308 18292
rect 12268 16988 12308 17872
rect 12268 16939 12308 16948
rect 12268 16316 12308 16325
rect 12172 16064 12212 16073
rect 12172 14804 12212 16024
rect 12268 15476 12308 16276
rect 12364 16232 12404 16241
rect 12364 15560 12404 16192
rect 12460 15728 12500 18712
rect 12556 17996 12596 23584
rect 12652 19508 12692 23668
rect 12748 20852 12788 24844
rect 12844 23036 12884 25348
rect 12940 23456 12980 25936
rect 12940 23407 12980 23416
rect 13036 23204 13076 26524
rect 13132 26312 13172 27532
rect 13132 26060 13172 26272
rect 13132 26011 13172 26020
rect 13132 25892 13172 25901
rect 13132 24212 13172 25852
rect 13228 25052 13268 32992
rect 13324 31268 13364 34840
rect 13516 32276 13556 37192
rect 13708 36728 13748 36737
rect 13612 36644 13652 36655
rect 13612 36560 13652 36604
rect 13708 36593 13748 36688
rect 13804 36644 13844 36653
rect 13612 36140 13652 36520
rect 13804 36509 13844 36604
rect 13612 36091 13652 36100
rect 13708 36476 13748 36485
rect 13708 33032 13748 36436
rect 13804 36224 13844 36233
rect 13804 33620 13844 36184
rect 13804 33116 13844 33580
rect 13804 33067 13844 33076
rect 13708 32983 13748 32992
rect 13804 32948 13844 32957
rect 13708 32864 13748 32873
rect 13708 32276 13748 32824
rect 13516 32236 13652 32276
rect 13516 32108 13556 32117
rect 13324 31228 13460 31268
rect 13324 30344 13364 30353
rect 13324 29756 13364 30304
rect 13324 29707 13364 29716
rect 13324 29168 13364 29177
rect 13324 29084 13364 29128
rect 13324 29033 13364 29044
rect 13228 24548 13268 25012
rect 13228 24499 13268 24508
rect 13132 24163 13172 24172
rect 13228 24380 13268 24389
rect 13036 23155 13076 23164
rect 12844 22987 12884 22996
rect 12844 22868 12884 22877
rect 12844 22364 12884 22828
rect 12940 22448 12980 22457
rect 12980 22408 13076 22448
rect 12940 22380 12980 22408
rect 12844 22315 12884 22324
rect 12748 20803 12788 20812
rect 12844 21272 12884 21281
rect 12844 20684 12884 21232
rect 12940 20684 12980 20693
rect 12844 20644 12940 20684
rect 12652 19468 12788 19508
rect 12556 17947 12596 17956
rect 12652 19340 12692 19349
rect 12460 15679 12500 15688
rect 12556 17828 12596 17837
rect 12364 15511 12404 15520
rect 12268 15427 12308 15436
rect 12172 13964 12212 14764
rect 12364 14804 12404 14813
rect 12172 13915 12212 13924
rect 12268 14552 12308 14561
rect 12076 12571 12116 12580
rect 11884 11143 11924 11152
rect 12076 12452 12116 12461
rect 12076 10856 12116 12412
rect 12116 10816 12212 10856
rect 12076 10807 12116 10816
rect 12172 10352 12212 10816
rect 12172 10303 12212 10312
rect 11788 10219 11828 10228
rect 12076 10268 12116 10277
rect 11980 10184 12020 10193
rect 11884 9428 11924 9437
rect 11884 8924 11924 9388
rect 11884 8875 11924 8884
rect 11980 8840 12020 10144
rect 11980 8791 12020 8800
rect 11596 7916 11636 8716
rect 11788 8756 11828 8765
rect 11788 8168 11828 8716
rect 11788 8119 11828 8128
rect 11980 8672 12020 8681
rect 11596 7244 11636 7876
rect 11596 7195 11636 7204
rect 11500 6320 11540 6329
rect 11500 5732 11540 6280
rect 11596 5732 11636 5741
rect 11500 5692 11596 5732
rect 11596 5683 11636 5692
rect 11404 5263 11444 5272
rect 11500 5564 11540 5573
rect 11404 5060 11444 5069
rect 11404 4808 11444 5020
rect 11500 4976 11540 5524
rect 11500 4927 11540 4936
rect 11884 4892 11924 4901
rect 11404 4768 11540 4808
rect 11500 4220 11540 4768
rect 11884 4556 11924 4852
rect 11884 4507 11924 4516
rect 11500 4171 11540 4180
rect 11980 3548 12020 8632
rect 12076 7076 12116 10228
rect 12076 7027 12116 7036
rect 12172 6992 12212 7001
rect 12172 6404 12212 6952
rect 12076 5480 12116 5489
rect 12076 5228 12116 5440
rect 12076 5179 12116 5188
rect 12076 4892 12116 4901
rect 12076 4472 12116 4852
rect 12076 4423 12116 4432
rect 12172 4220 12212 6364
rect 12172 4171 12212 4180
rect 11980 3499 12020 3508
rect 11020 2659 11060 2668
rect 11116 2860 11252 2900
rect 11116 2624 11156 2860
rect 11116 2575 11156 2584
rect 11692 2708 11732 2717
rect 10924 1903 10964 1912
rect 11308 2036 11348 2045
rect 11308 1901 11348 1996
rect 11500 1952 11540 1961
rect 11500 1817 11540 1912
rect 11212 1784 11252 1793
rect 11020 1700 11060 1709
rect 11020 80 11060 1660
rect 11212 80 11252 1744
rect 11404 1700 11444 1709
rect 11404 80 11444 1660
rect 11596 1700 11636 1709
rect 11596 80 11636 1660
rect 11692 1616 11732 2668
rect 12268 2624 12308 14512
rect 12364 14216 12404 14764
rect 12364 14167 12404 14176
rect 12460 14552 12500 14561
rect 12460 13964 12500 14512
rect 12460 13915 12500 13924
rect 12460 12452 12500 12461
rect 12460 10940 12500 12412
rect 12460 10436 12500 10900
rect 12460 10387 12500 10396
rect 12364 10352 12404 10361
rect 12364 9344 12404 10312
rect 12364 8756 12404 9304
rect 12364 8707 12404 8716
rect 12556 8588 12596 17788
rect 12652 17156 12692 19300
rect 12652 17107 12692 17116
rect 12556 7328 12596 8548
rect 12556 7279 12596 7288
rect 12652 14300 12692 14309
rect 12364 6992 12404 7001
rect 12364 6656 12404 6952
rect 12364 6607 12404 6616
rect 12460 5732 12500 5741
rect 12460 3968 12500 5692
rect 12556 5228 12596 5237
rect 12556 4892 12596 5188
rect 12556 4843 12596 4852
rect 12556 4724 12596 4733
rect 12556 4388 12596 4684
rect 12556 4339 12596 4348
rect 12460 3919 12500 3928
rect 12652 2900 12692 14260
rect 12748 13964 12788 19468
rect 12844 18920 12884 20644
rect 12940 20635 12980 20644
rect 13036 19088 13076 22408
rect 13036 19039 13076 19048
rect 13132 22364 13172 22373
rect 12844 18880 13076 18920
rect 12940 18416 12980 18425
rect 12940 16232 12980 18376
rect 13036 17072 13076 18880
rect 13132 18416 13172 22324
rect 13228 19424 13268 24340
rect 13324 24212 13364 24221
rect 13324 21188 13364 24172
rect 13324 21139 13364 21148
rect 13324 20096 13364 20105
rect 13324 19961 13364 20056
rect 13228 19375 13268 19384
rect 13132 18367 13172 18376
rect 13324 18584 13364 18593
rect 13324 17408 13364 18544
rect 13036 17032 13172 17072
rect 12940 14804 12980 16192
rect 12748 13924 12884 13964
rect 12748 13796 12788 13805
rect 12748 12032 12788 13756
rect 12844 13628 12884 13924
rect 12940 13880 12980 14764
rect 13036 15476 13076 15485
rect 13036 15056 13076 15436
rect 13036 14720 13076 15016
rect 13036 14671 13076 14680
rect 12940 13831 12980 13840
rect 12844 13579 12884 13588
rect 13036 13544 13076 13553
rect 12940 13208 12980 13217
rect 12940 12980 12980 13168
rect 12844 12940 12980 12980
rect 12844 12536 12884 12940
rect 12844 12487 12884 12496
rect 12940 12452 12980 12461
rect 12940 12317 12980 12412
rect 12940 12032 12980 12041
rect 12748 11992 12940 12032
rect 12844 11780 12884 11992
rect 12940 11983 12980 11992
rect 12940 11780 12980 11789
rect 12844 11740 12940 11780
rect 12940 11731 12980 11740
rect 12844 10436 12884 10445
rect 12748 10100 12788 10109
rect 12748 9512 12788 10060
rect 12748 8756 12788 9472
rect 12748 5396 12788 8716
rect 12844 9428 12884 10396
rect 12844 8672 12884 9388
rect 12844 8623 12884 8632
rect 13036 7832 13076 13504
rect 13132 13292 13172 17032
rect 13228 15728 13268 15737
rect 13228 15308 13268 15688
rect 13228 15259 13268 15268
rect 13132 13243 13172 13252
rect 13228 13796 13268 13805
rect 13132 13124 13172 13133
rect 13132 9176 13172 13084
rect 13132 9127 13172 9136
rect 13036 7783 13076 7792
rect 13132 8924 13172 8933
rect 13132 6404 13172 8884
rect 12844 6364 13172 6404
rect 12844 5564 12884 6364
rect 13036 6236 13076 6245
rect 13036 5816 13076 6196
rect 13036 5767 13076 5776
rect 13132 6152 13172 6161
rect 12844 5515 12884 5524
rect 12748 5356 12884 5396
rect 12268 2575 12308 2584
rect 12460 2860 12692 2900
rect 12748 3296 12788 3305
rect 12268 2456 12308 2465
rect 12268 1952 12308 2416
rect 12460 2036 12500 2860
rect 12460 1987 12500 1996
rect 12556 2456 12596 2465
rect 12268 1903 12308 1912
rect 11692 1567 11732 1576
rect 11788 1784 11828 1793
rect 11788 80 11828 1744
rect 11980 1700 12020 1709
rect 11980 80 12020 1660
rect 12172 1700 12212 1709
rect 12172 80 12212 1660
rect 12364 1616 12404 1625
rect 12364 80 12404 1576
rect 12556 80 12596 2416
rect 12748 2120 12788 3256
rect 12844 2708 12884 5356
rect 13132 5144 13172 6112
rect 13132 5095 13172 5104
rect 12844 2659 12884 2668
rect 13036 3464 13076 3473
rect 12940 2456 12980 2465
rect 12748 2071 12788 2080
rect 12844 2416 12940 2456
rect 12652 2036 12692 2047
rect 12652 1952 12692 1996
rect 12652 1903 12692 1912
rect 12748 1784 12788 1793
rect 12748 80 12788 1744
rect 12844 440 12884 2416
rect 12940 2407 12980 2416
rect 13036 1952 13076 3424
rect 13228 2900 13268 13756
rect 13324 9596 13364 17368
rect 13420 13208 13460 31228
rect 13516 29336 13556 32068
rect 13516 29287 13556 29296
rect 13516 29084 13556 29093
rect 13516 25892 13556 29044
rect 13612 28076 13652 32236
rect 13708 32227 13748 32236
rect 13804 32108 13844 32908
rect 13708 32024 13748 32033
rect 13708 31856 13748 31984
rect 13804 32024 13844 32068
rect 13804 31975 13844 31984
rect 13708 30596 13748 31816
rect 13900 31688 13940 39880
rect 13996 40592 14036 40601
rect 13996 39584 14036 40552
rect 14092 40340 14132 52060
rect 14188 49832 14228 52564
rect 14188 49783 14228 49792
rect 14284 48068 14324 52732
rect 14380 51260 14420 52816
rect 14380 51211 14420 51220
rect 14476 48908 14516 54160
rect 14572 53612 14612 53621
rect 14572 51008 14612 53572
rect 14572 50959 14612 50968
rect 14476 48859 14516 48868
rect 14284 48019 14324 48028
rect 14572 47228 14612 47237
rect 14188 47060 14228 47069
rect 14188 45800 14228 47020
rect 14476 46556 14516 46565
rect 14188 45751 14228 45760
rect 14380 46472 14420 46481
rect 14380 45800 14420 46432
rect 14188 44960 14228 44969
rect 14188 44825 14228 44920
rect 14380 44960 14420 45760
rect 14476 46388 14516 46516
rect 14476 45044 14516 46348
rect 14572 45464 14612 47188
rect 14572 45415 14612 45424
rect 14476 44995 14516 45004
rect 14380 44911 14420 44920
rect 14188 44540 14228 44549
rect 14188 43364 14228 44500
rect 14188 43315 14228 43324
rect 14284 43868 14324 43877
rect 14188 42692 14228 42701
rect 14284 42692 14324 43828
rect 14572 43532 14612 43541
rect 14476 43448 14516 43457
rect 14380 43280 14420 43289
rect 14380 42860 14420 43240
rect 14380 42811 14420 42820
rect 14284 42652 14420 42692
rect 14188 42020 14228 42652
rect 14188 41971 14228 41980
rect 14284 42524 14324 42533
rect 14188 41768 14228 41777
rect 14188 41633 14228 41728
rect 14188 41432 14228 41441
rect 14188 41297 14228 41392
rect 14188 41096 14228 41105
rect 14188 40961 14228 41056
rect 14092 40291 14132 40300
rect 14188 40424 14228 40433
rect 14092 40172 14132 40181
rect 14092 39836 14132 40132
rect 14092 39787 14132 39796
rect 14092 39584 14132 39593
rect 13996 39544 14092 39584
rect 13996 38912 14036 38921
rect 13996 38777 14036 38872
rect 13900 31639 13940 31648
rect 13996 36224 14036 36233
rect 13708 30547 13748 30556
rect 13900 31436 13940 31445
rect 13900 30596 13940 31396
rect 13900 30176 13940 30556
rect 13900 30127 13940 30136
rect 13900 30008 13940 30017
rect 13900 29840 13940 29968
rect 13900 29791 13940 29800
rect 13708 29756 13748 29765
rect 13708 29504 13748 29716
rect 13708 29455 13748 29464
rect 13708 29336 13748 29345
rect 13708 29252 13748 29296
rect 13996 29252 14036 36184
rect 14092 33788 14132 39544
rect 14188 39164 14228 40384
rect 14188 39115 14228 39124
rect 14092 33739 14132 33748
rect 14188 36728 14228 36737
rect 13708 29201 13748 29212
rect 13900 29212 14036 29252
rect 14092 32948 14132 32957
rect 13612 28027 13652 28036
rect 13804 29168 13844 29177
rect 13516 25843 13556 25852
rect 13708 27572 13748 27581
rect 13708 25808 13748 27532
rect 13804 27572 13844 29128
rect 13804 27523 13844 27532
rect 13804 26900 13844 26909
rect 13804 25976 13844 26860
rect 13804 25927 13844 25936
rect 13708 25768 13844 25808
rect 13516 25136 13556 25145
rect 13516 24548 13556 25096
rect 13516 23876 13556 24508
rect 13516 21524 13556 23836
rect 13612 23624 13652 23633
rect 13612 23036 13652 23584
rect 13612 22987 13652 22996
rect 13708 23204 13748 23213
rect 13516 20768 13556 21484
rect 13612 21440 13652 21449
rect 13612 21188 13652 21400
rect 13612 21139 13652 21148
rect 13516 20719 13556 20728
rect 13612 20936 13652 20945
rect 13612 20600 13652 20896
rect 13516 20560 13652 20600
rect 13516 20180 13556 20560
rect 13516 20131 13556 20140
rect 13612 20432 13652 20441
rect 13420 13159 13460 13168
rect 13516 19928 13556 19937
rect 13420 13040 13460 13049
rect 13420 12452 13460 13000
rect 13516 12788 13556 19888
rect 13612 18164 13652 20392
rect 13708 19928 13748 23164
rect 13708 19879 13748 19888
rect 13804 19172 13844 25768
rect 13900 25304 13940 29212
rect 13996 28412 14036 28421
rect 13996 26648 14036 28372
rect 13996 26599 14036 26608
rect 13996 26312 14036 26321
rect 13996 26177 14036 26272
rect 13900 25255 13940 25264
rect 13996 25976 14036 25985
rect 13996 24296 14036 25936
rect 13900 24256 14036 24296
rect 13900 23036 13940 24256
rect 13996 23792 14036 23801
rect 13996 23657 14036 23752
rect 13900 22987 13940 22996
rect 13900 22868 13940 22877
rect 13900 22532 13940 22828
rect 13940 22492 14036 22532
rect 13900 22483 13940 22492
rect 13996 22280 14036 22492
rect 13996 22231 14036 22240
rect 13900 22196 13940 22205
rect 13900 21524 13940 22156
rect 13900 21475 13940 21484
rect 13996 21356 14036 21365
rect 13900 20432 13940 20441
rect 13900 20012 13940 20392
rect 13900 19963 13940 19972
rect 13900 19844 13940 19853
rect 13900 19256 13940 19804
rect 13996 19340 14036 21316
rect 14092 20180 14132 32908
rect 14188 32108 14228 36688
rect 14284 35888 14324 42484
rect 14380 38996 14420 42652
rect 14476 42440 14516 43408
rect 14476 42391 14516 42400
rect 14476 42272 14516 42281
rect 14476 39836 14516 42232
rect 14572 41516 14612 43492
rect 14572 41467 14612 41476
rect 14572 41264 14612 41273
rect 14572 40760 14612 41224
rect 14572 40711 14612 40720
rect 14476 39500 14516 39796
rect 14476 39451 14516 39460
rect 14572 40592 14612 40601
rect 14380 38947 14420 38956
rect 14380 38828 14420 38837
rect 14380 36056 14420 38788
rect 14380 36007 14420 36016
rect 14476 38156 14516 38165
rect 14284 35848 14420 35888
rect 14380 35552 14420 35848
rect 14380 35503 14420 35512
rect 14380 35216 14420 35225
rect 14284 35048 14324 35057
rect 14284 34544 14324 35008
rect 14284 34495 14324 34504
rect 14380 34376 14420 35176
rect 14188 32059 14228 32068
rect 14284 32864 14324 32873
rect 14284 31856 14324 32824
rect 14380 32444 14420 34336
rect 14380 32276 14420 32404
rect 14380 32227 14420 32236
rect 14188 31816 14324 31856
rect 14188 31352 14228 31816
rect 14188 31303 14228 31312
rect 14284 31688 14324 31697
rect 14188 31184 14228 31193
rect 14188 30428 14228 31144
rect 14188 30092 14228 30388
rect 14188 30043 14228 30052
rect 14188 29924 14228 29933
rect 14188 29840 14228 29884
rect 14188 29789 14228 29800
rect 14284 29672 14324 31648
rect 14380 30764 14420 30773
rect 14380 30596 14420 30724
rect 14476 30680 14516 38116
rect 14572 36224 14612 40552
rect 14668 40508 14708 56176
rect 14764 54368 14804 58108
rect 14860 57812 14900 64492
rect 14956 63188 14996 68944
rect 15052 66884 15092 69280
rect 15052 66835 15092 66844
rect 15052 66716 15092 66725
rect 15052 65372 15092 66676
rect 15052 65323 15092 65332
rect 15052 64028 15092 64037
rect 15052 63524 15092 63988
rect 15052 63475 15092 63484
rect 14956 60080 14996 63148
rect 15052 63356 15092 63365
rect 15052 63104 15092 63316
rect 15052 63055 15092 63064
rect 15052 62852 15092 62861
rect 15052 62717 15092 62812
rect 14956 60031 14996 60040
rect 15052 61508 15092 61517
rect 14956 59324 14996 59333
rect 14956 59189 14996 59284
rect 14956 58736 14996 58745
rect 14956 58064 14996 58696
rect 14956 58015 14996 58024
rect 15052 58316 15092 61468
rect 15052 57980 15092 58276
rect 15052 57931 15092 57940
rect 14860 57772 14996 57812
rect 14860 57644 14900 57653
rect 14860 56300 14900 57604
rect 14860 56251 14900 56260
rect 14860 55376 14900 55385
rect 14860 54788 14900 55336
rect 14860 54739 14900 54748
rect 14764 54319 14804 54328
rect 14956 54284 14996 57772
rect 15052 56300 15092 56309
rect 15052 55040 15092 56260
rect 15052 54991 15092 55000
rect 14956 54235 14996 54244
rect 14956 47816 14996 47825
rect 14668 40459 14708 40468
rect 14764 46724 14804 46733
rect 14668 39584 14708 39593
rect 14668 38408 14708 39544
rect 14764 39164 14804 46684
rect 14956 46556 14996 47776
rect 14956 46507 14996 46516
rect 15052 45968 15092 45977
rect 14860 45716 14900 45725
rect 14860 45581 14900 45676
rect 15052 45212 15092 45928
rect 15052 45163 15092 45172
rect 15052 45044 15092 45053
rect 14860 44960 14900 44969
rect 14860 43364 14900 44920
rect 15052 44456 15092 45004
rect 15052 44407 15092 44416
rect 15052 44204 15092 44213
rect 14956 44036 14996 44045
rect 14956 43901 14996 43996
rect 15052 43700 15092 44164
rect 15052 43532 15092 43660
rect 14860 43315 14900 43324
rect 14956 43492 15052 43532
rect 14764 39115 14804 39124
rect 14860 43112 14900 43121
rect 14668 38359 14708 38368
rect 14860 38156 14900 43072
rect 14956 43028 14996 43492
rect 15052 43483 15092 43492
rect 15052 43364 15092 43373
rect 15052 43196 15092 43324
rect 15052 43147 15092 43156
rect 14956 42979 14996 42988
rect 15052 42944 15092 42953
rect 15052 42692 15092 42904
rect 14860 38107 14900 38116
rect 14956 42652 15092 42692
rect 14860 37988 14900 37997
rect 14764 37904 14804 37913
rect 14668 36644 14708 36653
rect 14668 36476 14708 36604
rect 14668 36427 14708 36436
rect 14572 36184 14708 36224
rect 14572 36056 14612 36065
rect 14572 35804 14612 36016
rect 14572 35755 14612 35764
rect 14668 35216 14708 36184
rect 14764 35384 14804 37864
rect 14860 37232 14900 37948
rect 14956 37316 14996 42652
rect 15052 42524 15092 42533
rect 15052 42020 15092 42484
rect 15052 41012 15092 41980
rect 15052 40963 15092 40972
rect 15052 40760 15092 40769
rect 15052 38408 15092 40720
rect 15052 38359 15092 38368
rect 15052 38240 15092 38249
rect 15052 37484 15092 38200
rect 15052 37435 15092 37444
rect 14956 37276 15092 37316
rect 14860 36812 14900 37192
rect 14860 36224 14900 36772
rect 14860 36175 14900 36184
rect 14956 36560 14996 36569
rect 14860 35804 14900 35813
rect 14860 35669 14900 35764
rect 14860 35552 14900 35561
rect 14860 35417 14900 35512
rect 14764 35335 14804 35344
rect 14572 35176 14708 35216
rect 14572 31520 14612 35176
rect 14764 35132 14804 35141
rect 14804 35092 14900 35132
rect 14764 35083 14804 35092
rect 14668 35048 14708 35057
rect 14668 34460 14708 35008
rect 14668 34411 14708 34420
rect 14764 34544 14804 34553
rect 14764 34292 14804 34504
rect 14668 34252 14804 34292
rect 14860 34376 14900 35092
rect 14956 34880 14996 36520
rect 14956 34544 14996 34840
rect 14956 34495 14996 34504
rect 14668 31856 14708 34252
rect 14764 32696 14804 32705
rect 14764 32108 14804 32656
rect 14764 31973 14804 32068
rect 14860 32276 14900 34336
rect 14668 31816 14804 31856
rect 14572 31480 14708 31520
rect 14572 31352 14612 31361
rect 14572 30848 14612 31312
rect 14572 30799 14612 30808
rect 14476 30631 14516 30640
rect 14380 30547 14420 30556
rect 14572 30512 14612 30521
rect 14476 30428 14516 30437
rect 14188 29632 14324 29672
rect 14380 30260 14420 30269
rect 14188 24044 14228 29632
rect 14380 29000 14420 30220
rect 14476 30176 14516 30388
rect 14476 30127 14516 30136
rect 14476 29756 14516 29796
rect 14476 29672 14516 29716
rect 14476 29420 14516 29632
rect 14476 29371 14516 29380
rect 14380 28951 14420 28960
rect 14572 28748 14612 30472
rect 14668 30344 14708 31480
rect 14764 31268 14804 31816
rect 14860 31520 14900 32236
rect 14860 31471 14900 31480
rect 14764 31219 14804 31228
rect 14956 31436 14996 31445
rect 14860 31184 14900 31193
rect 14668 30295 14708 30304
rect 14764 30680 14804 30689
rect 14764 29924 14804 30640
rect 14860 30008 14900 31144
rect 14956 30092 14996 31396
rect 15052 31352 15092 37276
rect 15052 31303 15092 31312
rect 14956 30043 14996 30052
rect 15052 31184 15092 31193
rect 14860 29959 14900 29968
rect 14572 28699 14612 28708
rect 14668 29884 14804 29924
rect 14668 28412 14708 29884
rect 14764 29756 14804 29765
rect 14764 28580 14804 29716
rect 14956 29756 14996 29765
rect 14860 29672 14900 29681
rect 14860 29084 14900 29632
rect 14956 29672 14996 29716
rect 14956 29621 14996 29632
rect 14860 29035 14900 29044
rect 14956 29336 14996 29345
rect 14764 28531 14804 28540
rect 14668 28363 14708 28372
rect 14764 27992 14804 28001
rect 14380 26984 14420 26993
rect 14188 24004 14324 24044
rect 14188 23876 14228 23885
rect 14188 23708 14228 23836
rect 14188 23036 14228 23668
rect 14284 23540 14324 24004
rect 14284 23491 14324 23500
rect 14188 22987 14228 22996
rect 14284 23288 14324 23297
rect 14284 23120 14324 23248
rect 14284 22616 14324 23080
rect 14284 22567 14324 22576
rect 14380 22448 14420 26944
rect 14668 26900 14708 26995
rect 14668 26851 14708 26860
rect 14668 26732 14708 26741
rect 14572 26648 14612 26657
rect 14476 26144 14516 26153
rect 14476 26009 14516 26104
rect 14572 26060 14612 26608
rect 14668 26228 14708 26692
rect 14668 26179 14708 26188
rect 14572 26011 14612 26020
rect 14668 25388 14708 25397
rect 14572 25136 14612 25145
rect 14476 24800 14516 24809
rect 14476 24716 14516 24760
rect 14476 24665 14516 24676
rect 14476 23876 14516 23885
rect 14476 23036 14516 23836
rect 14476 22987 14516 22996
rect 14092 20131 14132 20140
rect 14188 22408 14420 22448
rect 14476 22616 14516 22625
rect 13996 19291 14036 19300
rect 14092 20012 14132 20021
rect 13900 19207 13940 19216
rect 14092 19172 14132 19972
rect 13804 19123 13844 19132
rect 13996 19132 14132 19172
rect 13612 18115 13652 18124
rect 13900 18500 13940 18509
rect 13900 17996 13940 18460
rect 13900 17947 13940 17956
rect 13900 17492 13940 17501
rect 13612 17072 13652 17081
rect 13612 16316 13652 17032
rect 13708 16988 13748 16997
rect 13708 16400 13748 16948
rect 13708 16351 13748 16360
rect 13612 14804 13652 16276
rect 13612 14132 13652 14764
rect 13612 14083 13652 14092
rect 13804 16232 13844 16241
rect 13804 14720 13844 16192
rect 13804 13964 13844 14680
rect 13804 13915 13844 13924
rect 13516 12739 13556 12748
rect 13612 13880 13652 13889
rect 13420 12403 13460 12412
rect 13516 12620 13556 12629
rect 13516 11780 13556 12580
rect 13516 10100 13556 11740
rect 13516 10051 13556 10060
rect 13324 9547 13364 9556
rect 13324 9428 13364 9437
rect 13612 9428 13652 13840
rect 13324 8756 13364 9388
rect 13324 8707 13364 8716
rect 13516 9388 13652 9428
rect 13708 12788 13748 12797
rect 13708 10436 13748 12748
rect 13324 8420 13364 8429
rect 13324 7244 13364 8380
rect 13324 6404 13364 7204
rect 13324 5984 13364 6364
rect 13324 5935 13364 5944
rect 13420 5732 13460 5741
rect 13324 5480 13364 5489
rect 13324 4976 13364 5440
rect 13324 4927 13364 4936
rect 13420 5228 13460 5692
rect 13420 4724 13460 5188
rect 13420 4675 13460 4684
rect 13516 3968 13556 9388
rect 13516 3919 13556 3928
rect 13612 9260 13652 9269
rect 13612 3548 13652 9220
rect 13708 8924 13748 10396
rect 13804 11780 13844 11789
rect 13804 10352 13844 11740
rect 13804 9428 13844 10312
rect 13900 10016 13940 17452
rect 13996 15056 14036 19132
rect 13996 15007 14036 15016
rect 14092 17576 14132 17585
rect 13996 14804 14036 14813
rect 13996 14216 14036 14764
rect 13996 13964 14036 14176
rect 13996 13915 14036 13924
rect 13996 11360 14036 11369
rect 13996 11225 14036 11320
rect 13900 9967 13940 9976
rect 13996 10268 14036 10277
rect 13804 9379 13844 9388
rect 13900 9596 13940 9605
rect 13900 9092 13940 9556
rect 13900 9043 13940 9052
rect 13708 8884 13940 8924
rect 13708 8756 13748 8765
rect 13708 8000 13748 8716
rect 13804 8756 13844 8765
rect 13804 8168 13844 8716
rect 13804 8119 13844 8128
rect 13708 7960 13844 8000
rect 13612 3499 13652 3508
rect 13708 7832 13748 7841
rect 13228 2860 13460 2900
rect 13420 2708 13460 2860
rect 13420 2659 13460 2668
rect 13612 2792 13652 2801
rect 13612 2624 13652 2752
rect 13708 2708 13748 7792
rect 13804 3044 13844 7960
rect 13900 5648 13940 8884
rect 13996 8168 14036 10228
rect 13996 8119 14036 8128
rect 13996 5732 14036 5827
rect 13996 5683 14036 5692
rect 13900 4808 13940 5608
rect 13996 5564 14036 5573
rect 13996 5429 14036 5524
rect 13900 4759 13940 4768
rect 13804 2995 13844 3004
rect 14092 2900 14132 17536
rect 14188 17492 14228 22408
rect 14380 22280 14420 22289
rect 14188 17443 14228 17452
rect 14284 21776 14324 21785
rect 14284 21524 14324 21736
rect 14284 18668 14324 21484
rect 14380 21356 14420 22240
rect 14476 21608 14516 22576
rect 14572 22280 14612 25096
rect 14668 24548 14708 25348
rect 14668 24499 14708 24508
rect 14668 23876 14708 23885
rect 14668 23036 14708 23836
rect 14668 22532 14708 22996
rect 14668 22483 14708 22492
rect 14572 22231 14612 22240
rect 14476 21568 14708 21608
rect 14668 21440 14708 21568
rect 14668 21391 14708 21400
rect 14380 21307 14420 21316
rect 14572 21356 14612 21365
rect 14476 21272 14516 21281
rect 14380 20852 14420 20861
rect 14380 20348 14420 20812
rect 14476 20516 14516 21232
rect 14476 20467 14516 20476
rect 14380 20299 14420 20308
rect 14380 20012 14420 20021
rect 14420 19972 14516 20012
rect 14380 19963 14420 19972
rect 14380 19760 14420 19769
rect 14380 19088 14420 19720
rect 14476 19508 14516 19972
rect 14476 19459 14516 19468
rect 14572 19424 14612 21316
rect 14668 21272 14708 21281
rect 14668 20936 14708 21232
rect 14668 20264 14708 20896
rect 14668 20012 14708 20224
rect 14764 20180 14804 27952
rect 14764 20131 14804 20140
rect 14860 27992 14900 28001
rect 14764 20012 14804 20021
rect 14668 19972 14764 20012
rect 14764 19963 14804 19972
rect 14572 19375 14612 19384
rect 14668 19844 14708 19853
rect 14668 19256 14708 19804
rect 14764 19760 14804 19769
rect 14764 19424 14804 19720
rect 14764 19375 14804 19384
rect 14380 19039 14420 19048
rect 14572 19216 14708 19256
rect 14284 16988 14324 18628
rect 14572 17660 14612 19216
rect 14860 17996 14900 27952
rect 14956 25388 14996 29296
rect 15052 29000 15092 31144
rect 15052 28951 15092 28960
rect 14956 25339 14996 25348
rect 15052 28748 15092 28757
rect 14956 24632 14996 24641
rect 14956 24497 14996 24592
rect 14956 23792 14996 23801
rect 14956 23204 14996 23752
rect 14956 23155 14996 23164
rect 15052 23060 15092 28708
rect 15148 27656 15188 76924
rect 15244 73460 15284 81628
rect 15340 80408 15380 81964
rect 15340 80359 15380 80368
rect 15340 79820 15380 79829
rect 15340 76712 15380 79780
rect 15340 76124 15380 76672
rect 15340 76075 15380 76084
rect 15340 75704 15380 75713
rect 15340 75284 15380 75664
rect 15340 74696 15380 75244
rect 15340 74647 15380 74656
rect 15340 74444 15380 74453
rect 15340 74309 15380 74404
rect 15436 74276 15476 93640
rect 16300 93620 16340 94816
rect 16492 94856 16532 94865
rect 16492 94604 16532 94816
rect 16588 94688 16628 96688
rect 16588 94639 16628 94648
rect 16492 94555 16532 94564
rect 16780 94604 16820 96688
rect 16972 95024 17012 96688
rect 17164 95108 17204 96688
rect 17356 95612 17396 96688
rect 17356 95563 17396 95572
rect 17164 95068 17396 95108
rect 17356 95024 17396 95068
rect 16972 94984 17204 95024
rect 17164 94940 17204 94984
rect 17356 94975 17396 94984
rect 17164 94891 17204 94900
rect 16780 94555 16820 94564
rect 17068 94856 17108 94865
rect 16972 94184 17012 94193
rect 16972 94049 17012 94144
rect 16588 93932 16628 93941
rect 16588 93797 16628 93892
rect 16204 93580 16340 93620
rect 16396 93764 16436 93773
rect 15532 92504 15572 92513
rect 15532 86540 15572 92464
rect 16012 92420 16052 92429
rect 15628 90404 15668 90413
rect 15628 87968 15668 90364
rect 15628 87919 15668 87928
rect 15532 85868 15572 86500
rect 15532 83684 15572 85828
rect 15724 86288 15764 86297
rect 15628 85112 15668 85121
rect 15628 84692 15668 85072
rect 15628 84356 15668 84652
rect 15628 84307 15668 84316
rect 15724 85028 15764 86248
rect 15724 84272 15764 84988
rect 15820 85700 15860 85709
rect 15820 85112 15860 85660
rect 15820 84356 15860 85072
rect 16012 84776 16052 92380
rect 16108 90152 16148 90161
rect 16108 88892 16148 90112
rect 16108 88843 16148 88852
rect 16012 84727 16052 84736
rect 16108 84860 16148 84869
rect 16108 84608 16148 84820
rect 15820 84307 15860 84316
rect 16012 84568 16148 84608
rect 15724 83852 15764 84232
rect 15724 83803 15764 83812
rect 16012 83684 16052 84568
rect 15532 83644 15764 83684
rect 15628 83516 15668 83525
rect 15628 83012 15668 83476
rect 15532 82972 15668 83012
rect 15532 80576 15572 82972
rect 15628 82844 15668 82853
rect 15628 82004 15668 82804
rect 15628 81955 15668 81964
rect 15532 80072 15572 80536
rect 15628 81752 15668 81761
rect 15628 80408 15668 81712
rect 15724 81752 15764 83644
rect 15916 83600 15956 83609
rect 15724 81332 15764 81712
rect 15820 83516 15860 83525
rect 15820 81500 15860 83476
rect 15916 83012 15956 83560
rect 16012 83516 16052 83644
rect 16204 83540 16244 93580
rect 16300 89060 16340 89069
rect 16300 88925 16340 89020
rect 16012 83467 16052 83476
rect 16108 83500 16244 83540
rect 16300 84188 16340 84197
rect 16300 83768 16340 84148
rect 15916 82972 16052 83012
rect 15916 82844 15956 82853
rect 15916 81836 15956 82804
rect 16012 82676 16052 82972
rect 16012 82627 16052 82636
rect 16108 82676 16148 83500
rect 16108 82627 16148 82636
rect 16204 82760 16244 82769
rect 15916 81787 15956 81796
rect 16012 82004 16052 82013
rect 15820 81451 15860 81460
rect 15724 81283 15764 81292
rect 15628 80156 15668 80368
rect 15916 80492 15956 80501
rect 15628 80116 15764 80156
rect 15532 80032 15668 80072
rect 15628 79232 15668 80032
rect 15532 79192 15628 79232
rect 15532 77216 15572 79192
rect 15628 79183 15668 79192
rect 15628 79064 15668 79075
rect 15628 78980 15668 79024
rect 15628 78931 15668 78940
rect 15532 77167 15572 77176
rect 15628 78224 15668 78233
rect 15628 77468 15668 78184
rect 15724 78224 15764 80116
rect 15820 79820 15860 79915
rect 15820 79771 15860 79780
rect 15724 78175 15764 78184
rect 15820 79568 15860 79577
rect 15724 77972 15764 77981
rect 15724 77636 15764 77932
rect 15724 77587 15764 77596
rect 15820 77552 15860 79528
rect 15820 77503 15860 77512
rect 15628 76460 15668 77428
rect 15628 76411 15668 76420
rect 15724 77468 15764 77477
rect 15532 75788 15572 75797
rect 15532 74444 15572 75748
rect 15628 75200 15668 75209
rect 15628 74528 15668 75160
rect 15628 74479 15668 74488
rect 15532 74395 15572 74404
rect 15628 74360 15668 74369
rect 15436 74236 15572 74276
rect 15436 73940 15476 73949
rect 15244 73420 15380 73460
rect 15244 73268 15284 73277
rect 15244 73016 15284 73228
rect 15244 72967 15284 72976
rect 15244 72428 15284 72437
rect 15244 69236 15284 72388
rect 15244 68648 15284 69196
rect 15244 68599 15284 68608
rect 15340 71420 15380 73420
rect 15244 67724 15284 67733
rect 15244 66968 15284 67684
rect 15244 66919 15284 66928
rect 15244 66800 15284 66809
rect 15244 64364 15284 66760
rect 15340 66212 15380 71380
rect 15436 71588 15476 73900
rect 15436 71168 15476 71548
rect 15532 71672 15572 74236
rect 15628 74024 15668 74320
rect 15628 73975 15668 73984
rect 15628 73520 15668 73529
rect 15628 73016 15668 73480
rect 15628 72967 15668 72976
rect 15532 71504 15572 71632
rect 15532 71455 15572 71464
rect 15628 71840 15668 71849
rect 15532 71336 15572 71347
rect 15532 71252 15572 71296
rect 15532 71203 15572 71212
rect 15436 71119 15476 71128
rect 15436 70412 15476 70421
rect 15436 67808 15476 70372
rect 15532 69740 15572 69749
rect 15532 69236 15572 69700
rect 15532 69187 15572 69196
rect 15436 67759 15476 67768
rect 15532 68480 15572 68489
rect 15532 67892 15572 68440
rect 15340 65624 15380 66172
rect 15340 65575 15380 65584
rect 15436 67472 15476 67481
rect 15436 65456 15476 67432
rect 15244 64315 15284 64324
rect 15340 65416 15476 65456
rect 15244 63692 15284 63701
rect 15244 63557 15284 63652
rect 15340 63188 15380 65416
rect 15436 65288 15476 65297
rect 15436 64280 15476 65248
rect 15436 64231 15476 64240
rect 15244 63148 15380 63188
rect 15436 63944 15476 63953
rect 15244 62684 15284 63148
rect 15436 63104 15476 63904
rect 15244 62635 15284 62644
rect 15340 63064 15476 63104
rect 15532 63188 15572 67852
rect 15628 66212 15668 71800
rect 15724 71756 15764 77428
rect 15820 76964 15860 76973
rect 15820 76040 15860 76924
rect 15820 75991 15860 76000
rect 15820 74108 15860 74117
rect 15820 73772 15860 74068
rect 15820 73723 15860 73732
rect 15916 73688 15956 80452
rect 16012 75284 16052 81964
rect 16204 81416 16244 82720
rect 16204 81367 16244 81376
rect 16300 80324 16340 83728
rect 16300 80275 16340 80284
rect 16300 79736 16340 79745
rect 16204 79232 16244 79241
rect 16108 78224 16148 78233
rect 16108 78056 16148 78184
rect 16108 78007 16148 78016
rect 16108 77804 16148 77813
rect 16108 77468 16148 77764
rect 16108 77419 16148 77428
rect 16204 75368 16244 79192
rect 16300 78980 16340 79696
rect 16300 78931 16340 78940
rect 16300 78560 16340 78569
rect 16300 77384 16340 78520
rect 16300 77335 16340 77344
rect 16396 76376 16436 93724
rect 17068 90572 17108 94816
rect 17452 94856 17492 94865
rect 17452 94520 17492 94816
rect 17452 94471 17492 94480
rect 17356 94184 17396 94193
rect 17356 93680 17396 94144
rect 17356 93631 17396 93640
rect 17452 93932 17492 93941
rect 17452 93620 17492 93892
rect 17548 93848 17588 96688
rect 17548 93799 17588 93808
rect 17644 94856 17684 94865
rect 17452 93580 17588 93620
rect 17068 90523 17108 90532
rect 17260 90320 17300 90329
rect 17164 89732 17204 89741
rect 16780 89564 16820 89573
rect 16780 88892 16820 89524
rect 16588 88052 16628 88061
rect 16588 87380 16628 88012
rect 16588 87331 16628 87340
rect 16492 85952 16532 85961
rect 16492 82340 16532 85912
rect 16684 85700 16724 85709
rect 16492 82291 16532 82300
rect 16588 84440 16628 84449
rect 16492 82088 16532 82097
rect 16492 79904 16532 82048
rect 16492 79820 16532 79864
rect 16492 79771 16532 79780
rect 16492 79652 16532 79661
rect 16492 78476 16532 79612
rect 16492 78427 16532 78436
rect 16492 78308 16532 78317
rect 16492 77888 16532 78268
rect 16588 78140 16628 84400
rect 16684 83684 16724 85660
rect 16684 82004 16724 83644
rect 16780 82088 16820 88852
rect 16972 86456 17012 86465
rect 16876 84860 16916 84869
rect 16876 84725 16916 84820
rect 16780 82039 16820 82048
rect 16876 84524 16916 84533
rect 16684 81955 16724 81964
rect 16780 81920 16820 81929
rect 16588 78091 16628 78100
rect 16684 81836 16724 81845
rect 16492 77839 16532 77848
rect 16684 77804 16724 81796
rect 16780 81164 16820 81880
rect 16780 81115 16820 81124
rect 16780 80660 16820 80669
rect 16780 80492 16820 80620
rect 16780 80443 16820 80452
rect 16684 77755 16724 77764
rect 16780 80324 16820 80333
rect 16204 75319 16244 75328
rect 16300 76336 16436 76376
rect 16684 77468 16724 77477
rect 16012 75235 16052 75244
rect 16108 75200 16148 75209
rect 16108 74696 16148 75160
rect 16108 74647 16148 74656
rect 15916 73460 15956 73648
rect 16108 74528 16148 74537
rect 15916 73420 16052 73460
rect 15916 72932 15956 72941
rect 15724 71707 15764 71716
rect 15820 72260 15860 72269
rect 15820 71588 15860 72220
rect 15724 71548 15860 71588
rect 15724 70748 15764 71548
rect 15724 70699 15764 70708
rect 15820 71420 15860 71429
rect 15724 70580 15764 70589
rect 15724 66296 15764 70540
rect 15820 68396 15860 71380
rect 15820 68347 15860 68356
rect 15724 66247 15764 66256
rect 15820 67556 15860 67565
rect 15820 66968 15860 67516
rect 15628 66163 15668 66172
rect 15820 66212 15860 66928
rect 15820 66163 15860 66172
rect 15724 66128 15764 66137
rect 15244 62432 15284 62527
rect 15244 62383 15284 62392
rect 15244 62264 15284 62273
rect 15244 55712 15284 62224
rect 15340 55880 15380 63064
rect 15436 62936 15476 62945
rect 15436 61676 15476 62896
rect 15532 62432 15572 63148
rect 15532 62383 15572 62392
rect 15628 65456 15668 65465
rect 15436 61627 15476 61636
rect 15532 60164 15572 60173
rect 15436 60080 15476 60089
rect 15436 59324 15476 60040
rect 15532 59492 15572 60124
rect 15532 59443 15572 59452
rect 15436 59284 15572 59324
rect 15436 59156 15476 59165
rect 15436 57140 15476 59116
rect 15436 57091 15476 57100
rect 15340 55831 15380 55840
rect 15436 56300 15476 56309
rect 15244 55672 15380 55712
rect 15244 54116 15284 54125
rect 15244 53276 15284 54076
rect 15340 53300 15380 55672
rect 15436 55628 15476 56260
rect 15436 55579 15476 55588
rect 15340 53260 15476 53300
rect 15244 52184 15284 53236
rect 15244 52135 15284 52144
rect 15340 51596 15380 51605
rect 15340 51092 15380 51556
rect 15340 51043 15380 51052
rect 15340 50084 15380 50093
rect 15340 48740 15380 50044
rect 15340 48691 15380 48700
rect 15340 46304 15380 46313
rect 15340 45716 15380 46264
rect 15340 45667 15380 45676
rect 15340 45548 15380 45557
rect 15244 45464 15284 45473
rect 15244 43280 15284 45424
rect 15340 43532 15380 45508
rect 15340 43364 15380 43492
rect 15340 43315 15380 43324
rect 15244 43231 15284 43240
rect 15436 43220 15476 53260
rect 15532 51680 15572 59284
rect 15628 54116 15668 65416
rect 15724 65372 15764 66088
rect 15724 65323 15764 65332
rect 15820 66044 15860 66053
rect 15724 64700 15764 64709
rect 15724 64565 15764 64660
rect 15724 63944 15764 63953
rect 15724 63356 15764 63904
rect 15724 63307 15764 63316
rect 15820 63020 15860 66004
rect 15916 64028 15956 72892
rect 16012 71000 16052 73420
rect 16108 71420 16148 74488
rect 16108 71371 16148 71380
rect 16204 73520 16244 73529
rect 16012 70960 16148 71000
rect 16012 70832 16052 70841
rect 16012 70160 16052 70792
rect 16012 70111 16052 70120
rect 16108 70244 16148 70960
rect 16012 69908 16052 69917
rect 16108 69908 16148 70204
rect 16052 69868 16148 69908
rect 16012 69859 16052 69868
rect 15916 63979 15956 63988
rect 16012 69152 16052 69161
rect 15916 63860 15956 63869
rect 15916 63356 15956 63820
rect 16012 63608 16052 69112
rect 16204 68564 16244 73480
rect 16300 70496 16340 76336
rect 16588 75452 16628 75461
rect 16396 75284 16436 75293
rect 16436 75244 16532 75284
rect 16396 75235 16436 75244
rect 16396 74528 16436 74539
rect 16396 74444 16436 74488
rect 16396 74395 16436 74404
rect 16396 73940 16436 73949
rect 16396 73772 16436 73900
rect 16396 73723 16436 73732
rect 16492 73940 16532 75244
rect 16396 73520 16436 73529
rect 16396 72260 16436 73480
rect 16396 72211 16436 72220
rect 16396 71588 16436 71597
rect 16396 71453 16436 71548
rect 16300 70447 16340 70456
rect 16396 71336 16436 71345
rect 16396 70328 16436 71296
rect 16396 70279 16436 70288
rect 16492 68648 16532 73900
rect 16588 70580 16628 75412
rect 16684 72176 16724 77428
rect 16780 75284 16820 80284
rect 16780 75235 16820 75244
rect 16684 72136 16820 72176
rect 16684 72008 16724 72017
rect 16684 71420 16724 71968
rect 16684 71371 16724 71380
rect 16588 70531 16628 70540
rect 16684 71168 16724 71177
rect 16588 70412 16628 70421
rect 16588 69320 16628 70372
rect 16588 69271 16628 69280
rect 16396 68608 16492 68648
rect 16204 68524 16340 68564
rect 16204 68396 16244 68405
rect 16108 68312 16148 68321
rect 16108 67388 16148 68272
rect 16204 67892 16244 68356
rect 16204 67843 16244 67852
rect 16108 67348 16244 67388
rect 16012 63559 16052 63568
rect 16108 66716 16148 66725
rect 15916 63307 15956 63316
rect 15820 62980 15956 63020
rect 15820 62852 15860 62861
rect 15724 62348 15764 62357
rect 15820 62348 15860 62812
rect 15916 62432 15956 62980
rect 15916 62383 15956 62392
rect 16012 62936 16052 62945
rect 15764 62308 15860 62348
rect 16012 62348 16052 62896
rect 15724 62299 15764 62308
rect 16012 62299 16052 62308
rect 15916 62264 15956 62273
rect 15820 62180 15860 62189
rect 15724 61844 15764 61853
rect 15724 57308 15764 61804
rect 15820 61592 15860 62140
rect 15820 61543 15860 61552
rect 15916 60248 15956 62224
rect 15916 60199 15956 60208
rect 16012 61676 16052 61685
rect 15820 60080 15860 60089
rect 15820 58064 15860 60040
rect 15916 60080 15956 60089
rect 15916 59828 15956 60040
rect 15916 59779 15956 59788
rect 15916 59576 15956 59585
rect 15916 58736 15956 59536
rect 16012 59324 16052 61636
rect 16012 59275 16052 59284
rect 15916 58687 15956 58696
rect 16012 58904 16052 58913
rect 16012 58652 16052 58864
rect 15820 58015 15860 58024
rect 15916 58400 15956 58409
rect 15724 57259 15764 57268
rect 15628 54067 15668 54076
rect 15724 57140 15764 57149
rect 15724 54788 15764 57100
rect 15820 56384 15860 56393
rect 15820 55628 15860 56344
rect 15820 55579 15860 55588
rect 15724 53948 15764 54748
rect 15628 53276 15668 53285
rect 15628 53141 15668 53236
rect 15724 52604 15764 53908
rect 15820 54032 15860 54041
rect 15820 53897 15860 53992
rect 15724 52555 15764 52564
rect 15532 51640 15668 51680
rect 15340 43180 15476 43220
rect 15532 51008 15572 51017
rect 15532 48824 15572 50968
rect 15628 50420 15668 51640
rect 15628 50371 15668 50380
rect 15916 50336 15956 58360
rect 16012 56300 16052 58612
rect 16108 58400 16148 66676
rect 16204 61760 16244 67348
rect 16300 66884 16340 68524
rect 16300 66835 16340 66844
rect 16396 66380 16436 68608
rect 16492 68599 16532 68608
rect 16588 69152 16628 69161
rect 16588 68228 16628 69112
rect 16588 68179 16628 68188
rect 16492 68144 16532 68153
rect 16492 67640 16532 68104
rect 16492 67591 16532 67600
rect 16588 67724 16628 67733
rect 16588 67304 16628 67684
rect 16684 67472 16724 71128
rect 16684 67423 16724 67432
rect 16588 67264 16724 67304
rect 16588 66884 16628 66893
rect 16300 66340 16436 66380
rect 16492 66632 16532 66641
rect 16300 65372 16340 66340
rect 16396 66212 16436 66221
rect 16396 65540 16436 66172
rect 16492 65960 16532 66592
rect 16492 65911 16532 65920
rect 16396 65491 16436 65500
rect 16492 65792 16532 65801
rect 16300 65323 16340 65332
rect 16396 65120 16436 65129
rect 16396 64616 16436 65080
rect 16396 64567 16436 64576
rect 16396 63860 16436 63869
rect 16300 63524 16340 63533
rect 16300 61760 16340 63484
rect 16396 62432 16436 63820
rect 16396 62383 16436 62392
rect 16492 63860 16532 65752
rect 16492 62264 16532 63820
rect 16492 62215 16532 62224
rect 16300 61720 16532 61760
rect 16204 60500 16244 61720
rect 16204 60451 16244 60460
rect 16300 61592 16340 61601
rect 16204 60248 16244 60343
rect 16204 60199 16244 60208
rect 16108 58351 16148 58360
rect 16204 60080 16244 60089
rect 16204 58820 16244 60040
rect 16300 59072 16340 61552
rect 16396 61508 16436 61517
rect 16396 61088 16436 61468
rect 16396 61039 16436 61048
rect 16396 60164 16436 60173
rect 16396 59576 16436 60124
rect 16396 59527 16436 59536
rect 16300 59023 16340 59032
rect 16396 59324 16436 59333
rect 16012 55544 16052 56260
rect 16012 55495 16052 55504
rect 16108 58232 16148 58241
rect 16012 54116 16052 54125
rect 16012 53360 16052 54076
rect 16012 53311 16052 53320
rect 15916 50287 15956 50296
rect 15820 50084 15860 50093
rect 15244 43028 15284 43037
rect 15244 42692 15284 42988
rect 15244 41852 15284 42652
rect 15244 41348 15284 41812
rect 15244 41299 15284 41308
rect 15244 41096 15284 41105
rect 15244 37988 15284 41056
rect 15244 37939 15284 37948
rect 15244 37484 15284 37493
rect 15244 36476 15284 37444
rect 15244 36056 15284 36436
rect 15244 35636 15284 36016
rect 15244 35587 15284 35596
rect 15244 35384 15284 35393
rect 15244 34796 15284 35344
rect 15244 34747 15284 34756
rect 15244 34460 15284 34469
rect 15244 34325 15284 34420
rect 15244 33452 15284 33461
rect 15244 32948 15284 33412
rect 15244 32899 15284 32908
rect 15244 32108 15284 32117
rect 15244 27824 15284 32068
rect 15244 27775 15284 27784
rect 15148 27616 15284 27656
rect 14764 17956 14900 17996
rect 14956 23020 15092 23060
rect 15148 27488 15188 27497
rect 14572 17611 14612 17620
rect 14668 17744 14708 17755
rect 14668 17660 14708 17704
rect 14668 17611 14708 17620
rect 14284 16232 14324 16948
rect 14284 16183 14324 16192
rect 14380 17576 14420 17585
rect 14380 15812 14420 17536
rect 14380 15763 14420 15772
rect 14476 16988 14516 16997
rect 14476 16316 14516 16948
rect 14668 16988 14708 16997
rect 14668 16853 14708 16948
rect 14284 15560 14324 15569
rect 14188 15476 14228 15485
rect 14188 15224 14228 15436
rect 14188 13292 14228 15184
rect 14284 14972 14324 15520
rect 14284 14923 14324 14932
rect 14284 14804 14324 14813
rect 14476 14804 14516 16276
rect 14324 14764 14516 14804
rect 14668 16736 14708 16745
rect 14668 14972 14708 16696
rect 14284 14755 14324 14764
rect 14476 14636 14516 14645
rect 14380 14552 14420 14561
rect 14188 13243 14228 13252
rect 14284 14132 14324 14141
rect 14188 12032 14228 12041
rect 14188 11528 14228 11992
rect 14188 11479 14228 11488
rect 14284 9596 14324 14092
rect 14380 12704 14420 14512
rect 14380 12655 14420 12664
rect 14380 12452 14420 12461
rect 14380 11864 14420 12412
rect 14380 11815 14420 11824
rect 14380 11696 14420 11705
rect 14476 11696 14516 14596
rect 14668 14636 14708 14932
rect 14668 14587 14708 14596
rect 14764 12980 14804 17956
rect 14860 17828 14900 17837
rect 14860 16736 14900 17788
rect 14860 16687 14900 16696
rect 14860 16316 14900 16325
rect 14860 15728 14900 16276
rect 14860 15679 14900 15688
rect 14956 15560 14996 23020
rect 15052 22784 15092 22793
rect 15052 22364 15092 22744
rect 15052 19424 15092 22324
rect 15052 19375 15092 19384
rect 15052 19256 15092 19265
rect 15052 19004 15092 19216
rect 15052 18955 15092 18964
rect 15052 17912 15092 17921
rect 15052 16484 15092 17872
rect 15052 16435 15092 16444
rect 14668 12940 14804 12980
rect 14860 15520 14996 15560
rect 14860 14132 14900 15520
rect 14668 11864 14708 12940
rect 14668 11815 14708 11824
rect 14764 12872 14804 12881
rect 14764 12452 14804 12832
rect 14420 11656 14516 11696
rect 14380 11108 14420 11656
rect 14380 11059 14420 11068
rect 14476 11528 14516 11537
rect 14476 10940 14516 11488
rect 14284 9547 14324 9556
rect 14380 10772 14420 10781
rect 14380 9512 14420 10732
rect 14380 9463 14420 9472
rect 14476 10184 14516 10900
rect 14284 9428 14324 9437
rect 14188 9176 14228 9185
rect 14188 8756 14228 9136
rect 14188 8707 14228 8716
rect 14188 8588 14228 8597
rect 14188 6152 14228 8548
rect 14284 7076 14324 9388
rect 14284 7027 14324 7036
rect 14380 9344 14420 9353
rect 14188 6112 14324 6152
rect 14284 5732 14324 6112
rect 14284 5683 14324 5692
rect 14188 4892 14228 4901
rect 14188 4757 14228 4852
rect 13708 2659 13748 2668
rect 13996 2876 14036 2885
rect 14092 2876 14324 2900
rect 14092 2860 14284 2876
rect 13612 2575 13652 2584
rect 13996 2624 14036 2836
rect 14284 2827 14324 2836
rect 13996 2575 14036 2584
rect 14380 2624 14420 9304
rect 14476 9344 14516 10144
rect 14476 6404 14516 9304
rect 14476 6355 14516 6364
rect 14572 10100 14612 10109
rect 14476 6236 14516 6245
rect 14476 5816 14516 6196
rect 14476 5767 14516 5776
rect 14380 2575 14420 2584
rect 13036 1903 13076 1912
rect 13324 2456 13364 2465
rect 13132 1616 13172 1625
rect 12844 400 12980 440
rect 12940 80 12980 400
rect 13132 80 13172 1576
rect 13324 80 13364 2416
rect 13708 2456 13748 2465
rect 13420 1952 13460 1961
rect 13420 1817 13460 1912
rect 13516 1616 13556 1625
rect 13516 80 13556 1576
rect 13708 80 13748 2416
rect 14092 2456 14132 2465
rect 13900 2036 13940 2045
rect 13900 80 13940 1996
rect 14092 80 14132 2416
rect 14476 2456 14516 2465
rect 14188 2372 14228 2381
rect 14188 1952 14228 2332
rect 14188 1903 14228 1912
rect 14284 1616 14324 1625
rect 14284 80 14324 1576
rect 14476 80 14516 2416
rect 14572 1952 14612 10060
rect 14764 9512 14804 12412
rect 14764 9463 14804 9472
rect 14860 8924 14900 14092
rect 14956 15392 14996 15401
rect 14956 12032 14996 15352
rect 15148 14972 15188 27448
rect 15244 21776 15284 27616
rect 15340 27488 15380 43180
rect 15436 43112 15476 43121
rect 15436 42776 15476 43072
rect 15436 42727 15476 42736
rect 15436 42524 15476 42533
rect 15436 42104 15476 42484
rect 15436 42055 15476 42064
rect 15436 41936 15476 41945
rect 15436 41180 15476 41896
rect 15436 41131 15476 41140
rect 15436 41012 15476 41021
rect 15436 40877 15476 40972
rect 15436 40760 15476 40769
rect 15436 40424 15476 40720
rect 15436 40375 15476 40384
rect 15436 40004 15476 40013
rect 15436 38828 15476 39964
rect 15436 38240 15476 38788
rect 15436 38191 15476 38200
rect 15436 38072 15476 38081
rect 15436 37937 15476 38032
rect 15436 35972 15476 35981
rect 15436 35837 15476 35932
rect 15436 34292 15476 34301
rect 15436 33704 15476 34252
rect 15436 33655 15476 33664
rect 15532 31940 15572 48784
rect 15628 49580 15668 49589
rect 15628 47228 15668 49540
rect 15628 47093 15668 47188
rect 15724 49244 15764 49253
rect 15628 44204 15668 44213
rect 15628 44069 15668 44164
rect 15628 43448 15668 43457
rect 15628 42944 15668 43408
rect 15628 42895 15668 42904
rect 15628 42692 15668 42701
rect 15628 42188 15668 42652
rect 15628 41936 15668 42148
rect 15628 41887 15668 41896
rect 15628 41600 15668 41609
rect 15628 40676 15668 41560
rect 15628 40627 15668 40636
rect 15628 40508 15668 40517
rect 15628 38912 15668 40468
rect 15628 38863 15668 38872
rect 15724 38576 15764 49204
rect 15820 48992 15860 50044
rect 15820 48943 15860 48952
rect 15820 48740 15860 48835
rect 15820 48691 15860 48700
rect 15820 48572 15860 48581
rect 16108 48572 16148 58192
rect 16204 57812 16244 58780
rect 16204 57763 16244 57772
rect 16300 58568 16340 58577
rect 16300 57224 16340 58528
rect 16300 56384 16340 57184
rect 16300 56335 16340 56344
rect 16300 56216 16340 56225
rect 16300 55628 16340 56176
rect 16300 55579 16340 55588
rect 16300 54872 16340 54881
rect 16204 54032 16244 54041
rect 16204 53276 16244 53992
rect 16204 53227 16244 53236
rect 16204 51260 16244 51269
rect 16204 51092 16244 51220
rect 16300 51176 16340 54832
rect 16396 52184 16436 59284
rect 16492 59156 16532 61720
rect 16588 59324 16628 66844
rect 16684 65876 16724 67264
rect 16780 66044 16820 72136
rect 16876 69068 16916 84484
rect 16972 84356 17012 86416
rect 16972 84307 17012 84316
rect 17068 85196 17108 85205
rect 16972 84020 17012 84029
rect 16972 83684 17012 83980
rect 16972 83635 17012 83644
rect 17068 83516 17108 85156
rect 17164 83600 17204 89692
rect 17260 89480 17300 90280
rect 17260 88892 17300 89440
rect 17260 87380 17300 88852
rect 17260 87331 17300 87340
rect 17356 89564 17396 89573
rect 17260 86624 17300 86633
rect 17260 84020 17300 86584
rect 17260 83971 17300 83980
rect 17164 83551 17204 83560
rect 17260 83852 17300 83861
rect 17068 83467 17108 83476
rect 17260 83516 17300 83812
rect 17260 83467 17300 83476
rect 17164 83432 17204 83441
rect 16972 82844 17012 82853
rect 16972 82172 17012 82804
rect 16972 82123 17012 82132
rect 16972 82004 17012 82013
rect 16972 80576 17012 81964
rect 16972 80527 17012 80536
rect 17068 81920 17108 81929
rect 16972 78476 17012 78485
rect 16972 78341 17012 78436
rect 16972 76796 17012 76805
rect 16972 75872 17012 76756
rect 17068 76292 17108 81880
rect 17164 79148 17204 83392
rect 17260 83096 17300 83105
rect 17260 81248 17300 83056
rect 17260 81199 17300 81208
rect 17356 80156 17396 89524
rect 17452 87464 17492 87473
rect 17452 87329 17492 87424
rect 17452 86456 17492 86465
rect 17452 85952 17492 86416
rect 17452 85903 17492 85912
rect 17452 85784 17492 85793
rect 17452 80240 17492 85744
rect 17548 81500 17588 93580
rect 17644 89564 17684 94816
rect 17740 94604 17780 96688
rect 17836 94604 17876 94613
rect 17740 94564 17836 94604
rect 17836 94555 17876 94564
rect 17740 94436 17780 94445
rect 17740 94184 17780 94396
rect 17740 94135 17780 94144
rect 17932 94100 17972 96688
rect 18028 95612 18068 95621
rect 18028 94688 18068 95572
rect 18124 94940 18164 96688
rect 18124 94891 18164 94900
rect 18220 94856 18260 94865
rect 18220 94721 18260 94816
rect 18124 94688 18164 94697
rect 18028 94648 18124 94688
rect 18124 94639 18164 94648
rect 18220 94520 18260 94529
rect 18124 94184 18164 94193
rect 18028 94100 18068 94109
rect 17932 94060 18028 94100
rect 18028 94051 18068 94060
rect 18124 94049 18164 94144
rect 17740 93932 17780 93941
rect 17740 93797 17780 93892
rect 18220 93764 18260 94480
rect 18316 93848 18356 96688
rect 18316 93799 18356 93808
rect 18412 94856 18452 94865
rect 18220 93715 18260 93724
rect 18316 93680 18356 93689
rect 18412 93680 18452 94816
rect 18356 93640 18452 93680
rect 18316 93631 18356 93640
rect 18508 93596 18548 96688
rect 18604 94856 18644 94865
rect 18604 94520 18644 94816
rect 18604 94471 18644 94480
rect 18604 94184 18644 94193
rect 18604 94049 18644 94144
rect 18508 93547 18548 93556
rect 18700 93512 18740 96688
rect 18796 94856 18836 94865
rect 18796 94721 18836 94816
rect 18892 94688 18932 96688
rect 19084 94856 19124 96688
rect 19084 94807 19124 94816
rect 19276 94772 19316 96688
rect 19468 95024 19508 96688
rect 20048 95276 20416 95285
rect 20088 95236 20130 95276
rect 20170 95236 20212 95276
rect 20252 95236 20294 95276
rect 20334 95236 20376 95276
rect 20048 95227 20416 95236
rect 19468 94984 19604 95024
rect 19468 94856 19508 94865
rect 19276 94732 19412 94772
rect 18892 94648 19316 94688
rect 18808 94520 19176 94529
rect 18848 94480 18890 94520
rect 18930 94480 18972 94520
rect 19012 94480 19054 94520
rect 19094 94480 19136 94520
rect 18808 94471 19176 94480
rect 19084 94268 19124 94277
rect 18988 94184 19028 94193
rect 18700 93463 18740 93472
rect 18796 93848 18836 93857
rect 18796 93344 18836 93808
rect 18988 93764 19028 94144
rect 18988 93715 19028 93724
rect 18796 93295 18836 93304
rect 18988 93344 19028 93353
rect 18988 93209 19028 93304
rect 19084 93260 19124 94228
rect 19084 93211 19124 93220
rect 18700 93176 18740 93185
rect 18700 93041 18740 93136
rect 18808 93008 19176 93017
rect 18848 92968 18890 93008
rect 18930 92968 18972 93008
rect 19012 92968 19054 93008
rect 19094 92968 19136 93008
rect 18808 92959 19176 92968
rect 19276 92840 19316 94648
rect 19276 92791 19316 92800
rect 19180 92672 19220 92681
rect 19180 92420 19220 92632
rect 19180 92371 19220 92380
rect 19372 92084 19412 94732
rect 19468 92840 19508 94816
rect 19564 94268 19604 94984
rect 19948 94940 19988 94949
rect 19756 94856 19796 94865
rect 19564 94219 19604 94228
rect 19660 94772 19700 94781
rect 19564 93932 19604 93941
rect 19564 93428 19604 93892
rect 19660 93596 19700 94732
rect 19756 94100 19796 94816
rect 19756 94051 19796 94060
rect 19852 94184 19892 94193
rect 19852 94049 19892 94144
rect 19660 93547 19700 93556
rect 19756 93932 19796 93941
rect 19756 93428 19796 93892
rect 19564 93388 19700 93428
rect 19468 92791 19508 92800
rect 19564 93260 19604 93269
rect 19468 92672 19508 92681
rect 19468 92537 19508 92632
rect 19372 92035 19412 92044
rect 19564 91832 19604 93220
rect 19660 92588 19700 93388
rect 19756 93379 19796 93388
rect 19852 93764 19892 93773
rect 19660 92539 19700 92548
rect 19756 92672 19796 92681
rect 19756 92537 19796 92632
rect 19564 91783 19604 91792
rect 19756 91832 19796 91841
rect 19756 91697 19796 91792
rect 18508 91580 18548 91589
rect 17644 89515 17684 89524
rect 18028 89648 18068 89657
rect 17644 89396 17684 89405
rect 17644 87380 17684 89356
rect 17932 88220 17972 88229
rect 17644 87331 17684 87340
rect 17836 87716 17876 87725
rect 17740 87212 17780 87221
rect 17644 87128 17684 87137
rect 17644 83768 17684 87088
rect 17740 86540 17780 87172
rect 17836 87128 17876 87676
rect 17836 87079 17876 87088
rect 17740 86405 17780 86500
rect 17932 86456 17972 88180
rect 17932 86407 17972 86416
rect 17932 86120 17972 86129
rect 17836 85784 17876 85793
rect 17836 85649 17876 85744
rect 17932 84860 17972 86080
rect 17836 84820 17972 84860
rect 17740 84188 17780 84228
rect 17740 84104 17780 84148
rect 17740 83852 17780 84064
rect 17836 84020 17876 84820
rect 17836 83971 17876 83980
rect 17932 84692 17972 84701
rect 17932 84356 17972 84652
rect 17740 83812 17876 83852
rect 17836 83768 17876 83812
rect 17644 83728 17780 83768
rect 17548 81451 17588 81460
rect 17644 83600 17684 83609
rect 17548 80576 17588 80585
rect 17548 80441 17588 80536
rect 17452 80200 17588 80240
rect 17356 80116 17492 80156
rect 17164 78224 17204 79108
rect 17164 78175 17204 78184
rect 17260 79736 17300 79745
rect 17068 76243 17108 76252
rect 17164 78056 17204 78065
rect 17164 77804 17204 78016
rect 16972 75823 17012 75832
rect 17068 75956 17108 75965
rect 17068 75821 17108 75916
rect 17068 75284 17108 75293
rect 16876 69019 16916 69028
rect 16972 75200 17012 75209
rect 16972 69236 17012 75160
rect 17068 74948 17108 75244
rect 17068 74899 17108 74908
rect 17068 74696 17108 74705
rect 17068 74192 17108 74656
rect 17068 74143 17108 74152
rect 17164 73520 17204 77764
rect 17260 77300 17300 79696
rect 17260 77251 17300 77260
rect 17356 75956 17396 75965
rect 17260 75788 17300 75797
rect 17260 74528 17300 75748
rect 17356 74696 17396 75916
rect 17356 74647 17396 74656
rect 17260 74479 17300 74488
rect 17164 73471 17204 73480
rect 17068 73352 17108 73361
rect 17068 70916 17108 73312
rect 17164 72848 17204 72857
rect 17164 72428 17204 72808
rect 17260 72764 17300 72773
rect 17300 72724 17396 72764
rect 17260 72715 17300 72724
rect 17260 72428 17300 72437
rect 17164 72388 17260 72428
rect 17260 72379 17300 72388
rect 17164 72092 17204 72101
rect 17164 71588 17204 72052
rect 17164 71539 17204 71548
rect 17260 71504 17300 71513
rect 17260 71369 17300 71464
rect 17068 70876 17204 70916
rect 16876 68900 16916 68909
rect 16876 66884 16916 68860
rect 16876 66835 16916 66844
rect 16780 65995 16820 66004
rect 16684 65836 16820 65876
rect 16684 65372 16724 65381
rect 16684 64868 16724 65332
rect 16684 64819 16724 64828
rect 16780 64868 16820 65836
rect 16780 64819 16820 64828
rect 16876 65288 16916 65297
rect 16780 64700 16820 64709
rect 16684 64112 16724 64121
rect 16684 63608 16724 64072
rect 16684 63559 16724 63568
rect 16684 62432 16724 62441
rect 16684 62348 16724 62392
rect 16684 60836 16724 62308
rect 16684 60787 16724 60796
rect 16588 59275 16628 59284
rect 16684 60500 16724 60509
rect 16492 59116 16628 59156
rect 16396 52135 16436 52144
rect 16492 57812 16532 57821
rect 16492 51680 16532 57772
rect 16588 55460 16628 59116
rect 16684 58232 16724 60460
rect 16684 58183 16724 58192
rect 16684 57896 16724 57907
rect 16684 57812 16724 57856
rect 16684 57763 16724 57772
rect 16780 57812 16820 64660
rect 16876 62096 16916 65248
rect 16972 64700 17012 69196
rect 17068 70748 17108 70757
rect 17068 69236 17108 70708
rect 17164 70412 17204 70876
rect 17164 70363 17204 70372
rect 17260 70748 17300 70757
rect 17068 69187 17108 69196
rect 17164 70244 17204 70253
rect 17260 70244 17300 70708
rect 17356 70412 17396 72724
rect 17356 70363 17396 70372
rect 17260 70204 17396 70244
rect 17164 69992 17204 70204
rect 16972 64651 17012 64660
rect 17068 69068 17108 69077
rect 17068 64616 17108 69028
rect 17164 67052 17204 69952
rect 17260 68228 17300 68237
rect 17260 67640 17300 68188
rect 17260 67591 17300 67600
rect 17164 67003 17204 67012
rect 17260 67472 17300 67481
rect 17068 64567 17108 64576
rect 17164 66884 17204 66893
rect 16876 62047 16916 62056
rect 16972 64532 17012 64541
rect 16972 63188 17012 64492
rect 16780 57763 16820 57772
rect 16876 61928 16916 61937
rect 16876 61592 16916 61888
rect 16876 58652 16916 61552
rect 16972 60080 17012 63148
rect 17068 63020 17108 63029
rect 17068 61844 17108 62980
rect 17068 61795 17108 61804
rect 16972 60031 17012 60040
rect 17068 61676 17108 61687
rect 17068 61592 17108 61636
rect 17068 60164 17108 61552
rect 16876 57308 16916 58612
rect 16972 59912 17012 59921
rect 16972 57980 17012 59872
rect 16972 57931 17012 57940
rect 16876 57259 16916 57268
rect 16972 57644 17012 57653
rect 16876 56888 16916 56897
rect 16588 55411 16628 55420
rect 16780 56300 16820 56309
rect 16780 55040 16820 56260
rect 16876 55628 16916 56848
rect 16876 55579 16916 55588
rect 16780 54991 16820 55000
rect 16684 54704 16724 54713
rect 16588 54116 16628 54144
rect 16684 54116 16724 54664
rect 16628 54076 16724 54116
rect 16588 54067 16628 54076
rect 16684 53276 16724 54076
rect 16684 53227 16724 53236
rect 16972 53360 17012 57604
rect 17068 56384 17108 60124
rect 17068 56335 17108 56344
rect 17164 57140 17204 66844
rect 17260 65120 17300 67432
rect 17356 66716 17396 70204
rect 17452 70160 17492 80116
rect 17548 77720 17588 80200
rect 17644 78056 17684 83560
rect 17740 83012 17780 83728
rect 17836 83719 17876 83728
rect 17740 82963 17780 82972
rect 17836 83600 17876 83609
rect 17740 82844 17780 82853
rect 17836 82844 17876 83560
rect 17932 83516 17972 84316
rect 17932 83467 17972 83476
rect 17780 82804 17876 82844
rect 17740 78980 17780 82804
rect 17932 82760 17972 82769
rect 17740 78931 17780 78940
rect 17836 82720 17932 82760
rect 17836 80324 17876 82720
rect 17932 82711 17972 82720
rect 18028 81920 18068 89608
rect 18124 89564 18164 89573
rect 18124 88052 18164 89524
rect 18124 88003 18164 88012
rect 18220 88136 18260 88145
rect 18220 88001 18260 88096
rect 18508 88052 18548 91540
rect 18808 91496 19176 91505
rect 18848 91456 18890 91496
rect 18930 91456 18972 91496
rect 19012 91456 19054 91496
rect 19094 91456 19136 91496
rect 18808 91447 19176 91456
rect 19660 91160 19700 91169
rect 19276 90320 19316 90329
rect 18808 89984 19176 89993
rect 18848 89944 18890 89984
rect 18930 89944 18972 89984
rect 19012 89944 19054 89984
rect 19094 89944 19136 89984
rect 18808 89935 19176 89944
rect 18988 88892 19028 88903
rect 18604 88808 18644 88817
rect 18604 88673 18644 88768
rect 18988 88808 19028 88852
rect 18988 88759 19028 88768
rect 18316 87380 18356 87389
rect 18124 87128 18164 87137
rect 18124 86540 18164 87088
rect 18124 86120 18164 86500
rect 18124 86071 18164 86080
rect 18316 86540 18356 87340
rect 18412 87296 18452 87305
rect 18412 86624 18452 87256
rect 18412 86575 18452 86584
rect 18220 85700 18260 85709
rect 18124 85616 18164 85625
rect 18124 85028 18164 85576
rect 18124 84440 18164 84988
rect 18124 84391 18164 84400
rect 18124 84272 18164 84281
rect 18124 83852 18164 84232
rect 18124 83803 18164 83812
rect 18124 83684 18164 83693
rect 18124 82088 18164 83644
rect 18124 82039 18164 82048
rect 18028 81880 18164 81920
rect 18028 81752 18068 81761
rect 17932 81248 17972 81257
rect 17932 81113 17972 81208
rect 17644 78007 17684 78016
rect 17548 77671 17588 77680
rect 17836 77552 17876 80284
rect 17932 80996 17972 81005
rect 17932 78644 17972 80956
rect 18028 80492 18068 81712
rect 18028 80443 18068 80452
rect 18124 80576 18164 81880
rect 18220 81584 18260 85660
rect 18316 82760 18356 86500
rect 18508 85868 18548 88012
rect 18700 88640 18740 88649
rect 18604 87380 18644 87389
rect 18604 87128 18644 87340
rect 18604 87079 18644 87088
rect 18604 86960 18644 86969
rect 18604 86372 18644 86920
rect 18700 86540 18740 88600
rect 18808 88472 19176 88481
rect 18848 88432 18890 88472
rect 18930 88432 18972 88472
rect 19012 88432 19054 88472
rect 19094 88432 19136 88472
rect 18808 88423 19176 88432
rect 18796 88304 18836 88313
rect 18796 87128 18836 88264
rect 19276 88136 19316 90280
rect 19468 89648 19508 89657
rect 19372 88808 19412 88817
rect 19372 88724 19412 88768
rect 19372 88673 19412 88684
rect 19276 88096 19412 88136
rect 19276 87968 19316 87977
rect 19276 87380 19316 87928
rect 19276 87331 19316 87340
rect 18796 87079 18836 87088
rect 18808 86960 19176 86969
rect 19372 86960 19412 88096
rect 18848 86920 18890 86960
rect 18930 86920 18972 86960
rect 19012 86920 19054 86960
rect 19094 86920 19136 86960
rect 18808 86911 19176 86920
rect 19276 86920 19412 86960
rect 18700 86491 18740 86500
rect 18796 86456 18836 86465
rect 18604 86332 18740 86372
rect 18508 85819 18548 85828
rect 18316 82711 18356 82720
rect 18412 85784 18452 85793
rect 18316 82592 18356 82601
rect 18316 82004 18356 82552
rect 18316 81955 18356 81964
rect 18220 81535 18260 81544
rect 18316 81836 18356 81845
rect 17932 78595 17972 78604
rect 17836 77503 17876 77512
rect 17932 78476 17972 78485
rect 17932 78140 17972 78436
rect 18028 78392 18068 78401
rect 18028 78257 18068 78352
rect 17644 77468 17684 77477
rect 17644 77333 17684 77428
rect 17644 76544 17684 76553
rect 17644 76040 17684 76504
rect 17548 75788 17588 75797
rect 17548 75653 17588 75748
rect 17548 75536 17588 75545
rect 17548 73856 17588 75496
rect 17644 74528 17684 76000
rect 17836 75956 17876 75965
rect 17644 74479 17684 74488
rect 17740 75872 17780 75881
rect 17740 74276 17780 75832
rect 17836 74696 17876 75916
rect 17836 74647 17876 74656
rect 17836 74528 17876 74537
rect 17836 74393 17876 74488
rect 17740 74227 17780 74236
rect 17932 74360 17972 78100
rect 18124 76208 18164 80536
rect 18220 81416 18260 81425
rect 18220 79148 18260 81376
rect 18316 81332 18356 81796
rect 18316 80996 18356 81292
rect 18316 80947 18356 80956
rect 18220 79099 18260 79108
rect 18316 80660 18356 80669
rect 18220 78980 18260 78989
rect 18220 76796 18260 78940
rect 18220 76747 18260 76756
rect 18028 75032 18068 75041
rect 18028 74528 18068 74992
rect 18028 74479 18068 74488
rect 18124 74360 18164 76168
rect 17836 74024 17876 74033
rect 17644 73940 17684 73949
rect 17836 73940 17876 73984
rect 17684 73900 17876 73940
rect 17644 73891 17684 73900
rect 17932 73856 17972 74320
rect 17548 73807 17588 73816
rect 17740 73816 17972 73856
rect 18028 74320 18164 74360
rect 18220 76292 18260 76301
rect 18220 75956 18260 76252
rect 17548 72764 17588 72773
rect 17548 72344 17588 72724
rect 17548 72295 17588 72304
rect 17644 72764 17684 72773
rect 17644 72260 17684 72724
rect 17644 72211 17684 72220
rect 17644 72092 17684 72101
rect 17548 70916 17588 70925
rect 17548 70781 17588 70876
rect 17452 70111 17492 70120
rect 17548 70496 17588 70505
rect 17548 69908 17588 70456
rect 17548 69859 17588 69868
rect 17548 68900 17588 68909
rect 17548 68396 17588 68860
rect 17356 66667 17396 66676
rect 17452 67976 17492 67985
rect 17260 65071 17300 65080
rect 17356 66548 17396 66557
rect 17356 65372 17396 66508
rect 17356 65036 17396 65332
rect 17356 64987 17396 64996
rect 17260 64616 17300 64625
rect 17260 63860 17300 64576
rect 17260 63811 17300 63820
rect 17356 63944 17396 63953
rect 17260 63524 17300 63533
rect 17260 62684 17300 63484
rect 17260 62635 17300 62644
rect 17260 62516 17300 62525
rect 17260 62381 17300 62476
rect 17260 62096 17300 62105
rect 17260 60584 17300 62056
rect 17356 61844 17396 63904
rect 17356 61795 17396 61804
rect 17356 61508 17396 61517
rect 17356 61373 17396 61468
rect 17260 60535 17300 60544
rect 17260 60332 17300 60341
rect 17260 58736 17300 60292
rect 17260 58687 17300 58696
rect 17356 60164 17396 60173
rect 17068 56216 17108 56225
rect 17068 56081 17108 56176
rect 17164 55544 17204 57100
rect 16492 51631 16532 51640
rect 16300 51136 16532 51176
rect 16204 50168 16244 51052
rect 16204 50119 16244 50128
rect 16300 51008 16340 51017
rect 16300 50084 16340 50968
rect 16396 50336 16436 50345
rect 16396 50201 16436 50296
rect 16300 50035 16340 50044
rect 16204 49664 16244 49673
rect 16204 49529 16244 49624
rect 15860 48532 16148 48572
rect 16300 49412 16340 49421
rect 16300 48992 16340 49372
rect 15820 48523 15860 48532
rect 16204 48068 16244 48077
rect 15820 47984 15860 47993
rect 15820 47480 15860 47944
rect 16204 47933 16244 48028
rect 16300 47984 16340 48952
rect 16396 48908 16436 48917
rect 16396 48740 16436 48868
rect 16396 48068 16436 48700
rect 16396 48019 16436 48028
rect 16300 47935 16340 47944
rect 15820 47431 15860 47440
rect 15820 47228 15860 47237
rect 15820 46892 15860 47188
rect 15820 42944 15860 46852
rect 16492 45296 16532 51136
rect 16780 51092 16820 51101
rect 16780 50957 16820 51052
rect 16876 50252 16916 50261
rect 16972 50252 17012 53320
rect 17068 55292 17108 55301
rect 17068 52688 17108 55252
rect 17164 54788 17204 55504
rect 17164 54739 17204 54748
rect 17260 58568 17300 58577
rect 17260 54704 17300 58528
rect 17356 58400 17396 60124
rect 17452 60080 17492 67936
rect 17548 60164 17588 68356
rect 17644 65288 17684 72052
rect 17740 67976 17780 73816
rect 17836 73520 17876 73529
rect 17836 71420 17876 73480
rect 17836 71371 17876 71380
rect 17932 72848 17972 72857
rect 17836 71252 17876 71261
rect 17836 70496 17876 71212
rect 17932 70748 17972 72808
rect 18028 72596 18068 74320
rect 18028 72547 18068 72556
rect 18124 73772 18164 73781
rect 18124 72344 18164 73732
rect 18028 72304 18164 72344
rect 18028 71252 18068 72304
rect 18028 71203 18068 71212
rect 18124 72176 18164 72185
rect 18124 71336 18164 72136
rect 17932 70699 17972 70708
rect 18028 70664 18068 70673
rect 17836 69236 17876 70456
rect 17932 70580 17972 70589
rect 17932 69992 17972 70540
rect 17932 69943 17972 69952
rect 17836 69187 17876 69196
rect 17932 69488 17972 69497
rect 17740 67927 17780 67936
rect 17740 66884 17780 66893
rect 17740 66548 17780 66844
rect 17740 66499 17780 66508
rect 17836 66716 17876 66725
rect 17836 66212 17876 66676
rect 17836 66163 17876 66172
rect 17644 65239 17684 65248
rect 17740 66128 17780 66137
rect 17740 65204 17780 66088
rect 17932 66044 17972 69448
rect 18028 67136 18068 70624
rect 18028 67087 18068 67096
rect 18124 69824 18164 71296
rect 18220 70748 18260 75916
rect 18316 75200 18356 80620
rect 18412 80324 18452 85744
rect 18604 85532 18644 85541
rect 18508 84860 18548 84869
rect 18508 84440 18548 84820
rect 18508 84391 18548 84400
rect 18508 84272 18548 84281
rect 18508 82844 18548 84232
rect 18508 82795 18548 82804
rect 18508 82592 18548 82601
rect 18508 81416 18548 82552
rect 18604 81752 18644 85492
rect 18700 85280 18740 86332
rect 18796 86321 18836 86416
rect 18808 85448 19176 85457
rect 18848 85408 18890 85448
rect 18930 85408 18972 85448
rect 19012 85408 19054 85448
rect 19094 85408 19136 85448
rect 18808 85399 19176 85408
rect 18700 85240 18836 85280
rect 18700 84356 18740 84365
rect 18700 83684 18740 84316
rect 18796 84104 18836 85240
rect 18796 84055 18836 84064
rect 18808 83936 19176 83945
rect 18848 83896 18890 83936
rect 18930 83896 18972 83936
rect 19012 83896 19054 83936
rect 19094 83896 19136 83936
rect 18808 83887 19176 83896
rect 18700 83635 18740 83644
rect 18796 83768 18836 83777
rect 18796 83540 18836 83728
rect 18988 83768 19028 83777
rect 18988 83600 19028 83728
rect 18988 83551 19028 83560
rect 18604 81703 18644 81712
rect 18700 83500 18836 83540
rect 18508 81367 18548 81376
rect 18604 81332 18644 81427
rect 18604 81283 18644 81292
rect 18412 80275 18452 80284
rect 18508 81248 18548 81257
rect 18508 80156 18548 81208
rect 18316 75151 18356 75160
rect 18412 80116 18548 80156
rect 18604 81080 18644 81089
rect 18316 74864 18356 74873
rect 18316 72848 18356 74824
rect 18412 74444 18452 80116
rect 18508 79568 18548 79577
rect 18508 76460 18548 79528
rect 18604 76880 18644 81040
rect 18604 76831 18644 76840
rect 18508 76411 18548 76420
rect 18604 76712 18644 76721
rect 18508 75872 18548 75881
rect 18508 75284 18548 75832
rect 18508 75235 18548 75244
rect 18412 74395 18452 74404
rect 18508 75032 18548 75041
rect 18508 73856 18548 74992
rect 18508 73807 18548 73816
rect 18604 73772 18644 76672
rect 18604 73460 18644 73732
rect 18316 72799 18356 72808
rect 18412 73420 18644 73460
rect 18412 72932 18452 73420
rect 18316 72680 18356 72689
rect 18316 72260 18356 72640
rect 18316 72211 18356 72220
rect 18412 72092 18452 72892
rect 18604 73352 18644 73361
rect 18508 72848 18548 72857
rect 18508 72428 18548 72808
rect 18508 72379 18548 72388
rect 18604 72512 18644 73312
rect 18604 72260 18644 72472
rect 18220 70699 18260 70708
rect 18316 72052 18452 72092
rect 18508 72220 18644 72260
rect 18316 70580 18356 72052
rect 18124 69152 18164 69784
rect 18124 66800 18164 69112
rect 18028 66296 18068 66305
rect 18028 66161 18068 66256
rect 17740 65155 17780 65164
rect 17836 66004 17972 66044
rect 17548 60115 17588 60124
rect 17644 65120 17684 65129
rect 17452 60031 17492 60040
rect 17548 59996 17588 60005
rect 17452 59912 17492 59921
rect 17452 58736 17492 59872
rect 17452 58687 17492 58696
rect 17548 58652 17588 59956
rect 17548 58603 17588 58612
rect 17356 58351 17396 58360
rect 17644 56132 17684 65080
rect 17740 65036 17780 65045
rect 17740 60920 17780 64996
rect 17836 63380 17876 66004
rect 18028 64448 18068 64457
rect 17836 63340 17972 63380
rect 17836 63104 17876 63113
rect 17836 61508 17876 63064
rect 17932 61928 17972 63340
rect 18028 63188 18068 64408
rect 18124 63440 18164 66760
rect 18220 70540 18356 70580
rect 18412 71924 18452 71933
rect 18412 71420 18452 71884
rect 18508 71672 18548 72220
rect 18508 71623 18548 71632
rect 18604 72092 18644 72101
rect 18220 64700 18260 70540
rect 18316 69992 18356 70001
rect 18316 69320 18356 69952
rect 18412 69908 18452 71380
rect 18508 71504 18548 71513
rect 18604 71504 18644 72052
rect 18548 71464 18644 71504
rect 18508 70748 18548 71464
rect 18508 70699 18548 70708
rect 18604 70664 18644 70673
rect 18412 69859 18452 69868
rect 18508 70580 18548 70589
rect 18412 69320 18452 69329
rect 18316 69280 18412 69320
rect 18412 69271 18452 69280
rect 18412 69068 18452 69077
rect 18412 67136 18452 69028
rect 18412 67087 18452 67096
rect 18412 66884 18452 66893
rect 18220 64028 18260 64660
rect 18220 63979 18260 63988
rect 18316 66800 18356 66809
rect 18316 66212 18356 66760
rect 18124 63391 18164 63400
rect 18220 63860 18260 63869
rect 18028 63139 18068 63148
rect 18124 63272 18164 63281
rect 18028 62936 18068 62945
rect 18028 62600 18068 62896
rect 18028 62551 18068 62560
rect 18124 62348 18164 63232
rect 18220 63188 18260 63820
rect 18316 63524 18356 66172
rect 18412 63692 18452 66844
rect 18508 65540 18548 70540
rect 18604 66044 18644 70624
rect 18604 65995 18644 66004
rect 18508 65491 18548 65500
rect 18508 65372 18548 65381
rect 18508 64112 18548 65332
rect 18508 64063 18548 64072
rect 18412 63643 18452 63652
rect 18508 63944 18548 63953
rect 18316 63484 18452 63524
rect 18220 63139 18260 63148
rect 18316 63356 18356 63365
rect 17932 61879 17972 61888
rect 18028 62308 18164 62348
rect 18220 62348 18260 62357
rect 18028 61760 18068 62308
rect 17836 61459 17876 61468
rect 17932 61720 18068 61760
rect 18124 62180 18164 62189
rect 17932 61004 17972 61720
rect 18124 61676 18164 62140
rect 18124 61627 18164 61636
rect 17932 60955 17972 60964
rect 18028 61592 18068 61601
rect 17740 60871 17780 60880
rect 17932 60500 17972 60509
rect 17836 60164 17876 60173
rect 17740 60080 17780 60089
rect 17740 58652 17780 60040
rect 17836 58820 17876 60124
rect 17836 58771 17876 58780
rect 17740 58612 17876 58652
rect 17740 56384 17780 56393
rect 17740 56249 17780 56344
rect 17260 54655 17300 54664
rect 17548 56092 17684 56132
rect 17068 52639 17108 52648
rect 17164 53612 17204 53621
rect 16916 50212 17012 50252
rect 16876 50203 16916 50212
rect 17068 50084 17108 50093
rect 16876 49580 16916 49589
rect 16204 44792 16244 44801
rect 15820 42895 15860 42904
rect 15916 44372 15956 44381
rect 15820 42524 15860 42533
rect 15820 42389 15860 42484
rect 15820 42104 15860 42113
rect 15820 42020 15860 42064
rect 15820 41969 15860 41980
rect 15820 41852 15860 41861
rect 15820 41717 15860 41812
rect 15820 41516 15860 41525
rect 15820 41264 15860 41476
rect 15820 41215 15860 41224
rect 15916 41180 15956 44332
rect 16204 44204 16244 44752
rect 16492 44372 16532 45256
rect 16492 44323 16532 44332
rect 16780 47900 16820 47909
rect 16012 44164 16204 44204
rect 16012 42692 16052 44164
rect 16204 44155 16244 44164
rect 16780 43700 16820 47860
rect 16300 43448 16340 43457
rect 16012 42643 16052 42652
rect 16108 43364 16148 43373
rect 16108 42104 16148 43324
rect 16300 42692 16340 43408
rect 16108 42055 16148 42064
rect 16204 42272 16244 42281
rect 16108 41936 16148 41945
rect 16108 41684 16148 41896
rect 15916 41131 15956 41140
rect 16012 41348 16052 41357
rect 15916 41012 15956 41021
rect 15820 40508 15860 40519
rect 15820 40424 15860 40468
rect 15820 39752 15860 40384
rect 15820 39703 15860 39712
rect 15628 38536 15764 38576
rect 15820 38996 15860 39005
rect 15628 34964 15668 38536
rect 15724 38408 15764 38417
rect 15724 38273 15764 38368
rect 15820 38072 15860 38956
rect 15820 38023 15860 38032
rect 15724 36980 15764 36989
rect 15724 36140 15764 36940
rect 15724 36091 15764 36100
rect 15820 36896 15860 36905
rect 15820 35972 15860 36856
rect 15916 36812 15956 40972
rect 16012 40844 16052 41308
rect 16108 41180 16148 41644
rect 16108 41131 16148 41140
rect 16204 41432 16244 42232
rect 16300 42020 16340 42652
rect 16300 41971 16340 41980
rect 16396 42692 16436 42701
rect 16204 41012 16244 41392
rect 16204 40963 16244 40972
rect 16300 41852 16340 41861
rect 16012 40795 16052 40804
rect 16300 39080 16340 41812
rect 16204 39040 16340 39080
rect 16012 38744 16052 38753
rect 16012 38240 16052 38704
rect 16012 38191 16052 38200
rect 15916 36772 16052 36812
rect 15916 36644 15956 36653
rect 15916 36509 15956 36604
rect 15820 35923 15860 35932
rect 15628 34915 15668 34924
rect 15820 35636 15860 35645
rect 15532 31891 15572 31900
rect 15628 34796 15668 34805
rect 15436 31520 15476 31529
rect 15436 30092 15476 31480
rect 15436 30008 15476 30052
rect 15436 29959 15476 29968
rect 15532 31352 15572 31361
rect 15436 29672 15476 29681
rect 15436 29537 15476 29632
rect 15532 29000 15572 31312
rect 15628 29252 15668 34756
rect 15724 33536 15764 33545
rect 15724 30512 15764 33496
rect 15820 32864 15860 35596
rect 15916 35636 15956 35647
rect 15916 35552 15956 35596
rect 15916 35503 15956 35512
rect 15916 35132 15956 35143
rect 15916 35048 15956 35092
rect 15916 34999 15956 35008
rect 15916 34544 15956 34553
rect 15916 34376 15956 34504
rect 15916 34327 15956 34336
rect 16012 34460 16052 36772
rect 15820 32024 15860 32824
rect 15820 31975 15860 31984
rect 15916 33536 15956 33545
rect 15916 32024 15956 33496
rect 15724 30463 15764 30472
rect 15820 31268 15860 31277
rect 15628 29203 15668 29212
rect 15724 30344 15764 30353
rect 15724 29168 15764 30304
rect 15820 29924 15860 31228
rect 15916 30680 15956 31984
rect 15916 30631 15956 30640
rect 15820 29756 15860 29884
rect 15820 29707 15860 29716
rect 15724 29119 15764 29128
rect 15916 29672 15956 29681
rect 15916 29504 15956 29632
rect 15436 28960 15572 29000
rect 15724 29000 15764 29009
rect 15436 27572 15476 28960
rect 15436 27523 15476 27532
rect 15532 28832 15572 28841
rect 15340 27439 15380 27448
rect 15436 26228 15476 26237
rect 15436 26144 15476 26188
rect 15436 26093 15476 26104
rect 15340 25976 15380 25985
rect 15340 25304 15380 25936
rect 15340 25255 15380 25264
rect 15436 25724 15476 25733
rect 15340 24716 15380 24725
rect 15340 23036 15380 24676
rect 15436 24632 15476 25684
rect 15436 24583 15476 24592
rect 15340 22987 15380 22996
rect 15244 21727 15284 21736
rect 15340 22868 15380 22877
rect 15340 21608 15380 22828
rect 15340 21440 15380 21568
rect 15340 21391 15380 21400
rect 15436 21524 15476 21533
rect 15244 21356 15284 21365
rect 15244 20180 15284 21316
rect 15340 21104 15380 21113
rect 15340 20768 15380 21064
rect 15340 20719 15380 20728
rect 15244 20131 15284 20140
rect 15340 20600 15380 20609
rect 15244 20012 15284 20021
rect 15244 19508 15284 19972
rect 15340 19760 15380 20560
rect 15340 19711 15380 19720
rect 15436 19592 15476 21484
rect 15436 19543 15476 19552
rect 15244 19459 15284 19468
rect 15436 19424 15476 19433
rect 15340 18500 15380 18509
rect 15340 18365 15380 18460
rect 15244 18332 15284 18341
rect 15244 18080 15284 18292
rect 15244 18031 15284 18040
rect 15340 17996 15380 18005
rect 15244 17828 15284 17837
rect 15244 17492 15284 17788
rect 15244 17443 15284 17452
rect 15148 14923 15188 14932
rect 15148 14804 15188 14813
rect 15052 14636 15092 14645
rect 15052 12452 15092 14596
rect 15052 12403 15092 12412
rect 14956 11983 14996 11992
rect 14956 11780 14996 11789
rect 14956 11192 14996 11740
rect 14956 11143 14996 11152
rect 14860 8875 14900 8884
rect 15052 9512 15092 9521
rect 14668 8840 14708 8849
rect 14668 7244 14708 8800
rect 15052 8336 15092 9472
rect 15148 8924 15188 14764
rect 15244 13880 15284 13889
rect 15244 12704 15284 13840
rect 15244 12655 15284 12664
rect 15340 11444 15380 17956
rect 15436 16988 15476 19384
rect 15436 15476 15476 16948
rect 15436 15427 15476 15436
rect 15436 14804 15476 14813
rect 15436 13796 15476 14764
rect 15436 13747 15476 13756
rect 15436 13460 15476 13469
rect 15436 13325 15476 13420
rect 15340 10100 15380 11404
rect 15340 10051 15380 10060
rect 15436 12452 15476 12461
rect 15436 11864 15476 12412
rect 15340 9680 15380 9689
rect 15340 9545 15380 9640
rect 15148 8875 15188 8884
rect 15052 7412 15092 8296
rect 15340 8084 15380 8093
rect 15436 8084 15476 11824
rect 15380 8044 15476 8084
rect 15340 7664 15380 8044
rect 15340 7615 15380 7624
rect 15052 7363 15092 7372
rect 14668 7195 14708 7204
rect 15340 6992 15380 7001
rect 15052 6488 15092 6497
rect 14764 5984 14804 5993
rect 14764 5732 14804 5944
rect 15052 5900 15092 6448
rect 15340 6404 15380 6952
rect 15340 6355 15380 6364
rect 15052 5851 15092 5860
rect 14764 5683 14804 5692
rect 15052 5732 15092 5741
rect 14668 5648 14708 5657
rect 14668 5060 14708 5608
rect 15052 5597 15092 5692
rect 14668 5011 14708 5020
rect 14668 4892 14708 4901
rect 14668 4556 14708 4852
rect 14668 4507 14708 4516
rect 14764 2624 14804 2633
rect 14764 2489 14804 2584
rect 15532 2624 15572 28792
rect 15724 28832 15764 28960
rect 15724 28783 15764 28792
rect 15820 28916 15860 28925
rect 15820 28580 15860 28876
rect 15820 28531 15860 28540
rect 15820 28412 15860 28421
rect 15820 27572 15860 28372
rect 15724 27152 15764 27247
rect 15724 27103 15764 27112
rect 15724 26900 15764 26909
rect 15724 25388 15764 26860
rect 15724 25339 15764 25348
rect 15628 24548 15668 24557
rect 15628 17996 15668 24508
rect 15724 24044 15764 24053
rect 15724 23909 15764 24004
rect 15724 23792 15764 23801
rect 15724 23288 15764 23752
rect 15724 23239 15764 23248
rect 15724 21524 15764 21533
rect 15724 21020 15764 21484
rect 15820 21356 15860 27532
rect 15820 21307 15860 21316
rect 15724 19340 15764 20980
rect 15820 21104 15860 21113
rect 15820 20852 15860 21064
rect 15820 20803 15860 20812
rect 15724 19291 15764 19300
rect 15820 20180 15860 20189
rect 15820 19256 15860 20140
rect 15820 19207 15860 19216
rect 15820 19088 15860 19097
rect 15628 17947 15668 17956
rect 15724 18584 15764 18593
rect 15628 17744 15668 17753
rect 15628 17660 15668 17704
rect 15628 14804 15668 17620
rect 15628 14755 15668 14764
rect 15628 14216 15668 14225
rect 15628 14048 15668 14176
rect 15628 13999 15668 14008
rect 15628 12452 15668 12461
rect 15628 10268 15668 12412
rect 15628 10219 15668 10228
rect 15628 9260 15668 9269
rect 15628 8840 15668 9220
rect 15628 6320 15668 8800
rect 15628 6271 15668 6280
rect 15628 5900 15668 5909
rect 15628 4892 15668 5860
rect 15628 4843 15668 4852
rect 15532 2575 15572 2584
rect 14572 1903 14612 1912
rect 14860 2456 14900 2465
rect 14668 1784 14708 1793
rect 14668 80 14708 1744
rect 14860 80 14900 2416
rect 15244 2456 15284 2465
rect 15052 1616 15092 1625
rect 15052 80 15092 1576
rect 15244 80 15284 2416
rect 15340 1952 15380 1961
rect 15340 1817 15380 1912
rect 15724 1952 15764 18544
rect 15820 17828 15860 19048
rect 15820 17779 15860 17788
rect 15916 17660 15956 29464
rect 16012 27656 16052 34420
rect 16108 36728 16148 36737
rect 16108 31520 16148 36688
rect 16108 31471 16148 31480
rect 16204 31436 16244 39040
rect 16300 38912 16340 38921
rect 16300 38777 16340 38872
rect 16300 36644 16340 36653
rect 16300 36560 16340 36604
rect 16300 36509 16340 36520
rect 16300 36056 16340 36065
rect 16300 35972 16340 36016
rect 16300 35921 16340 35932
rect 16300 35804 16340 35813
rect 16300 35468 16340 35764
rect 16300 35419 16340 35428
rect 16300 35216 16340 35225
rect 16300 33620 16340 35176
rect 16300 33116 16340 33580
rect 16300 33067 16340 33076
rect 16300 32108 16340 32117
rect 16300 31772 16340 32068
rect 16300 31723 16340 31732
rect 16204 31387 16244 31396
rect 16300 31604 16340 31613
rect 16108 31268 16148 31277
rect 16108 30260 16148 31228
rect 16108 30211 16148 30220
rect 16204 31100 16244 31109
rect 16108 29420 16148 29429
rect 16108 29168 16148 29380
rect 16108 29119 16148 29128
rect 16108 29000 16148 29009
rect 16204 29000 16244 31060
rect 16300 30176 16340 31564
rect 16396 31016 16436 42652
rect 16588 42020 16628 42029
rect 16492 41684 16532 41779
rect 16492 41635 16532 41644
rect 16492 41432 16532 41441
rect 16492 41096 16532 41392
rect 16492 41047 16532 41056
rect 16492 40928 16532 40939
rect 16492 40844 16532 40888
rect 16492 40795 16532 40804
rect 16492 40508 16532 40517
rect 16492 40088 16532 40468
rect 16492 38240 16532 40048
rect 16492 38191 16532 38200
rect 16396 30848 16436 30976
rect 16396 30799 16436 30808
rect 16492 38072 16532 38081
rect 16300 30127 16340 30136
rect 16396 30512 16436 30521
rect 16396 29924 16436 30472
rect 16396 29756 16436 29884
rect 16300 29336 16340 29345
rect 16300 29168 16340 29296
rect 16300 29119 16340 29128
rect 16204 28960 16340 29000
rect 16108 27824 16148 28960
rect 16300 28496 16340 28960
rect 16300 28447 16340 28456
rect 16108 27775 16148 27784
rect 16204 28412 16244 28421
rect 16204 27656 16244 28372
rect 16012 27616 16148 27656
rect 16012 23624 16052 23633
rect 16012 21524 16052 23584
rect 16108 23288 16148 27616
rect 16204 27607 16244 27616
rect 16300 28076 16340 28085
rect 16204 26144 16244 26153
rect 16204 25556 16244 26104
rect 16204 25507 16244 25516
rect 16108 23239 16148 23248
rect 16204 25304 16244 25313
rect 16204 24800 16244 25264
rect 16012 21475 16052 21484
rect 16108 23036 16148 23045
rect 16204 23036 16244 24760
rect 16148 22996 16244 23036
rect 16012 21356 16052 21365
rect 16012 20012 16052 21316
rect 16108 20768 16148 22996
rect 16300 21692 16340 28036
rect 16396 27572 16436 29716
rect 16396 27523 16436 27532
rect 16492 26900 16532 38032
rect 16588 37484 16628 41980
rect 16684 42020 16724 42029
rect 16684 41852 16724 41980
rect 16684 41768 16724 41812
rect 16684 38408 16724 41728
rect 16780 38576 16820 43660
rect 16876 46556 16916 49540
rect 16876 40508 16916 46516
rect 16876 40459 16916 40468
rect 16972 48656 17012 48665
rect 16780 38527 16820 38536
rect 16876 39080 16916 39089
rect 16876 38996 16916 39040
rect 16684 38368 16820 38408
rect 16588 37435 16628 37444
rect 16684 38240 16724 38249
rect 16684 36980 16724 38200
rect 16684 36931 16724 36940
rect 16588 36896 16628 36905
rect 16588 36224 16628 36856
rect 16588 36175 16628 36184
rect 16780 35888 16820 38368
rect 16876 38240 16916 38956
rect 16876 37400 16916 38200
rect 16876 37351 16916 37360
rect 16780 35839 16820 35848
rect 16876 36980 16916 36989
rect 16780 35636 16820 35645
rect 16684 35300 16724 35309
rect 16588 35132 16628 35141
rect 16588 34997 16628 35092
rect 16684 35048 16724 35260
rect 16780 35132 16820 35596
rect 16780 35083 16820 35092
rect 16588 33620 16628 33631
rect 16588 33536 16628 33580
rect 16588 33487 16628 33496
rect 16588 32948 16628 32957
rect 16588 31352 16628 32908
rect 16684 32360 16724 35008
rect 16780 33620 16820 33629
rect 16780 32948 16820 33580
rect 16780 32899 16820 32908
rect 16684 32311 16724 32320
rect 16780 32612 16820 32621
rect 16780 31772 16820 32572
rect 16588 31303 16628 31312
rect 16684 31732 16820 31772
rect 16588 31184 16628 31193
rect 16588 31049 16628 31144
rect 16588 30848 16628 30857
rect 16588 28412 16628 30808
rect 16684 30092 16724 31732
rect 16780 31436 16820 31445
rect 16780 30260 16820 31396
rect 16780 30211 16820 30220
rect 16684 30052 16820 30092
rect 16684 29924 16724 29933
rect 16684 28916 16724 29884
rect 16684 28832 16724 28876
rect 16684 28752 16724 28792
rect 16588 28363 16628 28372
rect 16684 28496 16724 28505
rect 16588 27068 16628 27077
rect 16588 26933 16628 27028
rect 16492 26144 16532 26860
rect 16492 26095 16532 26104
rect 16588 26060 16628 26155
rect 16588 26011 16628 26020
rect 16684 25556 16724 28456
rect 16780 27908 16820 30052
rect 16876 28076 16916 36940
rect 16972 31352 17012 48616
rect 17068 39668 17108 50044
rect 17164 40004 17204 53572
rect 17452 53360 17492 53455
rect 17452 53311 17492 53320
rect 17260 52604 17300 52613
rect 17260 52184 17300 52564
rect 17260 51932 17300 52144
rect 17260 51883 17300 51892
rect 17452 52436 17492 52445
rect 17452 51260 17492 52396
rect 17452 51211 17492 51220
rect 17548 48824 17588 56092
rect 17836 52436 17876 58612
rect 17932 54116 17972 60460
rect 18028 59408 18068 61552
rect 18220 60920 18260 62308
rect 18220 60871 18260 60880
rect 18220 60668 18260 60677
rect 18028 59359 18068 59368
rect 18124 60164 18164 60173
rect 18028 59156 18068 59165
rect 18028 58652 18068 59116
rect 18028 58603 18068 58612
rect 18028 58484 18068 58493
rect 18028 57812 18068 58444
rect 18028 57763 18068 57772
rect 18124 57224 18164 60124
rect 18220 58904 18260 60628
rect 18316 60500 18356 63316
rect 18412 61676 18452 63484
rect 18508 63188 18548 63904
rect 18508 61844 18548 63148
rect 18604 63608 18644 63617
rect 18604 62516 18644 63568
rect 18604 62467 18644 62476
rect 18508 61795 18548 61804
rect 18604 61676 18644 61685
rect 18412 61636 18604 61676
rect 18316 60460 18452 60500
rect 18316 60080 18356 60089
rect 18316 59912 18356 60040
rect 18412 60080 18452 60460
rect 18412 60031 18452 60040
rect 18508 60164 18548 60173
rect 18316 59863 18356 59872
rect 18412 59912 18452 59921
rect 18220 58855 18260 58864
rect 18316 59744 18356 59753
rect 18220 58400 18260 58409
rect 18220 58265 18260 58360
rect 18124 55628 18164 57184
rect 18220 57896 18260 57905
rect 18220 56216 18260 57856
rect 18220 56081 18260 56176
rect 18316 56132 18356 59704
rect 18412 58568 18452 59872
rect 18412 58519 18452 58528
rect 18412 57896 18452 57905
rect 18412 57812 18452 57856
rect 18412 57761 18452 57772
rect 18508 57476 18548 60124
rect 18316 56083 18356 56092
rect 18412 57436 18548 57476
rect 18604 59324 18644 61636
rect 18124 55579 18164 55588
rect 18316 55628 18356 55637
rect 18316 54872 18356 55588
rect 18316 54823 18356 54832
rect 17932 54067 17972 54076
rect 18412 54788 18452 57436
rect 18508 57308 18548 57317
rect 18508 56300 18548 57268
rect 18508 56251 18548 56260
rect 17836 52387 17876 52396
rect 18316 53612 18356 53621
rect 17644 52352 17684 52361
rect 17644 51092 17684 52312
rect 18316 51848 18356 53572
rect 18412 52352 18452 54748
rect 18508 54620 18548 54629
rect 18508 54200 18548 54580
rect 18508 54151 18548 54160
rect 18604 54116 18644 59284
rect 18508 54032 18548 54041
rect 18508 53360 18548 53992
rect 18508 53311 18548 53320
rect 18412 52303 18452 52312
rect 18604 53276 18644 54076
rect 18604 51932 18644 53236
rect 18604 51883 18644 51892
rect 18316 51799 18356 51808
rect 17644 51043 17684 51052
rect 17644 49328 17684 49337
rect 17644 49193 17684 49288
rect 17548 48775 17588 48784
rect 18220 48908 18260 48917
rect 18220 48740 18260 48868
rect 18220 48488 18260 48700
rect 18316 48824 18356 48833
rect 18316 48656 18356 48784
rect 18316 48607 18356 48616
rect 18604 48824 18644 48833
rect 18220 48439 18260 48448
rect 18604 48404 18644 48784
rect 18604 48355 18644 48364
rect 17452 48236 17492 48245
rect 17260 48068 17300 48077
rect 17260 47480 17300 48028
rect 17260 47431 17300 47440
rect 17356 46472 17396 46481
rect 17260 46388 17300 46397
rect 17260 45632 17300 46348
rect 17260 45583 17300 45592
rect 17260 45044 17300 45053
rect 17356 45044 17396 46432
rect 17300 45004 17396 45044
rect 17260 44036 17300 45004
rect 17260 43532 17300 43996
rect 17260 43483 17300 43492
rect 17164 39955 17204 39964
rect 17260 40844 17300 40853
rect 17068 39619 17108 39628
rect 17260 39500 17300 40804
rect 17068 39460 17300 39500
rect 17068 35468 17108 39460
rect 17356 37400 17396 37409
rect 17164 37316 17204 37325
rect 17164 36560 17204 37276
rect 17356 37265 17396 37360
rect 17260 37232 17300 37241
rect 17260 37148 17300 37192
rect 17260 37097 17300 37108
rect 17356 37064 17396 37073
rect 17164 35636 17204 36520
rect 17260 36644 17300 36653
rect 17260 35804 17300 36604
rect 17260 35755 17300 35764
rect 17164 35587 17204 35596
rect 17068 35428 17204 35468
rect 17068 34460 17108 34469
rect 17068 34376 17108 34420
rect 17068 34325 17108 34336
rect 17164 32612 17204 35428
rect 17260 35216 17300 35225
rect 17260 35081 17300 35176
rect 17356 33536 17396 37024
rect 17452 35132 17492 48196
rect 18028 47228 18068 47237
rect 17548 46556 17588 46565
rect 17548 46220 17588 46516
rect 17548 45800 17588 46180
rect 17548 45751 17588 45760
rect 17740 45548 17780 45557
rect 17644 45044 17684 45053
rect 17644 44456 17684 45004
rect 17644 44407 17684 44416
rect 17740 44204 17780 45508
rect 18028 44456 18068 47188
rect 18412 46052 18452 46061
rect 18316 45800 18356 45809
rect 17740 44155 17780 44164
rect 17932 44204 17972 44213
rect 17644 44120 17684 44129
rect 17548 41432 17588 41441
rect 17548 40508 17588 41392
rect 17548 39668 17588 40468
rect 17548 39533 17588 39628
rect 17644 41096 17684 44080
rect 17836 42524 17876 42533
rect 17836 42020 17876 42484
rect 17836 41600 17876 41980
rect 17836 41551 17876 41560
rect 17644 39584 17684 41056
rect 17740 41180 17780 41189
rect 17740 39920 17780 41140
rect 17836 41012 17876 41021
rect 17836 40508 17876 40972
rect 17836 40459 17876 40468
rect 17740 39871 17780 39880
rect 17644 39332 17684 39544
rect 17644 39292 17780 39332
rect 17644 37400 17684 37409
rect 17548 37316 17588 37325
rect 17548 36812 17588 37276
rect 17548 36763 17588 36772
rect 17548 36560 17588 36569
rect 17548 36392 17588 36520
rect 17548 36343 17588 36352
rect 17644 36140 17684 37360
rect 17740 37064 17780 39292
rect 17836 37568 17876 37577
rect 17836 37433 17876 37528
rect 17740 37015 17780 37024
rect 17740 36644 17780 36653
rect 17740 36560 17780 36604
rect 17726 36520 17780 36560
rect 17726 36308 17766 36520
rect 17836 36308 17876 36317
rect 17726 36268 17780 36308
rect 17644 36091 17684 36100
rect 17452 35083 17492 35092
rect 17548 35972 17588 35981
rect 17740 35972 17780 36268
rect 17452 34964 17492 34973
rect 17452 34544 17492 34924
rect 17452 34495 17492 34504
rect 17356 33487 17396 33496
rect 17452 34208 17492 34217
rect 17452 33536 17492 34168
rect 17548 34208 17588 35932
rect 17644 35932 17780 35972
rect 17644 35300 17684 35932
rect 17644 35251 17684 35260
rect 17740 35804 17780 35813
rect 17548 34159 17588 34168
rect 17740 34124 17780 35764
rect 17836 35216 17876 36268
rect 17836 35167 17876 35176
rect 17740 34075 17780 34084
rect 17836 34964 17876 34973
rect 17836 33956 17876 34924
rect 17932 34712 17972 44164
rect 18028 41432 18068 44416
rect 18124 45716 18164 45725
rect 18124 45044 18164 45676
rect 18316 45044 18356 45760
rect 18412 45716 18452 46012
rect 18412 45212 18452 45676
rect 18412 45163 18452 45172
rect 18412 45044 18452 45053
rect 18316 45004 18412 45044
rect 18452 45004 18548 45044
rect 18124 43868 18164 45004
rect 18412 44995 18452 45004
rect 18412 44288 18452 44297
rect 18124 43532 18164 43828
rect 18124 42692 18164 43492
rect 18124 42643 18164 42652
rect 18316 44036 18356 44045
rect 18028 41383 18068 41392
rect 18220 41180 18260 41189
rect 18124 40424 18164 40433
rect 18124 40289 18164 40384
rect 18124 39752 18164 39761
rect 18124 39617 18164 39712
rect 18028 38996 18068 39005
rect 18028 36896 18068 38956
rect 18124 38828 18164 38837
rect 18124 37400 18164 38788
rect 18124 37351 18164 37360
rect 18028 36847 18068 36856
rect 18124 37232 18164 37241
rect 18124 36728 18164 37192
rect 18220 37148 18260 41140
rect 18220 37099 18260 37108
rect 18124 36679 18164 36688
rect 18220 36644 18260 36653
rect 18028 36392 18068 36401
rect 18028 35804 18068 36352
rect 18028 35132 18068 35764
rect 18028 35083 18068 35092
rect 18124 36392 18164 36401
rect 18124 34964 18164 36352
rect 18220 35384 18260 36604
rect 18316 35804 18356 43996
rect 18412 42020 18452 44248
rect 18508 43532 18548 45004
rect 18700 44456 18740 83500
rect 19084 83432 19124 83441
rect 19084 83297 19124 83392
rect 18808 82424 19176 82433
rect 18848 82384 18890 82424
rect 18930 82384 18972 82424
rect 19012 82384 19054 82424
rect 19094 82384 19136 82424
rect 18808 82375 19176 82384
rect 18988 82256 19028 82265
rect 18892 82088 18932 82097
rect 18892 81332 18932 82048
rect 18892 81283 18932 81292
rect 18988 82004 19028 82216
rect 18988 81248 19028 81964
rect 19180 82004 19220 82013
rect 19084 81500 19124 81509
rect 19084 81365 19124 81460
rect 19180 81332 19220 81964
rect 19180 81283 19220 81292
rect 18988 81199 19028 81208
rect 18808 80912 19176 80921
rect 18848 80872 18890 80912
rect 18930 80872 18972 80912
rect 19012 80872 19054 80912
rect 19094 80872 19136 80912
rect 18808 80863 19176 80872
rect 18988 80744 19028 80753
rect 18796 80492 18836 80501
rect 18796 79820 18836 80452
rect 18796 79568 18836 79780
rect 18796 79519 18836 79528
rect 18988 79568 19028 80704
rect 19084 80744 19124 80753
rect 19084 79652 19124 80704
rect 19084 79603 19124 79612
rect 18988 79519 19028 79528
rect 18808 79400 19176 79409
rect 18848 79360 18890 79400
rect 18930 79360 18972 79400
rect 19012 79360 19054 79400
rect 19094 79360 19136 79400
rect 18808 79351 19176 79360
rect 18796 79232 18836 79241
rect 18796 78392 18836 79192
rect 19180 79232 19220 79241
rect 19084 79148 19124 79157
rect 19084 78980 19124 79108
rect 18988 78812 19028 78821
rect 18796 78343 18836 78352
rect 18892 78644 18932 78653
rect 18892 78308 18932 78604
rect 18892 78259 18932 78268
rect 18796 78224 18836 78233
rect 18796 78056 18836 78184
rect 18796 78007 18836 78016
rect 18988 78056 19028 78772
rect 19084 78560 19124 78940
rect 19084 78511 19124 78520
rect 19180 78560 19220 79192
rect 19180 78511 19220 78520
rect 19180 78308 19220 78317
rect 19180 78173 19220 78268
rect 18988 78007 19028 78016
rect 19276 78056 19316 86920
rect 19372 85616 19412 85625
rect 19372 84356 19412 85576
rect 19372 84307 19412 84316
rect 19372 84188 19412 84197
rect 19372 84053 19412 84148
rect 19372 83936 19412 83945
rect 19372 82592 19412 83896
rect 19372 82543 19412 82552
rect 19372 82424 19412 82433
rect 19372 81164 19412 82384
rect 19372 81115 19412 81124
rect 19276 78007 19316 78016
rect 19372 79568 19412 79577
rect 19372 78392 19412 79528
rect 18808 77888 19176 77897
rect 18848 77848 18890 77888
rect 18930 77848 18972 77888
rect 19012 77848 19054 77888
rect 19094 77848 19136 77888
rect 18808 77839 19176 77848
rect 19276 77888 19316 77897
rect 18892 77468 18932 77477
rect 18892 76964 18932 77428
rect 18892 76915 18932 76924
rect 18808 76376 19176 76385
rect 18848 76336 18890 76376
rect 18930 76336 18972 76376
rect 19012 76336 19054 76376
rect 19094 76336 19136 76376
rect 18808 76327 19176 76336
rect 19276 76124 19316 77848
rect 19372 77636 19412 78352
rect 19372 77587 19412 77596
rect 19276 76075 19316 76084
rect 19372 77468 19412 77477
rect 18892 76040 18932 76049
rect 18796 75368 18836 75377
rect 18796 75032 18836 75328
rect 18892 75284 18932 76000
rect 18892 75235 18932 75244
rect 18796 74983 18836 74992
rect 19276 75032 19316 75041
rect 18808 74864 19176 74873
rect 18848 74824 18890 74864
rect 18930 74824 18972 74864
rect 19012 74824 19054 74864
rect 19094 74824 19136 74864
rect 18808 74815 19176 74824
rect 18988 74696 19028 74705
rect 18892 74444 18932 74453
rect 18892 73856 18932 74404
rect 18892 73807 18932 73816
rect 18988 73520 19028 74656
rect 19084 74612 19124 74621
rect 19084 74276 19124 74572
rect 19276 74276 19316 74992
rect 19372 74696 19412 77428
rect 19372 74647 19412 74656
rect 19468 74528 19508 89608
rect 19564 89564 19604 89573
rect 19564 83852 19604 89524
rect 19564 83803 19604 83812
rect 19564 83684 19604 83693
rect 19564 82424 19604 83644
rect 19564 82375 19604 82384
rect 19660 82172 19700 91120
rect 19756 89648 19796 89657
rect 19756 89513 19796 89608
rect 19756 88808 19796 88817
rect 19756 87968 19796 88768
rect 19852 88052 19892 93724
rect 19948 93680 19988 94900
rect 20236 94184 20276 94193
rect 20236 94049 20276 94144
rect 20048 93764 20416 93773
rect 20088 93724 20130 93764
rect 20170 93724 20212 93764
rect 20252 93724 20294 93764
rect 20334 93724 20376 93764
rect 20048 93715 20416 93724
rect 19948 93631 19988 93640
rect 19948 93344 19988 93353
rect 19948 93209 19988 93304
rect 20140 93344 20180 93353
rect 20140 93209 20180 93304
rect 21004 93176 21044 93185
rect 20524 92672 20564 92681
rect 20048 92252 20416 92261
rect 20088 92212 20130 92252
rect 20170 92212 20212 92252
rect 20252 92212 20294 92252
rect 20334 92212 20376 92252
rect 20048 92203 20416 92212
rect 20140 91160 20180 91169
rect 20140 91025 20180 91120
rect 20048 90740 20416 90749
rect 20088 90700 20130 90740
rect 20170 90700 20212 90740
rect 20252 90700 20294 90740
rect 20334 90700 20376 90740
rect 20048 90691 20416 90700
rect 20140 90320 20180 90329
rect 20140 90185 20180 90280
rect 20140 89648 20180 89657
rect 20140 89513 20180 89608
rect 20048 89228 20416 89237
rect 20088 89188 20130 89228
rect 20170 89188 20212 89228
rect 20252 89188 20294 89228
rect 20334 89188 20376 89228
rect 20048 89179 20416 89188
rect 20524 88892 20564 92632
rect 21004 92672 21044 93136
rect 21004 92623 21044 92632
rect 21004 92420 21044 92429
rect 20908 91832 20948 91841
rect 20812 91664 20852 91673
rect 20716 90992 20756 91001
rect 20716 90152 20756 90952
rect 20812 90656 20852 91624
rect 20812 90607 20852 90616
rect 20716 90103 20756 90112
rect 20812 90068 20852 90077
rect 20428 88852 20564 88892
rect 20620 89480 20660 89489
rect 19852 88003 19892 88012
rect 20140 88808 20180 88817
rect 19756 87919 19796 87928
rect 19852 87884 19892 87893
rect 19756 87296 19796 87305
rect 19756 87161 19796 87256
rect 19564 82132 19700 82172
rect 19756 86624 19796 86633
rect 19564 78980 19604 82132
rect 19660 82004 19700 82013
rect 19660 79148 19700 81964
rect 19660 79099 19700 79108
rect 19564 78940 19700 78980
rect 19564 78812 19604 78821
rect 19564 78224 19604 78772
rect 19564 78175 19604 78184
rect 19084 74227 19124 74236
rect 19180 74236 19316 74276
rect 19372 74488 19508 74528
rect 19564 78056 19604 78065
rect 18988 73471 19028 73480
rect 19180 73520 19220 74236
rect 19180 73471 19220 73480
rect 19276 73940 19316 73949
rect 18808 73352 19176 73361
rect 18848 73312 18890 73352
rect 18930 73312 18972 73352
rect 19012 73312 19054 73352
rect 19094 73312 19136 73352
rect 18808 73303 19176 73312
rect 19276 73184 19316 73900
rect 19276 73135 19316 73144
rect 19084 72932 19124 72941
rect 18892 72892 19084 72932
rect 18796 72260 18836 72269
rect 18796 72092 18836 72220
rect 18796 72043 18836 72052
rect 18892 72092 18932 72892
rect 19084 72883 19124 72892
rect 19180 72848 19220 72857
rect 19084 72764 19124 72773
rect 19084 72629 19124 72724
rect 18892 72043 18932 72052
rect 19084 72260 19124 72269
rect 19084 72008 19124 72220
rect 19180 72008 19220 72808
rect 19180 71968 19316 72008
rect 19084 71959 19124 71968
rect 18808 71840 19176 71849
rect 18848 71800 18890 71840
rect 18930 71800 18972 71840
rect 19012 71800 19054 71840
rect 19094 71800 19136 71840
rect 18808 71791 19176 71800
rect 18892 71672 18932 71681
rect 18892 70496 18932 71632
rect 18988 71252 19028 71261
rect 18988 70832 19028 71212
rect 19276 71000 19316 71968
rect 19276 70951 19316 70960
rect 18988 70783 19028 70792
rect 18892 70447 18932 70456
rect 19276 70748 19316 70757
rect 18808 70328 19176 70337
rect 18848 70288 18890 70328
rect 18930 70288 18972 70328
rect 19012 70288 19054 70328
rect 19094 70288 19136 70328
rect 18808 70279 19176 70288
rect 18796 70160 18836 70169
rect 18796 69908 18836 70120
rect 18796 69320 18836 69868
rect 19084 70160 19124 70169
rect 18796 69271 18836 69280
rect 18892 69740 18932 69749
rect 18892 69152 18932 69700
rect 18892 69103 18932 69112
rect 19084 69656 19124 70120
rect 19276 70076 19316 70708
rect 19276 70027 19316 70036
rect 19084 68984 19124 69616
rect 19084 68935 19124 68944
rect 19276 69908 19316 69917
rect 18808 68816 19176 68825
rect 18848 68776 18890 68816
rect 18930 68776 18972 68816
rect 19012 68776 19054 68816
rect 19094 68776 19136 68816
rect 18808 68767 19176 68776
rect 18796 68648 18836 68657
rect 18796 68396 18836 68608
rect 19276 68648 19316 69868
rect 19276 68599 19316 68608
rect 18796 67556 18836 68356
rect 18796 67507 18836 67516
rect 19276 68480 19316 68489
rect 18808 67304 19176 67313
rect 18848 67264 18890 67304
rect 18930 67264 18972 67304
rect 19012 67264 19054 67304
rect 19094 67264 19136 67304
rect 18808 67255 19176 67264
rect 18796 67136 18836 67145
rect 18796 66884 18836 67096
rect 18796 66835 18836 66844
rect 19276 66380 19316 68440
rect 19180 66340 19316 66380
rect 19180 66128 19220 66340
rect 19180 65993 19220 66088
rect 19276 66212 19316 66221
rect 18808 65792 19176 65801
rect 18848 65752 18890 65792
rect 18930 65752 18972 65792
rect 19012 65752 19054 65792
rect 19094 65752 19136 65792
rect 18808 65743 19176 65752
rect 19084 65372 19124 65381
rect 19084 65036 19124 65332
rect 19084 64987 19124 64996
rect 19180 65288 19220 65297
rect 19180 64868 19220 65248
rect 19180 64819 19220 64828
rect 18808 64280 19176 64289
rect 18848 64240 18890 64280
rect 18930 64240 18972 64280
rect 19012 64240 19054 64280
rect 19094 64240 19136 64280
rect 18808 64231 19176 64240
rect 19276 64028 19316 66172
rect 19276 63979 19316 63988
rect 18796 63860 18836 63869
rect 18796 63104 18836 63820
rect 18988 63860 19028 63869
rect 18988 63725 19028 63820
rect 19180 63860 19220 63869
rect 19180 63188 19220 63820
rect 19372 63440 19412 74488
rect 19564 74444 19604 78016
rect 19372 63391 19412 63400
rect 19468 74404 19604 74444
rect 19468 63272 19508 74404
rect 19660 73940 19700 78940
rect 19660 73891 19700 73900
rect 19756 73772 19796 86584
rect 19852 83600 19892 87844
rect 20140 87884 20180 88768
rect 20236 88724 20276 88733
rect 20236 87968 20276 88684
rect 20332 88640 20372 88649
rect 20332 88505 20372 88600
rect 20428 88136 20468 88852
rect 20620 88640 20660 89440
rect 20620 88591 20660 88600
rect 20716 89312 20756 89321
rect 20428 88096 20660 88136
rect 20236 87919 20276 87928
rect 20140 87835 20180 87844
rect 20048 87716 20416 87725
rect 20088 87676 20130 87716
rect 20170 87676 20212 87716
rect 20252 87676 20294 87716
rect 20334 87676 20376 87716
rect 20048 87667 20416 87676
rect 20236 87548 20276 87557
rect 20140 87296 20180 87305
rect 20140 87161 20180 87256
rect 20140 86624 20180 86633
rect 20140 86489 20180 86584
rect 19852 83551 19892 83560
rect 19948 86372 19988 86381
rect 19948 83516 19988 86332
rect 20236 86372 20276 87508
rect 20236 86323 20276 86332
rect 20524 87464 20564 87473
rect 20048 86204 20416 86213
rect 20088 86164 20130 86204
rect 20170 86164 20212 86204
rect 20252 86164 20294 86204
rect 20334 86164 20376 86204
rect 20048 86155 20416 86164
rect 20044 85868 20084 85877
rect 20044 85028 20084 85828
rect 20044 84979 20084 84988
rect 20048 84692 20416 84701
rect 20088 84652 20130 84692
rect 20170 84652 20212 84692
rect 20252 84652 20294 84692
rect 20334 84652 20376 84692
rect 20048 84643 20416 84652
rect 20140 84272 20180 84281
rect 20140 84137 20180 84232
rect 19948 83467 19988 83476
rect 20044 84104 20084 84113
rect 19852 83432 19892 83441
rect 19852 77720 19892 83392
rect 20044 83348 20084 84064
rect 20140 83600 20180 83695
rect 20140 83551 20180 83560
rect 19948 83308 20084 83348
rect 19948 79988 19988 83308
rect 20048 83180 20416 83189
rect 20088 83140 20130 83180
rect 20170 83140 20212 83180
rect 20252 83140 20294 83180
rect 20334 83140 20376 83180
rect 20048 83131 20416 83140
rect 20044 83012 20084 83021
rect 20044 81836 20084 82972
rect 20044 81787 20084 81796
rect 20048 81668 20416 81677
rect 20088 81628 20130 81668
rect 20170 81628 20212 81668
rect 20252 81628 20294 81668
rect 20334 81628 20376 81668
rect 20048 81619 20416 81628
rect 20044 81416 20084 81425
rect 20044 80408 20084 81376
rect 20044 80359 20084 80368
rect 20048 80156 20416 80165
rect 20088 80116 20130 80156
rect 20170 80116 20212 80156
rect 20252 80116 20294 80156
rect 20334 80116 20376 80156
rect 20048 80107 20416 80116
rect 19948 79948 20084 79988
rect 19948 79820 19988 79829
rect 19948 79232 19988 79780
rect 19948 79183 19988 79192
rect 20044 78896 20084 79948
rect 20140 79736 20180 79745
rect 20140 79316 20180 79696
rect 20140 79267 20180 79276
rect 20428 79568 20468 79577
rect 20044 78847 20084 78856
rect 19852 77671 19892 77680
rect 19948 78812 19988 78821
rect 19948 77468 19988 78772
rect 20428 78812 20468 79528
rect 20428 78763 20468 78772
rect 20048 78644 20416 78653
rect 20088 78604 20130 78644
rect 20170 78604 20212 78644
rect 20252 78604 20294 78644
rect 20334 78604 20376 78644
rect 20048 78595 20416 78604
rect 20044 78392 20084 78401
rect 20044 78257 20084 78352
rect 20140 78308 20180 78317
rect 20044 78140 20084 78149
rect 20044 78005 20084 78100
rect 20140 78056 20180 78268
rect 19948 77419 19988 77428
rect 19852 77384 19892 77393
rect 19852 76628 19892 77344
rect 20140 77300 20180 78016
rect 19948 77260 20180 77300
rect 19948 76796 19988 77260
rect 20048 77132 20416 77141
rect 20088 77092 20130 77132
rect 20170 77092 20212 77132
rect 20252 77092 20294 77132
rect 20334 77092 20376 77132
rect 20048 77083 20416 77092
rect 19948 76747 19988 76756
rect 20140 76796 20180 76891
rect 20140 76747 20180 76756
rect 20140 76628 20180 76637
rect 19852 76588 20140 76628
rect 20140 76579 20180 76588
rect 20428 76628 20468 76637
rect 19564 73732 19796 73772
rect 19852 76460 19892 76469
rect 19564 68396 19604 73732
rect 19660 73604 19700 73613
rect 19660 73016 19700 73564
rect 19660 72967 19700 72976
rect 19756 73520 19796 73529
rect 19660 72848 19700 72857
rect 19660 70328 19700 72808
rect 19756 71420 19796 73480
rect 19852 72932 19892 76420
rect 20140 76040 20180 76049
rect 20140 75905 20180 76000
rect 19948 75788 19988 75797
rect 19948 74444 19988 75748
rect 20428 75788 20468 76588
rect 20428 75739 20468 75748
rect 20048 75620 20416 75629
rect 20088 75580 20130 75620
rect 20170 75580 20212 75620
rect 20252 75580 20294 75620
rect 20334 75580 20376 75620
rect 20048 75571 20416 75580
rect 20428 75452 20468 75461
rect 20332 75116 20372 75125
rect 19948 74395 19988 74404
rect 20044 75032 20084 75041
rect 20044 74276 20084 74992
rect 20332 74528 20372 75076
rect 20332 74479 20372 74488
rect 19852 72883 19892 72892
rect 19948 74236 20084 74276
rect 20428 74276 20468 75412
rect 19756 71371 19796 71380
rect 19852 72764 19892 72773
rect 19660 70279 19700 70288
rect 19756 71168 19796 71177
rect 19756 70160 19796 71128
rect 19852 70748 19892 72724
rect 19948 72260 19988 74236
rect 20428 74227 20468 74236
rect 20048 74108 20416 74117
rect 20088 74068 20130 74108
rect 20170 74068 20212 74108
rect 20252 74068 20294 74108
rect 20334 74068 20376 74108
rect 20048 74059 20416 74068
rect 20044 73940 20084 73949
rect 20044 72764 20084 73900
rect 20428 73940 20468 73949
rect 20428 72848 20468 73900
rect 20428 72799 20468 72808
rect 20044 72715 20084 72724
rect 20048 72596 20416 72605
rect 20088 72556 20130 72596
rect 20170 72556 20212 72596
rect 20252 72556 20294 72596
rect 20334 72556 20376 72596
rect 20048 72547 20416 72556
rect 19948 72211 19988 72220
rect 20044 72428 20084 72437
rect 19948 71588 19988 71597
rect 19948 71504 19988 71548
rect 19948 71453 19988 71464
rect 20044 71252 20084 72388
rect 20332 72344 20372 72353
rect 20332 71504 20372 72304
rect 20332 71455 20372 71464
rect 19948 71212 20044 71252
rect 19948 70832 19988 71212
rect 20044 71203 20084 71212
rect 20048 71084 20416 71093
rect 20088 71044 20130 71084
rect 20170 71044 20212 71084
rect 20252 71044 20294 71084
rect 20334 71044 20376 71084
rect 20048 71035 20416 71044
rect 20332 70916 20372 70925
rect 19948 70792 20084 70832
rect 19852 70708 19988 70748
rect 19756 70111 19796 70120
rect 19852 70580 19892 70589
rect 19660 70076 19700 70085
rect 19660 68480 19700 70036
rect 19756 69992 19796 70001
rect 19756 69857 19796 69952
rect 19756 69740 19796 69749
rect 19756 68648 19796 69700
rect 19852 69236 19892 70540
rect 19852 69187 19892 69196
rect 19756 68599 19796 68608
rect 19852 68480 19892 68489
rect 19660 68440 19796 68480
rect 19564 68356 19700 68396
rect 19180 63139 19220 63148
rect 19372 63232 19508 63272
rect 19564 63944 19604 63953
rect 18796 63055 18836 63064
rect 18988 63020 19028 63115
rect 18988 62971 19028 62980
rect 19276 62852 19316 62861
rect 18808 62768 19176 62777
rect 18848 62728 18890 62768
rect 18930 62728 18972 62768
rect 19012 62728 19054 62768
rect 19094 62728 19136 62768
rect 18808 62719 19176 62728
rect 18796 62600 18836 62609
rect 18796 62012 18836 62560
rect 18796 61963 18836 61972
rect 19180 62600 19220 62609
rect 18988 61592 19028 61601
rect 18988 61457 19028 61552
rect 19180 61508 19220 62560
rect 19180 61459 19220 61468
rect 18808 61256 19176 61265
rect 18848 61216 18890 61256
rect 18930 61216 18972 61256
rect 19012 61216 19054 61256
rect 19094 61216 19136 61256
rect 18808 61207 19176 61216
rect 19180 60920 19220 60929
rect 19180 60080 19220 60880
rect 19180 60031 19220 60040
rect 18808 59744 19176 59753
rect 18848 59704 18890 59744
rect 18930 59704 18972 59744
rect 19012 59704 19054 59744
rect 19094 59704 19136 59744
rect 18808 59695 19176 59704
rect 18796 59492 18836 59501
rect 18796 58736 18836 59452
rect 18796 58484 18836 58696
rect 18796 58435 18836 58444
rect 18808 58232 19176 58241
rect 18848 58192 18890 58232
rect 18930 58192 18972 58232
rect 19012 58192 19054 58232
rect 19094 58192 19136 58232
rect 18808 58183 19176 58192
rect 18796 57896 18836 57905
rect 18796 56888 18836 57856
rect 18892 57812 18932 57821
rect 18892 57677 18932 57772
rect 18796 56839 18836 56848
rect 18808 56720 19176 56729
rect 18848 56680 18890 56720
rect 18930 56680 18972 56720
rect 19012 56680 19054 56720
rect 19094 56680 19136 56720
rect 18808 56671 19176 56680
rect 18796 56384 18836 56393
rect 18796 55376 18836 56344
rect 19180 56384 19220 56393
rect 19180 56300 19220 56344
rect 19180 56249 19220 56260
rect 18796 55327 18836 55336
rect 18808 55208 19176 55217
rect 18848 55168 18890 55208
rect 18930 55168 18972 55208
rect 19012 55168 19054 55208
rect 19094 55168 19136 55208
rect 18808 55159 19176 55168
rect 18796 55040 18836 55049
rect 18796 54116 18836 55000
rect 18892 55040 18932 55049
rect 18892 54368 18932 55000
rect 18892 54319 18932 54328
rect 19084 54536 19124 54545
rect 18796 53864 18836 54076
rect 19084 54116 19124 54496
rect 19084 54067 19124 54076
rect 18892 54032 18932 54041
rect 18892 53897 18932 53992
rect 18796 53815 18836 53824
rect 18808 53696 19176 53705
rect 18848 53656 18890 53696
rect 18930 53656 18972 53696
rect 19012 53656 19054 53696
rect 19094 53656 19136 53696
rect 18808 53647 19176 53656
rect 19084 53276 19124 53285
rect 19084 52772 19124 53236
rect 19084 52723 19124 52732
rect 18808 52184 19176 52193
rect 18848 52144 18890 52184
rect 18930 52144 18972 52184
rect 19012 52144 19054 52184
rect 19094 52144 19136 52184
rect 18808 52135 19176 52144
rect 18808 50672 19176 50681
rect 18848 50632 18890 50672
rect 18930 50632 18972 50672
rect 19012 50632 19054 50672
rect 19094 50632 19136 50672
rect 18808 50623 19176 50632
rect 19180 50252 19220 50261
rect 19180 50117 19220 50212
rect 18808 49160 19176 49169
rect 18848 49120 18890 49160
rect 18930 49120 18972 49160
rect 19012 49120 19054 49160
rect 19094 49120 19136 49160
rect 18808 49111 19176 49120
rect 19276 48236 19316 62812
rect 19372 58484 19412 63232
rect 19468 63104 19508 63113
rect 19468 61676 19508 63064
rect 19564 62348 19604 63904
rect 19660 63380 19700 68356
rect 19756 66716 19796 68440
rect 19756 66667 19796 66676
rect 19756 66128 19796 66137
rect 19756 63524 19796 66088
rect 19852 63692 19892 68440
rect 19852 63643 19892 63652
rect 19756 63475 19796 63484
rect 19852 63440 19892 63449
rect 19660 63340 19796 63380
rect 19564 62299 19604 62308
rect 19468 61627 19508 61636
rect 19564 62180 19604 62189
rect 19468 61508 19508 61517
rect 19468 60248 19508 61468
rect 19468 59492 19508 60208
rect 19468 59443 19508 59452
rect 19468 59324 19508 59333
rect 19468 59189 19508 59284
rect 19564 58652 19604 62140
rect 19660 61928 19700 61937
rect 19660 60164 19700 61888
rect 19660 60115 19700 60124
rect 19564 58603 19604 58612
rect 19660 59912 19700 59921
rect 19372 58435 19412 58444
rect 19564 58484 19604 58493
rect 19372 58316 19412 58325
rect 19372 53612 19412 58276
rect 19468 57728 19508 57737
rect 19468 54788 19508 57688
rect 19468 54284 19508 54748
rect 19468 54235 19508 54244
rect 19372 53563 19412 53572
rect 19468 54116 19508 54125
rect 19468 53444 19508 54076
rect 19372 53404 19508 53444
rect 19372 53276 19412 53404
rect 19372 53227 19412 53236
rect 19468 53276 19508 53285
rect 19372 51008 19412 51017
rect 19372 50873 19412 50968
rect 19468 50504 19508 53236
rect 19372 50464 19508 50504
rect 19372 49664 19412 50464
rect 19372 49615 19412 49624
rect 19468 50336 19508 50345
rect 19372 49496 19412 49505
rect 19372 49361 19412 49456
rect 19468 48992 19508 50296
rect 19468 48943 19508 48952
rect 19372 48824 19412 48833
rect 19372 48689 19412 48784
rect 19468 48740 19508 48749
rect 19276 48196 19412 48236
rect 19276 48068 19316 48077
rect 18808 47648 19176 47657
rect 18848 47608 18890 47648
rect 18930 47608 18972 47648
rect 19012 47608 19054 47648
rect 19094 47608 19136 47648
rect 18808 47599 19176 47608
rect 19276 47228 19316 48028
rect 19276 47179 19316 47188
rect 19276 46304 19316 46313
rect 18808 46136 19176 46145
rect 18848 46096 18890 46136
rect 18930 46096 18972 46136
rect 19012 46096 19054 46136
rect 19094 46096 19136 46136
rect 18808 46087 19176 46096
rect 18892 45716 18932 45725
rect 19276 45716 19316 46264
rect 18932 45676 19028 45716
rect 18892 45667 18932 45676
rect 18892 45212 18932 45221
rect 18892 45077 18932 45172
rect 18988 45044 19028 45676
rect 19276 45667 19316 45676
rect 18988 44995 19028 45004
rect 19276 45044 19316 45053
rect 18808 44624 19176 44633
rect 18848 44584 18890 44624
rect 18930 44584 18972 44624
rect 19012 44584 19054 44624
rect 19094 44584 19136 44624
rect 18808 44575 19176 44584
rect 19276 44540 19316 45004
rect 19276 44491 19316 44500
rect 18700 44416 18836 44456
rect 18508 42776 18548 43492
rect 18508 42727 18548 42736
rect 18604 43448 18644 43457
rect 18604 42692 18644 43408
rect 18604 42104 18644 42652
rect 18604 42055 18644 42064
rect 18700 43364 18740 43373
rect 18412 41971 18452 41980
rect 18700 42020 18740 43324
rect 18796 43280 18836 44416
rect 18796 43231 18836 43240
rect 19276 43532 19316 43541
rect 18808 43112 19176 43121
rect 18848 43072 18890 43112
rect 18930 43072 18972 43112
rect 19012 43072 19054 43112
rect 19094 43072 19136 43112
rect 18808 43063 19176 43072
rect 18700 41971 18740 41980
rect 18796 42944 18836 42953
rect 18412 41768 18452 41777
rect 18796 41768 18836 42904
rect 19276 42692 19316 43492
rect 19276 42643 19316 42652
rect 18412 40676 18452 41728
rect 18700 41728 18836 41768
rect 18412 40627 18452 40636
rect 18508 41684 18548 41693
rect 18508 41180 18548 41644
rect 18700 41348 18740 41728
rect 18808 41600 19176 41609
rect 18848 41560 18890 41600
rect 18930 41560 18972 41600
rect 19012 41560 19054 41600
rect 19094 41560 19136 41600
rect 18808 41551 19176 41560
rect 18700 41299 18740 41308
rect 18988 41264 19028 41273
rect 18508 40508 18548 41140
rect 18892 41180 18932 41189
rect 18892 41096 18932 41140
rect 18412 40468 18548 40508
rect 18700 41056 18932 41096
rect 18412 38912 18452 40468
rect 18604 40424 18644 40433
rect 18508 39920 18548 39929
rect 18508 39752 18548 39880
rect 18508 39703 18548 39712
rect 18412 38863 18452 38872
rect 18508 39164 18548 39173
rect 18508 38912 18548 39124
rect 18412 38744 18452 38753
rect 18412 38324 18452 38704
rect 18412 38275 18452 38284
rect 18508 38408 18548 38872
rect 18316 35755 18356 35764
rect 18412 38072 18452 38081
rect 18412 37568 18452 38032
rect 18412 36056 18452 37528
rect 18412 35636 18452 36016
rect 18220 35335 18260 35344
rect 18316 35596 18452 35636
rect 18124 34915 18164 34924
rect 18220 35048 18260 35057
rect 17932 34663 17972 34672
rect 18124 34712 18164 34721
rect 17452 33487 17492 33496
rect 17548 33916 17876 33956
rect 17932 34460 17972 34469
rect 17164 32563 17204 32572
rect 17356 32696 17396 32705
rect 16972 30428 17012 31312
rect 17260 32192 17300 32201
rect 17260 30932 17300 32152
rect 17260 30883 17300 30892
rect 17164 30680 17204 30689
rect 16972 30379 17012 30388
rect 17068 30596 17108 30605
rect 17068 30344 17108 30556
rect 17068 29672 17108 30304
rect 17068 29623 17108 29632
rect 17164 29084 17204 30640
rect 17260 29924 17300 29933
rect 17260 29789 17300 29884
rect 16876 28027 16916 28036
rect 16972 29044 17204 29084
rect 17260 29084 17300 29179
rect 16780 27859 16820 27868
rect 16780 27404 16820 27413
rect 16780 26900 16820 27364
rect 16780 26851 16820 26860
rect 16780 26648 16820 26657
rect 16780 26060 16820 26608
rect 16780 26011 16820 26020
rect 16876 26060 16916 26069
rect 16684 25516 16820 25556
rect 16684 25388 16724 25397
rect 16588 24884 16628 24893
rect 16588 24044 16628 24844
rect 16588 23995 16628 24004
rect 16684 24632 16724 25348
rect 16396 23792 16436 23801
rect 16396 23657 16436 23752
rect 16300 21643 16340 21652
rect 16396 23456 16436 23465
rect 16300 21524 16340 21533
rect 16108 20719 16148 20728
rect 16204 20852 16244 20861
rect 16012 19963 16052 19972
rect 16108 20516 16148 20525
rect 16012 19844 16052 19853
rect 16012 19592 16052 19804
rect 16012 19172 16052 19552
rect 16012 19123 16052 19132
rect 16108 19340 16148 20476
rect 15820 17576 15860 17585
rect 15820 12788 15860 17536
rect 15820 12739 15860 12748
rect 15820 11444 15860 11453
rect 15820 11360 15860 11404
rect 15820 11309 15860 11320
rect 15916 10016 15956 17620
rect 16012 19004 16052 19013
rect 16012 14384 16052 18964
rect 16108 18500 16148 19300
rect 16108 18451 16148 18460
rect 16012 14335 16052 14344
rect 16108 18164 16148 18173
rect 16012 14216 16052 14225
rect 16012 13124 16052 14176
rect 16108 13292 16148 18124
rect 16204 16148 16244 20812
rect 16300 20180 16340 21484
rect 16300 20131 16340 20140
rect 16204 14216 16244 16108
rect 16300 18500 16340 18509
rect 16300 15644 16340 18460
rect 16300 15595 16340 15604
rect 16204 14167 16244 14176
rect 16300 15476 16340 15485
rect 16108 13243 16148 13252
rect 16204 13964 16244 13973
rect 16012 13084 16148 13124
rect 16108 12980 16148 13084
rect 15820 9764 15860 9773
rect 15820 8588 15860 9724
rect 15916 8924 15956 9976
rect 15916 8875 15956 8884
rect 16012 12940 16148 12980
rect 15820 8539 15860 8548
rect 15916 8756 15956 8765
rect 15916 7832 15956 8716
rect 16012 8000 16052 12940
rect 16204 12284 16244 13924
rect 16300 13292 16340 15436
rect 16396 13964 16436 23416
rect 16588 23288 16628 23297
rect 16492 22952 16532 22961
rect 16492 21272 16532 22912
rect 16588 21524 16628 23248
rect 16684 23120 16724 24592
rect 16780 23288 16820 25516
rect 16780 23239 16820 23248
rect 16684 23071 16724 23080
rect 16876 23036 16916 26020
rect 16972 25304 17012 29044
rect 17260 29035 17300 29044
rect 17068 28916 17108 28925
rect 17068 26900 17108 28876
rect 17260 28916 17300 28925
rect 17068 26851 17108 26860
rect 17164 28412 17204 28421
rect 17164 27572 17204 28372
rect 16972 24884 17012 25264
rect 16972 24835 17012 24844
rect 17068 26732 17108 26741
rect 16876 22987 16916 22996
rect 16972 24716 17012 24725
rect 16684 22952 16724 22961
rect 16684 22364 16724 22912
rect 16684 22315 16724 22324
rect 16876 22364 16916 22373
rect 16588 21484 16724 21524
rect 16492 21223 16532 21232
rect 16588 21356 16628 21365
rect 16492 20936 16532 21031
rect 16492 20887 16532 20896
rect 16492 20768 16532 20777
rect 16492 20264 16532 20728
rect 16492 20215 16532 20224
rect 16588 19424 16628 21316
rect 16684 20012 16724 21484
rect 16724 19972 16820 20012
rect 16684 19963 16724 19972
rect 16588 19375 16628 19384
rect 16492 19088 16532 19097
rect 16492 17912 16532 19048
rect 16492 17863 16532 17872
rect 16588 18668 16628 18677
rect 16492 17744 16532 17755
rect 16492 17660 16532 17704
rect 16492 17611 16532 17620
rect 16588 17072 16628 18628
rect 16684 17828 16724 17837
rect 16684 17240 16724 17788
rect 16684 17191 16724 17200
rect 16588 17032 16724 17072
rect 16492 16820 16532 16829
rect 16492 15476 16532 16780
rect 16492 15427 16532 15436
rect 16588 14468 16628 14477
rect 16396 13915 16436 13924
rect 16492 14048 16532 14057
rect 16300 13243 16340 13252
rect 16396 13796 16436 13805
rect 16396 13124 16436 13756
rect 16108 12200 16148 12209
rect 16108 11696 16148 12160
rect 16108 11647 16148 11656
rect 16204 11276 16244 12244
rect 16108 11236 16244 11276
rect 16300 13084 16436 13124
rect 16108 8840 16148 11236
rect 16300 10352 16340 13084
rect 16492 12200 16532 14008
rect 16588 13208 16628 14428
rect 16684 13880 16724 17032
rect 16780 14048 16820 19972
rect 16876 18164 16916 22324
rect 16876 18115 16916 18124
rect 16876 16568 16916 16577
rect 16876 16484 16916 16528
rect 16876 16433 16916 16444
rect 16972 16316 17012 24676
rect 17068 18668 17108 26692
rect 17164 21188 17204 27532
rect 17260 26648 17300 28876
rect 17260 26599 17300 26608
rect 17260 26144 17300 26153
rect 17260 26060 17300 26104
rect 17260 26009 17300 26020
rect 17260 24632 17300 24641
rect 17260 24497 17300 24592
rect 17260 23624 17300 23633
rect 17260 23489 17300 23584
rect 17260 23036 17300 23045
rect 17260 22196 17300 22996
rect 17260 22147 17300 22156
rect 17164 19676 17204 21148
rect 17260 21524 17300 21533
rect 17260 20432 17300 21484
rect 17260 20383 17300 20392
rect 17164 19627 17204 19636
rect 17068 18619 17108 18628
rect 17164 18584 17204 18593
rect 17204 18544 17300 18584
rect 17164 18535 17204 18544
rect 17260 17828 17300 18544
rect 17260 17779 17300 17788
rect 17260 17240 17300 17249
rect 17260 17105 17300 17200
rect 17356 16988 17396 32656
rect 17452 32444 17492 32453
rect 17452 32108 17492 32404
rect 17452 32059 17492 32068
rect 17452 31436 17492 31445
rect 17452 30008 17492 31396
rect 17452 29959 17492 29968
rect 17452 29840 17492 29849
rect 17452 28580 17492 29800
rect 17452 28531 17492 28540
rect 17452 27740 17492 27749
rect 17452 23204 17492 27700
rect 17452 23155 17492 23164
rect 16972 16267 17012 16276
rect 17068 16948 17396 16988
rect 17452 22532 17492 22541
rect 16972 15476 17012 15485
rect 16876 15140 16916 15149
rect 16876 14804 16916 15100
rect 16876 14755 16916 14764
rect 16780 13999 16820 14008
rect 16876 13964 16916 13973
rect 16684 13840 16820 13880
rect 16588 13159 16628 13168
rect 16684 13292 16724 13301
rect 16492 12151 16532 12160
rect 16588 13040 16628 13049
rect 16492 10940 16532 10949
rect 16588 10940 16628 13000
rect 16684 12452 16724 13252
rect 16684 12403 16724 12412
rect 16532 10900 16628 10940
rect 16108 8791 16148 8800
rect 16204 10312 16300 10352
rect 16012 7951 16052 7960
rect 16108 8672 16148 8681
rect 15916 7792 16052 7832
rect 15820 7748 15860 7757
rect 15820 6656 15860 7708
rect 15820 6607 15860 6616
rect 15916 6488 15956 6497
rect 15820 5816 15860 5825
rect 15820 5144 15860 5776
rect 15820 5095 15860 5104
rect 15916 4724 15956 6448
rect 15916 4675 15956 4684
rect 16012 6404 16052 7792
rect 16108 7160 16148 8632
rect 16204 7916 16244 10312
rect 16300 10303 16340 10312
rect 16396 10772 16436 10781
rect 16300 9596 16340 9605
rect 16300 9092 16340 9556
rect 16300 8756 16340 9052
rect 16300 8707 16340 8716
rect 16300 8168 16340 8177
rect 16300 8033 16340 8128
rect 16204 7867 16244 7876
rect 16108 7111 16148 7120
rect 16300 7244 16340 7253
rect 16012 4556 16052 6364
rect 16300 5732 16340 7204
rect 16396 6824 16436 10732
rect 16492 9764 16532 10900
rect 16492 8756 16532 9724
rect 16492 8707 16532 8716
rect 16588 9260 16628 9269
rect 16396 6775 16436 6784
rect 16492 8588 16532 8597
rect 16300 5683 16340 5692
rect 16396 6320 16436 6329
rect 16396 5144 16436 6280
rect 16492 5732 16532 8548
rect 16588 6572 16628 9220
rect 16588 6523 16628 6532
rect 16684 8924 16724 8933
rect 16492 5683 16532 5692
rect 16684 6404 16724 8884
rect 16396 4892 16436 5104
rect 16396 4843 16436 4852
rect 16684 4808 16724 6364
rect 16684 4759 16724 4768
rect 16012 4507 16052 4516
rect 16780 2900 16820 13840
rect 16876 12704 16916 13924
rect 16972 13796 17012 15436
rect 16972 13747 17012 13756
rect 16972 13544 17012 13553
rect 16972 13208 17012 13504
rect 16972 13159 17012 13168
rect 16876 12655 16916 12664
rect 16972 13040 17012 13049
rect 16972 12620 17012 13000
rect 16972 12571 17012 12580
rect 16972 12200 17012 12209
rect 16972 11780 17012 12160
rect 16972 11528 17012 11740
rect 16876 10940 16916 10949
rect 16876 9680 16916 10900
rect 16876 9631 16916 9640
rect 16972 8924 17012 11488
rect 16972 8875 17012 8884
rect 16972 6404 17012 6413
rect 16972 5900 17012 6364
rect 16972 5851 17012 5860
rect 15724 1903 15764 1912
rect 16492 2860 16820 2900
rect 17068 2900 17108 16948
rect 17260 16148 17300 16157
rect 17260 16013 17300 16108
rect 17452 15476 17492 22492
rect 17452 15427 17492 15436
rect 17164 15392 17204 15401
rect 17164 14720 17204 15352
rect 17452 15308 17492 15317
rect 17164 12452 17204 14680
rect 17260 14804 17300 14813
rect 17260 14669 17300 14764
rect 17356 14636 17396 14645
rect 17260 14384 17300 14393
rect 17260 13124 17300 14344
rect 17356 13460 17396 14596
rect 17356 13411 17396 13420
rect 17260 13084 17396 13124
rect 17260 12956 17300 13084
rect 17356 13040 17396 13084
rect 17356 12991 17396 13000
rect 17260 12907 17300 12916
rect 17452 12872 17492 15268
rect 17452 12823 17492 12832
rect 17356 12704 17396 12713
rect 17356 12569 17396 12664
rect 17164 12412 17300 12452
rect 17164 12284 17204 12293
rect 17164 11780 17204 12244
rect 17164 11731 17204 11740
rect 17260 10688 17300 12412
rect 17452 12368 17492 12377
rect 17260 6572 17300 10648
rect 17356 12328 17452 12368
rect 17356 10268 17396 12328
rect 17452 12233 17492 12328
rect 17356 10219 17396 10228
rect 17452 11948 17492 11957
rect 17452 10268 17492 11908
rect 17356 8756 17396 8765
rect 17356 7160 17396 8716
rect 17452 8672 17492 10228
rect 17548 9428 17588 33916
rect 17740 33788 17780 33797
rect 17644 31940 17684 31949
rect 17644 25220 17684 31900
rect 17740 31856 17780 33748
rect 17836 33536 17876 33545
rect 17836 32024 17876 33496
rect 17932 32864 17972 34420
rect 18124 33116 18164 34672
rect 18220 33200 18260 35008
rect 18316 34880 18356 35596
rect 18316 34831 18356 34840
rect 18412 35132 18452 35141
rect 18220 33151 18260 33160
rect 18316 34208 18356 34217
rect 18124 33067 18164 33076
rect 18220 32948 18260 32957
rect 17932 32780 17972 32824
rect 17932 32731 17972 32740
rect 18028 32864 18068 32873
rect 17932 32192 17972 32201
rect 17932 32057 17972 32152
rect 17836 31975 17876 31984
rect 17740 31816 17876 31856
rect 17740 30596 17780 30605
rect 17740 29336 17780 30556
rect 17740 29287 17780 29296
rect 17836 30092 17876 31816
rect 17740 27152 17780 27161
rect 17740 26816 17780 27112
rect 17740 26767 17780 26776
rect 17740 26648 17780 26657
rect 17740 26513 17780 26608
rect 17740 25892 17780 25901
rect 17740 25388 17780 25852
rect 17740 25339 17780 25348
rect 17644 25180 17780 25220
rect 17644 25052 17684 25061
rect 17644 22364 17684 25012
rect 17740 22532 17780 25180
rect 17836 25052 17876 30052
rect 17932 29672 17972 29681
rect 17932 29168 17972 29632
rect 17932 29119 17972 29128
rect 17836 25003 17876 25012
rect 17932 29000 17972 29009
rect 17932 28244 17972 28960
rect 18028 28748 18068 32824
rect 18124 32528 18164 32537
rect 18124 30764 18164 32488
rect 18220 31436 18260 32908
rect 18220 31387 18260 31396
rect 18124 29000 18164 30724
rect 18124 28951 18164 28960
rect 18220 30764 18260 30773
rect 18028 28699 18068 28708
rect 17836 24884 17876 24893
rect 17836 24128 17876 24844
rect 17836 24079 17876 24088
rect 17836 23960 17876 23969
rect 17836 23792 17876 23920
rect 17836 23743 17876 23752
rect 17836 23624 17876 23633
rect 17836 23456 17876 23584
rect 17836 23407 17876 23416
rect 17836 23120 17876 23129
rect 17836 22616 17876 23080
rect 17836 22567 17876 22576
rect 17740 22483 17780 22492
rect 17836 22364 17876 22373
rect 17644 22324 17836 22364
rect 17740 21524 17780 21533
rect 17644 20936 17684 20945
rect 17644 13796 17684 20896
rect 17740 20852 17780 21484
rect 17740 20096 17780 20812
rect 17740 20047 17780 20056
rect 17836 20012 17876 22324
rect 17740 19928 17780 19937
rect 17740 19088 17780 19888
rect 17836 19340 17876 19972
rect 17836 19291 17876 19300
rect 17740 19048 17876 19088
rect 17836 18500 17876 19048
rect 17932 18584 17972 28204
rect 18028 28412 18068 28421
rect 18028 24464 18068 28372
rect 18220 27572 18260 30724
rect 18220 27523 18260 27532
rect 18220 27404 18260 27413
rect 18220 26900 18260 27364
rect 18220 26851 18260 26860
rect 18220 26732 18260 26741
rect 18220 25892 18260 26692
rect 18028 23792 18068 24424
rect 18028 23743 18068 23752
rect 18124 25852 18260 25892
rect 18124 25304 18164 25852
rect 18316 25640 18356 34168
rect 18412 30680 18452 35092
rect 18508 33620 18548 38368
rect 18604 38072 18644 40384
rect 18604 38023 18644 38032
rect 18604 37400 18644 37409
rect 18604 36728 18644 37360
rect 18604 36679 18644 36688
rect 18700 36056 18740 41056
rect 18988 40424 19028 41224
rect 18988 40375 19028 40384
rect 19276 40508 19316 40517
rect 18808 40088 19176 40097
rect 18848 40048 18890 40088
rect 18930 40048 18972 40088
rect 19012 40048 19054 40088
rect 19094 40048 19136 40088
rect 18808 40039 19176 40048
rect 18892 39836 18932 39845
rect 18892 39668 18932 39796
rect 18892 39619 18932 39628
rect 18808 38576 19176 38585
rect 18848 38536 18890 38576
rect 18930 38536 18972 38576
rect 19012 38536 19054 38576
rect 19094 38536 19136 38576
rect 18808 38527 19176 38536
rect 19180 38408 19220 38417
rect 19084 38156 19124 38165
rect 18892 37568 18932 37577
rect 18892 37433 18932 37528
rect 19084 37400 19124 38116
rect 19084 37351 19124 37360
rect 19180 37232 19220 38368
rect 19180 37183 19220 37192
rect 19276 38240 19316 40468
rect 19276 37484 19316 38200
rect 18808 37064 19176 37073
rect 18848 37024 18890 37064
rect 18930 37024 18972 37064
rect 19012 37024 19054 37064
rect 19094 37024 19136 37064
rect 18808 37015 19176 37024
rect 18892 36896 18932 36905
rect 18892 36644 18932 36856
rect 18892 36595 18932 36604
rect 19180 36896 19220 36905
rect 19084 36476 19124 36485
rect 18700 36016 18836 36056
rect 18508 33571 18548 33580
rect 18604 35972 18644 35981
rect 18508 33452 18548 33461
rect 18508 33032 18548 33412
rect 18508 32983 18548 32992
rect 18508 32864 18548 32873
rect 18508 32192 18548 32824
rect 18508 32143 18548 32152
rect 18508 32024 18548 32033
rect 18508 31604 18548 31984
rect 18508 31555 18548 31564
rect 18412 29924 18452 30640
rect 18412 29875 18452 29884
rect 18508 31436 18548 31445
rect 18412 29084 18452 29093
rect 18412 28949 18452 29044
rect 18124 23708 18164 25264
rect 18124 23540 18164 23668
rect 18220 25600 18356 25640
rect 18412 28244 18452 28253
rect 18220 23624 18260 25600
rect 18220 23575 18260 23584
rect 18316 25472 18356 25481
rect 18316 24548 18356 25432
rect 18124 23491 18164 23500
rect 18220 23372 18260 23381
rect 18028 23036 18068 23045
rect 18028 22532 18068 22996
rect 18028 22483 18068 22492
rect 18028 22196 18068 22205
rect 18028 21272 18068 22156
rect 18124 21524 18164 21619
rect 18124 21475 18164 21484
rect 18124 21272 18164 21281
rect 18028 21232 18124 21272
rect 17932 18535 17972 18544
rect 18028 21104 18068 21113
rect 18028 20096 18068 21064
rect 17836 18332 17876 18460
rect 17836 18292 17972 18332
rect 17836 18164 17876 18173
rect 17836 17996 17876 18124
rect 17932 18164 17972 18292
rect 17932 18115 17972 18124
rect 17644 11528 17684 13756
rect 17644 11479 17684 11488
rect 17740 17956 17876 17996
rect 18028 17996 18068 20056
rect 18124 19592 18164 21232
rect 18124 19543 18164 19552
rect 17740 11276 17780 17956
rect 18028 17947 18068 17956
rect 18124 18584 18164 18593
rect 17932 17912 17972 17921
rect 17836 17744 17876 17753
rect 17836 17324 17876 17704
rect 17836 17275 17876 17284
rect 17836 16484 17876 16493
rect 17836 16349 17876 16444
rect 17836 16064 17876 16073
rect 17836 13460 17876 16024
rect 17836 13411 17876 13420
rect 17740 10940 17780 11236
rect 17740 10891 17780 10900
rect 17836 12452 17876 12461
rect 17836 10436 17876 12412
rect 17836 10387 17876 10396
rect 17644 10352 17684 10361
rect 17644 9596 17684 10312
rect 17644 9547 17684 9556
rect 17836 10268 17876 10277
rect 17740 9428 17780 9437
rect 17548 9388 17684 9428
rect 17452 7916 17492 8632
rect 17452 7496 17492 7876
rect 17452 7328 17492 7456
rect 17452 7279 17492 7288
rect 17548 9260 17588 9269
rect 17356 7111 17396 7120
rect 17260 6523 17300 6532
rect 17356 6992 17396 7001
rect 17260 6236 17300 6245
rect 17260 3716 17300 6196
rect 17356 4304 17396 6952
rect 17548 4640 17588 9220
rect 17548 4591 17588 4600
rect 17356 4255 17396 4264
rect 17260 3667 17300 3676
rect 17356 4136 17396 4145
rect 17068 2860 17204 2900
rect 16492 1952 16532 2860
rect 17164 2792 17204 2860
rect 17164 2743 17204 2752
rect 17356 2120 17396 4096
rect 17644 3632 17684 9388
rect 17740 8168 17780 9388
rect 17740 8119 17780 8128
rect 17836 4052 17876 10228
rect 17836 4003 17876 4012
rect 17644 3583 17684 3592
rect 17932 2900 17972 17872
rect 18028 17828 18068 17837
rect 18028 17744 18068 17788
rect 18028 17693 18068 17704
rect 18124 17408 18164 18544
rect 18220 18164 18260 23332
rect 18316 22112 18356 24508
rect 18412 23372 18452 28204
rect 18508 27740 18548 31396
rect 18604 28244 18644 35932
rect 18700 35888 18740 35897
rect 18700 34544 18740 35848
rect 18796 35720 18836 36016
rect 19084 35888 19124 36436
rect 19180 36056 19220 36856
rect 19180 35921 19220 36016
rect 19276 35972 19316 37444
rect 19084 35839 19124 35848
rect 18796 35671 18836 35680
rect 18808 35552 19176 35561
rect 18848 35512 18890 35552
rect 18930 35512 18972 35552
rect 19012 35512 19054 35552
rect 19094 35512 19136 35552
rect 18808 35503 19176 35512
rect 18700 34495 18740 34504
rect 18796 35384 18836 35393
rect 18700 34292 18740 34301
rect 18700 33032 18740 34252
rect 18796 34208 18836 35344
rect 19180 35384 19220 35393
rect 18892 35216 18932 35225
rect 18892 35132 18932 35176
rect 18892 34628 18932 35092
rect 18892 34579 18932 34588
rect 18988 34544 19028 34553
rect 18988 34376 19028 34504
rect 18988 34327 19028 34336
rect 18796 34159 18836 34168
rect 19180 34208 19220 35344
rect 19180 34159 19220 34168
rect 18808 34040 19176 34049
rect 18848 34000 18890 34040
rect 18930 34000 18972 34040
rect 19012 34000 19054 34040
rect 19094 34000 19136 34040
rect 18808 33991 19176 34000
rect 19276 33872 19316 35932
rect 18892 33832 19316 33872
rect 18700 32983 18740 32992
rect 18796 33620 18836 33629
rect 18700 32864 18740 32873
rect 18700 32108 18740 32824
rect 18796 32696 18836 33580
rect 18796 32647 18836 32656
rect 18892 32696 18932 33832
rect 19276 33704 19316 33713
rect 18988 33536 19028 33545
rect 18988 33116 19028 33496
rect 18988 33067 19028 33076
rect 18892 32647 18932 32656
rect 18808 32528 19176 32537
rect 18848 32488 18890 32528
rect 18930 32488 18972 32528
rect 19012 32488 19054 32528
rect 19094 32488 19136 32528
rect 18808 32479 19176 32488
rect 18700 32059 18740 32068
rect 18796 32360 18836 32369
rect 18796 31184 18836 32320
rect 19180 32360 19220 32369
rect 19084 32024 19124 32033
rect 19084 31889 19124 31984
rect 18700 31144 18836 31184
rect 19180 31184 19220 32320
rect 18700 30260 18740 31144
rect 19180 31135 19220 31144
rect 18808 31016 19176 31025
rect 18848 30976 18890 31016
rect 18930 30976 18972 31016
rect 19012 30976 19054 31016
rect 19094 30976 19136 31016
rect 18808 30967 19176 30976
rect 18796 30848 18836 30857
rect 18796 30680 18836 30808
rect 18796 30631 18836 30640
rect 19180 30848 19220 30857
rect 19084 30512 19124 30521
rect 18700 30211 18740 30220
rect 18988 30428 19028 30437
rect 18604 28195 18644 28204
rect 18700 30092 18740 30101
rect 18508 27572 18548 27700
rect 18508 27523 18548 27532
rect 18604 27572 18644 27581
rect 18412 23323 18452 23332
rect 18508 26900 18548 26909
rect 18508 23708 18548 26860
rect 18604 26060 18644 27532
rect 18700 26816 18740 30052
rect 18988 30008 19028 30388
rect 18988 29873 19028 29968
rect 19084 29756 19124 30472
rect 19084 29707 19124 29716
rect 19180 29672 19220 30808
rect 19276 30008 19316 33664
rect 19372 30848 19412 48196
rect 19468 47480 19508 48700
rect 19468 47431 19508 47440
rect 19564 47312 19604 58444
rect 19660 55880 19700 59872
rect 19660 55831 19700 55840
rect 19660 55544 19700 55639
rect 19660 55495 19700 55504
rect 19660 55376 19700 55385
rect 19660 53276 19700 55336
rect 19756 53300 19796 63340
rect 19852 57728 19892 63400
rect 19852 57679 19892 57688
rect 19852 57560 19892 57569
rect 19852 56384 19892 57520
rect 19852 56335 19892 56344
rect 19852 55376 19892 55385
rect 19852 54116 19892 55336
rect 19948 55376 19988 70708
rect 20044 69740 20084 70792
rect 20044 69691 20084 69700
rect 20140 69992 20180 70001
rect 20140 69740 20180 69952
rect 20332 69824 20372 70876
rect 20332 69775 20372 69784
rect 20428 70832 20468 70841
rect 20140 69691 20180 69700
rect 20428 69740 20468 70792
rect 20428 69691 20468 69700
rect 20048 69572 20416 69581
rect 20088 69532 20130 69572
rect 20170 69532 20212 69572
rect 20252 69532 20294 69572
rect 20334 69532 20376 69572
rect 20048 69523 20416 69532
rect 20236 69320 20276 69329
rect 20236 68228 20276 69280
rect 20236 68179 20276 68188
rect 20048 68060 20416 68069
rect 20088 68020 20130 68060
rect 20170 68020 20212 68060
rect 20252 68020 20294 68060
rect 20334 68020 20376 68060
rect 20048 68011 20416 68020
rect 20428 67892 20468 67901
rect 20140 67724 20180 67733
rect 20140 66716 20180 67684
rect 20140 66667 20180 66676
rect 20428 66716 20468 67852
rect 20428 66667 20468 66676
rect 20048 66548 20416 66557
rect 20088 66508 20130 66548
rect 20170 66508 20212 66548
rect 20252 66508 20294 66548
rect 20334 66508 20376 66548
rect 20048 66499 20416 66508
rect 20044 65960 20084 65969
rect 20084 65920 20180 65960
rect 20044 65911 20084 65920
rect 20140 65204 20180 65920
rect 20140 65155 20180 65164
rect 20048 65036 20416 65045
rect 20088 64996 20130 65036
rect 20170 64996 20212 65036
rect 20252 64996 20294 65036
rect 20334 64996 20376 65036
rect 20048 64987 20416 64996
rect 20428 64868 20468 64877
rect 20140 64616 20180 64625
rect 20140 64481 20180 64576
rect 20044 64196 20084 64205
rect 20044 64112 20084 64156
rect 20044 64061 20084 64072
rect 20428 63692 20468 64828
rect 20428 63643 20468 63652
rect 20048 63524 20416 63533
rect 20088 63484 20130 63524
rect 20170 63484 20212 63524
rect 20252 63484 20294 63524
rect 20334 63484 20376 63524
rect 20048 63475 20416 63484
rect 20236 63356 20276 63365
rect 20044 62432 20084 62441
rect 20044 62264 20084 62392
rect 20044 62215 20084 62224
rect 20236 62180 20276 63316
rect 20236 62131 20276 62140
rect 20048 62012 20416 62021
rect 20088 61972 20130 62012
rect 20170 61972 20212 62012
rect 20252 61972 20294 62012
rect 20334 61972 20376 62012
rect 20048 61963 20416 61972
rect 20428 61760 20468 61769
rect 20428 61088 20468 61720
rect 20428 61039 20468 61048
rect 20048 60500 20416 60509
rect 20088 60460 20130 60500
rect 20170 60460 20212 60500
rect 20252 60460 20294 60500
rect 20334 60460 20376 60500
rect 20048 60451 20416 60460
rect 20044 60164 20084 60173
rect 20044 59576 20084 60124
rect 20044 59527 20084 59536
rect 20428 59996 20468 60005
rect 20428 59408 20468 59956
rect 20428 59359 20468 59368
rect 20048 58988 20416 58997
rect 20088 58948 20130 58988
rect 20170 58948 20212 58988
rect 20252 58948 20294 58988
rect 20334 58948 20376 58988
rect 20048 58939 20416 58948
rect 20044 58820 20084 58829
rect 20044 57812 20084 58780
rect 20044 57763 20084 57772
rect 20048 57476 20416 57485
rect 20088 57436 20130 57476
rect 20170 57436 20212 57476
rect 20252 57436 20294 57476
rect 20334 57436 20376 57476
rect 20048 57427 20416 57436
rect 20048 55964 20416 55973
rect 20088 55924 20130 55964
rect 20170 55924 20212 55964
rect 20252 55924 20294 55964
rect 20334 55924 20376 55964
rect 20048 55915 20416 55924
rect 19948 55327 19988 55336
rect 19852 54067 19892 54076
rect 19948 54956 19988 54965
rect 19756 53260 19892 53300
rect 19660 53227 19700 53236
rect 19660 53108 19700 53117
rect 19660 52520 19700 53068
rect 19660 52471 19700 52480
rect 19756 52436 19796 52445
rect 19660 51596 19700 51605
rect 19660 50420 19700 51556
rect 19756 51260 19796 52396
rect 19756 51211 19796 51220
rect 19660 50371 19700 50380
rect 19756 50252 19796 50263
rect 19756 50168 19796 50212
rect 19660 49664 19700 49673
rect 19660 47480 19700 49624
rect 19756 48908 19796 50128
rect 19756 48859 19796 48868
rect 19660 47431 19700 47440
rect 19756 47984 19796 47993
rect 19468 47272 19604 47312
rect 19660 47312 19700 47321
rect 19468 34292 19508 47272
rect 19564 47144 19604 47153
rect 19564 45968 19604 47104
rect 19564 45919 19604 45928
rect 19564 45800 19604 45809
rect 19564 44708 19604 45760
rect 19564 44659 19604 44668
rect 19564 43532 19604 43541
rect 19564 42188 19604 43492
rect 19564 42139 19604 42148
rect 19564 40508 19604 40517
rect 19564 38576 19604 40468
rect 19564 38527 19604 38536
rect 19660 38408 19700 47272
rect 19756 43700 19796 47944
rect 19756 43651 19796 43660
rect 19852 43220 19892 53260
rect 19948 53276 19988 54916
rect 20048 54452 20416 54461
rect 20088 54412 20130 54452
rect 20170 54412 20212 54452
rect 20252 54412 20294 54452
rect 20334 54412 20376 54452
rect 20048 54403 20416 54412
rect 19948 53227 19988 53236
rect 20044 54284 20084 54293
rect 20044 53108 20084 54244
rect 20524 53300 20564 87424
rect 20620 62516 20660 88096
rect 20716 87128 20756 89272
rect 20812 88136 20852 90028
rect 20812 88087 20852 88096
rect 20908 87464 20948 91792
rect 21004 91664 21044 92380
rect 21004 91615 21044 91624
rect 21004 90908 21044 90917
rect 21004 89144 21044 90868
rect 21292 90236 21332 90245
rect 21196 89732 21236 89741
rect 21004 89095 21044 89104
rect 21100 89396 21140 89405
rect 20908 87415 20948 87424
rect 21004 88556 21044 88565
rect 20716 87079 20756 87088
rect 20908 86792 20948 86801
rect 20716 86456 20756 86465
rect 20716 85112 20756 86416
rect 20908 85364 20948 86752
rect 21004 86120 21044 88516
rect 21004 86071 21044 86080
rect 20908 85324 21044 85364
rect 20716 85063 20756 85072
rect 20812 84944 20852 84953
rect 20716 84860 20756 84869
rect 20716 81332 20756 84820
rect 20716 81283 20756 81292
rect 20716 80660 20756 80669
rect 20716 68144 20756 80620
rect 20812 79064 20852 84904
rect 20908 84608 20948 84617
rect 20908 84473 20948 84568
rect 20812 79015 20852 79024
rect 20908 84104 20948 84113
rect 20812 78812 20852 78821
rect 20812 73604 20852 78772
rect 20908 78056 20948 84064
rect 21004 81080 21044 85324
rect 21100 84104 21140 89356
rect 21196 85616 21236 89692
rect 21292 86624 21332 90196
rect 21484 88976 21524 88985
rect 21292 86575 21332 86584
rect 21388 88808 21428 88817
rect 21196 85567 21236 85576
rect 21292 86372 21332 86381
rect 21100 84055 21140 84064
rect 21196 85448 21236 85457
rect 21196 83768 21236 85408
rect 21292 85112 21332 86332
rect 21292 85063 21332 85072
rect 21196 83719 21236 83728
rect 21292 84020 21332 84029
rect 21196 83600 21236 83609
rect 21004 81031 21044 81040
rect 21100 82676 21140 82685
rect 20908 78007 20948 78016
rect 21004 79652 21044 79661
rect 20908 77888 20948 77897
rect 20908 75956 20948 77848
rect 20908 75907 20948 75916
rect 20812 73555 20852 73564
rect 20908 75788 20948 75797
rect 20908 73460 20948 75748
rect 20812 73420 20948 73460
rect 20812 68984 20852 73420
rect 20812 68935 20852 68944
rect 20908 73352 20948 73361
rect 20716 68095 20756 68104
rect 20812 68816 20852 68825
rect 20812 67052 20852 68776
rect 20908 68564 20948 73312
rect 21004 72512 21044 79612
rect 21100 75536 21140 82636
rect 21196 77552 21236 83560
rect 21292 79904 21332 83980
rect 21388 83096 21428 88768
rect 21484 87464 21524 88936
rect 21484 87415 21524 87424
rect 21388 83047 21428 83056
rect 21484 87296 21524 87305
rect 21388 81836 21428 81845
rect 21388 80660 21428 81796
rect 21388 80611 21428 80620
rect 21484 80576 21524 87256
rect 21484 80527 21524 80536
rect 21292 79864 21524 79904
rect 21388 79736 21428 79745
rect 21196 77503 21236 77512
rect 21292 77720 21332 77729
rect 21100 75487 21140 75496
rect 21196 76712 21236 76721
rect 21100 74948 21140 74957
rect 21100 73016 21140 74908
rect 21196 74024 21236 76672
rect 21292 75032 21332 77680
rect 21388 76796 21428 79696
rect 21388 76747 21428 76756
rect 21292 74983 21332 74992
rect 21388 76628 21428 76637
rect 21196 73975 21236 73984
rect 21292 74276 21332 74285
rect 21100 72967 21140 72976
rect 21196 73436 21236 73445
rect 21004 72463 21044 72472
rect 21100 72848 21140 72857
rect 21100 72008 21140 72808
rect 21100 71959 21140 71968
rect 21100 71252 21140 71261
rect 20908 68515 20948 68524
rect 21004 69824 21044 69833
rect 21004 68396 21044 69784
rect 20812 67003 20852 67012
rect 20908 68356 21044 68396
rect 20620 62467 20660 62476
rect 20716 66968 20756 66977
rect 20620 62348 20660 62357
rect 20620 57392 20660 62308
rect 20716 61844 20756 66928
rect 20908 64616 20948 68356
rect 20908 64567 20948 64576
rect 21004 68144 21044 68153
rect 20908 64448 20948 64457
rect 20812 64028 20852 64037
rect 20812 63104 20852 63988
rect 20812 63055 20852 63064
rect 20716 61795 20756 61804
rect 20812 62936 20852 62945
rect 20716 60416 20756 60425
rect 20716 57896 20756 60376
rect 20716 57847 20756 57856
rect 20620 57343 20660 57352
rect 20716 56972 20756 56981
rect 20620 55292 20660 55301
rect 20620 54368 20660 55252
rect 20716 54872 20756 56932
rect 20812 56888 20852 62896
rect 20908 62348 20948 64408
rect 20908 62299 20948 62308
rect 20812 56839 20852 56848
rect 20908 62180 20948 62189
rect 20908 56384 20948 62140
rect 21004 61256 21044 68104
rect 21100 64952 21140 71212
rect 21196 69908 21236 73396
rect 21196 69859 21236 69868
rect 21100 64903 21140 64912
rect 21196 69740 21236 69749
rect 21100 64784 21140 64793
rect 21100 63944 21140 64744
rect 21100 63895 21140 63904
rect 21196 63440 21236 69700
rect 21292 67472 21332 74236
rect 21388 69488 21428 76588
rect 21484 73184 21524 79864
rect 21484 73135 21524 73144
rect 21388 69439 21428 69448
rect 21484 72764 21524 72773
rect 21292 67423 21332 67432
rect 21388 68228 21428 68237
rect 21196 63391 21236 63400
rect 21292 66380 21332 66389
rect 21100 63104 21140 63113
rect 21100 61928 21140 63064
rect 21100 61879 21140 61888
rect 21196 62516 21236 62525
rect 21004 61207 21044 61216
rect 21100 61760 21140 61769
rect 21004 61088 21044 61097
rect 21004 57812 21044 61048
rect 21100 58400 21140 61720
rect 21196 61424 21236 62476
rect 21196 61375 21236 61384
rect 21100 58351 21140 58360
rect 21196 61172 21236 61181
rect 21004 57772 21140 57812
rect 20908 56335 20948 56344
rect 21004 56216 21044 56225
rect 20716 54823 20756 54832
rect 20812 55460 20852 55469
rect 20620 54319 20660 54328
rect 20812 53360 20852 55420
rect 20812 53311 20852 53320
rect 20908 55376 20948 55385
rect 20524 53260 20660 53300
rect 19948 53068 20084 53108
rect 19948 52604 19988 53068
rect 20048 52940 20416 52949
rect 20088 52900 20130 52940
rect 20170 52900 20212 52940
rect 20252 52900 20294 52940
rect 20334 52900 20376 52940
rect 20048 52891 20416 52900
rect 19948 52555 19988 52564
rect 20140 52520 20180 52529
rect 20140 52385 20180 52480
rect 20428 52352 20468 52361
rect 20140 51848 20180 51857
rect 20140 51713 20180 51808
rect 20428 51848 20468 52312
rect 20428 51799 20468 51808
rect 20048 51428 20416 51437
rect 20088 51388 20130 51428
rect 20170 51388 20212 51428
rect 20252 51388 20294 51428
rect 20334 51388 20376 51428
rect 20048 51379 20416 51388
rect 20236 50756 20276 50765
rect 20236 50336 20276 50716
rect 20236 50287 20276 50296
rect 20524 50168 20564 50177
rect 20048 49916 20416 49925
rect 20088 49876 20130 49916
rect 20170 49876 20212 49916
rect 20252 49876 20294 49916
rect 20334 49876 20376 49916
rect 20048 49867 20416 49876
rect 19948 49496 19988 49505
rect 19948 44876 19988 49456
rect 20428 49328 20468 49337
rect 20428 48908 20468 49288
rect 20428 48859 20468 48868
rect 20524 48824 20564 50128
rect 20524 48775 20564 48784
rect 20048 48404 20416 48413
rect 20088 48364 20130 48404
rect 20170 48364 20212 48404
rect 20252 48364 20294 48404
rect 20334 48364 20376 48404
rect 20048 48355 20416 48364
rect 20140 47984 20180 47993
rect 20140 47849 20180 47944
rect 20524 47228 20564 47237
rect 20048 46892 20416 46901
rect 20088 46852 20130 46892
rect 20170 46852 20212 46892
rect 20252 46852 20294 46892
rect 20334 46852 20376 46892
rect 20048 46843 20416 46852
rect 20524 46640 20564 47188
rect 20428 46600 20564 46640
rect 20140 46472 20180 46481
rect 20140 46337 20180 46432
rect 20428 45632 20468 46600
rect 20620 46556 20660 53260
rect 20908 52856 20948 55336
rect 21004 53864 21044 56176
rect 21004 53815 21044 53824
rect 20908 52807 20948 52816
rect 21100 51008 21140 57772
rect 21196 51092 21236 61132
rect 21292 59912 21332 66340
rect 21388 65792 21428 68188
rect 21484 65960 21524 72724
rect 21484 65911 21524 65920
rect 21388 65752 21524 65792
rect 21388 65204 21428 65213
rect 21388 61424 21428 65164
rect 21388 61375 21428 61384
rect 21292 59863 21332 59872
rect 21388 61256 21428 61265
rect 21196 51043 21236 51052
rect 21292 59240 21332 59249
rect 21100 50959 21140 50968
rect 20716 50840 20756 50849
rect 20716 50336 20756 50800
rect 20716 50287 20756 50296
rect 21292 48992 21332 59200
rect 20524 46516 20660 46556
rect 20716 48952 21332 48992
rect 20524 45884 20564 46516
rect 20524 45835 20564 45844
rect 20620 46388 20660 46397
rect 20620 45800 20660 46348
rect 20620 45751 20660 45760
rect 20428 45592 20660 45632
rect 20524 45464 20564 45473
rect 20048 45380 20416 45389
rect 20088 45340 20130 45380
rect 20170 45340 20212 45380
rect 20252 45340 20294 45380
rect 20334 45340 20376 45380
rect 20048 45331 20416 45340
rect 19948 44827 19988 44836
rect 20140 45044 20180 45053
rect 20140 44456 20180 45004
rect 20140 44407 20180 44416
rect 20048 43868 20416 43877
rect 20088 43828 20130 43868
rect 20170 43828 20212 43868
rect 20252 43828 20294 43868
rect 20334 43828 20376 43868
rect 20048 43819 20416 43828
rect 20524 43448 20564 45424
rect 20524 43399 20564 43408
rect 20620 43280 20660 45592
rect 20620 43231 20660 43240
rect 19564 38368 19700 38408
rect 19756 43180 19892 43220
rect 19564 35468 19604 38368
rect 19564 35419 19604 35428
rect 19660 38240 19700 38249
rect 19468 34243 19508 34252
rect 19564 35300 19604 35309
rect 19468 34124 19508 34133
rect 19468 33284 19508 34084
rect 19564 33452 19604 35260
rect 19660 34544 19700 38200
rect 19660 34495 19700 34504
rect 19660 34376 19700 34385
rect 19660 33620 19700 34336
rect 19660 33571 19700 33580
rect 19564 33403 19604 33412
rect 19756 33368 19796 43180
rect 20524 42776 20564 42785
rect 20048 42356 20416 42365
rect 20088 42316 20130 42356
rect 20170 42316 20212 42356
rect 20252 42316 20294 42356
rect 20334 42316 20376 42356
rect 20048 42307 20416 42316
rect 20524 42188 20564 42736
rect 20524 42139 20564 42148
rect 20620 42272 20660 42281
rect 20524 41432 20564 41441
rect 20044 41180 20084 41189
rect 19948 41140 20044 41180
rect 19852 40340 19892 40349
rect 19852 39164 19892 40300
rect 19948 39920 19988 41140
rect 20044 41131 20084 41140
rect 20048 40844 20416 40853
rect 20088 40804 20130 40844
rect 20170 40804 20212 40844
rect 20252 40804 20294 40844
rect 20334 40804 20376 40844
rect 20048 40795 20416 40804
rect 19948 39871 19988 39880
rect 20044 40676 20084 40685
rect 20044 39836 20084 40636
rect 20140 40508 20180 40517
rect 20140 39920 20180 40468
rect 20140 39871 20180 39880
rect 20044 39787 20084 39796
rect 20048 39332 20416 39341
rect 20088 39292 20130 39332
rect 20170 39292 20212 39332
rect 20252 39292 20294 39332
rect 20334 39292 20376 39332
rect 20048 39283 20416 39292
rect 19852 39124 20084 39164
rect 19948 38744 19988 38753
rect 19852 38660 19892 38669
rect 19852 34544 19892 38620
rect 19948 37484 19988 38704
rect 20044 37988 20084 39124
rect 20524 38324 20564 41392
rect 20620 41348 20660 42232
rect 20620 41299 20660 41308
rect 20044 37939 20084 37948
rect 20428 38284 20564 38324
rect 20620 39248 20660 39257
rect 20428 37988 20468 38284
rect 20428 37939 20468 37948
rect 20524 38156 20564 38165
rect 20048 37820 20416 37829
rect 20088 37780 20130 37820
rect 20170 37780 20212 37820
rect 20252 37780 20294 37820
rect 20334 37780 20376 37820
rect 20048 37771 20416 37780
rect 19948 37435 19988 37444
rect 20044 37652 20084 37661
rect 19852 34495 19892 34504
rect 19948 37148 19988 37157
rect 19852 34124 19892 34133
rect 19852 33536 19892 34084
rect 19948 34124 19988 37108
rect 20044 36476 20084 37612
rect 20428 37652 20468 37661
rect 20428 36476 20468 37612
rect 20524 36896 20564 38116
rect 20524 36847 20564 36856
rect 20428 36436 20564 36476
rect 20044 36427 20084 36436
rect 20048 36308 20416 36317
rect 20088 36268 20130 36308
rect 20170 36268 20212 36308
rect 20252 36268 20294 36308
rect 20334 36268 20376 36308
rect 20048 36259 20416 36268
rect 20044 36140 20084 36149
rect 20044 34964 20084 36100
rect 20524 35384 20564 36436
rect 20044 34915 20084 34924
rect 20428 35344 20564 35384
rect 20428 34964 20468 35344
rect 20428 34915 20468 34924
rect 20524 35216 20564 35225
rect 20048 34796 20416 34805
rect 20088 34756 20130 34796
rect 20170 34756 20212 34796
rect 20252 34756 20294 34796
rect 20334 34756 20376 34796
rect 20048 34747 20416 34756
rect 19948 34075 19988 34084
rect 20044 34628 20084 34637
rect 20044 34460 20084 34588
rect 20140 34544 20180 34572
rect 20180 34504 20276 34544
rect 20140 34495 20180 34504
rect 19852 33487 19892 33496
rect 19948 33452 19988 33461
rect 19756 33319 19796 33328
rect 19852 33368 19892 33377
rect 19468 33244 19604 33284
rect 19372 30799 19412 30808
rect 19468 32696 19508 32705
rect 19468 31772 19508 32656
rect 19564 32360 19604 33244
rect 19756 33200 19796 33209
rect 19564 32311 19604 32320
rect 19660 32696 19700 32705
rect 19468 31436 19508 31732
rect 19372 30680 19412 30689
rect 19372 30545 19412 30640
rect 19276 29968 19412 30008
rect 19180 29623 19220 29632
rect 19276 29840 19316 29849
rect 18808 29504 19176 29513
rect 18848 29464 18890 29504
rect 18930 29464 18972 29504
rect 19012 29464 19054 29504
rect 19094 29464 19136 29504
rect 18808 29455 19176 29464
rect 19180 29336 19220 29345
rect 19180 28412 19220 29296
rect 19276 28580 19316 29800
rect 19276 28531 19316 28540
rect 19180 28372 19316 28412
rect 18808 27992 19176 28001
rect 18848 27952 18890 27992
rect 18930 27952 18972 27992
rect 19012 27952 19054 27992
rect 19094 27952 19136 27992
rect 18808 27943 19176 27952
rect 19276 27992 19316 28372
rect 19276 27943 19316 27952
rect 18892 27824 18932 27833
rect 18700 26767 18740 26776
rect 18796 27068 18836 27077
rect 18796 26648 18836 27028
rect 18892 26816 18932 27784
rect 18892 26767 18932 26776
rect 19180 27572 19220 27581
rect 19180 26732 19220 27532
rect 19180 26683 19220 26692
rect 19276 27404 19316 27413
rect 18604 25388 18644 26020
rect 18604 24632 18644 25348
rect 18604 24583 18644 24592
rect 18700 26608 18836 26648
rect 18700 23960 18740 26608
rect 18808 26480 19176 26489
rect 18848 26440 18890 26480
rect 18930 26440 18972 26480
rect 19012 26440 19054 26480
rect 19094 26440 19136 26480
rect 18808 26431 19176 26440
rect 18796 26312 18836 26321
rect 18796 26060 18836 26272
rect 18796 26011 18836 26020
rect 18796 25808 18836 25817
rect 18796 25472 18836 25768
rect 18796 25423 18836 25432
rect 18808 24968 19176 24977
rect 18848 24928 18890 24968
rect 18930 24928 18972 24968
rect 19012 24928 19054 24968
rect 19094 24928 19136 24968
rect 18808 24919 19176 24928
rect 19276 24800 19316 27364
rect 19372 26900 19412 29968
rect 19468 27404 19508 31396
rect 19564 32192 19604 32201
rect 19564 30848 19604 32152
rect 19564 30799 19604 30808
rect 19564 30680 19604 30689
rect 19564 29840 19604 30640
rect 19564 29791 19604 29800
rect 19660 29252 19700 32656
rect 19756 30848 19796 33160
rect 19756 30799 19796 30808
rect 19756 30680 19796 30689
rect 19756 30596 19796 30640
rect 19756 30545 19796 30556
rect 19756 30176 19796 30185
rect 19756 29840 19796 30136
rect 19852 30092 19892 33328
rect 19948 32948 19988 33412
rect 20044 33452 20084 34420
rect 20140 34376 20180 34385
rect 20140 34241 20180 34336
rect 20140 34124 20180 34133
rect 20236 34124 20276 34504
rect 20180 34084 20276 34124
rect 20140 34056 20180 34084
rect 20044 33403 20084 33412
rect 20048 33284 20416 33293
rect 20088 33244 20130 33284
rect 20170 33244 20212 33284
rect 20252 33244 20294 33284
rect 20334 33244 20376 33284
rect 20048 33235 20416 33244
rect 20524 33140 20564 35176
rect 20620 34544 20660 39208
rect 20620 34495 20660 34504
rect 20620 33788 20660 33797
rect 20620 33452 20660 33748
rect 20620 33403 20660 33412
rect 20140 33116 20276 33140
rect 20180 33100 20276 33116
rect 20140 33067 20180 33076
rect 19948 32899 19988 32908
rect 20044 33032 20084 33041
rect 19948 32780 19988 32789
rect 19948 32276 19988 32740
rect 19948 32227 19988 32236
rect 20044 31940 20084 32992
rect 20236 32024 20276 33100
rect 20236 31975 20276 31984
rect 20332 33116 20372 33125
rect 19948 31900 20084 31940
rect 20332 31940 20372 33076
rect 20428 33100 20564 33140
rect 20620 33200 20660 33209
rect 20428 32444 20468 33100
rect 20620 32864 20660 33160
rect 20428 32395 20468 32404
rect 20524 32824 20660 32864
rect 20524 32108 20564 32824
rect 20524 32059 20564 32068
rect 20620 32696 20660 32705
rect 20332 31900 20564 31940
rect 19948 30092 19988 31900
rect 20048 31772 20416 31781
rect 20088 31732 20130 31772
rect 20170 31732 20212 31772
rect 20252 31732 20294 31772
rect 20334 31732 20376 31772
rect 20048 31723 20416 31732
rect 20428 31604 20468 31613
rect 20044 31520 20084 31560
rect 20044 31436 20084 31480
rect 20044 30512 20084 31396
rect 20140 30680 20180 30689
rect 20140 30545 20180 30640
rect 20044 30463 20084 30472
rect 20428 30512 20468 31564
rect 20428 30463 20468 30472
rect 20048 30260 20416 30269
rect 20088 30220 20130 30260
rect 20170 30220 20212 30260
rect 20252 30220 20294 30260
rect 20334 30220 20376 30260
rect 20048 30211 20416 30220
rect 19948 30052 20084 30092
rect 19852 30043 19892 30052
rect 19756 29791 19796 29800
rect 19948 29924 19988 29933
rect 19564 29212 19700 29252
rect 19564 28160 19604 29212
rect 19564 28111 19604 28120
rect 19660 29084 19700 29093
rect 19468 27355 19508 27364
rect 19564 27992 19604 28001
rect 19372 26851 19412 26860
rect 19468 27236 19508 27245
rect 19276 24751 19316 24760
rect 19372 25892 19412 25901
rect 19276 24632 19316 24641
rect 18700 23911 18740 23920
rect 18796 24380 18836 24389
rect 18796 23876 18836 24340
rect 18988 24296 19028 24305
rect 18988 23960 19028 24256
rect 18988 23911 19028 23920
rect 18796 23827 18836 23836
rect 18316 19088 18356 22072
rect 18412 23204 18452 23213
rect 18412 20936 18452 23164
rect 18508 22448 18548 23668
rect 18604 23792 18644 23801
rect 18604 23657 18644 23752
rect 18700 23708 18740 23717
rect 18508 22399 18548 22408
rect 18604 23456 18644 23465
rect 18412 20887 18452 20896
rect 18508 22280 18548 22289
rect 18508 21608 18548 22240
rect 18316 19039 18356 19048
rect 18412 20348 18452 20357
rect 18220 18115 18260 18124
rect 18316 18416 18356 18425
rect 18412 18416 18452 20308
rect 18508 20264 18548 21568
rect 18508 20215 18548 20224
rect 18356 18376 18452 18416
rect 18508 20096 18548 20105
rect 18508 19340 18548 20056
rect 18508 18836 18548 19300
rect 18124 17359 18164 17368
rect 18220 17996 18260 18005
rect 18028 17324 18068 17333
rect 18028 14720 18068 17284
rect 18124 16316 18164 16325
rect 18124 15728 18164 16276
rect 18124 15679 18164 15688
rect 18028 10604 18068 14680
rect 18124 15476 18164 15485
rect 18124 14888 18164 15436
rect 18220 15308 18260 17956
rect 18220 15259 18260 15268
rect 18316 16988 18356 18376
rect 18124 13964 18164 14848
rect 18220 14972 18260 14981
rect 18220 14837 18260 14932
rect 18124 13915 18164 13924
rect 18220 14720 18260 14729
rect 18316 14720 18356 16948
rect 18412 18164 18452 18173
rect 18412 15140 18452 18124
rect 18508 16316 18548 18796
rect 18604 17912 18644 23416
rect 18700 22532 18740 23668
rect 18808 23456 19176 23465
rect 18848 23416 18890 23456
rect 18930 23416 18972 23456
rect 19012 23416 19054 23456
rect 19094 23416 19136 23456
rect 18808 23407 19176 23416
rect 18892 23288 18932 23297
rect 18796 23204 18836 23215
rect 18796 23120 18836 23164
rect 18796 23071 18836 23080
rect 18892 23036 18932 23248
rect 19180 23204 19220 23213
rect 18892 22616 18932 22996
rect 18892 22567 18932 22576
rect 19084 23120 19124 23129
rect 18700 22483 18740 22492
rect 18700 22364 18740 22373
rect 18700 21356 18740 22324
rect 18892 22364 18932 22373
rect 18796 22196 18836 22291
rect 18892 22229 18932 22324
rect 18796 22147 18836 22156
rect 19084 22196 19124 23080
rect 19180 22364 19220 23164
rect 19180 22315 19220 22324
rect 19084 22147 19124 22156
rect 18808 21944 19176 21953
rect 18848 21904 18890 21944
rect 18930 21904 18972 21944
rect 19012 21904 19054 21944
rect 19094 21904 19136 21944
rect 18808 21895 19176 21904
rect 18700 18584 18740 21316
rect 18988 21524 19028 21533
rect 18988 20600 19028 21484
rect 19180 21524 19220 21533
rect 19180 21389 19220 21484
rect 18988 20551 19028 20560
rect 18808 20432 19176 20441
rect 18848 20392 18890 20432
rect 18930 20392 18972 20432
rect 19012 20392 19054 20432
rect 19094 20392 19136 20432
rect 18808 20383 19176 20392
rect 19084 20264 19124 20273
rect 19084 20096 19124 20224
rect 18892 20012 18932 20021
rect 18892 19340 18932 19972
rect 19084 20012 19124 20056
rect 19084 19932 19124 19972
rect 19180 20264 19220 20273
rect 18892 19205 18932 19300
rect 19180 19340 19220 20224
rect 19180 19291 19220 19300
rect 18808 18920 19176 18929
rect 18848 18880 18890 18920
rect 18930 18880 18972 18920
rect 19012 18880 19054 18920
rect 19094 18880 19136 18920
rect 18808 18871 19176 18880
rect 18700 18535 18740 18544
rect 18796 18752 18836 18761
rect 18796 18416 18836 18712
rect 18604 17863 18644 17872
rect 18700 18376 18836 18416
rect 19180 18752 19220 18761
rect 18604 17744 18644 17753
rect 18604 17408 18644 17704
rect 18604 17359 18644 17368
rect 18508 15560 18548 16276
rect 18700 16232 18740 18376
rect 19180 17660 19220 18712
rect 19276 18500 19316 24592
rect 19372 24212 19412 25852
rect 19468 24548 19508 27196
rect 19564 27152 19604 27952
rect 19564 27103 19604 27112
rect 19660 27068 19700 29044
rect 19852 28664 19892 28673
rect 19660 27019 19700 27028
rect 19756 27152 19796 27161
rect 19468 24499 19508 24508
rect 19564 26984 19604 26993
rect 19372 24163 19412 24172
rect 19372 24044 19412 24053
rect 19412 24004 19508 24044
rect 19372 23995 19412 24004
rect 19372 23792 19412 23801
rect 19372 21860 19412 23752
rect 19372 21811 19412 21820
rect 19372 21608 19412 21617
rect 19372 19256 19412 21568
rect 19372 19207 19412 19216
rect 19468 18668 19508 24004
rect 19564 23288 19604 26944
rect 19660 26900 19700 26909
rect 19660 25052 19700 26860
rect 19660 25003 19700 25012
rect 19756 24296 19796 27112
rect 19852 24800 19892 28624
rect 19948 28580 19988 29884
rect 20044 28916 20084 30052
rect 20428 29672 20468 29681
rect 20428 28916 20468 29632
rect 20524 29168 20564 31900
rect 20620 29336 20660 32656
rect 20620 29287 20660 29296
rect 20524 29119 20564 29128
rect 20428 28876 20564 28916
rect 20044 28867 20084 28876
rect 20048 28748 20416 28757
rect 20088 28708 20130 28748
rect 20170 28708 20212 28748
rect 20252 28708 20294 28748
rect 20334 28708 20376 28748
rect 20048 28699 20416 28708
rect 19948 28531 19988 28540
rect 20140 28412 20180 28421
rect 19852 24751 19892 24760
rect 19948 28160 19988 28169
rect 19948 24548 19988 28120
rect 20140 27992 20180 28372
rect 20140 27943 20180 27952
rect 20044 27740 20084 27749
rect 20044 27404 20084 27700
rect 20524 27488 20564 28876
rect 20524 27439 20564 27448
rect 20620 28244 20660 28253
rect 20044 27355 20084 27364
rect 20048 27236 20416 27245
rect 20088 27196 20130 27236
rect 20170 27196 20212 27236
rect 20252 27196 20294 27236
rect 20334 27196 20376 27236
rect 20048 27187 20416 27196
rect 20044 27068 20084 27077
rect 20044 26060 20084 27028
rect 20044 25925 20084 26020
rect 20524 26228 20564 26237
rect 20048 25724 20416 25733
rect 20088 25684 20130 25724
rect 20170 25684 20212 25724
rect 20252 25684 20294 25724
rect 20334 25684 20376 25724
rect 20048 25675 20416 25684
rect 20524 25640 20564 26188
rect 20524 25591 20564 25600
rect 20524 25472 20564 25481
rect 19948 24499 19988 24508
rect 20044 25052 20084 25061
rect 19756 24247 19796 24256
rect 19852 24464 19892 24473
rect 19564 23239 19604 23248
rect 19660 23876 19700 23885
rect 19564 22868 19604 22877
rect 19564 22448 19604 22828
rect 19564 21524 19604 22408
rect 19660 22280 19700 23836
rect 19756 23624 19796 23633
rect 19756 22364 19796 23584
rect 19852 23624 19892 24424
rect 20044 24380 20084 25012
rect 20140 24884 20180 24893
rect 20140 24749 20180 24844
rect 19948 24340 20084 24380
rect 20524 24380 20564 25432
rect 20620 24632 20660 28204
rect 20716 28076 20756 48952
rect 21100 48824 21140 48833
rect 20812 48572 20852 48581
rect 20812 44120 20852 48532
rect 21004 45632 21044 45641
rect 21004 44288 21044 45592
rect 21004 44239 21044 44248
rect 20812 44080 21044 44120
rect 20908 43280 20948 43289
rect 20812 42692 20852 42701
rect 20812 35972 20852 42652
rect 20908 37988 20948 43240
rect 21004 41600 21044 44080
rect 21004 41551 21044 41560
rect 21100 41516 21140 48784
rect 21100 41467 21140 41476
rect 21196 45296 21236 45305
rect 21100 40676 21140 40685
rect 20908 37939 20948 37948
rect 21004 39080 21044 39089
rect 21004 37736 21044 39040
rect 21004 37687 21044 37696
rect 21004 37400 21044 37409
rect 20812 35923 20852 35932
rect 20908 36224 20948 36233
rect 20716 28027 20756 28036
rect 20812 35804 20852 35813
rect 20716 27908 20756 27917
rect 20716 25304 20756 27868
rect 20812 27320 20852 35764
rect 20908 30848 20948 36184
rect 21004 34880 21044 37360
rect 21100 35972 21140 40636
rect 21100 35923 21140 35932
rect 21196 35804 21236 45256
rect 21292 44960 21332 44969
rect 21292 44825 21332 44920
rect 21388 43220 21428 61216
rect 21484 60920 21524 65752
rect 21484 60871 21524 60880
rect 21292 43180 21428 43220
rect 21484 45632 21524 45641
rect 21292 40592 21332 43180
rect 21292 40543 21332 40552
rect 21388 41936 21428 41945
rect 21292 39500 21332 39509
rect 21292 37400 21332 39460
rect 21292 37351 21332 37360
rect 21196 35755 21236 35764
rect 21292 37232 21332 37241
rect 21100 35720 21140 35729
rect 21100 35300 21140 35680
rect 21100 35251 21140 35260
rect 21004 34840 21236 34880
rect 20908 30799 20948 30808
rect 21004 34712 21044 34721
rect 20908 30596 20948 30605
rect 20908 28244 20948 30556
rect 21004 30092 21044 34672
rect 21100 34208 21140 34217
rect 21100 30764 21140 34168
rect 21196 33452 21236 34840
rect 21292 34292 21332 37192
rect 21292 34243 21332 34252
rect 21196 33403 21236 33412
rect 21196 33284 21236 33293
rect 21196 31940 21236 33244
rect 21388 33140 21428 41896
rect 21484 33368 21524 45592
rect 21484 33319 21524 33328
rect 21196 31891 21236 31900
rect 21292 33100 21428 33140
rect 21484 33200 21524 33209
rect 21100 30715 21140 30724
rect 21004 30043 21044 30052
rect 21100 30176 21140 30185
rect 20908 28195 20948 28204
rect 21004 29168 21044 29177
rect 20812 27271 20852 27280
rect 20908 27992 20948 28001
rect 20716 25255 20756 25264
rect 20812 26060 20852 26069
rect 20620 24583 20660 24592
rect 20716 25136 20756 25145
rect 20524 24340 20660 24380
rect 19948 23792 19988 24340
rect 20048 24212 20416 24221
rect 20088 24172 20130 24212
rect 20170 24172 20212 24212
rect 20252 24172 20294 24212
rect 20334 24172 20376 24212
rect 20048 24163 20416 24172
rect 20524 23876 20564 23885
rect 19948 23752 20084 23792
rect 19852 23036 19892 23584
rect 19852 22987 19892 22996
rect 19948 23624 19988 23633
rect 19852 22784 19892 22793
rect 19852 22532 19892 22744
rect 19852 22483 19892 22492
rect 19948 22448 19988 23584
rect 20044 23372 20084 23752
rect 20044 23323 20084 23332
rect 20048 22700 20416 22709
rect 20088 22660 20130 22700
rect 20170 22660 20212 22700
rect 20252 22660 20294 22700
rect 20334 22660 20376 22700
rect 20048 22651 20416 22660
rect 19948 22399 19988 22408
rect 19852 22364 19892 22373
rect 19756 22324 19852 22364
rect 19852 22315 19892 22324
rect 19948 22280 19988 22291
rect 19660 22240 19796 22280
rect 19564 21475 19604 21484
rect 19660 22112 19700 22121
rect 19564 20852 19604 20861
rect 19564 20180 19604 20812
rect 19564 18752 19604 20140
rect 19564 18703 19604 18712
rect 19468 18619 19508 18628
rect 19276 18460 19604 18500
rect 19372 18080 19412 18089
rect 19180 17611 19220 17620
rect 19276 17828 19316 17837
rect 18808 17408 19176 17417
rect 18848 17368 18890 17408
rect 18930 17368 18972 17408
rect 19012 17368 19054 17408
rect 19094 17368 19136 17408
rect 18808 17359 19176 17368
rect 19276 17240 19316 17788
rect 19276 17191 19316 17200
rect 19372 16400 19412 18040
rect 19372 16351 19412 16360
rect 19468 17576 19508 17585
rect 18700 16183 18740 16192
rect 18892 16316 18932 16325
rect 18892 16064 18932 16276
rect 18508 15511 18548 15520
rect 18700 16024 18932 16064
rect 18700 15476 18740 16024
rect 18808 15896 19176 15905
rect 18848 15856 18890 15896
rect 18930 15856 18972 15896
rect 19012 15856 19054 15896
rect 19094 15856 19136 15896
rect 18808 15847 19176 15856
rect 18700 15427 18740 15436
rect 19372 15476 19412 15485
rect 18412 15091 18452 15100
rect 18508 15392 18548 15401
rect 18260 14680 18356 14720
rect 18124 13208 18164 13217
rect 18124 12452 18164 13168
rect 18220 13040 18260 14680
rect 18508 14216 18548 15352
rect 18508 14167 18548 14176
rect 18604 15140 18644 15149
rect 18508 14048 18548 14057
rect 18220 12991 18260 13000
rect 18316 13376 18356 13385
rect 18124 12403 18164 12412
rect 18220 12872 18260 12881
rect 18028 10436 18068 10564
rect 18028 10387 18068 10396
rect 18124 11528 18164 11537
rect 18124 10268 18164 11488
rect 18028 10228 18164 10268
rect 18028 7916 18068 10228
rect 18124 9848 18164 9857
rect 18124 9260 18164 9808
rect 18124 9211 18164 9220
rect 18220 9680 18260 12832
rect 18316 11948 18356 13336
rect 18316 11899 18356 11908
rect 18412 13292 18452 13301
rect 18412 12536 18452 13252
rect 18124 8924 18164 8933
rect 18124 8000 18164 8884
rect 18124 7951 18164 7960
rect 18028 7867 18068 7876
rect 17356 2071 17396 2080
rect 17644 2860 17972 2900
rect 18124 7160 18164 7169
rect 16492 1903 16532 1912
rect 17356 1952 17396 1961
rect 15436 1616 15476 1625
rect 15436 80 15476 1576
rect 16396 1448 16436 1457
rect 16012 1280 16052 1289
rect 15820 1196 15860 1205
rect 15628 608 15668 617
rect 15628 80 15668 568
rect 15820 80 15860 1156
rect 16012 80 16052 1240
rect 16204 272 16244 281
rect 16204 80 16244 232
rect 16396 80 16436 1408
rect 16780 1364 16820 1373
rect 16588 440 16628 449
rect 16588 80 16628 400
rect 16780 80 16820 1324
rect 17164 860 17204 869
rect 16972 188 17012 197
rect 16972 80 17012 148
rect 17164 80 17204 820
rect 17356 80 17396 1912
rect 17644 1532 17684 2860
rect 17644 1483 17684 1492
rect 17740 2204 17780 2213
rect 17548 356 17588 365
rect 17548 80 17588 316
rect 17740 80 17780 2164
rect 17932 1028 17972 1037
rect 17932 80 17972 988
rect 18124 80 18164 7120
rect 18220 6404 18260 9640
rect 18220 6355 18260 6364
rect 18316 11360 18356 11369
rect 18316 4304 18356 11320
rect 18412 10352 18452 12496
rect 18508 12452 18548 14008
rect 18604 12536 18644 15100
rect 18808 14384 19176 14393
rect 18848 14344 18890 14384
rect 18930 14344 18972 14384
rect 19012 14344 19054 14384
rect 19094 14344 19136 14384
rect 18808 14335 19176 14344
rect 19372 14048 19412 15436
rect 19372 13999 19412 14008
rect 18700 13544 18740 13553
rect 18700 12788 18740 13504
rect 19276 13544 19316 13553
rect 18808 12872 19176 12881
rect 18848 12832 18890 12872
rect 18930 12832 18972 12872
rect 19012 12832 19054 12872
rect 19094 12832 19136 12872
rect 18808 12823 19176 12832
rect 18700 12739 18740 12748
rect 19276 12620 19316 13504
rect 19276 12571 19316 12580
rect 18604 12487 18644 12496
rect 18508 12317 18548 12412
rect 19372 12452 19412 12461
rect 18508 11780 18548 11789
rect 18508 11528 18548 11740
rect 18508 11479 18548 11488
rect 18700 11612 18740 11621
rect 18700 10940 18740 11572
rect 18808 11360 19176 11369
rect 18848 11320 18890 11360
rect 18930 11320 18972 11360
rect 19012 11320 19054 11360
rect 19094 11320 19136 11360
rect 18808 11311 19176 11320
rect 19372 11192 19412 12412
rect 19372 11143 19412 11152
rect 18700 10891 18740 10900
rect 18412 9512 18452 10312
rect 18604 10436 18644 10445
rect 18412 8840 18452 9472
rect 18412 8791 18452 8800
rect 18508 10268 18548 10277
rect 18508 8168 18548 10228
rect 18508 8119 18548 8128
rect 18604 9344 18644 10396
rect 18700 10184 18740 10193
rect 18700 9428 18740 10144
rect 19276 10100 19316 10109
rect 18808 9848 19176 9857
rect 18848 9808 18890 9848
rect 18930 9808 18972 9848
rect 19012 9808 19054 9848
rect 19094 9808 19136 9848
rect 18808 9799 19176 9808
rect 18700 9379 18740 9388
rect 18604 5228 18644 9304
rect 19180 9260 19220 9269
rect 18700 9092 18740 9101
rect 18700 8084 18740 9052
rect 19180 8672 19220 9220
rect 19276 8924 19316 10060
rect 19276 8875 19316 8884
rect 19180 8623 19220 8632
rect 19372 8756 19412 8765
rect 18808 8336 19176 8345
rect 18848 8296 18890 8336
rect 18930 8296 18972 8336
rect 19012 8296 19054 8336
rect 19094 8296 19136 8336
rect 18808 8287 19176 8296
rect 18700 8035 18740 8044
rect 19372 7916 19412 8716
rect 18700 7664 18740 7673
rect 18700 7244 18740 7624
rect 18700 5732 18740 7204
rect 18808 6824 19176 6833
rect 18848 6784 18890 6824
rect 18930 6784 18972 6824
rect 19012 6784 19054 6824
rect 19094 6784 19136 6824
rect 18808 6775 19176 6784
rect 19372 6404 19412 7876
rect 19372 6355 19412 6364
rect 18700 5683 18740 5692
rect 18808 5312 19176 5321
rect 18848 5272 18890 5312
rect 18930 5272 18972 5312
rect 19012 5272 19054 5312
rect 19094 5272 19136 5312
rect 18808 5263 19176 5272
rect 18604 5179 18644 5188
rect 18316 4255 18356 4264
rect 18808 3800 19176 3809
rect 18848 3760 18890 3800
rect 18930 3760 18972 3800
rect 19012 3760 19054 3800
rect 19094 3760 19136 3800
rect 18808 3751 19176 3760
rect 18700 3212 18740 3221
rect 18700 3077 18740 3172
rect 18700 2540 18740 2549
rect 18700 1364 18740 2500
rect 18808 2288 19176 2297
rect 18848 2248 18890 2288
rect 18930 2248 18972 2288
rect 19012 2248 19054 2288
rect 19094 2248 19136 2288
rect 18808 2239 19176 2248
rect 19468 2036 19508 17536
rect 19564 16484 19604 18460
rect 19660 17744 19700 22072
rect 19756 21776 19796 22240
rect 19756 21727 19796 21736
rect 19852 22196 19892 22205
rect 19660 17695 19700 17704
rect 19756 21608 19796 21617
rect 19564 16435 19604 16444
rect 19660 17576 19700 17585
rect 19660 16316 19700 17536
rect 19756 17240 19796 21568
rect 19852 19424 19892 22156
rect 19948 22196 19988 22240
rect 20428 22280 20468 22289
rect 19948 22147 19988 22156
rect 20236 22196 20276 22205
rect 20044 21944 20084 21953
rect 20044 21524 20084 21904
rect 19948 21484 20044 21524
rect 19948 20768 19988 21484
rect 20044 21475 20084 21484
rect 20236 21356 20276 22156
rect 20428 21608 20468 22240
rect 20524 21776 20564 23836
rect 20524 21727 20564 21736
rect 20428 21568 20564 21608
rect 20236 21307 20276 21316
rect 20048 21188 20416 21197
rect 20088 21148 20130 21188
rect 20170 21148 20212 21188
rect 20252 21148 20294 21188
rect 20334 21148 20376 21188
rect 20048 21139 20416 21148
rect 20524 21020 20564 21568
rect 20428 20980 20564 21020
rect 20140 20768 20180 20777
rect 19948 20728 20084 20768
rect 19948 20600 19988 20609
rect 19948 20012 19988 20560
rect 20044 20096 20084 20728
rect 20140 20633 20180 20728
rect 20332 20684 20372 20693
rect 20044 20047 20084 20056
rect 19948 19963 19988 19972
rect 20332 20012 20372 20644
rect 20332 19963 20372 19972
rect 20044 19844 20084 19939
rect 20428 19928 20468 20980
rect 20428 19879 20468 19888
rect 20524 20600 20564 20609
rect 20044 19795 20084 19804
rect 20048 19676 20416 19685
rect 20088 19636 20130 19676
rect 20170 19636 20212 19676
rect 20252 19636 20294 19676
rect 20334 19636 20376 19676
rect 20048 19627 20416 19636
rect 20524 19592 20564 20560
rect 20524 19543 20564 19552
rect 19852 19375 19892 19384
rect 20140 19508 20180 19517
rect 20140 19373 20180 19468
rect 19948 19340 19988 19349
rect 19756 17191 19796 17200
rect 19852 19256 19892 19265
rect 19852 17072 19892 19216
rect 19948 18752 19988 19300
rect 19948 18703 19988 18712
rect 20524 19256 20564 19265
rect 20140 18584 20180 18593
rect 19660 16267 19700 16276
rect 19756 17032 19892 17072
rect 19948 18500 19988 18509
rect 19756 15896 19796 17032
rect 19756 15847 19796 15856
rect 19852 16736 19892 16745
rect 19852 14720 19892 16696
rect 19948 16064 19988 18460
rect 20140 18449 20180 18544
rect 20048 18164 20416 18173
rect 20088 18124 20130 18164
rect 20170 18124 20212 18164
rect 20252 18124 20294 18164
rect 20334 18124 20376 18164
rect 20048 18115 20416 18124
rect 20140 17744 20180 17753
rect 20140 17609 20180 17704
rect 20044 17240 20084 17249
rect 20044 17072 20084 17200
rect 20044 17023 20084 17032
rect 20140 17156 20180 17167
rect 20140 17072 20180 17116
rect 20140 17023 20180 17032
rect 20524 16820 20564 19216
rect 20524 16771 20564 16780
rect 20048 16652 20416 16661
rect 20088 16612 20130 16652
rect 20170 16612 20212 16652
rect 20252 16612 20294 16652
rect 20334 16612 20376 16652
rect 20048 16603 20416 16612
rect 19948 16015 19988 16024
rect 20524 16316 20564 16325
rect 19852 14671 19892 14680
rect 19948 15896 19988 15905
rect 19756 14552 19796 14561
rect 19564 13712 19604 13721
rect 19564 11192 19604 13672
rect 19660 13292 19700 13301
rect 19660 11612 19700 13252
rect 19660 11563 19700 11572
rect 19564 11143 19604 11152
rect 19756 11024 19796 14512
rect 19852 13460 19892 13469
rect 19852 12704 19892 13420
rect 19852 12655 19892 12664
rect 19852 11864 19892 11873
rect 19852 11729 19892 11824
rect 19948 11192 19988 15856
rect 20048 15140 20416 15149
rect 20088 15100 20130 15140
rect 20170 15100 20212 15140
rect 20252 15100 20294 15140
rect 20334 15100 20376 15140
rect 20048 15091 20416 15100
rect 20524 14972 20564 16276
rect 20620 15644 20660 24340
rect 20716 21020 20756 25096
rect 20812 24464 20852 26020
rect 20812 24415 20852 24424
rect 20716 20971 20756 20980
rect 20812 23624 20852 23633
rect 20716 19928 20756 19937
rect 20716 19256 20756 19888
rect 20716 19207 20756 19216
rect 20716 19088 20756 19097
rect 20716 16148 20756 19048
rect 20812 18668 20852 23584
rect 20908 22952 20948 27952
rect 21004 24800 21044 29128
rect 21100 25556 21140 30136
rect 21100 25507 21140 25516
rect 21196 29672 21236 29681
rect 21196 25472 21236 29632
rect 21292 27908 21332 33100
rect 21292 27859 21332 27868
rect 21388 33032 21428 33041
rect 21196 25423 21236 25432
rect 21292 27404 21332 27413
rect 21004 24751 21044 24760
rect 21100 24884 21140 24893
rect 20908 22903 20948 22912
rect 21004 24632 21044 24641
rect 21004 22784 21044 24592
rect 21100 24632 21140 24844
rect 21100 24583 21140 24592
rect 21196 23960 21236 23969
rect 20812 18619 20852 18628
rect 20908 22744 21044 22784
rect 21100 23120 21140 23129
rect 20908 17744 20948 22744
rect 20716 16099 20756 16108
rect 20812 17704 20948 17744
rect 21004 22616 21044 22625
rect 20620 15604 20756 15644
rect 20524 14923 20564 14932
rect 20620 15476 20660 15485
rect 20620 14216 20660 15436
rect 20620 14167 20660 14176
rect 20716 14048 20756 15604
rect 20812 15308 20852 17704
rect 20812 15259 20852 15268
rect 20908 17576 20948 17585
rect 20812 15056 20852 15065
rect 20812 14636 20852 15016
rect 20812 14587 20852 14596
rect 20524 14008 20756 14048
rect 20812 14048 20852 14057
rect 20048 13628 20416 13637
rect 20088 13588 20130 13628
rect 20170 13588 20212 13628
rect 20252 13588 20294 13628
rect 20334 13588 20376 13628
rect 20048 13579 20416 13588
rect 20048 12116 20416 12125
rect 20088 12076 20130 12116
rect 20170 12076 20212 12116
rect 20252 12076 20294 12116
rect 20334 12076 20376 12116
rect 20048 12067 20416 12076
rect 19948 11143 19988 11152
rect 20044 11444 20084 11453
rect 20044 11024 20084 11404
rect 19756 10975 19796 10984
rect 19948 10984 20084 11024
rect 19564 10520 19604 10529
rect 19564 8672 19604 10480
rect 19756 9428 19796 9437
rect 19564 8623 19604 8632
rect 19660 9260 19700 9269
rect 19660 7160 19700 9220
rect 19660 7111 19700 7120
rect 19564 6992 19604 7001
rect 19564 5648 19604 6952
rect 19756 6656 19796 9388
rect 19948 8672 19988 10984
rect 20048 10604 20416 10613
rect 20088 10564 20130 10604
rect 20170 10564 20212 10604
rect 20252 10564 20294 10604
rect 20334 10564 20376 10604
rect 20048 10555 20416 10564
rect 20524 10436 20564 14008
rect 20524 10387 20564 10396
rect 20812 10184 20852 14008
rect 20908 13208 20948 17536
rect 21004 17240 21044 22576
rect 21100 17996 21140 23080
rect 21196 20180 21236 23920
rect 21292 22280 21332 27364
rect 21388 24716 21428 32992
rect 21388 24667 21428 24676
rect 21388 24548 21428 24557
rect 21484 24548 21524 33160
rect 21428 24508 21524 24548
rect 21388 24499 21428 24508
rect 21292 22231 21332 22240
rect 21388 22952 21428 22961
rect 21196 20131 21236 20140
rect 21292 22112 21332 22121
rect 21100 17947 21140 17956
rect 21196 20012 21236 20021
rect 21004 17191 21044 17200
rect 21196 16904 21236 19972
rect 21292 17156 21332 22072
rect 21292 17107 21332 17116
rect 21196 16855 21236 16864
rect 20908 13159 20948 13168
rect 21004 16568 21044 16577
rect 20812 10135 20852 10144
rect 20908 13040 20948 13049
rect 20044 9764 20084 9773
rect 20044 9680 20084 9724
rect 20044 9629 20084 9640
rect 20908 9512 20948 13000
rect 21004 12536 21044 16528
rect 21388 16232 21428 22912
rect 21484 21104 21524 21113
rect 21484 18248 21524 21064
rect 21484 18199 21524 18208
rect 21292 16192 21428 16232
rect 21004 12487 21044 12496
rect 21196 15560 21236 15569
rect 20908 9463 20948 9472
rect 21004 12032 21044 12041
rect 20048 9092 20416 9101
rect 20088 9052 20130 9092
rect 20170 9052 20212 9092
rect 20252 9052 20294 9092
rect 20334 9052 20376 9092
rect 20048 9043 20416 9052
rect 19948 8623 19988 8632
rect 21004 8672 21044 11992
rect 21196 11024 21236 15520
rect 21292 13460 21332 16192
rect 21292 13411 21332 13420
rect 21388 16064 21428 16073
rect 21388 11696 21428 16024
rect 21388 11647 21428 11656
rect 21196 10975 21236 10984
rect 21388 11024 21428 11033
rect 21004 8623 21044 8632
rect 21100 10016 21140 10025
rect 20908 8504 20948 8513
rect 20716 7916 20756 7925
rect 20048 7580 20416 7589
rect 20088 7540 20130 7580
rect 20170 7540 20212 7580
rect 20252 7540 20294 7580
rect 20334 7540 20376 7580
rect 20048 7531 20416 7540
rect 19756 6607 19796 6616
rect 20524 7496 20564 7505
rect 19564 5599 19604 5608
rect 19948 6404 19988 6413
rect 19948 4976 19988 6364
rect 20048 6068 20416 6077
rect 20088 6028 20130 6068
rect 20170 6028 20212 6068
rect 20252 6028 20294 6068
rect 20334 6028 20376 6068
rect 20048 6019 20416 6028
rect 19948 4927 19988 4936
rect 20428 4976 20468 4985
rect 20524 4976 20564 7456
rect 20716 5732 20756 7876
rect 20716 5683 20756 5692
rect 20908 5648 20948 8464
rect 21100 7160 21140 9976
rect 21100 7111 21140 7120
rect 21196 9512 21236 9521
rect 21196 6572 21236 9472
rect 21388 8000 21428 10984
rect 21388 7951 21428 7960
rect 21196 6523 21236 6532
rect 20908 5599 20948 5608
rect 20468 4936 20564 4976
rect 21292 5480 21332 5489
rect 20428 4927 20468 4936
rect 20048 4556 20416 4565
rect 20088 4516 20130 4556
rect 20170 4516 20212 4556
rect 20252 4516 20294 4556
rect 20334 4516 20376 4556
rect 20048 4507 20416 4516
rect 21292 4136 21332 5440
rect 21292 4087 21332 4096
rect 20332 3968 20372 3977
rect 20332 3464 20372 3928
rect 20332 3415 20372 3424
rect 20048 3044 20416 3053
rect 20088 3004 20130 3044
rect 20170 3004 20212 3044
rect 20252 3004 20294 3044
rect 20334 3004 20376 3044
rect 20048 2995 20416 3004
rect 19468 1987 19508 1996
rect 20048 1532 20416 1541
rect 20088 1492 20130 1532
rect 20170 1492 20212 1532
rect 20252 1492 20294 1532
rect 20334 1492 20376 1532
rect 20048 1483 20416 1492
rect 19276 1448 19316 1457
rect 18700 1324 18932 1364
rect 18508 1280 18548 1289
rect 18316 524 18356 533
rect 18316 80 18356 484
rect 18508 80 18548 1240
rect 18700 1196 18740 1205
rect 18700 80 18740 1156
rect 18892 80 18932 1324
rect 19084 188 19124 197
rect 19084 80 19124 148
rect 19276 80 19316 1408
rect 19468 1448 19508 1457
rect 19468 80 19508 1408
rect 1784 0 1864 80
rect 1976 0 2056 80
rect 2168 0 2248 80
rect 2360 0 2440 80
rect 2552 0 2632 80
rect 2744 0 2824 80
rect 2936 0 3016 80
rect 3128 0 3208 80
rect 3320 0 3400 80
rect 3512 0 3592 80
rect 3704 0 3784 80
rect 3896 0 3976 80
rect 4088 0 4168 80
rect 4280 0 4360 80
rect 4472 0 4552 80
rect 4664 0 4744 80
rect 4856 0 4936 80
rect 5048 0 5128 80
rect 5240 0 5320 80
rect 5432 0 5512 80
rect 5624 0 5704 80
rect 5816 0 5896 80
rect 6008 0 6088 80
rect 6200 0 6280 80
rect 6392 0 6472 80
rect 6584 0 6664 80
rect 6776 0 6856 80
rect 6968 0 7048 80
rect 7160 0 7240 80
rect 7352 0 7432 80
rect 7544 0 7624 80
rect 7736 0 7816 80
rect 7928 0 8008 80
rect 8120 0 8200 80
rect 8312 0 8392 80
rect 8504 0 8584 80
rect 8696 0 8776 80
rect 8888 0 8968 80
rect 9080 0 9160 80
rect 9272 0 9352 80
rect 9464 0 9544 80
rect 9656 0 9736 80
rect 9848 0 9928 80
rect 10040 0 10120 80
rect 10232 0 10312 80
rect 10424 0 10504 80
rect 10616 0 10696 80
rect 10808 0 10888 80
rect 11000 0 11080 80
rect 11192 0 11272 80
rect 11384 0 11464 80
rect 11576 0 11656 80
rect 11768 0 11848 80
rect 11960 0 12040 80
rect 12152 0 12232 80
rect 12344 0 12424 80
rect 12536 0 12616 80
rect 12728 0 12808 80
rect 12920 0 13000 80
rect 13112 0 13192 80
rect 13304 0 13384 80
rect 13496 0 13576 80
rect 13688 0 13768 80
rect 13880 0 13960 80
rect 14072 0 14152 80
rect 14264 0 14344 80
rect 14456 0 14536 80
rect 14648 0 14728 80
rect 14840 0 14920 80
rect 15032 0 15112 80
rect 15224 0 15304 80
rect 15416 0 15496 80
rect 15608 0 15688 80
rect 15800 0 15880 80
rect 15992 0 16072 80
rect 16184 0 16264 80
rect 16376 0 16456 80
rect 16568 0 16648 80
rect 16760 0 16840 80
rect 16952 0 17032 80
rect 17144 0 17224 80
rect 17336 0 17416 80
rect 17528 0 17608 80
rect 17720 0 17800 80
rect 17912 0 17992 80
rect 18104 0 18184 80
rect 18296 0 18376 80
rect 18488 0 18568 80
rect 18680 0 18760 80
rect 18872 0 18952 80
rect 19064 0 19144 80
rect 19256 0 19336 80
rect 19448 0 19528 80
<< via3 >>
rect 1324 94816 1364 94856
rect 1708 94816 1748 94856
rect 364 79528 404 79568
rect 748 86164 788 86204
rect 652 80872 692 80912
rect 364 73816 404 73856
rect 556 75496 596 75536
rect 556 74404 596 74444
rect 460 69112 500 69152
rect 1420 90280 1460 90320
rect 1132 87424 1172 87464
rect 1420 89860 1460 89900
rect 1420 89440 1460 89480
rect 1324 87424 1364 87464
rect 1228 86164 1268 86204
rect 940 80872 980 80912
rect 844 76756 884 76796
rect 748 70708 788 70748
rect 1132 76756 1172 76796
rect 1612 89692 1652 89732
rect 1612 89356 1652 89396
rect 1420 85492 1460 85532
rect 1420 82048 1460 82088
rect 1228 76504 1268 76544
rect 1132 75748 1172 75788
rect 1036 72472 1076 72512
rect 1228 70960 1268 71000
rect 1420 74320 1460 74360
rect 1420 74152 1460 74192
rect 1228 68944 1268 68984
rect 1324 68188 1364 68228
rect 1420 67600 1460 67640
rect 1420 66928 1460 66968
rect 1612 84064 1652 84104
rect 2092 94816 2132 94856
rect 2476 94816 2516 94856
rect 2572 93556 2612 93596
rect 1612 80368 1652 80408
rect 1708 83392 1748 83432
rect 1612 79276 1652 79316
rect 1612 76924 1652 76964
rect 1612 76756 1652 76796
rect 1996 89776 2036 89816
rect 1996 89608 2036 89648
rect 1900 84232 1940 84272
rect 1900 84064 1940 84104
rect 1900 82636 1940 82676
rect 1900 82300 1940 82340
rect 1804 80536 1844 80576
rect 1900 82132 1940 82172
rect 1804 79864 1844 79904
rect 1804 79444 1844 79484
rect 1708 72052 1748 72092
rect 1612 68356 1652 68396
rect 1516 63316 1556 63356
rect 1420 63232 1460 63272
rect 1804 68440 1844 68480
rect 1804 66256 1844 66296
rect 1708 64408 1748 64448
rect 1420 59368 1460 59408
rect 2188 86332 2228 86372
rect 2188 85744 2228 85784
rect 3148 93808 3188 93848
rect 2860 93556 2900 93596
rect 2956 92632 2996 92672
rect 2764 92296 2804 92336
rect 2476 89272 2516 89312
rect 2476 87928 2516 87968
rect 3052 90868 3092 90908
rect 2764 89944 2804 89984
rect 2860 89692 2900 89732
rect 2860 89440 2900 89480
rect 3052 89356 3092 89396
rect 2956 88852 2996 88892
rect 2764 87844 2804 87884
rect 2572 85744 2612 85784
rect 2476 82132 2516 82172
rect 2476 81880 2516 81920
rect 2380 80872 2420 80912
rect 2092 80452 2132 80492
rect 2188 80200 2228 80240
rect 1996 76924 2036 76964
rect 1996 74068 2036 74108
rect 1996 73420 2036 73460
rect 1996 73312 2036 73352
rect 2380 79108 2420 79148
rect 2284 76924 2324 76964
rect 2284 76756 2324 76796
rect 2476 77008 2516 77048
rect 2284 73564 2324 73604
rect 2380 73420 2420 73460
rect 2668 84988 2708 85028
rect 2956 87256 2996 87296
rect 2956 85072 2996 85112
rect 2668 83980 2708 84020
rect 2668 83392 2708 83432
rect 3628 94900 3668 94940
rect 4012 94816 4052 94856
rect 3688 94480 3728 94520
rect 3770 94480 3810 94520
rect 3852 94480 3892 94520
rect 3934 94480 3974 94520
rect 4016 94480 4056 94520
rect 4396 94816 4436 94856
rect 4588 95572 4628 95612
rect 5260 95572 5300 95612
rect 4928 95236 4968 95276
rect 5010 95236 5050 95276
rect 5092 95236 5132 95276
rect 5174 95236 5214 95276
rect 5256 95236 5296 95276
rect 5548 94816 5588 94856
rect 4972 94144 5012 94184
rect 4588 93892 4628 93932
rect 5356 94144 5396 94184
rect 5740 94144 5780 94184
rect 4928 93724 4968 93764
rect 5010 93724 5050 93764
rect 5092 93724 5132 93764
rect 5174 93724 5214 93764
rect 5256 93724 5296 93764
rect 3688 92968 3728 93008
rect 3770 92968 3810 93008
rect 3852 92968 3892 93008
rect 3934 92968 3974 93008
rect 4016 92968 4056 93008
rect 3688 91456 3728 91496
rect 3770 91456 3810 91496
rect 3852 91456 3892 91496
rect 3934 91456 3974 91496
rect 4016 91456 4056 91496
rect 3244 89608 3284 89648
rect 3244 89020 3284 89060
rect 3244 88852 3284 88892
rect 3340 87256 3380 87296
rect 3244 84988 3284 85028
rect 4012 90112 4052 90152
rect 3688 89944 3728 89984
rect 3770 89944 3810 89984
rect 3852 89944 3892 89984
rect 3934 89944 3974 89984
rect 4016 89944 4056 89984
rect 3628 89776 3668 89816
rect 3628 89356 3668 89396
rect 3688 88432 3728 88472
rect 3770 88432 3810 88472
rect 3852 88432 3892 88472
rect 3934 88432 3974 88472
rect 4016 88432 4056 88472
rect 3628 87256 3668 87296
rect 3244 83560 3284 83600
rect 2668 81292 2708 81332
rect 2668 81040 2708 81080
rect 2668 80536 2708 80576
rect 3148 83224 3188 83264
rect 4012 87088 4052 87128
rect 3688 86920 3728 86960
rect 3770 86920 3810 86960
rect 3852 86920 3892 86960
rect 3934 86920 3974 86960
rect 4016 86920 4056 86960
rect 4012 86752 4052 86792
rect 3688 85408 3728 85448
rect 3770 85408 3810 85448
rect 3852 85408 3892 85448
rect 3934 85408 3974 85448
rect 4016 85408 4056 85448
rect 3628 84904 3668 84944
rect 3724 84568 3764 84608
rect 3724 84316 3764 84356
rect 4012 84064 4052 84104
rect 3688 83896 3728 83936
rect 3770 83896 3810 83936
rect 3852 83896 3892 83936
rect 3934 83896 3974 83936
rect 4016 83896 4056 83936
rect 3532 82972 3572 83012
rect 3724 83644 3764 83684
rect 2860 80704 2900 80744
rect 2668 79948 2708 79988
rect 2956 80200 2996 80240
rect 2956 80032 2996 80072
rect 3244 82468 3284 82508
rect 3724 82552 3764 82592
rect 3916 82552 3956 82592
rect 4108 83560 4148 83600
rect 3688 82384 3728 82424
rect 3770 82384 3810 82424
rect 3852 82384 3892 82424
rect 3934 82384 3974 82424
rect 4016 82384 4056 82424
rect 4012 82048 4052 82088
rect 3820 81964 3860 82004
rect 2668 79108 2708 79148
rect 2860 77176 2900 77216
rect 3340 80032 3380 80072
rect 3244 79444 3284 79484
rect 3244 78940 3284 78980
rect 2860 76588 2900 76628
rect 2956 76336 2996 76376
rect 2860 76000 2900 76040
rect 2572 73060 2612 73100
rect 2188 71716 2228 71756
rect 2284 71296 2324 71336
rect 2284 68440 2324 68480
rect 2092 67432 2132 67472
rect 2188 68356 2228 68396
rect 1996 66844 2036 66884
rect 1996 66676 2036 66716
rect 1900 63484 1940 63524
rect 2092 64072 2132 64112
rect 1900 59284 1940 59324
rect 1804 57352 1844 57392
rect 1708 53992 1748 54032
rect 3148 77680 3188 77720
rect 3052 73648 3092 73688
rect 3148 76588 3188 76628
rect 2956 73480 2996 73520
rect 2956 72892 2996 72932
rect 2860 72472 2900 72512
rect 2956 72220 2996 72260
rect 2956 71716 2996 71756
rect 2860 71464 2900 71504
rect 2764 70036 2804 70076
rect 2668 69112 2708 69152
rect 2956 69868 2996 69908
rect 2764 69196 2804 69236
rect 2860 69112 2900 69152
rect 2476 68776 2516 68816
rect 2956 68104 2996 68144
rect 2668 66844 2708 66884
rect 2572 65752 2612 65792
rect 2860 65920 2900 65960
rect 2764 65752 2804 65792
rect 3052 65836 3092 65876
rect 2284 64072 2324 64112
rect 2380 63400 2420 63440
rect 2476 64156 2516 64196
rect 2188 61468 2228 61508
rect 1996 54748 2036 54788
rect 1804 51808 1844 51848
rect 2284 60040 2324 60080
rect 2860 65416 2900 65456
rect 2956 65332 2996 65372
rect 2860 64576 2900 64616
rect 2860 63736 2900 63776
rect 2668 61804 2708 61844
rect 2860 62812 2900 62852
rect 3052 64660 3092 64700
rect 4396 88936 4436 88976
rect 4396 85072 4436 85112
rect 4300 84148 4340 84188
rect 4396 83644 4436 83684
rect 4300 83476 4340 83516
rect 4396 83308 4436 83348
rect 4204 82888 4244 82928
rect 4300 83056 4340 83096
rect 4300 82720 4340 82760
rect 3628 81040 3668 81080
rect 4300 81292 4340 81332
rect 3688 80872 3728 80912
rect 3770 80872 3810 80912
rect 3852 80872 3892 80912
rect 3934 80872 3974 80912
rect 4016 80872 4056 80912
rect 3724 79696 3764 79736
rect 4012 80704 4052 80744
rect 4012 79612 4052 79652
rect 3628 79528 3668 79568
rect 3688 79360 3728 79400
rect 3770 79360 3810 79400
rect 3852 79360 3892 79400
rect 3934 79360 3974 79400
rect 4016 79360 4056 79400
rect 3532 78268 3572 78308
rect 3148 63484 3188 63524
rect 3244 73648 3284 73688
rect 3052 63232 3092 63272
rect 3148 63316 3188 63356
rect 2668 60964 2708 61004
rect 2476 60292 2516 60332
rect 2956 62140 2996 62180
rect 2668 57856 2708 57896
rect 2860 58444 2900 58484
rect 2668 57268 2708 57308
rect 3148 58360 3188 58400
rect 3148 58192 3188 58232
rect 2572 54832 2612 54872
rect 2668 54916 2708 54956
rect 2188 53488 2228 53528
rect 2860 54916 2900 54956
rect 2668 53152 2708 53192
rect 2860 53152 2900 53192
rect 2572 50968 2612 51008
rect 2380 50800 2420 50840
rect 3052 53404 3092 53444
rect 3052 53236 3092 53276
rect 2668 48028 2708 48068
rect 1996 47188 2036 47228
rect 76 38200 116 38240
rect 76 32656 116 32696
rect 1996 43072 2036 43112
rect 1516 40720 1556 40760
rect 1324 38452 1364 38492
rect 1420 36520 1460 36560
rect 1420 35008 1460 35048
rect 1996 41896 2036 41936
rect 1612 36520 1652 36560
rect 1612 35008 1652 35048
rect 1612 34588 1652 34628
rect 1516 33664 1556 33704
rect 460 28288 500 28328
rect 172 25600 212 25640
rect 76 25516 116 25556
rect 268 19384 308 19424
rect 460 20644 500 20684
rect 1036 29884 1076 29924
rect 1516 33076 1556 33116
rect 1420 32152 1460 32192
rect 1132 28792 1172 28832
rect 748 19384 788 19424
rect 1324 29800 1364 29840
rect 1324 28540 1364 28580
rect 1132 22408 1172 22448
rect 1228 13840 1268 13880
rect 1708 33496 1748 33536
rect 1900 39544 1940 39584
rect 1804 33412 1844 33452
rect 1708 30892 1748 30932
rect 1708 30220 1748 30260
rect 1612 28372 1652 28412
rect 1612 28120 1652 28160
rect 1612 25180 1652 25220
rect 1612 21568 1652 21608
rect 1420 13840 1460 13880
rect 1420 12832 1460 12872
rect 2188 43240 2228 43280
rect 2860 45508 2900 45548
rect 2284 41896 2324 41936
rect 2284 41224 2324 41264
rect 2188 40804 2228 40844
rect 2476 41728 2516 41768
rect 2380 40804 2420 40844
rect 2284 36772 2324 36812
rect 3052 45592 3092 45632
rect 4012 78268 4052 78308
rect 3724 78184 3764 78224
rect 4108 78184 4148 78224
rect 3688 77848 3728 77888
rect 3770 77848 3810 77888
rect 3852 77848 3892 77888
rect 3934 77848 3974 77888
rect 4016 77848 4056 77888
rect 3820 77428 3860 77468
rect 3628 76588 3668 76628
rect 3688 76336 3728 76376
rect 3770 76336 3810 76376
rect 3852 76336 3892 76376
rect 3934 76336 3974 76376
rect 4016 76336 4056 76376
rect 3628 75832 3668 75872
rect 3688 74824 3728 74864
rect 3770 74824 3810 74864
rect 3852 74824 3892 74864
rect 3934 74824 3974 74864
rect 4016 74824 4056 74864
rect 3532 74320 3572 74360
rect 3916 74152 3956 74192
rect 3532 73816 3572 73856
rect 3688 73312 3728 73352
rect 3770 73312 3810 73352
rect 3852 73312 3892 73352
rect 3934 73312 3974 73352
rect 4016 73312 4056 73352
rect 3340 72388 3380 72428
rect 3340 69196 3380 69236
rect 3436 70456 3476 70496
rect 3340 68104 3380 68144
rect 3436 68776 3476 68816
rect 3340 67600 3380 67640
rect 3340 66256 3380 66296
rect 3340 66088 3380 66128
rect 3340 65164 3380 65204
rect 3340 64744 3380 64784
rect 3628 72052 3668 72092
rect 3688 71800 3728 71840
rect 3770 71800 3810 71840
rect 3852 71800 3892 71840
rect 3934 71800 3974 71840
rect 4016 71800 4056 71840
rect 3628 71632 3668 71672
rect 4396 79864 4436 79904
rect 4396 78520 4436 78560
rect 4684 88936 4724 88976
rect 4928 92212 4968 92252
rect 5010 92212 5050 92252
rect 5092 92212 5132 92252
rect 5174 92212 5214 92252
rect 5256 92212 5296 92252
rect 6316 94816 6356 94856
rect 6700 94816 6740 94856
rect 7084 94816 7124 94856
rect 6124 94144 6164 94184
rect 4928 90700 4968 90740
rect 5010 90700 5050 90740
rect 5092 90700 5132 90740
rect 5174 90700 5214 90740
rect 5256 90700 5296 90740
rect 4928 89188 4968 89228
rect 5010 89188 5050 89228
rect 5092 89188 5132 89228
rect 5174 89188 5214 89228
rect 5256 89188 5296 89228
rect 4928 87676 4968 87716
rect 5010 87676 5050 87716
rect 5092 87676 5132 87716
rect 5174 87676 5214 87716
rect 5256 87676 5296 87716
rect 5164 86584 5204 86624
rect 4928 86164 4968 86204
rect 5010 86164 5050 86204
rect 5092 86164 5132 86204
rect 5174 86164 5214 86204
rect 5256 86164 5296 86204
rect 4684 84484 4724 84524
rect 4928 84652 4968 84692
rect 5010 84652 5050 84692
rect 5092 84652 5132 84692
rect 5174 84652 5214 84692
rect 5256 84652 5296 84692
rect 4780 83308 4820 83348
rect 5644 87256 5684 87296
rect 5740 87088 5780 87128
rect 5644 86752 5684 86792
rect 5356 83476 5396 83516
rect 5452 85072 5492 85112
rect 5548 84484 5588 84524
rect 5836 86668 5876 86708
rect 5740 84484 5780 84524
rect 4684 82888 4724 82928
rect 4684 80956 4724 80996
rect 4928 83140 4968 83180
rect 5010 83140 5050 83180
rect 5092 83140 5132 83180
rect 5174 83140 5214 83180
rect 5256 83140 5296 83180
rect 4972 82972 5012 83012
rect 4780 82048 4820 82088
rect 4396 73984 4436 74024
rect 4300 73900 4340 73940
rect 4300 73648 4340 73688
rect 4204 72304 4244 72344
rect 3724 70624 3764 70664
rect 3916 70624 3956 70664
rect 3628 70456 3668 70496
rect 3916 70456 3956 70496
rect 3688 70288 3728 70328
rect 3770 70288 3810 70328
rect 3852 70288 3892 70328
rect 3934 70288 3974 70328
rect 4016 70288 4056 70328
rect 3628 69196 3668 69236
rect 3688 68776 3728 68816
rect 3770 68776 3810 68816
rect 3852 68776 3892 68816
rect 3934 68776 3974 68816
rect 4016 68776 4056 68816
rect 4012 68440 4052 68480
rect 3916 68272 3956 68312
rect 4300 70624 4340 70664
rect 4876 82636 4916 82676
rect 4876 81964 4916 82004
rect 4972 81796 5012 81836
rect 4928 81628 4968 81668
rect 5010 81628 5050 81668
rect 5092 81628 5132 81668
rect 5174 81628 5214 81668
rect 5256 81628 5296 81668
rect 5164 81460 5204 81500
rect 4972 81208 5012 81248
rect 5356 81292 5396 81332
rect 5164 80284 5204 80324
rect 5548 83224 5588 83264
rect 4928 80116 4968 80156
rect 5010 80116 5050 80156
rect 5092 80116 5132 80156
rect 5174 80116 5214 80156
rect 5256 80116 5296 80156
rect 5260 79528 5300 79568
rect 4928 78604 4968 78644
rect 5010 78604 5050 78644
rect 5092 78604 5132 78644
rect 5174 78604 5214 78644
rect 5256 78604 5296 78644
rect 5356 77512 5396 77552
rect 5452 78940 5492 78980
rect 5260 77428 5300 77468
rect 4928 77092 4968 77132
rect 5010 77092 5050 77132
rect 5092 77092 5132 77132
rect 5174 77092 5214 77132
rect 5256 77092 5296 77132
rect 5452 76336 5492 76376
rect 5260 75916 5300 75956
rect 4684 75748 4724 75788
rect 4928 75580 4968 75620
rect 5010 75580 5050 75620
rect 5092 75580 5132 75620
rect 5174 75580 5214 75620
rect 5256 75580 5296 75620
rect 4876 75244 4916 75284
rect 4588 72136 4628 72176
rect 4108 67852 4148 67892
rect 4012 67432 4052 67472
rect 3688 67264 3728 67304
rect 3770 67264 3810 67304
rect 3852 67264 3892 67304
rect 3934 67264 3974 67304
rect 4016 67264 4056 67304
rect 3628 67012 3668 67052
rect 3628 66088 3668 66128
rect 3820 66760 3860 66800
rect 3820 66172 3860 66212
rect 3688 65752 3728 65792
rect 3770 65752 3810 65792
rect 3852 65752 3892 65792
rect 3934 65752 3974 65792
rect 4016 65752 4056 65792
rect 4012 65332 4052 65372
rect 3436 63400 3476 63440
rect 3436 63232 3476 63272
rect 3628 65164 3668 65204
rect 3820 64912 3860 64952
rect 3688 64240 3728 64280
rect 3770 64240 3810 64280
rect 3852 64240 3892 64280
rect 3934 64240 3974 64280
rect 4016 64240 4056 64280
rect 4012 63988 4052 64028
rect 3688 62728 3728 62768
rect 3770 62728 3810 62768
rect 3852 62728 3892 62768
rect 3934 62728 3974 62768
rect 4016 62728 4056 62768
rect 3532 61636 3572 61676
rect 4012 62308 4052 62348
rect 4012 61552 4052 61592
rect 3628 61384 3668 61424
rect 3688 61216 3728 61256
rect 3770 61216 3810 61256
rect 3852 61216 3892 61256
rect 3934 61216 3974 61256
rect 4016 61216 4056 61256
rect 3628 61048 3668 61088
rect 3820 61048 3860 61088
rect 3724 60964 3764 61004
rect 4012 60880 4052 60920
rect 3916 60712 3956 60752
rect 3916 60292 3956 60332
rect 3916 59956 3956 59996
rect 3436 59536 3476 59576
rect 3340 58360 3380 58400
rect 3244 51892 3284 51932
rect 3688 59704 3728 59744
rect 3770 59704 3810 59744
rect 3852 59704 3892 59744
rect 3934 59704 3974 59744
rect 4016 59704 4056 59744
rect 3628 59536 3668 59576
rect 3532 58444 3572 58484
rect 3532 58276 3572 58316
rect 3436 56848 3476 56888
rect 3688 58192 3728 58232
rect 3770 58192 3810 58232
rect 3852 58192 3892 58232
rect 3934 58192 3974 58232
rect 4016 58192 4056 58232
rect 4012 57772 4052 57812
rect 3628 57604 3668 57644
rect 3628 56848 3668 56888
rect 3688 56680 3728 56720
rect 3770 56680 3810 56720
rect 3852 56680 3892 56720
rect 3934 56680 3974 56720
rect 4016 56680 4056 56720
rect 3688 55168 3728 55208
rect 3770 55168 3810 55208
rect 3852 55168 3892 55208
rect 3934 55168 3974 55208
rect 4016 55168 4056 55208
rect 3820 54664 3860 54704
rect 3724 53824 3764 53864
rect 3688 53656 3728 53696
rect 3770 53656 3810 53696
rect 3852 53656 3892 53696
rect 3934 53656 3974 53696
rect 4016 53656 4056 53696
rect 3436 53404 3476 53444
rect 3532 53320 3572 53360
rect 4492 67684 4532 67724
rect 5260 74656 5300 74696
rect 5164 74320 5204 74360
rect 4928 74068 4968 74108
rect 5010 74068 5050 74108
rect 5092 74068 5132 74108
rect 5174 74068 5214 74108
rect 5256 74068 5296 74108
rect 4972 73648 5012 73688
rect 5260 72724 5300 72764
rect 4928 72556 4968 72596
rect 5010 72556 5050 72596
rect 5092 72556 5132 72596
rect 5174 72556 5214 72596
rect 5256 72556 5296 72596
rect 5068 71464 5108 71504
rect 5260 71464 5300 71504
rect 4928 71044 4968 71084
rect 5010 71044 5050 71084
rect 5092 71044 5132 71084
rect 5174 71044 5214 71084
rect 5256 71044 5296 71084
rect 4972 70876 5012 70916
rect 4876 70708 4916 70748
rect 5164 70876 5204 70916
rect 5164 69700 5204 69740
rect 4928 69532 4968 69572
rect 5010 69532 5050 69572
rect 5092 69532 5132 69572
rect 5174 69532 5214 69572
rect 5256 69532 5296 69572
rect 5260 69364 5300 69404
rect 4684 68776 4724 68816
rect 4300 64576 4340 64616
rect 4204 63904 4244 63944
rect 4204 62728 4244 62768
rect 4300 63568 4340 63608
rect 3688 52144 3728 52184
rect 3770 52144 3810 52184
rect 3852 52144 3892 52184
rect 3934 52144 3974 52184
rect 4016 52144 4056 52184
rect 3688 50632 3728 50672
rect 3770 50632 3810 50672
rect 3852 50632 3892 50672
rect 3934 50632 3974 50672
rect 4016 50632 4056 50672
rect 3688 49120 3728 49160
rect 3770 49120 3810 49160
rect 3852 49120 3892 49160
rect 3934 49120 3974 49160
rect 4016 49120 4056 49160
rect 4492 64912 4532 64952
rect 4396 63064 4436 63104
rect 4876 68776 4916 68816
rect 4928 68020 4968 68060
rect 5010 68020 5050 68060
rect 5092 68020 5132 68060
rect 5174 68020 5214 68060
rect 5256 68020 5296 68060
rect 4876 67684 4916 67724
rect 5356 67768 5396 67808
rect 4876 66928 4916 66968
rect 4928 66508 4968 66548
rect 5010 66508 5050 66548
rect 5092 66508 5132 66548
rect 5174 66508 5214 66548
rect 5256 66508 5296 66548
rect 5356 66508 5396 66548
rect 5164 65332 5204 65372
rect 4928 64996 4968 65036
rect 5010 64996 5050 65036
rect 5092 64996 5132 65036
rect 5174 64996 5214 65036
rect 5256 64996 5296 65036
rect 4876 64492 4916 64532
rect 4780 64072 4820 64112
rect 4684 63484 4724 63524
rect 4780 63652 4820 63692
rect 4588 61552 4628 61592
rect 4684 63148 4724 63188
rect 4588 61384 4628 61424
rect 4396 59116 4436 59156
rect 4492 54748 4532 54788
rect 4492 53992 4532 54032
rect 4928 63484 4968 63524
rect 5010 63484 5050 63524
rect 5092 63484 5132 63524
rect 5174 63484 5214 63524
rect 5256 63484 5296 63524
rect 5260 63316 5300 63356
rect 4780 62896 4820 62936
rect 4972 62812 5012 62852
rect 4876 62140 4916 62180
rect 5836 82720 5876 82760
rect 6028 87844 6068 87884
rect 6316 89776 6356 89816
rect 6220 87844 6260 87884
rect 5932 82216 5972 82256
rect 6124 81460 6164 81500
rect 6220 82216 6260 82256
rect 6028 81208 6068 81248
rect 5932 81124 5972 81164
rect 5836 78940 5876 78980
rect 5740 75160 5780 75200
rect 6028 80704 6068 80744
rect 6028 80368 6068 80408
rect 6028 80116 6068 80156
rect 6028 79612 6068 79652
rect 6028 79192 6068 79232
rect 6028 76252 6068 76292
rect 5932 76168 5972 76208
rect 5836 74488 5876 74528
rect 6412 86584 6452 86624
rect 6412 82216 6452 82256
rect 6508 81628 6548 81668
rect 6508 80956 6548 80996
rect 6508 80536 6548 80576
rect 6508 80200 6548 80240
rect 6220 76252 6260 76292
rect 6220 76084 6260 76124
rect 6220 75580 6260 75620
rect 5932 74404 5972 74444
rect 5836 73900 5876 73940
rect 5932 74068 5972 74108
rect 6220 74488 6260 74528
rect 7180 93556 7220 93596
rect 8044 94144 8084 94184
rect 7564 88600 7604 88640
rect 7276 86668 7316 86708
rect 6796 86248 6836 86288
rect 7084 86248 7124 86288
rect 6700 84232 6740 84272
rect 6988 84568 7028 84608
rect 7180 85996 7220 86036
rect 7084 84232 7124 84272
rect 6988 83476 7028 83516
rect 8044 91792 8084 91832
rect 7948 91120 7988 91160
rect 8044 88600 8084 88640
rect 7852 87256 7892 87296
rect 7948 86752 7988 86792
rect 7948 86500 7988 86540
rect 8236 93892 8276 93932
rect 8332 91120 8372 91160
rect 8140 86332 8180 86372
rect 7756 85072 7796 85112
rect 7372 84064 7412 84104
rect 7468 83812 7508 83852
rect 7948 84064 7988 84104
rect 6988 83224 7028 83264
rect 6604 78436 6644 78476
rect 6700 80536 6740 80576
rect 6892 81628 6932 81668
rect 7660 83308 7700 83348
rect 6892 81460 6932 81500
rect 6988 79696 7028 79736
rect 6796 78688 6836 78728
rect 6796 78436 6836 78476
rect 6700 77512 6740 77552
rect 6604 76756 6644 76796
rect 6316 74068 6356 74108
rect 5740 73060 5780 73100
rect 6412 73480 6452 73520
rect 5548 70876 5588 70916
rect 5548 70540 5588 70580
rect 5548 69280 5588 69320
rect 5452 63148 5492 63188
rect 5548 67768 5588 67808
rect 4928 61972 4968 62012
rect 5010 61972 5050 62012
rect 5092 61972 5132 62012
rect 5174 61972 5214 62012
rect 5256 61972 5296 62012
rect 4928 60460 4968 60500
rect 5010 60460 5050 60500
rect 5092 60460 5132 60500
rect 5174 60460 5214 60500
rect 5256 60460 5296 60500
rect 5932 72220 5972 72260
rect 5836 72136 5876 72176
rect 5740 69112 5780 69152
rect 6220 70540 6260 70580
rect 5836 66088 5876 66128
rect 5740 63904 5780 63944
rect 5644 63652 5684 63692
rect 5740 61804 5780 61844
rect 5452 61468 5492 61508
rect 4876 60292 4916 60332
rect 4876 59116 4916 59156
rect 5356 60208 5396 60248
rect 4928 58948 4968 58988
rect 5010 58948 5050 58988
rect 5092 58948 5132 58988
rect 5174 58948 5214 58988
rect 5256 58948 5296 58988
rect 4876 57772 4916 57812
rect 4928 57436 4968 57476
rect 5010 57436 5050 57476
rect 5092 57436 5132 57476
rect 5174 57436 5214 57476
rect 5256 57436 5296 57476
rect 5644 58780 5684 58820
rect 5932 60124 5972 60164
rect 6220 66844 6260 66884
rect 6124 65836 6164 65876
rect 6604 73564 6644 73604
rect 6604 72892 6644 72932
rect 6316 65332 6356 65372
rect 6412 64744 6452 64784
rect 6316 64660 6356 64700
rect 6220 63652 6260 63692
rect 4928 55924 4968 55964
rect 5010 55924 5050 55964
rect 5092 55924 5132 55964
rect 5174 55924 5214 55964
rect 5256 55924 5296 55964
rect 5548 56932 5588 56972
rect 4928 54412 4968 54452
rect 5010 54412 5050 54452
rect 5092 54412 5132 54452
rect 5174 54412 5214 54452
rect 5256 54412 5296 54452
rect 4928 52900 4968 52940
rect 5010 52900 5050 52940
rect 5092 52900 5132 52940
rect 5174 52900 5214 52940
rect 5256 52900 5296 52940
rect 6316 62308 6356 62348
rect 6412 57772 6452 57812
rect 4928 51388 4968 51428
rect 5010 51388 5050 51428
rect 5092 51388 5132 51428
rect 5174 51388 5214 51428
rect 5256 51388 5296 51428
rect 4928 49876 4968 49916
rect 5010 49876 5050 49916
rect 5092 49876 5132 49916
rect 5174 49876 5214 49916
rect 5256 49876 5296 49916
rect 4204 48532 4244 48572
rect 3688 47608 3728 47648
rect 3770 47608 3810 47648
rect 3852 47608 3892 47648
rect 3934 47608 3974 47648
rect 4016 47608 4056 47648
rect 3340 46684 3380 46724
rect 3244 46600 3284 46640
rect 3916 47188 3956 47228
rect 3052 41308 3092 41348
rect 2860 38032 2900 38072
rect 2092 34252 2132 34292
rect 1900 29800 1940 29840
rect 2092 33160 2132 33200
rect 2092 33076 2132 33116
rect 2092 29296 2132 29336
rect 2092 29128 2132 29168
rect 1804 26776 1844 26816
rect 2188 26356 2228 26396
rect 1996 23920 2036 23960
rect 2092 25096 2132 25136
rect 1804 20896 1844 20936
rect 1900 21400 1940 21440
rect 1996 19972 2036 20012
rect 1900 14260 1940 14300
rect 1900 12940 1940 12980
rect 1708 9640 1748 9680
rect 1612 6112 1652 6152
rect 1804 8548 1844 8588
rect 2188 17956 2228 17996
rect 2188 15016 2228 15056
rect 2668 34672 2708 34712
rect 2764 34504 2804 34544
rect 2572 33664 2612 33704
rect 2476 33580 2516 33620
rect 2380 29716 2420 29756
rect 3148 40720 3188 40760
rect 3688 46096 3728 46136
rect 3770 46096 3810 46136
rect 3852 46096 3892 46136
rect 3934 46096 3974 46136
rect 4016 46096 4056 46136
rect 3916 45844 3956 45884
rect 4012 45760 4052 45800
rect 4108 45676 4148 45716
rect 3688 44584 3728 44624
rect 3770 44584 3810 44624
rect 3852 44584 3892 44624
rect 3934 44584 3974 44624
rect 4016 44584 4056 44624
rect 4012 44416 4052 44456
rect 3244 38284 3284 38324
rect 3052 38032 3092 38072
rect 2956 35176 2996 35216
rect 2956 35008 2996 35048
rect 2956 34504 2996 34544
rect 2860 33748 2900 33788
rect 3052 33664 3092 33704
rect 3916 43912 3956 43952
rect 3628 43492 3668 43532
rect 4012 43240 4052 43280
rect 3688 43072 3728 43112
rect 3770 43072 3810 43112
rect 3852 43072 3892 43112
rect 3934 43072 3974 43112
rect 4016 43072 4056 43112
rect 3688 41560 3728 41600
rect 3770 41560 3810 41600
rect 3852 41560 3892 41600
rect 3934 41560 3974 41600
rect 4016 41560 4056 41600
rect 3532 40720 3572 40760
rect 4108 40888 4148 40928
rect 3628 40216 3668 40256
rect 3688 40048 3728 40088
rect 3770 40048 3810 40088
rect 3852 40048 3892 40088
rect 3934 40048 3974 40088
rect 4016 40048 4056 40088
rect 4492 45592 4532 45632
rect 4492 45340 4532 45380
rect 4492 44080 4532 44120
rect 4928 48364 4968 48404
rect 5010 48364 5050 48404
rect 5092 48364 5132 48404
rect 5174 48364 5214 48404
rect 5256 48364 5296 48404
rect 4876 47944 4916 47984
rect 5356 47944 5396 47984
rect 4928 46852 4968 46892
rect 5010 46852 5050 46892
rect 5092 46852 5132 46892
rect 5174 46852 5214 46892
rect 5256 46852 5296 46892
rect 4684 46684 4724 46724
rect 5164 46684 5204 46724
rect 4780 45928 4820 45968
rect 4684 45676 4724 45716
rect 5068 46012 5108 46052
rect 6028 54244 6068 54284
rect 6412 56344 6452 56384
rect 6220 55336 6260 55376
rect 6220 54244 6260 54284
rect 6124 53908 6164 53948
rect 6124 53740 6164 53780
rect 5452 46684 5492 46724
rect 4588 43660 4628 43700
rect 4396 43072 4436 43112
rect 4928 45340 4968 45380
rect 5010 45340 5050 45380
rect 5092 45340 5132 45380
rect 5174 45340 5214 45380
rect 5256 45340 5296 45380
rect 5452 45844 5492 45884
rect 5452 45172 5492 45212
rect 5068 44332 5108 44372
rect 4876 43996 4916 44036
rect 5260 44584 5300 44624
rect 5452 44500 5492 44540
rect 5260 44248 5300 44288
rect 4928 43828 4968 43868
rect 5010 43828 5050 43868
rect 5092 43828 5132 43868
rect 5174 43828 5214 43868
rect 5256 43828 5296 43868
rect 5452 44080 5492 44120
rect 5452 43828 5492 43868
rect 5260 43660 5300 43700
rect 5356 43576 5396 43616
rect 4876 43240 4916 43280
rect 4588 42820 4628 42860
rect 4684 42652 4724 42692
rect 5164 42820 5204 42860
rect 4588 41560 4628 41600
rect 4588 41392 4628 41432
rect 4928 42316 4968 42356
rect 5010 42316 5050 42356
rect 5092 42316 5132 42356
rect 5174 42316 5214 42356
rect 5256 42316 5296 42356
rect 4492 39712 4532 39752
rect 4300 39292 4340 39332
rect 4396 39544 4436 39584
rect 3724 39208 3764 39248
rect 4300 38956 4340 38996
rect 4108 38872 4148 38912
rect 3688 38536 3728 38576
rect 3770 38536 3810 38576
rect 3852 38536 3892 38576
rect 3934 38536 3974 38576
rect 4016 38536 4056 38576
rect 3148 33496 3188 33536
rect 3532 38284 3572 38324
rect 2956 31900 2996 31940
rect 2668 30472 2708 30512
rect 2572 29800 2612 29840
rect 2860 29044 2900 29084
rect 2860 28792 2900 28832
rect 3052 30724 3092 30764
rect 3148 28456 3188 28496
rect 2476 25180 2516 25220
rect 2380 23248 2420 23288
rect 2380 22996 2420 23036
rect 2380 22156 2420 22196
rect 2380 21316 2420 21356
rect 2380 20812 2420 20852
rect 2380 16360 2420 16400
rect 2092 10480 2132 10520
rect 2092 10312 2132 10352
rect 2860 24844 2900 24884
rect 2956 25432 2996 25472
rect 2860 24340 2900 24380
rect 3052 24760 3092 24800
rect 3148 24676 3188 24716
rect 3820 37696 3860 37736
rect 3688 37024 3728 37064
rect 3770 37024 3810 37064
rect 3852 37024 3892 37064
rect 3934 37024 3974 37064
rect 4016 37024 4056 37064
rect 3628 36688 3668 36728
rect 3436 36520 3476 36560
rect 3340 34336 3380 34376
rect 3340 33328 3380 33368
rect 3724 35848 3764 35888
rect 4012 36100 4052 36140
rect 4108 35848 4148 35888
rect 3688 35512 3728 35552
rect 3770 35512 3810 35552
rect 3852 35512 3892 35552
rect 3934 35512 3974 35552
rect 4016 35512 4056 35552
rect 4012 34168 4052 34208
rect 3688 34000 3728 34040
rect 3770 34000 3810 34040
rect 3852 34000 3892 34040
rect 3934 34000 3974 34040
rect 4016 34000 4056 34040
rect 4300 38368 4340 38408
rect 4300 38200 4340 38240
rect 4492 39460 4532 39500
rect 4684 40972 4724 41012
rect 5164 41056 5204 41096
rect 5356 41812 5396 41852
rect 5356 41308 5396 41348
rect 4928 40804 4968 40844
rect 5010 40804 5050 40844
rect 5092 40804 5132 40844
rect 5174 40804 5214 40844
rect 5256 40804 5296 40844
rect 4876 40048 4916 40088
rect 4684 39124 4724 39164
rect 5068 40636 5108 40676
rect 5164 40468 5204 40508
rect 5260 40384 5300 40424
rect 5164 39796 5204 39836
rect 5068 39628 5108 39668
rect 4972 39544 5012 39584
rect 5164 39460 5204 39500
rect 4928 39292 4968 39332
rect 5010 39292 5050 39332
rect 5092 39292 5132 39332
rect 5174 39292 5214 39332
rect 5256 39292 5296 39332
rect 5356 39292 5396 39332
rect 4684 37444 4724 37484
rect 4928 37780 4968 37820
rect 5010 37780 5050 37820
rect 5092 37780 5132 37820
rect 5174 37780 5214 37820
rect 5256 37780 5296 37820
rect 4684 37276 4724 37316
rect 4396 35260 4436 35300
rect 3340 32068 3380 32108
rect 4204 35176 4244 35216
rect 3340 31732 3380 31772
rect 3340 23668 3380 23708
rect 3724 33664 3764 33704
rect 3820 33580 3860 33620
rect 4204 33580 4244 33620
rect 3916 32992 3956 33032
rect 3688 32488 3728 32528
rect 3770 32488 3810 32528
rect 3852 32488 3892 32528
rect 3934 32488 3974 32528
rect 4016 32488 4056 32528
rect 3532 32404 3572 32444
rect 3688 30976 3728 31016
rect 3770 30976 3810 31016
rect 3852 30976 3892 31016
rect 3934 30976 3974 31016
rect 4016 30976 4056 31016
rect 3916 30556 3956 30596
rect 4012 29632 4052 29672
rect 3688 29464 3728 29504
rect 3770 29464 3810 29504
rect 3852 29464 3892 29504
rect 3934 29464 3974 29504
rect 4016 29464 4056 29504
rect 4012 28792 4052 28832
rect 4012 28624 4052 28664
rect 3688 27952 3728 27992
rect 3770 27952 3810 27992
rect 3852 27952 3892 27992
rect 3934 27952 3974 27992
rect 4016 27952 4056 27992
rect 4012 27364 4052 27404
rect 3820 26860 3860 26900
rect 3688 26440 3728 26480
rect 3770 26440 3810 26480
rect 3852 26440 3892 26480
rect 3934 26440 3974 26480
rect 4016 26440 4056 26480
rect 3916 26272 3956 26312
rect 3436 23248 3476 23288
rect 3052 23020 3092 23060
rect 2668 18628 2708 18668
rect 2668 17956 2708 17996
rect 2860 20560 2900 20600
rect 2860 19384 2900 19424
rect 3052 19384 3092 19424
rect 2956 17788 2996 17828
rect 2668 14008 2708 14048
rect 2380 11656 2420 11696
rect 2284 10312 2324 10352
rect 2284 10144 2324 10184
rect 2188 10060 2228 10100
rect 1420 2920 1460 2960
rect 2476 10480 2516 10520
rect 3436 23080 3476 23120
rect 3628 25600 3668 25640
rect 3820 25600 3860 25640
rect 4012 25684 4052 25724
rect 3916 25432 3956 25472
rect 3688 24928 3728 24968
rect 3770 24928 3810 24968
rect 3852 24928 3892 24968
rect 3934 24928 3974 24968
rect 4016 24928 4056 24968
rect 3628 24760 3668 24800
rect 3916 24004 3956 24044
rect 3628 23752 3668 23792
rect 3724 23584 3764 23624
rect 4204 32992 4244 33032
rect 4492 33160 4532 33200
rect 4588 35848 4628 35888
rect 4396 32908 4436 32948
rect 4204 31060 4244 31100
rect 4300 29716 4340 29756
rect 4588 32824 4628 32864
rect 4492 30976 4532 31016
rect 4492 30640 4532 30680
rect 4492 28372 4532 28412
rect 4588 28120 4628 28160
rect 4204 25684 4244 25724
rect 4928 36268 4968 36308
rect 5010 36268 5050 36308
rect 5092 36268 5132 36308
rect 5174 36268 5214 36308
rect 5256 36268 5296 36308
rect 5644 48700 5684 48740
rect 6316 53908 6356 53948
rect 6124 48868 6164 48908
rect 5644 45928 5684 45968
rect 5548 43324 5588 43364
rect 5644 44500 5684 44540
rect 5548 43072 5588 43112
rect 6892 77428 6932 77468
rect 6892 76504 6932 76544
rect 6988 75916 7028 75956
rect 6796 73480 6836 73520
rect 6604 70876 6644 70916
rect 6700 71968 6740 72008
rect 6988 75076 7028 75116
rect 7660 81208 7700 81248
rect 7372 80200 7412 80240
rect 7276 79948 7316 79988
rect 7468 79696 7508 79736
rect 7372 78520 7412 78560
rect 7180 77512 7220 77552
rect 7276 77848 7316 77888
rect 7084 74572 7124 74612
rect 6988 73984 7028 74024
rect 6892 72052 6932 72092
rect 7084 73564 7124 73604
rect 7180 73396 7220 73436
rect 6604 66676 6644 66716
rect 6604 65920 6644 65960
rect 6700 63484 6740 63524
rect 6700 63316 6740 63356
rect 6700 61804 6740 61844
rect 6700 61468 6740 61508
rect 6700 53740 6740 53780
rect 6508 52564 6548 52604
rect 6988 69280 7028 69320
rect 8140 84148 8180 84188
rect 7948 78184 7988 78224
rect 8140 81292 8180 81332
rect 8812 94648 8852 94688
rect 9388 94648 9428 94688
rect 9772 94648 9812 94688
rect 10732 94732 10772 94772
rect 10540 94648 10580 94688
rect 11212 94648 11252 94688
rect 8428 85912 8468 85952
rect 8716 87508 8756 87548
rect 8620 85828 8660 85868
rect 8332 84148 8372 84188
rect 8332 83812 8372 83852
rect 8524 84904 8564 84944
rect 8524 83224 8564 83264
rect 8236 80116 8276 80156
rect 8332 80452 8372 80492
rect 7948 76084 7988 76124
rect 7660 74656 7700 74696
rect 7660 74236 7700 74276
rect 7948 75328 7988 75368
rect 8332 77344 8372 77384
rect 7948 74992 7988 75032
rect 8524 77428 8564 77468
rect 8428 76672 8468 76712
rect 8812 85996 8852 86036
rect 8716 83896 8756 83936
rect 8812 82216 8852 82256
rect 8908 84148 8948 84188
rect 8908 82552 8948 82592
rect 8716 81544 8756 81584
rect 8812 81964 8852 82004
rect 8716 81376 8756 81416
rect 8428 75328 8468 75368
rect 8236 75244 8276 75284
rect 7948 74572 7988 74612
rect 7276 72724 7316 72764
rect 7372 71464 7412 71504
rect 7276 71296 7316 71336
rect 7180 70792 7220 70832
rect 7372 70708 7412 70748
rect 7372 70540 7412 70580
rect 7660 70876 7700 70916
rect 7564 70708 7604 70748
rect 7660 70204 7700 70244
rect 7564 69364 7604 69404
rect 7180 68440 7220 68480
rect 7276 68524 7316 68564
rect 6988 67432 7028 67472
rect 6892 66424 6932 66464
rect 6892 66172 6932 66212
rect 7468 68440 7508 68480
rect 7372 66592 7412 66632
rect 7276 66172 7316 66212
rect 6988 63064 7028 63104
rect 7084 62812 7124 62852
rect 7084 61636 7124 61676
rect 7180 62476 7220 62516
rect 7084 61468 7124 61508
rect 7372 62476 7412 62516
rect 7372 61636 7412 61676
rect 7372 60880 7412 60920
rect 6988 53260 7028 53300
rect 6892 52396 6932 52436
rect 5932 45676 5972 45716
rect 6124 45676 6164 45716
rect 5932 44248 5972 44288
rect 5836 43828 5876 43868
rect 5740 43324 5780 43364
rect 5644 40468 5684 40508
rect 5644 40216 5684 40256
rect 5644 39292 5684 39332
rect 5836 42820 5876 42860
rect 6796 45676 6836 45716
rect 6700 45592 6740 45632
rect 6604 45424 6644 45464
rect 6124 43324 6164 43364
rect 6220 44584 6260 44624
rect 6412 44668 6452 44708
rect 6412 44500 6452 44540
rect 6508 44332 6548 44372
rect 6508 43576 6548 43616
rect 6412 43408 6452 43448
rect 6316 42904 6356 42944
rect 6124 41308 6164 41348
rect 6028 41140 6068 41180
rect 6124 41056 6164 41096
rect 6028 40720 6068 40760
rect 6028 40468 6068 40508
rect 6316 41056 6356 41096
rect 6124 39964 6164 40004
rect 5452 38452 5492 38492
rect 5452 36940 5492 36980
rect 5356 35848 5396 35888
rect 4780 35680 4820 35720
rect 5356 35680 5396 35720
rect 4780 35260 4820 35300
rect 4928 34756 4968 34796
rect 5010 34756 5050 34796
rect 5092 34756 5132 34796
rect 5174 34756 5214 34796
rect 5256 34756 5296 34796
rect 4972 34588 5012 34628
rect 4876 34420 4916 34460
rect 5260 34588 5300 34628
rect 4928 33244 4968 33284
rect 5010 33244 5050 33284
rect 5092 33244 5132 33284
rect 5174 33244 5214 33284
rect 5256 33244 5296 33284
rect 5260 32824 5300 32864
rect 5260 31900 5300 31940
rect 4928 31732 4968 31772
rect 5010 31732 5050 31772
rect 5092 31732 5132 31772
rect 5174 31732 5214 31772
rect 5256 31732 5296 31772
rect 5164 31564 5204 31604
rect 4876 30976 4916 31016
rect 5260 31480 5300 31520
rect 5164 30808 5204 30848
rect 5068 30556 5108 30596
rect 4928 30220 4968 30260
rect 5010 30220 5050 30260
rect 5092 30220 5132 30260
rect 5174 30220 5214 30260
rect 5256 30220 5296 30260
rect 5260 29968 5300 30008
rect 4876 28876 4916 28916
rect 5260 28876 5300 28916
rect 4928 28708 4968 28748
rect 5010 28708 5050 28748
rect 5092 28708 5132 28748
rect 5174 28708 5214 28748
rect 5256 28708 5296 28748
rect 4780 28624 4820 28664
rect 4780 28372 4820 28412
rect 5068 28540 5108 28580
rect 5260 28540 5300 28580
rect 4588 27112 4628 27152
rect 4492 26104 4532 26144
rect 4588 26020 4628 26060
rect 3688 23416 3728 23456
rect 3770 23416 3810 23456
rect 3852 23416 3892 23456
rect 3934 23416 3974 23456
rect 4016 23416 4056 23456
rect 3436 22324 3476 22364
rect 3532 22240 3572 22280
rect 3820 23248 3860 23288
rect 3436 22072 3476 22112
rect 3724 23164 3764 23204
rect 4012 23248 4052 23288
rect 3916 23080 3956 23120
rect 3916 22156 3956 22196
rect 4204 23248 4244 23288
rect 4396 23500 4436 23540
rect 3724 22072 3764 22112
rect 3688 21904 3728 21944
rect 3770 21904 3810 21944
rect 3852 21904 3892 21944
rect 3934 21904 3974 21944
rect 4016 21904 4056 21944
rect 3820 21736 3860 21776
rect 3436 19888 3476 19928
rect 4012 21568 4052 21608
rect 3916 20728 3956 20768
rect 3628 20644 3668 20684
rect 3688 20392 3728 20432
rect 3770 20392 3810 20432
rect 3852 20392 3892 20432
rect 3934 20392 3974 20432
rect 4016 20392 4056 20432
rect 3532 20224 3572 20264
rect 3244 18544 3284 18584
rect 3628 19888 3668 19928
rect 3532 19300 3572 19340
rect 3628 19216 3668 19256
rect 3688 18880 3728 18920
rect 3770 18880 3810 18920
rect 3852 18880 3892 18920
rect 3934 18880 3974 18920
rect 4016 18880 4056 18920
rect 3244 18292 3284 18332
rect 3148 15436 3188 15476
rect 2956 15352 2996 15392
rect 2860 13924 2900 13964
rect 2764 13504 2804 13544
rect 2860 11572 2900 11612
rect 3148 13504 3188 13544
rect 3628 18376 3668 18416
rect 3340 17452 3380 17492
rect 3916 17788 3956 17828
rect 4012 17704 4052 17744
rect 3436 17116 3476 17156
rect 3340 16444 3380 16484
rect 3052 13000 3092 13040
rect 3052 12328 3092 12368
rect 2092 2584 2132 2624
rect 2860 10480 2900 10520
rect 2956 9976 2996 10016
rect 2956 8464 2996 8504
rect 2860 6868 2900 6908
rect 2860 6280 2900 6320
rect 2380 3424 2420 3464
rect 3340 13336 3380 13376
rect 3688 17368 3728 17408
rect 3770 17368 3810 17408
rect 3852 17368 3892 17408
rect 3934 17368 3974 17408
rect 4016 17368 4056 17408
rect 3820 17116 3860 17156
rect 4396 21736 4436 21776
rect 4300 21400 4340 21440
rect 4300 18880 4340 18920
rect 4684 25852 4724 25892
rect 4588 24508 4628 24548
rect 4684 23584 4724 23624
rect 4588 21400 4628 21440
rect 4588 20728 4628 20768
rect 4204 18292 4244 18332
rect 4300 16948 4340 16988
rect 3688 15856 3728 15896
rect 3770 15856 3810 15896
rect 3852 15856 3892 15896
rect 3934 15856 3974 15896
rect 4016 15856 4056 15896
rect 3628 15604 3668 15644
rect 3688 14344 3728 14384
rect 3770 14344 3810 14384
rect 3852 14344 3892 14384
rect 3934 14344 3974 14384
rect 4016 14344 4056 14384
rect 3628 13924 3668 13964
rect 3340 13168 3380 13208
rect 3340 12832 3380 12872
rect 4012 13000 4052 13040
rect 3688 12832 3728 12872
rect 3770 12832 3810 12872
rect 3852 12832 3892 12872
rect 3934 12832 3974 12872
rect 4016 12832 4056 12872
rect 3916 12664 3956 12704
rect 3532 12580 3572 12620
rect 3724 12580 3764 12620
rect 3340 12496 3380 12536
rect 3244 12412 3284 12452
rect 3436 11152 3476 11192
rect 3436 10228 3476 10268
rect 3148 5524 3188 5564
rect 4928 27196 4968 27236
rect 5010 27196 5050 27236
rect 5092 27196 5132 27236
rect 5174 27196 5214 27236
rect 5256 27196 5296 27236
rect 5452 34000 5492 34040
rect 7180 54664 7220 54704
rect 7468 60460 7508 60500
rect 7084 52816 7124 52856
rect 7180 53152 7220 53192
rect 6988 51640 7028 51680
rect 7852 71464 7892 71504
rect 7852 68524 7892 68564
rect 8236 74152 8276 74192
rect 8140 72976 8180 73016
rect 8332 72892 8372 72932
rect 8428 73312 8468 73352
rect 8332 72724 8372 72764
rect 7756 63652 7796 63692
rect 8236 69280 8276 69320
rect 8236 68188 8276 68228
rect 8044 63904 8084 63944
rect 7948 63400 7988 63440
rect 8620 75244 8660 75284
rect 8908 81880 8948 81920
rect 8908 81124 8948 81164
rect 8812 80116 8852 80156
rect 8812 79528 8852 79568
rect 8908 74740 8948 74780
rect 8620 72892 8660 72932
rect 8812 72976 8852 73016
rect 8620 69448 8660 69488
rect 8716 68440 8756 68480
rect 8524 66592 8564 66632
rect 9196 83896 9236 83936
rect 9292 83728 9332 83768
rect 9196 83644 9236 83684
rect 9100 81544 9140 81584
rect 9100 78940 9140 78980
rect 9100 78268 9140 78308
rect 9100 78016 9140 78056
rect 9292 80536 9332 80576
rect 9292 80200 9332 80240
rect 9100 73480 9140 73520
rect 9964 93976 10004 94016
rect 11020 93976 11060 94016
rect 10156 93892 10196 93932
rect 10828 93892 10868 93932
rect 9676 83728 9716 83768
rect 9772 89356 9812 89396
rect 9772 81460 9812 81500
rect 9484 81124 9524 81164
rect 9484 78940 9524 78980
rect 9484 78688 9524 78728
rect 9292 73648 9332 73688
rect 9484 73816 9524 73856
rect 8908 70540 8948 70580
rect 8908 67096 8948 67136
rect 8620 64996 8660 65036
rect 8428 63904 8468 63944
rect 8140 63400 8180 63440
rect 8332 63232 8372 63272
rect 8236 63148 8276 63188
rect 7948 60124 7988 60164
rect 8044 60544 8084 60584
rect 8332 60712 8372 60752
rect 8620 63232 8660 63272
rect 8620 63064 8660 63104
rect 8524 62392 8564 62432
rect 8812 65164 8852 65204
rect 8812 64660 8852 64700
rect 8908 63988 8948 64028
rect 8908 63340 8948 63380
rect 9292 72052 9332 72092
rect 9292 69364 9332 69404
rect 9292 65584 9332 65624
rect 9292 64912 9332 64952
rect 9196 64072 9236 64112
rect 9484 71800 9524 71840
rect 9484 68608 9524 68648
rect 7564 48616 7604 48656
rect 6892 45340 6932 45380
rect 7948 54244 7988 54284
rect 7756 53908 7796 53948
rect 8140 56092 8180 56132
rect 8236 53908 8276 53948
rect 8428 51640 8468 51680
rect 6796 44080 6836 44120
rect 6796 43912 6836 43952
rect 6796 43660 6836 43700
rect 6700 43324 6740 43364
rect 6220 39460 6260 39500
rect 6028 39376 6068 39416
rect 5932 39040 5972 39080
rect 5836 38032 5876 38072
rect 5644 34000 5684 34040
rect 5548 32992 5588 33032
rect 5548 32488 5588 32528
rect 4928 25684 4968 25724
rect 5010 25684 5050 25724
rect 5092 25684 5132 25724
rect 5174 25684 5214 25724
rect 5256 25684 5296 25724
rect 4972 25516 5012 25556
rect 4876 25348 4916 25388
rect 5260 25012 5300 25052
rect 5932 34840 5972 34880
rect 5740 32320 5780 32360
rect 5836 31900 5876 31940
rect 5644 31396 5684 31436
rect 5548 30640 5588 30680
rect 4876 24424 4916 24464
rect 4928 24172 4968 24212
rect 5010 24172 5050 24212
rect 5092 24172 5132 24212
rect 5174 24172 5214 24212
rect 5256 24172 5296 24212
rect 4972 23920 5012 23960
rect 4780 22996 4820 23036
rect 4928 22660 4968 22700
rect 5010 22660 5050 22700
rect 5092 22660 5132 22700
rect 5174 22660 5214 22700
rect 5256 22660 5296 22700
rect 5548 28792 5588 28832
rect 5740 29968 5780 30008
rect 5836 28120 5876 28160
rect 5548 22828 5588 22868
rect 5644 25768 5684 25808
rect 4928 21148 4968 21188
rect 5010 21148 5050 21188
rect 5092 21148 5132 21188
rect 5174 21148 5214 21188
rect 5256 21148 5296 21188
rect 4780 20980 4820 21020
rect 5260 20896 5300 20936
rect 5164 20812 5204 20852
rect 5356 20812 5396 20852
rect 5164 20308 5204 20348
rect 4928 19636 4968 19676
rect 5010 19636 5050 19676
rect 5092 19636 5132 19676
rect 5174 19636 5214 19676
rect 5256 19636 5296 19676
rect 5548 20224 5588 20264
rect 5356 19636 5396 19676
rect 5452 19552 5492 19592
rect 4780 19384 4820 19424
rect 5164 19468 5204 19508
rect 5068 18544 5108 18584
rect 4972 18376 5012 18416
rect 4928 18124 4968 18164
rect 5010 18124 5050 18164
rect 5092 18124 5132 18164
rect 5174 18124 5214 18164
rect 5256 18124 5296 18164
rect 4492 15184 4532 15224
rect 4396 13840 4436 13880
rect 4684 14764 4724 14804
rect 3688 11320 3728 11360
rect 3770 11320 3810 11360
rect 3852 11320 3892 11360
rect 3934 11320 3974 11360
rect 4016 11320 4056 11360
rect 3724 11152 3764 11192
rect 3628 10312 3668 10352
rect 3724 9976 3764 10016
rect 3688 9808 3728 9848
rect 3770 9808 3810 9848
rect 3852 9808 3892 9848
rect 3934 9808 3974 9848
rect 4016 9808 4056 9848
rect 4012 9472 4052 9512
rect 3436 7960 3476 8000
rect 3916 8968 3956 9008
rect 3820 8632 3860 8672
rect 4588 13672 4628 13712
rect 4684 11824 4724 11864
rect 4300 10732 4340 10772
rect 3916 8548 3956 8588
rect 3688 8296 3728 8336
rect 3770 8296 3810 8336
rect 3852 8296 3892 8336
rect 3934 8296 3974 8336
rect 4016 8296 4056 8336
rect 3688 6784 3728 6824
rect 3770 6784 3810 6824
rect 3852 6784 3892 6824
rect 3934 6784 3974 6824
rect 4016 6784 4056 6824
rect 4300 8128 4340 8168
rect 4684 10228 4724 10268
rect 4588 8128 4628 8168
rect 4108 5692 4148 5732
rect 3688 5272 3728 5312
rect 3770 5272 3810 5312
rect 3852 5272 3892 5312
rect 3934 5272 3974 5312
rect 4016 5272 4056 5312
rect 3688 3760 3728 3800
rect 3770 3760 3810 3800
rect 3852 3760 3892 3800
rect 3934 3760 3974 3800
rect 4016 3760 4056 3800
rect 2764 2584 2804 2624
rect 2476 2332 2516 2372
rect 5548 17872 5588 17912
rect 5068 16864 5108 16904
rect 4928 16612 4968 16652
rect 5010 16612 5050 16652
rect 5092 16612 5132 16652
rect 5174 16612 5214 16652
rect 5256 16612 5296 16652
rect 4972 16276 5012 16316
rect 4928 15100 4968 15140
rect 5010 15100 5050 15140
rect 5092 15100 5132 15140
rect 5174 15100 5214 15140
rect 5256 15100 5296 15140
rect 6220 39124 6260 39164
rect 6220 38200 6260 38240
rect 6124 37780 6164 37820
rect 6316 37948 6356 37988
rect 7468 45424 7508 45464
rect 7564 45340 7604 45380
rect 7084 43660 7124 43700
rect 6892 42736 6932 42776
rect 6508 39124 6548 39164
rect 6796 39796 6836 39836
rect 6604 39040 6644 39080
rect 6700 39376 6740 39416
rect 6892 40216 6932 40256
rect 7180 42736 7220 42776
rect 7084 40804 7124 40844
rect 6988 39460 7028 39500
rect 7180 40552 7220 40592
rect 7084 39712 7124 39752
rect 6988 39208 7028 39248
rect 6892 39040 6932 39080
rect 6508 38032 6548 38072
rect 6412 37780 6452 37820
rect 6508 37864 6548 37904
rect 6220 32488 6260 32528
rect 6124 31900 6164 31940
rect 6124 31228 6164 31268
rect 6220 30724 6260 30764
rect 6124 29380 6164 29420
rect 6028 29296 6068 29336
rect 6124 28876 6164 28916
rect 6124 26356 6164 26396
rect 6220 28204 6260 28244
rect 6028 26272 6068 26312
rect 5932 25012 5972 25052
rect 5932 23164 5972 23204
rect 5740 23080 5780 23120
rect 6124 23164 6164 23204
rect 6028 22240 6068 22280
rect 6124 20644 6164 20684
rect 5932 19720 5972 19760
rect 5356 13840 5396 13880
rect 5740 17368 5780 17408
rect 4928 13588 4968 13628
rect 5010 13588 5050 13628
rect 5092 13588 5132 13628
rect 5174 13588 5214 13628
rect 5256 13588 5296 13628
rect 4876 12664 4916 12704
rect 4928 12076 4968 12116
rect 5010 12076 5050 12116
rect 5092 12076 5132 12116
rect 5174 12076 5214 12116
rect 5256 12076 5296 12116
rect 5260 11908 5300 11948
rect 4972 11572 5012 11612
rect 4928 10564 4968 10604
rect 5010 10564 5050 10604
rect 5092 10564 5132 10604
rect 5174 10564 5214 10604
rect 5256 10564 5296 10604
rect 5164 10396 5204 10436
rect 4928 9052 4968 9092
rect 5010 9052 5050 9092
rect 5092 9052 5132 9092
rect 5174 9052 5214 9092
rect 5256 9052 5296 9092
rect 5356 8968 5396 9008
rect 5068 8884 5108 8924
rect 5356 8800 5396 8840
rect 4928 7540 4968 7580
rect 5010 7540 5050 7580
rect 5092 7540 5132 7580
rect 5174 7540 5214 7580
rect 5256 7540 5296 7580
rect 5548 13672 5588 13712
rect 5644 11908 5684 11948
rect 6412 29380 6452 29420
rect 6796 38032 6836 38072
rect 6988 38368 7028 38408
rect 6892 37780 6932 37820
rect 6988 38116 7028 38156
rect 7372 40636 7412 40676
rect 7372 40468 7412 40508
rect 7276 38956 7316 38996
rect 7084 37948 7124 37988
rect 6604 28204 6644 28244
rect 7276 38116 7316 38156
rect 7372 38200 7412 38240
rect 7276 37276 7316 37316
rect 7084 32068 7124 32108
rect 6892 31816 6932 31856
rect 6892 31480 6932 31520
rect 6796 31060 6836 31100
rect 6796 28372 6836 28412
rect 6412 20980 6452 21020
rect 6124 19216 6164 19256
rect 6124 18796 6164 18836
rect 6220 17704 6260 17744
rect 6124 16948 6164 16988
rect 6124 16444 6164 16484
rect 5836 13840 5876 13880
rect 5932 12832 5972 12872
rect 5836 12496 5876 12536
rect 5836 10396 5876 10436
rect 5932 10228 5972 10268
rect 5836 9640 5876 9680
rect 4928 6028 4968 6068
rect 5010 6028 5050 6068
rect 5092 6028 5132 6068
rect 5174 6028 5214 6068
rect 5256 6028 5296 6068
rect 4876 5608 4916 5648
rect 4780 5440 4820 5480
rect 2284 2080 2324 2120
rect 2572 2080 2612 2120
rect 2476 1744 2516 1784
rect 4928 4516 4968 4556
rect 5010 4516 5050 4556
rect 5092 4516 5132 4556
rect 5174 4516 5214 4556
rect 5256 4516 5296 4556
rect 3532 2752 3572 2792
rect 3340 2080 3380 2120
rect 3688 2248 3728 2288
rect 3770 2248 3810 2288
rect 3852 2248 3892 2288
rect 3934 2248 3974 2288
rect 4016 2248 4056 2288
rect 4204 2164 4244 2204
rect 5356 4264 5396 4304
rect 4684 3760 4724 3800
rect 4928 3004 4968 3044
rect 5010 3004 5050 3044
rect 5092 3004 5132 3044
rect 5174 3004 5214 3044
rect 5256 3004 5296 3044
rect 4876 2836 4916 2876
rect 5548 3508 5588 3548
rect 4928 1492 4968 1532
rect 5010 1492 5050 1532
rect 5092 1492 5132 1532
rect 5174 1492 5214 1532
rect 5256 1492 5296 1532
rect 5260 988 5300 1028
rect 6124 15772 6164 15812
rect 6220 15100 6260 15140
rect 6220 14008 6260 14048
rect 6220 10228 6260 10268
rect 6508 18544 6548 18584
rect 6892 27952 6932 27992
rect 6700 25348 6740 25388
rect 6796 25600 6836 25640
rect 6508 16444 6548 16484
rect 6604 15604 6644 15644
rect 7084 25600 7124 25640
rect 7468 36268 7508 36308
rect 7372 33100 7412 33140
rect 7372 32992 7412 33032
rect 7276 32656 7316 32696
rect 7660 43492 7700 43532
rect 7756 42568 7796 42608
rect 8908 57268 8948 57308
rect 9004 54832 9044 54872
rect 9292 54832 9332 54872
rect 9100 51640 9140 51680
rect 8620 47188 8660 47228
rect 7756 41056 7796 41096
rect 7660 39964 7700 40004
rect 8044 41224 8084 41264
rect 8044 40048 8084 40088
rect 7468 32656 7508 32696
rect 7276 30724 7316 30764
rect 7660 36268 7700 36308
rect 7756 32824 7796 32864
rect 7276 30388 7316 30428
rect 7276 30220 7316 30260
rect 7372 29716 7412 29756
rect 7372 28960 7376 29000
rect 7376 28960 7412 29000
rect 7276 26440 7316 26480
rect 7276 25516 7316 25556
rect 6988 24928 7028 24968
rect 6988 24592 7028 24632
rect 6796 21820 6836 21860
rect 6796 21652 6836 21692
rect 6988 21652 7028 21692
rect 7084 22576 7124 22616
rect 6700 15184 6740 15224
rect 6604 15100 6644 15140
rect 6604 13756 6644 13796
rect 6604 12580 6644 12620
rect 6412 10312 6452 10352
rect 6604 11152 6644 11192
rect 7468 25936 7508 25976
rect 7468 24928 7508 24968
rect 7468 24508 7508 24548
rect 7756 30136 7796 30176
rect 8044 32404 8084 32444
rect 8428 43576 8468 43616
rect 8236 38872 8276 38912
rect 8236 35932 8276 35972
rect 8620 45592 8660 45632
rect 8716 44416 8756 44456
rect 8428 38956 8468 38996
rect 8428 34588 8468 34628
rect 8524 36016 8564 36056
rect 7948 31816 7988 31856
rect 7948 31312 7988 31352
rect 7948 30052 7988 30092
rect 7852 28372 7892 28412
rect 7948 27448 7988 27488
rect 7852 26776 7892 26816
rect 7660 25180 7700 25220
rect 7564 24340 7604 24380
rect 7084 20140 7124 20180
rect 7084 19972 7124 20012
rect 7372 23080 7412 23120
rect 7372 21568 7412 21608
rect 7372 18796 7412 18836
rect 7276 18628 7316 18668
rect 7180 17536 7220 17576
rect 6988 16192 7028 16232
rect 7180 16444 7220 16484
rect 6892 13420 6932 13460
rect 6988 14680 7028 14720
rect 7084 13756 7124 13796
rect 6892 11152 6932 11192
rect 6124 6868 6164 6908
rect 5836 5944 5876 5984
rect 6700 8800 6740 8840
rect 7564 16948 7604 16988
rect 7276 14680 7316 14720
rect 7372 13840 7412 13880
rect 7372 13420 7412 13460
rect 7180 12832 7220 12872
rect 6700 3088 6740 3128
rect 5548 988 5588 1028
rect 6028 2332 6068 2372
rect 6892 2080 6932 2120
rect 7084 1996 7124 2036
rect 7180 1156 7220 1196
rect 7948 26608 7988 26648
rect 7948 26020 7988 26060
rect 8236 31312 8276 31352
rect 8332 28540 8372 28580
rect 8140 26104 8180 26144
rect 7948 24592 7988 24632
rect 7852 23164 7892 23204
rect 7852 22912 7892 22952
rect 8140 23080 8180 23120
rect 8044 21820 8084 21860
rect 7852 19888 7892 19928
rect 7756 17956 7796 17996
rect 8140 18460 8180 18500
rect 8044 17956 8084 17996
rect 7852 16864 7892 16904
rect 7564 11824 7604 11864
rect 7948 9976 7988 10016
rect 7756 3340 7796 3380
rect 7756 1408 7796 1448
rect 7564 316 7604 356
rect 8332 23752 8372 23792
rect 8524 26020 8564 26060
rect 8332 22576 8372 22616
rect 8428 22240 8468 22280
rect 8332 20896 8372 20936
rect 8332 19300 8372 19340
rect 8428 18880 8468 18920
rect 8908 45760 8948 45800
rect 8812 40216 8852 40256
rect 8908 40300 8948 40340
rect 9292 51640 9332 51680
rect 9196 48700 9236 48740
rect 9676 79864 9716 79904
rect 9676 79612 9716 79652
rect 10060 89440 10100 89480
rect 9964 83644 10004 83684
rect 9964 83476 10004 83516
rect 10156 84988 10196 85028
rect 10156 80704 10196 80744
rect 10156 78688 10196 78728
rect 9868 77344 9908 77384
rect 10060 76420 10100 76460
rect 9772 70960 9812 71000
rect 9676 70540 9716 70580
rect 10060 75412 10100 75452
rect 10060 73312 10100 73352
rect 9964 72136 10004 72176
rect 10060 70624 10100 70664
rect 10060 70456 10100 70496
rect 9676 68608 9716 68648
rect 9676 66760 9716 66800
rect 9676 65248 9716 65288
rect 9580 61132 9620 61172
rect 9868 68188 9908 68228
rect 10060 68608 10100 68648
rect 10060 68104 10100 68144
rect 10444 85576 10484 85616
rect 10444 82048 10484 82088
rect 10636 84148 10676 84188
rect 10636 82048 10676 82088
rect 10636 79780 10676 79820
rect 10540 79024 10580 79064
rect 10540 78856 10580 78896
rect 10540 78268 10580 78308
rect 10444 78100 10484 78140
rect 10252 76924 10292 76964
rect 10252 76672 10292 76712
rect 10540 77428 10580 77468
rect 10444 76588 10484 76628
rect 10732 77260 10772 77300
rect 10732 76840 10772 76880
rect 10252 70456 10292 70496
rect 10252 69280 10292 69320
rect 10252 65500 10292 65540
rect 10348 67516 10388 67556
rect 10156 64744 10196 64784
rect 9964 63904 10004 63944
rect 9964 62728 10004 62768
rect 9964 62392 10004 62432
rect 10348 63652 10388 63692
rect 10540 76252 10580 76292
rect 10732 75916 10772 75956
rect 10540 70036 10580 70076
rect 10636 70792 10676 70832
rect 9868 61132 9908 61172
rect 9580 54160 9620 54200
rect 9388 45508 9428 45548
rect 9196 40216 9236 40256
rect 8908 34840 8948 34880
rect 8812 34672 8852 34712
rect 8908 33244 8948 33284
rect 9004 32404 9044 32444
rect 8716 29884 8756 29924
rect 8716 29380 8756 29420
rect 9004 30892 9044 30932
rect 8908 30472 8948 30512
rect 9196 34420 9236 34460
rect 9772 53068 9812 53108
rect 9772 49540 9812 49580
rect 9964 58696 10004 58736
rect 10060 56512 10100 56552
rect 10156 53320 10196 53360
rect 10060 50296 10100 50336
rect 10156 50212 10196 50252
rect 10156 49540 10196 49580
rect 10636 64324 10676 64364
rect 10924 78688 10964 78728
rect 12364 94732 12404 94772
rect 11596 94648 11636 94688
rect 12172 94648 12212 94688
rect 11500 94144 11540 94184
rect 11212 88012 11252 88052
rect 11020 78520 11060 78560
rect 10924 76588 10964 76628
rect 11212 80368 11252 80408
rect 11212 79948 11252 79988
rect 11212 78940 11252 78980
rect 11212 78436 11252 78476
rect 11116 73648 11156 73688
rect 11020 70372 11060 70412
rect 11500 84652 11540 84692
rect 10348 59368 10388 59408
rect 10444 58444 10484 58484
rect 10540 57772 10580 57812
rect 11212 65164 11252 65204
rect 10444 53824 10484 53864
rect 11116 61804 11156 61844
rect 13228 94732 13268 94772
rect 11980 84484 12020 84524
rect 11596 73396 11636 73436
rect 12076 83308 12116 83348
rect 11788 80620 11828 80660
rect 11500 72220 11540 72260
rect 11596 71968 11636 72008
rect 11116 59284 11156 59324
rect 11212 58948 11252 58988
rect 11020 58360 11060 58400
rect 10924 58108 10964 58148
rect 11212 58528 11252 58568
rect 10924 57940 10964 57980
rect 10924 57688 10964 57728
rect 10636 53824 10676 53864
rect 10636 53404 10676 53444
rect 10540 53068 10580 53108
rect 10348 52732 10388 52772
rect 10732 52732 10772 52772
rect 10924 53404 10964 53444
rect 11116 50464 11156 50504
rect 10732 49540 10772 49580
rect 9676 48784 9716 48824
rect 9484 39376 9524 39416
rect 9484 37696 9524 37736
rect 9484 33244 9524 33284
rect 9580 32992 9620 33032
rect 9100 29800 9140 29840
rect 8812 29044 8852 29084
rect 8812 24844 8852 24884
rect 8812 21148 8852 21188
rect 9292 32236 9332 32276
rect 9868 44164 9908 44204
rect 9772 40636 9812 40676
rect 9772 40384 9812 40424
rect 10636 47860 10676 47900
rect 10252 46516 10292 46556
rect 10156 46432 10196 46472
rect 10444 46600 10484 46640
rect 10252 41728 10292 41768
rect 10156 41140 10196 41180
rect 9964 40552 10004 40592
rect 10540 44080 10580 44120
rect 10444 42736 10484 42776
rect 10348 40804 10388 40844
rect 10060 40300 10100 40340
rect 10060 39712 10100 39752
rect 10252 39796 10292 39836
rect 10156 39544 10196 39584
rect 10060 39376 10100 39416
rect 9964 39040 10004 39080
rect 10060 37528 10100 37568
rect 9868 34420 9908 34460
rect 9388 31984 9428 32024
rect 9292 31228 9332 31268
rect 9292 29800 9332 29840
rect 9388 29716 9428 29756
rect 9292 29632 9332 29672
rect 9292 29380 9332 29420
rect 9580 31984 9620 32024
rect 9676 29884 9716 29924
rect 9292 27028 9332 27068
rect 9292 26272 9332 26312
rect 9100 25600 9140 25640
rect 9196 25852 9236 25892
rect 9100 25432 9140 25472
rect 9100 23668 9140 23708
rect 9004 23080 9044 23120
rect 8620 20812 8660 20852
rect 8524 18460 8564 18500
rect 8332 17452 8372 17492
rect 9196 20896 9236 20936
rect 8524 17452 8564 17492
rect 9100 20560 9140 20600
rect 8620 16192 8660 16232
rect 8620 15268 8660 15308
rect 8524 14008 8564 14048
rect 8908 17368 8948 17408
rect 8812 14848 8852 14888
rect 8812 14008 8852 14048
rect 9868 32992 9908 33032
rect 9676 25600 9716 25640
rect 9772 25348 9812 25388
rect 9676 23668 9716 23708
rect 9676 23164 9716 23204
rect 9292 19216 9332 19256
rect 9196 16360 9236 16400
rect 9004 14596 9044 14636
rect 8908 12664 8948 12704
rect 8812 12244 8852 12284
rect 8524 10480 8564 10520
rect 9484 14596 9524 14636
rect 9292 11656 9332 11696
rect 8812 7120 8852 7160
rect 8428 2836 8468 2876
rect 9100 7876 9140 7916
rect 8140 1408 8180 1448
rect 8332 1408 8372 1448
rect 8524 1408 8564 1448
rect 9004 1912 9044 1952
rect 9964 32236 10004 32276
rect 10348 37612 10388 37652
rect 10348 37276 10388 37316
rect 10732 44080 10772 44120
rect 10828 41476 10868 41516
rect 11500 66928 11540 66968
rect 11500 64324 11540 64364
rect 11788 79696 11828 79736
rect 11788 79192 11828 79232
rect 11788 77428 11828 77468
rect 11980 79948 12020 79988
rect 11980 79696 12020 79736
rect 11980 78268 12020 78308
rect 11884 73396 11924 73436
rect 11788 71296 11828 71336
rect 11788 69364 11828 69404
rect 12556 89188 12596 89228
rect 12460 86164 12500 86204
rect 12556 86080 12596 86120
rect 12364 85828 12404 85868
rect 12460 84904 12500 84944
rect 12268 83644 12308 83684
rect 12268 80452 12308 80492
rect 12556 84316 12596 84356
rect 12172 79192 12212 79232
rect 12172 78772 12212 78812
rect 12172 77428 12212 77468
rect 11980 73144 12020 73184
rect 12076 73396 12116 73436
rect 12076 71968 12116 72008
rect 11980 71296 12020 71336
rect 11788 63568 11828 63608
rect 11500 58360 11540 58400
rect 11404 50296 11444 50336
rect 11308 50044 11348 50084
rect 11020 43492 11060 43532
rect 11788 59620 11828 59660
rect 12172 66340 12212 66380
rect 12172 66172 12212 66212
rect 12076 63652 12116 63692
rect 12364 79864 12404 79904
rect 12460 78772 12500 78812
rect 12364 78100 12404 78140
rect 11788 57772 11828 57812
rect 11884 57688 11924 57728
rect 11596 50380 11636 50420
rect 11692 50464 11732 50504
rect 12172 62980 12212 63020
rect 12268 60208 12308 60248
rect 12172 60040 12212 60080
rect 12268 59200 12308 59240
rect 12172 58696 12212 58736
rect 12172 58444 12212 58484
rect 12172 58192 12212 58232
rect 12076 57940 12116 57980
rect 12076 57520 12116 57560
rect 11788 48196 11828 48236
rect 11500 46096 11540 46136
rect 11116 42064 11156 42104
rect 11020 41140 11060 41180
rect 10732 40972 10772 41012
rect 10540 38116 10580 38156
rect 10540 35008 10580 35048
rect 10444 34420 10484 34460
rect 10156 33244 10196 33284
rect 10060 28876 10100 28916
rect 10252 30052 10292 30092
rect 10060 28288 10100 28328
rect 10060 27952 10100 27992
rect 9964 26860 10004 26900
rect 10060 26524 10100 26564
rect 9964 26188 10004 26228
rect 10060 26104 10100 26144
rect 9964 26020 10004 26060
rect 10060 25768 10100 25808
rect 9964 25264 10004 25304
rect 9964 23584 10004 23624
rect 10540 32236 10580 32276
rect 10444 31984 10484 32024
rect 10444 30052 10484 30092
rect 10444 29884 10484 29924
rect 10444 28876 10484 28916
rect 10252 23752 10292 23792
rect 10348 28624 10388 28664
rect 10156 23332 10196 23372
rect 10252 23584 10292 23624
rect 9964 22408 10004 22448
rect 9964 20140 10004 20180
rect 10636 29800 10676 29840
rect 10636 28708 10676 28748
rect 10348 21484 10388 21524
rect 10348 21232 10388 21272
rect 9868 16948 9908 16988
rect 9772 12496 9812 12536
rect 9868 9304 9908 9344
rect 10060 9388 10100 9428
rect 10924 41056 10964 41096
rect 10924 39712 10964 39752
rect 11020 39544 11060 39584
rect 11116 38872 11156 38912
rect 11020 38116 11060 38156
rect 10924 33748 10964 33788
rect 10828 32068 10868 32108
rect 10924 32908 10964 32948
rect 10828 30808 10868 30848
rect 10924 29884 10964 29924
rect 10924 28876 10964 28916
rect 10828 27532 10868 27572
rect 10732 20224 10772 20264
rect 10348 11656 10388 11696
rect 10156 9220 10196 9260
rect 10060 8884 10100 8924
rect 9964 7876 10004 7916
rect 9484 5524 9524 5564
rect 9676 6028 9716 6068
rect 9196 2668 9236 2708
rect 10060 6112 10100 6152
rect 10060 5188 10100 5228
rect 11020 27616 11060 27656
rect 11020 20308 11060 20348
rect 10924 20056 10964 20096
rect 10828 10984 10868 11024
rect 10828 10816 10868 10856
rect 11212 33412 11252 33452
rect 11212 33244 11252 33284
rect 11596 42652 11636 42692
rect 11596 41056 11636 41096
rect 11596 40132 11636 40172
rect 11500 39796 11540 39836
rect 11500 37864 11540 37904
rect 11692 37864 11732 37904
rect 11500 36436 11540 36476
rect 11500 35008 11540 35048
rect 11692 37444 11732 37484
rect 12268 50296 12308 50336
rect 11980 40888 12020 40928
rect 11980 40216 12020 40256
rect 11980 39964 12020 40004
rect 11788 36856 11828 36896
rect 11788 36688 11828 36728
rect 11692 36436 11732 36476
rect 11308 29380 11348 29420
rect 11212 27616 11252 27656
rect 11692 32740 11732 32780
rect 11788 30304 11828 30344
rect 12268 48616 12308 48656
rect 12268 46096 12308 46136
rect 12556 73900 12596 73940
rect 12940 93892 12980 93932
rect 14284 95908 14324 95948
rect 14380 94732 14420 94772
rect 14668 96580 14708 96620
rect 13900 93892 13940 93932
rect 14284 93892 14324 93932
rect 13036 93724 13076 93764
rect 13228 89188 13268 89228
rect 12844 87928 12884 87968
rect 13132 87928 13172 87968
rect 12940 87340 12980 87380
rect 13036 86416 13076 86456
rect 12844 86164 12884 86204
rect 12748 85240 12788 85280
rect 12940 84988 12980 85028
rect 13324 87340 13364 87380
rect 13228 86080 13268 86120
rect 13228 83980 13268 84020
rect 13228 83560 13268 83600
rect 12748 82804 12788 82844
rect 12748 80536 12788 80576
rect 13036 80452 13076 80492
rect 12748 79864 12788 79904
rect 12940 79696 12980 79736
rect 13036 78520 13076 78560
rect 12844 76420 12884 76460
rect 14668 93892 14708 93932
rect 14476 90700 14516 90740
rect 13708 85240 13748 85280
rect 13324 81712 13364 81752
rect 13324 80536 13364 80576
rect 13132 76252 13172 76292
rect 12844 76084 12884 76124
rect 12748 74656 12788 74696
rect 12748 74404 12788 74444
rect 13324 76252 13364 76292
rect 13132 75748 13172 75788
rect 13132 73816 13172 73856
rect 12460 70792 12500 70832
rect 12652 73144 12692 73184
rect 12844 73312 12884 73352
rect 12940 73144 12980 73184
rect 13036 73564 13076 73604
rect 12844 72220 12884 72260
rect 12844 71380 12884 71420
rect 13132 70876 13172 70916
rect 13036 70792 13076 70832
rect 13516 83644 13556 83684
rect 13612 83980 13652 84020
rect 13516 81544 13556 81584
rect 13516 78772 13556 78812
rect 13708 83896 13748 83936
rect 14284 89020 14324 89060
rect 14188 85156 14228 85196
rect 14188 84988 14228 85028
rect 14188 84652 14228 84692
rect 14092 83896 14132 83936
rect 13804 81796 13844 81836
rect 14092 83728 14132 83768
rect 14284 83644 14324 83684
rect 14380 83140 14420 83180
rect 14476 84232 14516 84272
rect 14092 82720 14132 82760
rect 14092 82468 14132 82508
rect 14092 81796 14132 81836
rect 13900 79276 13940 79316
rect 13996 81712 14036 81752
rect 13612 78100 13652 78140
rect 13900 78856 13940 78896
rect 13324 75076 13364 75116
rect 13324 74488 13364 74528
rect 13804 78268 13844 78308
rect 13708 76084 13748 76124
rect 13612 75916 13652 75956
rect 13804 74236 13844 74276
rect 14380 82048 14420 82088
rect 14572 84148 14612 84188
rect 14092 78016 14132 78056
rect 14092 76672 14132 76712
rect 13900 74068 13940 74108
rect 13708 73144 13748 73184
rect 13420 71044 13460 71084
rect 13900 73732 13940 73772
rect 13324 69112 13364 69152
rect 12940 68272 12980 68312
rect 13132 67096 13172 67136
rect 12748 65332 12788 65372
rect 13612 70372 13652 70412
rect 13420 68356 13460 68396
rect 13420 67768 13460 67808
rect 13708 67180 13748 67220
rect 12556 64072 12596 64112
rect 12748 63568 12788 63608
rect 12652 63400 12692 63440
rect 12940 64996 12980 65036
rect 13132 64996 13172 65036
rect 12844 62476 12884 62516
rect 12556 61132 12596 61172
rect 12652 60292 12692 60332
rect 12652 60040 12692 60080
rect 12940 58948 12980 58988
rect 13420 63484 13460 63524
rect 13324 63232 13364 63272
rect 13228 63148 13268 63188
rect 12940 57856 12980 57896
rect 13036 58612 13076 58652
rect 13132 58528 13172 58568
rect 13132 58276 13172 58316
rect 13324 63064 13364 63104
rect 13612 64828 13652 64868
rect 13804 64660 13844 64700
rect 14188 75916 14228 75956
rect 15436 95656 15476 95696
rect 15148 93892 15188 93932
rect 14860 89356 14900 89396
rect 14860 84316 14900 84356
rect 14764 83056 14804 83096
rect 16204 94144 16244 94184
rect 15340 87844 15380 87884
rect 15052 84484 15092 84524
rect 15244 84904 15284 84944
rect 15052 83560 15092 83600
rect 14860 82132 14900 82172
rect 15244 82468 15284 82508
rect 15340 83140 15380 83180
rect 14764 81796 14804 81836
rect 14860 81964 14900 82004
rect 14188 74572 14228 74612
rect 14284 75076 14324 75116
rect 14092 74488 14132 74528
rect 14188 74236 14228 74276
rect 14092 74068 14132 74108
rect 14188 69112 14228 69152
rect 13996 68944 14036 68984
rect 14188 68944 14228 68984
rect 13996 68272 14036 68312
rect 14092 63904 14132 63944
rect 13900 63736 13940 63776
rect 13996 63652 14036 63692
rect 13612 63316 13652 63356
rect 13708 63232 13748 63272
rect 13516 62224 13556 62264
rect 13516 58444 13556 58484
rect 13228 57352 13268 57392
rect 13324 53320 13364 53360
rect 12748 48700 12788 48740
rect 12364 46012 12404 46052
rect 12460 48616 12500 48656
rect 12556 46264 12596 46304
rect 12556 46012 12596 46052
rect 12748 48196 12788 48236
rect 13900 63148 13940 63188
rect 14092 63400 14132 63440
rect 14092 62896 14132 62936
rect 13996 62392 14036 62432
rect 13804 56260 13844 56300
rect 14668 77428 14708 77468
rect 14380 68608 14420 68648
rect 14380 66508 14420 66548
rect 14284 63652 14324 63692
rect 14284 63484 14324 63524
rect 14092 53320 14132 53360
rect 14380 63316 14420 63356
rect 14380 63148 14420 63188
rect 14380 61720 14420 61760
rect 14380 60208 14420 60248
rect 14380 60040 14420 60080
rect 14284 57772 14324 57812
rect 14284 53488 14324 53528
rect 14860 78772 14900 78812
rect 14860 78184 14900 78224
rect 14860 76420 14900 76460
rect 14860 76168 14900 76208
rect 14764 76000 14804 76040
rect 14572 71380 14612 71420
rect 14572 71212 14612 71252
rect 15340 82132 15380 82172
rect 15052 79108 15092 79148
rect 15148 78772 15188 78812
rect 15052 76336 15092 76376
rect 14956 72388 14996 72428
rect 15052 73480 15092 73520
rect 14956 71380 14996 71420
rect 14860 71296 14900 71336
rect 14572 65920 14612 65960
rect 14668 65332 14708 65372
rect 14764 65920 14804 65960
rect 14860 64660 14900 64700
rect 14764 64324 14804 64364
rect 14668 60124 14708 60164
rect 14668 59788 14708 59828
rect 14668 59368 14708 59408
rect 14764 58108 14804 58148
rect 14476 54160 14516 54200
rect 14380 53320 14420 53360
rect 13036 43240 13076 43280
rect 12748 41896 12788 41936
rect 12364 40468 12404 40508
rect 12652 40804 12692 40844
rect 12268 39712 12308 39752
rect 12364 39544 12404 39584
rect 12556 40216 12596 40256
rect 13036 43072 13076 43112
rect 12940 41896 12980 41936
rect 12940 40804 12980 40844
rect 12844 40300 12884 40340
rect 13324 43072 13364 43112
rect 13612 44164 13652 44204
rect 13612 42316 13652 42356
rect 13804 42736 13844 42776
rect 13804 41644 13844 41684
rect 13228 40552 13268 40592
rect 12940 40132 12980 40172
rect 12652 39544 12692 39584
rect 12652 39208 12692 39248
rect 12748 38872 12788 38912
rect 12460 37276 12500 37316
rect 11980 36100 12020 36140
rect 11980 35932 12020 35972
rect 12364 36100 12404 36140
rect 12268 35848 12308 35888
rect 12172 35260 12212 35300
rect 11692 29296 11732 29336
rect 11692 28456 11732 28496
rect 11308 27112 11348 27152
rect 11404 26860 11444 26900
rect 11500 27364 11540 27404
rect 11212 21904 11252 21944
rect 11116 20224 11156 20264
rect 11020 14344 11060 14384
rect 11212 14344 11252 14384
rect 10924 4180 10964 4220
rect 10060 2920 10100 2960
rect 9388 2332 9428 2372
rect 9772 2416 9812 2456
rect 10348 2584 10388 2624
rect 11788 27616 11828 27656
rect 11596 26020 11636 26060
rect 11500 22324 11540 22364
rect 11500 22072 11540 22112
rect 12076 31060 12116 31100
rect 11980 27532 12020 27572
rect 11788 22996 11828 23036
rect 11788 21568 11828 21608
rect 11692 20224 11732 20264
rect 11404 13924 11444 13964
rect 11308 10816 11348 10856
rect 11404 10060 11444 10100
rect 12268 29212 12308 29252
rect 12940 39712 12980 39752
rect 13036 39544 13076 39584
rect 13228 40300 13268 40340
rect 13228 39376 13268 39416
rect 13132 39208 13172 39248
rect 13036 38200 13076 38240
rect 12556 36688 12596 36728
rect 12652 37276 12692 37316
rect 12460 35848 12500 35888
rect 12460 35680 12500 35720
rect 12748 36856 12788 36896
rect 13228 38956 13268 38996
rect 13516 39712 13556 39752
rect 13516 39376 13556 39416
rect 13516 38200 13556 38240
rect 13420 37612 13460 37652
rect 12748 35932 12788 35972
rect 13036 35932 13076 35972
rect 12460 34504 12500 34544
rect 12460 32488 12500 32528
rect 12172 27532 12212 27572
rect 12268 26608 12308 26648
rect 12076 20224 12116 20264
rect 12364 25012 12404 25052
rect 13804 39208 13844 39248
rect 13996 41980 14036 42020
rect 13804 38956 13844 38996
rect 13420 36184 13460 36224
rect 13228 33160 13268 33200
rect 13228 32992 13268 33032
rect 12844 30976 12884 31016
rect 12940 30724 12980 30764
rect 12844 29968 12884 30008
rect 12940 29800 12980 29840
rect 12556 29044 12596 29084
rect 12652 29212 12692 29252
rect 12844 29632 12884 29672
rect 12652 26944 12692 26984
rect 13132 31480 13172 31520
rect 13132 30892 13172 30932
rect 13132 30472 13172 30512
rect 13132 30304 13172 30344
rect 13132 29212 13172 29252
rect 13036 26944 13076 26984
rect 12940 26104 12980 26144
rect 12460 23416 12500 23456
rect 12364 21400 12404 21440
rect 12076 17956 12116 17996
rect 12940 23416 12980 23456
rect 13132 25852 13172 25892
rect 13708 36688 13748 36728
rect 13804 36604 13844 36644
rect 13612 36520 13652 36560
rect 13708 36436 13748 36476
rect 13804 36184 13844 36224
rect 13708 32992 13748 33032
rect 13324 29716 13364 29756
rect 13324 29128 13364 29168
rect 13132 24172 13172 24212
rect 13228 24340 13268 24380
rect 12844 22996 12884 23036
rect 12940 20644 12980 20684
rect 12556 17956 12596 17996
rect 12268 14512 12308 14552
rect 12076 12412 12116 12452
rect 11308 1996 11348 2036
rect 11500 1912 11540 1952
rect 12652 14260 12692 14300
rect 12556 5188 12596 5228
rect 13324 24172 13364 24212
rect 13324 20056 13364 20096
rect 13036 14680 13076 14720
rect 12940 13168 12980 13208
rect 12940 12412 12980 12452
rect 13228 13756 13268 13796
rect 13132 13084 13172 13124
rect 13036 7792 13076 7832
rect 12268 2416 12308 2456
rect 13036 3424 13076 3464
rect 12652 1996 12692 2036
rect 13516 29044 13556 29084
rect 13804 31984 13844 32024
rect 13996 40552 14036 40592
rect 14572 50968 14612 51008
rect 14188 44920 14228 44960
rect 14380 44920 14420 44960
rect 14188 42652 14228 42692
rect 14380 42820 14420 42860
rect 14188 41728 14228 41768
rect 14188 41392 14228 41432
rect 14188 41056 14228 41096
rect 14092 39544 14132 39584
rect 13996 38872 14036 38912
rect 13900 31648 13940 31688
rect 13900 29968 13940 30008
rect 13708 29464 13748 29504
rect 14188 36688 14228 36728
rect 13708 29212 13748 29252
rect 14092 32908 14132 32948
rect 13804 29128 13844 29168
rect 13516 25852 13556 25892
rect 13708 27532 13748 27572
rect 13804 26860 13844 26900
rect 13708 23164 13748 23204
rect 13612 21400 13652 21440
rect 13420 13168 13460 13208
rect 13996 26272 14036 26312
rect 13996 23752 14036 23792
rect 13900 22996 13940 23036
rect 13900 19972 13940 20012
rect 14476 42232 14516 42272
rect 14572 41476 14612 41516
rect 14572 40720 14612 40760
rect 14476 39460 14516 39500
rect 14380 38956 14420 38996
rect 14380 38788 14420 38828
rect 14380 36016 14420 36056
rect 14476 38116 14516 38156
rect 14380 35512 14420 35552
rect 14380 32236 14420 32276
rect 14188 31312 14228 31352
rect 14284 31648 14324 31688
rect 14188 29884 14228 29924
rect 14380 30724 14420 30764
rect 15052 66844 15092 66884
rect 15052 63316 15092 63356
rect 15052 62812 15092 62852
rect 15052 61468 15092 61508
rect 14956 59284 14996 59324
rect 14860 45676 14900 45716
rect 14956 43996 14996 44036
rect 14860 43324 14900 43364
rect 14764 39124 14804 39164
rect 14860 43072 14900 43112
rect 15052 43324 15092 43364
rect 14956 42988 14996 43028
rect 15052 42904 15092 42944
rect 14860 38116 14900 38156
rect 14764 37864 14804 37904
rect 14668 36436 14708 36476
rect 14572 36016 14612 36056
rect 15052 40972 15092 41012
rect 15052 40720 15092 40760
rect 15052 38368 15092 38408
rect 15052 38200 15092 38240
rect 14860 35764 14900 35804
rect 14860 35512 14900 35552
rect 14668 35008 14708 35048
rect 14668 34420 14708 34460
rect 14764 32068 14804 32108
rect 14476 30640 14516 30680
rect 14476 30388 14516 30428
rect 14476 29716 14516 29756
rect 14476 29380 14516 29420
rect 14668 30304 14708 30344
rect 14764 30640 14804 30680
rect 15052 31312 15092 31352
rect 14572 28708 14612 28748
rect 14956 29632 14996 29672
rect 14956 29296 14996 29336
rect 14764 27952 14804 27992
rect 14188 23668 14228 23708
rect 14284 23248 14324 23288
rect 14284 22576 14324 22616
rect 14668 26860 14708 26900
rect 14476 26104 14516 26144
rect 14476 24760 14516 24800
rect 14476 22576 14516 22616
rect 14092 19972 14132 20012
rect 13900 17452 13940 17492
rect 13516 12748 13556 12788
rect 13324 9556 13364 9596
rect 13708 12748 13748 12788
rect 13804 11740 13844 11780
rect 13996 11320 14036 11360
rect 13900 9556 13940 9596
rect 13900 9052 13940 9092
rect 13708 8716 13748 8756
rect 13708 7792 13748 7832
rect 13612 2752 13652 2792
rect 13996 5692 14036 5732
rect 13996 5524 14036 5564
rect 14188 17452 14228 17492
rect 14284 21736 14324 21776
rect 14764 20140 14804 20180
rect 14764 19720 14804 19760
rect 14380 19048 14420 19088
rect 15052 28708 15092 28748
rect 14956 24592 14996 24632
rect 14956 23164 14996 23204
rect 15340 74404 15380 74444
rect 17356 95572 17396 95612
rect 16972 94144 17012 94184
rect 16588 93892 16628 93932
rect 16012 84736 16052 84776
rect 15724 84232 15764 84272
rect 15628 83476 15668 83516
rect 15628 81712 15668 81752
rect 16012 83644 16052 83684
rect 16300 89020 16340 89060
rect 16108 82636 16148 82676
rect 15628 80368 15668 80408
rect 15628 79024 15668 79064
rect 15820 79780 15860 79820
rect 15724 78184 15764 78224
rect 15724 77428 15764 77468
rect 15244 73228 15284 73268
rect 15244 72388 15284 72428
rect 15244 66760 15284 66800
rect 15532 71212 15572 71252
rect 15436 71128 15476 71168
rect 15244 64324 15284 64364
rect 15244 63652 15284 63692
rect 15436 65248 15476 65288
rect 15244 62644 15284 62684
rect 15820 76000 15860 76040
rect 16204 79192 16244 79232
rect 16108 78016 16148 78056
rect 16300 78940 16340 78980
rect 16300 78520 16340 78560
rect 17356 93640 17396 93680
rect 16492 82048 16532 82088
rect 16492 79864 16532 79904
rect 16492 79612 16532 79652
rect 16876 84820 16916 84860
rect 16780 82048 16820 82088
rect 16588 78100 16628 78140
rect 16684 81796 16724 81836
rect 16780 80620 16820 80660
rect 16108 74656 16148 74696
rect 16108 74488 16148 74528
rect 15916 72892 15956 72932
rect 15724 71716 15764 71756
rect 15724 70540 15764 70580
rect 15724 66256 15764 66296
rect 15820 66172 15860 66212
rect 15532 63148 15572 63188
rect 15244 62392 15284 62432
rect 15532 62392 15572 62432
rect 15436 59116 15476 59156
rect 15436 56260 15476 56300
rect 15244 53236 15284 53276
rect 15244 52144 15284 52184
rect 15244 43240 15284 43280
rect 15724 64660 15764 64700
rect 16204 73480 16244 73520
rect 16012 70792 16052 70832
rect 16396 74488 16436 74528
rect 16396 73900 16436 73940
rect 16396 71548 16436 71588
rect 16300 70456 16340 70496
rect 16396 71296 16436 71336
rect 16588 70540 16628 70580
rect 16684 71128 16724 71168
rect 16588 70372 16628 70412
rect 16588 69280 16628 69320
rect 16012 63568 16052 63608
rect 15916 62392 15956 62432
rect 15724 61804 15764 61844
rect 15916 60208 15956 60248
rect 16012 61636 16052 61676
rect 15916 60040 15956 60080
rect 15916 59788 15956 59828
rect 16012 59284 16052 59324
rect 15916 58360 15956 58400
rect 15628 53236 15668 53276
rect 15820 53992 15860 54032
rect 16684 67432 16724 67472
rect 16492 65752 16532 65792
rect 16396 65080 16436 65120
rect 16396 62392 16436 62432
rect 16492 63820 16532 63860
rect 16204 60208 16244 60248
rect 16108 58360 16148 58400
rect 16108 58192 16148 58232
rect 16012 53320 16052 53360
rect 15244 42988 15284 43028
rect 15244 41812 15284 41852
rect 15244 35596 15284 35636
rect 15244 34420 15284 34460
rect 15148 27448 15188 27488
rect 14572 17620 14612 17660
rect 14668 17704 14708 17744
rect 14476 16948 14516 16988
rect 14668 16948 14708 16988
rect 14668 16696 14708 16736
rect 14476 14596 14516 14636
rect 14188 11488 14228 11528
rect 14380 12412 14420 12452
rect 14668 14596 14708 14636
rect 14860 17788 14900 17828
rect 14860 16696 14900 16736
rect 15052 19384 15092 19424
rect 14476 11488 14516 11528
rect 14284 9556 14324 9596
rect 14188 8548 14228 8588
rect 14380 9304 14420 9344
rect 14284 5692 14324 5732
rect 14188 4852 14228 4892
rect 13996 2836 14036 2876
rect 14572 10060 14612 10100
rect 13420 1912 13460 1952
rect 14956 15352 14996 15392
rect 15436 42484 15476 42524
rect 15436 40972 15476 41012
rect 15436 39964 15476 40004
rect 15436 38032 15476 38072
rect 15436 35932 15476 35972
rect 15628 47188 15668 47228
rect 15628 44164 15668 44204
rect 15628 41896 15668 41936
rect 15628 38872 15668 38912
rect 15820 48700 15860 48740
rect 16204 53992 16244 54032
rect 17356 89524 17396 89564
rect 17164 83560 17204 83600
rect 17260 83812 17300 83852
rect 17068 83476 17108 83516
rect 17164 83392 17204 83432
rect 16972 82132 17012 82172
rect 16972 78436 17012 78476
rect 17260 83056 17300 83096
rect 17452 87424 17492 87464
rect 17452 85912 17492 85952
rect 18028 95572 18068 95612
rect 18220 94816 18260 94856
rect 18124 94144 18164 94184
rect 17740 93892 17780 93932
rect 18412 94816 18452 94856
rect 18604 94144 18644 94184
rect 18796 94816 18836 94856
rect 19084 94816 19124 94856
rect 20048 95236 20088 95276
rect 20130 95236 20170 95276
rect 20212 95236 20252 95276
rect 20294 95236 20334 95276
rect 20376 95236 20416 95276
rect 19468 94816 19508 94856
rect 18808 94480 18848 94520
rect 18890 94480 18930 94520
rect 18972 94480 19012 94520
rect 19054 94480 19094 94520
rect 19136 94480 19176 94520
rect 19084 94228 19124 94268
rect 18988 94144 19028 94184
rect 18988 93304 19028 93344
rect 18700 93136 18740 93176
rect 18808 92968 18848 93008
rect 18890 92968 18930 93008
rect 18972 92968 19012 93008
rect 19054 92968 19094 93008
rect 19136 92968 19176 93008
rect 19564 94228 19604 94268
rect 19756 94060 19796 94100
rect 19852 94144 19892 94184
rect 19468 92632 19508 92672
rect 19756 92632 19796 92672
rect 19756 91792 19796 91832
rect 17644 89524 17684 89564
rect 17740 86500 17780 86540
rect 17836 85744 17876 85784
rect 17740 84064 17780 84104
rect 17836 83980 17876 84020
rect 17644 83560 17684 83600
rect 17548 80536 17588 80576
rect 17068 75916 17108 75956
rect 16876 69028 16916 69068
rect 17356 75916 17396 75956
rect 17164 73480 17204 73520
rect 17164 71548 17204 71588
rect 17260 71464 17300 71504
rect 16876 68860 16916 68900
rect 16876 66844 16916 66884
rect 16780 64828 16820 64868
rect 16684 62392 16724 62432
rect 16684 58192 16724 58232
rect 16684 57772 16724 57812
rect 17164 70372 17204 70412
rect 17068 69196 17108 69236
rect 17068 69028 17108 69068
rect 17260 67432 17300 67472
rect 17068 64576 17108 64616
rect 17164 66844 17204 66884
rect 16876 62056 16916 62096
rect 16972 64492 17012 64532
rect 17068 62980 17108 63020
rect 17068 61804 17108 61844
rect 16972 60040 17012 60080
rect 17068 61552 17108 61592
rect 16972 57604 17012 57644
rect 17932 82720 17972 82760
rect 18220 88096 18260 88136
rect 18808 91456 18848 91496
rect 18890 91456 18930 91496
rect 18972 91456 19012 91496
rect 19054 91456 19094 91496
rect 19136 91456 19176 91496
rect 18808 89944 18848 89984
rect 18890 89944 18930 89984
rect 18972 89944 19012 89984
rect 19054 89944 19094 89984
rect 19136 89944 19176 89984
rect 18988 88852 19028 88892
rect 18604 88768 18644 88808
rect 18124 84400 18164 84440
rect 17932 81208 17972 81248
rect 17644 78016 17684 78056
rect 17548 77680 17588 77720
rect 18604 86920 18644 86960
rect 18808 88432 18848 88472
rect 18890 88432 18930 88472
rect 18972 88432 19012 88472
rect 19054 88432 19094 88472
rect 19136 88432 19176 88472
rect 19372 88684 19412 88724
rect 18796 87088 18836 87128
rect 18808 86920 18848 86960
rect 18890 86920 18930 86960
rect 18972 86920 19012 86960
rect 19054 86920 19094 86960
rect 19136 86920 19176 86960
rect 18796 86416 18836 86456
rect 18316 82720 18356 82760
rect 18316 81796 18356 81836
rect 17932 78604 17972 78644
rect 18028 78352 18068 78392
rect 17644 77428 17684 77468
rect 17548 75748 17588 75788
rect 17836 74488 17876 74528
rect 18316 81292 18356 81332
rect 18220 79108 18260 79148
rect 17548 72724 17588 72764
rect 17644 72052 17684 72092
rect 17548 70876 17588 70916
rect 17452 67936 17492 67976
rect 17260 65080 17300 65120
rect 17356 66508 17396 66548
rect 17356 64996 17396 65036
rect 17260 62476 17300 62516
rect 17260 62056 17300 62096
rect 17356 61468 17396 61508
rect 17260 60544 17300 60584
rect 17068 56176 17108 56216
rect 16396 50296 16436 50336
rect 16204 49624 16244 49664
rect 16300 48952 16340 48992
rect 16204 48028 16244 48068
rect 16396 48868 16436 48908
rect 16780 51052 16820 51092
rect 17260 58528 17300 58568
rect 17836 71212 17876 71252
rect 18028 72556 18068 72596
rect 18028 71212 18068 71252
rect 17932 70540 17972 70580
rect 17740 67936 17780 67976
rect 17740 66508 17780 66548
rect 18508 84232 18548 84272
rect 18808 85408 18848 85448
rect 18890 85408 18930 85448
rect 18972 85408 19012 85448
rect 19054 85408 19094 85448
rect 19136 85408 19176 85448
rect 18796 84064 18836 84104
rect 18808 83896 18848 83936
rect 18890 83896 18930 83936
rect 18972 83896 19012 83936
rect 19054 83896 19094 83936
rect 19136 83896 19176 83936
rect 18796 83728 18836 83768
rect 18988 83560 19028 83600
rect 18604 81292 18644 81332
rect 18604 76672 18644 76712
rect 18508 74992 18548 75032
rect 18316 72640 18356 72680
rect 18604 73312 18644 73352
rect 18508 72388 18548 72428
rect 18028 66256 18068 66296
rect 17548 60124 17588 60164
rect 17644 65080 17684 65120
rect 17452 60040 17492 60080
rect 17740 64996 17780 65036
rect 18508 71632 18548 71672
rect 18604 72052 18644 72092
rect 18508 70708 18548 70748
rect 18412 67096 18452 67136
rect 18220 63988 18260 64028
rect 18124 63400 18164 63440
rect 18124 63232 18164 63272
rect 18508 64072 18548 64112
rect 18412 63652 18452 63692
rect 18316 63316 18356 63356
rect 17836 61468 17876 61508
rect 17932 60460 17972 60500
rect 17740 60040 17780 60080
rect 17740 56344 17780 56384
rect 15820 42904 15860 42944
rect 15820 42484 15860 42524
rect 15820 42064 15860 42104
rect 15820 41812 15860 41852
rect 15820 41476 15860 41516
rect 16012 42652 16052 42692
rect 16108 41896 16148 41936
rect 15916 40972 15956 41012
rect 15820 40468 15860 40508
rect 15724 38368 15764 38408
rect 16300 41980 16340 42020
rect 16396 42652 16436 42692
rect 15916 36604 15956 36644
rect 15820 35596 15860 35636
rect 15436 29968 15476 30008
rect 15532 31312 15572 31352
rect 15436 29632 15476 29672
rect 15916 35512 15956 35552
rect 15916 35092 15956 35132
rect 15916 34504 15956 34544
rect 15916 33496 15956 33536
rect 15916 31984 15956 32024
rect 15820 29884 15860 29924
rect 15724 29128 15764 29168
rect 15916 29464 15956 29504
rect 15340 27448 15380 27488
rect 15436 26188 15476 26228
rect 15340 25264 15380 25304
rect 15244 21736 15284 21776
rect 15340 21568 15380 21608
rect 15244 21316 15284 21356
rect 15340 20728 15380 20768
rect 15244 20140 15284 20180
rect 15340 19720 15380 19760
rect 15436 19384 15476 19424
rect 15340 18460 15380 18500
rect 15340 17956 15380 17996
rect 15148 14764 15188 14804
rect 15436 14764 15476 14804
rect 15436 13420 15476 13460
rect 15340 9640 15380 9680
rect 15052 5692 15092 5732
rect 14668 5608 14708 5648
rect 14764 2584 14804 2624
rect 15724 28792 15764 28832
rect 15820 28876 15860 28916
rect 15724 27112 15764 27152
rect 15724 26860 15764 26900
rect 15724 24004 15764 24044
rect 15820 21316 15860 21356
rect 15820 21064 15860 21104
rect 15820 20140 15860 20180
rect 15628 17956 15668 17996
rect 15724 18544 15764 18584
rect 15628 17620 15668 17660
rect 15628 14764 15668 14804
rect 15628 9220 15668 9260
rect 15340 1912 15380 1952
rect 15820 17788 15860 17828
rect 16108 36688 16148 36728
rect 16300 38872 16340 38912
rect 16300 36520 16340 36560
rect 16300 35932 16340 35972
rect 16300 35176 16340 35216
rect 16300 31564 16340 31604
rect 16108 30220 16148 30260
rect 16204 31060 16244 31100
rect 16108 29128 16148 29168
rect 16588 41980 16628 42020
rect 16492 41644 16532 41684
rect 16492 41056 16532 41096
rect 16492 40804 16532 40844
rect 16492 38200 16532 38240
rect 16396 30976 16436 31016
rect 16396 30808 16436 30848
rect 16300 29296 16340 29336
rect 16204 27616 16244 27656
rect 16300 28036 16340 28076
rect 16108 23248 16148 23288
rect 16204 25264 16244 25304
rect 16012 21484 16052 21524
rect 16396 27532 16436 27572
rect 16684 41728 16724 41768
rect 16876 39040 16916 39080
rect 16684 38200 16724 38240
rect 16684 36940 16724 36980
rect 16588 36856 16628 36896
rect 16876 36940 16916 36980
rect 16780 35596 16820 35636
rect 16588 35092 16628 35132
rect 16588 33496 16628 33536
rect 16588 31144 16628 31184
rect 16588 30808 16628 30848
rect 16780 31396 16820 31436
rect 16684 28876 16724 28916
rect 16588 27028 16628 27068
rect 16492 26860 16532 26900
rect 16492 26104 16532 26144
rect 16588 26020 16628 26060
rect 17452 53320 17492 53360
rect 18124 60124 18164 60164
rect 18028 58444 18068 58484
rect 18412 60040 18452 60080
rect 18316 59872 18356 59912
rect 18316 59704 18356 59744
rect 18220 58360 18260 58400
rect 18220 57856 18260 57896
rect 18220 56176 18260 56216
rect 18412 57856 18452 57896
rect 18316 56092 18356 56132
rect 18316 53572 18356 53612
rect 18508 53992 18548 54032
rect 18604 51892 18644 51932
rect 17644 49288 17684 49328
rect 18220 48448 18260 48488
rect 18604 48364 18644 48404
rect 17260 43996 17300 44036
rect 17164 39964 17204 40004
rect 17260 40804 17300 40844
rect 17068 39628 17108 39668
rect 17356 37360 17396 37400
rect 17260 37108 17300 37148
rect 17356 37024 17396 37064
rect 17164 35596 17204 35636
rect 17068 34420 17108 34460
rect 17260 35176 17300 35216
rect 17548 41392 17588 41432
rect 17548 39628 17588 39668
rect 17548 36352 17588 36392
rect 17836 37528 17876 37568
rect 17740 37024 17780 37064
rect 17452 35092 17492 35132
rect 17356 33496 17396 33536
rect 17452 34168 17492 34208
rect 17740 35764 17780 35804
rect 17740 34084 17780 34124
rect 18124 40384 18164 40424
rect 18124 39712 18164 39752
rect 18028 36856 18068 36896
rect 18124 36688 18164 36728
rect 18028 36352 18068 36392
rect 19084 83392 19124 83432
rect 18808 82384 18848 82424
rect 18890 82384 18930 82424
rect 18972 82384 19012 82424
rect 19054 82384 19094 82424
rect 19136 82384 19176 82424
rect 18988 82216 19028 82256
rect 19084 81460 19124 81500
rect 18808 80872 18848 80912
rect 18890 80872 18930 80912
rect 18972 80872 19012 80912
rect 19054 80872 19094 80912
rect 19136 80872 19176 80912
rect 18796 79528 18836 79568
rect 19084 80704 19124 80744
rect 19084 79612 19124 79652
rect 18988 79528 19028 79568
rect 18808 79360 18848 79400
rect 18890 79360 18930 79400
rect 18972 79360 19012 79400
rect 19054 79360 19094 79400
rect 19136 79360 19176 79400
rect 18796 79192 18836 79232
rect 19084 79108 19124 79148
rect 18892 78604 18932 78644
rect 18796 78016 18836 78056
rect 19084 78520 19124 78560
rect 19180 78268 19220 78308
rect 19372 84148 19412 84188
rect 19372 83896 19412 83936
rect 19372 82552 19412 82592
rect 19372 82384 19412 82424
rect 19276 78016 19316 78056
rect 19372 78352 19412 78392
rect 18808 77848 18848 77888
rect 18890 77848 18930 77888
rect 18972 77848 19012 77888
rect 19054 77848 19094 77888
rect 19136 77848 19176 77888
rect 18808 76336 18848 76376
rect 18890 76336 18930 76376
rect 18972 76336 19012 76376
rect 19054 76336 19094 76376
rect 19136 76336 19176 76376
rect 18796 74992 18836 75032
rect 18808 74824 18848 74864
rect 18890 74824 18930 74864
rect 18972 74824 19012 74864
rect 19054 74824 19094 74864
rect 19136 74824 19176 74864
rect 18988 74656 19028 74696
rect 19084 74572 19124 74612
rect 19372 74656 19412 74696
rect 19564 83812 19604 83852
rect 19564 82384 19604 82424
rect 19756 89608 19796 89648
rect 20236 94144 20276 94184
rect 20048 93724 20088 93764
rect 20130 93724 20170 93764
rect 20212 93724 20252 93764
rect 20294 93724 20334 93764
rect 20376 93724 20416 93764
rect 19948 93304 19988 93344
rect 20140 93304 20180 93344
rect 20048 92212 20088 92252
rect 20130 92212 20170 92252
rect 20212 92212 20252 92252
rect 20294 92212 20334 92252
rect 20376 92212 20416 92252
rect 20140 91120 20180 91160
rect 20048 90700 20088 90740
rect 20130 90700 20170 90740
rect 20212 90700 20252 90740
rect 20294 90700 20334 90740
rect 20376 90700 20416 90740
rect 20140 90280 20180 90320
rect 20140 89608 20180 89648
rect 20048 89188 20088 89228
rect 20130 89188 20170 89228
rect 20212 89188 20252 89228
rect 20294 89188 20334 89228
rect 20376 89188 20416 89228
rect 19852 88012 19892 88052
rect 19756 87928 19796 87968
rect 19756 87256 19796 87296
rect 19564 78016 19604 78056
rect 18988 73480 19028 73520
rect 19180 73480 19220 73520
rect 18808 73312 18848 73352
rect 18890 73312 18930 73352
rect 18972 73312 19012 73352
rect 19054 73312 19094 73352
rect 19136 73312 19176 73352
rect 18796 72052 18836 72092
rect 19084 72724 19124 72764
rect 18808 71800 18848 71840
rect 18890 71800 18930 71840
rect 18972 71800 19012 71840
rect 19054 71800 19094 71840
rect 19136 71800 19176 71840
rect 18892 71632 18932 71672
rect 18892 70456 18932 70496
rect 18808 70288 18848 70328
rect 18890 70288 18930 70328
rect 18972 70288 19012 70328
rect 19054 70288 19094 70328
rect 19136 70288 19176 70328
rect 19084 70120 19124 70160
rect 19276 70036 19316 70076
rect 19084 68944 19124 68984
rect 18808 68776 18848 68816
rect 18890 68776 18930 68816
rect 18972 68776 19012 68816
rect 19054 68776 19094 68816
rect 19136 68776 19176 68816
rect 18796 68608 18836 68648
rect 19276 68440 19316 68480
rect 18808 67264 18848 67304
rect 18890 67264 18930 67304
rect 18972 67264 19012 67304
rect 19054 67264 19094 67304
rect 19136 67264 19176 67304
rect 18796 67096 18836 67136
rect 19180 66088 19220 66128
rect 18808 65752 18848 65792
rect 18890 65752 18930 65792
rect 18972 65752 19012 65792
rect 19054 65752 19094 65792
rect 19136 65752 19176 65792
rect 19084 64996 19124 65036
rect 18808 64240 18848 64280
rect 18890 64240 18930 64280
rect 18972 64240 19012 64280
rect 19054 64240 19094 64280
rect 19136 64240 19176 64280
rect 18988 63820 19028 63860
rect 19372 63400 19412 63440
rect 19660 73900 19700 73940
rect 20332 88600 20372 88640
rect 20140 87844 20180 87884
rect 20048 87676 20088 87716
rect 20130 87676 20170 87716
rect 20212 87676 20252 87716
rect 20294 87676 20334 87716
rect 20376 87676 20416 87716
rect 20140 87256 20180 87296
rect 20140 86584 20180 86624
rect 20524 87424 20564 87464
rect 20048 86164 20088 86204
rect 20130 86164 20170 86204
rect 20212 86164 20252 86204
rect 20294 86164 20334 86204
rect 20376 86164 20416 86204
rect 20048 84652 20088 84692
rect 20130 84652 20170 84692
rect 20212 84652 20252 84692
rect 20294 84652 20334 84692
rect 20376 84652 20416 84692
rect 20140 84232 20180 84272
rect 19948 83476 19988 83516
rect 20140 83560 20180 83600
rect 20048 83140 20088 83180
rect 20130 83140 20170 83180
rect 20212 83140 20252 83180
rect 20294 83140 20334 83180
rect 20376 83140 20416 83180
rect 20044 82972 20084 83012
rect 20044 81796 20084 81836
rect 20048 81628 20088 81668
rect 20130 81628 20170 81668
rect 20212 81628 20252 81668
rect 20294 81628 20334 81668
rect 20376 81628 20416 81668
rect 20044 81376 20084 81416
rect 20048 80116 20088 80156
rect 20130 80116 20170 80156
rect 20212 80116 20252 80156
rect 20294 80116 20334 80156
rect 20376 80116 20416 80156
rect 20428 78772 20468 78812
rect 20048 78604 20088 78644
rect 20130 78604 20170 78644
rect 20212 78604 20252 78644
rect 20294 78604 20334 78644
rect 20376 78604 20416 78644
rect 20044 78352 20084 78392
rect 20044 78100 20084 78140
rect 20048 77092 20088 77132
rect 20130 77092 20170 77132
rect 20212 77092 20252 77132
rect 20294 77092 20334 77132
rect 20376 77092 20416 77132
rect 20140 76756 20180 76796
rect 20140 76588 20180 76628
rect 19660 72808 19700 72848
rect 20140 76000 20180 76040
rect 20428 75748 20468 75788
rect 20048 75580 20088 75620
rect 20130 75580 20170 75620
rect 20212 75580 20252 75620
rect 20294 75580 20334 75620
rect 20376 75580 20416 75620
rect 20428 75412 20468 75452
rect 19852 72892 19892 72932
rect 20428 74236 20468 74276
rect 19852 72724 19892 72764
rect 20048 74068 20088 74108
rect 20130 74068 20170 74108
rect 20212 74068 20252 74108
rect 20294 74068 20334 74108
rect 20376 74068 20416 74108
rect 20044 73900 20084 73940
rect 20428 73900 20468 73940
rect 20428 72808 20468 72848
rect 20044 72724 20084 72764
rect 20048 72556 20088 72596
rect 20130 72556 20170 72596
rect 20212 72556 20252 72596
rect 20294 72556 20334 72596
rect 20376 72556 20416 72596
rect 20044 72388 20084 72428
rect 19948 71548 19988 71588
rect 20048 71044 20088 71084
rect 20130 71044 20170 71084
rect 20212 71044 20252 71084
rect 20294 71044 20334 71084
rect 20376 71044 20416 71084
rect 19756 69952 19796 69992
rect 19756 68608 19796 68648
rect 18988 62980 19028 63020
rect 19276 62812 19316 62852
rect 18808 62728 18848 62768
rect 18890 62728 18930 62768
rect 18972 62728 19012 62768
rect 19054 62728 19094 62768
rect 19136 62728 19176 62768
rect 19180 62560 19220 62600
rect 18988 61552 19028 61592
rect 19180 61468 19220 61508
rect 18808 61216 18848 61256
rect 18890 61216 18930 61256
rect 18972 61216 19012 61256
rect 19054 61216 19094 61256
rect 19136 61216 19176 61256
rect 18808 59704 18848 59744
rect 18890 59704 18930 59744
rect 18972 59704 19012 59744
rect 19054 59704 19094 59744
rect 19136 59704 19176 59744
rect 18796 58444 18836 58484
rect 18808 58192 18848 58232
rect 18890 58192 18930 58232
rect 18972 58192 19012 58232
rect 19054 58192 19094 58232
rect 19136 58192 19176 58232
rect 18892 57772 18932 57812
rect 18808 56680 18848 56720
rect 18890 56680 18930 56720
rect 18972 56680 19012 56720
rect 19054 56680 19094 56720
rect 19136 56680 19176 56720
rect 19180 56344 19220 56384
rect 18796 55336 18836 55376
rect 18808 55168 18848 55208
rect 18890 55168 18930 55208
rect 18972 55168 19012 55208
rect 19054 55168 19094 55208
rect 19136 55168 19176 55208
rect 18796 55000 18836 55040
rect 18892 53992 18932 54032
rect 18808 53656 18848 53696
rect 18890 53656 18930 53696
rect 18972 53656 19012 53696
rect 19054 53656 19094 53696
rect 19136 53656 19176 53696
rect 18808 52144 18848 52184
rect 18890 52144 18930 52184
rect 18972 52144 19012 52184
rect 19054 52144 19094 52184
rect 19136 52144 19176 52184
rect 18808 50632 18848 50672
rect 18890 50632 18930 50672
rect 18972 50632 19012 50672
rect 19054 50632 19094 50672
rect 19136 50632 19176 50672
rect 19180 50212 19220 50252
rect 18808 49120 18848 49160
rect 18890 49120 18930 49160
rect 18972 49120 19012 49160
rect 19054 49120 19094 49160
rect 19136 49120 19176 49160
rect 19756 66088 19796 66128
rect 19756 63484 19796 63524
rect 19852 63400 19892 63440
rect 19468 61468 19508 61508
rect 19468 59284 19508 59324
rect 19660 61888 19700 61928
rect 19372 58444 19412 58484
rect 19564 58444 19604 58484
rect 19468 57688 19508 57728
rect 19468 54244 19508 54284
rect 19372 53572 19412 53612
rect 19468 53236 19508 53276
rect 19372 50968 19412 51008
rect 19372 49624 19412 49664
rect 19372 49456 19412 49496
rect 19372 48784 19412 48824
rect 18808 47608 18848 47648
rect 18890 47608 18930 47648
rect 18972 47608 19012 47648
rect 19054 47608 19094 47648
rect 19136 47608 19176 47648
rect 18808 46096 18848 46136
rect 18890 46096 18930 46136
rect 18972 46096 19012 46136
rect 19054 46096 19094 46136
rect 19136 46096 19176 46136
rect 18892 45172 18932 45212
rect 18808 44584 18848 44624
rect 18890 44584 18930 44624
rect 18972 44584 19012 44624
rect 19054 44584 19094 44624
rect 19136 44584 19176 44624
rect 18604 42064 18644 42104
rect 18796 43240 18836 43280
rect 18808 43072 18848 43112
rect 18890 43072 18930 43112
rect 18972 43072 19012 43112
rect 19054 43072 19094 43112
rect 19136 43072 19176 43112
rect 18796 42904 18836 42944
rect 18808 41560 18848 41600
rect 18890 41560 18930 41600
rect 18972 41560 19012 41600
rect 19054 41560 19094 41600
rect 19136 41560 19176 41600
rect 18508 39880 18548 39920
rect 18412 38872 18452 38912
rect 18316 35764 18356 35804
rect 17932 34672 17972 34712
rect 18124 34672 18164 34712
rect 17260 30892 17300 30932
rect 17068 30304 17108 30344
rect 17260 29884 17300 29924
rect 16876 28036 16916 28076
rect 17260 29044 17300 29084
rect 16876 26020 16916 26060
rect 16588 24844 16628 24884
rect 16684 24592 16724 24632
rect 16396 23752 16436 23792
rect 16396 23416 16436 23456
rect 16204 20812 16244 20852
rect 15916 17620 15956 17660
rect 15820 11320 15860 11360
rect 16012 14176 16052 14216
rect 16204 14176 16244 14216
rect 15916 8716 15956 8756
rect 16972 24676 17012 24716
rect 16684 22912 16724 22952
rect 16492 21232 16532 21272
rect 16492 20896 16532 20936
rect 16492 19048 16532 19088
rect 16588 18628 16628 18668
rect 16492 17620 16532 17660
rect 16492 15436 16532 15476
rect 16396 13756 16436 13796
rect 16876 16528 16916 16568
rect 17260 26104 17300 26144
rect 17260 24592 17300 24632
rect 17260 23584 17300 23624
rect 17260 17200 17300 17240
rect 17452 29968 17492 30008
rect 17452 23164 17492 23204
rect 17452 22492 17492 22532
rect 16588 13168 16628 13208
rect 16300 8128 16340 8168
rect 16492 8716 16532 8756
rect 16396 4852 16436 4892
rect 16972 13756 17012 13796
rect 16972 13000 17012 13040
rect 17260 16108 17300 16148
rect 17260 14764 17300 14804
rect 17356 12664 17396 12704
rect 17452 12328 17492 12368
rect 17356 10228 17396 10268
rect 17740 33748 17780 33788
rect 17836 33496 17876 33536
rect 18412 35092 18452 35132
rect 18220 33160 18260 33200
rect 18124 33076 18164 33116
rect 18220 32908 18260 32948
rect 17932 32740 17972 32780
rect 18028 32824 18068 32864
rect 17932 32152 17972 32192
rect 17740 26608 17780 26648
rect 17644 25012 17684 25052
rect 17836 25012 17876 25052
rect 17932 28960 17972 29000
rect 18124 32488 18164 32528
rect 18220 30724 18260 30764
rect 17836 23416 17876 23456
rect 17836 22576 17876 22616
rect 17740 22492 17780 22532
rect 17740 19888 17780 19928
rect 18220 27532 18260 27572
rect 18220 26692 18260 26732
rect 18808 40048 18848 40088
rect 18890 40048 18930 40088
rect 18972 40048 19012 40088
rect 19054 40048 19094 40088
rect 19136 40048 19176 40088
rect 18892 39796 18932 39836
rect 18808 38536 18848 38576
rect 18890 38536 18930 38576
rect 18972 38536 19012 38576
rect 19054 38536 19094 38576
rect 19136 38536 19176 38576
rect 19180 38368 19220 38408
rect 18892 37528 18932 37568
rect 19180 37192 19220 37232
rect 18808 37024 18848 37064
rect 18890 37024 18930 37064
rect 18972 37024 19012 37064
rect 19054 37024 19094 37064
rect 19136 37024 19176 37064
rect 18892 36856 18932 36896
rect 19180 36856 19220 36896
rect 19084 36436 19124 36476
rect 18604 35932 18644 35972
rect 18508 31396 18548 31436
rect 18412 29044 18452 29084
rect 18412 28204 18452 28244
rect 18124 23500 18164 23540
rect 18220 23332 18260 23372
rect 18124 21484 18164 21524
rect 18028 21064 18068 21104
rect 17836 18124 17876 18164
rect 18028 17956 18068 17996
rect 17932 17872 17972 17912
rect 17836 16444 17876 16484
rect 17836 10228 17876 10268
rect 17356 4096 17396 4136
rect 18028 17788 18068 17828
rect 19180 36016 19220 36056
rect 18796 35680 18836 35720
rect 18808 35512 18848 35552
rect 18890 35512 18930 35552
rect 18972 35512 19012 35552
rect 19054 35512 19094 35552
rect 19136 35512 19176 35552
rect 18796 35344 18836 35384
rect 18700 34252 18740 34292
rect 19180 35344 19220 35384
rect 18892 35176 18932 35216
rect 18892 34588 18932 34628
rect 18988 34504 19028 34544
rect 18796 34168 18836 34208
rect 18808 34000 18848 34040
rect 18890 34000 18930 34040
rect 18972 34000 19012 34040
rect 19054 34000 19094 34040
rect 19136 34000 19176 34040
rect 18700 32992 18740 33032
rect 19276 33664 19316 33704
rect 18988 33496 19028 33536
rect 18988 33076 19028 33116
rect 18892 32656 18932 32696
rect 18808 32488 18848 32528
rect 18890 32488 18930 32528
rect 18972 32488 19012 32528
rect 19054 32488 19094 32528
rect 19136 32488 19176 32528
rect 18796 32320 18836 32360
rect 19180 32320 19220 32360
rect 19084 31984 19124 32024
rect 19180 31144 19220 31184
rect 18808 30976 18848 31016
rect 18890 30976 18930 31016
rect 18972 30976 19012 31016
rect 19054 30976 19094 31016
rect 19136 30976 19176 31016
rect 18796 30808 18836 30848
rect 19180 30808 19220 30848
rect 19084 30472 19124 30512
rect 18700 30220 18740 30260
rect 18988 30388 19028 30428
rect 18604 28204 18644 28244
rect 18604 27532 18644 27572
rect 18412 23332 18452 23372
rect 18988 29968 19028 30008
rect 19084 29716 19124 29756
rect 19660 55504 19700 55544
rect 19660 55336 19700 55376
rect 19660 53236 19700 53276
rect 19852 57688 19892 57728
rect 20332 69784 20372 69824
rect 20140 69700 20180 69740
rect 20428 69700 20468 69740
rect 20048 69532 20088 69572
rect 20130 69532 20170 69572
rect 20212 69532 20252 69572
rect 20294 69532 20334 69572
rect 20376 69532 20416 69572
rect 20048 68020 20088 68060
rect 20130 68020 20170 68060
rect 20212 68020 20252 68060
rect 20294 68020 20334 68060
rect 20376 68020 20416 68060
rect 20428 67852 20468 67892
rect 20140 66676 20180 66716
rect 20048 66508 20088 66548
rect 20130 66508 20170 66548
rect 20212 66508 20252 66548
rect 20294 66508 20334 66548
rect 20376 66508 20416 66548
rect 20048 64996 20088 65036
rect 20130 64996 20170 65036
rect 20212 64996 20252 65036
rect 20294 64996 20334 65036
rect 20376 64996 20416 65036
rect 20140 64576 20180 64616
rect 20044 64156 20084 64196
rect 20048 63484 20088 63524
rect 20130 63484 20170 63524
rect 20212 63484 20252 63524
rect 20294 63484 20334 63524
rect 20376 63484 20416 63524
rect 20044 62224 20084 62264
rect 20236 62140 20276 62180
rect 20048 61972 20088 62012
rect 20130 61972 20170 62012
rect 20212 61972 20252 62012
rect 20294 61972 20334 62012
rect 20376 61972 20416 62012
rect 20428 61720 20468 61760
rect 20428 61048 20468 61088
rect 20048 60460 20088 60500
rect 20130 60460 20170 60500
rect 20212 60460 20252 60500
rect 20294 60460 20334 60500
rect 20376 60460 20416 60500
rect 20048 58948 20088 58988
rect 20130 58948 20170 58988
rect 20212 58948 20252 58988
rect 20294 58948 20334 58988
rect 20376 58948 20416 58988
rect 20044 58780 20084 58820
rect 20044 57772 20084 57812
rect 20048 57436 20088 57476
rect 20130 57436 20170 57476
rect 20212 57436 20252 57476
rect 20294 57436 20334 57476
rect 20376 57436 20416 57476
rect 20048 55924 20088 55964
rect 20130 55924 20170 55964
rect 20212 55924 20252 55964
rect 20294 55924 20334 55964
rect 20376 55924 20416 55964
rect 19948 55336 19988 55376
rect 19756 50128 19796 50168
rect 19660 49624 19700 49664
rect 19660 47440 19700 47480
rect 19564 47104 19604 47144
rect 19564 38536 19604 38576
rect 20048 54412 20088 54452
rect 20130 54412 20170 54452
rect 20212 54412 20252 54452
rect 20294 54412 20334 54452
rect 20376 54412 20416 54452
rect 20044 54244 20084 54284
rect 20908 87424 20948 87464
rect 20716 85072 20756 85112
rect 20812 84904 20852 84944
rect 20908 84568 20948 84608
rect 20812 78772 20852 78812
rect 21196 85408 21236 85448
rect 20908 75916 20948 75956
rect 20716 68104 20756 68144
rect 20812 68776 20852 68816
rect 21484 87424 21524 87464
rect 21196 76672 21236 76712
rect 21388 76756 21428 76796
rect 21196 73396 21236 73436
rect 21100 72808 21140 72848
rect 20620 62476 20660 62516
rect 20620 62308 20660 62348
rect 21004 68104 21044 68144
rect 20812 63064 20852 63104
rect 20908 62308 20948 62348
rect 21100 63064 21140 63104
rect 21196 62476 21236 62516
rect 21004 61216 21044 61256
rect 21004 61048 21044 61088
rect 21196 61384 21236 61424
rect 21196 61132 21236 61172
rect 20048 52900 20088 52940
rect 20130 52900 20170 52940
rect 20212 52900 20252 52940
rect 20294 52900 20334 52940
rect 20376 52900 20416 52940
rect 20140 52480 20180 52520
rect 20140 51808 20180 51848
rect 20048 51388 20088 51428
rect 20130 51388 20170 51428
rect 20212 51388 20252 51428
rect 20294 51388 20334 51428
rect 20376 51388 20416 51428
rect 20048 49876 20088 49916
rect 20130 49876 20170 49916
rect 20212 49876 20252 49916
rect 20294 49876 20334 49916
rect 20376 49876 20416 49916
rect 20048 48364 20088 48404
rect 20130 48364 20170 48404
rect 20212 48364 20252 48404
rect 20294 48364 20334 48404
rect 20376 48364 20416 48404
rect 20140 47944 20180 47984
rect 20048 46852 20088 46892
rect 20130 46852 20170 46892
rect 20212 46852 20252 46892
rect 20294 46852 20334 46892
rect 20376 46852 20416 46892
rect 20140 46432 20180 46472
rect 21388 61216 21428 61256
rect 20048 45340 20088 45380
rect 20130 45340 20170 45380
rect 20212 45340 20252 45380
rect 20294 45340 20334 45380
rect 20376 45340 20416 45380
rect 20048 43828 20088 43868
rect 20130 43828 20170 43868
rect 20212 43828 20252 43868
rect 20294 43828 20334 43868
rect 20376 43828 20416 43868
rect 20620 43240 20660 43280
rect 19564 35428 19604 35468
rect 19468 34252 19508 34292
rect 19468 34084 19508 34124
rect 19660 33580 19700 33620
rect 20048 42316 20088 42356
rect 20130 42316 20170 42356
rect 20212 42316 20252 42356
rect 20294 42316 20334 42356
rect 20376 42316 20416 42356
rect 20048 40804 20088 40844
rect 20130 40804 20170 40844
rect 20212 40804 20252 40844
rect 20294 40804 20334 40844
rect 20376 40804 20416 40844
rect 20048 39292 20088 39332
rect 20130 39292 20170 39332
rect 20212 39292 20252 39332
rect 20294 39292 20334 39332
rect 20376 39292 20416 39332
rect 20044 37948 20084 37988
rect 20428 37948 20468 37988
rect 20048 37780 20088 37820
rect 20130 37780 20170 37820
rect 20212 37780 20252 37820
rect 20294 37780 20334 37820
rect 20376 37780 20416 37820
rect 20044 37612 20084 37652
rect 20044 36436 20084 36476
rect 20428 37612 20468 37652
rect 20048 36268 20088 36308
rect 20130 36268 20170 36308
rect 20212 36268 20252 36308
rect 20294 36268 20334 36308
rect 20376 36268 20416 36308
rect 20428 34924 20468 34964
rect 20048 34756 20088 34796
rect 20130 34756 20170 34796
rect 20212 34756 20252 34796
rect 20294 34756 20334 34796
rect 20376 34756 20416 34796
rect 19948 34084 19988 34124
rect 20140 34504 20180 34544
rect 19852 33496 19892 33536
rect 19756 33328 19796 33368
rect 19372 30808 19412 30848
rect 19564 32320 19604 32360
rect 19660 32656 19700 32696
rect 19372 30640 19412 30680
rect 19180 29632 19220 29672
rect 18808 29464 18848 29504
rect 18890 29464 18930 29504
rect 18972 29464 19012 29504
rect 19054 29464 19094 29504
rect 19136 29464 19176 29504
rect 19180 29296 19220 29336
rect 18808 27952 18848 27992
rect 18890 27952 18930 27992
rect 18972 27952 19012 27992
rect 19054 27952 19094 27992
rect 19136 27952 19176 27992
rect 19276 27952 19316 27992
rect 18892 27784 18932 27824
rect 19180 26692 19220 26732
rect 18604 24592 18644 24632
rect 18808 26440 18848 26480
rect 18890 26440 18930 26480
rect 18972 26440 19012 26480
rect 19054 26440 19094 26480
rect 19136 26440 19176 26480
rect 18796 26272 18836 26312
rect 18796 25768 18836 25808
rect 18808 24928 18848 24968
rect 18890 24928 18930 24968
rect 18972 24928 19012 24968
rect 19054 24928 19094 24968
rect 19136 24928 19176 24968
rect 19564 30640 19604 30680
rect 19564 29800 19604 29840
rect 19756 30556 19796 30596
rect 20140 34336 20180 34376
rect 20044 33412 20084 33452
rect 20048 33244 20088 33284
rect 20130 33244 20170 33284
rect 20212 33244 20252 33284
rect 20294 33244 20334 33284
rect 20376 33244 20416 33284
rect 20620 33412 20660 33452
rect 20140 33076 20180 33116
rect 20044 32992 20084 33032
rect 20236 31984 20276 32024
rect 20332 33076 20372 33116
rect 20524 32068 20564 32108
rect 20048 31732 20088 31772
rect 20130 31732 20170 31772
rect 20212 31732 20252 31772
rect 20294 31732 20334 31772
rect 20376 31732 20416 31772
rect 20428 31564 20468 31604
rect 20044 31480 20084 31520
rect 20140 30640 20180 30680
rect 20044 30472 20084 30512
rect 20048 30220 20088 30260
rect 20130 30220 20170 30260
rect 20212 30220 20252 30260
rect 20294 30220 20334 30260
rect 20376 30220 20416 30260
rect 19468 27364 19508 27404
rect 19564 27952 19604 27992
rect 18508 23668 18548 23708
rect 18412 23164 18452 23204
rect 18604 23752 18644 23792
rect 18508 22408 18548 22448
rect 18604 23416 18644 23456
rect 18508 21568 18548 21608
rect 18316 19048 18356 19088
rect 18220 18124 18260 18164
rect 18508 20224 18548 20264
rect 18220 17956 18260 17996
rect 18220 14932 18260 14972
rect 18808 23416 18848 23456
rect 18890 23416 18930 23456
rect 18972 23416 19012 23456
rect 19054 23416 19094 23456
rect 19136 23416 19176 23456
rect 18892 23248 18932 23288
rect 18796 23164 18836 23204
rect 19084 23080 19124 23120
rect 18700 22324 18740 22364
rect 18892 22324 18932 22364
rect 18796 22156 18836 22196
rect 18808 21904 18848 21944
rect 18890 21904 18930 21944
rect 18972 21904 19012 21944
rect 19054 21904 19094 21944
rect 19136 21904 19176 21944
rect 19180 21484 19220 21524
rect 18808 20392 18848 20432
rect 18890 20392 18930 20432
rect 18972 20392 19012 20432
rect 19054 20392 19094 20432
rect 19136 20392 19176 20432
rect 19084 20224 19124 20264
rect 19084 20056 19124 20096
rect 18892 19972 18932 20012
rect 18892 19300 18932 19340
rect 18808 18880 18848 18920
rect 18890 18880 18930 18920
rect 18972 18880 19012 18920
rect 19054 18880 19094 18920
rect 19136 18880 19176 18920
rect 18604 17872 18644 17912
rect 19660 27028 19700 27068
rect 19372 21568 19412 21608
rect 19372 19216 19412 19256
rect 19660 25012 19700 25052
rect 20048 28708 20088 28748
rect 20130 28708 20170 28748
rect 20212 28708 20252 28748
rect 20294 28708 20334 28748
rect 20376 28708 20416 28748
rect 20140 27952 20180 27992
rect 20620 28204 20660 28244
rect 20048 27196 20088 27236
rect 20130 27196 20170 27236
rect 20212 27196 20252 27236
rect 20294 27196 20334 27236
rect 20376 27196 20416 27236
rect 20044 27028 20084 27068
rect 20044 26020 20084 26060
rect 20048 25684 20088 25724
rect 20130 25684 20170 25724
rect 20212 25684 20252 25724
rect 20294 25684 20334 25724
rect 20376 25684 20416 25724
rect 20524 25432 20564 25472
rect 20044 25012 20084 25052
rect 20140 24844 20180 24884
rect 20908 43240 20948 43280
rect 21196 45256 21236 45296
rect 21004 37360 21044 37400
rect 20716 28036 20756 28076
rect 20812 35764 20852 35804
rect 20716 27868 20756 27908
rect 21100 35932 21140 35972
rect 21292 44920 21332 44960
rect 21292 37360 21332 37400
rect 21196 35764 21236 35804
rect 21196 33412 21236 33452
rect 21196 33244 21236 33284
rect 21484 33328 21524 33368
rect 21484 33160 21524 33200
rect 20908 28204 20948 28244
rect 20812 27280 20852 27320
rect 20908 27952 20948 27992
rect 20812 26020 20852 26060
rect 20620 24592 20660 24632
rect 20048 24172 20088 24212
rect 20130 24172 20170 24212
rect 20212 24172 20252 24212
rect 20294 24172 20334 24212
rect 20376 24172 20416 24212
rect 19852 23584 19892 23624
rect 20048 22660 20088 22700
rect 20130 22660 20170 22700
rect 20212 22660 20252 22700
rect 20294 22660 20334 22700
rect 20376 22660 20416 22700
rect 18808 17368 18848 17408
rect 18890 17368 18930 17408
rect 18972 17368 19012 17408
rect 19054 17368 19094 17408
rect 19136 17368 19176 17408
rect 18892 16276 18932 16316
rect 18808 15856 18848 15896
rect 18890 15856 18930 15896
rect 18972 15856 19012 15896
rect 19054 15856 19094 15896
rect 19136 15856 19176 15896
rect 19372 15436 19412 15476
rect 18508 14008 18548 14048
rect 18220 13000 18260 13040
rect 18220 12832 18260 12872
rect 18124 7120 18164 7160
rect 16396 1408 16436 1448
rect 16012 1240 16052 1280
rect 15820 1156 15860 1196
rect 15628 568 15668 608
rect 16204 232 16244 272
rect 16780 1324 16820 1364
rect 16588 400 16628 440
rect 17164 820 17204 860
rect 16972 148 17012 188
rect 17548 316 17588 356
rect 17932 988 17972 1028
rect 18808 14344 18848 14384
rect 18890 14344 18930 14384
rect 18972 14344 19012 14384
rect 19054 14344 19094 14384
rect 19136 14344 19176 14384
rect 19372 14008 19412 14048
rect 18808 12832 18848 12872
rect 18890 12832 18930 12872
rect 18972 12832 19012 12872
rect 19054 12832 19094 12872
rect 19136 12832 19176 12872
rect 18508 12412 18548 12452
rect 18808 11320 18848 11360
rect 18890 11320 18930 11360
rect 18972 11320 19012 11360
rect 19054 11320 19094 11360
rect 19136 11320 19176 11360
rect 18808 9808 18848 9848
rect 18890 9808 18930 9848
rect 18972 9808 19012 9848
rect 19054 9808 19094 9848
rect 19136 9808 19176 9848
rect 18808 8296 18848 8336
rect 18890 8296 18930 8336
rect 18972 8296 19012 8336
rect 19054 8296 19094 8336
rect 19136 8296 19176 8336
rect 18808 6784 18848 6824
rect 18890 6784 18930 6824
rect 18972 6784 19012 6824
rect 19054 6784 19094 6824
rect 19136 6784 19176 6824
rect 18808 5272 18848 5312
rect 18890 5272 18930 5312
rect 18972 5272 19012 5312
rect 19054 5272 19094 5312
rect 19136 5272 19176 5312
rect 18808 3760 18848 3800
rect 18890 3760 18930 3800
rect 18972 3760 19012 3800
rect 19054 3760 19094 3800
rect 19136 3760 19176 3800
rect 18700 3172 18740 3212
rect 18808 2248 18848 2288
rect 18890 2248 18930 2288
rect 18972 2248 19012 2288
rect 19054 2248 19094 2288
rect 19136 2248 19176 2288
rect 20428 22240 20468 22280
rect 19948 22156 19988 22196
rect 20048 21148 20088 21188
rect 20130 21148 20170 21188
rect 20212 21148 20252 21188
rect 20294 21148 20334 21188
rect 20376 21148 20416 21188
rect 20140 20728 20180 20768
rect 20044 20056 20084 20096
rect 20428 19888 20468 19928
rect 20044 19804 20084 19844
rect 20048 19636 20088 19676
rect 20130 19636 20170 19676
rect 20212 19636 20252 19676
rect 20294 19636 20334 19676
rect 20376 19636 20416 19676
rect 20140 19468 20180 19508
rect 19852 19216 19892 19256
rect 20524 19216 20564 19256
rect 20140 18544 20180 18584
rect 19756 15856 19796 15896
rect 20048 18124 20088 18164
rect 20130 18124 20170 18164
rect 20212 18124 20252 18164
rect 20294 18124 20334 18164
rect 20376 18124 20416 18164
rect 20140 17704 20180 17744
rect 20044 17032 20084 17072
rect 20140 17116 20180 17156
rect 20048 16612 20088 16652
rect 20130 16612 20170 16652
rect 20212 16612 20252 16652
rect 20294 16612 20334 16652
rect 20376 16612 20416 16652
rect 19948 15856 19988 15896
rect 19564 13672 19604 13712
rect 19852 11824 19892 11864
rect 20048 15100 20088 15140
rect 20130 15100 20170 15140
rect 20212 15100 20252 15140
rect 20294 15100 20334 15140
rect 20376 15100 20416 15140
rect 20716 19888 20756 19928
rect 20716 19216 20756 19256
rect 21292 27868 21332 27908
rect 20908 22912 20948 22952
rect 21004 24592 21044 24632
rect 20048 13588 20088 13628
rect 20130 13588 20170 13628
rect 20212 13588 20252 13628
rect 20294 13588 20334 13628
rect 20376 13588 20416 13628
rect 20048 12076 20088 12116
rect 20130 12076 20170 12116
rect 20212 12076 20252 12116
rect 20294 12076 20334 12116
rect 20376 12076 20416 12116
rect 20048 10564 20088 10604
rect 20130 10564 20170 10604
rect 20212 10564 20252 10604
rect 20294 10564 20334 10604
rect 20376 10564 20416 10604
rect 21292 22240 21332 22280
rect 21388 22912 21428 22952
rect 20044 9724 20084 9764
rect 20048 9052 20088 9092
rect 20130 9052 20170 9092
rect 20212 9052 20252 9092
rect 20294 9052 20334 9092
rect 20376 9052 20416 9092
rect 20048 7540 20088 7580
rect 20130 7540 20170 7580
rect 20212 7540 20252 7580
rect 20294 7540 20334 7580
rect 20376 7540 20416 7580
rect 20048 6028 20088 6068
rect 20130 6028 20170 6068
rect 20212 6028 20252 6068
rect 20294 6028 20334 6068
rect 20376 6028 20416 6068
rect 20048 4516 20088 4556
rect 20130 4516 20170 4556
rect 20212 4516 20252 4556
rect 20294 4516 20334 4556
rect 20376 4516 20416 4556
rect 20048 3004 20088 3044
rect 20130 3004 20170 3044
rect 20212 3004 20252 3044
rect 20294 3004 20334 3044
rect 20376 3004 20416 3044
rect 20048 1492 20088 1532
rect 20130 1492 20170 1532
rect 20212 1492 20252 1532
rect 20294 1492 20334 1532
rect 20376 1492 20416 1532
rect 19276 1408 19316 1448
rect 18508 1240 18548 1280
rect 18316 484 18356 524
rect 18700 1156 18740 1196
rect 19084 148 19124 188
rect 19468 1408 19508 1448
<< metal4 >>
rect 9091 96580 9100 96620
rect 9140 96580 14668 96620
rect 14708 96580 14717 96620
rect 12547 95908 12556 95948
rect 12596 95908 14284 95948
rect 14324 95908 14333 95948
rect 9475 95656 9484 95696
rect 9524 95656 15436 95696
rect 15476 95656 15485 95696
rect 4579 95572 4588 95612
rect 4628 95572 5260 95612
rect 5300 95572 5309 95612
rect 17347 95572 17356 95612
rect 17396 95572 18028 95612
rect 18068 95572 18077 95612
rect 4919 95236 4928 95276
rect 4968 95236 5010 95276
rect 5050 95236 5092 95276
rect 5132 95236 5174 95276
rect 5214 95236 5256 95276
rect 5296 95236 5305 95276
rect 20039 95236 20048 95276
rect 20088 95236 20130 95276
rect 20170 95236 20212 95276
rect 20252 95236 20294 95276
rect 20334 95236 20376 95276
rect 20416 95236 20425 95276
rect 3619 94900 3628 94940
rect 3668 94900 10636 94940
rect 10676 94900 10685 94940
rect 1229 94816 1324 94856
rect 1364 94816 1373 94856
rect 1699 94816 1708 94856
rect 1748 94816 1804 94856
rect 1844 94816 1853 94856
rect 1997 94816 2092 94856
rect 2132 94816 2141 94856
rect 2381 94816 2476 94856
rect 2516 94816 2525 94856
rect 3331 94816 3340 94856
rect 3380 94816 4012 94856
rect 4052 94816 4061 94856
rect 4301 94816 4396 94856
rect 4436 94816 4445 94856
rect 4675 94816 4684 94856
rect 4724 94816 5548 94856
rect 5588 94816 5597 94856
rect 6221 94816 6316 94856
rect 6356 94816 6365 94856
rect 6605 94816 6700 94856
rect 6740 94816 6749 94856
rect 6989 94816 7084 94856
rect 7124 94816 7133 94856
rect 18125 94816 18220 94856
rect 18260 94816 18269 94856
rect 18403 94816 18412 94856
rect 18452 94816 18796 94856
rect 18836 94816 18845 94856
rect 19075 94816 19084 94856
rect 19124 94816 19468 94856
rect 19508 94816 19517 94856
rect 10637 94732 10732 94772
rect 10772 94732 10781 94772
rect 12269 94732 12364 94772
rect 12404 94732 12413 94772
rect 13219 94732 13228 94772
rect 13268 94732 13420 94772
rect 13460 94732 13469 94772
rect 14285 94732 14380 94772
rect 14420 94732 14429 94772
rect 8717 94648 8812 94688
rect 8852 94648 8861 94688
rect 9293 94648 9388 94688
rect 9428 94648 9437 94688
rect 9677 94648 9772 94688
rect 9812 94648 9821 94688
rect 10445 94648 10540 94688
rect 10580 94648 10589 94688
rect 11117 94648 11212 94688
rect 11252 94648 11261 94688
rect 11501 94648 11596 94688
rect 11636 94648 11645 94688
rect 12077 94648 12172 94688
rect 12212 94648 12221 94688
rect 3679 94480 3688 94520
rect 3728 94480 3770 94520
rect 3810 94480 3852 94520
rect 3892 94480 3934 94520
rect 3974 94480 4016 94520
rect 4056 94480 4065 94520
rect 18799 94480 18808 94520
rect 18848 94480 18890 94520
rect 18930 94480 18972 94520
rect 19012 94480 19054 94520
rect 19094 94480 19136 94520
rect 19176 94480 19185 94520
rect 19075 94228 19084 94268
rect 19124 94228 19564 94268
rect 19604 94228 19613 94268
rect 4483 94144 4492 94184
rect 4532 94144 4972 94184
rect 5012 94144 5021 94184
rect 5347 94144 5356 94184
rect 5396 94144 5548 94184
rect 5588 94144 5597 94184
rect 5645 94144 5740 94184
rect 5780 94144 5789 94184
rect 6029 94144 6124 94184
rect 6164 94144 6173 94184
rect 7949 94144 8044 94184
rect 8084 94144 8093 94184
rect 11491 94144 11500 94184
rect 11540 94144 12748 94184
rect 12788 94144 12797 94184
rect 16109 94144 16204 94184
rect 16244 94144 16253 94184
rect 16877 94144 16972 94184
rect 17012 94144 17021 94184
rect 18019 94144 18028 94184
rect 18068 94144 18124 94184
rect 18164 94144 18173 94184
rect 18595 94144 18604 94184
rect 18644 94144 18988 94184
rect 19028 94144 19037 94184
rect 19363 94144 19372 94184
rect 19412 94144 19852 94184
rect 19892 94144 19901 94184
rect 20227 94144 20236 94184
rect 20276 94144 21484 94184
rect 21524 94144 21533 94184
rect 12451 94060 12460 94100
rect 12500 94060 19756 94100
rect 19796 94060 19805 94100
rect 9869 93976 9964 94016
rect 10004 93976 10013 94016
rect 10925 93976 11020 94016
rect 11060 93976 11069 94016
rect 4579 93892 4588 93932
rect 4628 93892 5932 93932
rect 5972 93892 5981 93932
rect 7747 93892 7756 93932
rect 7796 93892 8236 93932
rect 8276 93892 8285 93932
rect 10061 93892 10156 93932
rect 10196 93892 10205 93932
rect 10733 93892 10828 93932
rect 10868 93892 10877 93932
rect 11107 93892 11116 93932
rect 11156 93892 12940 93932
rect 12980 93892 12989 93932
rect 13805 93892 13900 93932
rect 13940 93892 13949 93932
rect 14189 93892 14284 93932
rect 14324 93892 14333 93932
rect 14573 93892 14668 93932
rect 14708 93892 14717 93932
rect 15053 93892 15148 93932
rect 15188 93892 15197 93932
rect 16493 93892 16588 93932
rect 16628 93892 16637 93932
rect 17645 93892 17740 93932
rect 17780 93892 17789 93932
rect 3139 93808 3148 93848
rect 3188 93808 6892 93848
rect 6932 93808 6941 93848
rect 4919 93724 4928 93764
rect 4968 93724 5010 93764
rect 5050 93724 5092 93764
rect 5132 93724 5174 93764
rect 5214 93724 5256 93764
rect 5296 93724 5305 93764
rect 11875 93724 11884 93764
rect 11924 93724 13036 93764
rect 13076 93724 13085 93764
rect 20039 93724 20048 93764
rect 20088 93724 20130 93764
rect 20170 93724 20212 93764
rect 20252 93724 20294 93764
rect 20334 93724 20376 93764
rect 20416 93724 20425 93764
rect 16771 93640 16780 93680
rect 16820 93640 17356 93680
rect 17396 93640 17405 93680
rect 2563 93556 2572 93596
rect 2612 93556 2860 93596
rect 2900 93556 2909 93596
rect 7085 93556 7180 93596
rect 7220 93556 7229 93596
rect 17155 93304 17164 93344
rect 17204 93304 18988 93344
rect 19028 93304 19037 93344
rect 19843 93304 19852 93344
rect 19892 93304 19948 93344
rect 19988 93304 19997 93344
rect 20131 93304 20140 93344
rect 20180 93304 21388 93344
rect 21428 93304 21437 93344
rect 18115 93136 18124 93176
rect 18164 93136 18700 93176
rect 18740 93136 18749 93176
rect 3679 92968 3688 93008
rect 3728 92968 3770 93008
rect 3810 92968 3852 93008
rect 3892 92968 3934 93008
rect 3974 92968 4016 93008
rect 4056 92968 4065 93008
rect 18799 92968 18808 93008
rect 18848 92968 18890 93008
rect 18930 92968 18972 93008
rect 19012 92968 19054 93008
rect 19094 92968 19136 93008
rect 19176 92968 19185 93008
rect 2947 92632 2956 92672
rect 2996 92632 9292 92672
rect 9332 92632 9341 92672
rect 19373 92632 19468 92672
rect 19508 92632 19517 92672
rect 19651 92632 19660 92672
rect 19700 92632 19756 92672
rect 19796 92632 19805 92672
rect 2755 92296 2764 92336
rect 2804 92296 6604 92336
rect 6644 92296 6653 92336
rect 4919 92212 4928 92252
rect 4968 92212 5010 92252
rect 5050 92212 5092 92252
rect 5132 92212 5174 92252
rect 5214 92212 5256 92252
rect 5296 92212 5305 92252
rect 20039 92212 20048 92252
rect 20088 92212 20130 92252
rect 20170 92212 20212 92252
rect 20252 92212 20294 92252
rect 20334 92212 20376 92252
rect 20416 92212 20425 92252
rect 8035 91792 8044 91832
rect 8084 91792 8332 91832
rect 8372 91792 8381 91832
rect 19555 91792 19564 91832
rect 19604 91792 19756 91832
rect 19796 91792 19805 91832
rect 3679 91456 3688 91496
rect 3728 91456 3770 91496
rect 3810 91456 3852 91496
rect 3892 91456 3934 91496
rect 3974 91456 4016 91496
rect 4056 91456 4065 91496
rect 18799 91456 18808 91496
rect 18848 91456 18890 91496
rect 18930 91456 18972 91496
rect 19012 91456 19054 91496
rect 19094 91456 19136 91496
rect 19176 91456 19185 91496
rect 7939 91120 7948 91160
rect 7988 91120 8140 91160
rect 8180 91120 8189 91160
rect 8323 91120 8332 91160
rect 8372 91120 8524 91160
rect 8564 91120 8573 91160
rect 20131 91120 20140 91160
rect 20180 91120 20908 91160
rect 20948 91120 20957 91160
rect 2957 90868 3052 90908
rect 3092 90868 3101 90908
rect 4919 90700 4928 90740
rect 4968 90700 5010 90740
rect 5050 90700 5092 90740
rect 5132 90700 5174 90740
rect 5214 90700 5256 90740
rect 5296 90700 5305 90740
rect 14381 90700 14476 90740
rect 14516 90700 14525 90740
rect 20039 90700 20048 90740
rect 20088 90700 20130 90740
rect 20170 90700 20212 90740
rect 20252 90700 20294 90740
rect 20334 90700 20376 90740
rect 20416 90700 20425 90740
rect 1411 90280 1420 90320
rect 1460 90280 2380 90320
rect 2420 90280 2429 90320
rect 20131 90280 20140 90320
rect 20180 90280 21292 90320
rect 21332 90280 21341 90320
rect 4003 90112 4012 90152
rect 4052 90112 4204 90152
rect 4244 90112 4253 90152
rect 2755 89944 2764 89984
rect 2804 89944 3532 89984
rect 3572 89944 3581 89984
rect 3679 89944 3688 89984
rect 3728 89944 3770 89984
rect 3810 89944 3852 89984
rect 3892 89944 3934 89984
rect 3974 89944 4016 89984
rect 4056 89944 4065 89984
rect 18799 89944 18808 89984
rect 18848 89944 18890 89984
rect 18930 89944 18972 89984
rect 19012 89944 19054 89984
rect 19094 89944 19136 89984
rect 19176 89944 19185 89984
rect 1411 89860 1420 89900
rect 1460 89860 10924 89900
rect 10964 89860 10973 89900
rect 1699 89776 1708 89816
rect 1748 89776 1996 89816
rect 2036 89776 2045 89816
rect 3619 89776 3628 89816
rect 3668 89776 6316 89816
rect 6356 89776 6365 89816
rect 1603 89692 1612 89732
rect 1652 89692 2860 89732
rect 2900 89692 2909 89732
rect 1411 89608 1420 89648
rect 1460 89608 1996 89648
rect 2036 89608 2045 89648
rect 3235 89608 3244 89648
rect 3284 89608 4588 89648
rect 4628 89608 4637 89648
rect 16483 89608 16492 89648
rect 16532 89608 19756 89648
rect 19796 89608 19805 89648
rect 20131 89608 20140 89648
rect 20180 89608 20812 89648
rect 20852 89608 20861 89648
rect 17347 89524 17356 89564
rect 17396 89524 17644 89564
rect 17684 89524 17693 89564
rect 1411 89440 1420 89480
rect 1460 89440 2860 89480
rect 2900 89440 2909 89480
rect 10051 89440 10060 89480
rect 10100 89440 13804 89480
rect 13844 89440 13853 89480
rect 1603 89356 1612 89396
rect 1652 89356 1996 89396
rect 2036 89356 2045 89396
rect 3043 89356 3052 89396
rect 3092 89356 3148 89396
rect 3188 89356 3197 89396
rect 3619 89356 3628 89396
rect 3668 89356 9772 89396
rect 9812 89356 9821 89396
rect 14765 89356 14860 89396
rect 14900 89356 14909 89396
rect 3628 89312 3668 89356
rect 2467 89272 2476 89312
rect 2516 89272 3668 89312
rect 4919 89188 4928 89228
rect 4968 89188 5010 89228
rect 5050 89188 5092 89228
rect 5132 89188 5174 89228
rect 5214 89188 5256 89228
rect 5296 89188 5305 89228
rect 12547 89188 12556 89228
rect 12596 89188 13228 89228
rect 13268 89188 13277 89228
rect 20039 89188 20048 89228
rect 20088 89188 20130 89228
rect 20170 89188 20212 89228
rect 20252 89188 20294 89228
rect 20334 89188 20376 89228
rect 20416 89188 20425 89228
rect 2851 89020 2860 89060
rect 2900 89020 3244 89060
rect 3284 89020 3293 89060
rect 14179 89020 14188 89060
rect 14228 89020 14284 89060
rect 14324 89020 14333 89060
rect 16291 89020 16300 89060
rect 16340 89020 16396 89060
rect 16436 89020 16445 89060
rect 4387 88936 4396 88976
rect 4436 88936 4684 88976
rect 4724 88936 4733 88976
rect 2947 88852 2956 88892
rect 2996 88852 3244 88892
rect 3284 88852 3293 88892
rect 12259 88852 12268 88892
rect 12308 88852 18988 88892
rect 19028 88852 19037 88892
rect 18509 88768 18604 88808
rect 18644 88768 18653 88808
rect 7651 88684 7660 88724
rect 7700 88684 19372 88724
rect 19412 88684 19421 88724
rect 7555 88600 7564 88640
rect 7604 88600 8044 88640
rect 8084 88600 8093 88640
rect 20323 88600 20332 88640
rect 20372 88600 20524 88640
rect 20564 88600 20573 88640
rect 3679 88432 3688 88472
rect 3728 88432 3770 88472
rect 3810 88432 3852 88472
rect 3892 88432 3934 88472
rect 3974 88432 4016 88472
rect 4056 88432 4065 88472
rect 18799 88432 18808 88472
rect 18848 88432 18890 88472
rect 18930 88432 18972 88472
rect 19012 88432 19054 88472
rect 19094 88432 19136 88472
rect 19176 88432 19185 88472
rect 17347 88096 17356 88136
rect 17396 88096 18220 88136
rect 18260 88096 18269 88136
rect 2860 88012 9676 88052
rect 9716 88012 9725 88052
rect 11203 88012 11212 88052
rect 11252 88012 19852 88052
rect 19892 88012 19901 88052
rect 2860 87968 2900 88012
rect 2467 87928 2476 87968
rect 2516 87928 2900 87968
rect 5548 87928 8236 87968
rect 8276 87928 8285 87968
rect 12835 87928 12844 87968
rect 12884 87928 13132 87968
rect 13172 87928 13181 87968
rect 13699 87928 13708 87968
rect 13748 87928 19756 87968
rect 19796 87928 19805 87968
rect 5548 87884 5588 87928
rect 2755 87844 2764 87884
rect 2804 87844 5588 87884
rect 6019 87844 6028 87884
rect 6068 87844 6220 87884
rect 6260 87844 6269 87884
rect 15245 87844 15340 87884
rect 15380 87844 15389 87884
rect 15523 87844 15532 87884
rect 15572 87844 20140 87884
rect 20180 87844 20189 87884
rect 4919 87676 4928 87716
rect 4968 87676 5010 87716
rect 5050 87676 5092 87716
rect 5132 87676 5174 87716
rect 5214 87676 5256 87716
rect 5296 87676 5305 87716
rect 20039 87676 20048 87716
rect 20088 87676 20130 87716
rect 20170 87676 20212 87716
rect 20252 87676 20294 87716
rect 20334 87676 20376 87716
rect 20416 87676 20425 87716
rect 8621 87508 8716 87548
rect 8756 87508 8765 87548
rect 1123 87424 1132 87464
rect 1172 87424 1324 87464
rect 1364 87424 1373 87464
rect 17443 87424 17452 87464
rect 17492 87424 17644 87464
rect 17684 87424 17693 87464
rect 20515 87424 20524 87464
rect 20564 87424 20908 87464
rect 20948 87424 20957 87464
rect 21187 87424 21196 87464
rect 21236 87424 21484 87464
rect 21524 87424 21533 87464
rect 12931 87340 12940 87380
rect 12980 87340 13324 87380
rect 13364 87340 13373 87380
rect 2947 87256 2956 87296
rect 2996 87256 3340 87296
rect 3380 87256 3389 87296
rect 3523 87256 3532 87296
rect 3572 87256 3628 87296
rect 3668 87256 3677 87296
rect 5635 87256 5644 87296
rect 5684 87256 7852 87296
rect 7892 87256 7901 87296
rect 19661 87256 19756 87296
rect 19796 87256 19805 87296
rect 20131 87256 20140 87296
rect 20180 87256 21100 87296
rect 21140 87256 21149 87296
rect 4003 87088 4012 87128
rect 4052 87088 4148 87128
rect 5443 87088 5452 87128
rect 5492 87088 5740 87128
rect 5780 87088 5789 87128
rect 18604 87088 18796 87128
rect 18836 87088 18845 87128
rect 3679 86920 3688 86960
rect 3728 86920 3770 86960
rect 3810 86920 3852 86960
rect 3892 86920 3934 86960
rect 3974 86920 4016 86960
rect 4056 86920 4065 86960
rect 4108 86876 4148 87088
rect 18604 86960 18644 87088
rect 18595 86920 18604 86960
rect 18644 86920 18653 86960
rect 18799 86920 18808 86960
rect 18848 86920 18890 86960
rect 18930 86920 18972 86960
rect 19012 86920 19054 86960
rect 19094 86920 19136 86960
rect 19176 86920 19185 86960
rect 4012 86836 4148 86876
rect 4012 86792 4052 86836
rect 4003 86752 4012 86792
rect 4052 86752 4061 86792
rect 5635 86752 5644 86792
rect 5684 86752 7948 86792
rect 7988 86752 7997 86792
rect 5827 86668 5836 86708
rect 5876 86668 7276 86708
rect 7316 86668 7325 86708
rect 5155 86584 5164 86624
rect 5204 86584 6412 86624
rect 6452 86584 6461 86624
rect 20131 86584 20140 86624
rect 20180 86584 20716 86624
rect 20756 86584 20765 86624
rect 7853 86500 7948 86540
rect 7988 86500 7997 86540
rect 17731 86500 17740 86540
rect 17780 86500 17932 86540
rect 17972 86500 17981 86540
rect 13027 86416 13036 86456
rect 13076 86416 13171 86456
rect 16675 86416 16684 86456
rect 16724 86416 18796 86456
rect 18836 86416 18845 86456
rect 2179 86332 2188 86372
rect 2228 86332 2668 86372
rect 2708 86332 2717 86372
rect 8131 86332 8140 86372
rect 8180 86332 10252 86372
rect 10292 86332 10301 86372
rect 6787 86248 6796 86288
rect 6836 86248 7084 86288
rect 7124 86248 7133 86288
rect 739 86164 748 86204
rect 788 86164 1228 86204
rect 1268 86164 1277 86204
rect 4919 86164 4928 86204
rect 4968 86164 5010 86204
rect 5050 86164 5092 86204
rect 5132 86164 5174 86204
rect 5214 86164 5256 86204
rect 5296 86164 5305 86204
rect 12451 86164 12460 86204
rect 12500 86164 12844 86204
rect 12884 86164 12893 86204
rect 20039 86164 20048 86204
rect 20088 86164 20130 86204
rect 20170 86164 20212 86204
rect 20252 86164 20294 86204
rect 20334 86164 20376 86204
rect 20416 86164 20425 86204
rect 12547 86080 12556 86120
rect 12596 86080 13228 86120
rect 13268 86080 13277 86120
rect 7171 85996 7180 86036
rect 7220 85996 8812 86036
rect 8852 85996 8861 86036
rect 8419 85912 8428 85952
rect 8468 85912 8477 85952
rect 17251 85912 17260 85952
rect 17300 85912 17452 85952
rect 17492 85912 17501 85952
rect 8428 85868 8468 85912
rect 8428 85828 8620 85868
rect 8660 85828 8669 85868
rect 12355 85828 12364 85868
rect 12404 85828 13996 85868
rect 14036 85828 14045 85868
rect 2179 85744 2188 85784
rect 2228 85744 2572 85784
rect 2612 85744 2621 85784
rect 17741 85744 17836 85784
rect 17876 85744 17885 85784
rect 10349 85576 10444 85616
rect 10484 85576 10493 85616
rect 1411 85492 1420 85532
rect 1460 85492 1516 85532
rect 1556 85492 1565 85532
rect 3679 85408 3688 85448
rect 3728 85408 3770 85448
rect 3810 85408 3852 85448
rect 3892 85408 3934 85448
rect 3974 85408 4016 85448
rect 4056 85408 4065 85448
rect 18799 85408 18808 85448
rect 18848 85408 18890 85448
rect 18930 85408 18972 85448
rect 19012 85408 19054 85448
rect 19094 85408 19136 85448
rect 19176 85408 19185 85448
rect 21101 85408 21196 85448
rect 21236 85408 21245 85448
rect 12739 85240 12748 85280
rect 12788 85240 13708 85280
rect 13748 85240 13757 85280
rect 14083 85156 14092 85196
rect 14132 85156 14188 85196
rect 14228 85156 14237 85196
rect 2947 85072 2956 85112
rect 2996 85072 3244 85112
rect 3284 85072 3293 85112
rect 4387 85072 4396 85112
rect 4436 85072 4780 85112
rect 4820 85072 4829 85112
rect 5357 85072 5452 85112
rect 5492 85072 5501 85112
rect 7747 85072 7756 85112
rect 7796 85072 7852 85112
rect 7892 85072 7901 85112
rect 20707 85072 20716 85112
rect 20756 85072 20852 85112
rect 2659 84988 2668 85028
rect 2708 84988 3244 85028
rect 3284 84988 3293 85028
rect 10147 84988 10156 85028
rect 10196 84988 12940 85028
rect 12980 84988 13132 85028
rect 13172 84988 13181 85028
rect 13987 84988 13996 85028
rect 14036 84988 14188 85028
rect 14228 84988 14237 85028
rect 20812 84944 20852 85072
rect 3619 84904 3628 84944
rect 3668 84904 8524 84944
rect 8564 84904 8573 84944
rect 12451 84904 12460 84944
rect 12500 84904 15244 84944
rect 15284 84904 15293 84944
rect 20803 84904 20812 84944
rect 20852 84904 20861 84944
rect 16781 84820 16876 84860
rect 16916 84820 16925 84860
rect 8419 84736 8428 84776
rect 8468 84736 16012 84776
rect 16052 84736 16061 84776
rect 4919 84652 4928 84692
rect 4968 84652 5010 84692
rect 5050 84652 5092 84692
rect 5132 84652 5174 84692
rect 5214 84652 5256 84692
rect 5296 84652 5305 84692
rect 11491 84652 11500 84692
rect 11540 84652 14188 84692
rect 14228 84652 14237 84692
rect 20039 84652 20048 84692
rect 20088 84652 20130 84692
rect 20170 84652 20212 84692
rect 20252 84652 20294 84692
rect 20334 84652 20376 84692
rect 20416 84652 20425 84692
rect 3715 84568 3724 84608
rect 3764 84568 6988 84608
rect 7028 84568 7037 84608
rect 20515 84568 20524 84608
rect 20564 84568 20908 84608
rect 20948 84568 20957 84608
rect 4675 84484 4684 84524
rect 4724 84484 4733 84524
rect 5453 84484 5548 84524
rect 5588 84484 5597 84524
rect 5731 84484 5740 84524
rect 5780 84484 5836 84524
rect 5876 84484 5885 84524
rect 11971 84484 11980 84524
rect 12020 84484 15052 84524
rect 15092 84484 15101 84524
rect 3427 84316 3436 84356
rect 3476 84316 3724 84356
rect 3764 84316 3773 84356
rect 1891 84232 1900 84272
rect 1940 84232 2764 84272
rect 2804 84232 2813 84272
rect 4684 84188 4724 84484
rect 18115 84400 18124 84440
rect 18164 84400 18173 84440
rect 12547 84316 12556 84356
rect 12596 84316 14860 84356
rect 14900 84316 14909 84356
rect 18124 84272 18164 84400
rect 6691 84232 6700 84272
rect 6740 84232 7084 84272
rect 7124 84232 7133 84272
rect 14467 84232 14476 84272
rect 14516 84232 15724 84272
rect 15764 84232 15773 84272
rect 18124 84232 18508 84272
rect 18548 84232 18557 84272
rect 20131 84232 20140 84272
rect 20180 84232 21004 84272
rect 21044 84232 21053 84272
rect 4291 84148 4300 84188
rect 4340 84148 4724 84188
rect 8131 84148 8140 84188
rect 8180 84148 8332 84188
rect 8372 84148 8381 84188
rect 8899 84148 8908 84188
rect 8948 84148 10636 84188
rect 10676 84148 10685 84188
rect 14467 84148 14476 84188
rect 14516 84148 14572 84188
rect 14612 84148 14621 84188
rect 19267 84148 19276 84188
rect 19316 84148 19372 84188
rect 19412 84148 19421 84188
rect 1517 84064 1612 84104
rect 1652 84064 1661 84104
rect 1805 84064 1900 84104
rect 1940 84064 1949 84104
rect 4003 84064 4012 84104
rect 4052 84064 4061 84104
rect 7363 84064 7372 84104
rect 7412 84064 7948 84104
rect 7988 84064 7997 84104
rect 13795 84064 13804 84104
rect 13844 84064 17740 84104
rect 17780 84064 17789 84104
rect 18787 84064 18796 84104
rect 18836 84064 19412 84104
rect 4012 84020 4052 84064
rect 2659 83980 2668 84020
rect 2708 83980 2860 84020
rect 2900 83980 2909 84020
rect 4012 83980 4148 84020
rect 13219 83980 13228 84020
rect 13268 83980 13612 84020
rect 13652 83980 13661 84020
rect 17644 83980 17836 84020
rect 17876 83980 17885 84020
rect 3679 83896 3688 83936
rect 3728 83896 3770 83936
rect 3810 83896 3852 83936
rect 3892 83896 3934 83936
rect 3974 83896 4016 83936
rect 4056 83896 4065 83936
rect 2371 83644 2380 83684
rect 2420 83644 3724 83684
rect 3764 83644 3773 83684
rect 4108 83600 4148 83980
rect 8707 83896 8716 83936
rect 8756 83896 9196 83936
rect 9236 83896 9245 83936
rect 13699 83896 13708 83936
rect 13748 83896 14092 83936
rect 14132 83896 14141 83936
rect 7459 83812 7468 83852
rect 7508 83812 8332 83852
rect 8372 83812 8381 83852
rect 17165 83812 17260 83852
rect 17300 83812 17309 83852
rect 9283 83728 9292 83768
rect 9332 83728 9676 83768
rect 9716 83728 9725 83768
rect 13997 83728 14092 83768
rect 14132 83728 14141 83768
rect 4204 83644 4396 83684
rect 4436 83644 4445 83684
rect 9187 83644 9196 83684
rect 9236 83644 9964 83684
rect 10004 83644 10013 83684
rect 12076 83644 12268 83684
rect 12308 83644 12317 83684
rect 13507 83644 13516 83684
rect 13556 83644 13565 83684
rect 14275 83644 14284 83684
rect 14324 83644 16012 83684
rect 16052 83644 16061 83684
rect 3149 83560 3244 83600
rect 3284 83560 3293 83600
rect 4099 83560 4108 83600
rect 4148 83560 4157 83600
rect 1507 83392 1516 83432
rect 1556 83392 1708 83432
rect 1748 83392 1757 83432
rect 2659 83392 2668 83432
rect 2708 83392 2764 83432
rect 2804 83392 2813 83432
rect 4204 83264 4244 83644
rect 4291 83476 4300 83516
rect 4340 83476 4349 83516
rect 5347 83476 5356 83516
rect 5396 83476 5452 83516
rect 5492 83476 5501 83516
rect 6979 83476 6988 83516
rect 7028 83476 9964 83516
rect 10004 83476 10013 83516
rect 4300 83432 4340 83476
rect 4300 83392 9004 83432
rect 9044 83392 9053 83432
rect 12076 83348 12116 83644
rect 13516 83600 13556 83644
rect 17644 83600 17684 83980
rect 19372 83936 19412 84064
rect 18799 83896 18808 83936
rect 18848 83896 18890 83936
rect 18930 83896 18972 83936
rect 19012 83896 19054 83936
rect 19094 83896 19136 83936
rect 19176 83896 19185 83936
rect 19363 83896 19372 83936
rect 19412 83896 19421 83936
rect 18796 83812 19564 83852
rect 19604 83812 19613 83852
rect 18796 83768 18836 83812
rect 18787 83728 18796 83768
rect 18836 83728 18845 83768
rect 13219 83560 13228 83600
rect 13268 83560 13556 83600
rect 14755 83560 14764 83600
rect 14804 83560 15052 83600
rect 15092 83560 15101 83600
rect 17155 83560 17164 83600
rect 17204 83560 17452 83600
rect 17492 83560 17501 83600
rect 17635 83560 17644 83600
rect 17684 83560 17693 83600
rect 18403 83560 18412 83600
rect 18452 83560 18988 83600
rect 19028 83560 19037 83600
rect 20131 83560 20140 83600
rect 20180 83560 21292 83600
rect 21332 83560 21341 83600
rect 15619 83476 15628 83516
rect 15668 83476 17068 83516
rect 17108 83476 17117 83516
rect 19939 83476 19948 83516
rect 19988 83476 19997 83516
rect 17155 83392 17164 83432
rect 17204 83392 17452 83432
rect 17492 83392 17501 83432
rect 18307 83392 18316 83432
rect 18356 83392 19084 83432
rect 19124 83392 19133 83432
rect 4387 83308 4396 83348
rect 4436 83308 4780 83348
rect 4820 83308 7660 83348
rect 7700 83308 7709 83348
rect 12067 83308 12076 83348
rect 12116 83308 12125 83348
rect 3139 83224 3148 83264
rect 3188 83224 4244 83264
rect 5539 83224 5548 83264
rect 5588 83224 5836 83264
rect 5876 83224 5885 83264
rect 6979 83224 6988 83264
rect 7028 83224 7948 83264
rect 7988 83224 8524 83264
rect 8564 83224 8573 83264
rect 4919 83140 4928 83180
rect 4968 83140 5010 83180
rect 5050 83140 5092 83180
rect 5132 83140 5174 83180
rect 5214 83140 5256 83180
rect 5296 83140 5305 83180
rect 14371 83140 14380 83180
rect 14420 83140 15340 83180
rect 15380 83140 15389 83180
rect 3427 83056 3436 83096
rect 3476 83056 4300 83096
rect 4340 83056 4349 83096
rect 14755 83056 14764 83096
rect 14804 83056 17260 83096
rect 17300 83056 17309 83096
rect 19948 83012 19988 83476
rect 20039 83140 20048 83180
rect 20088 83140 20130 83180
rect 20170 83140 20212 83180
rect 20252 83140 20294 83180
rect 20334 83140 20376 83180
rect 20416 83140 20425 83180
rect 3523 82972 3532 83012
rect 3572 82972 4300 83012
rect 4340 82972 4349 83012
rect 4771 82972 4780 83012
rect 4820 82972 4829 83012
rect 4963 82972 4972 83012
rect 5012 82972 11980 83012
rect 12020 82972 12029 83012
rect 19948 82972 20044 83012
rect 20084 82972 20093 83012
rect 4780 82928 4820 82972
rect 4195 82888 4204 82928
rect 4244 82888 4253 82928
rect 4675 82888 4684 82928
rect 4724 82888 4820 82928
rect 4204 82844 4244 82888
rect 4204 82804 4780 82844
rect 4820 82804 4829 82844
rect 10435 82804 10444 82844
rect 10484 82804 12748 82844
rect 12788 82804 12797 82844
rect 3523 82720 3532 82760
rect 3572 82720 3612 82760
rect 4291 82720 4300 82760
rect 4340 82720 5836 82760
rect 5876 82720 5885 82760
rect 13997 82720 14092 82760
rect 14132 82720 14141 82760
rect 17923 82720 17932 82760
rect 17972 82720 18316 82760
rect 18356 82720 18365 82760
rect 3532 82676 3572 82720
rect 1891 82636 1900 82676
rect 1940 82636 4876 82676
rect 4916 82636 4925 82676
rect 16013 82636 16108 82676
rect 16148 82636 16157 82676
rect 3523 82552 3532 82592
rect 3572 82552 3724 82592
rect 3764 82552 3773 82592
rect 3907 82552 3916 82592
rect 3956 82552 8908 82592
rect 8948 82552 8957 82592
rect 19276 82552 19372 82592
rect 19412 82552 19421 82592
rect 3916 82508 3956 82552
rect 3235 82468 3244 82508
rect 3284 82468 3956 82508
rect 14083 82468 14092 82508
rect 14132 82468 15244 82508
rect 15284 82468 15293 82508
rect 3679 82384 3688 82424
rect 3728 82384 3770 82424
rect 3810 82384 3852 82424
rect 3892 82384 3934 82424
rect 3974 82384 4016 82424
rect 4056 82384 4065 82424
rect 18799 82384 18808 82424
rect 18848 82384 18890 82424
rect 18930 82384 18972 82424
rect 19012 82384 19054 82424
rect 19094 82384 19136 82424
rect 19176 82384 19185 82424
rect 19276 82340 19316 82552
rect 19363 82384 19372 82424
rect 19412 82384 19564 82424
rect 19604 82384 19613 82424
rect 1315 82300 1324 82340
rect 1364 82300 1900 82340
rect 1940 82300 1949 82340
rect 18988 82300 19316 82340
rect 18988 82256 19028 82300
rect 5827 82216 5836 82256
rect 5876 82216 5932 82256
rect 5972 82216 5981 82256
rect 6211 82216 6220 82256
rect 6260 82216 6412 82256
rect 6452 82216 6461 82256
rect 8803 82216 8812 82256
rect 8852 82216 8948 82256
rect 18979 82216 18988 82256
rect 19028 82216 19037 82256
rect 1891 82132 1900 82172
rect 1940 82132 2476 82172
rect 2516 82132 2525 82172
rect 1325 82048 1420 82088
rect 1460 82048 1469 82088
rect 4003 82048 4012 82088
rect 4052 82048 4780 82088
rect 4820 82048 4829 82088
rect 3523 81964 3532 82004
rect 3572 81964 3820 82004
rect 3860 81964 3869 82004
rect 4867 81964 4876 82004
rect 4916 81964 8812 82004
rect 8852 81964 8861 82004
rect 8908 81920 8948 82216
rect 13603 82132 13612 82172
rect 13652 82132 14860 82172
rect 14900 82132 14909 82172
rect 15331 82132 15340 82172
rect 15380 82132 15389 82172
rect 16963 82132 16972 82172
rect 17012 82132 17021 82172
rect 15340 82088 15380 82132
rect 10435 82048 10444 82088
rect 10484 82048 10636 82088
rect 10676 82048 10685 82088
rect 13795 82048 13804 82088
rect 13844 82048 14380 82088
rect 14420 82048 14429 82088
rect 14860 82048 15380 82088
rect 16483 82048 16492 82088
rect 16532 82048 16780 82088
rect 16820 82048 16829 82088
rect 14860 82004 14900 82048
rect 14851 81964 14860 82004
rect 14900 81964 14909 82004
rect 2467 81880 2476 81920
rect 2516 81880 8908 81920
rect 8948 81880 8957 81920
rect 4963 81796 4972 81836
rect 5012 81796 7468 81836
rect 7508 81796 7517 81836
rect 13795 81796 13804 81836
rect 13844 81796 14092 81836
rect 14132 81796 14141 81836
rect 14755 81796 14764 81836
rect 14804 81796 16684 81836
rect 16724 81796 16733 81836
rect 16972 81752 17012 82132
rect 17923 81796 17932 81836
rect 17972 81796 18316 81836
rect 18356 81796 18365 81836
rect 20035 81796 20044 81836
rect 20084 81796 20093 81836
rect 20044 81752 20084 81796
rect 13315 81712 13324 81752
rect 13364 81712 13996 81752
rect 14036 81712 14045 81752
rect 15619 81712 15628 81752
rect 15668 81712 17012 81752
rect 19948 81712 20084 81752
rect 4919 81628 4928 81668
rect 4968 81628 5010 81668
rect 5050 81628 5092 81668
rect 5132 81628 5174 81668
rect 5214 81628 5256 81668
rect 5296 81628 5305 81668
rect 6499 81628 6508 81668
rect 6548 81628 6892 81668
rect 6932 81628 6941 81668
rect 8707 81544 8716 81584
rect 8756 81544 9100 81584
rect 9140 81544 9149 81584
rect 13507 81544 13516 81584
rect 13556 81544 16108 81584
rect 16148 81544 16157 81584
rect 5155 81460 5164 81500
rect 5204 81460 5548 81500
rect 5588 81460 5597 81500
rect 6019 81460 6028 81500
rect 6068 81460 6124 81500
rect 6164 81460 6173 81500
rect 6883 81460 6892 81500
rect 6932 81460 9772 81500
rect 9812 81460 9821 81500
rect 18499 81460 18508 81500
rect 18548 81460 19084 81500
rect 19124 81460 19133 81500
rect 19948 81416 19988 81712
rect 20039 81628 20048 81668
rect 20088 81628 20130 81668
rect 20170 81628 20212 81668
rect 20252 81628 20294 81668
rect 20334 81628 20376 81668
rect 20416 81628 20425 81668
rect 3139 81376 3148 81416
rect 3188 81376 8716 81416
rect 8756 81376 8765 81416
rect 19948 81376 20044 81416
rect 20084 81376 20093 81416
rect 2659 81292 2668 81332
rect 2708 81292 4300 81332
rect 4340 81292 4349 81332
rect 5347 81292 5356 81332
rect 5396 81292 8140 81332
rect 8180 81292 8189 81332
rect 18307 81292 18316 81332
rect 18356 81292 18604 81332
rect 18644 81292 18653 81332
rect 4963 81208 4972 81248
rect 5012 81208 6028 81248
rect 6068 81208 7660 81248
rect 7700 81208 7709 81248
rect 12940 81208 17932 81248
rect 17972 81208 17981 81248
rect 5827 81124 5836 81164
rect 5876 81124 5932 81164
rect 5972 81124 5981 81164
rect 8899 81124 8908 81164
rect 8948 81124 9484 81164
rect 9524 81124 9533 81164
rect 12940 81080 12980 81208
rect 2659 81040 2668 81080
rect 2708 81040 3628 81080
rect 3668 81040 3677 81080
rect 6403 81040 6412 81080
rect 6452 81040 12980 81080
rect 4675 80956 4684 80996
rect 4724 80956 6508 80996
rect 6548 80956 6557 80996
rect 643 80872 652 80912
rect 692 80872 940 80912
rect 980 80872 989 80912
rect 2371 80872 2380 80912
rect 2420 80872 2429 80912
rect 3679 80872 3688 80912
rect 3728 80872 3770 80912
rect 3810 80872 3852 80912
rect 3892 80872 3934 80912
rect 3974 80872 4016 80912
rect 4056 80872 4065 80912
rect 18799 80872 18808 80912
rect 18848 80872 18890 80912
rect 18930 80872 18972 80912
rect 19012 80872 19054 80912
rect 19094 80872 19136 80912
rect 19176 80872 19185 80912
rect 2380 80744 2420 80872
rect 2188 80704 2420 80744
rect 2851 80704 2860 80744
rect 2900 80704 4012 80744
rect 4052 80704 4061 80744
rect 6019 80704 6028 80744
rect 6068 80704 10156 80744
rect 10196 80704 10205 80744
rect 18307 80704 18316 80744
rect 18356 80704 19084 80744
rect 19124 80704 19133 80744
rect 1507 80536 1516 80576
rect 1556 80536 1804 80576
rect 1844 80536 1853 80576
rect 2188 80492 2228 80704
rect 11779 80620 11788 80660
rect 11828 80620 12076 80660
rect 12116 80620 16780 80660
rect 16820 80620 16829 80660
rect 2563 80536 2572 80576
rect 2612 80536 2668 80576
rect 2708 80536 2717 80576
rect 6499 80536 6508 80576
rect 6548 80536 6700 80576
rect 6740 80536 6749 80576
rect 9283 80536 9292 80576
rect 9332 80536 12748 80576
rect 12788 80536 13324 80576
rect 13364 80536 13373 80576
rect 17443 80536 17452 80576
rect 17492 80536 17548 80576
rect 17588 80536 17597 80576
rect 2064 80452 2092 80492
rect 2132 80452 8332 80492
rect 8372 80452 8381 80492
rect 12259 80452 12268 80492
rect 12308 80452 13036 80492
rect 13076 80452 13085 80492
rect 1603 80368 1612 80408
rect 1652 80368 5972 80408
rect 6019 80368 6028 80408
rect 6068 80368 7372 80408
rect 7412 80368 7421 80408
rect 11203 80368 11212 80408
rect 11252 80368 15628 80408
rect 15668 80368 15677 80408
rect 5155 80284 5164 80324
rect 5204 80284 5548 80324
rect 5588 80284 5597 80324
rect 2179 80200 2188 80240
rect 2228 80200 2956 80240
rect 2996 80200 3005 80240
rect 5932 80156 5972 80368
rect 6499 80200 6508 80240
rect 6548 80200 7372 80240
rect 7412 80200 9292 80240
rect 9332 80200 9341 80240
rect 4919 80116 4928 80156
rect 4968 80116 5010 80156
rect 5050 80116 5092 80156
rect 5132 80116 5174 80156
rect 5214 80116 5256 80156
rect 5296 80116 5305 80156
rect 5932 80116 6028 80156
rect 6068 80116 6077 80156
rect 8227 80116 8236 80156
rect 8276 80116 8812 80156
rect 8852 80116 8861 80156
rect 20039 80116 20048 80156
rect 20088 80116 20130 80156
rect 20170 80116 20212 80156
rect 20252 80116 20294 80156
rect 20334 80116 20376 80156
rect 20416 80116 20425 80156
rect 2947 80032 2956 80072
rect 2996 80032 3340 80072
rect 3380 80032 3389 80072
rect 7660 80032 12460 80072
rect 12500 80032 12509 80072
rect 2659 79948 2668 79988
rect 2708 79948 7276 79988
rect 7316 79948 7325 79988
rect 1680 79864 1708 79904
rect 1748 79864 1804 79904
rect 1844 79864 4396 79904
rect 4436 79864 4445 79904
rect 7660 79820 7700 80032
rect 11203 79948 11212 79988
rect 11252 79948 11980 79988
rect 12020 79948 12652 79988
rect 12692 79948 12701 79988
rect 7939 79864 7948 79904
rect 7988 79864 9676 79904
rect 9716 79864 9725 79904
rect 12355 79864 12364 79904
rect 12404 79864 12748 79904
rect 12788 79864 12797 79904
rect 13507 79864 13516 79904
rect 13556 79864 16492 79904
rect 16532 79864 16541 79904
rect 2755 79780 2764 79820
rect 2804 79780 7700 79820
rect 10627 79780 10636 79820
rect 10676 79780 13324 79820
rect 13364 79780 15820 79820
rect 15860 79780 17548 79820
rect 17588 79780 17597 79820
rect 3235 79696 3244 79736
rect 3284 79696 3724 79736
rect 3764 79696 3773 79736
rect 6979 79696 6988 79736
rect 7028 79696 7468 79736
rect 7508 79696 7517 79736
rect 11693 79696 11788 79736
rect 11828 79696 11837 79736
rect 11971 79696 11980 79736
rect 12020 79696 12940 79736
rect 12980 79696 12989 79736
rect 3523 79612 3532 79652
rect 3572 79612 4012 79652
rect 4052 79612 4061 79652
rect 6019 79612 6028 79652
rect 6068 79612 9676 79652
rect 9716 79612 9725 79652
rect 16483 79612 16492 79652
rect 16532 79612 19084 79652
rect 19124 79612 19133 79652
rect 355 79528 364 79568
rect 404 79528 3628 79568
rect 3668 79528 3677 79568
rect 5251 79528 5260 79568
rect 5300 79528 8812 79568
rect 8852 79528 8861 79568
rect 18604 79528 18796 79568
rect 18836 79528 18845 79568
rect 18979 79528 18988 79568
rect 19028 79528 19037 79568
rect 1795 79444 1804 79484
rect 1844 79444 3244 79484
rect 3284 79444 3293 79484
rect 3679 79360 3688 79400
rect 3728 79360 3770 79400
rect 3810 79360 3852 79400
rect 3892 79360 3934 79400
rect 3974 79360 4016 79400
rect 4056 79360 4065 79400
rect 1603 79276 1612 79316
rect 1652 79276 6508 79316
rect 6548 79276 6557 79316
rect 13891 79276 13900 79316
rect 13940 79276 15916 79316
rect 15956 79276 15965 79316
rect 5933 79192 6028 79232
rect 6068 79192 11788 79232
rect 11828 79192 11837 79232
rect 12163 79192 12172 79232
rect 12212 79192 16204 79232
rect 16244 79192 16253 79232
rect 18604 79148 18644 79528
rect 18988 79484 19028 79528
rect 18700 79444 19028 79484
rect 18700 79232 18740 79444
rect 18799 79360 18808 79400
rect 18848 79360 18890 79400
rect 18930 79360 18972 79400
rect 19012 79360 19054 79400
rect 19094 79360 19136 79400
rect 19176 79360 19185 79400
rect 18700 79192 18796 79232
rect 18836 79192 18845 79232
rect 2371 79108 2380 79148
rect 2420 79108 2668 79148
rect 2708 79108 2717 79148
rect 10915 79108 10924 79148
rect 10964 79108 15052 79148
rect 15092 79108 15101 79148
rect 18211 79108 18220 79148
rect 18260 79108 18316 79148
rect 18356 79108 18365 79148
rect 18604 79108 19084 79148
rect 19124 79108 19133 79148
rect 10531 79024 10540 79064
rect 10580 79024 15628 79064
rect 15668 79024 15677 79064
rect 3235 78940 3244 78980
rect 3284 78940 3436 78980
rect 3476 78940 3485 78980
rect 5357 78940 5452 78980
rect 5492 78940 5501 78980
rect 5827 78940 5836 78980
rect 5876 78940 9100 78980
rect 9140 78940 9149 78980
rect 9475 78940 9484 78980
rect 9524 78940 9868 78980
rect 9908 78940 9917 78980
rect 11203 78940 11212 78980
rect 11252 78940 16300 78980
rect 16340 78940 16349 78980
rect 10531 78856 10540 78896
rect 10580 78856 13900 78896
rect 13940 78856 13949 78896
rect 5539 78772 5548 78812
rect 5588 78772 10444 78812
rect 10484 78772 10493 78812
rect 12163 78772 12172 78812
rect 12212 78772 12460 78812
rect 12500 78772 12509 78812
rect 13507 78772 13516 78812
rect 13556 78772 13565 78812
rect 14851 78772 14860 78812
rect 14900 78772 15148 78812
rect 15188 78772 15197 78812
rect 20419 78772 20428 78812
rect 20468 78772 20812 78812
rect 20852 78772 20861 78812
rect 6787 78688 6796 78728
rect 6836 78688 9484 78728
rect 9524 78688 9533 78728
rect 10147 78688 10156 78728
rect 10196 78688 10924 78728
rect 10964 78688 10973 78728
rect 4919 78604 4928 78644
rect 4968 78604 5010 78644
rect 5050 78604 5092 78644
rect 5132 78604 5174 78644
rect 5214 78604 5256 78644
rect 5296 78604 5305 78644
rect 13516 78560 13556 78772
rect 17923 78604 17932 78644
rect 17972 78604 18892 78644
rect 18932 78604 18941 78644
rect 20039 78604 20048 78644
rect 20088 78604 20130 78644
rect 20170 78604 20212 78644
rect 20252 78604 20294 78644
rect 20334 78604 20376 78644
rect 20416 78604 20425 78644
rect 4387 78520 4396 78560
rect 4436 78520 7372 78560
rect 7412 78520 7421 78560
rect 11011 78520 11020 78560
rect 11060 78520 11069 78560
rect 13027 78520 13036 78560
rect 13076 78520 13556 78560
rect 16291 78520 16300 78560
rect 16340 78520 19084 78560
rect 19124 78520 19133 78560
rect 11020 78476 11060 78520
rect 6595 78436 6604 78476
rect 6644 78436 6796 78476
rect 6836 78436 6845 78476
rect 11020 78436 11212 78476
rect 11252 78436 11261 78476
rect 16963 78436 16972 78476
rect 17012 78436 17068 78476
rect 17108 78436 17117 78476
rect 18019 78352 18028 78392
rect 18068 78352 19372 78392
rect 19412 78352 20044 78392
rect 20084 78352 20093 78392
rect 3523 78268 3532 78308
rect 3572 78268 4012 78308
rect 4052 78268 4061 78308
rect 9091 78268 9100 78308
rect 9140 78268 9580 78308
rect 9620 78268 9629 78308
rect 10531 78268 10540 78308
rect 10580 78268 11980 78308
rect 12020 78268 13516 78308
rect 13556 78268 13565 78308
rect 13795 78268 13804 78308
rect 13844 78268 19180 78308
rect 19220 78268 19229 78308
rect 3427 78184 3436 78224
rect 3476 78184 3724 78224
rect 3764 78184 3773 78224
rect 4099 78184 4108 78224
rect 4148 78184 7948 78224
rect 7988 78184 7997 78224
rect 14851 78184 14860 78224
rect 14900 78184 15724 78224
rect 15764 78184 15773 78224
rect 8899 78100 8908 78140
rect 8948 78100 10444 78140
rect 10484 78100 10493 78140
rect 12355 78100 12364 78140
rect 12404 78100 13612 78140
rect 13652 78100 13661 78140
rect 14947 78100 14956 78140
rect 14996 78100 16588 78140
rect 16628 78100 16637 78140
rect 17443 78100 17452 78140
rect 17492 78100 20044 78140
rect 20084 78100 20093 78140
rect 5539 78016 5548 78056
rect 5588 78016 9100 78056
rect 9140 78016 9149 78056
rect 14083 78016 14092 78056
rect 14132 78016 16108 78056
rect 16148 78016 17644 78056
rect 17684 78016 18796 78056
rect 18836 78016 18845 78056
rect 19267 78016 19276 78056
rect 19316 78016 19564 78056
rect 19604 78016 19613 78056
rect 3679 77848 3688 77888
rect 3728 77848 3770 77888
rect 3810 77848 3852 77888
rect 3892 77848 3934 77888
rect 3974 77848 4016 77888
rect 4056 77848 4065 77888
rect 4291 77848 4300 77888
rect 4340 77848 7276 77888
rect 7316 77848 7325 77888
rect 18799 77848 18808 77888
rect 18848 77848 18890 77888
rect 18930 77848 18972 77888
rect 19012 77848 19054 77888
rect 19094 77848 19136 77888
rect 19176 77848 19185 77888
rect 3139 77680 3148 77720
rect 3188 77680 7948 77720
rect 7988 77680 7997 77720
rect 16291 77680 16300 77720
rect 16340 77680 17548 77720
rect 17588 77680 17597 77720
rect 2275 77512 2284 77552
rect 2324 77512 5356 77552
rect 5396 77512 5405 77552
rect 6691 77512 6700 77552
rect 6740 77512 7180 77552
rect 7220 77512 7229 77552
rect 2659 77428 2668 77468
rect 2708 77428 3820 77468
rect 3860 77428 3869 77468
rect 3916 77428 5260 77468
rect 5300 77428 5309 77468
rect 6883 77428 6892 77468
rect 6932 77428 8524 77468
rect 8564 77428 8573 77468
rect 10339 77428 10348 77468
rect 10388 77428 10540 77468
rect 10580 77428 10589 77468
rect 11779 77428 11788 77468
rect 11828 77428 12172 77468
rect 12212 77428 12221 77468
rect 14659 77428 14668 77468
rect 14708 77428 15724 77468
rect 15764 77428 15773 77468
rect 17539 77428 17548 77468
rect 17588 77428 17644 77468
rect 17684 77428 17693 77468
rect 3916 77216 3956 77428
rect 8323 77344 8332 77384
rect 8372 77344 9196 77384
rect 9236 77344 9868 77384
rect 9908 77344 9917 77384
rect 2851 77176 2860 77216
rect 2900 77176 3532 77216
rect 3572 77176 3956 77216
rect 10348 77260 10732 77300
rect 10772 77260 10781 77300
rect 4919 77092 4928 77132
rect 4968 77092 5010 77132
rect 5050 77092 5092 77132
rect 5132 77092 5174 77132
rect 5214 77092 5256 77132
rect 5296 77092 5305 77132
rect 2467 77008 2476 77048
rect 2516 77008 2572 77048
rect 2612 77008 2621 77048
rect 1603 76924 1612 76964
rect 1652 76924 1996 76964
rect 2036 76924 2045 76964
rect 2275 76924 2284 76964
rect 2324 76924 5548 76964
rect 5588 76924 5597 76964
rect 10157 76924 10252 76964
rect 10292 76924 10301 76964
rect 10348 76880 10388 77260
rect 20039 77092 20048 77132
rect 20088 77092 20130 77132
rect 20170 77092 20212 77132
rect 20252 77092 20294 77132
rect 20334 77092 20376 77132
rect 20416 77092 20425 77132
rect 10252 76840 10388 76880
rect 10636 76840 10732 76880
rect 10772 76840 10781 76880
rect 835 76756 844 76796
rect 884 76756 1132 76796
rect 1172 76756 1181 76796
rect 1507 76756 1516 76796
rect 1556 76756 1612 76796
rect 1652 76756 1661 76796
rect 2275 76756 2284 76796
rect 2324 76756 3244 76796
rect 3284 76756 6604 76796
rect 6644 76756 6653 76796
rect 10252 76712 10292 76840
rect 8419 76672 8428 76712
rect 8468 76672 10252 76712
rect 10292 76672 10301 76712
rect 2851 76588 2860 76628
rect 2900 76588 3148 76628
rect 3188 76588 3197 76628
rect 3523 76588 3532 76628
rect 3572 76588 3628 76628
rect 3668 76588 3677 76628
rect 10339 76588 10348 76628
rect 10388 76588 10444 76628
rect 10484 76588 10493 76628
rect 1219 76504 1228 76544
rect 1268 76504 6892 76544
rect 6932 76504 6941 76544
rect 10051 76420 10060 76460
rect 10100 76420 10109 76460
rect 2659 76336 2668 76376
rect 2708 76336 2956 76376
rect 2996 76336 3005 76376
rect 3679 76336 3688 76376
rect 3728 76336 3770 76376
rect 3810 76336 3852 76376
rect 3892 76336 3934 76376
rect 3974 76336 4016 76376
rect 4056 76336 4065 76376
rect 5357 76336 5452 76376
rect 5492 76336 5501 76376
rect 5933 76252 6028 76292
rect 6068 76252 6077 76292
rect 6211 76252 6220 76292
rect 6260 76252 8620 76292
rect 8660 76252 8669 76292
rect 10060 76208 10100 76420
rect 10636 76292 10676 76840
rect 17923 76756 17932 76796
rect 17972 76756 20140 76796
rect 20180 76756 20189 76796
rect 21196 76756 21388 76796
rect 21428 76756 21437 76796
rect 21196 76712 21236 76756
rect 14083 76672 14092 76712
rect 14132 76672 14476 76712
rect 14516 76672 14525 76712
rect 18307 76672 18316 76712
rect 18356 76672 18604 76712
rect 18644 76672 18653 76712
rect 21187 76672 21196 76712
rect 21236 76672 21245 76712
rect 10829 76588 10924 76628
rect 10964 76588 10973 76628
rect 20131 76588 20140 76628
rect 20180 76588 20524 76628
rect 20564 76588 20573 76628
rect 12749 76420 12844 76460
rect 12884 76420 12893 76460
rect 14851 76420 14860 76460
rect 14900 76420 15820 76460
rect 15860 76420 15869 76460
rect 14957 76336 15052 76376
rect 15092 76336 15101 76376
rect 18799 76336 18808 76376
rect 18848 76336 18890 76376
rect 18930 76336 18972 76376
rect 19012 76336 19054 76376
rect 19094 76336 19136 76376
rect 19176 76336 19185 76376
rect 10531 76252 10540 76292
rect 10580 76252 10676 76292
rect 13123 76252 13132 76292
rect 13172 76252 13324 76292
rect 13364 76252 13373 76292
rect 15715 76252 15724 76292
rect 15764 76252 16492 76292
rect 16532 76252 16541 76292
rect 5923 76168 5932 76208
rect 5972 76168 5981 76208
rect 10060 76168 14860 76208
rect 14900 76168 14909 76208
rect 5932 76124 5972 76168
rect 5932 76084 6220 76124
rect 6260 76084 6269 76124
rect 7853 76084 7948 76124
rect 7988 76084 7997 76124
rect 12835 76084 12844 76124
rect 12884 76084 13708 76124
rect 13748 76084 13757 76124
rect 1219 76000 1228 76040
rect 1268 76000 2860 76040
rect 2900 76000 2909 76040
rect 14755 76000 14764 76040
rect 14804 76000 15820 76040
rect 15860 76000 15869 76040
rect 18307 76000 18316 76040
rect 18356 76000 20140 76040
rect 20180 76000 20189 76040
rect 739 75916 748 75956
rect 788 75916 5260 75956
rect 5300 75916 5309 75956
rect 6893 75916 6988 75956
rect 7028 75916 7037 75956
rect 10723 75916 10732 75956
rect 10772 75916 13612 75956
rect 13652 75916 13661 75956
rect 14179 75916 14188 75956
rect 14228 75916 14237 75956
rect 17059 75916 17068 75956
rect 17108 75916 17356 75956
rect 17396 75916 17405 75956
rect 20611 75916 20620 75956
rect 20660 75916 20908 75956
rect 20948 75916 20957 75956
rect 3523 75832 3532 75872
rect 3572 75832 3628 75872
rect 3668 75832 3677 75872
rect 1123 75748 1132 75788
rect 1172 75748 4684 75788
rect 4724 75748 4733 75788
rect 13123 75748 13132 75788
rect 13172 75748 13996 75788
rect 14036 75748 14045 75788
rect 4919 75580 4928 75620
rect 4968 75580 5010 75620
rect 5050 75580 5092 75620
rect 5132 75580 5174 75620
rect 5214 75580 5256 75620
rect 5296 75580 5305 75620
rect 6211 75580 6220 75620
rect 6260 75580 13804 75620
rect 13844 75580 13853 75620
rect 355 75496 364 75536
rect 404 75496 556 75536
rect 596 75496 605 75536
rect 14188 75452 14228 75916
rect 17453 75748 17548 75788
rect 17588 75748 17597 75788
rect 20419 75748 20428 75788
rect 20468 75748 20564 75788
rect 20039 75580 20048 75620
rect 20088 75580 20130 75620
rect 20170 75580 20212 75620
rect 20252 75580 20294 75620
rect 20334 75580 20376 75620
rect 20416 75580 20425 75620
rect 20524 75452 20564 75748
rect 4771 75412 4780 75452
rect 4820 75412 10060 75452
rect 10100 75412 10109 75452
rect 14188 75412 14324 75452
rect 20419 75412 20428 75452
rect 20468 75412 20564 75452
rect 7939 75328 7948 75368
rect 7988 75328 8428 75368
rect 8468 75328 8477 75368
rect 4771 75244 4780 75284
rect 4820 75244 4876 75284
rect 4916 75244 4925 75284
rect 8227 75244 8236 75284
rect 8276 75244 8620 75284
rect 8660 75244 8669 75284
rect 5731 75160 5740 75200
rect 5780 75160 6796 75200
rect 6836 75160 6845 75200
rect 14284 75116 14324 75412
rect 6893 75076 6988 75116
rect 7028 75076 7037 75116
rect 13229 75076 13324 75116
rect 13364 75076 13373 75116
rect 14275 75076 14284 75116
rect 14324 75076 14333 75116
rect 7267 74992 7276 75032
rect 7316 74992 7948 75032
rect 7988 74992 7997 75032
rect 18499 74992 18508 75032
rect 18548 74992 18796 75032
rect 18836 74992 18845 75032
rect 3679 74824 3688 74864
rect 3728 74824 3770 74864
rect 3810 74824 3852 74864
rect 3892 74824 3934 74864
rect 3974 74824 4016 74864
rect 4056 74824 4065 74864
rect 18799 74824 18808 74864
rect 18848 74824 18890 74864
rect 18930 74824 18972 74864
rect 19012 74824 19054 74864
rect 19094 74824 19136 74864
rect 19176 74824 19185 74864
rect 5443 74740 5452 74780
rect 5492 74740 8908 74780
rect 8948 74740 8957 74780
rect 5251 74656 5260 74696
rect 5300 74656 7660 74696
rect 7700 74656 7709 74696
rect 12739 74656 12748 74696
rect 12788 74656 16108 74696
rect 16148 74656 16157 74696
rect 18979 74656 18988 74696
rect 19028 74656 19372 74696
rect 19412 74656 19421 74696
rect 5443 74572 5452 74612
rect 5492 74572 7084 74612
rect 7124 74572 7133 74612
rect 7939 74572 7948 74612
rect 7988 74572 8908 74612
rect 8948 74572 8957 74612
rect 14179 74572 14188 74612
rect 14228 74572 19084 74612
rect 19124 74572 19133 74612
rect 5827 74488 5836 74528
rect 5876 74488 6220 74528
rect 6260 74488 6269 74528
rect 13123 74488 13132 74528
rect 13172 74488 13324 74528
rect 13364 74488 13373 74528
rect 14083 74488 14092 74528
rect 14132 74488 16108 74528
rect 16148 74488 16157 74528
rect 16387 74488 16396 74528
rect 16436 74488 17836 74528
rect 17876 74488 17885 74528
rect 547 74404 556 74444
rect 596 74404 5932 74444
rect 5972 74404 5981 74444
rect 12643 74404 12652 74444
rect 12692 74404 12748 74444
rect 12788 74404 12797 74444
rect 14467 74404 14476 74444
rect 14516 74404 15340 74444
rect 15380 74404 17452 74444
rect 17492 74404 17501 74444
rect 1325 74320 1420 74360
rect 1460 74320 1469 74360
rect 3437 74320 3532 74360
rect 3572 74320 3581 74360
rect 5155 74320 5164 74360
rect 5204 74320 5452 74360
rect 5492 74320 5501 74360
rect 1123 74236 1132 74276
rect 1172 74236 7660 74276
rect 7700 74236 7709 74276
rect 13795 74236 13804 74276
rect 13844 74236 14188 74276
rect 14228 74236 14237 74276
rect 20419 74236 20428 74276
rect 20468 74236 20564 74276
rect 1315 74152 1324 74192
rect 1364 74152 1420 74192
rect 1460 74152 1469 74192
rect 3427 74152 3436 74192
rect 3476 74152 3916 74192
rect 3956 74152 3965 74192
rect 4771 74152 4780 74192
rect 4820 74152 8236 74192
rect 8276 74152 8285 74192
rect 1987 74068 1996 74108
rect 2036 74068 2324 74108
rect 4919 74068 4928 74108
rect 4968 74068 5010 74108
rect 5050 74068 5092 74108
rect 5132 74068 5174 74108
rect 5214 74068 5256 74108
rect 5296 74068 5305 74108
rect 5923 74068 5932 74108
rect 5972 74068 6316 74108
rect 6356 74068 6365 74108
rect 13891 74068 13900 74108
rect 13940 74068 14092 74108
rect 14132 74068 14141 74108
rect 20039 74068 20048 74108
rect 20088 74068 20130 74108
rect 20170 74068 20212 74108
rect 20252 74068 20294 74108
rect 20334 74068 20376 74108
rect 20416 74068 20425 74108
rect 269 73816 364 73856
rect 404 73816 413 73856
rect 2284 73604 2324 74068
rect 4387 73984 4396 74024
rect 4436 73984 6988 74024
rect 7028 73984 7037 74024
rect 20524 73940 20564 74236
rect 4291 73900 4300 73940
rect 4340 73900 5836 73940
rect 5876 73900 5885 73940
rect 12547 73900 12556 73940
rect 12596 73900 16012 73940
rect 16052 73900 16396 73940
rect 16436 73900 16445 73940
rect 19651 73900 19660 73940
rect 19700 73900 20044 73940
rect 20084 73900 20093 73940
rect 20419 73900 20428 73940
rect 20468 73900 20564 73940
rect 3523 73816 3532 73856
rect 3572 73816 9484 73856
rect 9524 73816 9533 73856
rect 13123 73816 13132 73856
rect 13172 73816 13181 73856
rect 3043 73648 3052 73688
rect 3092 73648 3244 73688
rect 3284 73648 3293 73688
rect 4291 73648 4300 73688
rect 4340 73648 4349 73688
rect 4963 73648 4972 73688
rect 5012 73648 9292 73688
rect 9332 73648 9341 73688
rect 10339 73648 10348 73688
rect 10388 73648 11116 73688
rect 11156 73648 11165 73688
rect 4300 73604 4340 73648
rect 13132 73604 13172 73816
rect 13891 73732 13900 73772
rect 13940 73732 18316 73772
rect 18356 73732 18365 73772
rect 2275 73564 2284 73604
rect 2324 73564 2333 73604
rect 4291 73564 4300 73604
rect 4340 73564 4351 73604
rect 6595 73564 6604 73604
rect 6644 73564 7084 73604
rect 7124 73564 7133 73604
rect 12076 73564 12844 73604
rect 12884 73564 12893 73604
rect 13027 73564 13036 73604
rect 13076 73564 13172 73604
rect 2947 73480 2956 73520
rect 2996 73480 3091 73520
rect 6019 73480 6028 73520
rect 6068 73480 6412 73520
rect 6452 73480 6461 73520
rect 6787 73480 6796 73520
rect 6836 73480 6845 73520
rect 8995 73480 9004 73520
rect 9044 73480 9100 73520
rect 9140 73480 9149 73520
rect 1987 73420 1996 73460
rect 2036 73436 2045 73460
rect 2036 73420 2188 73436
rect 1996 73396 2188 73420
rect 2228 73396 2237 73436
rect 2371 73420 2380 73460
rect 2420 73420 2429 73460
rect 6796 73436 6836 73480
rect 12076 73436 12116 73564
rect 14957 73480 15052 73520
rect 15092 73480 15101 73520
rect 16195 73480 16204 73520
rect 16244 73480 17164 73520
rect 17204 73480 17213 73520
rect 18979 73480 18988 73520
rect 19028 73480 19037 73520
rect 19171 73480 19180 73520
rect 19220 73480 19229 73520
rect 18988 73436 19028 73480
rect 2380 73352 2420 73420
rect 6796 73396 7180 73436
rect 7220 73396 7229 73436
rect 11587 73396 11596 73436
rect 11636 73396 11884 73436
rect 11924 73396 11933 73436
rect 12067 73396 12076 73436
rect 12116 73396 12125 73436
rect 18604 73396 19028 73436
rect 19180 73436 19220 73480
rect 19180 73396 19700 73436
rect 20611 73396 20620 73436
rect 20660 73396 21196 73436
rect 21236 73396 21245 73436
rect 18604 73352 18644 73396
rect 1987 73312 1996 73352
rect 2036 73312 2420 73352
rect 3679 73312 3688 73352
rect 3728 73312 3770 73352
rect 3810 73312 3852 73352
rect 3892 73312 3934 73352
rect 3974 73312 4016 73352
rect 4056 73312 4065 73352
rect 8419 73312 8428 73352
rect 8468 73312 9196 73352
rect 9236 73312 9245 73352
rect 10051 73312 10060 73352
rect 10100 73312 12844 73352
rect 12884 73312 13324 73352
rect 13364 73312 13373 73352
rect 18595 73312 18604 73352
rect 18644 73312 18653 73352
rect 18799 73312 18808 73352
rect 18848 73312 18890 73352
rect 18930 73312 18972 73352
rect 19012 73312 19054 73352
rect 19094 73312 19136 73352
rect 19176 73312 19185 73352
rect 8227 73228 8236 73268
rect 8276 73228 15244 73268
rect 15284 73228 15293 73268
rect 11971 73144 11980 73184
rect 12020 73144 12652 73184
rect 12692 73144 12701 73184
rect 12931 73144 12940 73184
rect 12980 73144 13708 73184
rect 13748 73144 13757 73184
rect 2477 73060 2572 73100
rect 2612 73060 2621 73100
rect 5731 73060 5740 73100
rect 5780 73060 12844 73100
rect 12884 73060 12893 73100
rect 8131 72976 8140 73016
rect 8180 72976 8812 73016
rect 8852 72976 8861 73016
rect 2947 72892 2956 72932
rect 2996 72892 6604 72932
rect 6644 72892 6653 72932
rect 8323 72892 8332 72932
rect 8372 72892 8620 72932
rect 8660 72892 8669 72932
rect 15907 72892 15916 72932
rect 15956 72892 16012 72932
rect 16052 72892 16061 72932
rect 19660 72848 19700 73396
rect 19756 72892 19852 72932
rect 19892 72892 19901 72932
rect 19651 72808 19660 72848
rect 19700 72808 19709 72848
rect 5251 72724 5260 72764
rect 5300 72724 6988 72764
rect 7028 72724 7037 72764
rect 7267 72724 7276 72764
rect 7316 72724 8332 72764
rect 8372 72724 8381 72764
rect 17539 72724 17548 72764
rect 17588 72724 19084 72764
rect 19124 72724 19133 72764
rect 19756 72680 19796 72892
rect 20419 72808 20428 72848
rect 20468 72808 21100 72848
rect 21140 72808 21149 72848
rect 19843 72724 19852 72764
rect 19892 72724 20044 72764
rect 20084 72724 20093 72764
rect 18307 72640 18316 72680
rect 18356 72640 19796 72680
rect 19948 72640 20524 72680
rect 20564 72640 20573 72680
rect 4919 72556 4928 72596
rect 4968 72556 5010 72596
rect 5050 72556 5092 72596
rect 5132 72556 5174 72596
rect 5214 72556 5256 72596
rect 5296 72556 5305 72596
rect 18019 72556 18028 72596
rect 18068 72556 18077 72596
rect 1027 72472 1036 72512
rect 1076 72472 2860 72512
rect 2900 72472 2909 72512
rect 3235 72472 3244 72512
rect 3284 72472 4204 72512
rect 4244 72472 4253 72512
rect 3139 72388 3148 72428
rect 3188 72388 3340 72428
rect 3380 72388 3389 72428
rect 14947 72388 14956 72428
rect 14996 72388 15244 72428
rect 15284 72388 15293 72428
rect 4109 72304 4204 72344
rect 4244 72304 4253 72344
rect 2947 72220 2956 72260
rect 2996 72220 3532 72260
rect 3572 72220 5932 72260
rect 5972 72220 5981 72260
rect 11491 72220 11500 72260
rect 11540 72220 12844 72260
rect 12884 72220 12893 72260
rect 4579 72136 4588 72176
rect 4628 72136 5836 72176
rect 5876 72136 5885 72176
rect 9859 72136 9868 72176
rect 9908 72136 9964 72176
rect 10004 72136 10013 72176
rect 18028 72092 18068 72556
rect 19948 72428 19988 72640
rect 20039 72556 20048 72596
rect 20088 72556 20130 72596
rect 20170 72556 20212 72596
rect 20252 72556 20294 72596
rect 20334 72556 20376 72596
rect 20416 72556 20425 72596
rect 18307 72388 18316 72428
rect 18356 72388 18508 72428
rect 18548 72388 18557 72428
rect 19948 72388 20044 72428
rect 20084 72388 20093 72428
rect 1613 72052 1708 72092
rect 1748 72052 1757 72092
rect 3619 72052 3628 72092
rect 3668 72052 6892 72092
rect 6932 72052 6941 72092
rect 9283 72052 9292 72092
rect 9332 72052 9341 72092
rect 17635 72052 17644 72092
rect 17684 72052 18068 72092
rect 18595 72052 18604 72092
rect 18644 72052 18796 72092
rect 18836 72052 18845 72092
rect 5443 71968 5452 72008
rect 5492 71968 6700 72008
rect 6740 71968 6749 72008
rect 9292 71840 9332 72052
rect 11587 71968 11596 72008
rect 11636 71968 12076 72008
rect 12116 71968 12125 72008
rect 3679 71800 3688 71840
rect 3728 71800 3770 71840
rect 3810 71800 3852 71840
rect 3892 71800 3934 71840
rect 3974 71800 4016 71840
rect 4056 71800 4065 71840
rect 9292 71800 9484 71840
rect 9524 71800 9533 71840
rect 18799 71800 18808 71840
rect 18848 71800 18890 71840
rect 18930 71800 18972 71840
rect 19012 71800 19054 71840
rect 19094 71800 19136 71840
rect 19176 71800 19185 71840
rect 2093 71716 2188 71756
rect 2228 71716 2237 71756
rect 2947 71716 2956 71756
rect 2996 71716 3091 71756
rect 15619 71716 15628 71756
rect 15668 71716 15724 71756
rect 15764 71716 15773 71756
rect 3523 71632 3532 71672
rect 3572 71632 3628 71672
rect 3668 71632 3677 71672
rect 18499 71632 18508 71672
rect 18548 71632 18892 71672
rect 18932 71632 18941 71672
rect 5635 71548 5644 71588
rect 5684 71548 10060 71588
rect 10100 71548 10109 71588
rect 15907 71548 15916 71588
rect 15956 71548 16396 71588
rect 16436 71548 16445 71588
rect 17155 71548 17164 71588
rect 17204 71548 19948 71588
rect 19988 71548 19997 71588
rect 2851 71464 2860 71504
rect 2900 71464 5068 71504
rect 5108 71464 5117 71504
rect 5251 71464 5260 71504
rect 5300 71464 7372 71504
rect 7412 71464 7421 71504
rect 7843 71464 7852 71504
rect 7892 71464 7948 71504
rect 7988 71464 7997 71504
rect 9667 71464 9676 71504
rect 9716 71464 17260 71504
rect 17300 71464 17309 71504
rect 1987 71380 1996 71420
rect 2036 71380 12844 71420
rect 12884 71380 12893 71420
rect 14563 71380 14572 71420
rect 14612 71380 14956 71420
rect 14996 71380 15005 71420
rect 2275 71296 2284 71336
rect 2324 71296 7276 71336
rect 7316 71296 7325 71336
rect 11779 71296 11788 71336
rect 11828 71296 11980 71336
rect 12020 71296 12029 71336
rect 14851 71296 14860 71336
rect 14900 71296 15820 71336
rect 15860 71296 15869 71336
rect 16387 71296 16396 71336
rect 16436 71296 17932 71336
rect 17972 71296 17981 71336
rect 14477 71212 14572 71252
rect 14612 71212 14621 71252
rect 15043 71212 15052 71252
rect 15092 71212 15532 71252
rect 15572 71212 15581 71252
rect 17827 71212 17836 71252
rect 17876 71212 18028 71252
rect 18068 71212 18077 71252
rect 1795 71128 1804 71168
rect 1844 71128 12980 71168
rect 15427 71128 15436 71168
rect 15476 71128 16684 71168
rect 16724 71128 16733 71168
rect 12940 71084 12980 71128
rect 4919 71044 4928 71084
rect 4968 71044 5010 71084
rect 5050 71044 5092 71084
rect 5132 71044 5174 71084
rect 5214 71044 5256 71084
rect 5296 71044 5305 71084
rect 12940 71044 13420 71084
rect 13460 71044 13469 71084
rect 20039 71044 20048 71084
rect 20088 71044 20130 71084
rect 20170 71044 20212 71084
rect 20252 71044 20294 71084
rect 20334 71044 20376 71084
rect 20416 71044 20425 71084
rect 1219 70960 1228 71000
rect 1268 70960 9772 71000
rect 9812 70960 9821 71000
rect 4771 70876 4780 70916
rect 4820 70876 4972 70916
rect 5012 70876 5021 70916
rect 5155 70876 5164 70916
rect 5204 70876 5548 70916
rect 5588 70876 5597 70916
rect 6595 70876 6604 70916
rect 6644 70876 7660 70916
rect 7700 70876 7709 70916
rect 13123 70876 13132 70916
rect 13172 70876 17548 70916
rect 17588 70876 17597 70916
rect 6979 70792 6988 70832
rect 7028 70792 7180 70832
rect 7220 70792 7229 70832
rect 10627 70792 10636 70832
rect 10676 70792 12460 70832
rect 12500 70792 12509 70832
rect 13027 70792 13036 70832
rect 13076 70792 16012 70832
rect 16052 70792 16061 70832
rect 653 70708 748 70748
rect 788 70708 797 70748
rect 4771 70708 4780 70748
rect 4820 70708 4876 70748
rect 4916 70708 4925 70748
rect 6499 70708 6508 70748
rect 6548 70708 7372 70748
rect 7412 70708 7564 70748
rect 7604 70708 7613 70748
rect 17932 70708 18508 70748
rect 18548 70708 18557 70748
rect 17932 70664 17972 70708
rect 3715 70624 3724 70664
rect 3764 70624 3916 70664
rect 3956 70624 4300 70664
rect 4340 70624 4349 70664
rect 9571 70624 9580 70664
rect 9620 70624 10060 70664
rect 10100 70624 10109 70664
rect 15043 70624 15052 70664
rect 15092 70624 17972 70664
rect 17932 70580 17972 70624
rect 5453 70540 5548 70580
rect 5588 70540 5597 70580
rect 6125 70540 6220 70580
rect 6260 70540 6269 70580
rect 7277 70540 7372 70580
rect 7412 70540 7421 70580
rect 8813 70540 8908 70580
rect 8948 70540 8957 70580
rect 9581 70540 9676 70580
rect 9716 70540 9725 70580
rect 15619 70540 15628 70580
rect 15668 70540 15724 70580
rect 15764 70540 15773 70580
rect 15907 70540 15916 70580
rect 15956 70540 16588 70580
rect 16628 70540 16637 70580
rect 17923 70540 17932 70580
rect 17972 70540 17981 70580
rect 3427 70456 3436 70496
rect 3476 70456 3628 70496
rect 3668 70456 3677 70496
rect 3907 70456 3916 70496
rect 3956 70456 5644 70496
rect 5684 70456 5693 70496
rect 10051 70456 10060 70496
rect 10100 70456 10252 70496
rect 10292 70456 10301 70496
rect 12643 70456 12652 70496
rect 12692 70456 16300 70496
rect 16340 70456 16349 70496
rect 17923 70456 17932 70496
rect 17972 70456 18892 70496
rect 18932 70456 18941 70496
rect 11011 70372 11020 70412
rect 11060 70372 13612 70412
rect 13652 70372 13661 70412
rect 16579 70372 16588 70412
rect 16628 70372 17164 70412
rect 17204 70372 17213 70412
rect 3679 70288 3688 70328
rect 3728 70288 3770 70328
rect 3810 70288 3852 70328
rect 3892 70288 3934 70328
rect 3974 70288 4016 70328
rect 4056 70288 4065 70328
rect 18799 70288 18808 70328
rect 18848 70288 18890 70328
rect 18930 70288 18972 70328
rect 19012 70288 19054 70328
rect 19094 70288 19136 70328
rect 19176 70288 19185 70328
rect 7651 70204 7660 70244
rect 7700 70204 7948 70244
rect 7988 70204 7997 70244
rect 17443 70120 17452 70160
rect 17492 70120 19084 70160
rect 19124 70120 19133 70160
rect 1987 70036 1996 70076
rect 2036 70036 2764 70076
rect 2804 70036 5836 70076
rect 5876 70036 5885 70076
rect 10243 70036 10252 70076
rect 10292 70036 10540 70076
rect 10580 70036 10589 70076
rect 17251 70036 17260 70076
rect 17300 70036 19276 70076
rect 19316 70036 19325 70076
rect 2371 69952 2380 69992
rect 2420 69952 19756 69992
rect 19796 69952 19805 69992
rect 2947 69868 2956 69908
rect 2996 69868 4300 69908
rect 4340 69868 4349 69908
rect 20323 69784 20332 69824
rect 20372 69784 20620 69824
rect 20660 69784 20669 69824
rect 5155 69700 5164 69740
rect 5204 69700 5548 69740
rect 5588 69700 5597 69740
rect 11395 69700 11404 69740
rect 11444 69700 20140 69740
rect 20180 69700 20189 69740
rect 20419 69700 20428 69740
rect 20468 69700 20524 69740
rect 20564 69700 20573 69740
rect 4919 69532 4928 69572
rect 4968 69532 5010 69572
rect 5050 69532 5092 69572
rect 5132 69532 5174 69572
rect 5214 69532 5256 69572
rect 5296 69532 5305 69572
rect 20039 69532 20048 69572
rect 20088 69532 20130 69572
rect 20170 69532 20212 69572
rect 20252 69532 20294 69572
rect 20334 69532 20376 69572
rect 20416 69532 20425 69572
rect 5260 69448 8620 69488
rect 8660 69448 8669 69488
rect 5260 69404 5300 69448
rect 5251 69364 5260 69404
rect 5300 69364 5309 69404
rect 7469 69364 7564 69404
rect 7604 69364 7613 69404
rect 9283 69364 9292 69404
rect 9332 69364 11788 69404
rect 11828 69364 11837 69404
rect 5539 69280 5548 69320
rect 5588 69280 5597 69320
rect 5827 69280 5836 69320
rect 5876 69280 6988 69320
rect 7028 69280 8236 69320
rect 8276 69280 8285 69320
rect 10060 69280 10252 69320
rect 10292 69280 10301 69320
rect 16483 69280 16492 69320
rect 16532 69280 16588 69320
rect 16628 69280 16637 69320
rect 2755 69196 2764 69236
rect 2804 69196 2860 69236
rect 2900 69196 2909 69236
rect 3331 69196 3340 69236
rect 3380 69196 3532 69236
rect 3572 69196 3628 69236
rect 3668 69196 3677 69236
rect 5548 69152 5588 69280
rect 451 69112 460 69152
rect 500 69112 1708 69152
rect 1748 69112 1757 69152
rect 2659 69112 2668 69152
rect 2708 69112 2860 69152
rect 2900 69112 2909 69152
rect 5548 69112 5740 69152
rect 5780 69112 5789 69152
rect 10060 68984 10100 69280
rect 17059 69196 17068 69236
rect 17108 69196 17204 69236
rect 10339 69112 10348 69152
rect 10388 69112 11884 69152
rect 11924 69112 11933 69152
rect 13229 69112 13324 69152
rect 13364 69112 13373 69152
rect 14179 69112 14188 69152
rect 14228 69112 14476 69152
rect 14516 69112 14525 69152
rect 16867 69028 16876 69068
rect 16916 69028 17068 69068
rect 17108 69028 17117 69068
rect 17164 68984 17204 69196
rect 20611 69112 20620 69152
rect 20660 69112 20852 69152
rect 1133 68944 1228 68984
rect 1268 68944 1277 68984
rect 9868 68944 10100 68984
rect 13987 68944 13996 68984
rect 14036 68944 14188 68984
rect 14228 68944 14237 68984
rect 16876 68944 17204 68984
rect 19075 68944 19084 68984
rect 19124 68944 20620 68984
rect 20660 68944 20669 68984
rect 2467 68776 2476 68816
rect 2516 68776 3436 68816
rect 3476 68776 3485 68816
rect 3679 68776 3688 68816
rect 3728 68776 3770 68816
rect 3810 68776 3852 68816
rect 3892 68776 3934 68816
rect 3974 68776 4016 68816
rect 4056 68776 4065 68816
rect 4675 68776 4684 68816
rect 4724 68776 4876 68816
rect 4916 68776 4925 68816
rect 9475 68608 9484 68648
rect 9524 68608 9676 68648
rect 9716 68608 9725 68648
rect 7267 68524 7276 68564
rect 7316 68524 7852 68564
rect 7892 68524 7901 68564
rect 1795 68440 1804 68480
rect 1844 68440 2284 68480
rect 2324 68440 2333 68480
rect 4003 68440 4012 68480
rect 4052 68440 4780 68480
rect 4820 68440 4829 68480
rect 6499 68440 6508 68480
rect 6548 68440 7180 68480
rect 7220 68440 7229 68480
rect 7459 68440 7468 68480
rect 7508 68440 8716 68480
rect 8756 68440 8765 68480
rect 1603 68356 1612 68396
rect 1652 68356 2188 68396
rect 2228 68356 2237 68396
rect 5443 68356 5452 68396
rect 5492 68356 7660 68396
rect 7700 68356 7709 68396
rect 3907 68272 3916 68312
rect 3956 68272 5644 68312
rect 5684 68272 9004 68312
rect 9044 68272 9053 68312
rect 9868 68228 9908 68944
rect 16876 68900 16916 68944
rect 16867 68860 16876 68900
rect 16916 68860 16925 68900
rect 20812 68816 20852 69112
rect 18799 68776 18808 68816
rect 18848 68776 18890 68816
rect 18930 68776 18972 68816
rect 19012 68776 19054 68816
rect 19094 68776 19136 68816
rect 19176 68776 19185 68816
rect 20803 68776 20812 68816
rect 20852 68776 20861 68816
rect 10051 68608 10060 68648
rect 10100 68608 14380 68648
rect 14420 68608 14429 68648
rect 18307 68608 18316 68648
rect 18356 68608 18796 68648
rect 18836 68608 18845 68648
rect 19747 68608 19756 68648
rect 19796 68608 19805 68648
rect 19756 68480 19796 68608
rect 19267 68440 19276 68480
rect 19316 68440 19796 68480
rect 10060 68356 13420 68396
rect 13460 68356 13996 68396
rect 14036 68356 14045 68396
rect 1315 68188 1324 68228
rect 1364 68188 7948 68228
rect 7988 68188 7997 68228
rect 8141 68188 8236 68228
rect 8276 68188 8285 68228
rect 9859 68188 9868 68228
rect 9908 68188 9917 68228
rect 10060 68144 10100 68356
rect 12931 68272 12940 68312
rect 12980 68272 13996 68312
rect 14036 68272 14045 68312
rect 2947 68104 2956 68144
rect 2996 68104 3340 68144
rect 3380 68104 3389 68144
rect 10051 68104 10060 68144
rect 10100 68104 10109 68144
rect 4919 68020 4928 68060
rect 4968 68020 5010 68060
rect 5050 68020 5092 68060
rect 5132 68020 5174 68060
rect 5214 68020 5256 68060
rect 5296 68020 5305 68060
rect 4099 67852 4108 67892
rect 4148 67852 4780 67892
rect 4820 67852 4829 67892
rect 13420 67808 13460 68272
rect 20707 68104 20716 68144
rect 20756 68104 21004 68144
rect 21044 68104 21053 68144
rect 20039 68020 20048 68060
rect 20088 68020 20130 68060
rect 20170 68020 20212 68060
rect 20252 68020 20294 68060
rect 20334 68020 20376 68060
rect 20416 68020 20425 68060
rect 17443 67936 17452 67976
rect 17492 67936 17740 67976
rect 17780 67936 17789 67976
rect 20419 67852 20428 67892
rect 20468 67852 20524 67892
rect 20564 67852 20573 67892
rect 5347 67768 5356 67808
rect 5396 67768 5548 67808
rect 5588 67768 5597 67808
rect 13411 67768 13420 67808
rect 13460 67768 13469 67808
rect 4483 67684 4492 67724
rect 4532 67684 4876 67724
rect 4916 67684 4925 67724
rect 1325 67600 1420 67640
rect 1460 67600 1469 67640
rect 3331 67600 3340 67640
rect 3380 67600 3532 67640
rect 3572 67600 3581 67640
rect 6787 67600 6796 67640
rect 6836 67600 7372 67640
rect 7412 67600 7421 67640
rect 10243 67516 10252 67556
rect 10292 67516 10348 67556
rect 10388 67516 10397 67556
rect 2083 67432 2092 67472
rect 2132 67432 2188 67472
rect 2228 67432 2237 67472
rect 3523 67432 3532 67472
rect 3572 67432 4012 67472
rect 4052 67432 4061 67472
rect 6787 67432 6796 67472
rect 6836 67432 6988 67472
rect 7028 67432 7037 67472
rect 16675 67432 16684 67472
rect 16724 67432 17260 67472
rect 17300 67432 17309 67472
rect 3679 67264 3688 67304
rect 3728 67264 3770 67304
rect 3810 67264 3852 67304
rect 3892 67264 3934 67304
rect 3974 67264 4016 67304
rect 4056 67264 4065 67304
rect 18799 67264 18808 67304
rect 18848 67264 18890 67304
rect 18930 67264 18972 67304
rect 19012 67264 19054 67304
rect 19094 67264 19136 67304
rect 19176 67264 19185 67304
rect 1795 67180 1804 67220
rect 1844 67180 13708 67220
rect 13748 67180 13757 67220
rect 2083 67096 2092 67136
rect 2132 67096 8908 67136
rect 8948 67096 8957 67136
rect 13037 67096 13132 67136
rect 13172 67096 13181 67136
rect 18403 67096 18412 67136
rect 18452 67096 18796 67136
rect 18836 67096 18845 67136
rect 3523 67012 3532 67052
rect 3572 67012 3628 67052
rect 3668 67012 3677 67052
rect 1325 66928 1420 66968
rect 1460 66928 1469 66968
rect 4867 66928 4876 66968
rect 4916 66928 5548 66968
rect 5588 66928 6028 66968
rect 6068 66928 6077 66968
rect 11491 66928 11500 66968
rect 11540 66928 11692 66968
rect 11732 66928 11741 66968
rect 1901 66844 1996 66884
rect 2036 66844 2045 66884
rect 2659 66844 2668 66884
rect 2708 66844 6220 66884
rect 6260 66844 6269 66884
rect 15043 66844 15052 66884
rect 15092 66844 15284 66884
rect 16867 66844 16876 66884
rect 16916 66844 17164 66884
rect 17204 66844 17213 66884
rect 15244 66800 15284 66844
rect 3811 66760 3820 66800
rect 3860 66760 9676 66800
rect 9716 66760 9725 66800
rect 15235 66760 15244 66800
rect 15284 66760 15293 66800
rect 1987 66676 1996 66716
rect 2036 66676 6604 66716
rect 6644 66676 6653 66716
rect 20131 66676 20140 66716
rect 20180 66676 20620 66716
rect 20660 66676 20669 66716
rect 7363 66592 7372 66632
rect 7412 66592 8524 66632
rect 8564 66592 8573 66632
rect 4919 66508 4928 66548
rect 4968 66508 5010 66548
rect 5050 66508 5092 66548
rect 5132 66508 5174 66548
rect 5214 66508 5256 66548
rect 5296 66508 5305 66548
rect 5347 66508 5356 66548
rect 5396 66508 11692 66548
rect 11732 66508 11741 66548
rect 14371 66508 14380 66548
rect 14420 66508 17356 66548
rect 17396 66508 17740 66548
rect 17780 66508 17789 66548
rect 20039 66508 20048 66548
rect 20088 66508 20130 66548
rect 20170 66508 20212 66548
rect 20252 66508 20294 66548
rect 20334 66508 20376 66548
rect 20416 66508 20425 66548
rect 6883 66424 6892 66464
rect 6932 66424 7316 66464
rect 1699 66256 1708 66296
rect 1748 66256 1804 66296
rect 1844 66256 1853 66296
rect 2659 66256 2668 66296
rect 2708 66256 3340 66296
rect 3380 66256 3389 66296
rect 7276 66212 7316 66424
rect 12163 66340 12172 66380
rect 12212 66340 12460 66380
rect 12500 66340 12509 66380
rect 15427 66256 15436 66296
rect 15476 66256 15724 66296
rect 15764 66256 15773 66296
rect 17923 66256 17932 66296
rect 17972 66256 18028 66296
rect 18068 66256 18077 66296
rect 3523 66172 3532 66212
rect 3572 66172 3820 66212
rect 3860 66172 3869 66212
rect 4291 66172 4300 66212
rect 4340 66172 6892 66212
rect 6932 66172 6941 66212
rect 7267 66172 7276 66212
rect 7316 66172 7325 66212
rect 10627 66172 10636 66212
rect 10676 66172 12172 66212
rect 12212 66172 12221 66212
rect 15619 66172 15628 66212
rect 15668 66172 15820 66212
rect 15860 66172 15869 66212
rect 3331 66088 3340 66128
rect 3380 66088 3628 66128
rect 3668 66088 3677 66128
rect 5827 66088 5836 66128
rect 5876 66088 6988 66128
rect 7028 66088 7037 66128
rect 19171 66088 19180 66128
rect 19220 66088 19756 66128
rect 19796 66088 19805 66128
rect 6604 65960 6644 66088
rect 2765 65920 2860 65960
rect 2900 65920 2909 65960
rect 6595 65920 6604 65960
rect 6644 65920 6653 65960
rect 14563 65920 14572 65960
rect 14612 65920 14764 65960
rect 14804 65920 14813 65960
rect 3043 65836 3052 65876
rect 3092 65836 6124 65876
rect 6164 65836 6173 65876
rect 2563 65752 2572 65792
rect 2612 65752 2764 65792
rect 2804 65752 2813 65792
rect 3679 65752 3688 65792
rect 3728 65752 3770 65792
rect 3810 65752 3852 65792
rect 3892 65752 3934 65792
rect 3974 65752 4016 65792
rect 4056 65752 4065 65792
rect 16397 65752 16492 65792
rect 16532 65752 16541 65792
rect 18799 65752 18808 65792
rect 18848 65752 18890 65792
rect 18930 65752 18972 65792
rect 19012 65752 19054 65792
rect 19094 65752 19136 65792
rect 19176 65752 19185 65792
rect 4195 65584 4204 65624
rect 4244 65584 9292 65624
rect 9332 65584 9341 65624
rect 2083 65500 2092 65540
rect 2132 65500 10252 65540
rect 10292 65500 10301 65540
rect 2851 65416 2860 65456
rect 2900 65416 3148 65456
rect 3188 65416 3197 65456
rect 2947 65332 2956 65372
rect 2996 65332 4012 65372
rect 4052 65332 4061 65372
rect 5155 65332 5164 65372
rect 5204 65332 6316 65372
rect 6356 65332 6365 65372
rect 12739 65332 12748 65372
rect 12788 65332 14668 65372
rect 14708 65332 14717 65372
rect 2563 65248 2572 65288
rect 2612 65248 9676 65288
rect 9716 65248 9725 65288
rect 15341 65248 15436 65288
rect 15476 65248 15485 65288
rect 3331 65164 3340 65204
rect 3380 65164 3628 65204
rect 3668 65164 8812 65204
rect 8852 65164 8861 65204
rect 11203 65164 11212 65204
rect 11252 65164 11308 65204
rect 11348 65164 11357 65204
rect 3235 65080 3244 65120
rect 3284 65080 8564 65120
rect 4919 64996 4928 65036
rect 4968 64996 5010 65036
rect 5050 64996 5092 65036
rect 5132 64996 5174 65036
rect 5214 64996 5256 65036
rect 5296 64996 5305 65036
rect 3811 64912 3820 64952
rect 3860 64912 4492 64952
rect 4532 64912 4541 64952
rect 8524 64868 8564 65080
rect 10060 65080 13132 65120
rect 13172 65080 16396 65120
rect 16436 65080 16445 65120
rect 17251 65080 17260 65120
rect 17300 65080 17644 65120
rect 17684 65080 17693 65120
rect 10060 65036 10100 65080
rect 8611 64996 8620 65036
rect 8660 64996 10100 65036
rect 12931 64996 12940 65036
rect 12980 64996 13132 65036
rect 13172 64996 13228 65036
rect 13268 64996 13277 65036
rect 17347 64996 17356 65036
rect 17396 64996 17740 65036
rect 17780 64996 19084 65036
rect 19124 64996 19133 65036
rect 20039 64996 20048 65036
rect 20088 64996 20130 65036
rect 20170 64996 20212 65036
rect 20252 64996 20294 65036
rect 20334 64996 20376 65036
rect 20416 64996 20425 65036
rect 9187 64912 9196 64952
rect 9236 64912 9292 64952
rect 9332 64912 9341 64952
rect 5068 64828 6260 64868
rect 8524 64828 10100 64868
rect 13507 64828 13516 64868
rect 13556 64828 13612 64868
rect 13652 64828 13661 64868
rect 16771 64828 16780 64868
rect 16820 64828 17012 64868
rect 5068 64784 5108 64828
rect 6220 64784 6260 64828
rect 10060 64784 10100 64828
rect 2851 64744 2860 64784
rect 2900 64744 3340 64784
rect 3380 64744 5108 64784
rect 5539 64744 5548 64784
rect 5588 64744 6124 64784
rect 6164 64744 6173 64784
rect 6220 64744 6412 64784
rect 6452 64744 8852 64784
rect 10060 64744 10156 64784
rect 10196 64744 10205 64784
rect 8812 64700 8852 64744
rect 3043 64660 3052 64700
rect 3092 64660 3532 64700
rect 3572 64660 6316 64700
rect 6356 64660 6365 64700
rect 8803 64660 8812 64700
rect 8852 64660 8908 64700
rect 8948 64660 8957 64700
rect 13795 64660 13804 64700
rect 13844 64660 14860 64700
rect 14900 64660 15724 64700
rect 15764 64660 15773 64700
rect 2851 64576 2860 64616
rect 2900 64576 2956 64616
rect 2996 64576 3005 64616
rect 3427 64576 3436 64616
rect 3476 64576 4300 64616
rect 4340 64576 5836 64616
rect 5876 64576 5885 64616
rect 16972 64532 17012 64828
rect 17059 64576 17068 64616
rect 17108 64576 20140 64616
rect 20180 64576 20189 64616
rect 4867 64492 4876 64532
rect 4916 64492 6124 64532
rect 6164 64492 6173 64532
rect 16963 64492 16972 64532
rect 17012 64492 17021 64532
rect 1613 64408 1708 64448
rect 1748 64408 1757 64448
rect 10627 64324 10636 64364
rect 10676 64324 11500 64364
rect 11540 64324 11549 64364
rect 14755 64324 14764 64364
rect 14804 64324 15244 64364
rect 15284 64324 15293 64364
rect 3679 64240 3688 64280
rect 3728 64240 3770 64280
rect 3810 64240 3852 64280
rect 3892 64240 3934 64280
rect 3974 64240 4016 64280
rect 4056 64240 4065 64280
rect 18799 64240 18808 64280
rect 18848 64240 18890 64280
rect 18930 64240 18972 64280
rect 19012 64240 19054 64280
rect 19094 64240 19136 64280
rect 19176 64240 19185 64280
rect 2179 64156 2188 64196
rect 2228 64156 2476 64196
rect 2516 64156 2525 64196
rect 3436 64156 12556 64196
rect 12596 64156 12605 64196
rect 18211 64156 18220 64196
rect 18260 64156 20044 64196
rect 20084 64156 20093 64196
rect 2083 64072 2092 64112
rect 2132 64072 2284 64112
rect 2324 64072 2333 64112
rect 2179 63988 2188 64028
rect 2228 63988 2380 64028
rect 2420 63988 2429 64028
rect 2659 63904 2668 63944
rect 2708 63904 2956 63944
rect 2996 63904 3005 63944
rect 3436 63860 3476 64156
rect 4685 64072 4780 64112
rect 4820 64072 4829 64112
rect 7075 64072 7084 64112
rect 7124 64072 9196 64112
rect 9236 64072 9245 64112
rect 12547 64072 12556 64112
rect 12596 64072 18508 64112
rect 18548 64072 18557 64112
rect 4003 63988 4012 64028
rect 4052 63988 8756 64028
rect 8813 63988 8908 64028
rect 8948 63988 8957 64028
rect 18125 63988 18220 64028
rect 18260 63988 18269 64028
rect 8716 63944 8756 63988
rect 4109 63904 4204 63944
rect 4244 63904 4253 63944
rect 4771 63904 4780 63944
rect 4820 63904 5740 63944
rect 5780 63904 5789 63944
rect 8035 63904 8044 63944
rect 8084 63904 8428 63944
rect 8468 63904 8477 63944
rect 8716 63904 9964 63944
rect 10004 63904 10013 63944
rect 10060 63904 14092 63944
rect 14132 63904 14141 63944
rect 1987 63820 1996 63860
rect 2036 63820 3476 63860
rect 10060 63776 10100 63904
rect 16483 63820 16492 63860
rect 16532 63820 18988 63860
rect 19028 63820 19037 63860
rect 2851 63736 2860 63776
rect 2900 63736 2909 63776
rect 3235 63736 3244 63776
rect 3284 63736 10100 63776
rect 13891 63736 13900 63776
rect 13940 63736 14420 63776
rect 2860 63692 2900 63736
rect 2563 63652 2572 63692
rect 2612 63652 4780 63692
rect 4820 63652 4829 63692
rect 5635 63652 5644 63692
rect 5684 63652 5779 63692
rect 6211 63652 6220 63692
rect 6260 63652 6796 63692
rect 6836 63652 6845 63692
rect 7747 63652 7756 63692
rect 7796 63652 10348 63692
rect 10388 63652 10397 63692
rect 11491 63652 11500 63692
rect 11540 63652 12076 63692
rect 12116 63652 12125 63692
rect 13987 63652 13996 63692
rect 14036 63652 14284 63692
rect 14324 63652 14333 63692
rect 14380 63608 14420 63736
rect 14467 63652 14476 63692
rect 14516 63652 15244 63692
rect 15284 63652 15293 63692
rect 18307 63652 18316 63692
rect 18356 63652 18412 63692
rect 18452 63652 18461 63692
rect 4205 63568 4300 63608
rect 4340 63568 4349 63608
rect 11779 63568 11788 63608
rect 11828 63568 12748 63608
rect 12788 63568 12797 63608
rect 14284 63568 14420 63608
rect 15235 63568 15244 63608
rect 15284 63568 16012 63608
rect 16052 63568 16061 63608
rect 14284 63524 14324 63568
rect 1804 63484 1900 63524
rect 1940 63484 1949 63524
rect 3053 63484 3148 63524
rect 3188 63484 3197 63524
rect 3427 63484 3436 63524
rect 3476 63484 4684 63524
rect 4724 63484 4733 63524
rect 4919 63484 4928 63524
rect 4968 63484 5010 63524
rect 5050 63484 5092 63524
rect 5132 63484 5174 63524
rect 5214 63484 5256 63524
rect 5296 63484 5305 63524
rect 6691 63484 6700 63524
rect 6740 63484 6932 63524
rect 8899 63484 8908 63524
rect 8948 63484 8957 63524
rect 13411 63484 13420 63524
rect 13460 63484 13469 63524
rect 14275 63484 14284 63524
rect 14324 63484 14333 63524
rect 19747 63484 19756 63524
rect 19796 63484 19805 63524
rect 20039 63484 20048 63524
rect 20088 63484 20130 63524
rect 20170 63484 20212 63524
rect 20252 63484 20294 63524
rect 20334 63484 20376 63524
rect 20416 63484 20425 63524
rect 1804 63380 1844 63484
rect 2371 63400 2380 63440
rect 2420 63400 2429 63440
rect 3427 63400 3436 63440
rect 3476 63400 3485 63440
rect 1804 63356 1940 63380
rect 1421 63316 1516 63356
rect 1556 63316 1565 63356
rect 1699 63316 1708 63356
rect 1748 63316 1940 63356
rect 2380 63272 2420 63400
rect 3436 63356 3476 63400
rect 2659 63316 2668 63356
rect 2708 63316 2860 63356
rect 2900 63316 2909 63356
rect 3139 63316 3148 63356
rect 3188 63316 3476 63356
rect 5251 63316 5260 63356
rect 5300 63316 5644 63356
rect 5684 63316 5693 63356
rect 6115 63316 6124 63356
rect 6164 63316 6700 63356
rect 6740 63316 6749 63356
rect 1411 63232 1420 63272
rect 1460 63232 2420 63272
rect 2957 63232 3052 63272
rect 3092 63232 3101 63272
rect 3427 63232 3436 63272
rect 3476 63232 3532 63272
rect 3572 63232 3581 63272
rect 4675 63148 4684 63188
rect 4724 63148 5452 63188
rect 5492 63148 5501 63188
rect 6892 63104 6932 63484
rect 7939 63400 7948 63440
rect 7988 63400 8140 63440
rect 8180 63400 8189 63440
rect 8908 63380 8948 63484
rect 13420 63440 13460 63484
rect 12451 63400 12460 63440
rect 12500 63400 12652 63440
rect 12692 63400 12701 63440
rect 13420 63400 14092 63440
rect 14132 63400 14141 63440
rect 18115 63400 18124 63440
rect 18164 63400 18173 63440
rect 19363 63400 19372 63440
rect 19412 63400 19421 63440
rect 8899 63340 8908 63380
rect 8948 63340 8957 63380
rect 18124 63356 18164 63400
rect 13228 63316 13612 63356
rect 13652 63316 13661 63356
rect 14371 63316 14380 63356
rect 14420 63316 15052 63356
rect 15092 63316 15101 63356
rect 18124 63316 18316 63356
rect 18356 63316 18365 63356
rect 8323 63232 8332 63272
rect 8372 63232 8620 63272
rect 8660 63232 8669 63272
rect 13228 63188 13268 63316
rect 13315 63232 13324 63272
rect 13364 63232 13373 63272
rect 13507 63232 13516 63272
rect 13556 63232 13708 63272
rect 13748 63232 13757 63272
rect 18115 63232 18124 63272
rect 18164 63232 18220 63272
rect 18260 63232 18269 63272
rect 13324 63188 13364 63232
rect 8227 63148 8236 63188
rect 8276 63148 9676 63188
rect 9716 63148 9725 63188
rect 13219 63148 13228 63188
rect 13268 63148 13277 63188
rect 13324 63148 13900 63188
rect 13940 63148 13949 63188
rect 14371 63148 14380 63188
rect 14420 63148 15532 63188
rect 15572 63148 15581 63188
rect 4387 63064 4396 63104
rect 4436 63064 4780 63104
rect 4820 63064 4829 63104
rect 6892 63064 6988 63104
rect 7028 63064 7037 63104
rect 7939 63064 7948 63104
rect 7988 63064 8620 63104
rect 8660 63064 8669 63104
rect 13229 63064 13324 63104
rect 13364 63064 13373 63104
rect 17923 63064 17932 63104
rect 17972 63064 18220 63104
rect 18260 63064 18269 63104
rect 2947 62980 2956 63020
rect 2996 62980 12172 63020
rect 12212 62980 12221 63020
rect 17059 62980 17068 63020
rect 17108 62980 18988 63020
rect 19028 62980 19037 63020
rect 1411 62896 1420 62936
rect 1460 62896 4780 62936
rect 4820 62896 4829 62936
rect 13987 62896 13996 62936
rect 14036 62896 14092 62936
rect 14132 62896 14141 62936
rect 19372 62852 19412 63400
rect 2851 62812 2860 62852
rect 2900 62812 4972 62852
rect 5012 62812 5021 62852
rect 6989 62812 7084 62852
rect 7124 62812 7133 62852
rect 11875 62812 11884 62852
rect 11924 62812 12268 62852
rect 12308 62812 12317 62852
rect 15043 62812 15052 62852
rect 15092 62812 15244 62852
rect 15284 62812 15293 62852
rect 17923 62812 17932 62852
rect 17972 62812 18316 62852
rect 18356 62812 18365 62852
rect 19267 62812 19276 62852
rect 19316 62812 19412 62852
rect 3679 62728 3688 62768
rect 3728 62728 3770 62768
rect 3810 62728 3852 62768
rect 3892 62728 3934 62768
rect 3974 62728 4016 62768
rect 4056 62728 4065 62768
rect 4195 62728 4204 62768
rect 4244 62728 9964 62768
rect 10004 62728 10013 62768
rect 18799 62728 18808 62768
rect 18848 62728 18890 62768
rect 18930 62728 18972 62768
rect 19012 62728 19054 62768
rect 19094 62728 19136 62768
rect 19176 62728 19185 62768
rect 15235 62644 15244 62684
rect 15284 62644 15436 62684
rect 15476 62644 15485 62684
rect 19756 62600 19796 63484
rect 19843 63400 19852 63440
rect 19892 63400 20620 63440
rect 20660 63400 20669 63440
rect 20803 63064 20812 63104
rect 20852 63064 21100 63104
rect 21140 63064 21149 63104
rect 19171 62560 19180 62600
rect 19220 62560 19796 62600
rect 7171 62476 7180 62516
rect 7220 62476 7372 62516
rect 7412 62476 7421 62516
rect 12835 62476 12844 62516
rect 12884 62476 13132 62516
rect 13172 62476 13181 62516
rect 13996 62476 16436 62516
rect 17165 62476 17260 62516
rect 17300 62476 17309 62516
rect 20611 62476 20620 62516
rect 20660 62476 21196 62516
rect 21236 62476 21245 62516
rect 13996 62432 14036 62476
rect 16396 62432 16436 62476
rect 8515 62392 8524 62432
rect 8564 62392 9196 62432
rect 9236 62392 9964 62432
rect 10004 62392 10013 62432
rect 13987 62392 13996 62432
rect 14036 62392 14045 62432
rect 15149 62392 15244 62432
rect 15284 62392 15532 62432
rect 15572 62392 15581 62432
rect 15907 62392 15916 62432
rect 15956 62392 16012 62432
rect 16052 62392 16061 62432
rect 16387 62392 16396 62432
rect 16436 62392 16684 62432
rect 16724 62392 16733 62432
rect 4003 62308 4012 62348
rect 4052 62308 4204 62348
rect 4244 62308 4253 62348
rect 6307 62308 6316 62348
rect 6356 62308 17932 62348
rect 17972 62308 17981 62348
rect 20611 62308 20620 62348
rect 20660 62308 20908 62348
rect 20948 62308 20957 62348
rect 13507 62224 13516 62264
rect 13556 62224 20044 62264
rect 20084 62224 20093 62264
rect 2947 62140 2956 62180
rect 2996 62140 3148 62180
rect 3188 62140 3197 62180
rect 4771 62140 4780 62180
rect 4820 62140 4876 62180
rect 4916 62140 4925 62180
rect 20140 62140 20236 62180
rect 20276 62140 20285 62180
rect 20140 62096 20180 62140
rect 8995 62056 9004 62096
rect 9044 62056 11116 62096
rect 11156 62056 11165 62096
rect 16867 62056 16876 62096
rect 16916 62056 17260 62096
rect 17300 62056 17309 62096
rect 19660 62056 20180 62096
rect 4919 61972 4928 62012
rect 4968 61972 5010 62012
rect 5050 61972 5092 62012
rect 5132 61972 5174 62012
rect 5214 61972 5256 62012
rect 5296 61972 5305 62012
rect 9187 61972 9196 62012
rect 9236 61972 10156 62012
rect 10196 61972 10205 62012
rect 19660 61928 19700 62056
rect 20039 61972 20048 62012
rect 20088 61972 20130 62012
rect 20170 61972 20212 62012
rect 20252 61972 20294 62012
rect 20334 61972 20376 62012
rect 20416 61972 20425 62012
rect 19651 61888 19660 61928
rect 19700 61888 19709 61928
rect 2659 61804 2668 61844
rect 2708 61804 5740 61844
rect 5780 61804 6700 61844
rect 6740 61804 6749 61844
rect 11021 61804 11116 61844
rect 11156 61804 11165 61844
rect 15715 61804 15724 61844
rect 15764 61804 17068 61844
rect 17108 61804 17117 61844
rect 14371 61720 14380 61760
rect 14420 61720 20428 61760
rect 20468 61720 20477 61760
rect 3437 61636 3532 61676
rect 3572 61636 3581 61676
rect 7075 61636 7084 61676
rect 7124 61636 7372 61676
rect 7412 61636 7421 61676
rect 15917 61636 16012 61676
rect 16052 61636 16061 61676
rect 4003 61552 4012 61592
rect 4052 61552 4300 61592
rect 4340 61552 4349 61592
rect 4579 61552 4588 61592
rect 4628 61552 4637 61592
rect 17059 61552 17068 61592
rect 17108 61552 18220 61592
rect 18260 61552 18988 61592
rect 19028 61552 19037 61592
rect 2179 61468 2188 61508
rect 2228 61468 2572 61508
rect 2612 61468 2621 61508
rect 4300 61424 4340 61552
rect 4588 61508 4628 61552
rect 4588 61468 5452 61508
rect 5492 61468 5501 61508
rect 6019 61468 6028 61508
rect 6068 61468 6700 61508
rect 6740 61468 6749 61508
rect 6989 61468 7084 61508
rect 7124 61468 7133 61508
rect 15043 61468 15052 61508
rect 15092 61468 15628 61508
rect 15668 61468 15677 61508
rect 17347 61468 17356 61508
rect 17396 61468 17452 61508
rect 17492 61468 17836 61508
rect 17876 61468 17885 61508
rect 19171 61468 19180 61508
rect 19220 61468 19468 61508
rect 19508 61468 19517 61508
rect 3619 61384 3628 61424
rect 3668 61384 3677 61424
rect 4300 61384 4588 61424
rect 4628 61384 4637 61424
rect 21187 61384 21196 61424
rect 21236 61384 21428 61424
rect 3628 61340 3668 61384
rect 3532 61300 3668 61340
rect 3532 61172 3572 61300
rect 21388 61256 21428 61384
rect 3679 61216 3688 61256
rect 3728 61216 3770 61256
rect 3810 61216 3852 61256
rect 3892 61216 3934 61256
rect 3974 61216 4016 61256
rect 4056 61216 4065 61256
rect 18799 61216 18808 61256
rect 18848 61216 18890 61256
rect 18930 61216 18972 61256
rect 19012 61216 19054 61256
rect 19094 61216 19136 61256
rect 19176 61216 19185 61256
rect 20995 61216 21004 61256
rect 21044 61216 21053 61256
rect 21379 61216 21388 61256
rect 21428 61216 21437 61256
rect 21004 61172 21044 61216
rect 3532 61132 3860 61172
rect 9571 61132 9580 61172
rect 9620 61132 9868 61172
rect 9908 61132 9917 61172
rect 12259 61132 12268 61172
rect 12308 61132 12556 61172
rect 12596 61132 12605 61172
rect 21004 61132 21196 61172
rect 21236 61132 21245 61172
rect 3820 61088 3860 61132
rect 3523 61048 3532 61088
rect 3572 61048 3628 61088
rect 3668 61048 3677 61088
rect 3811 61048 3820 61088
rect 3860 61048 3869 61088
rect 20419 61048 20428 61088
rect 20468 61048 21004 61088
rect 21044 61048 21053 61088
rect 2659 60964 2668 61004
rect 2708 60964 3436 61004
rect 3476 60964 3724 61004
rect 3764 60964 3773 61004
rect 4003 60880 4012 60920
rect 4052 60880 4204 60920
rect 4244 60880 7372 60920
rect 7412 60880 7421 60920
rect 3907 60712 3916 60752
rect 3956 60712 4204 60752
rect 4244 60712 6124 60752
rect 6164 60712 6173 60752
rect 7363 60712 7372 60752
rect 7412 60712 8332 60752
rect 8372 60712 8381 60752
rect 8035 60544 8044 60584
rect 8084 60544 12172 60584
rect 12212 60544 12221 60584
rect 17165 60544 17260 60584
rect 17300 60544 17309 60584
rect 4919 60460 4928 60500
rect 4968 60460 5010 60500
rect 5050 60460 5092 60500
rect 5132 60460 5174 60500
rect 5214 60460 5256 60500
rect 5296 60460 5305 60500
rect 7459 60460 7468 60500
rect 7508 60460 11596 60500
rect 11636 60460 11645 60500
rect 12451 60460 12460 60500
rect 12500 60460 15532 60500
rect 15572 60460 15581 60500
rect 16387 60460 16396 60500
rect 16436 60460 17932 60500
rect 17972 60460 17981 60500
rect 20039 60460 20048 60500
rect 20088 60460 20130 60500
rect 20170 60460 20212 60500
rect 20252 60460 20294 60500
rect 20334 60460 20376 60500
rect 20416 60460 20425 60500
rect 2467 60376 2476 60416
rect 2516 60376 4916 60416
rect 4876 60332 4916 60376
rect 2467 60292 2476 60332
rect 2516 60292 3916 60332
rect 3956 60292 3965 60332
rect 4867 60292 4876 60332
rect 4916 60292 4925 60332
rect 12557 60292 12652 60332
rect 12692 60292 12701 60332
rect 1891 60208 1900 60248
rect 1940 60208 5356 60248
rect 5396 60208 5405 60248
rect 5452 60208 11884 60248
rect 11924 60208 11933 60248
rect 12259 60208 12268 60248
rect 12308 60208 14380 60248
rect 14420 60208 14429 60248
rect 15907 60208 15916 60248
rect 15956 60208 16204 60248
rect 16244 60208 16253 60248
rect 5452 60164 5492 60208
rect 3427 60124 3436 60164
rect 3476 60124 5492 60164
rect 5923 60124 5932 60164
rect 5972 60124 7948 60164
rect 7988 60124 7997 60164
rect 8707 60124 8716 60164
rect 8756 60124 14668 60164
rect 14708 60124 14717 60164
rect 17539 60124 17548 60164
rect 17588 60124 18124 60164
rect 18164 60124 18173 60164
rect 5932 60080 5972 60124
rect 2275 60040 2284 60080
rect 2324 60040 5972 60080
rect 12163 60040 12172 60080
rect 12212 60040 12652 60080
rect 12692 60040 12701 60080
rect 14371 60040 14380 60080
rect 14420 60040 14476 60080
rect 14516 60040 14525 60080
rect 15907 60040 15916 60080
rect 15956 60040 16972 60080
rect 17012 60040 17021 60080
rect 17443 60040 17452 60080
rect 17492 60040 17740 60080
rect 17780 60040 17789 60080
rect 18403 60040 18412 60080
rect 18452 60040 18461 60080
rect 3907 59956 3916 59996
rect 3956 59956 11884 59996
rect 11924 59956 11933 59996
rect 12835 59872 12844 59912
rect 12884 59872 18316 59912
rect 18356 59872 18365 59912
rect 14659 59788 14668 59828
rect 14708 59788 15916 59828
rect 15956 59788 15965 59828
rect 18412 59744 18452 60040
rect 3679 59704 3688 59744
rect 3728 59704 3770 59744
rect 3810 59704 3852 59744
rect 3892 59704 3934 59744
rect 3974 59704 4016 59744
rect 4056 59704 4065 59744
rect 6979 59704 6988 59744
rect 7028 59704 17836 59744
rect 17876 59704 17885 59744
rect 18307 59704 18316 59744
rect 18356 59704 18452 59744
rect 18799 59704 18808 59744
rect 18848 59704 18890 59744
rect 18930 59704 18972 59744
rect 19012 59704 19054 59744
rect 19094 59704 19136 59744
rect 19176 59704 19185 59744
rect 11779 59620 11788 59660
rect 11828 59620 12172 59660
rect 12212 59620 12221 59660
rect 3427 59536 3436 59576
rect 3476 59536 3628 59576
rect 3668 59536 3677 59576
rect 1411 59368 1420 59408
rect 1460 59368 2092 59408
rect 2132 59368 2141 59408
rect 10339 59368 10348 59408
rect 10388 59368 14668 59408
rect 14708 59368 14717 59408
rect 1507 59284 1516 59324
rect 1556 59284 1900 59324
rect 1940 59284 1949 59324
rect 11107 59284 11116 59324
rect 11156 59284 14956 59324
rect 14996 59284 15005 59324
rect 16003 59284 16012 59324
rect 16052 59284 18316 59324
rect 18356 59284 19468 59324
rect 19508 59284 19517 59324
rect 11875 59200 11884 59240
rect 11924 59200 12268 59240
rect 12308 59200 12317 59240
rect 4387 59116 4396 59156
rect 4436 59116 4876 59156
rect 4916 59116 4925 59156
rect 15341 59116 15436 59156
rect 15476 59116 15485 59156
rect 4919 58948 4928 58988
rect 4968 58948 5010 58988
rect 5050 58948 5092 58988
rect 5132 58948 5174 58988
rect 5214 58948 5256 58988
rect 5296 58948 5305 58988
rect 11203 58948 11212 58988
rect 11252 58948 12940 58988
rect 12980 58948 12989 58988
rect 20039 58948 20048 58988
rect 20088 58948 20130 58988
rect 20170 58948 20212 58988
rect 20252 58948 20294 58988
rect 20334 58948 20376 58988
rect 20416 58948 20425 58988
rect 5549 58780 5644 58820
rect 5684 58780 5693 58820
rect 20035 58780 20044 58820
rect 20084 58780 20524 58820
rect 20564 58780 20573 58820
rect 9955 58696 9964 58736
rect 10004 58696 12172 58736
rect 12212 58696 12221 58736
rect 13036 58696 13132 58736
rect 13172 58696 13181 58736
rect 13036 58652 13076 58696
rect 13027 58612 13036 58652
rect 13076 58612 13085 58652
rect 11203 58528 11212 58568
rect 11252 58528 11596 58568
rect 11636 58528 11645 58568
rect 13037 58528 13132 58568
rect 13172 58528 13181 58568
rect 17165 58528 17260 58568
rect 17300 58528 17309 58568
rect 2851 58444 2860 58484
rect 2900 58444 3532 58484
rect 3572 58444 3581 58484
rect 10435 58444 10444 58484
rect 10484 58444 12172 58484
rect 12212 58444 12221 58484
rect 13507 58444 13516 58484
rect 13556 58444 13565 58484
rect 18019 58444 18028 58484
rect 18068 58444 18796 58484
rect 18836 58444 18845 58484
rect 19363 58444 19372 58484
rect 19412 58444 19564 58484
rect 19604 58444 19613 58484
rect 3139 58360 3148 58400
rect 3188 58360 3340 58400
rect 3380 58360 3389 58400
rect 11011 58360 11020 58400
rect 11060 58360 11500 58400
rect 11540 58360 11549 58400
rect 13516 58316 13556 58444
rect 15907 58360 15916 58400
rect 15956 58360 16108 58400
rect 16148 58360 16157 58400
rect 18125 58360 18220 58400
rect 18260 58360 18269 58400
rect 3523 58276 3532 58316
rect 3572 58276 6412 58316
rect 6452 58276 6461 58316
rect 13123 58276 13132 58316
rect 13172 58276 13556 58316
rect 3043 58192 3052 58232
rect 3092 58192 3148 58232
rect 3188 58192 3197 58232
rect 3679 58192 3688 58232
rect 3728 58192 3770 58232
rect 3810 58192 3852 58232
rect 3892 58192 3934 58232
rect 3974 58192 4016 58232
rect 4056 58192 4065 58232
rect 12077 58192 12172 58232
rect 12212 58192 12221 58232
rect 16099 58192 16108 58232
rect 16148 58192 16684 58232
rect 16724 58192 16733 58232
rect 18799 58192 18808 58232
rect 18848 58192 18890 58232
rect 18930 58192 18972 58232
rect 19012 58192 19054 58232
rect 19094 58192 19136 58232
rect 19176 58192 19185 58232
rect 10915 58108 10924 58148
rect 10964 58108 14764 58148
rect 14804 58108 14813 58148
rect 10915 57940 10924 57980
rect 10964 57940 12076 57980
rect 12116 57940 12268 57980
rect 12308 57940 12317 57980
rect 2659 57856 2668 57896
rect 2708 57856 4916 57896
rect 12931 57856 12940 57896
rect 12980 57856 17452 57896
rect 17492 57856 18220 57896
rect 18260 57856 18412 57896
rect 18452 57856 18461 57896
rect 4876 57812 4916 57856
rect 4003 57772 4012 57812
rect 4052 57772 4204 57812
rect 4244 57772 4253 57812
rect 4867 57772 4876 57812
rect 4916 57772 6412 57812
rect 6452 57772 6461 57812
rect 10531 57772 10540 57812
rect 10580 57772 11788 57812
rect 11828 57772 11837 57812
rect 14275 57772 14284 57812
rect 14324 57772 16684 57812
rect 16724 57772 18892 57812
rect 18932 57772 20044 57812
rect 20084 57772 20093 57812
rect 10915 57688 10924 57728
rect 10964 57688 11884 57728
rect 11924 57688 11933 57728
rect 19459 57688 19468 57728
rect 19508 57688 19852 57728
rect 19892 57688 19901 57728
rect 3619 57604 3628 57644
rect 3668 57604 11404 57644
rect 11444 57604 11453 57644
rect 16963 57604 16972 57644
rect 17012 57604 17068 57644
rect 17108 57604 17117 57644
rect 11587 57520 11596 57560
rect 11636 57520 12076 57560
rect 12116 57520 12125 57560
rect 4919 57436 4928 57476
rect 4968 57436 5010 57476
rect 5050 57436 5092 57476
rect 5132 57436 5174 57476
rect 5214 57436 5256 57476
rect 5296 57436 5305 57476
rect 20039 57436 20048 57476
rect 20088 57436 20130 57476
rect 20170 57436 20212 57476
rect 20252 57436 20294 57476
rect 20334 57436 20376 57476
rect 20416 57436 20425 57476
rect 1795 57352 1804 57392
rect 1844 57352 13228 57392
rect 13268 57352 13277 57392
rect 2659 57268 2668 57308
rect 2708 57268 8908 57308
rect 8948 57268 8957 57308
rect 5539 56932 5548 56972
rect 5588 56932 5644 56972
rect 5684 56932 5693 56972
rect 3427 56848 3436 56888
rect 3476 56848 3628 56888
rect 3668 56848 3677 56888
rect 3679 56680 3688 56720
rect 3728 56680 3770 56720
rect 3810 56680 3852 56720
rect 3892 56680 3934 56720
rect 3974 56680 4016 56720
rect 4056 56680 4065 56720
rect 18799 56680 18808 56720
rect 18848 56680 18890 56720
rect 18930 56680 18972 56720
rect 19012 56680 19054 56720
rect 19094 56680 19136 56720
rect 19176 56680 19185 56720
rect 9283 56512 9292 56552
rect 9332 56512 10060 56552
rect 10100 56512 10109 56552
rect 6317 56344 6412 56384
rect 6452 56344 6461 56384
rect 17635 56344 17644 56384
rect 17684 56344 17740 56384
rect 17780 56344 17789 56384
rect 18307 56344 18316 56384
rect 18356 56344 19180 56384
rect 19220 56344 19229 56384
rect 13795 56260 13804 56300
rect 13844 56260 15436 56300
rect 15476 56260 15485 56300
rect 16973 56176 17068 56216
rect 17108 56176 17117 56216
rect 17827 56176 17836 56216
rect 17876 56176 18220 56216
rect 18260 56176 18269 56216
rect 8131 56092 8140 56132
rect 8180 56092 8812 56132
rect 8852 56092 8861 56132
rect 16483 56092 16492 56132
rect 16532 56092 18316 56132
rect 18356 56092 18365 56132
rect 4919 55924 4928 55964
rect 4968 55924 5010 55964
rect 5050 55924 5092 55964
rect 5132 55924 5174 55964
rect 5214 55924 5256 55964
rect 5296 55924 5305 55964
rect 20039 55924 20048 55964
rect 20088 55924 20130 55964
rect 20170 55924 20212 55964
rect 20252 55924 20294 55964
rect 20334 55924 20376 55964
rect 20416 55924 20425 55964
rect 18403 55504 18412 55544
rect 18452 55504 19660 55544
rect 19700 55504 19709 55544
rect 6125 55336 6220 55376
rect 6260 55336 6269 55376
rect 18700 55336 18796 55376
rect 18836 55336 18845 55376
rect 19651 55336 19660 55376
rect 19700 55336 19948 55376
rect 19988 55336 19997 55376
rect 3679 55168 3688 55208
rect 3728 55168 3770 55208
rect 3810 55168 3852 55208
rect 3892 55168 3934 55208
rect 3974 55168 4016 55208
rect 4056 55168 4065 55208
rect 18700 55124 18740 55336
rect 18799 55168 18808 55208
rect 18848 55168 18890 55208
rect 18930 55168 18972 55208
rect 19012 55168 19054 55208
rect 19094 55168 19136 55208
rect 19176 55168 19185 55208
rect 18700 55084 18836 55124
rect 18796 55040 18836 55084
rect 18787 55000 18796 55040
rect 18836 55000 18845 55040
rect 1699 54916 1708 54956
rect 1748 54916 2668 54956
rect 2708 54916 2860 54956
rect 2900 54916 2909 54956
rect 2563 54832 2572 54872
rect 2612 54832 9004 54872
rect 9044 54832 9292 54872
rect 9332 54832 9341 54872
rect 1987 54748 1996 54788
rect 2036 54748 3244 54788
rect 3284 54748 3293 54788
rect 4483 54748 4492 54788
rect 4532 54748 4780 54788
rect 4820 54748 4829 54788
rect 3811 54664 3820 54704
rect 3860 54664 7180 54704
rect 7220 54664 7229 54704
rect 4919 54412 4928 54452
rect 4968 54412 5010 54452
rect 5050 54412 5092 54452
rect 5132 54412 5174 54452
rect 5214 54412 5256 54452
rect 5296 54412 5305 54452
rect 20039 54412 20048 54452
rect 20088 54412 20130 54452
rect 20170 54412 20212 54452
rect 20252 54412 20294 54452
rect 20334 54412 20376 54452
rect 20416 54412 20425 54452
rect 5923 54328 5932 54368
rect 5972 54328 12980 54368
rect 1603 54244 1612 54284
rect 1652 54244 6028 54284
rect 6068 54244 6220 54284
rect 6260 54244 6269 54284
rect 7853 54244 7948 54284
rect 7988 54244 7997 54284
rect 12940 54200 12980 54328
rect 19459 54244 19468 54284
rect 19508 54244 20044 54284
rect 20084 54244 20093 54284
rect 9571 54160 9580 54200
rect 9620 54160 9868 54200
rect 9908 54160 9917 54200
rect 12940 54160 14476 54200
rect 14516 54160 14525 54200
rect 1699 53992 1708 54032
rect 1748 53992 4492 54032
rect 4532 53992 4541 54032
rect 15811 53992 15820 54032
rect 15860 53992 16204 54032
rect 16244 53992 18316 54032
rect 18356 53992 18508 54032
rect 18548 53992 18892 54032
rect 18932 53992 18941 54032
rect 6115 53908 6124 53948
rect 6164 53908 6316 53948
rect 6356 53908 6365 53948
rect 7747 53908 7756 53948
rect 7796 53908 8236 53948
rect 8276 53908 8285 53948
rect 3235 53824 3244 53864
rect 3284 53824 3724 53864
rect 3764 53824 3773 53864
rect 10435 53824 10444 53864
rect 10484 53824 10636 53864
rect 10676 53824 10685 53864
rect 6115 53740 6124 53780
rect 6164 53740 6700 53780
rect 6740 53740 6749 53780
rect 3679 53656 3688 53696
rect 3728 53656 3770 53696
rect 3810 53656 3852 53696
rect 3892 53656 3934 53696
rect 3974 53656 4016 53696
rect 4056 53656 4065 53696
rect 18799 53656 18808 53696
rect 18848 53656 18890 53696
rect 18930 53656 18972 53696
rect 19012 53656 19054 53696
rect 19094 53656 19136 53696
rect 19176 53656 19185 53696
rect 18307 53572 18316 53612
rect 18356 53572 19372 53612
rect 19412 53572 19421 53612
rect 2093 53488 2188 53528
rect 2228 53488 2237 53528
rect 9955 53488 9964 53528
rect 10004 53488 14284 53528
rect 14324 53488 14333 53528
rect 3043 53404 3052 53444
rect 3092 53404 3436 53444
rect 3476 53404 3485 53444
rect 10541 53404 10636 53444
rect 10676 53404 10685 53444
rect 10915 53404 10924 53444
rect 10964 53404 10973 53444
rect 10924 53360 10964 53404
rect 2659 53320 2668 53360
rect 2708 53320 2860 53360
rect 2900 53320 2909 53360
rect 3148 53320 3532 53360
rect 3572 53320 3581 53360
rect 10147 53320 10156 53360
rect 10196 53320 10964 53360
rect 13229 53320 13324 53360
rect 13364 53320 13373 53360
rect 14083 53320 14092 53360
rect 14132 53320 14380 53360
rect 14420 53320 14429 53360
rect 15917 53320 16012 53360
rect 16052 53320 16061 53360
rect 17357 53320 17452 53360
rect 17492 53320 17501 53360
rect 3148 53276 3188 53320
rect 3043 53236 3052 53276
rect 3092 53236 3188 53276
rect 6979 53260 6988 53300
rect 7028 53260 7037 53300
rect 6988 53192 7028 53260
rect 15235 53236 15244 53276
rect 15284 53236 15628 53276
rect 15668 53236 15677 53276
rect 19459 53236 19468 53276
rect 19508 53236 19660 53276
rect 19700 53236 19709 53276
rect 2659 53152 2668 53192
rect 2708 53152 2860 53192
rect 2900 53152 2909 53192
rect 6988 53152 7180 53192
rect 7220 53152 7229 53192
rect 2659 53068 2668 53108
rect 2708 53068 2860 53108
rect 2900 53068 2909 53108
rect 9763 53068 9772 53108
rect 9812 53068 10540 53108
rect 10580 53068 10589 53108
rect 4919 52900 4928 52940
rect 4968 52900 5010 52940
rect 5050 52900 5092 52940
rect 5132 52900 5174 52940
rect 5214 52900 5256 52940
rect 5296 52900 5305 52940
rect 20039 52900 20048 52940
rect 20088 52900 20130 52940
rect 20170 52900 20212 52940
rect 20252 52900 20294 52940
rect 20334 52900 20376 52940
rect 20416 52900 20425 52940
rect 7075 52816 7084 52856
rect 7124 52816 8812 52856
rect 8852 52816 8861 52856
rect 10339 52732 10348 52772
rect 10388 52732 10732 52772
rect 10772 52732 10781 52772
rect 6499 52564 6508 52604
rect 6548 52564 6557 52604
rect 6508 52436 6548 52564
rect 10435 52480 10444 52520
rect 10484 52480 20140 52520
rect 20180 52480 20189 52520
rect 6508 52396 6892 52436
rect 6932 52396 6941 52436
rect 3679 52144 3688 52184
rect 3728 52144 3770 52184
rect 3810 52144 3852 52184
rect 3892 52144 3934 52184
rect 3974 52144 4016 52184
rect 4056 52144 4065 52184
rect 15235 52144 15244 52184
rect 15284 52144 15628 52184
rect 15668 52144 15677 52184
rect 18799 52144 18808 52184
rect 18848 52144 18890 52184
rect 18930 52144 18972 52184
rect 19012 52144 19054 52184
rect 19094 52144 19136 52184
rect 19176 52144 19185 52184
rect 3235 51892 3244 51932
rect 3284 51892 9772 51932
rect 9812 51892 9821 51932
rect 16387 51892 16396 51932
rect 16436 51892 18028 51932
rect 18068 51892 18077 51932
rect 18403 51892 18412 51932
rect 18452 51892 18604 51932
rect 18644 51892 18653 51932
rect 1709 51808 1804 51848
rect 1844 51808 1853 51848
rect 15331 51808 15340 51848
rect 15380 51808 20140 51848
rect 20180 51808 20189 51848
rect 6979 51640 6988 51680
rect 7028 51640 8428 51680
rect 8468 51640 8477 51680
rect 9091 51640 9100 51680
rect 9140 51640 9292 51680
rect 9332 51640 9341 51680
rect 4919 51388 4928 51428
rect 4968 51388 5010 51428
rect 5050 51388 5092 51428
rect 5132 51388 5174 51428
rect 5214 51388 5256 51428
rect 5296 51388 5305 51428
rect 20039 51388 20048 51428
rect 20088 51388 20130 51428
rect 20170 51388 20212 51428
rect 20252 51388 20294 51428
rect 20334 51388 20376 51428
rect 20416 51388 20425 51428
rect 11203 51052 11212 51092
rect 11252 51052 16780 51092
rect 16820 51052 16829 51092
rect 2477 50968 2572 51008
rect 2612 50968 2621 51008
rect 14563 50968 14572 51008
rect 14612 50968 19372 51008
rect 19412 50968 19421 51008
rect 2285 50800 2380 50840
rect 2420 50800 2429 50840
rect 3679 50632 3688 50672
rect 3728 50632 3770 50672
rect 3810 50632 3852 50672
rect 3892 50632 3934 50672
rect 3974 50632 4016 50672
rect 4056 50632 4065 50672
rect 18799 50632 18808 50672
rect 18848 50632 18890 50672
rect 18930 50632 18972 50672
rect 19012 50632 19054 50672
rect 19094 50632 19136 50672
rect 19176 50632 19185 50672
rect 11107 50464 11116 50504
rect 11156 50464 11692 50504
rect 11732 50464 11741 50504
rect 6787 50380 6796 50420
rect 6836 50380 11596 50420
rect 11636 50380 11645 50420
rect 10051 50296 10060 50336
rect 10100 50296 10828 50336
rect 10868 50296 10877 50336
rect 11309 50296 11404 50336
rect 11444 50296 11453 50336
rect 12173 50296 12268 50336
rect 12308 50296 12317 50336
rect 12643 50296 12652 50336
rect 12692 50296 16396 50336
rect 16436 50296 16445 50336
rect 10147 50212 10156 50252
rect 10196 50212 10348 50252
rect 10388 50212 10397 50252
rect 12355 50212 12364 50252
rect 12404 50212 19180 50252
rect 19220 50212 19229 50252
rect 11011 50128 11020 50168
rect 11060 50128 19756 50168
rect 19796 50128 19805 50168
rect 11203 50044 11212 50084
rect 11252 50044 11308 50084
rect 11348 50044 11357 50084
rect 4919 49876 4928 49916
rect 4968 49876 5010 49916
rect 5050 49876 5092 49916
rect 5132 49876 5174 49916
rect 5214 49876 5256 49916
rect 5296 49876 5305 49916
rect 20039 49876 20048 49916
rect 20088 49876 20130 49916
rect 20170 49876 20212 49916
rect 20252 49876 20294 49916
rect 20334 49876 20376 49916
rect 20416 49876 20425 49916
rect 16099 49624 16108 49664
rect 16148 49624 16204 49664
rect 16244 49624 16253 49664
rect 19363 49624 19372 49664
rect 19412 49624 19660 49664
rect 19700 49624 19709 49664
rect 9571 49540 9580 49580
rect 9620 49540 9772 49580
rect 9812 49540 9821 49580
rect 10061 49540 10156 49580
rect 10196 49540 10205 49580
rect 10723 49540 10732 49580
rect 10772 49540 10828 49580
rect 10868 49540 10877 49580
rect 19363 49456 19372 49496
rect 19412 49456 20620 49496
rect 20660 49456 20669 49496
rect 17549 49288 17644 49328
rect 17684 49288 17693 49328
rect 3679 49120 3688 49160
rect 3728 49120 3770 49160
rect 3810 49120 3852 49160
rect 3892 49120 3934 49160
rect 3974 49120 4016 49160
rect 4056 49120 4065 49160
rect 18799 49120 18808 49160
rect 18848 49120 18890 49160
rect 18930 49120 18972 49160
rect 19012 49120 19054 49160
rect 19094 49120 19136 49160
rect 19176 49120 19185 49160
rect 15907 48952 15916 48992
rect 15956 48952 16300 48992
rect 16340 48952 16349 48992
rect 6115 48868 6124 48908
rect 6164 48868 10540 48908
rect 10580 48868 10589 48908
rect 10723 48868 10732 48908
rect 10772 48868 16396 48908
rect 16436 48868 16445 48908
rect 9581 48784 9676 48824
rect 9716 48784 9725 48824
rect 10051 48784 10060 48824
rect 10100 48784 19372 48824
rect 19412 48784 19421 48824
rect 5635 48700 5644 48740
rect 5684 48700 6124 48740
rect 6164 48700 6173 48740
rect 9187 48700 9196 48740
rect 9236 48700 9772 48740
rect 9812 48700 9821 48740
rect 12653 48700 12748 48740
rect 12788 48700 12797 48740
rect 13411 48700 13420 48740
rect 13460 48700 15820 48740
rect 15860 48700 15869 48740
rect 7555 48616 7564 48656
rect 7604 48616 9388 48656
rect 9428 48616 12268 48656
rect 12308 48616 12460 48656
rect 12500 48616 12509 48656
rect 4109 48532 4204 48572
rect 4244 48532 4253 48572
rect 7363 48448 7372 48488
rect 7412 48448 18220 48488
rect 18260 48448 18269 48488
rect 4919 48364 4928 48404
rect 4968 48364 5010 48404
rect 5050 48364 5092 48404
rect 5132 48364 5174 48404
rect 5214 48364 5256 48404
rect 5296 48364 5305 48404
rect 8707 48364 8716 48404
rect 8756 48364 18604 48404
rect 18644 48364 18653 48404
rect 19747 48364 19756 48404
rect 19796 48364 19805 48404
rect 20039 48364 20048 48404
rect 20088 48364 20130 48404
rect 20170 48364 20212 48404
rect 20252 48364 20294 48404
rect 20334 48364 20376 48404
rect 20416 48364 20425 48404
rect 19756 48320 19796 48364
rect 19756 48280 19892 48320
rect 11779 48196 11788 48236
rect 11828 48196 12748 48236
rect 12788 48196 12797 48236
rect 19267 48196 19276 48236
rect 19316 48196 19756 48236
rect 19796 48196 19805 48236
rect 19852 48068 19892 48280
rect 2467 48028 2476 48068
rect 2516 48028 2668 48068
rect 2708 48028 2717 48068
rect 10243 48028 10252 48068
rect 10292 48028 16204 48068
rect 16244 48028 16253 48068
rect 19267 48028 19276 48068
rect 19316 48028 19892 48068
rect 4867 47944 4876 47984
rect 4916 47944 5356 47984
rect 5396 47944 9196 47984
rect 9236 47944 9245 47984
rect 12163 47944 12172 47984
rect 12212 47944 20140 47984
rect 20180 47944 20189 47984
rect 10531 47860 10540 47900
rect 10580 47860 10636 47900
rect 10676 47860 10685 47900
rect 3679 47608 3688 47648
rect 3728 47608 3770 47648
rect 3810 47608 3852 47648
rect 3892 47608 3934 47648
rect 3974 47608 4016 47648
rect 4056 47608 4065 47648
rect 18799 47608 18808 47648
rect 18848 47608 18890 47648
rect 18930 47608 18972 47648
rect 19012 47608 19054 47648
rect 19094 47608 19136 47648
rect 19176 47608 19185 47648
rect 19651 47440 19660 47480
rect 19700 47440 19709 47480
rect 1987 47188 1996 47228
rect 2036 47188 3916 47228
rect 3956 47188 3965 47228
rect 8611 47188 8620 47228
rect 8660 47188 9196 47228
rect 9236 47188 9245 47228
rect 10531 47188 10540 47228
rect 10580 47188 15628 47228
rect 15668 47188 15677 47228
rect 19660 47144 19700 47440
rect 19555 47104 19564 47144
rect 19604 47104 19700 47144
rect 4919 46852 4928 46892
rect 4968 46852 5010 46892
rect 5050 46852 5092 46892
rect 5132 46852 5174 46892
rect 5214 46852 5256 46892
rect 5296 46852 5305 46892
rect 20039 46852 20048 46892
rect 20088 46852 20130 46892
rect 20170 46852 20212 46892
rect 20252 46852 20294 46892
rect 20334 46852 20376 46892
rect 20416 46852 20425 46892
rect 3245 46684 3340 46724
rect 3380 46684 3389 46724
rect 4483 46684 4492 46724
rect 4532 46684 4684 46724
rect 4724 46684 4733 46724
rect 5155 46684 5164 46724
rect 5204 46684 5452 46724
rect 5492 46684 5501 46724
rect 3235 46600 3244 46640
rect 3284 46600 10444 46640
rect 10484 46600 10493 46640
rect 10156 46472 10196 46600
rect 10243 46516 10252 46556
rect 10292 46516 10444 46556
rect 10484 46516 10493 46556
rect 10147 46432 10156 46472
rect 10196 46432 10205 46472
rect 13507 46432 13516 46472
rect 13556 46432 20140 46472
rect 20180 46432 20189 46472
rect 12461 46264 12556 46304
rect 12596 46264 12605 46304
rect 3679 46096 3688 46136
rect 3728 46096 3770 46136
rect 3810 46096 3852 46136
rect 3892 46096 3934 46136
rect 3974 46096 4016 46136
rect 4056 46096 4065 46136
rect 11491 46096 11500 46136
rect 11540 46096 12268 46136
rect 12308 46096 12317 46136
rect 18799 46096 18808 46136
rect 18848 46096 18890 46136
rect 18930 46096 18972 46136
rect 19012 46096 19054 46136
rect 19094 46096 19136 46136
rect 19176 46096 19185 46136
rect 5059 46012 5068 46052
rect 5108 46012 5644 46052
rect 5684 46012 5693 46052
rect 12355 46012 12364 46052
rect 12404 46012 12556 46052
rect 12596 46012 12605 46052
rect 4771 45928 4780 45968
rect 4820 45928 5644 45968
rect 5684 45928 5693 45968
rect 3907 45844 3916 45884
rect 3956 45844 5452 45884
rect 5492 45844 5501 45884
rect 4003 45760 4012 45800
rect 4052 45760 8908 45800
rect 8948 45760 8957 45800
rect 4099 45676 4108 45716
rect 4148 45676 4684 45716
rect 4724 45676 5932 45716
rect 5972 45676 5981 45716
rect 6115 45676 6124 45716
rect 6164 45676 6796 45716
rect 6836 45676 6845 45716
rect 9187 45676 9196 45716
rect 9236 45676 14860 45716
rect 14900 45676 14909 45716
rect 6124 45632 6164 45676
rect 3043 45592 3052 45632
rect 3092 45592 4492 45632
rect 4532 45592 6164 45632
rect 6691 45592 6700 45632
rect 6740 45592 8620 45632
rect 8660 45592 8669 45632
rect 2851 45508 2860 45548
rect 2900 45508 9388 45548
rect 9428 45508 9437 45548
rect 6595 45424 6604 45464
rect 6644 45424 7468 45464
rect 7508 45424 7517 45464
rect 4397 45340 4492 45380
rect 4532 45340 4541 45380
rect 4919 45340 4928 45380
rect 4968 45340 5010 45380
rect 5050 45340 5092 45380
rect 5132 45340 5174 45380
rect 5214 45340 5256 45380
rect 5296 45340 5305 45380
rect 6883 45340 6892 45380
rect 6932 45340 7564 45380
rect 7604 45340 7613 45380
rect 20039 45340 20048 45380
rect 20088 45340 20130 45380
rect 20170 45340 20212 45380
rect 20252 45340 20294 45380
rect 20334 45340 20376 45380
rect 20416 45340 20425 45380
rect 21187 45256 21196 45296
rect 21236 45256 21388 45296
rect 21428 45256 21437 45296
rect 5443 45172 5452 45212
rect 5492 45172 5644 45212
rect 5684 45172 5693 45212
rect 18019 45172 18028 45212
rect 18068 45172 18892 45212
rect 18932 45172 18941 45212
rect 13987 44920 13996 44960
rect 14036 44920 14188 44960
rect 14228 44920 14380 44960
rect 14420 44920 14429 44960
rect 21283 44920 21292 44960
rect 21332 44920 21388 44960
rect 21428 44920 21437 44960
rect 1987 44752 1996 44792
rect 2036 44752 2668 44792
rect 2708 44752 2717 44792
rect 5260 44668 6412 44708
rect 6452 44668 6461 44708
rect 5260 44624 5300 44668
rect 3679 44584 3688 44624
rect 3728 44584 3770 44624
rect 3810 44584 3852 44624
rect 3892 44584 3934 44624
rect 3974 44584 4016 44624
rect 4056 44584 4065 44624
rect 5251 44584 5260 44624
rect 5300 44584 5309 44624
rect 6211 44584 6220 44624
rect 6260 44584 6508 44624
rect 6548 44584 6557 44624
rect 18799 44584 18808 44624
rect 18848 44584 18890 44624
rect 18930 44584 18972 44624
rect 19012 44584 19054 44624
rect 19094 44584 19136 44624
rect 19176 44584 19185 44624
rect 5443 44500 5452 44540
rect 5492 44500 5644 44540
rect 5684 44500 6412 44540
rect 6452 44500 6461 44540
rect 4003 44416 4012 44456
rect 4052 44416 8716 44456
rect 8756 44416 8765 44456
rect 5059 44332 5068 44372
rect 5108 44332 5644 44372
rect 5684 44332 5693 44372
rect 5923 44332 5932 44372
rect 5972 44332 6508 44372
rect 6548 44332 6557 44372
rect 5251 44248 5260 44288
rect 5300 44248 5932 44288
rect 5972 44248 5981 44288
rect 9859 44164 9868 44204
rect 9908 44164 9964 44204
rect 10004 44164 10013 44204
rect 13603 44164 13612 44204
rect 13652 44164 15628 44204
rect 15668 44164 15677 44204
rect 4483 44080 4492 44120
rect 4532 44080 5452 44120
rect 5492 44080 5501 44120
rect 6499 44080 6508 44120
rect 6548 44080 6796 44120
rect 6836 44080 6845 44120
rect 10531 44080 10540 44120
rect 10580 44080 10732 44120
rect 10772 44080 10781 44120
rect 4291 43996 4300 44036
rect 4340 43996 4876 44036
rect 4916 43996 4925 44036
rect 14947 43996 14956 44036
rect 14996 43996 17260 44036
rect 17300 43996 17309 44036
rect 3907 43912 3916 43952
rect 3956 43912 6796 43952
rect 6836 43912 6845 43952
rect 4919 43828 4928 43868
rect 4968 43828 5010 43868
rect 5050 43828 5092 43868
rect 5132 43828 5174 43868
rect 5214 43828 5256 43868
rect 5296 43828 5305 43868
rect 5443 43828 5452 43868
rect 5492 43828 5836 43868
rect 5876 43828 5885 43868
rect 20039 43828 20048 43868
rect 20088 43828 20130 43868
rect 20170 43828 20212 43868
rect 20252 43828 20294 43868
rect 20334 43828 20376 43868
rect 20416 43828 20425 43868
rect 4579 43660 4588 43700
rect 4628 43660 4780 43700
rect 4820 43660 4829 43700
rect 5251 43660 5260 43700
rect 5300 43660 5644 43700
rect 5684 43660 5693 43700
rect 6787 43660 6796 43700
rect 6836 43660 7084 43700
rect 7124 43660 7133 43700
rect 4483 43576 4492 43616
rect 4532 43576 5356 43616
rect 5396 43576 5405 43616
rect 6499 43576 6508 43616
rect 6548 43576 8428 43616
rect 8468 43576 8477 43616
rect 3619 43492 3628 43532
rect 3668 43492 7660 43532
rect 7700 43492 7709 43532
rect 10925 43492 11020 43532
rect 11060 43492 11069 43532
rect 6403 43408 6412 43448
rect 6452 43408 6508 43448
rect 6548 43408 6557 43448
rect 5539 43324 5548 43364
rect 5588 43324 5740 43364
rect 5780 43324 5789 43364
rect 6115 43324 6124 43364
rect 6164 43324 6700 43364
rect 6740 43324 6749 43364
rect 14851 43324 14860 43364
rect 14900 43324 15052 43364
rect 15092 43324 15101 43364
rect 2093 43240 2188 43280
rect 2228 43240 2237 43280
rect 4003 43240 4012 43280
rect 4052 43240 4436 43280
rect 4867 43240 4876 43280
rect 4916 43240 5932 43280
rect 5972 43240 5981 43280
rect 12912 43240 12940 43280
rect 12980 43240 13036 43280
rect 13076 43240 13085 43280
rect 15235 43240 15244 43280
rect 15284 43240 15476 43280
rect 18787 43240 18796 43280
rect 18836 43240 18876 43280
rect 20611 43240 20620 43280
rect 20660 43240 20908 43280
rect 20948 43240 20957 43280
rect 4396 43196 4436 43240
rect 4396 43156 4628 43196
rect 1987 43072 1996 43112
rect 2036 43072 2572 43112
rect 2612 43072 2621 43112
rect 3679 43072 3688 43112
rect 3728 43072 3770 43112
rect 3810 43072 3852 43112
rect 3892 43072 3934 43112
rect 3974 43072 4016 43112
rect 4056 43072 4065 43112
rect 4291 43072 4300 43112
rect 4340 43072 4396 43112
rect 4436 43072 4445 43112
rect 4588 42860 4628 43156
rect 15436 43112 15476 43240
rect 18796 43196 18836 43240
rect 5539 43072 5548 43112
rect 5588 43072 5932 43112
rect 5972 43072 5981 43112
rect 13027 43072 13036 43112
rect 13076 43072 13324 43112
rect 13364 43072 13373 43112
rect 14851 43072 14860 43112
rect 14900 43072 15476 43112
rect 18700 43156 18836 43196
rect 14947 42988 14956 43028
rect 14996 42988 15244 43028
rect 15284 42988 15293 43028
rect 18700 42944 18740 43156
rect 18799 43072 18808 43112
rect 18848 43072 18890 43112
rect 18930 43072 18972 43112
rect 19012 43072 19054 43112
rect 19094 43072 19136 43112
rect 19176 43072 19185 43112
rect 5923 42904 5932 42944
rect 5972 42904 6316 42944
rect 6356 42904 6365 42944
rect 15043 42904 15052 42944
rect 15092 42904 15820 42944
rect 15860 42904 15869 42944
rect 18700 42904 18796 42944
rect 18836 42904 18845 42944
rect 4579 42820 4588 42860
rect 4628 42820 4637 42860
rect 5155 42820 5164 42860
rect 5204 42820 5836 42860
rect 5876 42820 5885 42860
rect 13027 42820 13036 42860
rect 13076 42820 13420 42860
rect 13460 42820 13469 42860
rect 14371 42820 14380 42860
rect 14420 42820 14429 42860
rect 6883 42736 6892 42776
rect 6932 42736 7180 42776
rect 7220 42736 7229 42776
rect 10435 42736 10444 42776
rect 10484 42736 13804 42776
rect 13844 42736 13853 42776
rect 4675 42652 4684 42692
rect 4724 42652 4733 42692
rect 11587 42652 11596 42692
rect 11636 42652 14188 42692
rect 14228 42652 14237 42692
rect 4684 42608 4724 42652
rect 4684 42568 7756 42608
rect 7796 42568 7805 42608
rect 10819 42400 10828 42440
rect 10868 42400 13708 42440
rect 13748 42400 13757 42440
rect 4919 42316 4928 42356
rect 4968 42316 5010 42356
rect 5050 42316 5092 42356
rect 5132 42316 5174 42356
rect 5214 42316 5256 42356
rect 5296 42316 5305 42356
rect 13603 42316 13612 42356
rect 13652 42316 13661 42356
rect 13612 42272 13652 42316
rect 14380 42272 14420 42820
rect 16003 42652 16012 42692
rect 16052 42652 16396 42692
rect 16436 42652 16445 42692
rect 15427 42484 15436 42524
rect 15476 42484 15820 42524
rect 15860 42484 15869 42524
rect 20039 42316 20048 42356
rect 20088 42316 20130 42356
rect 20170 42316 20212 42356
rect 20252 42316 20294 42356
rect 20334 42316 20376 42356
rect 20416 42316 20425 42356
rect 13612 42232 13708 42272
rect 13748 42232 13757 42272
rect 14380 42232 14476 42272
rect 14516 42232 14525 42272
rect 11107 42064 11116 42104
rect 11156 42064 15820 42104
rect 15860 42064 18604 42104
rect 18644 42064 18653 42104
rect 13987 41980 13996 42020
rect 14036 41980 16300 42020
rect 16340 41980 16588 42020
rect 16628 41980 16637 42020
rect 1987 41896 1996 41936
rect 2036 41896 2284 41936
rect 2324 41896 2333 41936
rect 12739 41896 12748 41936
rect 12788 41896 12940 41936
rect 12980 41896 12989 41936
rect 15619 41896 15628 41936
rect 15668 41896 16108 41936
rect 16148 41896 16157 41936
rect 4483 41812 4492 41852
rect 4532 41812 4780 41852
rect 4820 41812 5356 41852
rect 5396 41812 5405 41852
rect 15235 41812 15244 41852
rect 15284 41812 15820 41852
rect 15860 41812 15869 41852
rect 2467 41728 2476 41768
rect 2516 41728 10252 41768
rect 10292 41728 10301 41768
rect 14179 41728 14188 41768
rect 14228 41728 16684 41768
rect 16724 41728 16733 41768
rect 13795 41644 13804 41684
rect 13844 41644 16492 41684
rect 16532 41644 16541 41684
rect 3679 41560 3688 41600
rect 3728 41560 3770 41600
rect 3810 41560 3852 41600
rect 3892 41560 3934 41600
rect 3974 41560 4016 41600
rect 4056 41560 4065 41600
rect 4291 41560 4300 41600
rect 4340 41560 4588 41600
rect 4628 41560 4637 41600
rect 18799 41560 18808 41600
rect 18848 41560 18890 41600
rect 18930 41560 18972 41600
rect 19012 41560 19054 41600
rect 19094 41560 19136 41600
rect 19176 41560 19185 41600
rect 9283 41476 9292 41516
rect 9332 41476 10828 41516
rect 10868 41476 10877 41516
rect 14563 41476 14572 41516
rect 14612 41476 15820 41516
rect 15860 41476 15869 41516
rect 4493 41392 4588 41432
rect 4628 41392 4637 41432
rect 14179 41392 14188 41432
rect 14228 41392 17548 41432
rect 17588 41392 17597 41432
rect 3043 41308 3052 41348
rect 3092 41308 3148 41348
rect 3188 41308 3197 41348
rect 4771 41308 4780 41348
rect 4820 41308 5356 41348
rect 5396 41308 6124 41348
rect 6164 41308 6173 41348
rect 2275 41224 2284 41264
rect 2324 41224 8044 41264
rect 8084 41224 8093 41264
rect 5933 41140 6028 41180
rect 6068 41140 6077 41180
rect 10147 41140 10156 41180
rect 10196 41140 11020 41180
rect 11060 41140 11069 41180
rect 5155 41056 5164 41096
rect 5204 41056 6124 41096
rect 6164 41056 6173 41096
rect 6307 41056 6316 41096
rect 6356 41056 7756 41096
rect 7796 41056 7805 41096
rect 10723 41056 10732 41096
rect 10772 41056 10924 41096
rect 10964 41056 11596 41096
rect 11636 41056 11645 41096
rect 14179 41056 14188 41096
rect 14228 41056 16492 41096
rect 16532 41056 16541 41096
rect 15916 41012 15956 41056
rect 4675 40972 4684 41012
rect 4724 40972 6124 41012
rect 6164 40972 6173 41012
rect 10531 40972 10540 41012
rect 10580 40972 10732 41012
rect 10772 40972 10781 41012
rect 15043 40972 15052 41012
rect 15092 40972 15436 41012
rect 15476 40972 15485 41012
rect 15907 40972 15916 41012
rect 15956 40972 15996 41012
rect 4099 40888 4108 40928
rect 4148 40888 9196 40928
rect 9236 40888 11980 40928
rect 12020 40888 12029 40928
rect 2179 40804 2188 40844
rect 2228 40804 2380 40844
rect 2420 40804 2429 40844
rect 4919 40804 4928 40844
rect 4968 40804 5010 40844
rect 5050 40804 5092 40844
rect 5132 40804 5174 40844
rect 5214 40804 5256 40844
rect 5296 40804 5305 40844
rect 6115 40804 6124 40844
rect 6164 40804 7084 40844
rect 7124 40804 7133 40844
rect 10339 40804 10348 40844
rect 10388 40804 10540 40844
rect 10580 40804 10589 40844
rect 11299 40804 11308 40844
rect 11348 40804 12652 40844
rect 12692 40804 12701 40844
rect 12931 40804 12940 40844
rect 12980 40804 16492 40844
rect 16532 40804 17260 40844
rect 17300 40804 17309 40844
rect 20039 40804 20048 40844
rect 20088 40804 20130 40844
rect 20170 40804 20212 40844
rect 20252 40804 20294 40844
rect 20334 40804 20376 40844
rect 20416 40804 20425 40844
rect 1421 40720 1516 40760
rect 1556 40720 1565 40760
rect 3139 40720 3148 40760
rect 3188 40720 3532 40760
rect 3572 40720 6028 40760
rect 6068 40720 6077 40760
rect 14563 40720 14572 40760
rect 14612 40720 15052 40760
rect 15092 40720 15101 40760
rect 5059 40636 5068 40676
rect 5108 40636 7372 40676
rect 7412 40636 7421 40676
rect 9763 40636 9772 40676
rect 9812 40636 9821 40676
rect 9772 40592 9812 40636
rect 7171 40552 7180 40592
rect 7220 40552 7229 40592
rect 9772 40552 9964 40592
rect 10004 40552 10013 40592
rect 13219 40552 13228 40592
rect 13268 40552 13996 40592
rect 14036 40552 14045 40592
rect 7180 40508 7220 40552
rect 4579 40468 4588 40508
rect 4628 40468 5164 40508
rect 5204 40468 5644 40508
rect 5684 40468 5693 40508
rect 6019 40468 6028 40508
rect 6068 40468 7124 40508
rect 7180 40468 7372 40508
rect 7412 40468 7421 40508
rect 12355 40468 12364 40508
rect 12404 40468 15820 40508
rect 15860 40468 15869 40508
rect 7084 40424 7124 40468
rect 5251 40384 5260 40424
rect 5300 40384 6124 40424
rect 6164 40384 6173 40424
rect 7084 40384 9772 40424
rect 9812 40384 9821 40424
rect 13228 40384 13996 40424
rect 14036 40384 14045 40424
rect 18029 40384 18124 40424
rect 18164 40384 18173 40424
rect 13228 40340 13268 40384
rect 5731 40300 5740 40340
rect 5780 40300 8908 40340
rect 8948 40300 8957 40340
rect 10051 40300 10060 40340
rect 10100 40300 10196 40340
rect 12749 40300 12844 40340
rect 12884 40300 12893 40340
rect 13188 40300 13228 40340
rect 13268 40300 13277 40340
rect 13411 40300 13420 40340
rect 13460 40300 15436 40340
rect 15476 40300 15485 40340
rect 3523 40216 3532 40256
rect 3572 40216 3628 40256
rect 3668 40216 3677 40256
rect 5635 40216 5644 40256
rect 5684 40216 6892 40256
rect 6932 40216 6941 40256
rect 8803 40216 8812 40256
rect 8852 40216 9196 40256
rect 9236 40216 9245 40256
rect 10156 40172 10196 40300
rect 11971 40216 11980 40256
rect 12020 40216 12556 40256
rect 12596 40216 12605 40256
rect 6691 40132 6700 40172
rect 6740 40132 7084 40172
rect 7124 40132 7133 40172
rect 10060 40132 10196 40172
rect 11587 40132 11596 40172
rect 11636 40132 12940 40172
rect 12980 40132 12989 40172
rect 3679 40048 3688 40088
rect 3728 40048 3770 40088
rect 3810 40048 3852 40088
rect 3892 40048 3934 40088
rect 3974 40048 4016 40088
rect 4056 40048 4065 40088
rect 4867 40048 4876 40088
rect 4916 40048 8044 40088
rect 8084 40048 8093 40088
rect 10060 40004 10100 40132
rect 18799 40048 18808 40088
rect 18848 40048 18890 40088
rect 18930 40048 18972 40088
rect 19012 40048 19054 40088
rect 19094 40048 19136 40088
rect 19176 40048 19185 40088
rect 6115 39964 6124 40004
rect 6164 39964 7660 40004
rect 7700 39964 7709 40004
rect 10060 39964 10348 40004
rect 10388 39964 10397 40004
rect 11971 39964 11980 40004
rect 12020 39964 15436 40004
rect 15476 39964 15485 40004
rect 15811 39964 15820 40004
rect 15860 39964 17164 40004
rect 17204 39964 17213 40004
rect 8611 39880 8620 39920
rect 8660 39880 18508 39920
rect 18548 39880 18557 39920
rect 5155 39796 5164 39836
rect 5204 39796 6796 39836
rect 6836 39796 6845 39836
rect 10243 39796 10252 39836
rect 10292 39796 10444 39836
rect 10484 39796 10493 39836
rect 11491 39796 11500 39836
rect 11540 39796 18124 39836
rect 18164 39796 18892 39836
rect 18932 39796 18941 39836
rect 4483 39712 4492 39752
rect 4532 39712 7084 39752
rect 7124 39712 7133 39752
rect 10051 39712 10060 39752
rect 10100 39712 10924 39752
rect 10964 39712 10973 39752
rect 12259 39712 12268 39752
rect 12308 39712 12364 39752
rect 12404 39712 12413 39752
rect 12845 39712 12940 39752
rect 12980 39712 12989 39752
rect 13411 39712 13420 39752
rect 13460 39712 13516 39752
rect 13556 39712 13565 39752
rect 16867 39712 16876 39752
rect 16916 39712 18124 39752
rect 18164 39712 18173 39752
rect 2947 39628 2956 39668
rect 2996 39628 5068 39668
rect 5108 39628 5117 39668
rect 6499 39628 6508 39668
rect 6548 39628 17068 39668
rect 17108 39628 17117 39668
rect 17251 39628 17260 39668
rect 17300 39628 17548 39668
rect 17588 39628 17597 39668
rect 1891 39544 1900 39584
rect 1940 39544 2284 39584
rect 2324 39544 2333 39584
rect 4387 39544 4396 39584
rect 4436 39544 4972 39584
rect 5012 39544 5021 39584
rect 10147 39544 10156 39584
rect 10196 39544 11020 39584
rect 11060 39544 11069 39584
rect 12355 39544 12364 39584
rect 12404 39544 12652 39584
rect 12692 39544 12701 39584
rect 13027 39544 13036 39584
rect 13076 39544 14092 39584
rect 14132 39544 14141 39584
rect 12652 39500 12692 39544
rect 4291 39460 4300 39500
rect 4340 39460 4492 39500
rect 4532 39460 4541 39500
rect 5155 39460 5164 39500
rect 5204 39460 6220 39500
rect 6260 39460 6269 39500
rect 6691 39460 6700 39500
rect 6740 39460 6988 39500
rect 7028 39460 7037 39500
rect 12652 39460 14476 39500
rect 14516 39460 14525 39500
rect 6019 39376 6028 39416
rect 6068 39376 6700 39416
rect 6740 39376 6749 39416
rect 9187 39376 9196 39416
rect 9236 39376 9484 39416
rect 9524 39376 9533 39416
rect 10051 39376 10060 39416
rect 10100 39376 13228 39416
rect 13268 39376 13277 39416
rect 13507 39376 13516 39416
rect 13556 39376 13708 39416
rect 13748 39376 13757 39416
rect 4205 39292 4300 39332
rect 4340 39292 4349 39332
rect 4919 39292 4928 39332
rect 4968 39292 5010 39332
rect 5050 39292 5092 39332
rect 5132 39292 5174 39332
rect 5214 39292 5256 39332
rect 5296 39292 5305 39332
rect 5347 39292 5356 39332
rect 5396 39292 5644 39332
rect 5684 39292 5693 39332
rect 20039 39292 20048 39332
rect 20088 39292 20130 39332
rect 20170 39292 20212 39332
rect 20252 39292 20294 39332
rect 20334 39292 20376 39332
rect 20416 39292 20425 39332
rect 3715 39208 3724 39248
rect 3764 39208 6988 39248
rect 7028 39208 7037 39248
rect 12643 39208 12652 39248
rect 12692 39208 13132 39248
rect 13172 39208 13804 39248
rect 13844 39208 13853 39248
rect 4300 39124 4684 39164
rect 4724 39124 4733 39164
rect 6211 39124 6220 39164
rect 6260 39124 6508 39164
rect 6548 39124 6557 39164
rect 14755 39124 14764 39164
rect 14804 39124 16876 39164
rect 16916 39124 16925 39164
rect 4300 38996 4340 39124
rect 5923 39040 5932 39080
rect 5972 39040 6604 39080
rect 6644 39040 6653 39080
rect 6883 39040 6892 39080
rect 6932 39040 7316 39080
rect 9955 39040 9964 39080
rect 10004 39040 16876 39080
rect 16916 39040 16925 39080
rect 7276 38996 7316 39040
rect 3043 38956 3052 38996
rect 3092 38956 4300 38996
rect 4340 38956 4349 38996
rect 7267 38956 7276 38996
rect 7316 38956 7325 38996
rect 7651 38956 7660 38996
rect 7700 38956 8428 38996
rect 8468 38956 8477 38996
rect 12931 38956 12940 38996
rect 12980 38956 13228 38996
rect 13268 38956 13277 38996
rect 13795 38956 13804 38996
rect 13844 38956 14380 38996
rect 14420 38956 14429 38996
rect 14476 38956 18604 38996
rect 18644 38956 18653 38996
rect 4099 38872 4108 38912
rect 4148 38872 8236 38912
rect 8276 38872 8285 38912
rect 11107 38872 11116 38912
rect 11156 38872 11308 38912
rect 11348 38872 11357 38912
rect 12739 38872 12748 38912
rect 12788 38872 13996 38912
rect 14036 38872 14045 38912
rect 8035 38788 8044 38828
rect 8084 38788 14380 38828
rect 14420 38788 14429 38828
rect 14476 38744 14516 38956
rect 15619 38872 15628 38912
rect 15668 38872 16300 38912
rect 16340 38872 16349 38912
rect 18403 38872 18412 38912
rect 18452 38872 18461 38912
rect 18412 38828 18452 38872
rect 18412 38788 18604 38828
rect 18644 38788 18653 38828
rect 13987 38704 13996 38744
rect 14036 38704 14516 38744
rect 3679 38536 3688 38576
rect 3728 38536 3770 38576
rect 3810 38536 3852 38576
rect 3892 38536 3934 38576
rect 3974 38536 4016 38576
rect 4056 38536 4065 38576
rect 18799 38536 18808 38576
rect 18848 38536 18890 38576
rect 18930 38536 18972 38576
rect 19012 38536 19054 38576
rect 19094 38536 19136 38576
rect 19176 38536 19185 38576
rect 19555 38536 19564 38576
rect 19604 38536 19613 38576
rect 19564 38492 19604 38536
rect 1315 38452 1324 38492
rect 1364 38452 5452 38492
rect 5492 38452 5644 38492
rect 5684 38452 5693 38492
rect 19180 38452 19604 38492
rect 19180 38408 19220 38452
rect 4291 38368 4300 38408
rect 4340 38368 6988 38408
rect 7028 38368 7037 38408
rect 15043 38368 15052 38408
rect 15092 38368 15101 38408
rect 15629 38368 15724 38408
rect 15764 38368 15773 38408
rect 19171 38368 19180 38408
rect 19220 38368 19229 38408
rect 15052 38324 15092 38368
rect 3235 38284 3244 38324
rect 3284 38284 3532 38324
rect 3572 38284 3581 38324
rect 15052 38284 15188 38324
rect 19459 38284 19468 38324
rect 19508 38284 19517 38324
rect 67 38200 76 38240
rect 116 38200 4300 38240
rect 4340 38200 4349 38240
rect 6211 38200 6220 38240
rect 6260 38200 7372 38240
rect 7412 38200 7421 38240
rect 13027 38200 13036 38240
rect 13076 38200 13516 38240
rect 13556 38200 13565 38240
rect 14467 38200 14476 38240
rect 14516 38200 15052 38240
rect 15092 38200 15101 38240
rect 4387 38116 4396 38156
rect 4436 38116 5740 38156
rect 5780 38116 5789 38156
rect 6979 38116 6988 38156
rect 7028 38116 7276 38156
rect 7316 38116 7325 38156
rect 10531 38116 10540 38156
rect 10580 38116 11020 38156
rect 11060 38116 11069 38156
rect 14467 38116 14476 38156
rect 14516 38116 14860 38156
rect 14900 38116 14909 38156
rect 2851 38032 2860 38072
rect 2900 38032 3052 38072
rect 3092 38032 3101 38072
rect 5827 38032 5836 38072
rect 5876 38032 6508 38072
rect 6548 38032 6557 38072
rect 6701 38032 6796 38072
rect 6836 38032 6845 38072
rect 6307 37948 6316 37988
rect 6356 37948 7084 37988
rect 7124 37948 7133 37988
rect 6508 37904 6548 37948
rect 15148 37904 15188 38284
rect 19468 38240 19508 38284
rect 16483 38200 16492 38240
rect 16532 38200 16684 38240
rect 16724 38200 16733 38240
rect 19468 38200 19604 38240
rect 18019 38116 18028 38156
rect 18068 38116 18316 38156
rect 18356 38116 18365 38156
rect 19267 38116 19276 38156
rect 19316 38116 19468 38156
rect 19508 38116 19517 38156
rect 15427 38032 15436 38072
rect 15476 38032 15532 38072
rect 15572 38032 15581 38072
rect 19564 37988 19604 38200
rect 19267 37948 19276 37988
rect 19316 37948 19604 37988
rect 19948 37948 20044 37988
rect 20084 37948 20093 37988
rect 20419 37948 20428 37988
rect 20468 37948 20564 37988
rect 6499 37864 6508 37904
rect 6548 37864 6588 37904
rect 11491 37864 11500 37904
rect 11540 37864 11692 37904
rect 11732 37864 12748 37904
rect 12788 37864 12797 37904
rect 14755 37864 14764 37904
rect 14804 37864 15188 37904
rect 4919 37780 4928 37820
rect 4968 37780 5010 37820
rect 5050 37780 5092 37820
rect 5132 37780 5174 37820
rect 5214 37780 5256 37820
rect 5296 37780 5305 37820
rect 6115 37780 6124 37820
rect 6164 37780 6412 37820
rect 6452 37780 6892 37820
rect 6932 37780 6941 37820
rect 19948 37736 19988 37948
rect 20039 37780 20048 37820
rect 20088 37780 20130 37820
rect 20170 37780 20212 37820
rect 20252 37780 20294 37820
rect 20334 37780 20376 37820
rect 20416 37780 20425 37820
rect 3811 37696 3820 37736
rect 3860 37696 9484 37736
rect 9524 37696 9533 37736
rect 19948 37696 20084 37736
rect 20044 37652 20084 37696
rect 20524 37652 20564 37948
rect 10339 37612 10348 37652
rect 10388 37612 13420 37652
rect 13460 37612 13469 37652
rect 20035 37612 20044 37652
rect 20084 37612 20093 37652
rect 20419 37612 20428 37652
rect 20468 37612 20564 37652
rect 10051 37528 10060 37568
rect 10100 37528 10540 37568
rect 10580 37528 10589 37568
rect 11299 37528 11308 37568
rect 11348 37528 17836 37568
rect 17876 37528 17885 37568
rect 18115 37528 18124 37568
rect 18164 37528 18892 37568
rect 18932 37528 18941 37568
rect 10540 37484 10580 37528
rect 3331 37444 3340 37484
rect 3380 37444 4684 37484
rect 4724 37444 4733 37484
rect 10540 37444 11692 37484
rect 11732 37444 11741 37484
rect 17261 37360 17356 37400
rect 17396 37360 17405 37400
rect 20995 37360 21004 37400
rect 21044 37360 21292 37400
rect 21332 37360 21341 37400
rect 4675 37276 4684 37316
rect 4724 37276 7276 37316
rect 7316 37276 7325 37316
rect 10253 37276 10348 37316
rect 10388 37276 10397 37316
rect 12451 37276 12460 37316
rect 12500 37276 12652 37316
rect 12692 37276 12701 37316
rect 17347 37192 17356 37232
rect 17396 37192 17836 37232
rect 17876 37192 17885 37232
rect 19171 37192 19180 37232
rect 19220 37192 19316 37232
rect 7075 37108 7084 37148
rect 7124 37108 17260 37148
rect 17300 37108 17309 37148
rect 3679 37024 3688 37064
rect 3728 37024 3770 37064
rect 3810 37024 3852 37064
rect 3892 37024 3934 37064
rect 3974 37024 4016 37064
rect 4056 37024 4065 37064
rect 17347 37024 17356 37064
rect 17396 37024 17740 37064
rect 17780 37024 17789 37064
rect 18799 37024 18808 37064
rect 18848 37024 18890 37064
rect 18930 37024 18972 37064
rect 19012 37024 19054 37064
rect 19094 37024 19136 37064
rect 19176 37024 19185 37064
rect 19276 36980 19316 37192
rect 5443 36940 5452 36980
rect 5492 36940 5932 36980
rect 5972 36940 5981 36980
rect 16675 36940 16684 36980
rect 16724 36940 16876 36980
rect 16916 36940 16925 36980
rect 19180 36940 19316 36980
rect 19180 36896 19220 36940
rect 11779 36856 11788 36896
rect 11828 36856 12748 36896
rect 12788 36856 12797 36896
rect 16579 36856 16588 36896
rect 16628 36856 18028 36896
rect 18068 36856 18892 36896
rect 18932 36856 18941 36896
rect 19171 36856 19180 36896
rect 19220 36856 19229 36896
rect 2189 36772 2284 36812
rect 2324 36772 2333 36812
rect 3523 36688 3532 36728
rect 3572 36688 3628 36728
rect 3668 36688 3677 36728
rect 11779 36688 11788 36728
rect 11828 36688 12364 36728
rect 12404 36688 12413 36728
rect 12547 36688 12556 36728
rect 12596 36688 13708 36728
rect 13748 36688 14188 36728
rect 14228 36688 14237 36728
rect 16099 36688 16108 36728
rect 16148 36688 18124 36728
rect 18164 36688 18173 36728
rect 13699 36604 13708 36644
rect 13748 36604 13804 36644
rect 13844 36604 15916 36644
rect 15956 36604 15965 36644
rect 1411 36520 1420 36560
rect 1460 36520 1612 36560
rect 1652 36520 1661 36560
rect 3427 36520 3436 36560
rect 3476 36520 3532 36560
rect 3572 36520 3581 36560
rect 13603 36520 13612 36560
rect 13652 36520 16300 36560
rect 16340 36520 16349 36560
rect 11491 36436 11500 36476
rect 11540 36436 11692 36476
rect 11732 36436 11741 36476
rect 13699 36436 13708 36476
rect 13748 36436 14668 36476
rect 14708 36436 19084 36476
rect 19124 36436 20044 36476
rect 20084 36436 20093 36476
rect 17539 36352 17548 36392
rect 17588 36352 18028 36392
rect 18068 36352 18077 36392
rect 4919 36268 4928 36308
rect 4968 36268 5010 36308
rect 5050 36268 5092 36308
rect 5132 36268 5174 36308
rect 5214 36268 5256 36308
rect 5296 36268 5305 36308
rect 7459 36268 7468 36308
rect 7508 36268 7660 36308
rect 7700 36268 7709 36308
rect 20039 36268 20048 36308
rect 20088 36268 20130 36308
rect 20170 36268 20212 36308
rect 20252 36268 20294 36308
rect 20334 36268 20376 36308
rect 20416 36268 20425 36308
rect 13411 36184 13420 36224
rect 13460 36184 13804 36224
rect 13844 36184 13853 36224
rect 4003 36100 4012 36140
rect 4052 36100 4300 36140
rect 4340 36100 4349 36140
rect 11971 36100 11980 36140
rect 12020 36100 12364 36140
rect 12404 36100 12413 36140
rect 8515 36016 8524 36056
rect 8564 36016 13516 36056
rect 13556 36016 13565 36056
rect 14371 36016 14380 36056
rect 14420 36016 14572 36056
rect 14612 36016 14621 36056
rect 15907 36016 15916 36056
rect 15956 36016 19180 36056
rect 19220 36016 19229 36056
rect 3523 35932 3532 35972
rect 3572 35932 8236 35972
rect 8276 35932 8285 35972
rect 11971 35932 11980 35972
rect 12020 35932 12748 35972
rect 12788 35932 13036 35972
rect 13076 35932 13085 35972
rect 15427 35932 15436 35972
rect 15476 35932 16300 35972
rect 16340 35932 16349 35972
rect 18595 35932 18604 35972
rect 18644 35932 21100 35972
rect 21140 35932 21149 35972
rect 3715 35848 3724 35888
rect 3764 35848 4108 35888
rect 4148 35848 4157 35888
rect 4579 35848 4588 35888
rect 4628 35848 5356 35888
rect 5396 35848 5405 35888
rect 12259 35848 12268 35888
rect 12308 35848 12460 35888
rect 12500 35848 12509 35888
rect 14851 35764 14860 35804
rect 14900 35764 14956 35804
rect 14996 35764 15005 35804
rect 17731 35764 17740 35804
rect 17780 35764 18316 35804
rect 18356 35764 18365 35804
rect 20803 35764 20812 35804
rect 20852 35764 21196 35804
rect 21236 35764 21245 35804
rect 4771 35680 4780 35720
rect 4820 35680 5356 35720
rect 5396 35680 5405 35720
rect 12355 35680 12364 35720
rect 12404 35680 12460 35720
rect 12500 35680 12509 35720
rect 18700 35680 18796 35720
rect 18836 35680 18845 35720
rect 15235 35596 15244 35636
rect 15284 35596 15820 35636
rect 15860 35596 15869 35636
rect 16771 35596 16780 35636
rect 16820 35596 17164 35636
rect 17204 35596 17213 35636
rect 3679 35512 3688 35552
rect 3728 35512 3770 35552
rect 3810 35512 3852 35552
rect 3892 35512 3934 35552
rect 3974 35512 4016 35552
rect 4056 35512 4065 35552
rect 14371 35512 14380 35552
rect 14420 35512 14860 35552
rect 14900 35512 14909 35552
rect 15821 35512 15916 35552
rect 15956 35512 15965 35552
rect 18700 35468 18740 35680
rect 18799 35512 18808 35552
rect 18848 35512 18890 35552
rect 18930 35512 18972 35552
rect 19012 35512 19054 35552
rect 19094 35512 19136 35552
rect 19176 35512 19185 35552
rect 7171 35428 7180 35468
rect 7220 35428 12980 35468
rect 18700 35428 18836 35468
rect 12940 35384 12980 35428
rect 18796 35384 18836 35428
rect 19180 35428 19564 35468
rect 19604 35428 19613 35468
rect 19180 35384 19220 35428
rect 12940 35344 15340 35384
rect 15380 35344 15389 35384
rect 18787 35344 18796 35384
rect 18836 35344 18845 35384
rect 19171 35344 19180 35384
rect 19220 35344 19229 35384
rect 1603 35260 1612 35300
rect 1652 35260 2092 35300
rect 2132 35260 2141 35300
rect 4387 35260 4396 35300
rect 4436 35260 4780 35300
rect 4820 35260 4829 35300
rect 12163 35260 12172 35300
rect 12212 35260 13420 35300
rect 13460 35260 13469 35300
rect 2947 35176 2956 35216
rect 2996 35176 4204 35216
rect 4244 35176 4253 35216
rect 16291 35176 16300 35216
rect 16340 35176 17260 35216
rect 17300 35176 17309 35216
rect 18019 35176 18028 35216
rect 18068 35176 18892 35216
rect 18932 35176 18941 35216
rect 15907 35092 15916 35132
rect 15956 35092 16588 35132
rect 16628 35092 16637 35132
rect 17443 35092 17452 35132
rect 17492 35092 18412 35132
rect 18452 35092 18461 35132
rect 1411 35008 1420 35048
rect 1460 35008 1612 35048
rect 1652 35008 1661 35048
rect 2861 35008 2956 35048
rect 2996 35008 3005 35048
rect 10531 35008 10540 35048
rect 10580 35008 11500 35048
rect 11540 35008 11549 35048
rect 13699 35008 13708 35048
rect 13748 35008 14668 35048
rect 14708 35008 14717 35048
rect 17827 34924 17836 34964
rect 17876 34924 20428 34964
rect 20468 34924 20477 34964
rect 5923 34840 5932 34880
rect 5972 34840 8908 34880
rect 8948 34840 8957 34880
rect 4919 34756 4928 34796
rect 4968 34756 5010 34796
rect 5050 34756 5092 34796
rect 5132 34756 5174 34796
rect 5214 34756 5256 34796
rect 5296 34756 5305 34796
rect 20039 34756 20048 34796
rect 20088 34756 20130 34796
rect 20170 34756 20212 34796
rect 20252 34756 20294 34796
rect 20334 34756 20376 34796
rect 20416 34756 20425 34796
rect 2659 34672 2668 34712
rect 2708 34672 7084 34712
rect 7124 34672 8812 34712
rect 8852 34672 8861 34712
rect 17923 34672 17932 34712
rect 17972 34672 18124 34712
rect 18164 34672 18173 34712
rect 1603 34588 1612 34628
rect 1652 34588 4972 34628
rect 5012 34588 5021 34628
rect 5251 34588 5260 34628
rect 5300 34588 5932 34628
rect 5972 34588 5981 34628
rect 8419 34588 8428 34628
rect 8468 34588 13516 34628
rect 13556 34588 13565 34628
rect 18883 34588 18892 34628
rect 18932 34588 20180 34628
rect 20140 34544 20180 34588
rect 2755 34504 2764 34544
rect 2804 34504 2956 34544
rect 2996 34504 4244 34544
rect 4291 34504 4300 34544
rect 4340 34504 4780 34544
rect 4820 34504 4829 34544
rect 6691 34504 6700 34544
rect 6740 34504 10732 34544
rect 10772 34504 10781 34544
rect 12365 34504 12460 34544
rect 12500 34504 12509 34544
rect 13795 34504 13804 34544
rect 13844 34504 15916 34544
rect 15956 34504 15965 34544
rect 16675 34504 16684 34544
rect 16724 34504 18988 34544
rect 19028 34504 19037 34544
rect 20131 34504 20140 34544
rect 20180 34504 20189 34544
rect 4204 34460 4244 34504
rect 3139 34420 3148 34460
rect 3188 34420 3476 34460
rect 4204 34420 4876 34460
rect 4916 34420 4925 34460
rect 9187 34420 9196 34460
rect 9236 34420 9868 34460
rect 9908 34420 9917 34460
rect 10435 34420 10444 34460
rect 10484 34420 13612 34460
rect 13652 34420 13661 34460
rect 14659 34420 14668 34460
rect 14708 34420 14956 34460
rect 14996 34420 15244 34460
rect 15284 34420 15293 34460
rect 17059 34420 17068 34460
rect 17108 34420 21196 34460
rect 21236 34420 21245 34460
rect 3331 34336 3340 34376
rect 3380 34336 3389 34376
rect 1699 34252 1708 34292
rect 1748 34252 2092 34292
rect 2132 34252 2141 34292
rect 2851 33748 2860 33788
rect 2900 33748 2909 33788
rect 1507 33664 1516 33704
rect 1556 33664 2572 33704
rect 2612 33664 2621 33704
rect 2860 33620 2900 33748
rect 3340 33704 3380 34336
rect 3436 34292 3476 34420
rect 7459 34336 7468 34376
rect 7508 34336 20140 34376
rect 20180 34336 20189 34376
rect 3436 34252 12980 34292
rect 18691 34252 18700 34292
rect 18740 34252 19468 34292
rect 19508 34252 19517 34292
rect 4003 34168 4012 34208
rect 4052 34168 4244 34208
rect 3679 34000 3688 34040
rect 3728 34000 3770 34040
rect 3810 34000 3852 34040
rect 3892 34000 3934 34040
rect 3974 34000 4016 34040
rect 4056 34000 4065 34040
rect 2947 33664 2956 33704
rect 2996 33664 3052 33704
rect 3092 33664 3101 33704
rect 3340 33664 3724 33704
rect 3764 33664 3773 33704
rect 4204 33620 4244 34168
rect 5443 34000 5452 34040
rect 5492 34000 5644 34040
rect 5684 34000 5693 34040
rect 12940 33872 12980 34252
rect 17443 34168 17452 34208
rect 17492 34168 18124 34208
rect 18164 34168 18173 34208
rect 18787 34168 18796 34208
rect 18836 34168 19316 34208
rect 17731 34084 17740 34124
rect 17780 34084 17789 34124
rect 12940 33832 13036 33872
rect 13076 33832 13085 33872
rect 17740 33788 17780 34084
rect 18799 34000 18808 34040
rect 18848 34000 18890 34040
rect 18930 34000 18972 34040
rect 19012 34000 19054 34040
rect 19094 34000 19136 34040
rect 19176 34000 19185 34040
rect 10915 33748 10924 33788
rect 10964 33748 10973 33788
rect 17731 33748 17740 33788
rect 17780 33748 17789 33788
rect 2275 33580 2284 33620
rect 2324 33580 2476 33620
rect 2516 33580 2525 33620
rect 2860 33580 3820 33620
rect 3860 33580 3869 33620
rect 4195 33580 4204 33620
rect 4244 33580 4253 33620
rect 10924 33536 10964 33748
rect 19276 33704 19316 34168
rect 19459 34084 19468 34124
rect 19508 34084 19948 34124
rect 19988 34084 19997 34124
rect 19267 33664 19276 33704
rect 19316 33664 19325 33704
rect 14851 33580 14860 33620
rect 14900 33580 19660 33620
rect 19700 33580 19709 33620
rect 1699 33496 1708 33536
rect 1748 33496 1757 33536
rect 1987 33496 1996 33536
rect 2036 33496 2860 33536
rect 2900 33496 2909 33536
rect 3139 33496 3148 33536
rect 3188 33496 3197 33536
rect 10924 33496 11348 33536
rect 15907 33496 15916 33536
rect 15956 33496 16588 33536
rect 16628 33496 16637 33536
rect 17347 33496 17356 33536
rect 17396 33496 17836 33536
rect 17876 33496 17885 33536
rect 18979 33496 18988 33536
rect 19028 33496 19852 33536
rect 19892 33496 19901 33536
rect 1708 33200 1748 33496
rect 1795 33412 1804 33452
rect 1844 33412 2228 33452
rect 2188 33284 2228 33412
rect 3148 33368 3188 33496
rect 10444 33412 11212 33452
rect 11252 33412 11261 33452
rect 2275 33328 2284 33368
rect 2324 33328 3052 33368
rect 3092 33328 3101 33368
rect 3148 33328 3340 33368
rect 3380 33328 3389 33368
rect 10444 33284 10484 33412
rect 11308 33284 11348 33496
rect 19660 33412 20044 33452
rect 20084 33412 20093 33452
rect 20611 33412 20620 33452
rect 20660 33412 20669 33452
rect 21100 33412 21196 33452
rect 21236 33412 21245 33452
rect 11587 33328 11596 33368
rect 11636 33328 12364 33368
rect 12404 33328 12413 33368
rect 2188 33244 3148 33284
rect 3188 33244 3197 33284
rect 4291 33244 4300 33284
rect 4340 33244 4349 33284
rect 4919 33244 4928 33284
rect 4968 33244 5010 33284
rect 5050 33244 5092 33284
rect 5132 33244 5174 33284
rect 5214 33244 5256 33284
rect 5296 33244 5305 33284
rect 8899 33244 8908 33284
rect 8948 33244 9484 33284
rect 9524 33244 9533 33284
rect 10147 33244 10156 33284
rect 10196 33244 10484 33284
rect 11203 33244 11212 33284
rect 11252 33244 11348 33284
rect 11395 33244 11404 33284
rect 11444 33244 13708 33284
rect 13748 33244 13757 33284
rect 18412 33244 18604 33284
rect 18644 33244 18653 33284
rect 4300 33200 4340 33244
rect 1708 33160 2092 33200
rect 2132 33160 2141 33200
rect 3043 33160 3052 33200
rect 3092 33160 4340 33200
rect 4387 33160 4396 33200
rect 4436 33160 4492 33200
rect 4532 33160 4541 33200
rect 12355 33160 12364 33200
rect 12404 33160 13228 33200
rect 13268 33160 13277 33200
rect 18115 33160 18124 33200
rect 18164 33160 18220 33200
rect 18260 33160 18269 33200
rect 1421 33076 1516 33116
rect 1556 33076 1565 33116
rect 1804 33076 2092 33116
rect 2132 33076 2141 33116
rect 7363 33100 7372 33140
rect 7412 33116 7421 33140
rect 7412 33100 7508 33116
rect 7372 33076 7508 33100
rect 12931 33076 12940 33116
rect 12980 33076 13420 33116
rect 13460 33076 13469 33116
rect 18019 33076 18028 33116
rect 18068 33076 18124 33116
rect 18164 33076 18173 33116
rect 1804 32948 1844 33076
rect 2179 32992 2188 33032
rect 2228 32992 2860 33032
rect 2900 32992 2909 33032
rect 3907 32992 3916 33032
rect 3956 32992 4204 33032
rect 4244 32992 5548 33032
rect 5588 32992 7372 33032
rect 7412 32992 7421 33032
rect 1795 32908 1804 32948
rect 1844 32908 1853 32948
rect 4301 32908 4396 32948
rect 4436 32908 4445 32948
rect 7468 32864 7508 33076
rect 9571 32992 9580 33032
rect 9620 32992 9868 33032
rect 9908 32992 9917 33032
rect 11299 32992 11308 33032
rect 11348 32992 13228 33032
rect 13268 32992 13277 33032
rect 13699 32992 13708 33032
rect 13748 32992 13757 33032
rect 13708 32948 13748 32992
rect 10915 32908 10924 32948
rect 10964 32908 13748 32948
rect 14083 32908 14092 32948
rect 14132 32908 15820 32948
rect 15860 32908 15869 32948
rect 18115 32908 18124 32948
rect 18164 32908 18220 32948
rect 18260 32908 18269 32948
rect 1603 32824 1612 32864
rect 1652 32824 2092 32864
rect 2132 32824 2141 32864
rect 4579 32824 4588 32864
rect 4628 32824 4637 32864
rect 5251 32824 5260 32864
rect 5300 32824 7084 32864
rect 7124 32824 7133 32864
rect 7468 32824 7756 32864
rect 7796 32824 7805 32864
rect 17827 32824 17836 32864
rect 17876 32824 18028 32864
rect 18068 32824 18077 32864
rect 4588 32780 4628 32824
rect 18412 32780 18452 33244
rect 19660 33200 19700 33412
rect 19747 33328 19756 33368
rect 19796 33328 20524 33368
rect 20564 33328 20573 33368
rect 20039 33244 20048 33284
rect 20088 33244 20130 33284
rect 20170 33244 20212 33284
rect 20252 33244 20294 33284
rect 20334 33244 20376 33284
rect 20416 33244 20425 33284
rect 19660 33160 20180 33200
rect 20140 33116 20180 33160
rect 20620 33116 20660 33412
rect 21100 33200 21140 33412
rect 21196 33328 21484 33368
rect 21524 33328 21533 33368
rect 21196 33284 21236 33328
rect 21187 33244 21196 33284
rect 21236 33244 21245 33284
rect 21100 33160 21484 33200
rect 21524 33160 21533 33200
rect 18595 33076 18604 33116
rect 18644 33076 18988 33116
rect 19028 33076 19037 33116
rect 20131 33076 20140 33116
rect 20180 33076 20189 33116
rect 20323 33076 20332 33116
rect 20372 33076 20660 33116
rect 18691 32992 18700 33032
rect 18740 32992 18749 33032
rect 20035 32992 20044 33032
rect 20084 32992 20524 33032
rect 20564 32992 20573 33032
rect 4387 32740 4396 32780
rect 4436 32740 4628 32780
rect 11683 32740 11692 32780
rect 11732 32740 17932 32780
rect 17972 32740 17981 32780
rect 18115 32740 18124 32780
rect 18164 32740 18452 32780
rect 67 32656 76 32696
rect 116 32656 7276 32696
rect 7316 32656 7325 32696
rect 7459 32656 7468 32696
rect 7508 32656 7660 32696
rect 7700 32656 7709 32696
rect 3679 32488 3688 32528
rect 3728 32488 3770 32528
rect 3810 32488 3852 32528
rect 3892 32488 3934 32528
rect 3974 32488 4016 32528
rect 4056 32488 4065 32528
rect 5539 32488 5548 32528
rect 5588 32488 6220 32528
rect 6260 32488 6269 32528
rect 12451 32488 12460 32528
rect 12500 32488 17260 32528
rect 17300 32488 18124 32528
rect 18164 32488 18173 32528
rect 3523 32404 3532 32444
rect 3572 32404 8044 32444
rect 8084 32404 8093 32444
rect 8611 32404 8620 32444
rect 8660 32404 9004 32444
rect 9044 32404 9053 32444
rect 18700 32360 18740 32992
rect 18883 32656 18892 32696
rect 18932 32656 19660 32696
rect 19700 32656 19709 32696
rect 18799 32488 18808 32528
rect 18848 32488 18890 32528
rect 18930 32488 18972 32528
rect 19012 32488 19054 32528
rect 19094 32488 19136 32528
rect 19176 32488 19185 32528
rect 5731 32320 5740 32360
rect 5780 32320 8044 32360
rect 8084 32320 8093 32360
rect 18700 32320 18796 32360
rect 18836 32320 18845 32360
rect 19171 32320 19180 32360
rect 19220 32320 19564 32360
rect 19604 32320 19613 32360
rect 3235 32236 3244 32276
rect 3284 32236 4300 32276
rect 4340 32236 4349 32276
rect 9283 32236 9292 32276
rect 9332 32236 9964 32276
rect 10004 32236 10013 32276
rect 10531 32236 10540 32276
rect 10580 32236 10732 32276
rect 10772 32236 10781 32276
rect 13603 32236 13612 32276
rect 13652 32236 14380 32276
rect 14420 32236 14429 32276
rect 1411 32152 1420 32192
rect 1460 32152 7028 32192
rect 11971 32152 11980 32192
rect 12020 32152 17932 32192
rect 17972 32152 17981 32192
rect 3235 32068 3244 32108
rect 3284 32068 3340 32108
rect 3380 32068 3389 32108
rect 6988 32024 7028 32152
rect 7075 32068 7084 32108
rect 7124 32068 9196 32108
rect 9236 32068 9245 32108
rect 10435 32068 10444 32108
rect 10484 32068 10828 32108
rect 10868 32068 10877 32108
rect 14755 32068 14764 32108
rect 14804 32068 15820 32108
rect 15860 32068 16108 32108
rect 16148 32068 16157 32108
rect 20515 32068 20524 32108
rect 20564 32068 20573 32108
rect 1603 31984 1612 32024
rect 1652 31984 6836 32024
rect 6988 31984 9388 32024
rect 9428 31984 9580 32024
rect 9620 31984 9629 32024
rect 10435 31984 10444 32024
rect 10484 31984 10540 32024
rect 10580 31984 10589 32024
rect 12940 31984 13804 32024
rect 13844 31984 13853 32024
rect 15907 31984 15916 32024
rect 15956 31984 19084 32024
rect 19124 31984 19133 32024
rect 19948 31984 20236 32024
rect 20276 31984 20285 32024
rect 6796 31940 6836 31984
rect 12940 31940 12980 31984
rect 2947 31900 2956 31940
rect 2996 31900 3091 31940
rect 5251 31900 5260 31940
rect 5300 31900 5309 31940
rect 5827 31900 5836 31940
rect 5876 31900 6124 31940
rect 6164 31900 6173 31940
rect 6787 31900 6796 31940
rect 6836 31900 12980 31940
rect 5260 31856 5300 31900
rect 5260 31816 5396 31856
rect 6883 31816 6892 31856
rect 6932 31816 7948 31856
rect 7988 31816 7997 31856
rect 3331 31732 3340 31772
rect 3380 31732 4780 31772
rect 4820 31732 4829 31772
rect 4919 31732 4928 31772
rect 4968 31732 5010 31772
rect 5050 31732 5092 31772
rect 5132 31732 5174 31772
rect 5214 31732 5256 31772
rect 5296 31732 5305 31772
rect 5356 31604 5396 31816
rect 13891 31648 13900 31688
rect 13940 31648 14284 31688
rect 14324 31648 14333 31688
rect 5155 31564 5164 31604
rect 5204 31564 5396 31604
rect 11107 31564 11116 31604
rect 11156 31564 16300 31604
rect 16340 31564 16349 31604
rect 19948 31520 19988 31984
rect 20039 31732 20048 31772
rect 20088 31732 20130 31772
rect 20170 31732 20212 31772
rect 20252 31732 20294 31772
rect 20334 31732 20376 31772
rect 20416 31732 20425 31772
rect 20524 31604 20564 32068
rect 20419 31564 20428 31604
rect 20468 31564 20564 31604
rect 5251 31480 5260 31520
rect 5300 31480 6892 31520
rect 6932 31480 6941 31520
rect 13123 31480 13132 31520
rect 13172 31480 18548 31520
rect 19948 31480 20044 31520
rect 20084 31480 20093 31520
rect 18508 31436 18548 31480
rect 5635 31396 5644 31436
rect 5684 31396 11308 31436
rect 11348 31396 11357 31436
rect 14179 31396 14188 31436
rect 14228 31396 16780 31436
rect 16820 31396 16829 31436
rect 18499 31396 18508 31436
rect 18548 31396 18557 31436
rect 7939 31312 7948 31352
rect 7988 31312 8236 31352
rect 8276 31312 8285 31352
rect 13795 31312 13804 31352
rect 13844 31312 14188 31352
rect 14228 31312 14237 31352
rect 15043 31312 15052 31352
rect 15092 31312 15532 31352
rect 15572 31312 15581 31352
rect 6115 31228 6124 31268
rect 6164 31228 9292 31268
rect 9332 31228 9341 31268
rect 17059 31228 17068 31268
rect 17108 31228 20180 31268
rect 5731 31144 5740 31184
rect 5780 31144 16588 31184
rect 16628 31144 16637 31184
rect 19171 31144 19180 31184
rect 19220 31144 19316 31184
rect 4195 31060 4204 31100
rect 4244 31060 4396 31100
rect 4436 31060 6796 31100
rect 6836 31060 6845 31100
rect 12067 31060 12076 31100
rect 12116 31060 16204 31100
rect 16244 31060 16253 31100
rect 3679 30976 3688 31016
rect 3728 30976 3770 31016
rect 3810 30976 3852 31016
rect 3892 30976 3934 31016
rect 3974 30976 4016 31016
rect 4056 30976 4065 31016
rect 4483 30976 4492 31016
rect 4532 30976 4876 31016
rect 4916 30976 4925 31016
rect 12835 30976 12844 31016
rect 12884 30976 16396 31016
rect 16436 30976 16445 31016
rect 18799 30976 18808 31016
rect 18848 30976 18890 31016
rect 18930 30976 18972 31016
rect 19012 30976 19054 31016
rect 19094 30976 19136 31016
rect 19176 30976 19185 31016
rect 19276 30932 19316 31144
rect 1699 30892 1708 30932
rect 1748 30892 9004 30932
rect 9044 30892 9053 30932
rect 13123 30892 13132 30932
rect 13172 30892 15532 30932
rect 15572 30892 17260 30932
rect 17300 30892 17309 30932
rect 19180 30892 19316 30932
rect 19180 30848 19220 30892
rect 4387 30808 4396 30848
rect 4436 30808 5164 30848
rect 5204 30808 5213 30848
rect 10733 30808 10828 30848
rect 10868 30808 10877 30848
rect 16387 30808 16396 30848
rect 16436 30808 16588 30848
rect 16628 30808 16637 30848
rect 16867 30808 16876 30848
rect 16916 30808 18796 30848
rect 18836 30808 18845 30848
rect 19171 30808 19180 30848
rect 19220 30808 19229 30848
rect 19363 30808 19372 30848
rect 19412 30808 19421 30848
rect 19372 30764 19412 30808
rect 3043 30724 3052 30764
rect 3092 30724 6220 30764
rect 6260 30724 7276 30764
rect 7316 30724 7325 30764
rect 12931 30724 12940 30764
rect 12980 30724 14380 30764
rect 14420 30724 18220 30764
rect 18260 30724 18269 30764
rect 19372 30724 19604 30764
rect 19564 30680 19604 30724
rect 20140 30680 20180 31228
rect 4483 30640 4492 30680
rect 4532 30640 5548 30680
rect 5588 30640 5597 30680
rect 14467 30640 14476 30680
rect 14516 30640 14764 30680
rect 14804 30640 14813 30680
rect 18499 30640 18508 30680
rect 18548 30640 19372 30680
rect 19412 30640 19421 30680
rect 19555 30640 19564 30680
rect 19604 30640 19613 30680
rect 20131 30640 20140 30680
rect 20180 30640 20189 30680
rect 3907 30556 3916 30596
rect 3956 30556 5068 30596
rect 5108 30556 5117 30596
rect 7939 30556 7948 30596
rect 7988 30556 19756 30596
rect 19796 30556 19805 30596
rect 2659 30472 2668 30512
rect 2708 30472 8908 30512
rect 8948 30472 8957 30512
rect 13123 30472 13132 30512
rect 13172 30472 13181 30512
rect 19075 30472 19084 30512
rect 19124 30472 20044 30512
rect 20084 30472 20093 30512
rect 13132 30428 13172 30472
rect 7267 30388 7276 30428
rect 7316 30388 8620 30428
rect 8660 30388 8669 30428
rect 13132 30388 14476 30428
rect 14516 30388 14525 30428
rect 18115 30388 18124 30428
rect 18164 30388 18988 30428
rect 19028 30388 19037 30428
rect 6115 30304 6124 30344
rect 6164 30304 8660 30344
rect 11779 30304 11788 30344
rect 11828 30304 12364 30344
rect 12404 30304 12413 30344
rect 13123 30304 13132 30344
rect 13172 30304 14668 30344
rect 14708 30304 14717 30344
rect 15916 30304 17068 30344
rect 17108 30304 17117 30344
rect 17923 30304 17932 30344
rect 17972 30304 20524 30344
rect 20564 30304 20573 30344
rect 1613 30220 1708 30260
rect 1748 30220 1757 30260
rect 4919 30220 4928 30260
rect 4968 30220 5010 30260
rect 5050 30220 5092 30260
rect 5132 30220 5174 30260
rect 5214 30220 5256 30260
rect 5296 30220 5305 30260
rect 7236 30220 7276 30260
rect 7316 30220 7325 30260
rect 7276 30176 7316 30220
rect 8620 30176 8660 30304
rect 15916 30260 15956 30304
rect 12259 30220 12268 30260
rect 12308 30220 14188 30260
rect 14228 30220 14237 30260
rect 14668 30220 15956 30260
rect 16013 30220 16108 30260
rect 16148 30220 16157 30260
rect 18691 30220 18700 30260
rect 18740 30220 18749 30260
rect 20039 30220 20048 30260
rect 20088 30220 20130 30260
rect 20170 30220 20212 30260
rect 20252 30220 20294 30260
rect 20334 30220 20376 30260
rect 20416 30220 20425 30260
rect 14668 30176 14708 30220
rect 18700 30176 18740 30220
rect 2860 30136 7316 30176
rect 7459 30136 7468 30176
rect 7508 30136 7756 30176
rect 7796 30136 7805 30176
rect 8620 30136 14708 30176
rect 14764 30136 15916 30176
rect 15956 30136 15965 30176
rect 18115 30136 18124 30176
rect 18164 30136 18740 30176
rect 2860 29924 2900 30136
rect 7853 30052 7948 30092
rect 7988 30052 7997 30092
rect 10243 30052 10252 30092
rect 10292 30052 10444 30092
rect 10484 30052 10493 30092
rect 12451 30052 12460 30092
rect 12500 30052 13420 30092
rect 13460 30052 13469 30092
rect 14764 30008 14804 30136
rect 5251 29968 5260 30008
rect 5300 29968 5740 30008
rect 5780 29968 5789 30008
rect 12835 29968 12844 30008
rect 12884 29968 13900 30008
rect 13940 29968 13949 30008
rect 14188 29968 14804 30008
rect 14860 30052 18028 30092
rect 18068 30052 18077 30092
rect 14188 29924 14228 29968
rect 1027 29884 1036 29924
rect 1076 29884 2900 29924
rect 8707 29884 8716 29924
rect 8756 29884 9676 29924
rect 9716 29884 9725 29924
rect 10349 29884 10444 29924
rect 10484 29884 10924 29924
rect 10964 29884 10973 29924
rect 12931 29884 12940 29924
rect 12980 29884 14188 29924
rect 14228 29884 14237 29924
rect 14860 29840 14900 30052
rect 14947 29968 14956 30008
rect 14996 29968 15436 30008
rect 15476 29968 15485 30008
rect 15715 29968 15724 30008
rect 15764 29968 17452 30008
rect 17492 29968 17501 30008
rect 18499 29968 18508 30008
rect 18548 29968 18988 30008
rect 19028 29968 19037 30008
rect 15811 29884 15820 29924
rect 15860 29884 17260 29924
rect 17300 29884 17309 29924
rect 1229 29800 1324 29840
rect 1364 29800 1373 29840
rect 1891 29800 1900 29840
rect 1940 29800 1949 29840
rect 2563 29800 2572 29840
rect 2612 29800 9100 29840
rect 9140 29800 9149 29840
rect 9283 29800 9292 29840
rect 9332 29800 10348 29840
rect 10388 29800 10636 29840
rect 10676 29800 10685 29840
rect 12931 29800 12940 29840
rect 12980 29800 14900 29840
rect 15523 29800 15532 29840
rect 15572 29800 19564 29840
rect 19604 29800 19613 29840
rect 1900 29252 1940 29800
rect 2371 29716 2380 29756
rect 2420 29716 2860 29756
rect 2900 29716 4300 29756
rect 4340 29716 4349 29756
rect 7363 29716 7372 29756
rect 7412 29716 9388 29756
rect 9428 29716 9437 29756
rect 13315 29716 13324 29756
rect 13364 29716 13420 29756
rect 13460 29716 13469 29756
rect 14467 29716 14476 29756
rect 14516 29716 14860 29756
rect 14900 29716 14909 29756
rect 17827 29716 17836 29756
rect 17876 29716 19084 29756
rect 19124 29716 19133 29756
rect 4003 29632 4012 29672
rect 4052 29632 9292 29672
rect 9332 29632 9341 29672
rect 12835 29632 12844 29672
rect 12884 29632 14956 29672
rect 14996 29632 15005 29672
rect 15427 29632 15436 29672
rect 15476 29632 15724 29672
rect 15764 29632 15773 29672
rect 19171 29632 19180 29672
rect 19220 29632 19316 29672
rect 4291 29548 4300 29588
rect 4340 29548 14860 29588
rect 14900 29548 14909 29588
rect 3679 29464 3688 29504
rect 3728 29464 3770 29504
rect 3810 29464 3852 29504
rect 3892 29464 3934 29504
rect 3974 29464 4016 29504
rect 4056 29464 4065 29504
rect 13699 29464 13708 29504
rect 13748 29464 15916 29504
rect 15956 29464 15965 29504
rect 18799 29464 18808 29504
rect 18848 29464 18890 29504
rect 18930 29464 18972 29504
rect 19012 29464 19054 29504
rect 19094 29464 19136 29504
rect 19176 29464 19185 29504
rect 19276 29420 19316 29632
rect 6115 29380 6124 29420
rect 6164 29380 6412 29420
rect 6452 29380 6461 29420
rect 8707 29380 8716 29420
rect 8756 29380 9292 29420
rect 9332 29380 9341 29420
rect 11299 29380 11308 29420
rect 11348 29380 13804 29420
rect 13844 29380 13853 29420
rect 14467 29380 14476 29420
rect 14516 29380 15916 29420
rect 15956 29380 15965 29420
rect 19180 29380 19316 29420
rect 19180 29336 19220 29380
rect 2083 29296 2092 29336
rect 2132 29296 6028 29336
rect 6068 29296 6077 29336
rect 11683 29296 11692 29336
rect 11732 29296 14956 29336
rect 14996 29296 16300 29336
rect 16340 29296 16349 29336
rect 19171 29296 19180 29336
rect 19220 29296 19229 29336
rect 1900 29212 2132 29252
rect 11971 29212 11980 29252
rect 12020 29212 12268 29252
rect 12308 29212 12317 29252
rect 12643 29212 12652 29252
rect 12692 29212 13132 29252
rect 13172 29212 13181 29252
rect 13699 29212 13708 29252
rect 13748 29212 14956 29252
rect 14996 29212 15005 29252
rect 2092 29168 2132 29212
rect 2083 29128 2092 29168
rect 2132 29128 2141 29168
rect 13315 29128 13324 29168
rect 13364 29128 13804 29168
rect 13844 29128 15724 29168
rect 15764 29128 15773 29168
rect 16099 29128 16108 29168
rect 16148 29128 21292 29168
rect 21332 29128 21341 29168
rect 2851 29044 2860 29084
rect 2900 29044 8812 29084
rect 8852 29044 8861 29084
rect 12259 29044 12268 29084
rect 12308 29044 12556 29084
rect 12596 29044 12605 29084
rect 13507 29044 13516 29084
rect 13556 29044 13612 29084
rect 13652 29044 13661 29084
rect 17251 29044 17260 29084
rect 17300 29044 17309 29084
rect 18019 29044 18028 29084
rect 18068 29044 18412 29084
rect 18452 29044 18461 29084
rect 17260 29000 17300 29044
rect 4876 28960 7372 29000
rect 7412 28960 7421 29000
rect 17260 28960 17932 29000
rect 17972 28960 17981 29000
rect 4876 28916 4916 28960
rect 4387 28876 4396 28916
rect 4436 28876 4876 28916
rect 4916 28876 4925 28916
rect 5251 28876 5260 28916
rect 5300 28876 5309 28916
rect 6115 28876 6124 28916
rect 6164 28876 10060 28916
rect 10100 28876 10109 28916
rect 10435 28876 10444 28916
rect 10484 28876 10540 28916
rect 10580 28876 10924 28916
rect 10964 28876 10973 28916
rect 15811 28876 15820 28916
rect 15860 28876 16684 28916
rect 16724 28876 16733 28916
rect 5260 28832 5300 28876
rect 1123 28792 1132 28832
rect 1172 28792 1364 28832
rect 2851 28792 2860 28832
rect 2900 28792 4012 28832
rect 4052 28792 4061 28832
rect 5260 28792 5396 28832
rect 5539 28792 5548 28832
rect 5588 28792 5644 28832
rect 5684 28792 5693 28832
rect 15715 28792 15724 28832
rect 15764 28792 15820 28832
rect 15860 28792 15869 28832
rect 1324 28580 1364 28792
rect 4919 28708 4928 28748
rect 4968 28708 5010 28748
rect 5050 28708 5092 28748
rect 5132 28708 5174 28748
rect 5214 28708 5256 28748
rect 5296 28708 5305 28748
rect 5356 28664 5396 28792
rect 5731 28708 5740 28748
rect 5780 28708 10636 28748
rect 10676 28708 10685 28748
rect 14563 28708 14572 28748
rect 14612 28708 15052 28748
rect 15092 28708 15101 28748
rect 20039 28708 20048 28748
rect 20088 28708 20130 28748
rect 20170 28708 20212 28748
rect 20252 28708 20294 28748
rect 20334 28708 20376 28748
rect 20416 28708 20425 28748
rect 4003 28624 4012 28664
rect 4052 28624 4780 28664
rect 4820 28624 4829 28664
rect 5068 28624 5396 28664
rect 10253 28624 10348 28664
rect 10388 28624 10397 28664
rect 5068 28580 5108 28624
rect 1315 28540 1324 28580
rect 1364 28540 1373 28580
rect 5059 28540 5068 28580
rect 5108 28540 5117 28580
rect 5251 28540 5260 28580
rect 5300 28540 6316 28580
rect 6356 28540 6365 28580
rect 8323 28540 8332 28580
rect 8372 28540 9196 28580
rect 9236 28540 9245 28580
rect 3139 28456 3148 28496
rect 3188 28456 11692 28496
rect 11732 28456 11741 28496
rect 1603 28372 1612 28412
rect 1652 28372 1804 28412
rect 1844 28372 1853 28412
rect 4483 28372 4492 28412
rect 4532 28372 4780 28412
rect 4820 28372 4829 28412
rect 6787 28372 6796 28412
rect 6836 28372 7852 28412
rect 7892 28372 7901 28412
rect 1804 28328 1844 28372
rect 365 28288 460 28328
rect 500 28288 509 28328
rect 1804 28288 10060 28328
rect 10100 28288 10109 28328
rect 6211 28204 6220 28244
rect 6260 28204 6604 28244
rect 6644 28204 6653 28244
rect 18403 28204 18412 28244
rect 18452 28204 18604 28244
rect 18644 28204 18653 28244
rect 20611 28204 20620 28244
rect 20660 28204 20908 28244
rect 20948 28204 20957 28244
rect 1517 28120 1612 28160
rect 1652 28120 1661 28160
rect 4579 28120 4588 28160
rect 4628 28120 5836 28160
rect 5876 28120 5885 28160
rect 16291 28036 16300 28076
rect 16340 28036 16876 28076
rect 16916 28036 16925 28076
rect 20707 28036 20716 28076
rect 20756 28036 20765 28076
rect 20716 27992 20756 28036
rect 3679 27952 3688 27992
rect 3728 27952 3770 27992
rect 3810 27952 3852 27992
rect 3892 27952 3934 27992
rect 3974 27952 4016 27992
rect 4056 27952 4065 27992
rect 6883 27952 6892 27992
rect 6932 27952 7660 27992
rect 7700 27952 10060 27992
rect 10100 27952 10109 27992
rect 14755 27952 14764 27992
rect 14804 27952 16588 27992
rect 16628 27952 16637 27992
rect 18799 27952 18808 27992
rect 18848 27952 18890 27992
rect 18930 27952 18972 27992
rect 19012 27952 19054 27992
rect 19094 27952 19136 27992
rect 19176 27952 19185 27992
rect 19267 27952 19276 27992
rect 19316 27952 19564 27992
rect 19604 27952 20140 27992
rect 20180 27952 20189 27992
rect 20716 27952 20908 27992
rect 20948 27952 20957 27992
rect 20707 27868 20716 27908
rect 20756 27868 21292 27908
rect 21332 27868 21341 27908
rect 18499 27784 18508 27824
rect 18548 27784 18892 27824
rect 18932 27784 18941 27824
rect 11011 27616 11020 27656
rect 11060 27616 11212 27656
rect 11252 27616 11261 27656
rect 11779 27616 11788 27656
rect 11828 27616 16204 27656
rect 16244 27616 16253 27656
rect 10723 27532 10732 27572
rect 10772 27532 10828 27572
rect 10868 27532 10877 27572
rect 11971 27532 11980 27572
rect 12020 27532 12172 27572
rect 12212 27532 12221 27572
rect 13699 27532 13708 27572
rect 13748 27532 16396 27572
rect 16436 27532 16445 27572
rect 18211 27532 18220 27572
rect 18260 27532 18604 27572
rect 18644 27532 18653 27572
rect 4771 27448 4780 27488
rect 4820 27448 5644 27488
rect 5684 27448 5693 27488
rect 7939 27448 7948 27488
rect 7988 27448 11788 27488
rect 11828 27448 11837 27488
rect 15139 27448 15148 27488
rect 15188 27448 15340 27488
rect 15380 27448 15389 27488
rect 4003 27364 4012 27404
rect 4052 27364 4396 27404
rect 4436 27364 5932 27404
rect 5972 27364 5981 27404
rect 11491 27364 11500 27404
rect 11540 27364 12172 27404
rect 12212 27364 12221 27404
rect 18595 27364 18604 27404
rect 18644 27364 19468 27404
rect 19508 27364 19517 27404
rect 20803 27280 20812 27320
rect 20852 27280 21292 27320
rect 21332 27280 21341 27320
rect 4919 27196 4928 27236
rect 4968 27196 5010 27236
rect 5050 27196 5092 27236
rect 5132 27196 5174 27236
rect 5214 27196 5256 27236
rect 5296 27196 5305 27236
rect 20039 27196 20048 27236
rect 20088 27196 20130 27236
rect 20170 27196 20212 27236
rect 20252 27196 20294 27236
rect 20334 27196 20376 27236
rect 20416 27196 20425 27236
rect 4387 27112 4396 27152
rect 4436 27112 4588 27152
rect 4628 27112 4637 27152
rect 11299 27112 11308 27152
rect 11348 27112 15532 27152
rect 15572 27112 15581 27152
rect 15629 27112 15724 27152
rect 15764 27112 15773 27152
rect 9283 27028 9292 27068
rect 9332 27028 16588 27068
rect 16628 27028 16637 27068
rect 19651 27028 19660 27068
rect 19700 27028 20044 27068
rect 20084 27028 20093 27068
rect 12643 26944 12652 26984
rect 12692 26944 13036 26984
rect 13076 26944 13085 26984
rect 3811 26860 3820 26900
rect 3860 26860 4300 26900
rect 4340 26860 9964 26900
rect 10004 26860 10013 26900
rect 11395 26860 11404 26900
rect 11444 26860 13804 26900
rect 13844 26860 13853 26900
rect 14659 26860 14668 26900
rect 14708 26860 15724 26900
rect 15764 26860 16492 26900
rect 16532 26860 16541 26900
rect 1795 26776 1804 26816
rect 1844 26776 7852 26816
rect 7892 26776 7901 26816
rect 4300 26732 4340 26776
rect 4291 26692 4300 26732
rect 4340 26692 4380 26732
rect 18211 26692 18220 26732
rect 18260 26692 19180 26732
rect 19220 26692 19229 26732
rect 7939 26608 7948 26648
rect 7988 26608 7997 26648
rect 12259 26608 12268 26648
rect 12308 26608 17740 26648
rect 17780 26608 17836 26648
rect 17876 26608 17885 26648
rect 7948 26564 7988 26608
rect 7276 26524 7988 26564
rect 10051 26524 10060 26564
rect 10100 26524 16108 26564
rect 16148 26524 16157 26564
rect 7276 26480 7316 26524
rect 3679 26440 3688 26480
rect 3728 26440 3770 26480
rect 3810 26440 3852 26480
rect 3892 26440 3934 26480
rect 3974 26440 4016 26480
rect 4056 26440 4065 26480
rect 7267 26440 7276 26480
rect 7316 26440 7325 26480
rect 18799 26440 18808 26480
rect 18848 26440 18890 26480
rect 18930 26440 18972 26480
rect 19012 26440 19054 26480
rect 19094 26440 19136 26480
rect 19176 26440 19185 26480
rect 2179 26356 2188 26396
rect 2228 26356 6124 26396
rect 6164 26356 6173 26396
rect 3907 26272 3916 26312
rect 3956 26272 6028 26312
rect 6068 26272 6077 26312
rect 9197 26272 9292 26312
rect 9332 26272 9341 26312
rect 13901 26272 13996 26312
rect 14036 26272 14045 26312
rect 18499 26272 18508 26312
rect 18548 26272 18796 26312
rect 18836 26272 18845 26312
rect 2860 26188 9484 26228
rect 9524 26188 9533 26228
rect 9955 26188 9964 26228
rect 10004 26188 10060 26228
rect 10100 26188 10109 26228
rect 13795 26188 13804 26228
rect 13844 26188 15436 26228
rect 15476 26188 15485 26228
rect 2860 26060 2900 26188
rect 4483 26104 4492 26144
rect 4532 26104 4541 26144
rect 8131 26104 8140 26144
rect 8180 26104 9388 26144
rect 9428 26104 10060 26144
rect 10100 26104 10109 26144
rect 12931 26104 12940 26144
rect 12980 26104 14476 26144
rect 14516 26104 14525 26144
rect 16483 26104 16492 26144
rect 16532 26104 17260 26144
rect 17300 26104 17309 26144
rect 1987 26020 1996 26060
rect 2036 26020 2900 26060
rect 4492 25892 4532 26104
rect 4579 26020 4588 26060
rect 4628 26020 7948 26060
rect 7988 26020 8524 26060
rect 8564 26020 9964 26060
rect 10004 26020 10013 26060
rect 11587 26020 11596 26060
rect 11636 26020 12268 26060
rect 12308 26020 12317 26060
rect 16579 26020 16588 26060
rect 16628 26020 16876 26060
rect 16916 26020 16925 26060
rect 20035 26020 20044 26060
rect 20084 26020 20812 26060
rect 20852 26020 20861 26060
rect 7171 25936 7180 25976
rect 7220 25936 7468 25976
rect 7508 25936 7517 25976
rect 4492 25852 4684 25892
rect 4724 25852 4733 25892
rect 7555 25852 7564 25892
rect 7604 25852 9196 25892
rect 9236 25852 9245 25892
rect 13123 25852 13132 25892
rect 13172 25852 13516 25892
rect 13556 25852 13565 25892
rect 4195 25768 4204 25808
rect 4244 25768 5644 25808
rect 5684 25768 5693 25808
rect 10051 25768 10060 25808
rect 10100 25768 18796 25808
rect 18836 25768 18845 25808
rect 4003 25684 4012 25724
rect 4052 25684 4204 25724
rect 4244 25684 4253 25724
rect 4919 25684 4928 25724
rect 4968 25684 5010 25724
rect 5050 25684 5092 25724
rect 5132 25684 5174 25724
rect 5214 25684 5256 25724
rect 5296 25684 5305 25724
rect 20039 25684 20048 25724
rect 20088 25684 20130 25724
rect 20170 25684 20212 25724
rect 20252 25684 20294 25724
rect 20334 25684 20376 25724
rect 20416 25684 20425 25724
rect 163 25600 172 25640
rect 212 25600 3628 25640
rect 3668 25600 3677 25640
rect 3811 25600 3820 25640
rect 3860 25600 5740 25640
rect 5780 25600 5789 25640
rect 6787 25600 6796 25640
rect 6836 25600 7084 25640
rect 7124 25600 7133 25640
rect 9091 25600 9100 25640
rect 9140 25600 9676 25640
rect 9716 25600 9725 25640
rect 67 25516 76 25556
rect 116 25516 4972 25556
rect 5012 25516 5021 25556
rect 7267 25516 7276 25556
rect 7316 25516 9140 25556
rect 9100 25472 9140 25516
rect 2947 25432 2956 25472
rect 2996 25432 3916 25472
rect 3956 25432 3965 25472
rect 9091 25432 9100 25472
rect 9140 25432 9149 25472
rect 20429 25432 20524 25472
rect 20564 25432 20573 25472
rect 2851 25348 2860 25388
rect 2900 25348 4876 25388
rect 4916 25348 6700 25388
rect 6740 25348 6749 25388
rect 9379 25348 9388 25388
rect 9428 25348 9772 25388
rect 9812 25348 9821 25388
rect 19180 25348 19276 25388
rect 19316 25348 19325 25388
rect 1891 25264 1900 25304
rect 1940 25264 9292 25304
rect 9332 25264 9341 25304
rect 9955 25264 9964 25304
rect 10004 25264 10060 25304
rect 10100 25264 10109 25304
rect 15331 25264 15340 25304
rect 15380 25264 16204 25304
rect 16244 25264 16253 25304
rect 1603 25180 1612 25220
rect 1652 25180 2476 25220
rect 2516 25180 2525 25220
rect 7565 25180 7660 25220
rect 7700 25180 7709 25220
rect 19180 25136 19220 25348
rect 19267 25180 19276 25220
rect 19316 25180 19468 25220
rect 19508 25180 19517 25220
rect 1315 25096 1324 25136
rect 1364 25096 2092 25136
rect 2132 25096 2141 25136
rect 3235 25096 3244 25136
rect 3284 25096 5972 25136
rect 19180 25096 19508 25136
rect 5932 25052 5972 25096
rect 19468 25052 19508 25096
rect 1795 25012 1804 25052
rect 1844 25012 5260 25052
rect 5300 25012 5309 25052
rect 5923 25012 5932 25052
rect 5972 25012 5981 25052
rect 11971 25012 11980 25052
rect 12020 25012 12364 25052
rect 12404 25012 12413 25052
rect 17635 25012 17644 25052
rect 17684 25012 17836 25052
rect 17876 25012 17885 25052
rect 19459 25012 19468 25052
rect 19508 25012 19517 25052
rect 19651 25012 19660 25052
rect 19700 25012 20044 25052
rect 20084 25012 20093 25052
rect 3679 24928 3688 24968
rect 3728 24928 3770 24968
rect 3810 24928 3852 24968
rect 3892 24928 3934 24968
rect 3974 24928 4016 24968
rect 4056 24928 4065 24968
rect 6979 24928 6988 24968
rect 7028 24928 7084 24968
rect 7124 24928 7133 24968
rect 7459 24928 7468 24968
rect 7508 24928 11596 24968
rect 11636 24928 11645 24968
rect 18799 24928 18808 24968
rect 18848 24928 18890 24968
rect 18930 24928 18972 24968
rect 19012 24928 19054 24968
rect 19094 24928 19136 24968
rect 19176 24928 19185 24968
rect 2851 24844 2860 24884
rect 2900 24844 4204 24884
rect 4244 24844 4253 24884
rect 8611 24844 8620 24884
rect 8660 24844 8812 24884
rect 8852 24844 8861 24884
rect 16579 24844 16588 24884
rect 16628 24844 20140 24884
rect 20180 24844 20189 24884
rect 3043 24760 3052 24800
rect 3092 24760 3628 24800
rect 3668 24760 3677 24800
rect 14467 24760 14476 24800
rect 14516 24760 18124 24800
rect 18164 24760 18173 24800
rect 3139 24676 3148 24716
rect 3188 24676 3244 24716
rect 3284 24676 3293 24716
rect 16963 24676 16972 24716
rect 17012 24676 18028 24716
rect 18068 24676 18077 24716
rect 6979 24592 6988 24632
rect 7028 24592 7948 24632
rect 7988 24592 7997 24632
rect 14947 24592 14956 24632
rect 14996 24592 15436 24632
rect 15476 24592 15485 24632
rect 16675 24592 16684 24632
rect 16724 24592 17260 24632
rect 17300 24592 17309 24632
rect 18115 24592 18124 24632
rect 18164 24592 18604 24632
rect 18644 24592 18653 24632
rect 20611 24592 20620 24632
rect 20660 24592 21004 24632
rect 21044 24592 21053 24632
rect 4579 24508 4588 24548
rect 4628 24508 6028 24548
rect 6068 24508 6077 24548
rect 7373 24508 7468 24548
rect 7508 24508 7517 24548
rect 7468 24464 7508 24508
rect 4867 24424 4876 24464
rect 4916 24424 7508 24464
rect 17539 24424 17548 24464
rect 17588 24424 20524 24464
rect 20564 24424 20573 24464
rect 2851 24340 2860 24380
rect 2900 24340 7564 24380
rect 7604 24340 7613 24380
rect 12931 24340 12940 24380
rect 12980 24340 13228 24380
rect 13268 24340 13277 24380
rect 4919 24172 4928 24212
rect 4968 24172 5010 24212
rect 5050 24172 5092 24212
rect 5132 24172 5174 24212
rect 5214 24172 5256 24212
rect 5296 24172 5305 24212
rect 13123 24172 13132 24212
rect 13172 24172 13324 24212
rect 13364 24172 13373 24212
rect 20039 24172 20048 24212
rect 20088 24172 20130 24212
rect 20170 24172 20212 24212
rect 20252 24172 20294 24212
rect 20334 24172 20376 24212
rect 20416 24172 20425 24212
rect 3523 24004 3532 24044
rect 3572 24004 3916 24044
rect 3956 24004 3965 24044
rect 15715 24004 15724 24044
rect 15764 24004 16492 24044
rect 16532 24004 16541 24044
rect 1987 23920 1996 23960
rect 2036 23920 4972 23960
rect 5012 23920 5021 23960
rect 3619 23752 3628 23792
rect 3668 23752 8332 23792
rect 8372 23752 8381 23792
rect 10243 23752 10252 23792
rect 10292 23752 13996 23792
rect 14036 23752 14045 23792
rect 14851 23752 14860 23792
rect 14900 23752 16396 23792
rect 16436 23752 16445 23792
rect 18307 23752 18316 23792
rect 18356 23752 18604 23792
rect 18644 23752 18653 23792
rect 3331 23668 3340 23708
rect 3380 23668 3532 23708
rect 3572 23668 3581 23708
rect 9091 23668 9100 23708
rect 9140 23668 9676 23708
rect 9716 23668 9725 23708
rect 14179 23668 14188 23708
rect 14228 23668 18508 23708
rect 18548 23668 18557 23708
rect 3715 23584 3724 23624
rect 3764 23584 4684 23624
rect 4724 23584 4733 23624
rect 9955 23584 9964 23624
rect 10004 23584 10252 23624
rect 10292 23584 10301 23624
rect 17251 23584 17260 23624
rect 17300 23584 18028 23624
rect 18068 23584 19852 23624
rect 19892 23584 19901 23624
rect 4301 23500 4396 23540
rect 4436 23500 4445 23540
rect 12940 23500 18124 23540
rect 18164 23500 18173 23540
rect 12940 23456 12980 23500
rect 3679 23416 3688 23456
rect 3728 23416 3770 23456
rect 3810 23416 3852 23456
rect 3892 23416 3934 23456
rect 3974 23416 4016 23456
rect 4056 23416 4065 23456
rect 12451 23416 12460 23456
rect 12500 23416 12940 23456
rect 12980 23416 12989 23456
rect 15907 23416 15916 23456
rect 15956 23416 16396 23456
rect 16436 23416 16445 23456
rect 17827 23416 17836 23456
rect 17876 23416 18604 23456
rect 18644 23416 18653 23456
rect 18799 23416 18808 23456
rect 18848 23416 18890 23456
rect 18930 23416 18972 23456
rect 19012 23416 19054 23456
rect 19094 23416 19136 23456
rect 19176 23416 19185 23456
rect 3052 23332 10156 23372
rect 10196 23332 10205 23372
rect 18115 23332 18124 23372
rect 18164 23332 18220 23372
rect 18260 23332 18269 23372
rect 18403 23332 18412 23372
rect 18452 23332 18548 23372
rect 2285 23248 2380 23288
rect 2420 23248 2429 23288
rect 2179 23164 2188 23204
rect 2228 23164 2860 23204
rect 2900 23164 2909 23204
rect 3052 23060 3092 23332
rect 3427 23248 3436 23288
rect 3476 23248 3820 23288
rect 3860 23248 3869 23288
rect 4003 23248 4012 23288
rect 4052 23248 4204 23288
rect 4244 23248 4253 23288
rect 13795 23248 13804 23288
rect 13844 23248 14284 23288
rect 14324 23248 14333 23288
rect 16013 23248 16108 23288
rect 16148 23248 16157 23288
rect 18508 23204 18548 23332
rect 18595 23248 18604 23288
rect 18644 23248 18892 23288
rect 18932 23248 18941 23288
rect 3523 23164 3532 23204
rect 3572 23164 3724 23204
rect 3764 23164 3773 23204
rect 5923 23164 5932 23204
rect 5972 23164 6124 23204
rect 6164 23164 6173 23204
rect 7843 23164 7852 23204
rect 7892 23164 8620 23204
rect 8660 23164 9004 23204
rect 9044 23164 9676 23204
rect 9716 23164 9725 23204
rect 13411 23164 13420 23204
rect 13460 23164 13708 23204
rect 13748 23164 13757 23204
rect 14947 23164 14956 23204
rect 14996 23164 17396 23204
rect 17443 23164 17452 23204
rect 17492 23164 18412 23204
rect 18452 23164 18461 23204
rect 18508 23164 18796 23204
rect 18836 23164 18845 23204
rect 17356 23120 17396 23164
rect 3235 23080 3244 23120
rect 3284 23080 3436 23120
rect 3476 23080 3485 23120
rect 3907 23080 3916 23120
rect 3956 23080 4204 23120
rect 4244 23080 4253 23120
rect 5731 23080 5740 23120
rect 5780 23080 6124 23120
rect 6164 23080 6173 23120
rect 7363 23080 7372 23120
rect 7412 23080 8140 23120
rect 8180 23080 9004 23120
rect 9044 23080 9196 23120
rect 9236 23080 9245 23120
rect 10723 23080 10732 23120
rect 10772 23080 15052 23120
rect 15092 23080 15101 23120
rect 17356 23080 19084 23120
rect 19124 23080 19133 23120
rect 2179 22996 2188 23036
rect 2228 22996 2380 23036
rect 2420 22996 2429 23036
rect 3043 23020 3052 23060
rect 3092 23020 3101 23060
rect 4685 22996 4780 23036
rect 4820 22996 4829 23036
rect 11779 22996 11788 23036
rect 11828 22996 12844 23036
rect 12884 22996 12893 23036
rect 13891 22996 13900 23036
rect 13940 22996 16724 23036
rect 16684 22952 16724 22996
rect 2371 22912 2380 22952
rect 2420 22912 2860 22952
rect 2900 22912 2909 22952
rect 7651 22912 7660 22952
rect 7700 22912 7852 22952
rect 7892 22912 7901 22952
rect 16675 22912 16684 22952
rect 16724 22912 16733 22952
rect 20899 22912 20908 22952
rect 20948 22912 21388 22952
rect 21428 22912 21437 22952
rect 5539 22828 5548 22868
rect 5588 22828 5740 22868
rect 5780 22828 5789 22868
rect 4919 22660 4928 22700
rect 4968 22660 5010 22700
rect 5050 22660 5092 22700
rect 5132 22660 5174 22700
rect 5214 22660 5256 22700
rect 5296 22660 5305 22700
rect 20039 22660 20048 22700
rect 20088 22660 20130 22700
rect 20170 22660 20212 22700
rect 20252 22660 20294 22700
rect 20334 22660 20376 22700
rect 20416 22660 20425 22700
rect 7075 22576 7084 22616
rect 7124 22576 8332 22616
rect 8372 22576 8381 22616
rect 14275 22576 14284 22616
rect 14324 22576 14476 22616
rect 14516 22576 14525 22616
rect 17741 22576 17836 22616
rect 17876 22576 17885 22616
rect 17443 22492 17452 22532
rect 17492 22492 17740 22532
rect 17780 22492 17789 22532
rect 1123 22408 1132 22448
rect 1172 22408 9964 22448
rect 10004 22408 10013 22448
rect 18413 22408 18508 22448
rect 18548 22408 18557 22448
rect 3427 22324 3436 22364
rect 3476 22324 4204 22364
rect 4244 22324 4253 22364
rect 11395 22324 11404 22364
rect 11444 22324 11500 22364
rect 11540 22324 11549 22364
rect 18691 22324 18700 22364
rect 18740 22324 18892 22364
rect 18932 22324 18941 22364
rect 3437 22240 3532 22280
rect 3572 22240 3581 22280
rect 6019 22240 6028 22280
rect 6068 22240 8428 22280
rect 8468 22240 8477 22280
rect 20419 22240 20428 22280
rect 20468 22240 21292 22280
rect 21332 22240 21341 22280
rect 2371 22156 2380 22196
rect 2420 22156 3916 22196
rect 3956 22156 3965 22196
rect 18787 22156 18796 22196
rect 18836 22156 19948 22196
rect 19988 22156 19997 22196
rect 3427 22072 3436 22112
rect 3476 22072 3724 22112
rect 3764 22072 3773 22112
rect 11491 22072 11500 22112
rect 11540 22072 20908 22112
rect 20948 22072 20957 22112
rect 3679 21904 3688 21944
rect 3728 21904 3770 21944
rect 3810 21904 3852 21944
rect 3892 21904 3934 21944
rect 3974 21904 4016 21944
rect 4056 21904 4065 21944
rect 11203 21904 11212 21944
rect 11252 21904 11404 21944
rect 11444 21904 11453 21944
rect 18799 21904 18808 21944
rect 18848 21904 18890 21944
rect 18930 21904 18972 21944
rect 19012 21904 19054 21944
rect 19094 21904 19136 21944
rect 19176 21904 19185 21944
rect 6787 21820 6796 21860
rect 6836 21820 8044 21860
rect 8084 21820 8093 21860
rect 3523 21736 3532 21776
rect 3572 21736 3820 21776
rect 3860 21736 3869 21776
rect 4291 21736 4300 21776
rect 4340 21736 4396 21776
rect 4436 21736 4445 21776
rect 14275 21736 14284 21776
rect 14324 21736 15244 21776
rect 15284 21736 15293 21776
rect 6787 21652 6796 21692
rect 6836 21652 6988 21692
rect 7028 21652 7037 21692
rect 13603 21652 13612 21692
rect 13652 21652 14572 21692
rect 14612 21652 14621 21692
rect 18403 21652 18412 21692
rect 18452 21652 19412 21692
rect 19372 21608 19412 21652
rect 451 21568 460 21608
rect 500 21568 1612 21608
rect 1652 21568 1661 21608
rect 4003 21568 4012 21608
rect 4052 21568 7180 21608
rect 7220 21568 7229 21608
rect 7363 21568 7372 21608
rect 7412 21568 7468 21608
rect 7508 21568 7517 21608
rect 10348 21568 11788 21608
rect 11828 21568 11837 21608
rect 15331 21568 15340 21608
rect 15380 21568 18508 21608
rect 18548 21568 18557 21608
rect 19363 21568 19372 21608
rect 19412 21568 19421 21608
rect 10348 21524 10388 21568
rect 4012 21484 10348 21524
rect 10388 21484 10397 21524
rect 10819 21484 10828 21524
rect 10868 21484 16012 21524
rect 16052 21484 16061 21524
rect 18019 21484 18028 21524
rect 18068 21484 18124 21524
rect 18164 21484 18173 21524
rect 18499 21484 18508 21524
rect 18548 21484 19180 21524
rect 19220 21484 19229 21524
rect 4012 21440 4052 21484
rect 1891 21400 1900 21440
rect 1940 21400 4052 21440
rect 4291 21400 4300 21440
rect 4340 21400 4588 21440
rect 4628 21400 4637 21440
rect 12355 21400 12364 21440
rect 12404 21400 13612 21440
rect 13652 21400 13661 21440
rect 15148 21400 21100 21440
rect 21140 21400 21149 21440
rect 15148 21356 15188 21400
rect 2371 21316 2380 21356
rect 2420 21316 15188 21356
rect 15235 21316 15244 21356
rect 15284 21316 15820 21356
rect 15860 21316 15869 21356
rect 10339 21232 10348 21272
rect 10388 21232 16492 21272
rect 16532 21232 16541 21272
rect 4919 21148 4928 21188
rect 4968 21148 5010 21188
rect 5050 21148 5092 21188
rect 5132 21148 5174 21188
rect 5214 21148 5256 21188
rect 5296 21148 5305 21188
rect 8803 21148 8812 21188
rect 8852 21148 8861 21188
rect 20039 21148 20048 21188
rect 20088 21148 20130 21188
rect 20170 21148 20212 21188
rect 20252 21148 20294 21188
rect 20334 21148 20376 21188
rect 20416 21148 20425 21188
rect 4771 20980 4780 21020
rect 4820 20980 6412 21020
rect 6452 20980 6461 21020
rect 8812 20936 8852 21148
rect 15811 21064 15820 21104
rect 15860 21064 18028 21104
rect 18068 21064 18508 21104
rect 18548 21064 18557 21104
rect 1795 20896 1804 20936
rect 1844 20896 5260 20936
rect 5300 20896 5309 20936
rect 8323 20896 8332 20936
rect 8372 20896 9196 20936
rect 9236 20896 9245 20936
rect 15331 20896 15340 20936
rect 15380 20896 16492 20936
rect 16532 20896 16541 20936
rect 2179 20812 2188 20852
rect 2228 20812 2380 20852
rect 2420 20812 2429 20852
rect 4195 20812 4204 20852
rect 4244 20812 5164 20852
rect 5204 20812 5213 20852
rect 5347 20812 5356 20852
rect 5396 20812 5740 20852
rect 5780 20812 5789 20852
rect 8525 20812 8620 20852
rect 8660 20812 8669 20852
rect 12739 20812 12748 20852
rect 12788 20812 16204 20852
rect 16244 20812 16253 20852
rect 3907 20728 3916 20768
rect 3956 20728 4588 20768
rect 4628 20728 4637 20768
rect 15331 20728 15340 20768
rect 15380 20728 20140 20768
rect 20180 20728 20189 20768
rect 451 20644 460 20684
rect 500 20644 3628 20684
rect 3668 20644 3677 20684
rect 5923 20644 5932 20684
rect 5972 20644 6124 20684
rect 6164 20644 6173 20684
rect 12931 20644 12940 20684
rect 12980 20644 16108 20684
rect 16148 20644 16157 20684
rect 2851 20560 2860 20600
rect 2900 20560 9100 20600
rect 9140 20560 9149 20600
rect 3679 20392 3688 20432
rect 3728 20392 3770 20432
rect 3810 20392 3852 20432
rect 3892 20392 3934 20432
rect 3974 20392 4016 20432
rect 4056 20392 4065 20432
rect 18799 20392 18808 20432
rect 18848 20392 18890 20432
rect 18930 20392 18972 20432
rect 19012 20392 19054 20432
rect 19094 20392 19136 20432
rect 19176 20392 19185 20432
rect 5155 20308 5164 20348
rect 5204 20308 11020 20348
rect 11060 20308 11212 20348
rect 11252 20308 11261 20348
rect 3523 20224 3532 20264
rect 3572 20224 4780 20264
rect 4820 20224 5548 20264
rect 5588 20224 5597 20264
rect 10723 20224 10732 20264
rect 10772 20224 11116 20264
rect 11156 20224 11165 20264
rect 11683 20224 11692 20264
rect 11732 20224 12076 20264
rect 12116 20224 12125 20264
rect 18499 20224 18508 20264
rect 18548 20224 19084 20264
rect 19124 20224 19133 20264
rect 7075 20140 7084 20180
rect 7124 20140 7133 20180
rect 7267 20140 7276 20180
rect 7316 20140 9964 20180
rect 10004 20140 10013 20180
rect 10915 20140 10924 20180
rect 10964 20140 13420 20180
rect 13460 20140 13469 20180
rect 14563 20140 14572 20180
rect 14612 20140 14764 20180
rect 14804 20140 14813 20180
rect 15235 20140 15244 20180
rect 15284 20140 15293 20180
rect 15725 20140 15820 20180
rect 15860 20140 15869 20180
rect 7084 20096 7124 20140
rect 15244 20096 15284 20140
rect 6787 20056 6796 20096
rect 6836 20056 7124 20096
rect 10915 20056 10924 20096
rect 10964 20056 13324 20096
rect 13364 20056 15340 20096
rect 15380 20056 15389 20096
rect 18595 20056 18604 20096
rect 18644 20056 19084 20096
rect 19124 20056 19133 20096
rect 20035 20056 20044 20096
rect 20084 20056 20093 20096
rect 20044 20012 20084 20056
rect 1987 19972 1996 20012
rect 2036 19972 7084 20012
rect 7124 19972 7133 20012
rect 13891 19972 13900 20012
rect 13940 19972 14092 20012
rect 14132 19972 14141 20012
rect 18883 19972 18892 20012
rect 18932 19972 20084 20012
rect 3427 19888 3436 19928
rect 3476 19888 3628 19928
rect 3668 19888 3677 19928
rect 7843 19888 7852 19928
rect 7892 19888 10348 19928
rect 10388 19888 10397 19928
rect 17731 19888 17740 19928
rect 17780 19888 17836 19928
rect 17876 19888 17885 19928
rect 20419 19888 20428 19928
rect 20468 19888 20716 19928
rect 20756 19888 20765 19928
rect 20035 19804 20044 19844
rect 20084 19804 20620 19844
rect 20660 19804 20669 19844
rect 5923 19720 5932 19760
rect 5972 19720 5981 19760
rect 14755 19720 14764 19760
rect 14804 19720 15340 19760
rect 15380 19720 15389 19760
rect 4919 19636 4928 19676
rect 4968 19636 5010 19676
rect 5050 19636 5092 19676
rect 5132 19636 5174 19676
rect 5214 19636 5256 19676
rect 5296 19636 5305 19676
rect 5347 19636 5356 19676
rect 5396 19636 5405 19676
rect 5356 19592 5396 19636
rect 5932 19592 5972 19720
rect 20039 19636 20048 19676
rect 20088 19636 20130 19676
rect 20170 19636 20212 19676
rect 20252 19636 20294 19676
rect 20334 19636 20376 19676
rect 20416 19636 20425 19676
rect 5164 19552 5396 19592
rect 5443 19552 5452 19592
rect 5492 19552 5972 19592
rect 5164 19508 5204 19552
rect 5155 19468 5164 19508
rect 5204 19468 5213 19508
rect 20131 19468 20140 19508
rect 20180 19468 21388 19508
rect 21428 19468 21437 19508
rect 259 19384 268 19424
rect 308 19384 748 19424
rect 788 19384 797 19424
rect 2851 19384 2860 19424
rect 2900 19384 3052 19424
rect 3092 19384 3101 19424
rect 4387 19384 4396 19424
rect 4436 19384 4780 19424
rect 4820 19384 4829 19424
rect 15043 19384 15052 19424
rect 15092 19384 15436 19424
rect 15476 19384 15485 19424
rect 3523 19300 3532 19340
rect 3572 19300 8332 19340
rect 8372 19300 8381 19340
rect 18499 19300 18508 19340
rect 18548 19300 18892 19340
rect 18932 19300 18941 19340
rect 3619 19216 3628 19256
rect 3668 19216 6124 19256
rect 6164 19216 9292 19256
rect 9332 19216 9341 19256
rect 19363 19216 19372 19256
rect 19412 19216 19852 19256
rect 19892 19216 19901 19256
rect 20515 19216 20524 19256
rect 20564 19216 20716 19256
rect 20756 19216 20765 19256
rect 14371 19048 14380 19088
rect 14420 19048 16492 19088
rect 16532 19048 18316 19088
rect 18356 19048 18365 19088
rect 3679 18880 3688 18920
rect 3728 18880 3770 18920
rect 3810 18880 3852 18920
rect 3892 18880 3934 18920
rect 3974 18880 4016 18920
rect 4056 18880 4065 18920
rect 4291 18880 4300 18920
rect 4340 18880 8428 18920
rect 8468 18880 8477 18920
rect 18799 18880 18808 18920
rect 18848 18880 18890 18920
rect 18930 18880 18972 18920
rect 19012 18880 19054 18920
rect 19094 18880 19136 18920
rect 19176 18880 19185 18920
rect 6115 18796 6124 18836
rect 6164 18796 7372 18836
rect 7412 18796 7421 18836
rect 2659 18628 2668 18668
rect 2708 18628 7276 18668
rect 7316 18628 7325 18668
rect 12835 18628 12844 18668
rect 12884 18628 16588 18668
rect 16628 18628 16637 18668
rect 3235 18544 3244 18584
rect 3284 18544 5068 18584
rect 5108 18544 5117 18584
rect 6499 18544 6508 18584
rect 6548 18544 6796 18584
rect 6836 18544 6845 18584
rect 7843 18544 7852 18584
rect 7892 18544 15724 18584
rect 15764 18544 15773 18584
rect 20131 18544 20140 18584
rect 20180 18544 20524 18584
rect 20564 18544 20573 18584
rect 8131 18460 8140 18500
rect 8180 18460 8524 18500
rect 8564 18460 8573 18500
rect 15245 18460 15340 18500
rect 15380 18460 15389 18500
rect 2179 18376 2188 18416
rect 2228 18376 3628 18416
rect 3668 18376 3677 18416
rect 4963 18376 4972 18416
rect 5012 18376 5452 18416
rect 5492 18376 5501 18416
rect 3149 18292 3244 18332
rect 3284 18292 4204 18332
rect 4244 18292 4253 18332
rect 19747 18208 19756 18248
rect 19796 18208 19805 18248
rect 4919 18124 4928 18164
rect 4968 18124 5010 18164
rect 5050 18124 5092 18164
rect 5132 18124 5174 18164
rect 5214 18124 5256 18164
rect 5296 18124 5305 18164
rect 17827 18124 17836 18164
rect 17876 18124 18220 18164
rect 18260 18124 18269 18164
rect 19756 17996 19796 18208
rect 20039 18124 20048 18164
rect 20088 18124 20130 18164
rect 20170 18124 20212 18164
rect 20252 18124 20294 18164
rect 20334 18124 20376 18164
rect 20416 18124 20425 18164
rect 2179 17956 2188 17996
rect 2228 17956 2668 17996
rect 2708 17956 2717 17996
rect 7747 17956 7756 17996
rect 7796 17956 8044 17996
rect 8084 17956 8093 17996
rect 12067 17956 12076 17996
rect 12116 17956 12556 17996
rect 12596 17956 12605 17996
rect 15331 17956 15340 17996
rect 15380 17956 15628 17996
rect 15668 17956 15677 17996
rect 18019 17956 18028 17996
rect 18068 17956 18220 17996
rect 18260 17956 18269 17996
rect 19651 17956 19660 17996
rect 19700 17956 19796 17996
rect 3139 17872 3148 17912
rect 3188 17872 5548 17912
rect 5588 17872 5597 17912
rect 17923 17872 17932 17912
rect 17972 17872 18604 17912
rect 18644 17872 18653 17912
rect 2947 17788 2956 17828
rect 2996 17788 3916 17828
rect 3956 17788 4300 17828
rect 4340 17788 4349 17828
rect 14851 17788 14860 17828
rect 14900 17788 15820 17828
rect 15860 17788 18028 17828
rect 18068 17788 18077 17828
rect 4003 17704 4012 17744
rect 4052 17704 6220 17744
rect 6260 17704 6269 17744
rect 14659 17704 14668 17744
rect 14708 17704 20140 17744
rect 20180 17704 20189 17744
rect 14563 17620 14572 17660
rect 14612 17620 15628 17660
rect 15668 17620 15677 17660
rect 15907 17620 15916 17660
rect 15956 17620 16492 17660
rect 16532 17620 16541 17660
rect 7171 17536 7180 17576
rect 7220 17536 21004 17576
rect 21044 17536 21053 17576
rect 2851 17452 2860 17492
rect 2900 17452 3340 17492
rect 3380 17452 3389 17492
rect 8323 17452 8332 17492
rect 8372 17452 8524 17492
rect 8564 17452 8573 17492
rect 13891 17452 13900 17492
rect 13940 17452 14188 17492
rect 14228 17452 14237 17492
rect 3679 17368 3688 17408
rect 3728 17368 3770 17408
rect 3810 17368 3852 17408
rect 3892 17368 3934 17408
rect 3974 17368 4016 17408
rect 4056 17368 4065 17408
rect 5731 17368 5740 17408
rect 5780 17368 8908 17408
rect 8948 17368 8957 17408
rect 18799 17368 18808 17408
rect 18848 17368 18890 17408
rect 18930 17368 18972 17408
rect 19012 17368 19054 17408
rect 19094 17368 19136 17408
rect 19176 17368 19185 17408
rect 11299 17200 11308 17240
rect 11348 17200 17260 17240
rect 17300 17200 17309 17240
rect 3427 17116 3436 17156
rect 3476 17116 3820 17156
rect 3860 17116 3869 17156
rect 5635 17116 5644 17156
rect 5684 17116 20140 17156
rect 20180 17116 20189 17156
rect 13507 17032 13516 17072
rect 13556 17032 20044 17072
rect 20084 17032 20093 17072
rect 4291 16948 4300 16988
rect 4340 16948 4780 16988
rect 4820 16948 6124 16988
rect 6164 16948 6173 16988
rect 7555 16948 7564 16988
rect 7604 16948 9868 16988
rect 9908 16948 9917 16988
rect 14371 16948 14380 16988
rect 14420 16948 14476 16988
rect 14516 16948 14668 16988
rect 14708 16948 14717 16988
rect 6124 16904 6164 16948
rect 4387 16864 4396 16904
rect 4436 16864 5068 16904
rect 5108 16864 5117 16904
rect 6124 16864 7852 16904
rect 7892 16864 7901 16904
rect 14659 16696 14668 16736
rect 14708 16696 14860 16736
rect 14900 16696 14909 16736
rect 4919 16612 4928 16652
rect 4968 16612 5010 16652
rect 5050 16612 5092 16652
rect 5132 16612 5174 16652
rect 5214 16612 5256 16652
rect 5296 16612 5305 16652
rect 20039 16612 20048 16652
rect 20088 16612 20130 16652
rect 20170 16612 20212 16652
rect 20252 16612 20294 16652
rect 20334 16612 20376 16652
rect 20416 16612 20425 16652
rect 13027 16528 13036 16568
rect 13076 16528 16876 16568
rect 16916 16528 16925 16568
rect 3331 16444 3340 16484
rect 3380 16444 3532 16484
rect 3572 16444 3581 16484
rect 6115 16444 6124 16484
rect 6164 16444 6508 16484
rect 6548 16444 6557 16484
rect 6979 16444 6988 16484
rect 7028 16444 7180 16484
rect 7220 16444 7229 16484
rect 15235 16444 15244 16484
rect 15284 16444 17836 16484
rect 17876 16444 17885 16484
rect 2371 16360 2380 16400
rect 2420 16360 9196 16400
rect 9236 16360 9245 16400
rect 4771 16276 4780 16316
rect 4820 16276 4972 16316
rect 5012 16276 5021 16316
rect 18499 16276 18508 16316
rect 18548 16276 18892 16316
rect 18932 16276 18941 16316
rect 6787 16192 6796 16232
rect 6836 16192 6988 16232
rect 7028 16192 7037 16232
rect 8611 16192 8620 16232
rect 8660 16192 11404 16232
rect 11444 16192 11453 16232
rect 2371 16108 2380 16148
rect 2420 16108 17260 16148
rect 17300 16108 17309 16148
rect 3679 15856 3688 15896
rect 3728 15856 3770 15896
rect 3810 15856 3852 15896
rect 3892 15856 3934 15896
rect 3974 15856 4016 15896
rect 4056 15856 4065 15896
rect 18799 15856 18808 15896
rect 18848 15856 18890 15896
rect 18930 15856 18972 15896
rect 19012 15856 19054 15896
rect 19094 15856 19136 15896
rect 19176 15856 19185 15896
rect 19747 15856 19756 15896
rect 19796 15856 19948 15896
rect 19988 15856 19997 15896
rect 6115 15772 6124 15812
rect 6164 15772 9580 15812
rect 9620 15772 9629 15812
rect 3619 15604 3628 15644
rect 3668 15604 6604 15644
rect 6644 15604 6796 15644
rect 6836 15604 6845 15644
rect 2956 15436 3148 15476
rect 3188 15436 3197 15476
rect 16483 15436 16492 15476
rect 16532 15436 18604 15476
rect 18644 15436 19372 15476
rect 19412 15436 19421 15476
rect 2956 15392 2996 15436
rect 2947 15352 2956 15392
rect 2996 15352 3005 15392
rect 13219 15352 13228 15392
rect 13268 15352 14956 15392
rect 14996 15352 15005 15392
rect 8611 15268 8620 15308
rect 8660 15268 20812 15308
rect 20852 15268 20861 15308
rect 4483 15184 4492 15224
rect 4532 15184 6700 15224
rect 6740 15184 6749 15224
rect 4919 15100 4928 15140
rect 4968 15100 5010 15140
rect 5050 15100 5092 15140
rect 5132 15100 5174 15140
rect 5214 15100 5256 15140
rect 5296 15100 5305 15140
rect 6211 15100 6220 15140
rect 6260 15100 6604 15140
rect 6644 15100 6653 15140
rect 20039 15100 20048 15140
rect 20088 15100 20130 15140
rect 20170 15100 20212 15140
rect 20252 15100 20294 15140
rect 20334 15100 20376 15140
rect 20416 15100 20425 15140
rect 2179 15016 2188 15056
rect 2228 15016 9100 15056
rect 9140 15016 9149 15056
rect 16003 14932 16012 14972
rect 16052 14932 18220 14972
rect 18260 14932 18269 14972
rect 8803 14848 8812 14888
rect 8852 14848 9580 14888
rect 9620 14848 9629 14888
rect 4387 14764 4396 14804
rect 4436 14764 4684 14804
rect 4724 14764 4733 14804
rect 14083 14764 14092 14804
rect 14132 14764 15148 14804
rect 15188 14764 15197 14804
rect 15427 14764 15436 14804
rect 15476 14764 15628 14804
rect 15668 14764 17260 14804
rect 17300 14764 17309 14804
rect 6979 14680 6988 14720
rect 7028 14680 7276 14720
rect 7316 14680 7325 14720
rect 13027 14680 13036 14720
rect 13076 14680 13171 14720
rect 8995 14596 9004 14636
rect 9044 14596 9484 14636
rect 9524 14596 9533 14636
rect 14467 14596 14476 14636
rect 14516 14596 14668 14636
rect 14708 14596 14717 14636
rect 12259 14512 12268 14552
rect 12308 14512 14284 14552
rect 14324 14512 14333 14552
rect 3679 14344 3688 14384
rect 3728 14344 3770 14384
rect 3810 14344 3852 14384
rect 3892 14344 3934 14384
rect 3974 14344 4016 14384
rect 4056 14344 4065 14384
rect 11011 14344 11020 14384
rect 11060 14344 11212 14384
rect 11252 14344 11261 14384
rect 18799 14344 18808 14384
rect 18848 14344 18890 14384
rect 18930 14344 18972 14384
rect 19012 14344 19054 14384
rect 19094 14344 19136 14384
rect 19176 14344 19185 14384
rect 1891 14260 1900 14300
rect 1940 14260 6700 14300
rect 6740 14260 6749 14300
rect 8227 14260 8236 14300
rect 8276 14260 12652 14300
rect 12692 14260 12701 14300
rect 16003 14176 16012 14216
rect 16052 14176 16204 14216
rect 16244 14176 16253 14216
rect 2659 14008 2668 14048
rect 2708 14008 2804 14048
rect 6211 14008 6220 14048
rect 6260 14008 8524 14048
rect 8564 14008 8812 14048
rect 8852 14008 8861 14048
rect 18499 14008 18508 14048
rect 18548 14008 19372 14048
rect 19412 14008 19421 14048
rect 1219 13840 1228 13880
rect 1268 13840 1420 13880
rect 1460 13840 1469 13880
rect 2764 13544 2804 14008
rect 2851 13924 2860 13964
rect 2900 13924 2995 13964
rect 3235 13924 3244 13964
rect 3284 13924 3628 13964
rect 3668 13924 3677 13964
rect 11309 13924 11404 13964
rect 11444 13924 11453 13964
rect 4387 13840 4396 13880
rect 4436 13840 5356 13880
rect 5396 13840 5405 13880
rect 5827 13840 5836 13880
rect 5876 13840 7372 13880
rect 7412 13840 7421 13880
rect 6595 13756 6604 13796
rect 6644 13756 7084 13796
rect 7124 13756 7133 13796
rect 13219 13756 13228 13796
rect 13268 13756 14668 13796
rect 14708 13756 14717 13796
rect 16387 13756 16396 13796
rect 16436 13756 16972 13796
rect 17012 13756 17021 13796
rect 4579 13672 4588 13712
rect 4628 13672 5548 13712
rect 5588 13672 5597 13712
rect 8899 13672 8908 13712
rect 8948 13672 19564 13712
rect 19604 13672 19613 13712
rect 4919 13588 4928 13628
rect 4968 13588 5010 13628
rect 5050 13588 5092 13628
rect 5132 13588 5174 13628
rect 5214 13588 5256 13628
rect 5296 13588 5305 13628
rect 20039 13588 20048 13628
rect 20088 13588 20130 13628
rect 20170 13588 20212 13628
rect 20252 13588 20294 13628
rect 20334 13588 20376 13628
rect 20416 13588 20425 13628
rect 2755 13504 2764 13544
rect 2804 13504 2813 13544
rect 3139 13504 3148 13544
rect 3188 13504 3244 13544
rect 3284 13504 3293 13544
rect 6883 13420 6892 13460
rect 6932 13420 7372 13460
rect 7412 13420 7421 13460
rect 11683 13420 11692 13460
rect 11732 13420 15436 13460
rect 15476 13420 15485 13460
rect 3148 13336 3340 13376
rect 3380 13336 3389 13376
rect 3148 13292 3188 13336
rect 2956 13252 3188 13292
rect 2956 13040 2996 13252
rect 3331 13168 3340 13208
rect 3380 13168 3532 13208
rect 3572 13168 3581 13208
rect 12931 13168 12940 13208
rect 12980 13168 13420 13208
rect 13460 13168 13469 13208
rect 16579 13168 16588 13208
rect 16628 13168 17012 13208
rect 13027 13084 13036 13124
rect 13076 13084 13132 13124
rect 13172 13084 13181 13124
rect 16972 13040 17012 13168
rect 2956 13000 3052 13040
rect 3092 13000 3101 13040
rect 4003 13000 4012 13040
rect 4052 13000 4204 13040
rect 4244 13000 4253 13040
rect 16963 13000 16972 13040
rect 17012 13000 17021 13040
rect 18211 13000 18220 13040
rect 18260 13000 18316 13040
rect 18356 13000 18365 13040
rect 1891 12940 1900 12980
rect 1940 12940 1949 12980
rect 1900 12872 1940 12940
rect 1411 12832 1420 12872
rect 1460 12832 1940 12872
rect 3331 12832 3340 12872
rect 3380 12832 3389 12872
rect 3679 12832 3688 12872
rect 3728 12832 3770 12872
rect 3810 12832 3852 12872
rect 3892 12832 3934 12872
rect 3974 12832 4016 12872
rect 4056 12832 4065 12872
rect 5923 12832 5932 12872
rect 5972 12832 7180 12872
rect 7220 12832 7229 12872
rect 18211 12832 18220 12872
rect 18260 12832 18316 12872
rect 18356 12832 18365 12872
rect 18799 12832 18808 12872
rect 18848 12832 18890 12872
rect 18930 12832 18972 12872
rect 19012 12832 19054 12872
rect 19094 12832 19136 12872
rect 19176 12832 19185 12872
rect 3340 12536 3380 12832
rect 13507 12748 13516 12788
rect 13556 12748 13708 12788
rect 13748 12748 13757 12788
rect 3907 12664 3916 12704
rect 3956 12664 4204 12704
rect 4244 12664 4253 12704
rect 4867 12664 4876 12704
rect 4916 12664 8908 12704
rect 8948 12664 8957 12704
rect 17261 12664 17356 12704
rect 17396 12664 17405 12704
rect 3523 12580 3532 12620
rect 3572 12580 3724 12620
rect 3764 12580 6604 12620
rect 6644 12580 6653 12620
rect 3331 12496 3340 12536
rect 3380 12496 3389 12536
rect 5827 12496 5836 12536
rect 5876 12496 9772 12536
rect 9812 12496 9821 12536
rect 2851 12412 2860 12452
rect 2900 12412 3244 12452
rect 3284 12412 3293 12452
rect 9571 12412 9580 12452
rect 9620 12412 10100 12452
rect 12067 12412 12076 12452
rect 12116 12412 12364 12452
rect 12404 12412 12413 12452
rect 12931 12412 12940 12452
rect 12980 12412 13900 12452
rect 13940 12412 13949 12452
rect 14371 12412 14380 12452
rect 14420 12412 18508 12452
rect 18548 12412 18557 12452
rect 3043 12328 3052 12368
rect 3092 12328 3244 12368
rect 3284 12328 3293 12368
rect 9580 12284 9620 12412
rect 10060 12368 10100 12412
rect 10060 12328 17452 12368
rect 17492 12328 17501 12368
rect 8803 12244 8812 12284
rect 8852 12244 9620 12284
rect 4919 12076 4928 12116
rect 4968 12076 5010 12116
rect 5050 12076 5092 12116
rect 5132 12076 5174 12116
rect 5214 12076 5256 12116
rect 5296 12076 5305 12116
rect 20039 12076 20048 12116
rect 20088 12076 20130 12116
rect 20170 12076 20212 12116
rect 20252 12076 20294 12116
rect 20334 12076 20376 12116
rect 20416 12076 20425 12116
rect 5251 11908 5260 11948
rect 5300 11908 5644 11948
rect 5684 11908 5693 11948
rect 4675 11824 4684 11864
rect 4724 11824 7564 11864
rect 7604 11824 7613 11864
rect 11875 11824 11884 11864
rect 11924 11824 19852 11864
rect 19892 11824 19901 11864
rect 13795 11740 13804 11780
rect 13844 11740 13900 11780
rect 13940 11740 13949 11780
rect 2371 11656 2380 11696
rect 2420 11656 3532 11696
rect 3572 11656 3581 11696
rect 9283 11656 9292 11696
rect 9332 11656 10348 11696
rect 10388 11656 10397 11696
rect 2851 11572 2860 11612
rect 2900 11572 4972 11612
rect 5012 11572 5021 11612
rect 14179 11488 14188 11528
rect 14228 11488 14476 11528
rect 14516 11488 14525 11528
rect 3679 11320 3688 11360
rect 3728 11320 3770 11360
rect 3810 11320 3852 11360
rect 3892 11320 3934 11360
rect 3974 11320 4016 11360
rect 4056 11320 4065 11360
rect 13987 11320 13996 11360
rect 14036 11320 15820 11360
rect 15860 11320 15869 11360
rect 18799 11320 18808 11360
rect 18848 11320 18890 11360
rect 18930 11320 18972 11360
rect 19012 11320 19054 11360
rect 19094 11320 19136 11360
rect 19176 11320 19185 11360
rect 3341 11152 3436 11192
rect 3476 11152 3485 11192
rect 3715 11152 3724 11192
rect 3764 11152 4300 11192
rect 4340 11152 4349 11192
rect 6595 11152 6604 11192
rect 6644 11152 6892 11192
rect 6932 11152 6941 11192
rect 10819 10984 10828 11024
rect 10868 10984 11404 11024
rect 11444 10984 11453 11024
rect 10819 10816 10828 10856
rect 10868 10816 11308 10856
rect 11348 10816 11357 10856
rect 4291 10732 4300 10772
rect 4340 10732 19756 10772
rect 19796 10732 19805 10772
rect 4919 10564 4928 10604
rect 4968 10564 5010 10604
rect 5050 10564 5092 10604
rect 5132 10564 5174 10604
rect 5214 10564 5256 10604
rect 5296 10564 5305 10604
rect 20039 10564 20048 10604
rect 20088 10564 20130 10604
rect 20170 10564 20212 10604
rect 20252 10564 20294 10604
rect 20334 10564 20376 10604
rect 20416 10564 20425 10604
rect 2083 10480 2092 10520
rect 2132 10480 2476 10520
rect 2516 10480 2525 10520
rect 2851 10480 2860 10520
rect 2900 10480 8524 10520
rect 8564 10480 8573 10520
rect 5155 10396 5164 10436
rect 5204 10396 5836 10436
rect 5876 10396 5885 10436
rect 2083 10312 2092 10352
rect 2132 10312 2284 10352
rect 2324 10312 2333 10352
rect 3619 10312 3628 10352
rect 3668 10312 6412 10352
rect 6452 10312 6461 10352
rect 3427 10228 3436 10268
rect 3476 10228 4684 10268
rect 4724 10228 4733 10268
rect 5923 10228 5932 10268
rect 5972 10228 6220 10268
rect 6260 10228 6269 10268
rect 17347 10228 17356 10268
rect 17396 10228 17836 10268
rect 17876 10228 17885 10268
rect 2275 10144 2284 10184
rect 2324 10144 19276 10184
rect 19316 10144 19325 10184
rect 2093 10060 2188 10100
rect 2228 10060 2237 10100
rect 3396 10060 3436 10100
rect 3476 10060 3485 10100
rect 11309 10060 11404 10100
rect 11444 10060 11453 10100
rect 14477 10060 14572 10100
rect 14612 10060 14621 10100
rect 3436 10016 3476 10060
rect 2947 9976 2956 10016
rect 2996 9976 3476 10016
rect 3715 9976 3724 10016
rect 3764 9976 7948 10016
rect 7988 9976 7997 10016
rect 3679 9808 3688 9848
rect 3728 9808 3770 9848
rect 3810 9808 3852 9848
rect 3892 9808 3934 9848
rect 3974 9808 4016 9848
rect 4056 9808 4065 9848
rect 18799 9808 18808 9848
rect 18848 9808 18890 9848
rect 18930 9808 18972 9848
rect 19012 9808 19054 9848
rect 19094 9808 19136 9848
rect 19176 9808 19185 9848
rect 15619 9724 15628 9764
rect 15668 9724 20044 9764
rect 20084 9724 20093 9764
rect 1699 9640 1708 9680
rect 1748 9640 5836 9680
rect 5876 9640 5885 9680
rect 15331 9640 15340 9680
rect 15380 9640 19564 9680
rect 19604 9640 19613 9680
rect 13315 9556 13324 9596
rect 13364 9556 13516 9596
rect 13556 9556 13565 9596
rect 13891 9556 13900 9596
rect 13940 9556 14284 9596
rect 14324 9556 14333 9596
rect 3427 9472 3436 9512
rect 3476 9472 4012 9512
rect 4052 9472 4061 9512
rect 10051 9388 10060 9428
rect 10100 9388 10109 9428
rect 10060 9344 10100 9388
rect 9859 9304 9868 9344
rect 9908 9304 10100 9344
rect 10627 9304 10636 9344
rect 10676 9304 14380 9344
rect 14420 9304 14429 9344
rect 10147 9220 10156 9260
rect 10196 9220 15628 9260
rect 15668 9220 15677 9260
rect 4919 9052 4928 9092
rect 4968 9052 5010 9092
rect 5050 9052 5092 9092
rect 5132 9052 5174 9092
rect 5214 9052 5256 9092
rect 5296 9052 5305 9092
rect 13891 9052 13900 9092
rect 13940 9052 13949 9092
rect 20039 9052 20048 9092
rect 20088 9052 20130 9092
rect 20170 9052 20212 9092
rect 20252 9052 20294 9092
rect 20334 9052 20376 9092
rect 20416 9052 20425 9092
rect 3907 8968 3916 9008
rect 3956 8968 5356 9008
rect 5396 8968 5405 9008
rect 5059 8884 5068 8924
rect 5108 8884 10060 8924
rect 10100 8884 10109 8924
rect 5347 8800 5356 8840
rect 5396 8800 6700 8840
rect 6740 8800 6749 8840
rect 13900 8756 13940 9052
rect 13699 8716 13708 8756
rect 13748 8716 13940 8756
rect 15907 8716 15916 8756
rect 15956 8716 16492 8756
rect 16532 8716 16541 8756
rect 3811 8632 3820 8672
rect 3860 8632 21292 8672
rect 21332 8632 21341 8672
rect 1795 8548 1804 8588
rect 1844 8548 3916 8588
rect 3956 8548 3965 8588
rect 13507 8548 13516 8588
rect 13556 8548 14188 8588
rect 14228 8548 14237 8588
rect 2467 8464 2476 8504
rect 2516 8464 2956 8504
rect 2996 8464 3005 8504
rect 3679 8296 3688 8336
rect 3728 8296 3770 8336
rect 3810 8296 3852 8336
rect 3892 8296 3934 8336
rect 3974 8296 4016 8336
rect 4056 8296 4065 8336
rect 18799 8296 18808 8336
rect 18848 8296 18890 8336
rect 18930 8296 18972 8336
rect 19012 8296 19054 8336
rect 19094 8296 19136 8336
rect 19176 8296 19185 8336
rect 4291 8128 4300 8168
rect 4340 8128 4588 8168
rect 4628 8128 4637 8168
rect 16205 8128 16300 8168
rect 16340 8128 16349 8168
rect 3427 7960 3436 8000
rect 3476 7960 11020 8000
rect 11060 7960 11069 8000
rect 9091 7876 9100 7916
rect 9140 7876 9964 7916
rect 10004 7876 10013 7916
rect 13027 7792 13036 7832
rect 13076 7792 13708 7832
rect 13748 7792 13757 7832
rect 4919 7540 4928 7580
rect 4968 7540 5010 7580
rect 5050 7540 5092 7580
rect 5132 7540 5174 7580
rect 5214 7540 5256 7580
rect 5296 7540 5305 7580
rect 20039 7540 20048 7580
rect 20088 7540 20130 7580
rect 20170 7540 20212 7580
rect 20252 7540 20294 7580
rect 20334 7540 20376 7580
rect 20416 7540 20425 7580
rect 6211 7120 6220 7160
rect 6260 7120 8812 7160
rect 8852 7120 8861 7160
rect 16771 7120 16780 7160
rect 16820 7120 18124 7160
rect 18164 7120 18173 7160
rect 2851 6868 2860 6908
rect 2900 6868 6124 6908
rect 6164 6868 6173 6908
rect 3679 6784 3688 6824
rect 3728 6784 3770 6824
rect 3810 6784 3852 6824
rect 3892 6784 3934 6824
rect 3974 6784 4016 6824
rect 4056 6784 4065 6824
rect 18799 6784 18808 6824
rect 18848 6784 18890 6824
rect 18930 6784 18972 6824
rect 19012 6784 19054 6824
rect 19094 6784 19136 6824
rect 19176 6784 19185 6824
rect 2851 6280 2860 6320
rect 2900 6280 19660 6320
rect 19700 6280 19709 6320
rect 1603 6112 1612 6152
rect 1652 6112 10060 6152
rect 10100 6112 10109 6152
rect 4919 6028 4928 6068
rect 4968 6028 5010 6068
rect 5050 6028 5092 6068
rect 5132 6028 5174 6068
rect 5214 6028 5256 6068
rect 5296 6028 5305 6068
rect 9667 6028 9676 6068
rect 9716 6028 12556 6068
rect 12596 6028 12605 6068
rect 20039 6028 20048 6068
rect 20088 6028 20130 6068
rect 20170 6028 20212 6068
rect 20252 6028 20294 6068
rect 20334 6028 20376 6068
rect 20416 6028 20425 6068
rect 5827 5944 5836 5984
rect 5876 5944 10156 5984
rect 10196 5944 10205 5984
rect 4099 5692 4108 5732
rect 4148 5692 7372 5732
rect 7412 5692 7421 5732
rect 13987 5692 13996 5732
rect 14036 5692 14045 5732
rect 14275 5692 14284 5732
rect 14324 5692 15052 5732
rect 15092 5692 15101 5732
rect 13996 5648 14036 5692
rect 4675 5608 4684 5648
rect 4724 5608 4876 5648
rect 4916 5608 4925 5648
rect 13996 5608 14668 5648
rect 14708 5608 14717 5648
rect 3139 5524 3148 5564
rect 3188 5524 5548 5564
rect 5588 5524 5597 5564
rect 9475 5524 9484 5564
rect 9524 5524 13996 5564
rect 14036 5524 14045 5564
rect 4771 5440 4780 5480
rect 4820 5440 20716 5480
rect 20756 5440 20765 5480
rect 3679 5272 3688 5312
rect 3728 5272 3770 5312
rect 3810 5272 3852 5312
rect 3892 5272 3934 5312
rect 3974 5272 4016 5312
rect 4056 5272 4065 5312
rect 18799 5272 18808 5312
rect 18848 5272 18890 5312
rect 18930 5272 18972 5312
rect 19012 5272 19054 5312
rect 19094 5272 19136 5312
rect 19176 5272 19185 5312
rect 10051 5188 10060 5228
rect 10100 5188 12556 5228
rect 12596 5188 12605 5228
rect 14179 4852 14188 4892
rect 14228 4852 16396 4892
rect 16436 4852 16445 4892
rect 4919 4516 4928 4556
rect 4968 4516 5010 4556
rect 5050 4516 5092 4556
rect 5132 4516 5174 4556
rect 5214 4516 5256 4556
rect 5296 4516 5305 4556
rect 20039 4516 20048 4556
rect 20088 4516 20130 4556
rect 20170 4516 20212 4556
rect 20252 4516 20294 4556
rect 20334 4516 20376 4556
rect 20416 4516 20425 4556
rect 5347 4264 5356 4304
rect 5396 4264 8716 4304
rect 8756 4264 8765 4304
rect 10915 4180 10924 4220
rect 10964 4180 17452 4220
rect 17492 4180 17501 4220
rect 14467 4096 14476 4136
rect 14516 4096 17356 4136
rect 17396 4096 17405 4136
rect 3679 3760 3688 3800
rect 3728 3760 3770 3800
rect 3810 3760 3852 3800
rect 3892 3760 3934 3800
rect 3974 3760 4016 3800
rect 4056 3760 4065 3800
rect 4675 3760 4684 3800
rect 4724 3760 12652 3800
rect 12692 3760 12701 3800
rect 18799 3760 18808 3800
rect 18848 3760 18890 3800
rect 18930 3760 18972 3800
rect 19012 3760 19054 3800
rect 19094 3760 19136 3800
rect 19176 3760 19185 3800
rect 5539 3508 5548 3548
rect 5588 3508 10252 3548
rect 10292 3508 10301 3548
rect 1987 3424 1996 3464
rect 2036 3424 2380 3464
rect 2420 3424 2429 3464
rect 13027 3424 13036 3464
rect 13076 3424 17644 3464
rect 17684 3424 17693 3464
rect 7747 3340 7756 3380
rect 7796 3340 12076 3380
rect 12116 3340 12125 3380
rect 9955 3172 9964 3212
rect 10004 3172 18700 3212
rect 18740 3172 18749 3212
rect 6691 3088 6700 3128
rect 6740 3088 9868 3128
rect 9908 3088 9917 3128
rect 4919 3004 4928 3044
rect 4968 3004 5010 3044
rect 5050 3004 5092 3044
rect 5132 3004 5174 3044
rect 5214 3004 5256 3044
rect 5296 3004 5305 3044
rect 20039 3004 20048 3044
rect 20088 3004 20130 3044
rect 20170 3004 20212 3044
rect 20252 3004 20294 3044
rect 20334 3004 20376 3044
rect 20416 3004 20425 3044
rect 1411 2920 1420 2960
rect 1460 2920 10060 2960
rect 10100 2920 10109 2960
rect 4579 2836 4588 2876
rect 4628 2836 4876 2876
rect 4916 2836 4925 2876
rect 8333 2836 8428 2876
rect 8468 2836 8477 2876
rect 13987 2836 13996 2876
rect 14036 2836 15148 2876
rect 15188 2836 15197 2876
rect 3523 2752 3532 2792
rect 3572 2752 4492 2792
rect 4532 2752 4541 2792
rect 13603 2752 13612 2792
rect 13652 2752 17740 2792
rect 17780 2752 17789 2792
rect 9187 2668 9196 2708
rect 9236 2668 10828 2708
rect 10868 2668 10877 2708
rect 1997 2584 2092 2624
rect 2132 2584 2141 2624
rect 2669 2584 2764 2624
rect 2804 2584 2813 2624
rect 10253 2584 10348 2624
rect 10388 2584 10397 2624
rect 14669 2584 14764 2624
rect 14804 2584 14813 2624
rect 8035 2416 8044 2456
rect 8084 2416 9772 2456
rect 9812 2416 9821 2456
rect 12259 2416 12268 2456
rect 12308 2416 13612 2456
rect 13652 2416 13661 2456
rect 2467 2332 2476 2372
rect 2516 2332 6028 2372
rect 6068 2332 6077 2372
rect 9379 2332 9388 2372
rect 9428 2332 12460 2372
rect 12500 2332 12509 2372
rect 3679 2248 3688 2288
rect 3728 2248 3770 2288
rect 3810 2248 3852 2288
rect 3892 2248 3934 2288
rect 3974 2248 4016 2288
rect 4056 2248 4065 2288
rect 18799 2248 18808 2288
rect 18848 2248 18890 2288
rect 18930 2248 18972 2288
rect 19012 2248 19054 2288
rect 19094 2248 19136 2288
rect 19176 2248 19185 2288
rect 2947 2164 2956 2204
rect 2996 2164 4204 2204
rect 4244 2164 4253 2204
rect 2189 2080 2284 2120
rect 2324 2080 2333 2120
rect 2477 2080 2572 2120
rect 2612 2080 2621 2120
rect 3245 2080 3340 2120
rect 3380 2080 3389 2120
rect 5827 2080 5836 2120
rect 5876 2080 6892 2120
rect 6932 2080 6941 2120
rect 7075 1996 7084 2036
rect 7124 1996 10732 2036
rect 10772 1996 10781 2036
rect 11299 1996 11308 2036
rect 11348 1996 12652 2036
rect 12692 1996 12701 2036
rect 8995 1912 9004 1952
rect 9044 1912 9292 1952
rect 9332 1912 9341 1952
rect 11405 1912 11500 1952
rect 11540 1912 11549 1952
rect 13325 1912 13420 1952
rect 13460 1912 13469 1952
rect 15331 1912 15340 1952
rect 15380 1912 18220 1952
rect 18260 1912 18269 1952
rect 2467 1744 2476 1784
rect 2516 1744 6508 1784
rect 6548 1744 6557 1784
rect 4919 1492 4928 1532
rect 4968 1492 5010 1532
rect 5050 1492 5092 1532
rect 5132 1492 5174 1532
rect 5214 1492 5256 1532
rect 5296 1492 5305 1532
rect 20039 1492 20048 1532
rect 20088 1492 20130 1532
rect 20170 1492 20212 1532
rect 20252 1492 20294 1532
rect 20334 1492 20376 1532
rect 20416 1492 20425 1532
rect 7661 1408 7756 1448
rect 7796 1408 7805 1448
rect 8045 1408 8140 1448
rect 8180 1408 8189 1448
rect 8237 1408 8332 1448
rect 8372 1408 8381 1448
rect 8429 1408 8524 1448
rect 8564 1408 8573 1448
rect 13123 1408 13132 1448
rect 13172 1408 16396 1448
rect 16436 1408 16445 1448
rect 17155 1408 17164 1448
rect 17204 1408 19276 1448
rect 19316 1408 19325 1448
rect 19373 1408 19468 1448
rect 19508 1408 19517 1448
rect 13699 1324 13708 1364
rect 13748 1324 16780 1364
rect 16820 1324 16829 1364
rect 8803 1240 8812 1280
rect 8852 1240 16012 1280
rect 16052 1240 16061 1280
rect 16387 1240 16396 1280
rect 16436 1240 18508 1280
rect 18548 1240 18557 1280
rect 6595 1156 6604 1196
rect 6644 1156 7180 1196
rect 7220 1156 7229 1196
rect 9667 1156 9676 1196
rect 9716 1156 15820 1196
rect 15860 1156 15869 1196
rect 18691 1156 18700 1196
rect 18740 1156 21484 1196
rect 21524 1156 21533 1196
rect 5251 988 5260 1028
rect 5300 988 5548 1028
rect 5588 988 5597 1028
rect 16963 988 16972 1028
rect 17012 988 17932 1028
rect 17972 988 17981 1028
rect 14179 820 14188 860
rect 14228 820 17164 860
rect 17204 820 17213 860
rect 15619 568 15628 608
rect 15668 568 19852 608
rect 19892 568 19901 608
rect 16195 484 16204 524
rect 16244 484 18316 524
rect 18356 484 18365 524
rect 13315 400 13324 440
rect 13364 400 16588 440
rect 16628 400 16637 440
rect 6883 316 6892 356
rect 6932 316 7564 356
rect 7604 316 7613 356
rect 9763 316 9772 356
rect 9812 316 17548 356
rect 17588 316 17597 356
rect 6403 232 6412 272
rect 6452 232 16204 272
rect 16244 232 16253 272
rect 2659 148 2668 188
rect 2708 148 16972 188
rect 17012 148 17021 188
rect 19075 148 19084 188
rect 19124 148 19372 188
rect 19412 148 19421 188
<< via4 >>
rect 9100 96580 9140 96620
rect 12556 95908 12596 95948
rect 9484 95656 9524 95696
rect 4928 95236 4968 95276
rect 5010 95236 5050 95276
rect 5092 95236 5132 95276
rect 5174 95236 5214 95276
rect 5256 95236 5296 95276
rect 20048 95236 20088 95276
rect 20130 95236 20170 95276
rect 20212 95236 20252 95276
rect 20294 95236 20334 95276
rect 20376 95236 20416 95276
rect 10636 94900 10676 94940
rect 1324 94816 1364 94856
rect 1804 94816 1844 94856
rect 2092 94816 2132 94856
rect 2476 94816 2516 94856
rect 3340 94816 3380 94856
rect 4396 94816 4436 94856
rect 4684 94816 4724 94856
rect 6316 94816 6356 94856
rect 6700 94816 6740 94856
rect 7084 94816 7124 94856
rect 18220 94816 18260 94856
rect 10732 94732 10772 94772
rect 12364 94732 12404 94772
rect 13420 94732 13460 94772
rect 14380 94732 14420 94772
rect 8812 94648 8852 94688
rect 9388 94648 9428 94688
rect 9772 94648 9812 94688
rect 10540 94648 10580 94688
rect 11212 94648 11252 94688
rect 11596 94648 11636 94688
rect 12172 94648 12212 94688
rect 3688 94480 3728 94520
rect 3770 94480 3810 94520
rect 3852 94480 3892 94520
rect 3934 94480 3974 94520
rect 4016 94480 4056 94520
rect 18808 94480 18848 94520
rect 18890 94480 18930 94520
rect 18972 94480 19012 94520
rect 19054 94480 19094 94520
rect 19136 94480 19176 94520
rect 4492 94144 4532 94184
rect 5548 94144 5588 94184
rect 5740 94144 5780 94184
rect 6124 94144 6164 94184
rect 8044 94144 8084 94184
rect 12748 94144 12788 94184
rect 16204 94144 16244 94184
rect 16972 94144 17012 94184
rect 18028 94144 18068 94184
rect 19372 94144 19412 94184
rect 21484 94144 21524 94184
rect 12460 94060 12500 94100
rect 9964 93976 10004 94016
rect 11020 93976 11060 94016
rect 5932 93892 5972 93932
rect 7756 93892 7796 93932
rect 10156 93892 10196 93932
rect 10828 93892 10868 93932
rect 11116 93892 11156 93932
rect 13900 93892 13940 93932
rect 14284 93892 14324 93932
rect 14668 93892 14708 93932
rect 15148 93892 15188 93932
rect 16588 93892 16628 93932
rect 17740 93892 17780 93932
rect 6892 93808 6932 93848
rect 4928 93724 4968 93764
rect 5010 93724 5050 93764
rect 5092 93724 5132 93764
rect 5174 93724 5214 93764
rect 5256 93724 5296 93764
rect 11884 93724 11924 93764
rect 20048 93724 20088 93764
rect 20130 93724 20170 93764
rect 20212 93724 20252 93764
rect 20294 93724 20334 93764
rect 20376 93724 20416 93764
rect 16780 93640 16820 93680
rect 7180 93556 7220 93596
rect 17164 93304 17204 93344
rect 19852 93304 19892 93344
rect 21388 93304 21428 93344
rect 18124 93136 18164 93176
rect 3688 92968 3728 93008
rect 3770 92968 3810 93008
rect 3852 92968 3892 93008
rect 3934 92968 3974 93008
rect 4016 92968 4056 93008
rect 18808 92968 18848 93008
rect 18890 92968 18930 93008
rect 18972 92968 19012 93008
rect 19054 92968 19094 93008
rect 19136 92968 19176 93008
rect 9292 92632 9332 92672
rect 19468 92632 19508 92672
rect 19660 92632 19700 92672
rect 6604 92296 6644 92336
rect 4928 92212 4968 92252
rect 5010 92212 5050 92252
rect 5092 92212 5132 92252
rect 5174 92212 5214 92252
rect 5256 92212 5296 92252
rect 20048 92212 20088 92252
rect 20130 92212 20170 92252
rect 20212 92212 20252 92252
rect 20294 92212 20334 92252
rect 20376 92212 20416 92252
rect 8332 91792 8372 91832
rect 19564 91792 19604 91832
rect 3688 91456 3728 91496
rect 3770 91456 3810 91496
rect 3852 91456 3892 91496
rect 3934 91456 3974 91496
rect 4016 91456 4056 91496
rect 18808 91456 18848 91496
rect 18890 91456 18930 91496
rect 18972 91456 19012 91496
rect 19054 91456 19094 91496
rect 19136 91456 19176 91496
rect 8140 91120 8180 91160
rect 8524 91120 8564 91160
rect 20908 91120 20948 91160
rect 3052 90868 3092 90908
rect 4928 90700 4968 90740
rect 5010 90700 5050 90740
rect 5092 90700 5132 90740
rect 5174 90700 5214 90740
rect 5256 90700 5296 90740
rect 14476 90700 14516 90740
rect 20048 90700 20088 90740
rect 20130 90700 20170 90740
rect 20212 90700 20252 90740
rect 20294 90700 20334 90740
rect 20376 90700 20416 90740
rect 2380 90280 2420 90320
rect 21292 90280 21332 90320
rect 4204 90112 4244 90152
rect 3532 89944 3572 89984
rect 3688 89944 3728 89984
rect 3770 89944 3810 89984
rect 3852 89944 3892 89984
rect 3934 89944 3974 89984
rect 4016 89944 4056 89984
rect 18808 89944 18848 89984
rect 18890 89944 18930 89984
rect 18972 89944 19012 89984
rect 19054 89944 19094 89984
rect 19136 89944 19176 89984
rect 10924 89860 10964 89900
rect 1708 89776 1748 89816
rect 1420 89608 1460 89648
rect 4588 89608 4628 89648
rect 16492 89608 16532 89648
rect 20812 89608 20852 89648
rect 13804 89440 13844 89480
rect 1996 89356 2036 89396
rect 3148 89356 3188 89396
rect 14860 89356 14900 89396
rect 4928 89188 4968 89228
rect 5010 89188 5050 89228
rect 5092 89188 5132 89228
rect 5174 89188 5214 89228
rect 5256 89188 5296 89228
rect 20048 89188 20088 89228
rect 20130 89188 20170 89228
rect 20212 89188 20252 89228
rect 20294 89188 20334 89228
rect 20376 89188 20416 89228
rect 2860 89020 2900 89060
rect 14188 89020 14228 89060
rect 16396 89020 16436 89060
rect 12268 88852 12308 88892
rect 18604 88768 18644 88808
rect 7660 88684 7700 88724
rect 20524 88600 20564 88640
rect 3688 88432 3728 88472
rect 3770 88432 3810 88472
rect 3852 88432 3892 88472
rect 3934 88432 3974 88472
rect 4016 88432 4056 88472
rect 18808 88432 18848 88472
rect 18890 88432 18930 88472
rect 18972 88432 19012 88472
rect 19054 88432 19094 88472
rect 19136 88432 19176 88472
rect 17356 88096 17396 88136
rect 9676 88012 9716 88052
rect 8236 87928 8276 87968
rect 13132 87928 13172 87968
rect 13708 87928 13748 87968
rect 15340 87844 15380 87884
rect 15532 87844 15572 87884
rect 4928 87676 4968 87716
rect 5010 87676 5050 87716
rect 5092 87676 5132 87716
rect 5174 87676 5214 87716
rect 5256 87676 5296 87716
rect 20048 87676 20088 87716
rect 20130 87676 20170 87716
rect 20212 87676 20252 87716
rect 20294 87676 20334 87716
rect 20376 87676 20416 87716
rect 8716 87508 8756 87548
rect 17644 87424 17684 87464
rect 21196 87424 21236 87464
rect 3532 87256 3572 87296
rect 19756 87256 19796 87296
rect 21100 87256 21140 87296
rect 5452 87088 5492 87128
rect 3688 86920 3728 86960
rect 3770 86920 3810 86960
rect 3852 86920 3892 86960
rect 3934 86920 3974 86960
rect 4016 86920 4056 86960
rect 18808 86920 18848 86960
rect 18890 86920 18930 86960
rect 18972 86920 19012 86960
rect 19054 86920 19094 86960
rect 19136 86920 19176 86960
rect 20716 86584 20756 86624
rect 7948 86500 7988 86540
rect 17932 86500 17972 86540
rect 13036 86416 13076 86456
rect 16684 86416 16724 86456
rect 2668 86332 2708 86372
rect 10252 86332 10292 86372
rect 4928 86164 4968 86204
rect 5010 86164 5050 86204
rect 5092 86164 5132 86204
rect 5174 86164 5214 86204
rect 5256 86164 5296 86204
rect 20048 86164 20088 86204
rect 20130 86164 20170 86204
rect 20212 86164 20252 86204
rect 20294 86164 20334 86204
rect 20376 86164 20416 86204
rect 17260 85912 17300 85952
rect 13996 85828 14036 85868
rect 17836 85744 17876 85784
rect 10444 85576 10484 85616
rect 1516 85492 1556 85532
rect 3688 85408 3728 85448
rect 3770 85408 3810 85448
rect 3852 85408 3892 85448
rect 3934 85408 3974 85448
rect 4016 85408 4056 85448
rect 18808 85408 18848 85448
rect 18890 85408 18930 85448
rect 18972 85408 19012 85448
rect 19054 85408 19094 85448
rect 19136 85408 19176 85448
rect 21196 85408 21236 85448
rect 14092 85156 14132 85196
rect 3244 85072 3284 85112
rect 4780 85072 4820 85112
rect 5452 85072 5492 85112
rect 7852 85072 7892 85112
rect 13132 84988 13172 85028
rect 13996 84988 14036 85028
rect 16876 84820 16916 84860
rect 8428 84736 8468 84776
rect 4928 84652 4968 84692
rect 5010 84652 5050 84692
rect 5092 84652 5132 84692
rect 5174 84652 5214 84692
rect 5256 84652 5296 84692
rect 20048 84652 20088 84692
rect 20130 84652 20170 84692
rect 20212 84652 20252 84692
rect 20294 84652 20334 84692
rect 20376 84652 20416 84692
rect 20524 84568 20564 84608
rect 5548 84484 5588 84524
rect 5836 84484 5876 84524
rect 3436 84316 3476 84356
rect 2764 84232 2804 84272
rect 21004 84232 21044 84272
rect 14476 84148 14516 84188
rect 19276 84148 19316 84188
rect 1612 84064 1652 84104
rect 1900 84064 1940 84104
rect 13804 84064 13844 84104
rect 2860 83980 2900 84020
rect 3688 83896 3728 83936
rect 3770 83896 3810 83936
rect 3852 83896 3892 83936
rect 3934 83896 3974 83936
rect 4016 83896 4056 83936
rect 2380 83644 2420 83684
rect 17260 83812 17300 83852
rect 14092 83728 14132 83768
rect 3244 83560 3284 83600
rect 1516 83392 1556 83432
rect 2764 83392 2804 83432
rect 5452 83476 5492 83516
rect 9004 83392 9044 83432
rect 18808 83896 18848 83936
rect 18890 83896 18930 83936
rect 18972 83896 19012 83936
rect 19054 83896 19094 83936
rect 19136 83896 19176 83936
rect 14764 83560 14804 83600
rect 17452 83560 17492 83600
rect 18412 83560 18452 83600
rect 21292 83560 21332 83600
rect 17452 83392 17492 83432
rect 18316 83392 18356 83432
rect 5836 83224 5876 83264
rect 7948 83224 7988 83264
rect 4928 83140 4968 83180
rect 5010 83140 5050 83180
rect 5092 83140 5132 83180
rect 5174 83140 5214 83180
rect 5256 83140 5296 83180
rect 3436 83056 3476 83096
rect 20048 83140 20088 83180
rect 20130 83140 20170 83180
rect 20212 83140 20252 83180
rect 20294 83140 20334 83180
rect 20376 83140 20416 83180
rect 4300 82972 4340 83012
rect 4780 82972 4820 83012
rect 11980 82972 12020 83012
rect 4780 82804 4820 82844
rect 10444 82804 10484 82844
rect 3532 82720 3572 82760
rect 14092 82720 14132 82760
rect 16108 82636 16148 82676
rect 3532 82552 3572 82592
rect 3688 82384 3728 82424
rect 3770 82384 3810 82424
rect 3852 82384 3892 82424
rect 3934 82384 3974 82424
rect 4016 82384 4056 82424
rect 18808 82384 18848 82424
rect 18890 82384 18930 82424
rect 18972 82384 19012 82424
rect 19054 82384 19094 82424
rect 19136 82384 19176 82424
rect 1324 82300 1364 82340
rect 5836 82216 5876 82256
rect 1420 82048 1460 82088
rect 3532 81964 3572 82004
rect 13612 82132 13652 82172
rect 13804 82048 13844 82088
rect 7468 81796 7508 81836
rect 17932 81796 17972 81836
rect 4928 81628 4968 81668
rect 5010 81628 5050 81668
rect 5092 81628 5132 81668
rect 5174 81628 5214 81668
rect 5256 81628 5296 81668
rect 16108 81544 16148 81584
rect 5548 81460 5588 81500
rect 6028 81460 6068 81500
rect 18508 81460 18548 81500
rect 20048 81628 20088 81668
rect 20130 81628 20170 81668
rect 20212 81628 20252 81668
rect 20294 81628 20334 81668
rect 20376 81628 20416 81668
rect 3148 81376 3188 81416
rect 5836 81124 5876 81164
rect 6412 81040 6452 81080
rect 3688 80872 3728 80912
rect 3770 80872 3810 80912
rect 3852 80872 3892 80912
rect 3934 80872 3974 80912
rect 4016 80872 4056 80912
rect 18808 80872 18848 80912
rect 18890 80872 18930 80912
rect 18972 80872 19012 80912
rect 19054 80872 19094 80912
rect 19136 80872 19176 80912
rect 18316 80704 18356 80744
rect 1516 80536 1556 80576
rect 12076 80620 12116 80660
rect 2572 80536 2612 80576
rect 17452 80536 17492 80576
rect 7372 80368 7412 80408
rect 5548 80284 5588 80324
rect 4928 80116 4968 80156
rect 5010 80116 5050 80156
rect 5092 80116 5132 80156
rect 5174 80116 5214 80156
rect 5256 80116 5296 80156
rect 20048 80116 20088 80156
rect 20130 80116 20170 80156
rect 20212 80116 20252 80156
rect 20294 80116 20334 80156
rect 20376 80116 20416 80156
rect 12460 80032 12500 80072
rect 1708 79864 1748 79904
rect 12652 79948 12692 79988
rect 7948 79864 7988 79904
rect 13516 79864 13556 79904
rect 2764 79780 2804 79820
rect 13324 79780 13364 79820
rect 17548 79780 17588 79820
rect 3244 79696 3284 79736
rect 11788 79696 11828 79736
rect 3532 79612 3572 79652
rect 3688 79360 3728 79400
rect 3770 79360 3810 79400
rect 3852 79360 3892 79400
rect 3934 79360 3974 79400
rect 4016 79360 4056 79400
rect 6508 79276 6548 79316
rect 15916 79276 15956 79316
rect 6028 79192 6068 79232
rect 18808 79360 18848 79400
rect 18890 79360 18930 79400
rect 18972 79360 19012 79400
rect 19054 79360 19094 79400
rect 19136 79360 19176 79400
rect 10924 79108 10964 79148
rect 18316 79108 18356 79148
rect 3436 78940 3476 78980
rect 5452 78940 5492 78980
rect 9868 78940 9908 78980
rect 5548 78772 5588 78812
rect 10444 78772 10484 78812
rect 4928 78604 4968 78644
rect 5010 78604 5050 78644
rect 5092 78604 5132 78644
rect 5174 78604 5214 78644
rect 5256 78604 5296 78644
rect 20048 78604 20088 78644
rect 20130 78604 20170 78644
rect 20212 78604 20252 78644
rect 20294 78604 20334 78644
rect 20376 78604 20416 78644
rect 17068 78436 17108 78476
rect 9580 78268 9620 78308
rect 13516 78268 13556 78308
rect 3436 78184 3476 78224
rect 8908 78100 8948 78140
rect 14956 78100 14996 78140
rect 17452 78100 17492 78140
rect 5548 78016 5588 78056
rect 3688 77848 3728 77888
rect 3770 77848 3810 77888
rect 3852 77848 3892 77888
rect 3934 77848 3974 77888
rect 4016 77848 4056 77888
rect 4300 77848 4340 77888
rect 18808 77848 18848 77888
rect 18890 77848 18930 77888
rect 18972 77848 19012 77888
rect 19054 77848 19094 77888
rect 19136 77848 19176 77888
rect 7948 77680 7988 77720
rect 16300 77680 16340 77720
rect 2284 77512 2324 77552
rect 2668 77428 2708 77468
rect 10348 77428 10388 77468
rect 17548 77428 17588 77468
rect 9196 77344 9236 77384
rect 3532 77176 3572 77216
rect 4928 77092 4968 77132
rect 5010 77092 5050 77132
rect 5092 77092 5132 77132
rect 5174 77092 5214 77132
rect 5256 77092 5296 77132
rect 2572 77008 2612 77048
rect 5548 76924 5588 76964
rect 10252 76924 10292 76964
rect 20048 77092 20088 77132
rect 20130 77092 20170 77132
rect 20212 77092 20252 77132
rect 20294 77092 20334 77132
rect 20376 77092 20416 77132
rect 1516 76756 1556 76796
rect 3244 76756 3284 76796
rect 3532 76588 3572 76628
rect 10348 76588 10388 76628
rect 2668 76336 2708 76376
rect 3688 76336 3728 76376
rect 3770 76336 3810 76376
rect 3852 76336 3892 76376
rect 3934 76336 3974 76376
rect 4016 76336 4056 76376
rect 5452 76336 5492 76376
rect 6028 76252 6068 76292
rect 8620 76252 8660 76292
rect 17932 76756 17972 76796
rect 14476 76672 14516 76712
rect 18316 76672 18356 76712
rect 10924 76588 10964 76628
rect 20524 76588 20564 76628
rect 12844 76420 12884 76460
rect 15820 76420 15860 76460
rect 15052 76336 15092 76376
rect 18808 76336 18848 76376
rect 18890 76336 18930 76376
rect 18972 76336 19012 76376
rect 19054 76336 19094 76376
rect 19136 76336 19176 76376
rect 15724 76252 15764 76292
rect 16492 76252 16532 76292
rect 7948 76084 7988 76124
rect 1228 76000 1268 76040
rect 18316 76000 18356 76040
rect 748 75916 788 75956
rect 6988 75916 7028 75956
rect 20620 75916 20660 75956
rect 3532 75832 3572 75872
rect 13996 75748 14036 75788
rect 4928 75580 4968 75620
rect 5010 75580 5050 75620
rect 5092 75580 5132 75620
rect 5174 75580 5214 75620
rect 5256 75580 5296 75620
rect 13804 75580 13844 75620
rect 364 75496 404 75536
rect 17548 75748 17588 75788
rect 20048 75580 20088 75620
rect 20130 75580 20170 75620
rect 20212 75580 20252 75620
rect 20294 75580 20334 75620
rect 20376 75580 20416 75620
rect 4780 75412 4820 75452
rect 4780 75244 4820 75284
rect 6796 75160 6836 75200
rect 6988 75076 7028 75116
rect 13324 75076 13364 75116
rect 7276 74992 7316 75032
rect 3688 74824 3728 74864
rect 3770 74824 3810 74864
rect 3852 74824 3892 74864
rect 3934 74824 3974 74864
rect 4016 74824 4056 74864
rect 18808 74824 18848 74864
rect 18890 74824 18930 74864
rect 18972 74824 19012 74864
rect 19054 74824 19094 74864
rect 19136 74824 19176 74864
rect 5452 74740 5492 74780
rect 5452 74572 5492 74612
rect 8908 74572 8948 74612
rect 6220 74488 6260 74528
rect 13132 74488 13172 74528
rect 12652 74404 12692 74444
rect 14476 74404 14516 74444
rect 17452 74404 17492 74444
rect 1420 74320 1460 74360
rect 3532 74320 3572 74360
rect 5452 74320 5492 74360
rect 1132 74236 1172 74276
rect 1324 74152 1364 74192
rect 3436 74152 3476 74192
rect 4780 74152 4820 74192
rect 4928 74068 4968 74108
rect 5010 74068 5050 74108
rect 5092 74068 5132 74108
rect 5174 74068 5214 74108
rect 5256 74068 5296 74108
rect 20048 74068 20088 74108
rect 20130 74068 20170 74108
rect 20212 74068 20252 74108
rect 20294 74068 20334 74108
rect 20376 74068 20416 74108
rect 364 73816 404 73856
rect 16012 73900 16052 73940
rect 10348 73648 10388 73688
rect 18316 73732 18356 73772
rect 4300 73564 4340 73604
rect 12844 73564 12884 73604
rect 2956 73480 2996 73520
rect 6028 73480 6068 73520
rect 9004 73480 9044 73520
rect 2188 73396 2228 73436
rect 15052 73480 15092 73520
rect 20620 73396 20660 73436
rect 3688 73312 3728 73352
rect 3770 73312 3810 73352
rect 3852 73312 3892 73352
rect 3934 73312 3974 73352
rect 4016 73312 4056 73352
rect 9196 73312 9236 73352
rect 13324 73312 13364 73352
rect 18808 73312 18848 73352
rect 18890 73312 18930 73352
rect 18972 73312 19012 73352
rect 19054 73312 19094 73352
rect 19136 73312 19176 73352
rect 8236 73228 8276 73268
rect 2572 73060 2612 73100
rect 12844 73060 12884 73100
rect 16012 72892 16052 72932
rect 6988 72724 7028 72764
rect 20524 72640 20564 72680
rect 4928 72556 4968 72596
rect 5010 72556 5050 72596
rect 5092 72556 5132 72596
rect 5174 72556 5214 72596
rect 5256 72556 5296 72596
rect 3244 72472 3284 72512
rect 4204 72472 4244 72512
rect 3148 72388 3188 72428
rect 4204 72304 4244 72344
rect 3532 72220 3572 72260
rect 9868 72136 9908 72176
rect 20048 72556 20088 72596
rect 20130 72556 20170 72596
rect 20212 72556 20252 72596
rect 20294 72556 20334 72596
rect 20376 72556 20416 72596
rect 18316 72388 18356 72428
rect 1708 72052 1748 72092
rect 5452 71968 5492 72008
rect 3688 71800 3728 71840
rect 3770 71800 3810 71840
rect 3852 71800 3892 71840
rect 3934 71800 3974 71840
rect 4016 71800 4056 71840
rect 18808 71800 18848 71840
rect 18890 71800 18930 71840
rect 18972 71800 19012 71840
rect 19054 71800 19094 71840
rect 19136 71800 19176 71840
rect 2188 71716 2228 71756
rect 2956 71716 2996 71756
rect 15628 71716 15668 71756
rect 3532 71632 3572 71672
rect 5644 71548 5684 71588
rect 10060 71548 10100 71588
rect 15916 71548 15956 71588
rect 7948 71464 7988 71504
rect 9676 71464 9716 71504
rect 1996 71380 2036 71420
rect 15820 71296 15860 71336
rect 17932 71296 17972 71336
rect 14572 71212 14612 71252
rect 15052 71212 15092 71252
rect 1804 71128 1844 71168
rect 4928 71044 4968 71084
rect 5010 71044 5050 71084
rect 5092 71044 5132 71084
rect 5174 71044 5214 71084
rect 5256 71044 5296 71084
rect 20048 71044 20088 71084
rect 20130 71044 20170 71084
rect 20212 71044 20252 71084
rect 20294 71044 20334 71084
rect 20376 71044 20416 71084
rect 4780 70876 4820 70916
rect 6988 70792 7028 70832
rect 748 70708 788 70748
rect 4780 70708 4820 70748
rect 6508 70708 6548 70748
rect 4300 70624 4340 70664
rect 9580 70624 9620 70664
rect 15052 70624 15092 70664
rect 5548 70540 5588 70580
rect 6220 70540 6260 70580
rect 7372 70540 7412 70580
rect 8908 70540 8948 70580
rect 9676 70540 9716 70580
rect 15628 70540 15668 70580
rect 15916 70540 15956 70580
rect 5644 70456 5684 70496
rect 12652 70456 12692 70496
rect 17932 70456 17972 70496
rect 3688 70288 3728 70328
rect 3770 70288 3810 70328
rect 3852 70288 3892 70328
rect 3934 70288 3974 70328
rect 4016 70288 4056 70328
rect 18808 70288 18848 70328
rect 18890 70288 18930 70328
rect 18972 70288 19012 70328
rect 19054 70288 19094 70328
rect 19136 70288 19176 70328
rect 7948 70204 7988 70244
rect 17452 70120 17492 70160
rect 1996 70036 2036 70076
rect 5836 70036 5876 70076
rect 10252 70036 10292 70076
rect 17260 70036 17300 70076
rect 2380 69952 2420 69992
rect 4300 69868 4340 69908
rect 20620 69784 20660 69824
rect 5548 69700 5588 69740
rect 11404 69700 11444 69740
rect 20524 69700 20564 69740
rect 4928 69532 4968 69572
rect 5010 69532 5050 69572
rect 5092 69532 5132 69572
rect 5174 69532 5214 69572
rect 5256 69532 5296 69572
rect 20048 69532 20088 69572
rect 20130 69532 20170 69572
rect 20212 69532 20252 69572
rect 20294 69532 20334 69572
rect 20376 69532 20416 69572
rect 7564 69364 7604 69404
rect 5836 69280 5876 69320
rect 16492 69280 16532 69320
rect 2860 69196 2900 69236
rect 3532 69196 3572 69236
rect 1708 69112 1748 69152
rect 10348 69112 10388 69152
rect 11884 69112 11924 69152
rect 13324 69112 13364 69152
rect 14476 69112 14516 69152
rect 20620 69112 20660 69152
rect 1228 68944 1268 68984
rect 20620 68944 20660 68984
rect 3688 68776 3728 68816
rect 3770 68776 3810 68816
rect 3852 68776 3892 68816
rect 3934 68776 3974 68816
rect 4016 68776 4056 68816
rect 4780 68440 4820 68480
rect 6508 68440 6548 68480
rect 5452 68356 5492 68396
rect 7660 68356 7700 68396
rect 5644 68272 5684 68312
rect 9004 68272 9044 68312
rect 18808 68776 18848 68816
rect 18890 68776 18930 68816
rect 18972 68776 19012 68816
rect 19054 68776 19094 68816
rect 19136 68776 19176 68816
rect 18316 68608 18356 68648
rect 13996 68356 14036 68396
rect 7948 68188 7988 68228
rect 8236 68188 8276 68228
rect 4928 68020 4968 68060
rect 5010 68020 5050 68060
rect 5092 68020 5132 68060
rect 5174 68020 5214 68060
rect 5256 68020 5296 68060
rect 4780 67852 4820 67892
rect 20048 68020 20088 68060
rect 20130 68020 20170 68060
rect 20212 68020 20252 68060
rect 20294 68020 20334 68060
rect 20376 68020 20416 68060
rect 20524 67852 20564 67892
rect 1420 67600 1460 67640
rect 3532 67600 3572 67640
rect 6796 67600 6836 67640
rect 7372 67600 7412 67640
rect 10252 67516 10292 67556
rect 2188 67432 2228 67472
rect 3532 67432 3572 67472
rect 6796 67432 6836 67472
rect 3688 67264 3728 67304
rect 3770 67264 3810 67304
rect 3852 67264 3892 67304
rect 3934 67264 3974 67304
rect 4016 67264 4056 67304
rect 18808 67264 18848 67304
rect 18890 67264 18930 67304
rect 18972 67264 19012 67304
rect 19054 67264 19094 67304
rect 19136 67264 19176 67304
rect 1804 67180 1844 67220
rect 2092 67096 2132 67136
rect 13132 67096 13172 67136
rect 3532 67012 3572 67052
rect 1420 66928 1460 66968
rect 5548 66928 5588 66968
rect 6028 66928 6068 66968
rect 11692 66928 11732 66968
rect 1996 66844 2036 66884
rect 20620 66676 20660 66716
rect 4928 66508 4968 66548
rect 5010 66508 5050 66548
rect 5092 66508 5132 66548
rect 5174 66508 5214 66548
rect 5256 66508 5296 66548
rect 11692 66508 11732 66548
rect 20048 66508 20088 66548
rect 20130 66508 20170 66548
rect 20212 66508 20252 66548
rect 20294 66508 20334 66548
rect 20376 66508 20416 66548
rect 1708 66256 1748 66296
rect 2668 66256 2708 66296
rect 12460 66340 12500 66380
rect 15436 66256 15476 66296
rect 17932 66256 17972 66296
rect 3532 66172 3572 66212
rect 4300 66172 4340 66212
rect 10636 66172 10676 66212
rect 15628 66172 15668 66212
rect 6988 66088 7028 66128
rect 2860 65920 2900 65960
rect 3688 65752 3728 65792
rect 3770 65752 3810 65792
rect 3852 65752 3892 65792
rect 3934 65752 3974 65792
rect 4016 65752 4056 65792
rect 16492 65752 16532 65792
rect 18808 65752 18848 65792
rect 18890 65752 18930 65792
rect 18972 65752 19012 65792
rect 19054 65752 19094 65792
rect 19136 65752 19176 65792
rect 4204 65584 4244 65624
rect 2092 65500 2132 65540
rect 3148 65416 3188 65456
rect 2572 65248 2612 65288
rect 15436 65248 15476 65288
rect 11308 65164 11348 65204
rect 3244 65080 3284 65120
rect 4928 64996 4968 65036
rect 5010 64996 5050 65036
rect 5092 64996 5132 65036
rect 5174 64996 5214 65036
rect 5256 64996 5296 65036
rect 13132 65080 13172 65120
rect 13228 64996 13268 65036
rect 20048 64996 20088 65036
rect 20130 64996 20170 65036
rect 20212 64996 20252 65036
rect 20294 64996 20334 65036
rect 20376 64996 20416 65036
rect 9196 64912 9236 64952
rect 13516 64828 13556 64868
rect 2860 64744 2900 64784
rect 5548 64744 5588 64784
rect 6124 64744 6164 64784
rect 3532 64660 3572 64700
rect 8908 64660 8948 64700
rect 2956 64576 2996 64616
rect 3436 64576 3476 64616
rect 5836 64576 5876 64616
rect 6124 64492 6164 64532
rect 1708 64408 1748 64448
rect 3688 64240 3728 64280
rect 3770 64240 3810 64280
rect 3852 64240 3892 64280
rect 3934 64240 3974 64280
rect 4016 64240 4056 64280
rect 18808 64240 18848 64280
rect 18890 64240 18930 64280
rect 18972 64240 19012 64280
rect 19054 64240 19094 64280
rect 19136 64240 19176 64280
rect 2188 64156 2228 64196
rect 12556 64156 12596 64196
rect 18220 64156 18260 64196
rect 2188 63988 2228 64028
rect 2380 63988 2420 64028
rect 2668 63904 2708 63944
rect 2956 63904 2996 63944
rect 4780 64072 4820 64112
rect 7084 64072 7124 64112
rect 8908 63988 8948 64028
rect 18220 63988 18260 64028
rect 4204 63904 4244 63944
rect 4780 63904 4820 63944
rect 1996 63820 2036 63860
rect 3244 63736 3284 63776
rect 2572 63652 2612 63692
rect 5644 63652 5684 63692
rect 6796 63652 6836 63692
rect 11500 63652 11540 63692
rect 14476 63652 14516 63692
rect 18316 63652 18356 63692
rect 4300 63568 4340 63608
rect 15244 63568 15284 63608
rect 3148 63484 3188 63524
rect 3436 63484 3476 63524
rect 4928 63484 4968 63524
rect 5010 63484 5050 63524
rect 5092 63484 5132 63524
rect 5174 63484 5214 63524
rect 5256 63484 5296 63524
rect 8908 63484 8948 63524
rect 20048 63484 20088 63524
rect 20130 63484 20170 63524
rect 20212 63484 20252 63524
rect 20294 63484 20334 63524
rect 20376 63484 20416 63524
rect 1516 63316 1556 63356
rect 1708 63316 1748 63356
rect 2668 63316 2708 63356
rect 2860 63316 2900 63356
rect 5644 63316 5684 63356
rect 6124 63316 6164 63356
rect 3052 63232 3092 63272
rect 3532 63232 3572 63272
rect 12460 63400 12500 63440
rect 13516 63232 13556 63272
rect 18220 63232 18260 63272
rect 9676 63148 9716 63188
rect 4780 63064 4820 63104
rect 7948 63064 7988 63104
rect 13324 63064 13364 63104
rect 17932 63064 17972 63104
rect 18220 63064 18260 63104
rect 2956 62980 2996 63020
rect 1420 62896 1460 62936
rect 13996 62896 14036 62936
rect 7084 62812 7124 62852
rect 11884 62812 11924 62852
rect 12268 62812 12308 62852
rect 15244 62812 15284 62852
rect 17932 62812 17972 62852
rect 18316 62812 18356 62852
rect 3688 62728 3728 62768
rect 3770 62728 3810 62768
rect 3852 62728 3892 62768
rect 3934 62728 3974 62768
rect 4016 62728 4056 62768
rect 18808 62728 18848 62768
rect 18890 62728 18930 62768
rect 18972 62728 19012 62768
rect 19054 62728 19094 62768
rect 19136 62728 19176 62768
rect 15436 62644 15476 62684
rect 20620 63400 20660 63440
rect 13132 62476 13172 62516
rect 17260 62476 17300 62516
rect 9196 62392 9236 62432
rect 15244 62392 15284 62432
rect 16012 62392 16052 62432
rect 4204 62308 4244 62348
rect 17932 62308 17972 62348
rect 3148 62140 3188 62180
rect 4780 62140 4820 62180
rect 9004 62056 9044 62096
rect 11116 62056 11156 62096
rect 4928 61972 4968 62012
rect 5010 61972 5050 62012
rect 5092 61972 5132 62012
rect 5174 61972 5214 62012
rect 5256 61972 5296 62012
rect 9196 61972 9236 62012
rect 10156 61972 10196 62012
rect 20048 61972 20088 62012
rect 20130 61972 20170 62012
rect 20212 61972 20252 62012
rect 20294 61972 20334 62012
rect 20376 61972 20416 62012
rect 11116 61804 11156 61844
rect 3532 61636 3572 61676
rect 16012 61636 16052 61676
rect 4300 61552 4340 61592
rect 18220 61552 18260 61592
rect 2572 61468 2612 61508
rect 6028 61468 6068 61508
rect 7084 61468 7124 61508
rect 15628 61468 15668 61508
rect 17452 61468 17492 61508
rect 3688 61216 3728 61256
rect 3770 61216 3810 61256
rect 3852 61216 3892 61256
rect 3934 61216 3974 61256
rect 4016 61216 4056 61256
rect 18808 61216 18848 61256
rect 18890 61216 18930 61256
rect 18972 61216 19012 61256
rect 19054 61216 19094 61256
rect 19136 61216 19176 61256
rect 12268 61132 12308 61172
rect 3532 61048 3572 61088
rect 3436 60964 3476 61004
rect 4204 60880 4244 60920
rect 4204 60712 4244 60752
rect 6124 60712 6164 60752
rect 7372 60712 7412 60752
rect 12172 60544 12212 60584
rect 17260 60544 17300 60584
rect 4928 60460 4968 60500
rect 5010 60460 5050 60500
rect 5092 60460 5132 60500
rect 5174 60460 5214 60500
rect 5256 60460 5296 60500
rect 11596 60460 11636 60500
rect 12460 60460 12500 60500
rect 15532 60460 15572 60500
rect 16396 60460 16436 60500
rect 20048 60460 20088 60500
rect 20130 60460 20170 60500
rect 20212 60460 20252 60500
rect 20294 60460 20334 60500
rect 20376 60460 20416 60500
rect 2476 60376 2516 60416
rect 12652 60292 12692 60332
rect 1900 60208 1940 60248
rect 11884 60208 11924 60248
rect 3436 60124 3476 60164
rect 8716 60124 8756 60164
rect 14476 60040 14516 60080
rect 11884 59956 11924 59996
rect 12844 59872 12884 59912
rect 3688 59704 3728 59744
rect 3770 59704 3810 59744
rect 3852 59704 3892 59744
rect 3934 59704 3974 59744
rect 4016 59704 4056 59744
rect 6988 59704 7028 59744
rect 17836 59704 17876 59744
rect 18808 59704 18848 59744
rect 18890 59704 18930 59744
rect 18972 59704 19012 59744
rect 19054 59704 19094 59744
rect 19136 59704 19176 59744
rect 12172 59620 12212 59660
rect 2092 59368 2132 59408
rect 1516 59284 1556 59324
rect 18316 59284 18356 59324
rect 11884 59200 11924 59240
rect 15436 59116 15476 59156
rect 4928 58948 4968 58988
rect 5010 58948 5050 58988
rect 5092 58948 5132 58988
rect 5174 58948 5214 58988
rect 5256 58948 5296 58988
rect 20048 58948 20088 58988
rect 20130 58948 20170 58988
rect 20212 58948 20252 58988
rect 20294 58948 20334 58988
rect 20376 58948 20416 58988
rect 5644 58780 5684 58820
rect 20524 58780 20564 58820
rect 13132 58696 13172 58736
rect 11596 58528 11636 58568
rect 13132 58528 13172 58568
rect 17260 58528 17300 58568
rect 18220 58360 18260 58400
rect 6412 58276 6452 58316
rect 3052 58192 3092 58232
rect 3688 58192 3728 58232
rect 3770 58192 3810 58232
rect 3852 58192 3892 58232
rect 3934 58192 3974 58232
rect 4016 58192 4056 58232
rect 12172 58192 12212 58232
rect 18808 58192 18848 58232
rect 18890 58192 18930 58232
rect 18972 58192 19012 58232
rect 19054 58192 19094 58232
rect 19136 58192 19176 58232
rect 12268 57940 12308 57980
rect 17452 57856 17492 57896
rect 4204 57772 4244 57812
rect 11404 57604 11444 57644
rect 17068 57604 17108 57644
rect 11596 57520 11636 57560
rect 4928 57436 4968 57476
rect 5010 57436 5050 57476
rect 5092 57436 5132 57476
rect 5174 57436 5214 57476
rect 5256 57436 5296 57476
rect 20048 57436 20088 57476
rect 20130 57436 20170 57476
rect 20212 57436 20252 57476
rect 20294 57436 20334 57476
rect 20376 57436 20416 57476
rect 5644 56932 5684 56972
rect 3688 56680 3728 56720
rect 3770 56680 3810 56720
rect 3852 56680 3892 56720
rect 3934 56680 3974 56720
rect 4016 56680 4056 56720
rect 18808 56680 18848 56720
rect 18890 56680 18930 56720
rect 18972 56680 19012 56720
rect 19054 56680 19094 56720
rect 19136 56680 19176 56720
rect 9292 56512 9332 56552
rect 6412 56344 6452 56384
rect 17644 56344 17684 56384
rect 18316 56344 18356 56384
rect 17068 56176 17108 56216
rect 17836 56176 17876 56216
rect 8812 56092 8852 56132
rect 16492 56092 16532 56132
rect 4928 55924 4968 55964
rect 5010 55924 5050 55964
rect 5092 55924 5132 55964
rect 5174 55924 5214 55964
rect 5256 55924 5296 55964
rect 20048 55924 20088 55964
rect 20130 55924 20170 55964
rect 20212 55924 20252 55964
rect 20294 55924 20334 55964
rect 20376 55924 20416 55964
rect 18412 55504 18452 55544
rect 6220 55336 6260 55376
rect 3688 55168 3728 55208
rect 3770 55168 3810 55208
rect 3852 55168 3892 55208
rect 3934 55168 3974 55208
rect 4016 55168 4056 55208
rect 18808 55168 18848 55208
rect 18890 55168 18930 55208
rect 18972 55168 19012 55208
rect 19054 55168 19094 55208
rect 19136 55168 19176 55208
rect 1708 54916 1748 54956
rect 3244 54748 3284 54788
rect 4780 54748 4820 54788
rect 4928 54412 4968 54452
rect 5010 54412 5050 54452
rect 5092 54412 5132 54452
rect 5174 54412 5214 54452
rect 5256 54412 5296 54452
rect 20048 54412 20088 54452
rect 20130 54412 20170 54452
rect 20212 54412 20252 54452
rect 20294 54412 20334 54452
rect 20376 54412 20416 54452
rect 5932 54328 5972 54368
rect 1612 54244 1652 54284
rect 7948 54244 7988 54284
rect 9868 54160 9908 54200
rect 18316 53992 18356 54032
rect 3244 53824 3284 53864
rect 3688 53656 3728 53696
rect 3770 53656 3810 53696
rect 3852 53656 3892 53696
rect 3934 53656 3974 53696
rect 4016 53656 4056 53696
rect 18808 53656 18848 53696
rect 18890 53656 18930 53696
rect 18972 53656 19012 53696
rect 19054 53656 19094 53696
rect 19136 53656 19176 53696
rect 2188 53488 2228 53528
rect 9964 53488 10004 53528
rect 10636 53404 10676 53444
rect 2668 53320 2708 53360
rect 2860 53320 2900 53360
rect 13324 53320 13364 53360
rect 16012 53320 16052 53360
rect 17452 53320 17492 53360
rect 2668 53068 2708 53108
rect 2860 53068 2900 53108
rect 4928 52900 4968 52940
rect 5010 52900 5050 52940
rect 5092 52900 5132 52940
rect 5174 52900 5214 52940
rect 5256 52900 5296 52940
rect 20048 52900 20088 52940
rect 20130 52900 20170 52940
rect 20212 52900 20252 52940
rect 20294 52900 20334 52940
rect 20376 52900 20416 52940
rect 8812 52816 8852 52856
rect 10444 52480 10484 52520
rect 3688 52144 3728 52184
rect 3770 52144 3810 52184
rect 3852 52144 3892 52184
rect 3934 52144 3974 52184
rect 4016 52144 4056 52184
rect 15628 52144 15668 52184
rect 18808 52144 18848 52184
rect 18890 52144 18930 52184
rect 18972 52144 19012 52184
rect 19054 52144 19094 52184
rect 19136 52144 19176 52184
rect 9772 51892 9812 51932
rect 16396 51892 16436 51932
rect 18028 51892 18068 51932
rect 18412 51892 18452 51932
rect 1804 51808 1844 51848
rect 15340 51808 15380 51848
rect 4928 51388 4968 51428
rect 5010 51388 5050 51428
rect 5092 51388 5132 51428
rect 5174 51388 5214 51428
rect 5256 51388 5296 51428
rect 20048 51388 20088 51428
rect 20130 51388 20170 51428
rect 20212 51388 20252 51428
rect 20294 51388 20334 51428
rect 20376 51388 20416 51428
rect 11212 51052 11252 51092
rect 2572 50968 2612 51008
rect 2380 50800 2420 50840
rect 3688 50632 3728 50672
rect 3770 50632 3810 50672
rect 3852 50632 3892 50672
rect 3934 50632 3974 50672
rect 4016 50632 4056 50672
rect 18808 50632 18848 50672
rect 18890 50632 18930 50672
rect 18972 50632 19012 50672
rect 19054 50632 19094 50672
rect 19136 50632 19176 50672
rect 6796 50380 6836 50420
rect 10828 50296 10868 50336
rect 11404 50296 11444 50336
rect 12268 50296 12308 50336
rect 12652 50296 12692 50336
rect 10348 50212 10388 50252
rect 12364 50212 12404 50252
rect 11020 50128 11060 50168
rect 11212 50044 11252 50084
rect 4928 49876 4968 49916
rect 5010 49876 5050 49916
rect 5092 49876 5132 49916
rect 5174 49876 5214 49916
rect 5256 49876 5296 49916
rect 20048 49876 20088 49916
rect 20130 49876 20170 49916
rect 20212 49876 20252 49916
rect 20294 49876 20334 49916
rect 20376 49876 20416 49916
rect 16108 49624 16148 49664
rect 9580 49540 9620 49580
rect 10156 49540 10196 49580
rect 10828 49540 10868 49580
rect 20620 49456 20660 49496
rect 17644 49288 17684 49328
rect 3688 49120 3728 49160
rect 3770 49120 3810 49160
rect 3852 49120 3892 49160
rect 3934 49120 3974 49160
rect 4016 49120 4056 49160
rect 18808 49120 18848 49160
rect 18890 49120 18930 49160
rect 18972 49120 19012 49160
rect 19054 49120 19094 49160
rect 19136 49120 19176 49160
rect 15916 48952 15956 48992
rect 10540 48868 10580 48908
rect 10732 48868 10772 48908
rect 9676 48784 9716 48824
rect 10060 48784 10100 48824
rect 6124 48700 6164 48740
rect 9772 48700 9812 48740
rect 12748 48700 12788 48740
rect 13420 48700 13460 48740
rect 9388 48616 9428 48656
rect 4204 48532 4244 48572
rect 7372 48448 7412 48488
rect 4928 48364 4968 48404
rect 5010 48364 5050 48404
rect 5092 48364 5132 48404
rect 5174 48364 5214 48404
rect 5256 48364 5296 48404
rect 8716 48364 8756 48404
rect 19756 48364 19796 48404
rect 20048 48364 20088 48404
rect 20130 48364 20170 48404
rect 20212 48364 20252 48404
rect 20294 48364 20334 48404
rect 20376 48364 20416 48404
rect 19276 48196 19316 48236
rect 19756 48196 19796 48236
rect 2476 48028 2516 48068
rect 10252 48028 10292 48068
rect 19276 48028 19316 48068
rect 9196 47944 9236 47984
rect 12172 47944 12212 47984
rect 10540 47860 10580 47900
rect 3688 47608 3728 47648
rect 3770 47608 3810 47648
rect 3852 47608 3892 47648
rect 3934 47608 3974 47648
rect 4016 47608 4056 47648
rect 18808 47608 18848 47648
rect 18890 47608 18930 47648
rect 18972 47608 19012 47648
rect 19054 47608 19094 47648
rect 19136 47608 19176 47648
rect 9196 47188 9236 47228
rect 10540 47188 10580 47228
rect 4928 46852 4968 46892
rect 5010 46852 5050 46892
rect 5092 46852 5132 46892
rect 5174 46852 5214 46892
rect 5256 46852 5296 46892
rect 20048 46852 20088 46892
rect 20130 46852 20170 46892
rect 20212 46852 20252 46892
rect 20294 46852 20334 46892
rect 20376 46852 20416 46892
rect 3340 46684 3380 46724
rect 4492 46684 4532 46724
rect 10444 46516 10484 46556
rect 13516 46432 13556 46472
rect 12556 46264 12596 46304
rect 3688 46096 3728 46136
rect 3770 46096 3810 46136
rect 3852 46096 3892 46136
rect 3934 46096 3974 46136
rect 4016 46096 4056 46136
rect 18808 46096 18848 46136
rect 18890 46096 18930 46136
rect 18972 46096 19012 46136
rect 19054 46096 19094 46136
rect 19136 46096 19176 46136
rect 5644 46012 5684 46052
rect 9196 45676 9236 45716
rect 4492 45340 4532 45380
rect 4928 45340 4968 45380
rect 5010 45340 5050 45380
rect 5092 45340 5132 45380
rect 5174 45340 5214 45380
rect 5256 45340 5296 45380
rect 20048 45340 20088 45380
rect 20130 45340 20170 45380
rect 20212 45340 20252 45380
rect 20294 45340 20334 45380
rect 20376 45340 20416 45380
rect 21388 45256 21428 45296
rect 5644 45172 5684 45212
rect 18028 45172 18068 45212
rect 13996 44920 14036 44960
rect 21388 44920 21428 44960
rect 1996 44752 2036 44792
rect 2668 44752 2708 44792
rect 3688 44584 3728 44624
rect 3770 44584 3810 44624
rect 3852 44584 3892 44624
rect 3934 44584 3974 44624
rect 4016 44584 4056 44624
rect 6508 44584 6548 44624
rect 18808 44584 18848 44624
rect 18890 44584 18930 44624
rect 18972 44584 19012 44624
rect 19054 44584 19094 44624
rect 19136 44584 19176 44624
rect 5644 44332 5684 44372
rect 5932 44332 5972 44372
rect 9964 44164 10004 44204
rect 6508 44080 6548 44120
rect 4300 43996 4340 44036
rect 4928 43828 4968 43868
rect 5010 43828 5050 43868
rect 5092 43828 5132 43868
rect 5174 43828 5214 43868
rect 5256 43828 5296 43868
rect 20048 43828 20088 43868
rect 20130 43828 20170 43868
rect 20212 43828 20252 43868
rect 20294 43828 20334 43868
rect 20376 43828 20416 43868
rect 4780 43660 4820 43700
rect 5644 43660 5684 43700
rect 4492 43576 4532 43616
rect 11020 43492 11060 43532
rect 6508 43408 6548 43448
rect 2188 43240 2228 43280
rect 5932 43240 5972 43280
rect 12940 43240 12980 43280
rect 2572 43072 2612 43112
rect 3688 43072 3728 43112
rect 3770 43072 3810 43112
rect 3852 43072 3892 43112
rect 3934 43072 3974 43112
rect 4016 43072 4056 43112
rect 4300 43072 4340 43112
rect 5932 43072 5972 43112
rect 18808 43072 18848 43112
rect 18890 43072 18930 43112
rect 18972 43072 19012 43112
rect 19054 43072 19094 43112
rect 19136 43072 19176 43112
rect 5932 42904 5972 42944
rect 13036 42820 13076 42860
rect 13420 42820 13460 42860
rect 10828 42400 10868 42440
rect 13708 42400 13748 42440
rect 4928 42316 4968 42356
rect 5010 42316 5050 42356
rect 5092 42316 5132 42356
rect 5174 42316 5214 42356
rect 5256 42316 5296 42356
rect 20048 42316 20088 42356
rect 20130 42316 20170 42356
rect 20212 42316 20252 42356
rect 20294 42316 20334 42356
rect 20376 42316 20416 42356
rect 13708 42232 13748 42272
rect 4492 41812 4532 41852
rect 4780 41812 4820 41852
rect 3688 41560 3728 41600
rect 3770 41560 3810 41600
rect 3852 41560 3892 41600
rect 3934 41560 3974 41600
rect 4016 41560 4056 41600
rect 4300 41560 4340 41600
rect 18808 41560 18848 41600
rect 18890 41560 18930 41600
rect 18972 41560 19012 41600
rect 19054 41560 19094 41600
rect 19136 41560 19176 41600
rect 9292 41476 9332 41516
rect 4588 41392 4628 41432
rect 3148 41308 3188 41348
rect 4780 41308 4820 41348
rect 6028 41140 6068 41180
rect 10732 41056 10772 41096
rect 6124 40972 6164 41012
rect 10540 40972 10580 41012
rect 9196 40888 9236 40928
rect 4928 40804 4968 40844
rect 5010 40804 5050 40844
rect 5092 40804 5132 40844
rect 5174 40804 5214 40844
rect 5256 40804 5296 40844
rect 6124 40804 6164 40844
rect 10540 40804 10580 40844
rect 11308 40804 11348 40844
rect 20048 40804 20088 40844
rect 20130 40804 20170 40844
rect 20212 40804 20252 40844
rect 20294 40804 20334 40844
rect 20376 40804 20416 40844
rect 1516 40720 1556 40760
rect 4588 40468 4628 40508
rect 6124 40384 6164 40424
rect 13996 40384 14036 40424
rect 18124 40384 18164 40424
rect 5740 40300 5780 40340
rect 12844 40300 12884 40340
rect 13420 40300 13460 40340
rect 15436 40300 15476 40340
rect 3532 40216 3572 40256
rect 6700 40132 6740 40172
rect 7084 40132 7124 40172
rect 3688 40048 3728 40088
rect 3770 40048 3810 40088
rect 3852 40048 3892 40088
rect 3934 40048 3974 40088
rect 4016 40048 4056 40088
rect 18808 40048 18848 40088
rect 18890 40048 18930 40088
rect 18972 40048 19012 40088
rect 19054 40048 19094 40088
rect 19136 40048 19176 40088
rect 10348 39964 10388 40004
rect 15820 39964 15860 40004
rect 8620 39880 8660 39920
rect 10444 39796 10484 39836
rect 18124 39796 18164 39836
rect 12364 39712 12404 39752
rect 12940 39712 12980 39752
rect 13420 39712 13460 39752
rect 16876 39712 16916 39752
rect 2956 39628 2996 39668
rect 6508 39628 6548 39668
rect 17260 39628 17300 39668
rect 2284 39544 2324 39584
rect 4300 39460 4340 39500
rect 6700 39460 6740 39500
rect 9196 39376 9236 39416
rect 13708 39376 13748 39416
rect 4300 39292 4340 39332
rect 4928 39292 4968 39332
rect 5010 39292 5050 39332
rect 5092 39292 5132 39332
rect 5174 39292 5214 39332
rect 5256 39292 5296 39332
rect 20048 39292 20088 39332
rect 20130 39292 20170 39332
rect 20212 39292 20252 39332
rect 20294 39292 20334 39332
rect 20376 39292 20416 39332
rect 16876 39124 16916 39164
rect 3052 38956 3092 38996
rect 7660 38956 7700 38996
rect 12940 38956 12980 38996
rect 18604 38956 18644 38996
rect 11308 38872 11348 38912
rect 8044 38788 8084 38828
rect 18604 38788 18644 38828
rect 13996 38704 14036 38744
rect 3688 38536 3728 38576
rect 3770 38536 3810 38576
rect 3852 38536 3892 38576
rect 3934 38536 3974 38576
rect 4016 38536 4056 38576
rect 18808 38536 18848 38576
rect 18890 38536 18930 38576
rect 18972 38536 19012 38576
rect 19054 38536 19094 38576
rect 19136 38536 19176 38576
rect 5644 38452 5684 38492
rect 15724 38368 15764 38408
rect 19468 38284 19508 38324
rect 14476 38200 14516 38240
rect 4396 38116 4436 38156
rect 5740 38116 5780 38156
rect 6796 38032 6836 38072
rect 18028 38116 18068 38156
rect 18316 38116 18356 38156
rect 19276 38116 19316 38156
rect 19468 38116 19508 38156
rect 15532 38032 15572 38072
rect 19276 37948 19316 37988
rect 12748 37864 12788 37904
rect 4928 37780 4968 37820
rect 5010 37780 5050 37820
rect 5092 37780 5132 37820
rect 5174 37780 5214 37820
rect 5256 37780 5296 37820
rect 20048 37780 20088 37820
rect 20130 37780 20170 37820
rect 20212 37780 20252 37820
rect 20294 37780 20334 37820
rect 20376 37780 20416 37820
rect 10540 37528 10580 37568
rect 11308 37528 11348 37568
rect 18124 37528 18164 37568
rect 3340 37444 3380 37484
rect 17356 37360 17396 37400
rect 10348 37276 10388 37316
rect 17356 37192 17396 37232
rect 17836 37192 17876 37232
rect 7084 37108 7124 37148
rect 3688 37024 3728 37064
rect 3770 37024 3810 37064
rect 3852 37024 3892 37064
rect 3934 37024 3974 37064
rect 4016 37024 4056 37064
rect 18808 37024 18848 37064
rect 18890 37024 18930 37064
rect 18972 37024 19012 37064
rect 19054 37024 19094 37064
rect 19136 37024 19176 37064
rect 5932 36940 5972 36980
rect 2284 36772 2324 36812
rect 3532 36688 3572 36728
rect 12364 36688 12404 36728
rect 13708 36604 13748 36644
rect 3532 36520 3572 36560
rect 4928 36268 4968 36308
rect 5010 36268 5050 36308
rect 5092 36268 5132 36308
rect 5174 36268 5214 36308
rect 5256 36268 5296 36308
rect 20048 36268 20088 36308
rect 20130 36268 20170 36308
rect 20212 36268 20252 36308
rect 20294 36268 20334 36308
rect 20376 36268 20416 36308
rect 4300 36100 4340 36140
rect 13516 36016 13556 36056
rect 15916 36016 15956 36056
rect 3532 35932 3572 35972
rect 14956 35764 14996 35804
rect 12364 35680 12404 35720
rect 3688 35512 3728 35552
rect 3770 35512 3810 35552
rect 3852 35512 3892 35552
rect 3934 35512 3974 35552
rect 4016 35512 4056 35552
rect 15916 35512 15956 35552
rect 18808 35512 18848 35552
rect 18890 35512 18930 35552
rect 18972 35512 19012 35552
rect 19054 35512 19094 35552
rect 19136 35512 19176 35552
rect 7180 35428 7220 35468
rect 15340 35344 15380 35384
rect 1612 35260 1652 35300
rect 2092 35260 2132 35300
rect 13420 35260 13460 35300
rect 18028 35176 18068 35216
rect 2956 35008 2996 35048
rect 13708 35008 13748 35048
rect 17836 34924 17876 34964
rect 4928 34756 4968 34796
rect 5010 34756 5050 34796
rect 5092 34756 5132 34796
rect 5174 34756 5214 34796
rect 5256 34756 5296 34796
rect 20048 34756 20088 34796
rect 20130 34756 20170 34796
rect 20212 34756 20252 34796
rect 20294 34756 20334 34796
rect 20376 34756 20416 34796
rect 7084 34672 7124 34712
rect 5932 34588 5972 34628
rect 13516 34588 13556 34628
rect 4300 34504 4340 34544
rect 4780 34504 4820 34544
rect 6700 34504 6740 34544
rect 10732 34504 10772 34544
rect 12460 34504 12500 34544
rect 13804 34504 13844 34544
rect 16684 34504 16724 34544
rect 3148 34420 3188 34460
rect 13612 34420 13652 34460
rect 14956 34420 14996 34460
rect 21196 34420 21236 34460
rect 1708 34252 1748 34292
rect 7468 34336 7508 34376
rect 3688 34000 3728 34040
rect 3770 34000 3810 34040
rect 3852 34000 3892 34040
rect 3934 34000 3974 34040
rect 4016 34000 4056 34040
rect 2956 33664 2996 33704
rect 18124 34168 18164 34208
rect 13036 33832 13076 33872
rect 18808 34000 18848 34040
rect 18890 34000 18930 34040
rect 18972 34000 19012 34040
rect 19054 34000 19094 34040
rect 19136 34000 19176 34040
rect 2284 33580 2324 33620
rect 14860 33580 14900 33620
rect 1996 33496 2036 33536
rect 2860 33496 2900 33536
rect 2284 33328 2324 33368
rect 3052 33328 3092 33368
rect 11596 33328 11636 33368
rect 12364 33328 12404 33368
rect 3148 33244 3188 33284
rect 4300 33244 4340 33284
rect 4928 33244 4968 33284
rect 5010 33244 5050 33284
rect 5092 33244 5132 33284
rect 5174 33244 5214 33284
rect 5256 33244 5296 33284
rect 11404 33244 11444 33284
rect 13708 33244 13748 33284
rect 18604 33244 18644 33284
rect 3052 33160 3092 33200
rect 4396 33160 4436 33200
rect 12364 33160 12404 33200
rect 18124 33160 18164 33200
rect 1516 33076 1556 33116
rect 12940 33076 12980 33116
rect 13420 33076 13460 33116
rect 18028 33076 18068 33116
rect 2188 32992 2228 33032
rect 2860 32992 2900 33032
rect 1804 32908 1844 32948
rect 4396 32908 4436 32948
rect 11308 32992 11348 33032
rect 15820 32908 15860 32948
rect 18124 32908 18164 32948
rect 1612 32824 1652 32864
rect 2092 32824 2132 32864
rect 7084 32824 7124 32864
rect 17836 32824 17876 32864
rect 20524 33328 20564 33368
rect 20048 33244 20088 33284
rect 20130 33244 20170 33284
rect 20212 33244 20252 33284
rect 20294 33244 20334 33284
rect 20376 33244 20416 33284
rect 18604 33076 18644 33116
rect 20524 32992 20564 33032
rect 4396 32740 4436 32780
rect 18124 32740 18164 32780
rect 7660 32656 7700 32696
rect 3688 32488 3728 32528
rect 3770 32488 3810 32528
rect 3852 32488 3892 32528
rect 3934 32488 3974 32528
rect 4016 32488 4056 32528
rect 17260 32488 17300 32528
rect 8620 32404 8660 32444
rect 18808 32488 18848 32528
rect 18890 32488 18930 32528
rect 18972 32488 19012 32528
rect 19054 32488 19094 32528
rect 19136 32488 19176 32528
rect 8044 32320 8084 32360
rect 3244 32236 3284 32276
rect 4300 32236 4340 32276
rect 10732 32236 10772 32276
rect 13612 32236 13652 32276
rect 11980 32152 12020 32192
rect 3244 32068 3284 32108
rect 9196 32068 9236 32108
rect 10444 32068 10484 32108
rect 15820 32068 15860 32108
rect 16108 32068 16148 32108
rect 1612 31984 1652 32024
rect 10540 31984 10580 32024
rect 2956 31900 2996 31940
rect 6796 31900 6836 31940
rect 4780 31732 4820 31772
rect 4928 31732 4968 31772
rect 5010 31732 5050 31772
rect 5092 31732 5132 31772
rect 5174 31732 5214 31772
rect 5256 31732 5296 31772
rect 11116 31564 11156 31604
rect 20048 31732 20088 31772
rect 20130 31732 20170 31772
rect 20212 31732 20252 31772
rect 20294 31732 20334 31772
rect 20376 31732 20416 31772
rect 11308 31396 11348 31436
rect 14188 31396 14228 31436
rect 13804 31312 13844 31352
rect 17068 31228 17108 31268
rect 5740 31144 5780 31184
rect 4396 31060 4436 31100
rect 3688 30976 3728 31016
rect 3770 30976 3810 31016
rect 3852 30976 3892 31016
rect 3934 30976 3974 31016
rect 4016 30976 4056 31016
rect 18808 30976 18848 31016
rect 18890 30976 18930 31016
rect 18972 30976 19012 31016
rect 19054 30976 19094 31016
rect 19136 30976 19176 31016
rect 15532 30892 15572 30932
rect 4396 30808 4436 30848
rect 10828 30808 10868 30848
rect 16876 30808 16916 30848
rect 18508 30640 18548 30680
rect 7948 30556 7988 30596
rect 8620 30388 8660 30428
rect 18124 30388 18164 30428
rect 6124 30304 6164 30344
rect 12364 30304 12404 30344
rect 17932 30304 17972 30344
rect 20524 30304 20564 30344
rect 1708 30220 1748 30260
rect 4928 30220 4968 30260
rect 5010 30220 5050 30260
rect 5092 30220 5132 30260
rect 5174 30220 5214 30260
rect 5256 30220 5296 30260
rect 12268 30220 12308 30260
rect 14188 30220 14228 30260
rect 16108 30220 16148 30260
rect 20048 30220 20088 30260
rect 20130 30220 20170 30260
rect 20212 30220 20252 30260
rect 20294 30220 20334 30260
rect 20376 30220 20416 30260
rect 7468 30136 7508 30176
rect 15916 30136 15956 30176
rect 18124 30136 18164 30176
rect 7948 30052 7988 30092
rect 12460 30052 12500 30092
rect 13420 30052 13460 30092
rect 18028 30052 18068 30092
rect 10444 29884 10484 29924
rect 12940 29884 12980 29924
rect 14956 29968 14996 30008
rect 15724 29968 15764 30008
rect 18508 29968 18548 30008
rect 1324 29800 1364 29840
rect 10348 29800 10388 29840
rect 15532 29800 15572 29840
rect 2860 29716 2900 29756
rect 13420 29716 13460 29756
rect 14860 29716 14900 29756
rect 17836 29716 17876 29756
rect 15724 29632 15764 29672
rect 4300 29548 4340 29588
rect 14860 29548 14900 29588
rect 3688 29464 3728 29504
rect 3770 29464 3810 29504
rect 3852 29464 3892 29504
rect 3934 29464 3974 29504
rect 4016 29464 4056 29504
rect 18808 29464 18848 29504
rect 18890 29464 18930 29504
rect 18972 29464 19012 29504
rect 19054 29464 19094 29504
rect 19136 29464 19176 29504
rect 13804 29380 13844 29420
rect 15916 29380 15956 29420
rect 11980 29212 12020 29252
rect 14956 29212 14996 29252
rect 21292 29128 21332 29168
rect 12268 29044 12308 29084
rect 13612 29044 13652 29084
rect 18028 29044 18068 29084
rect 4396 28876 4436 28916
rect 10540 28876 10580 28916
rect 5644 28792 5684 28832
rect 15820 28792 15860 28832
rect 4928 28708 4968 28748
rect 5010 28708 5050 28748
rect 5092 28708 5132 28748
rect 5174 28708 5214 28748
rect 5256 28708 5296 28748
rect 5740 28708 5780 28748
rect 20048 28708 20088 28748
rect 20130 28708 20170 28748
rect 20212 28708 20252 28748
rect 20294 28708 20334 28748
rect 20376 28708 20416 28748
rect 10348 28624 10388 28664
rect 6316 28540 6356 28580
rect 9196 28540 9236 28580
rect 1804 28372 1844 28412
rect 460 28288 500 28328
rect 1612 28120 1652 28160
rect 3688 27952 3728 27992
rect 3770 27952 3810 27992
rect 3852 27952 3892 27992
rect 3934 27952 3974 27992
rect 4016 27952 4056 27992
rect 7660 27952 7700 27992
rect 16588 27952 16628 27992
rect 18808 27952 18848 27992
rect 18890 27952 18930 27992
rect 18972 27952 19012 27992
rect 19054 27952 19094 27992
rect 19136 27952 19176 27992
rect 18508 27784 18548 27824
rect 10732 27532 10772 27572
rect 4780 27448 4820 27488
rect 5644 27448 5684 27488
rect 11788 27448 11828 27488
rect 4396 27364 4436 27404
rect 5932 27364 5972 27404
rect 12172 27364 12212 27404
rect 18604 27364 18644 27404
rect 21292 27280 21332 27320
rect 4928 27196 4968 27236
rect 5010 27196 5050 27236
rect 5092 27196 5132 27236
rect 5174 27196 5214 27236
rect 5256 27196 5296 27236
rect 20048 27196 20088 27236
rect 20130 27196 20170 27236
rect 20212 27196 20252 27236
rect 20294 27196 20334 27236
rect 20376 27196 20416 27236
rect 4396 27112 4436 27152
rect 15532 27112 15572 27152
rect 15724 27112 15764 27152
rect 4300 26860 4340 26900
rect 4300 26692 4340 26732
rect 17836 26608 17876 26648
rect 16108 26524 16148 26564
rect 3688 26440 3728 26480
rect 3770 26440 3810 26480
rect 3852 26440 3892 26480
rect 3934 26440 3974 26480
rect 4016 26440 4056 26480
rect 18808 26440 18848 26480
rect 18890 26440 18930 26480
rect 18972 26440 19012 26480
rect 19054 26440 19094 26480
rect 19136 26440 19176 26480
rect 9292 26272 9332 26312
rect 13996 26272 14036 26312
rect 18508 26272 18548 26312
rect 9484 26188 9524 26228
rect 10060 26188 10100 26228
rect 13804 26188 13844 26228
rect 9388 26104 9428 26144
rect 1996 26020 2036 26060
rect 12268 26020 12308 26060
rect 7180 25936 7220 25976
rect 7564 25852 7604 25892
rect 4204 25768 4244 25808
rect 4928 25684 4968 25724
rect 5010 25684 5050 25724
rect 5092 25684 5132 25724
rect 5174 25684 5214 25724
rect 5256 25684 5296 25724
rect 20048 25684 20088 25724
rect 20130 25684 20170 25724
rect 20212 25684 20252 25724
rect 20294 25684 20334 25724
rect 20376 25684 20416 25724
rect 5740 25600 5780 25640
rect 20524 25432 20564 25472
rect 2860 25348 2900 25388
rect 9388 25348 9428 25388
rect 19276 25348 19316 25388
rect 1900 25264 1940 25304
rect 9292 25264 9332 25304
rect 10060 25264 10100 25304
rect 7660 25180 7700 25220
rect 19276 25180 19316 25220
rect 19468 25180 19508 25220
rect 1324 25096 1364 25136
rect 3244 25096 3284 25136
rect 1804 25012 1844 25052
rect 11980 25012 12020 25052
rect 19468 25012 19508 25052
rect 3688 24928 3728 24968
rect 3770 24928 3810 24968
rect 3852 24928 3892 24968
rect 3934 24928 3974 24968
rect 4016 24928 4056 24968
rect 7084 24928 7124 24968
rect 11596 24928 11636 24968
rect 18808 24928 18848 24968
rect 18890 24928 18930 24968
rect 18972 24928 19012 24968
rect 19054 24928 19094 24968
rect 19136 24928 19176 24968
rect 4204 24844 4244 24884
rect 8620 24844 8660 24884
rect 18124 24760 18164 24800
rect 3244 24676 3284 24716
rect 18028 24676 18068 24716
rect 7948 24592 7988 24632
rect 15436 24592 15476 24632
rect 18124 24592 18164 24632
rect 6028 24508 6068 24548
rect 7468 24508 7508 24548
rect 17548 24424 17588 24464
rect 20524 24424 20564 24464
rect 12940 24340 12980 24380
rect 4928 24172 4968 24212
rect 5010 24172 5050 24212
rect 5092 24172 5132 24212
rect 5174 24172 5214 24212
rect 5256 24172 5296 24212
rect 20048 24172 20088 24212
rect 20130 24172 20170 24212
rect 20212 24172 20252 24212
rect 20294 24172 20334 24212
rect 20376 24172 20416 24212
rect 3532 24004 3572 24044
rect 16492 24004 16532 24044
rect 14860 23752 14900 23792
rect 18316 23752 18356 23792
rect 3532 23668 3572 23708
rect 18028 23584 18068 23624
rect 4396 23500 4436 23540
rect 3688 23416 3728 23456
rect 3770 23416 3810 23456
rect 3852 23416 3892 23456
rect 3934 23416 3974 23456
rect 4016 23416 4056 23456
rect 15916 23416 15956 23456
rect 18808 23416 18848 23456
rect 18890 23416 18930 23456
rect 18972 23416 19012 23456
rect 19054 23416 19094 23456
rect 19136 23416 19176 23456
rect 18124 23332 18164 23372
rect 2380 23248 2420 23288
rect 2188 23164 2228 23204
rect 2860 23164 2900 23204
rect 13804 23248 13844 23288
rect 16108 23248 16148 23288
rect 18604 23248 18644 23288
rect 3532 23164 3572 23204
rect 8620 23164 8660 23204
rect 9004 23164 9044 23204
rect 13420 23164 13460 23204
rect 3244 23080 3284 23120
rect 4204 23080 4244 23120
rect 6124 23080 6164 23120
rect 9196 23080 9236 23120
rect 10732 23080 10772 23120
rect 15052 23080 15092 23120
rect 2188 22996 2228 23036
rect 4780 22996 4820 23036
rect 2380 22912 2420 22952
rect 2860 22912 2900 22952
rect 7660 22912 7700 22952
rect 5740 22828 5780 22868
rect 4928 22660 4968 22700
rect 5010 22660 5050 22700
rect 5092 22660 5132 22700
rect 5174 22660 5214 22700
rect 5256 22660 5296 22700
rect 20048 22660 20088 22700
rect 20130 22660 20170 22700
rect 20212 22660 20252 22700
rect 20294 22660 20334 22700
rect 20376 22660 20416 22700
rect 17836 22576 17876 22616
rect 18508 22408 18548 22448
rect 4204 22324 4244 22364
rect 11404 22324 11444 22364
rect 3532 22240 3572 22280
rect 20908 22072 20948 22112
rect 3688 21904 3728 21944
rect 3770 21904 3810 21944
rect 3852 21904 3892 21944
rect 3934 21904 3974 21944
rect 4016 21904 4056 21944
rect 11404 21904 11444 21944
rect 18808 21904 18848 21944
rect 18890 21904 18930 21944
rect 18972 21904 19012 21944
rect 19054 21904 19094 21944
rect 19136 21904 19176 21944
rect 3532 21736 3572 21776
rect 4300 21736 4340 21776
rect 13612 21652 13652 21692
rect 14572 21652 14612 21692
rect 18412 21652 18452 21692
rect 460 21568 500 21608
rect 7180 21568 7220 21608
rect 7468 21568 7508 21608
rect 10828 21484 10868 21524
rect 18028 21484 18068 21524
rect 18508 21484 18548 21524
rect 21100 21400 21140 21440
rect 4928 21148 4968 21188
rect 5010 21148 5050 21188
rect 5092 21148 5132 21188
rect 5174 21148 5214 21188
rect 5256 21148 5296 21188
rect 20048 21148 20088 21188
rect 20130 21148 20170 21188
rect 20212 21148 20252 21188
rect 20294 21148 20334 21188
rect 20376 21148 20416 21188
rect 18508 21064 18548 21104
rect 15340 20896 15380 20936
rect 2188 20812 2228 20852
rect 4204 20812 4244 20852
rect 5740 20812 5780 20852
rect 8620 20812 8660 20852
rect 12748 20812 12788 20852
rect 5932 20644 5972 20684
rect 16108 20644 16148 20684
rect 3688 20392 3728 20432
rect 3770 20392 3810 20432
rect 3852 20392 3892 20432
rect 3934 20392 3974 20432
rect 4016 20392 4056 20432
rect 18808 20392 18848 20432
rect 18890 20392 18930 20432
rect 18972 20392 19012 20432
rect 19054 20392 19094 20432
rect 19136 20392 19176 20432
rect 11212 20308 11252 20348
rect 4780 20224 4820 20264
rect 7276 20140 7316 20180
rect 10924 20140 10964 20180
rect 13420 20140 13460 20180
rect 14572 20140 14612 20180
rect 15820 20140 15860 20180
rect 6796 20056 6836 20096
rect 15340 20056 15380 20096
rect 18604 20056 18644 20096
rect 7084 19972 7124 20012
rect 10348 19888 10388 19928
rect 17836 19888 17876 19928
rect 20620 19804 20660 19844
rect 4928 19636 4968 19676
rect 5010 19636 5050 19676
rect 5092 19636 5132 19676
rect 5174 19636 5214 19676
rect 5256 19636 5296 19676
rect 20048 19636 20088 19676
rect 20130 19636 20170 19676
rect 20212 19636 20252 19676
rect 20294 19636 20334 19676
rect 20376 19636 20416 19676
rect 21388 19468 21428 19508
rect 4396 19384 4436 19424
rect 18508 19300 18548 19340
rect 3688 18880 3728 18920
rect 3770 18880 3810 18920
rect 3852 18880 3892 18920
rect 3934 18880 3974 18920
rect 4016 18880 4056 18920
rect 18808 18880 18848 18920
rect 18890 18880 18930 18920
rect 18972 18880 19012 18920
rect 19054 18880 19094 18920
rect 19136 18880 19176 18920
rect 12844 18628 12884 18668
rect 6796 18544 6836 18584
rect 7852 18544 7892 18584
rect 20524 18544 20564 18584
rect 15340 18460 15380 18500
rect 2188 18376 2228 18416
rect 5452 18376 5492 18416
rect 3244 18292 3284 18332
rect 19756 18208 19796 18248
rect 4928 18124 4968 18164
rect 5010 18124 5050 18164
rect 5092 18124 5132 18164
rect 5174 18124 5214 18164
rect 5256 18124 5296 18164
rect 20048 18124 20088 18164
rect 20130 18124 20170 18164
rect 20212 18124 20252 18164
rect 20294 18124 20334 18164
rect 20376 18124 20416 18164
rect 19660 17956 19700 17996
rect 3148 17872 3188 17912
rect 4300 17788 4340 17828
rect 21004 17536 21044 17576
rect 2860 17452 2900 17492
rect 3688 17368 3728 17408
rect 3770 17368 3810 17408
rect 3852 17368 3892 17408
rect 3934 17368 3974 17408
rect 4016 17368 4056 17408
rect 18808 17368 18848 17408
rect 18890 17368 18930 17408
rect 18972 17368 19012 17408
rect 19054 17368 19094 17408
rect 19136 17368 19176 17408
rect 11308 17200 11348 17240
rect 5644 17116 5684 17156
rect 13516 17032 13556 17072
rect 4780 16948 4820 16988
rect 14380 16948 14420 16988
rect 4396 16864 4436 16904
rect 4928 16612 4968 16652
rect 5010 16612 5050 16652
rect 5092 16612 5132 16652
rect 5174 16612 5214 16652
rect 5256 16612 5296 16652
rect 20048 16612 20088 16652
rect 20130 16612 20170 16652
rect 20212 16612 20252 16652
rect 20294 16612 20334 16652
rect 20376 16612 20416 16652
rect 13036 16528 13076 16568
rect 3532 16444 3572 16484
rect 6988 16444 7028 16484
rect 15244 16444 15284 16484
rect 4780 16276 4820 16316
rect 18508 16276 18548 16316
rect 6796 16192 6836 16232
rect 11404 16192 11444 16232
rect 2380 16108 2420 16148
rect 3688 15856 3728 15896
rect 3770 15856 3810 15896
rect 3852 15856 3892 15896
rect 3934 15856 3974 15896
rect 4016 15856 4056 15896
rect 18808 15856 18848 15896
rect 18890 15856 18930 15896
rect 18972 15856 19012 15896
rect 19054 15856 19094 15896
rect 19136 15856 19176 15896
rect 9580 15772 9620 15812
rect 6796 15604 6836 15644
rect 18604 15436 18644 15476
rect 13228 15352 13268 15392
rect 20812 15268 20852 15308
rect 4928 15100 4968 15140
rect 5010 15100 5050 15140
rect 5092 15100 5132 15140
rect 5174 15100 5214 15140
rect 5256 15100 5296 15140
rect 20048 15100 20088 15140
rect 20130 15100 20170 15140
rect 20212 15100 20252 15140
rect 20294 15100 20334 15140
rect 20376 15100 20416 15140
rect 9100 15016 9140 15056
rect 16012 14932 16052 14972
rect 9580 14848 9620 14888
rect 4396 14764 4436 14804
rect 14092 14764 14132 14804
rect 13036 14680 13076 14720
rect 14284 14512 14324 14552
rect 3688 14344 3728 14384
rect 3770 14344 3810 14384
rect 3852 14344 3892 14384
rect 3934 14344 3974 14384
rect 4016 14344 4056 14384
rect 18808 14344 18848 14384
rect 18890 14344 18930 14384
rect 18972 14344 19012 14384
rect 19054 14344 19094 14384
rect 19136 14344 19176 14384
rect 6700 14260 6740 14300
rect 8236 14260 8276 14300
rect 2860 13924 2900 13964
rect 3244 13924 3284 13964
rect 11404 13924 11444 13964
rect 14668 13756 14708 13796
rect 8908 13672 8948 13712
rect 4928 13588 4968 13628
rect 5010 13588 5050 13628
rect 5092 13588 5132 13628
rect 5174 13588 5214 13628
rect 5256 13588 5296 13628
rect 20048 13588 20088 13628
rect 20130 13588 20170 13628
rect 20212 13588 20252 13628
rect 20294 13588 20334 13628
rect 20376 13588 20416 13628
rect 3244 13504 3284 13544
rect 11692 13420 11732 13460
rect 3532 13168 3572 13208
rect 13036 13084 13076 13124
rect 4204 13000 4244 13040
rect 18316 13000 18356 13040
rect 3688 12832 3728 12872
rect 3770 12832 3810 12872
rect 3852 12832 3892 12872
rect 3934 12832 3974 12872
rect 4016 12832 4056 12872
rect 18316 12832 18356 12872
rect 18808 12832 18848 12872
rect 18890 12832 18930 12872
rect 18972 12832 19012 12872
rect 19054 12832 19094 12872
rect 19136 12832 19176 12872
rect 4204 12664 4244 12704
rect 17356 12664 17396 12704
rect 2860 12412 2900 12452
rect 9580 12412 9620 12452
rect 12364 12412 12404 12452
rect 13900 12412 13940 12452
rect 3244 12328 3284 12368
rect 4928 12076 4968 12116
rect 5010 12076 5050 12116
rect 5092 12076 5132 12116
rect 5174 12076 5214 12116
rect 5256 12076 5296 12116
rect 20048 12076 20088 12116
rect 20130 12076 20170 12116
rect 20212 12076 20252 12116
rect 20294 12076 20334 12116
rect 20376 12076 20416 12116
rect 11884 11824 11924 11864
rect 13900 11740 13940 11780
rect 3532 11656 3572 11696
rect 3688 11320 3728 11360
rect 3770 11320 3810 11360
rect 3852 11320 3892 11360
rect 3934 11320 3974 11360
rect 4016 11320 4056 11360
rect 18808 11320 18848 11360
rect 18890 11320 18930 11360
rect 18972 11320 19012 11360
rect 19054 11320 19094 11360
rect 19136 11320 19176 11360
rect 3436 11152 3476 11192
rect 4300 11152 4340 11192
rect 11404 10984 11444 11024
rect 19756 10732 19796 10772
rect 4928 10564 4968 10604
rect 5010 10564 5050 10604
rect 5092 10564 5132 10604
rect 5174 10564 5214 10604
rect 5256 10564 5296 10604
rect 20048 10564 20088 10604
rect 20130 10564 20170 10604
rect 20212 10564 20252 10604
rect 20294 10564 20334 10604
rect 20376 10564 20416 10604
rect 19276 10144 19316 10184
rect 2188 10060 2228 10100
rect 3436 10060 3476 10100
rect 11404 10060 11444 10100
rect 14572 10060 14612 10100
rect 3688 9808 3728 9848
rect 3770 9808 3810 9848
rect 3852 9808 3892 9848
rect 3934 9808 3974 9848
rect 4016 9808 4056 9848
rect 18808 9808 18848 9848
rect 18890 9808 18930 9848
rect 18972 9808 19012 9848
rect 19054 9808 19094 9848
rect 19136 9808 19176 9848
rect 15628 9724 15668 9764
rect 19564 9640 19604 9680
rect 13516 9556 13556 9596
rect 3436 9472 3476 9512
rect 10636 9304 10676 9344
rect 4928 9052 4968 9092
rect 5010 9052 5050 9092
rect 5092 9052 5132 9092
rect 5174 9052 5214 9092
rect 5256 9052 5296 9092
rect 20048 9052 20088 9092
rect 20130 9052 20170 9092
rect 20212 9052 20252 9092
rect 20294 9052 20334 9092
rect 20376 9052 20416 9092
rect 21292 8632 21332 8672
rect 13516 8548 13556 8588
rect 2476 8464 2516 8504
rect 3688 8296 3728 8336
rect 3770 8296 3810 8336
rect 3852 8296 3892 8336
rect 3934 8296 3974 8336
rect 4016 8296 4056 8336
rect 18808 8296 18848 8336
rect 18890 8296 18930 8336
rect 18972 8296 19012 8336
rect 19054 8296 19094 8336
rect 19136 8296 19176 8336
rect 16300 8128 16340 8168
rect 11020 7960 11060 8000
rect 4928 7540 4968 7580
rect 5010 7540 5050 7580
rect 5092 7540 5132 7580
rect 5174 7540 5214 7580
rect 5256 7540 5296 7580
rect 20048 7540 20088 7580
rect 20130 7540 20170 7580
rect 20212 7540 20252 7580
rect 20294 7540 20334 7580
rect 20376 7540 20416 7580
rect 6220 7120 6260 7160
rect 16780 7120 16820 7160
rect 3688 6784 3728 6824
rect 3770 6784 3810 6824
rect 3852 6784 3892 6824
rect 3934 6784 3974 6824
rect 4016 6784 4056 6824
rect 18808 6784 18848 6824
rect 18890 6784 18930 6824
rect 18972 6784 19012 6824
rect 19054 6784 19094 6824
rect 19136 6784 19176 6824
rect 19660 6280 19700 6320
rect 4928 6028 4968 6068
rect 5010 6028 5050 6068
rect 5092 6028 5132 6068
rect 5174 6028 5214 6068
rect 5256 6028 5296 6068
rect 12556 6028 12596 6068
rect 20048 6028 20088 6068
rect 20130 6028 20170 6068
rect 20212 6028 20252 6068
rect 20294 6028 20334 6068
rect 20376 6028 20416 6068
rect 10156 5944 10196 5984
rect 7372 5692 7412 5732
rect 4684 5608 4724 5648
rect 5548 5524 5588 5564
rect 20716 5440 20756 5480
rect 3688 5272 3728 5312
rect 3770 5272 3810 5312
rect 3852 5272 3892 5312
rect 3934 5272 3974 5312
rect 4016 5272 4056 5312
rect 18808 5272 18848 5312
rect 18890 5272 18930 5312
rect 18972 5272 19012 5312
rect 19054 5272 19094 5312
rect 19136 5272 19176 5312
rect 4928 4516 4968 4556
rect 5010 4516 5050 4556
rect 5092 4516 5132 4556
rect 5174 4516 5214 4556
rect 5256 4516 5296 4556
rect 20048 4516 20088 4556
rect 20130 4516 20170 4556
rect 20212 4516 20252 4556
rect 20294 4516 20334 4556
rect 20376 4516 20416 4556
rect 8716 4264 8756 4304
rect 17452 4180 17492 4220
rect 14476 4096 14516 4136
rect 3688 3760 3728 3800
rect 3770 3760 3810 3800
rect 3852 3760 3892 3800
rect 3934 3760 3974 3800
rect 4016 3760 4056 3800
rect 12652 3760 12692 3800
rect 18808 3760 18848 3800
rect 18890 3760 18930 3800
rect 18972 3760 19012 3800
rect 19054 3760 19094 3800
rect 19136 3760 19176 3800
rect 10252 3508 10292 3548
rect 1996 3424 2036 3464
rect 17644 3424 17684 3464
rect 12076 3340 12116 3380
rect 9964 3172 10004 3212
rect 9868 3088 9908 3128
rect 4928 3004 4968 3044
rect 5010 3004 5050 3044
rect 5092 3004 5132 3044
rect 5174 3004 5214 3044
rect 5256 3004 5296 3044
rect 20048 3004 20088 3044
rect 20130 3004 20170 3044
rect 20212 3004 20252 3044
rect 20294 3004 20334 3044
rect 20376 3004 20416 3044
rect 4588 2836 4628 2876
rect 8428 2836 8468 2876
rect 15148 2836 15188 2876
rect 4492 2752 4532 2792
rect 17740 2752 17780 2792
rect 10828 2668 10868 2708
rect 2092 2584 2132 2624
rect 2764 2584 2804 2624
rect 10348 2584 10388 2624
rect 14764 2584 14804 2624
rect 8044 2416 8084 2456
rect 13612 2416 13652 2456
rect 12460 2332 12500 2372
rect 3688 2248 3728 2288
rect 3770 2248 3810 2288
rect 3852 2248 3892 2288
rect 3934 2248 3974 2288
rect 4016 2248 4056 2288
rect 18808 2248 18848 2288
rect 18890 2248 18930 2288
rect 18972 2248 19012 2288
rect 19054 2248 19094 2288
rect 19136 2248 19176 2288
rect 2956 2164 2996 2204
rect 2284 2080 2324 2120
rect 2572 2080 2612 2120
rect 3340 2080 3380 2120
rect 5836 2080 5876 2120
rect 10732 1996 10772 2036
rect 9292 1912 9332 1952
rect 11500 1912 11540 1952
rect 13420 1912 13460 1952
rect 18220 1912 18260 1952
rect 6508 1744 6548 1784
rect 4928 1492 4968 1532
rect 5010 1492 5050 1532
rect 5092 1492 5132 1532
rect 5174 1492 5214 1532
rect 5256 1492 5296 1532
rect 20048 1492 20088 1532
rect 20130 1492 20170 1532
rect 20212 1492 20252 1532
rect 20294 1492 20334 1532
rect 20376 1492 20416 1532
rect 7756 1408 7796 1448
rect 8140 1408 8180 1448
rect 8332 1408 8372 1448
rect 8524 1408 8564 1448
rect 13132 1408 13172 1448
rect 17164 1408 17204 1448
rect 19468 1408 19508 1448
rect 13708 1324 13748 1364
rect 8812 1240 8852 1280
rect 16396 1240 16436 1280
rect 6604 1156 6644 1196
rect 9676 1156 9716 1196
rect 21484 1156 21524 1196
rect 16972 988 17012 1028
rect 14188 820 14228 860
rect 19852 568 19892 608
rect 16204 484 16244 524
rect 13324 400 13364 440
rect 6892 316 6932 356
rect 9772 316 9812 356
rect 6412 232 6452 272
rect 2668 148 2708 188
rect 19372 148 19412 188
<< metal5 >>
rect 1324 94856 1364 94865
rect 1324 83540 1364 94816
rect 1804 94856 1844 94865
rect 1708 89816 1748 89825
rect 1132 83500 1364 83540
rect 1420 89648 1460 89657
rect 748 75956 788 75965
rect 364 75536 404 75545
rect 364 73856 404 75496
rect 364 73807 404 73816
rect 748 70748 788 75916
rect 1132 74276 1172 83500
rect 1324 82340 1364 82349
rect 1132 74227 1172 74236
rect 1228 76040 1268 76049
rect 748 70699 788 70708
rect 1228 68984 1268 76000
rect 1324 74192 1364 82300
rect 1420 82088 1460 89608
rect 1516 85532 1556 85541
rect 1516 83432 1556 85492
rect 1516 83383 1556 83392
rect 1612 84104 1652 84113
rect 1420 82039 1460 82048
rect 1516 80576 1556 80585
rect 1516 76796 1556 80536
rect 1516 76747 1556 76756
rect 1324 74143 1364 74152
rect 1420 74360 1460 74369
rect 1228 68935 1268 68944
rect 1420 67640 1460 74320
rect 1420 67591 1460 67600
rect 1420 66968 1460 66977
rect 1420 62936 1460 66928
rect 1420 62887 1460 62896
rect 1516 63356 1556 63365
rect 1516 59324 1556 63316
rect 1516 59275 1556 59284
rect 1612 54284 1652 84064
rect 1708 79904 1748 89776
rect 1708 79855 1748 79864
rect 1708 72092 1748 72101
rect 1708 69152 1748 72052
rect 1804 71168 1844 94816
rect 2092 94856 2132 94865
rect 1996 89396 2036 89405
rect 1804 71119 1844 71128
rect 1900 84104 1940 84113
rect 1708 69103 1748 69112
rect 1804 67220 1844 67229
rect 1708 66296 1748 66305
rect 1708 64448 1748 66256
rect 1708 64399 1748 64408
rect 1708 63356 1748 63365
rect 1708 54956 1748 63316
rect 1708 54907 1748 54916
rect 1612 54235 1652 54244
rect 1804 51848 1844 67180
rect 1900 60248 1940 84064
rect 1996 71420 2036 89356
rect 1996 71371 2036 71380
rect 1996 70076 2036 70085
rect 1996 66884 2036 70036
rect 2092 67136 2132 94816
rect 2476 94856 2516 94865
rect 2380 90320 2420 90329
rect 2380 83684 2420 90280
rect 2380 83635 2420 83644
rect 2284 77552 2324 77561
rect 2188 73436 2228 73445
rect 2188 71756 2228 73396
rect 2188 71707 2228 71716
rect 2092 67087 2132 67096
rect 2188 67472 2228 67481
rect 1996 66835 2036 66844
rect 2092 65540 2132 65549
rect 1900 60199 1940 60208
rect 1996 63860 2036 63869
rect 1996 53300 2036 63820
rect 2092 59408 2132 65500
rect 2188 64196 2228 67432
rect 2188 64147 2228 64156
rect 2092 59359 2132 59368
rect 2188 64028 2228 64037
rect 2188 53528 2228 63988
rect 2188 53479 2228 53488
rect 1996 53260 2132 53300
rect 1804 51799 1844 51808
rect 1996 44792 2036 44801
rect 1516 40760 1556 40769
rect 1516 33116 1556 40720
rect 1516 33067 1556 33076
rect 1612 35300 1652 35309
rect 1612 32864 1652 35260
rect 1612 32815 1652 32824
rect 1708 34292 1748 34301
rect 1612 32024 1652 32033
rect 1324 29840 1364 29849
rect 460 28328 500 28337
rect 460 21608 500 28288
rect 1324 25136 1364 29800
rect 1612 28160 1652 31984
rect 1708 30260 1748 34252
rect 1996 33536 2036 44752
rect 2092 35300 2132 53260
rect 2092 35251 2132 35260
rect 2188 43280 2228 43289
rect 1996 33487 2036 33496
rect 2188 33144 2228 43240
rect 2284 39584 2324 77512
rect 2380 69992 2420 70001
rect 2380 64028 2420 69952
rect 2380 63979 2420 63988
rect 2476 60416 2516 94816
rect 3340 94856 3380 94865
rect 3052 90908 3092 90917
rect 2860 89060 2900 89069
rect 2668 86372 2708 86381
rect 2572 80576 2612 80585
rect 2572 77048 2612 80536
rect 2572 76999 2612 77008
rect 2668 77468 2708 86332
rect 2764 84272 2804 84281
rect 2764 83432 2804 84232
rect 2860 84020 2900 89020
rect 2860 83971 2900 83980
rect 2764 83383 2804 83392
rect 2668 76376 2708 77428
rect 2668 76327 2708 76336
rect 2764 79820 2804 79829
rect 2572 73100 2612 73109
rect 2572 65288 2612 73060
rect 2572 65239 2612 65248
rect 2668 66296 2708 66305
rect 2668 63944 2708 66256
rect 2668 63895 2708 63904
rect 2572 63692 2612 63701
rect 2572 61508 2612 63652
rect 2572 61459 2612 61468
rect 2668 63356 2708 63365
rect 2476 60367 2516 60376
rect 2668 53360 2708 63316
rect 2668 53311 2708 53320
rect 2668 53108 2708 53117
rect 2572 51008 2612 51017
rect 2284 39535 2324 39544
rect 2380 50840 2420 50849
rect 2284 36812 2324 36821
rect 2284 33620 2324 36772
rect 2284 33571 2324 33580
rect 2092 33104 2228 33144
rect 2284 33368 2324 33377
rect 2092 33032 2132 33104
rect 1900 32992 2132 33032
rect 2188 33032 2228 33041
rect 1708 30211 1748 30220
rect 1804 32948 1844 32957
rect 1612 28111 1652 28120
rect 1804 28412 1844 32908
rect 1324 25087 1364 25096
rect 1804 25052 1844 28372
rect 1900 25304 1940 32992
rect 2092 32864 2132 32873
rect 1900 25255 1940 25264
rect 1996 26060 2036 26069
rect 1804 25003 1844 25012
rect 460 21559 500 21568
rect 1996 3464 2036 26020
rect 1996 3415 2036 3424
rect 2092 2624 2132 32824
rect 2188 23204 2228 32992
rect 2188 23155 2228 23164
rect 2188 23036 2228 23045
rect 2188 20852 2228 22996
rect 2188 20803 2228 20812
rect 2188 18416 2228 18425
rect 2188 10100 2228 18376
rect 2188 10051 2228 10060
rect 2092 2575 2132 2584
rect 2284 2120 2324 33328
rect 2380 23288 2420 50800
rect 2380 23239 2420 23248
rect 2476 48068 2516 48077
rect 2380 22952 2420 22961
rect 2380 16148 2420 22912
rect 2380 16099 2420 16108
rect 2476 8504 2516 48028
rect 2572 43280 2612 50968
rect 2668 44792 2708 53068
rect 2668 44743 2708 44752
rect 2572 43240 2708 43280
rect 2476 8455 2516 8464
rect 2572 43112 2612 43121
rect 2284 2071 2324 2080
rect 2572 2120 2612 43072
rect 2572 2071 2612 2080
rect 2668 188 2708 43240
rect 2764 2624 2804 79780
rect 2956 73520 2996 73529
rect 2956 71756 2996 73480
rect 2956 71707 2996 71716
rect 2860 69236 2900 69245
rect 2860 66432 2900 69196
rect 2860 66392 2996 66432
rect 2860 65960 2900 65969
rect 2860 64784 2900 65920
rect 2860 64735 2900 64744
rect 2956 64616 2996 66392
rect 2956 64567 2996 64576
rect 2956 63944 2996 63953
rect 2956 63696 2996 63904
rect 2860 63656 2996 63696
rect 2860 63356 2900 63656
rect 3052 63380 3092 90868
rect 3148 89396 3188 89405
rect 3148 81416 3188 89356
rect 3244 85112 3284 85121
rect 3244 83600 3284 85072
rect 3244 83551 3284 83560
rect 3148 81367 3188 81376
rect 3244 79736 3284 79745
rect 3244 76796 3284 79696
rect 3244 76747 3284 76756
rect 3244 72512 3284 72521
rect 3148 72428 3188 72437
rect 3148 65456 3188 72388
rect 3148 65407 3188 65416
rect 3244 65120 3284 72472
rect 3244 65071 3284 65080
rect 3244 63776 3284 63785
rect 2860 63307 2900 63316
rect 2956 63340 3092 63380
rect 3148 63524 3188 63533
rect 2956 63020 2996 63340
rect 2956 62971 2996 62980
rect 3052 63272 3092 63281
rect 3052 58232 3092 63232
rect 3148 62180 3188 63484
rect 3148 62131 3188 62140
rect 3052 58183 3092 58192
rect 3244 54788 3284 63736
rect 3244 54739 3284 54748
rect 3244 53864 3284 53873
rect 2860 53360 2900 53369
rect 2860 53108 2900 53320
rect 2860 53059 2900 53068
rect 3148 41348 3188 41357
rect 2956 39668 2996 39677
rect 2956 35048 2996 39628
rect 2956 34999 2996 35008
rect 3052 38996 3092 39005
rect 2956 33704 2996 33713
rect 2860 33536 2900 33545
rect 2860 33032 2900 33496
rect 2860 32983 2900 32992
rect 2956 31940 2996 33664
rect 3052 33368 3092 38956
rect 3148 34460 3188 41308
rect 3148 34411 3188 34420
rect 3052 33319 3092 33328
rect 3148 33284 3188 33293
rect 2956 31891 2996 31900
rect 3052 33200 3092 33209
rect 2860 29756 2900 29765
rect 2860 25388 2900 29716
rect 2860 25339 2900 25348
rect 2860 23204 2900 23213
rect 2860 22952 2900 23164
rect 3052 23060 3092 33160
rect 2860 22903 2900 22912
rect 2956 23020 3092 23060
rect 2860 17492 2900 17501
rect 2860 13964 2900 17452
rect 2860 12452 2900 13924
rect 2860 12403 2900 12412
rect 2764 2575 2804 2584
rect 2956 2204 2996 23020
rect 3148 17912 3188 33244
rect 3244 32276 3284 53824
rect 3340 46724 3380 94816
rect 3652 94520 4092 96768
rect 4892 95276 5332 96768
rect 4892 95236 4928 95276
rect 4968 95236 5010 95276
rect 5050 95236 5092 95276
rect 5132 95236 5174 95276
rect 5214 95236 5256 95276
rect 5296 95236 5332 95276
rect 3652 94480 3688 94520
rect 3728 94480 3770 94520
rect 3810 94480 3852 94520
rect 3892 94480 3934 94520
rect 3974 94480 4016 94520
rect 4056 94480 4092 94520
rect 3652 93008 4092 94480
rect 3652 92968 3688 93008
rect 3728 92968 3770 93008
rect 3810 92968 3852 93008
rect 3892 92968 3934 93008
rect 3974 92968 4016 93008
rect 4056 92968 4092 93008
rect 3652 91496 4092 92968
rect 3652 91456 3688 91496
rect 3728 91456 3770 91496
rect 3810 91456 3852 91496
rect 3892 91456 3934 91496
rect 3974 91456 4016 91496
rect 4056 91456 4092 91496
rect 3532 89984 3572 89993
rect 3532 87296 3572 89944
rect 3436 84356 3476 84365
rect 3436 83096 3476 84316
rect 3436 83047 3476 83056
rect 3532 82760 3572 87256
rect 3532 82711 3572 82720
rect 3652 89984 4092 91456
rect 4396 94856 4436 94865
rect 3652 89944 3688 89984
rect 3728 89944 3770 89984
rect 3810 89944 3852 89984
rect 3892 89944 3934 89984
rect 3974 89944 4016 89984
rect 4056 89944 4092 89984
rect 3652 88472 4092 89944
rect 3652 88432 3688 88472
rect 3728 88432 3770 88472
rect 3810 88432 3852 88472
rect 3892 88432 3934 88472
rect 3974 88432 4016 88472
rect 4056 88432 4092 88472
rect 3652 86960 4092 88432
rect 3652 86920 3688 86960
rect 3728 86920 3770 86960
rect 3810 86920 3852 86960
rect 3892 86920 3934 86960
rect 3974 86920 4016 86960
rect 4056 86920 4092 86960
rect 3652 85448 4092 86920
rect 3652 85408 3688 85448
rect 3728 85408 3770 85448
rect 3810 85408 3852 85448
rect 3892 85408 3934 85448
rect 3974 85408 4016 85448
rect 4056 85408 4092 85448
rect 3652 83936 4092 85408
rect 3652 83896 3688 83936
rect 3728 83896 3770 83936
rect 3810 83896 3852 83936
rect 3892 83896 3934 83936
rect 3974 83896 4016 83936
rect 4056 83896 4092 83936
rect 3532 82592 3572 82601
rect 3532 82004 3572 82552
rect 3532 81955 3572 81964
rect 3652 82424 4092 83896
rect 3652 82384 3688 82424
rect 3728 82384 3770 82424
rect 3810 82384 3852 82424
rect 3892 82384 3934 82424
rect 3974 82384 4016 82424
rect 4056 82384 4092 82424
rect 3652 80912 4092 82384
rect 3652 80872 3688 80912
rect 3728 80872 3770 80912
rect 3810 80872 3852 80912
rect 3892 80872 3934 80912
rect 3974 80872 4016 80912
rect 4056 80872 4092 80912
rect 3532 79652 3572 79661
rect 3436 78980 3476 78989
rect 3436 78224 3476 78940
rect 3436 77048 3476 78184
rect 3532 77216 3572 79612
rect 3532 77167 3572 77176
rect 3652 79400 4092 80872
rect 3652 79360 3688 79400
rect 3728 79360 3770 79400
rect 3810 79360 3852 79400
rect 3892 79360 3934 79400
rect 3974 79360 4016 79400
rect 4056 79360 4092 79400
rect 3652 77888 4092 79360
rect 3652 77848 3688 77888
rect 3728 77848 3770 77888
rect 3810 77848 3852 77888
rect 3892 77848 3934 77888
rect 3974 77848 4016 77888
rect 4056 77848 4092 77888
rect 3436 77008 3572 77048
rect 3532 76628 3572 77008
rect 3532 75872 3572 76588
rect 3532 74360 3572 75832
rect 3532 74311 3572 74320
rect 3652 76376 4092 77848
rect 3652 76336 3688 76376
rect 3728 76336 3770 76376
rect 3810 76336 3852 76376
rect 3892 76336 3934 76376
rect 3974 76336 4016 76376
rect 4056 76336 4092 76376
rect 3652 74864 4092 76336
rect 3652 74824 3688 74864
rect 3728 74824 3770 74864
rect 3810 74824 3852 74864
rect 3892 74824 3934 74864
rect 3974 74824 4016 74864
rect 4056 74824 4092 74864
rect 3436 74192 3476 74201
rect 3436 64616 3476 74152
rect 3652 73352 4092 74824
rect 3652 73312 3688 73352
rect 3728 73312 3770 73352
rect 3810 73312 3852 73352
rect 3892 73312 3934 73352
rect 3974 73312 4016 73352
rect 4056 73312 4092 73352
rect 3532 72260 3572 72269
rect 3532 71672 3572 72220
rect 3532 71623 3572 71632
rect 3652 71840 4092 73312
rect 4204 90152 4244 90161
rect 4204 72512 4244 90112
rect 4300 83012 4340 83021
rect 4300 77888 4340 82972
rect 4300 77839 4340 77848
rect 4204 72463 4244 72472
rect 4300 73604 4340 73613
rect 3652 71800 3688 71840
rect 3728 71800 3770 71840
rect 3810 71800 3852 71840
rect 3892 71800 3934 71840
rect 3974 71800 4016 71840
rect 4056 71800 4092 71840
rect 3652 70328 4092 71800
rect 3652 70288 3688 70328
rect 3728 70288 3770 70328
rect 3810 70288 3852 70328
rect 3892 70288 3934 70328
rect 3974 70288 4016 70328
rect 4056 70288 4092 70328
rect 3532 69236 3572 69245
rect 3532 67640 3572 69196
rect 3532 67591 3572 67600
rect 3652 68816 4092 70288
rect 3652 68776 3688 68816
rect 3728 68776 3770 68816
rect 3810 68776 3852 68816
rect 3892 68776 3934 68816
rect 3974 68776 4016 68816
rect 4056 68776 4092 68816
rect 3532 67472 3572 67481
rect 3532 67052 3572 67432
rect 3532 67003 3572 67012
rect 3652 67304 4092 68776
rect 3652 67264 3688 67304
rect 3728 67264 3770 67304
rect 3810 67264 3852 67304
rect 3892 67264 3934 67304
rect 3974 67264 4016 67304
rect 4056 67264 4092 67304
rect 3436 64567 3476 64576
rect 3532 66212 3572 66221
rect 3532 64700 3572 66172
rect 3436 63524 3476 63533
rect 3436 61004 3476 63484
rect 3532 63272 3572 64660
rect 3532 63223 3572 63232
rect 3652 65792 4092 67264
rect 3652 65752 3688 65792
rect 3728 65752 3770 65792
rect 3810 65752 3852 65792
rect 3892 65752 3934 65792
rect 3974 65752 4016 65792
rect 4056 65752 4092 65792
rect 3652 64280 4092 65752
rect 4204 72344 4244 72353
rect 4204 65624 4244 72304
rect 4300 70664 4340 73564
rect 4300 70615 4340 70624
rect 4204 65575 4244 65584
rect 4300 69908 4340 69917
rect 4300 66212 4340 69868
rect 3652 64240 3688 64280
rect 3728 64240 3770 64280
rect 3810 64240 3852 64280
rect 3892 64240 3934 64280
rect 3974 64240 4016 64280
rect 4056 64240 4092 64280
rect 3652 62768 4092 64240
rect 3652 62728 3688 62768
rect 3728 62728 3770 62768
rect 3810 62728 3852 62768
rect 3892 62728 3934 62768
rect 3974 62728 4016 62768
rect 4056 62728 4092 62768
rect 4204 63944 4244 63953
rect 4204 62784 4244 63904
rect 4300 63608 4340 66172
rect 4300 63559 4340 63568
rect 4204 62744 4340 62784
rect 3532 61676 3572 61685
rect 3532 61088 3572 61636
rect 3532 61039 3572 61048
rect 3652 61256 4092 62728
rect 3652 61216 3688 61256
rect 3728 61216 3770 61256
rect 3810 61216 3852 61256
rect 3892 61216 3934 61256
rect 3974 61216 4016 61256
rect 4056 61216 4092 61256
rect 3436 60955 3476 60964
rect 3340 46675 3380 46684
rect 3436 60164 3476 60173
rect 3244 32227 3284 32236
rect 3340 37484 3380 37493
rect 3244 32108 3284 32117
rect 3244 25136 3284 32068
rect 3244 25087 3284 25096
rect 3244 24716 3284 24725
rect 3244 23120 3284 24676
rect 3244 23071 3284 23080
rect 3148 17863 3188 17872
rect 3244 18332 3284 18341
rect 3244 13964 3284 18292
rect 3244 13915 3284 13924
rect 3244 13544 3284 13553
rect 3244 12368 3284 13504
rect 3244 12319 3284 12328
rect 2956 2155 2996 2164
rect 3340 2120 3380 37444
rect 3436 11192 3476 60124
rect 3652 59744 4092 61216
rect 4204 62348 4244 62357
rect 4204 60920 4244 62308
rect 4300 61592 4340 62744
rect 4300 61543 4340 61552
rect 4204 60871 4244 60880
rect 3652 59704 3688 59744
rect 3728 59704 3770 59744
rect 3810 59704 3852 59744
rect 3892 59704 3934 59744
rect 3974 59704 4016 59744
rect 4056 59704 4092 59744
rect 3652 58232 4092 59704
rect 3652 58192 3688 58232
rect 3728 58192 3770 58232
rect 3810 58192 3852 58232
rect 3892 58192 3934 58232
rect 3974 58192 4016 58232
rect 4056 58192 4092 58232
rect 3652 56720 4092 58192
rect 4204 60752 4244 60761
rect 4204 57812 4244 60712
rect 4204 57763 4244 57772
rect 3652 56680 3688 56720
rect 3728 56680 3770 56720
rect 3810 56680 3852 56720
rect 3892 56680 3934 56720
rect 3974 56680 4016 56720
rect 4056 56680 4092 56720
rect 3652 55208 4092 56680
rect 3652 55168 3688 55208
rect 3728 55168 3770 55208
rect 3810 55168 3852 55208
rect 3892 55168 3934 55208
rect 3974 55168 4016 55208
rect 4056 55168 4092 55208
rect 3652 53696 4092 55168
rect 3652 53656 3688 53696
rect 3728 53656 3770 53696
rect 3810 53656 3852 53696
rect 3892 53656 3934 53696
rect 3974 53656 4016 53696
rect 4056 53656 4092 53696
rect 3652 52184 4092 53656
rect 3652 52144 3688 52184
rect 3728 52144 3770 52184
rect 3810 52144 3852 52184
rect 3892 52144 3934 52184
rect 3974 52144 4016 52184
rect 4056 52144 4092 52184
rect 3652 50672 4092 52144
rect 3652 50632 3688 50672
rect 3728 50632 3770 50672
rect 3810 50632 3852 50672
rect 3892 50632 3934 50672
rect 3974 50632 4016 50672
rect 4056 50632 4092 50672
rect 3652 49160 4092 50632
rect 3652 49120 3688 49160
rect 3728 49120 3770 49160
rect 3810 49120 3852 49160
rect 3892 49120 3934 49160
rect 3974 49120 4016 49160
rect 4056 49120 4092 49160
rect 3652 47648 4092 49120
rect 3652 47608 3688 47648
rect 3728 47608 3770 47648
rect 3810 47608 3852 47648
rect 3892 47608 3934 47648
rect 3974 47608 4016 47648
rect 4056 47608 4092 47648
rect 3652 46136 4092 47608
rect 3652 46096 3688 46136
rect 3728 46096 3770 46136
rect 3810 46096 3852 46136
rect 3892 46096 3934 46136
rect 3974 46096 4016 46136
rect 4056 46096 4092 46136
rect 3652 44624 4092 46096
rect 3652 44584 3688 44624
rect 3728 44584 3770 44624
rect 3810 44584 3852 44624
rect 3892 44584 3934 44624
rect 3974 44584 4016 44624
rect 4056 44584 4092 44624
rect 3652 43112 4092 44584
rect 3652 43072 3688 43112
rect 3728 43072 3770 43112
rect 3810 43072 3852 43112
rect 3892 43072 3934 43112
rect 3974 43072 4016 43112
rect 4056 43072 4092 43112
rect 3652 41600 4092 43072
rect 3652 41560 3688 41600
rect 3728 41560 3770 41600
rect 3810 41560 3852 41600
rect 3892 41560 3934 41600
rect 3974 41560 4016 41600
rect 4056 41560 4092 41600
rect 3532 40256 3572 40265
rect 3532 36728 3572 40216
rect 3532 36679 3572 36688
rect 3652 40088 4092 41560
rect 3652 40048 3688 40088
rect 3728 40048 3770 40088
rect 3810 40048 3852 40088
rect 3892 40048 3934 40088
rect 3974 40048 4016 40088
rect 4056 40048 4092 40088
rect 3652 38576 4092 40048
rect 3652 38536 3688 38576
rect 3728 38536 3770 38576
rect 3810 38536 3852 38576
rect 3892 38536 3934 38576
rect 3974 38536 4016 38576
rect 4056 38536 4092 38576
rect 3652 37064 4092 38536
rect 3652 37024 3688 37064
rect 3728 37024 3770 37064
rect 3810 37024 3852 37064
rect 3892 37024 3934 37064
rect 3974 37024 4016 37064
rect 4056 37024 4092 37064
rect 3532 36560 3572 36569
rect 3532 35972 3572 36520
rect 3532 24044 3572 35932
rect 3532 23995 3572 24004
rect 3652 35552 4092 37024
rect 3652 35512 3688 35552
rect 3728 35512 3770 35552
rect 3810 35512 3852 35552
rect 3892 35512 3934 35552
rect 3974 35512 4016 35552
rect 4056 35512 4092 35552
rect 3652 34040 4092 35512
rect 3652 34000 3688 34040
rect 3728 34000 3770 34040
rect 3810 34000 3852 34040
rect 3892 34000 3934 34040
rect 3974 34000 4016 34040
rect 4056 34000 4092 34040
rect 3652 32528 4092 34000
rect 3652 32488 3688 32528
rect 3728 32488 3770 32528
rect 3810 32488 3852 32528
rect 3892 32488 3934 32528
rect 3974 32488 4016 32528
rect 4056 32488 4092 32528
rect 3652 31016 4092 32488
rect 3652 30976 3688 31016
rect 3728 30976 3770 31016
rect 3810 30976 3852 31016
rect 3892 30976 3934 31016
rect 3974 30976 4016 31016
rect 4056 30976 4092 31016
rect 3652 29504 4092 30976
rect 3652 29464 3688 29504
rect 3728 29464 3770 29504
rect 3810 29464 3852 29504
rect 3892 29464 3934 29504
rect 3974 29464 4016 29504
rect 4056 29464 4092 29504
rect 3652 27992 4092 29464
rect 3652 27952 3688 27992
rect 3728 27952 3770 27992
rect 3810 27952 3852 27992
rect 3892 27952 3934 27992
rect 3974 27952 4016 27992
rect 4056 27952 4092 27992
rect 3652 26480 4092 27952
rect 3652 26440 3688 26480
rect 3728 26440 3770 26480
rect 3810 26440 3852 26480
rect 3892 26440 3934 26480
rect 3974 26440 4016 26480
rect 4056 26440 4092 26480
rect 3652 24968 4092 26440
rect 4204 48572 4244 48581
rect 4204 25808 4244 48532
rect 4300 44036 4340 44045
rect 4300 43112 4340 43996
rect 4300 43063 4340 43072
rect 4300 41600 4340 41609
rect 4300 39500 4340 41560
rect 4300 39451 4340 39460
rect 4300 39332 4340 39341
rect 4300 36140 4340 39292
rect 4396 38156 4436 94816
rect 4684 94856 4724 94865
rect 4492 94184 4532 94193
rect 4492 46724 4532 94144
rect 4492 46675 4532 46684
rect 4588 89648 4628 89657
rect 4492 45380 4532 45389
rect 4492 43616 4532 45340
rect 4492 43567 4532 43576
rect 4396 38107 4436 38116
rect 4492 41852 4532 41861
rect 4300 36091 4340 36100
rect 4300 34544 4340 34553
rect 4300 33284 4340 34504
rect 4300 33235 4340 33244
rect 4396 33200 4436 33209
rect 4396 32948 4436 33160
rect 4396 32899 4436 32908
rect 4396 32780 4436 32789
rect 4300 32276 4340 32285
rect 4300 29588 4340 32236
rect 4396 31100 4436 32740
rect 4396 31051 4436 31060
rect 4300 29539 4340 29548
rect 4396 30848 4436 30857
rect 4396 29040 4436 30808
rect 4300 29000 4436 29040
rect 4300 26900 4340 29000
rect 4396 28916 4436 28925
rect 4396 27404 4436 28876
rect 4396 27355 4436 27364
rect 4300 26851 4340 26860
rect 4396 27152 4436 27161
rect 4204 25759 4244 25768
rect 4300 26732 4340 26741
rect 3652 24928 3688 24968
rect 3728 24928 3770 24968
rect 3810 24928 3852 24968
rect 3892 24928 3934 24968
rect 3974 24928 4016 24968
rect 4056 24928 4092 24968
rect 3532 23708 3572 23717
rect 3532 23204 3572 23668
rect 3532 23155 3572 23164
rect 3652 23456 4092 24928
rect 3652 23416 3688 23456
rect 3728 23416 3770 23456
rect 3810 23416 3852 23456
rect 3892 23416 3934 23456
rect 3974 23416 4016 23456
rect 4056 23416 4092 23456
rect 3532 22280 3572 22289
rect 3532 21776 3572 22240
rect 3532 21727 3572 21736
rect 3652 21944 4092 23416
rect 4204 24884 4244 24893
rect 4204 23120 4244 24844
rect 4204 23071 4244 23080
rect 3652 21904 3688 21944
rect 3728 21904 3770 21944
rect 3810 21904 3852 21944
rect 3892 21904 3934 21944
rect 3974 21904 4016 21944
rect 4056 21904 4092 21944
rect 3652 20432 4092 21904
rect 4204 22364 4244 22373
rect 4204 20852 4244 22324
rect 4300 21776 4340 26692
rect 4396 23540 4436 27112
rect 4396 23491 4436 23500
rect 4300 21727 4340 21736
rect 4204 20803 4244 20812
rect 3652 20392 3688 20432
rect 3728 20392 3770 20432
rect 3810 20392 3852 20432
rect 3892 20392 3934 20432
rect 3974 20392 4016 20432
rect 4056 20392 4092 20432
rect 3652 18920 4092 20392
rect 3652 18880 3688 18920
rect 3728 18880 3770 18920
rect 3810 18880 3852 18920
rect 3892 18880 3934 18920
rect 3974 18880 4016 18920
rect 4056 18880 4092 18920
rect 3652 17408 4092 18880
rect 4396 19424 4436 19433
rect 3652 17368 3688 17408
rect 3728 17368 3770 17408
rect 3810 17368 3852 17408
rect 3892 17368 3934 17408
rect 3974 17368 4016 17408
rect 4056 17368 4092 17408
rect 3532 16484 3572 16493
rect 3532 13208 3572 16444
rect 3532 13159 3572 13168
rect 3652 15896 4092 17368
rect 3652 15856 3688 15896
rect 3728 15856 3770 15896
rect 3810 15856 3852 15896
rect 3892 15856 3934 15896
rect 3974 15856 4016 15896
rect 4056 15856 4092 15896
rect 3652 14384 4092 15856
rect 3652 14344 3688 14384
rect 3728 14344 3770 14384
rect 3810 14344 3852 14384
rect 3892 14344 3934 14384
rect 3974 14344 4016 14384
rect 4056 14344 4092 14384
rect 3652 12872 4092 14344
rect 4300 17828 4340 17837
rect 3652 12832 3688 12872
rect 3728 12832 3770 12872
rect 3810 12832 3852 12872
rect 3892 12832 3934 12872
rect 3974 12832 4016 12872
rect 4056 12832 4092 12872
rect 3436 11143 3476 11152
rect 3532 11696 3572 11705
rect 3436 10100 3476 10109
rect 3532 10100 3572 11656
rect 3476 10060 3572 10100
rect 3652 11360 4092 12832
rect 4204 13040 4244 13049
rect 4204 12704 4244 13000
rect 4204 12655 4244 12664
rect 3652 11320 3688 11360
rect 3728 11320 3770 11360
rect 3810 11320 3852 11360
rect 3892 11320 3934 11360
rect 3974 11320 4016 11360
rect 4056 11320 4092 11360
rect 3436 9512 3476 10060
rect 3436 9463 3476 9472
rect 3652 9848 4092 11320
rect 4300 11192 4340 17788
rect 4396 16904 4436 19384
rect 4396 14804 4436 16864
rect 4396 14755 4436 14764
rect 4300 11143 4340 11152
rect 3652 9808 3688 9848
rect 3728 9808 3770 9848
rect 3810 9808 3852 9848
rect 3892 9808 3934 9848
rect 3974 9808 4016 9848
rect 4056 9808 4092 9848
rect 3340 2071 3380 2080
rect 3652 8336 4092 9808
rect 3652 8296 3688 8336
rect 3728 8296 3770 8336
rect 3810 8296 3852 8336
rect 3892 8296 3934 8336
rect 3974 8296 4016 8336
rect 4056 8296 4092 8336
rect 3652 6824 4092 8296
rect 3652 6784 3688 6824
rect 3728 6784 3770 6824
rect 3810 6784 3852 6824
rect 3892 6784 3934 6824
rect 3974 6784 4016 6824
rect 4056 6784 4092 6824
rect 3652 5312 4092 6784
rect 3652 5272 3688 5312
rect 3728 5272 3770 5312
rect 3810 5272 3852 5312
rect 3892 5272 3934 5312
rect 3974 5272 4016 5312
rect 4056 5272 4092 5312
rect 3652 3800 4092 5272
rect 3652 3760 3688 3800
rect 3728 3760 3770 3800
rect 3810 3760 3852 3800
rect 3892 3760 3934 3800
rect 3974 3760 4016 3800
rect 4056 3760 4092 3800
rect 3652 2288 4092 3760
rect 4492 2792 4532 41812
rect 4588 41432 4628 89608
rect 4588 41383 4628 41392
rect 4588 40508 4628 40517
rect 4588 2876 4628 40468
rect 4684 5648 4724 94816
rect 4892 93764 5332 95236
rect 9100 96620 9140 96629
rect 6316 94856 6356 94865
rect 4892 93724 4928 93764
rect 4968 93724 5010 93764
rect 5050 93724 5092 93764
rect 5132 93724 5174 93764
rect 5214 93724 5256 93764
rect 5296 93724 5332 93764
rect 4892 92252 5332 93724
rect 5548 94184 5588 94193
rect 5548 93620 5588 94144
rect 5740 94184 5780 94193
rect 5548 93580 5684 93620
rect 4892 92212 4928 92252
rect 4968 92212 5010 92252
rect 5050 92212 5092 92252
rect 5132 92212 5174 92252
rect 5214 92212 5256 92252
rect 5296 92212 5332 92252
rect 4892 90740 5332 92212
rect 4892 90700 4928 90740
rect 4968 90700 5010 90740
rect 5050 90700 5092 90740
rect 5132 90700 5174 90740
rect 5214 90700 5256 90740
rect 5296 90700 5332 90740
rect 4892 89228 5332 90700
rect 4892 89188 4928 89228
rect 4968 89188 5010 89228
rect 5050 89188 5092 89228
rect 5132 89188 5174 89228
rect 5214 89188 5256 89228
rect 5296 89188 5332 89228
rect 4892 87716 5332 89188
rect 4892 87676 4928 87716
rect 4968 87676 5010 87716
rect 5050 87676 5092 87716
rect 5132 87676 5174 87716
rect 5214 87676 5256 87716
rect 5296 87676 5332 87716
rect 4892 86204 5332 87676
rect 4892 86164 4928 86204
rect 4968 86164 5010 86204
rect 5050 86164 5092 86204
rect 5132 86164 5174 86204
rect 5214 86164 5256 86204
rect 5296 86164 5332 86204
rect 4780 85112 4820 85121
rect 4780 83012 4820 85072
rect 4780 82963 4820 82972
rect 4892 84692 5332 86164
rect 5452 87128 5492 87137
rect 5452 85112 5492 87088
rect 5452 85063 5492 85072
rect 4892 84652 4928 84692
rect 4968 84652 5010 84692
rect 5050 84652 5092 84692
rect 5132 84652 5174 84692
rect 5214 84652 5256 84692
rect 5296 84652 5332 84692
rect 4892 83180 5332 84652
rect 5548 84524 5588 84533
rect 4892 83140 4928 83180
rect 4968 83140 5010 83180
rect 5050 83140 5092 83180
rect 5132 83140 5174 83180
rect 5214 83140 5256 83180
rect 5296 83140 5332 83180
rect 4780 82844 4820 82853
rect 4780 75452 4820 82804
rect 4780 75403 4820 75412
rect 4892 81668 5332 83140
rect 4892 81628 4928 81668
rect 4968 81628 5010 81668
rect 5050 81628 5092 81668
rect 5132 81628 5174 81668
rect 5214 81628 5256 81668
rect 5296 81628 5332 81668
rect 4892 80156 5332 81628
rect 4892 80116 4928 80156
rect 4968 80116 5010 80156
rect 5050 80116 5092 80156
rect 5132 80116 5174 80156
rect 5214 80116 5256 80156
rect 5296 80116 5332 80156
rect 4892 78644 5332 80116
rect 5452 83516 5492 83525
rect 5452 78980 5492 83476
rect 5548 81500 5588 84484
rect 5548 81451 5588 81460
rect 5452 78931 5492 78940
rect 5548 80324 5588 80333
rect 5548 78812 5588 80284
rect 5548 78763 5588 78772
rect 4892 78604 4928 78644
rect 4968 78604 5010 78644
rect 5050 78604 5092 78644
rect 5132 78604 5174 78644
rect 5214 78604 5256 78644
rect 5296 78604 5332 78644
rect 4892 77132 5332 78604
rect 4892 77092 4928 77132
rect 4968 77092 5010 77132
rect 5050 77092 5092 77132
rect 5132 77092 5174 77132
rect 5214 77092 5256 77132
rect 5296 77092 5332 77132
rect 4892 75620 5332 77092
rect 5548 78056 5588 78065
rect 5548 76964 5588 78016
rect 4892 75580 4928 75620
rect 4968 75580 5010 75620
rect 5050 75580 5092 75620
rect 5132 75580 5174 75620
rect 5214 75580 5256 75620
rect 5296 75580 5332 75620
rect 4780 75284 4820 75293
rect 4780 74192 4820 75244
rect 4780 70916 4820 74152
rect 4780 70867 4820 70876
rect 4892 74108 5332 75580
rect 5452 76376 5492 76385
rect 5452 74780 5492 76336
rect 5452 74731 5492 74740
rect 4892 74068 4928 74108
rect 4968 74068 5010 74108
rect 5050 74068 5092 74108
rect 5132 74068 5174 74108
rect 5214 74068 5256 74108
rect 5296 74068 5332 74108
rect 4892 72596 5332 74068
rect 4892 72556 4928 72596
rect 4968 72556 5010 72596
rect 5050 72556 5092 72596
rect 5132 72556 5174 72596
rect 5214 72556 5256 72596
rect 5296 72556 5332 72596
rect 4892 71084 5332 72556
rect 5452 74612 5492 74621
rect 5452 74360 5492 74572
rect 5452 72008 5492 74320
rect 5452 71959 5492 71968
rect 4892 71044 4928 71084
rect 4968 71044 5010 71084
rect 5050 71044 5092 71084
rect 5132 71044 5174 71084
rect 5214 71044 5256 71084
rect 5296 71044 5332 71084
rect 4780 70748 4820 70757
rect 4780 68480 4820 70708
rect 4780 68431 4820 68440
rect 4892 69572 5332 71044
rect 5548 70580 5588 76924
rect 5644 71588 5684 93580
rect 5644 71539 5684 71548
rect 5548 70531 5588 70540
rect 5644 70496 5684 70505
rect 4892 69532 4928 69572
rect 4968 69532 5010 69572
rect 5050 69532 5092 69572
rect 5132 69532 5174 69572
rect 5214 69532 5256 69572
rect 5296 69532 5332 69572
rect 4892 68060 5332 69532
rect 5548 69740 5588 69749
rect 4892 68020 4928 68060
rect 4968 68020 5010 68060
rect 5050 68020 5092 68060
rect 5132 68020 5174 68060
rect 5214 68020 5256 68060
rect 5296 68020 5332 68060
rect 4780 67892 4820 67901
rect 4780 64112 4820 67852
rect 4780 64063 4820 64072
rect 4892 66548 5332 68020
rect 4892 66508 4928 66548
rect 4968 66508 5010 66548
rect 5050 66508 5092 66548
rect 5132 66508 5174 66548
rect 5214 66508 5256 66548
rect 5296 66508 5332 66548
rect 4892 65036 5332 66508
rect 4892 64996 4928 65036
rect 4968 64996 5010 65036
rect 5050 64996 5092 65036
rect 5132 64996 5174 65036
rect 5214 64996 5256 65036
rect 5296 64996 5332 65036
rect 4780 63944 4820 63953
rect 4780 63104 4820 63904
rect 4780 63055 4820 63064
rect 4892 63524 5332 64996
rect 4892 63484 4928 63524
rect 4968 63484 5010 63524
rect 5050 63484 5092 63524
rect 5132 63484 5174 63524
rect 5214 63484 5256 63524
rect 5296 63484 5332 63524
rect 4780 62180 4820 62189
rect 4780 54788 4820 62140
rect 4780 54739 4820 54748
rect 4892 62012 5332 63484
rect 4892 61972 4928 62012
rect 4968 61972 5010 62012
rect 5050 61972 5092 62012
rect 5132 61972 5174 62012
rect 5214 61972 5256 62012
rect 5296 61972 5332 62012
rect 4892 60500 5332 61972
rect 4892 60460 4928 60500
rect 4968 60460 5010 60500
rect 5050 60460 5092 60500
rect 5132 60460 5174 60500
rect 5214 60460 5256 60500
rect 5296 60460 5332 60500
rect 4892 58988 5332 60460
rect 4892 58948 4928 58988
rect 4968 58948 5010 58988
rect 5050 58948 5092 58988
rect 5132 58948 5174 58988
rect 5214 58948 5256 58988
rect 5296 58948 5332 58988
rect 4892 57476 5332 58948
rect 4892 57436 4928 57476
rect 4968 57436 5010 57476
rect 5050 57436 5092 57476
rect 5132 57436 5174 57476
rect 5214 57436 5256 57476
rect 5296 57436 5332 57476
rect 4892 55964 5332 57436
rect 4892 55924 4928 55964
rect 4968 55924 5010 55964
rect 5050 55924 5092 55964
rect 5132 55924 5174 55964
rect 5214 55924 5256 55964
rect 5296 55924 5332 55964
rect 4892 54452 5332 55924
rect 4892 54412 4928 54452
rect 4968 54412 5010 54452
rect 5050 54412 5092 54452
rect 5132 54412 5174 54452
rect 5214 54412 5256 54452
rect 5296 54412 5332 54452
rect 4892 52940 5332 54412
rect 4892 52900 4928 52940
rect 4968 52900 5010 52940
rect 5050 52900 5092 52940
rect 5132 52900 5174 52940
rect 5214 52900 5256 52940
rect 5296 52900 5332 52940
rect 4892 51428 5332 52900
rect 4892 51388 4928 51428
rect 4968 51388 5010 51428
rect 5050 51388 5092 51428
rect 5132 51388 5174 51428
rect 5214 51388 5256 51428
rect 5296 51388 5332 51428
rect 4892 49916 5332 51388
rect 4892 49876 4928 49916
rect 4968 49876 5010 49916
rect 5050 49876 5092 49916
rect 5132 49876 5174 49916
rect 5214 49876 5256 49916
rect 5296 49876 5332 49916
rect 4892 48404 5332 49876
rect 4892 48364 4928 48404
rect 4968 48364 5010 48404
rect 5050 48364 5092 48404
rect 5132 48364 5174 48404
rect 5214 48364 5256 48404
rect 5296 48364 5332 48404
rect 4892 46892 5332 48364
rect 4892 46852 4928 46892
rect 4968 46852 5010 46892
rect 5050 46852 5092 46892
rect 5132 46852 5174 46892
rect 5214 46852 5256 46892
rect 5296 46852 5332 46892
rect 4892 45380 5332 46852
rect 4892 45340 4928 45380
rect 4968 45340 5010 45380
rect 5050 45340 5092 45380
rect 5132 45340 5174 45380
rect 5214 45340 5256 45380
rect 5296 45340 5332 45380
rect 4892 43868 5332 45340
rect 4892 43828 4928 43868
rect 4968 43828 5010 43868
rect 5050 43828 5092 43868
rect 5132 43828 5174 43868
rect 5214 43828 5256 43868
rect 5296 43828 5332 43868
rect 4780 43700 4820 43709
rect 4780 41852 4820 43660
rect 4780 41803 4820 41812
rect 4892 42356 5332 43828
rect 4892 42316 4928 42356
rect 4968 42316 5010 42356
rect 5050 42316 5092 42356
rect 5132 42316 5174 42356
rect 5214 42316 5256 42356
rect 5296 42316 5332 42356
rect 4780 41348 4820 41357
rect 4780 34544 4820 41308
rect 4780 34495 4820 34504
rect 4892 40844 5332 42316
rect 4892 40804 4928 40844
rect 4968 40804 5010 40844
rect 5050 40804 5092 40844
rect 5132 40804 5174 40844
rect 5214 40804 5256 40844
rect 5296 40804 5332 40844
rect 4892 39332 5332 40804
rect 4892 39292 4928 39332
rect 4968 39292 5010 39332
rect 5050 39292 5092 39332
rect 5132 39292 5174 39332
rect 5214 39292 5256 39332
rect 5296 39292 5332 39332
rect 4892 37820 5332 39292
rect 4892 37780 4928 37820
rect 4968 37780 5010 37820
rect 5050 37780 5092 37820
rect 5132 37780 5174 37820
rect 5214 37780 5256 37820
rect 5296 37780 5332 37820
rect 4892 36308 5332 37780
rect 4892 36268 4928 36308
rect 4968 36268 5010 36308
rect 5050 36268 5092 36308
rect 5132 36268 5174 36308
rect 5214 36268 5256 36308
rect 5296 36268 5332 36308
rect 4892 34796 5332 36268
rect 4892 34756 4928 34796
rect 4968 34756 5010 34796
rect 5050 34756 5092 34796
rect 5132 34756 5174 34796
rect 5214 34756 5256 34796
rect 5296 34756 5332 34796
rect 4892 33284 5332 34756
rect 4892 33244 4928 33284
rect 4968 33244 5010 33284
rect 5050 33244 5092 33284
rect 5132 33244 5174 33284
rect 5214 33244 5256 33284
rect 5296 33244 5332 33284
rect 4780 31772 4820 31781
rect 4780 27488 4820 31732
rect 4780 27439 4820 27448
rect 4892 31772 5332 33244
rect 4892 31732 4928 31772
rect 4968 31732 5010 31772
rect 5050 31732 5092 31772
rect 5132 31732 5174 31772
rect 5214 31732 5256 31772
rect 5296 31732 5332 31772
rect 4892 30260 5332 31732
rect 4892 30220 4928 30260
rect 4968 30220 5010 30260
rect 5050 30220 5092 30260
rect 5132 30220 5174 30260
rect 5214 30220 5256 30260
rect 5296 30220 5332 30260
rect 4892 28748 5332 30220
rect 4892 28708 4928 28748
rect 4968 28708 5010 28748
rect 5050 28708 5092 28748
rect 5132 28708 5174 28748
rect 5214 28708 5256 28748
rect 5296 28708 5332 28748
rect 4892 27236 5332 28708
rect 4892 27196 4928 27236
rect 4968 27196 5010 27236
rect 5050 27196 5092 27236
rect 5132 27196 5174 27236
rect 5214 27196 5256 27236
rect 5296 27196 5332 27236
rect 4892 25724 5332 27196
rect 4892 25684 4928 25724
rect 4968 25684 5010 25724
rect 5050 25684 5092 25724
rect 5132 25684 5174 25724
rect 5214 25684 5256 25724
rect 5296 25684 5332 25724
rect 4892 24212 5332 25684
rect 4892 24172 4928 24212
rect 4968 24172 5010 24212
rect 5050 24172 5092 24212
rect 5132 24172 5174 24212
rect 5214 24172 5256 24212
rect 5296 24172 5332 24212
rect 4780 23036 4820 23045
rect 4780 20264 4820 22996
rect 4780 20215 4820 20224
rect 4892 22700 5332 24172
rect 4892 22660 4928 22700
rect 4968 22660 5010 22700
rect 5050 22660 5092 22700
rect 5132 22660 5174 22700
rect 5214 22660 5256 22700
rect 5296 22660 5332 22700
rect 4892 21188 5332 22660
rect 4892 21148 4928 21188
rect 4968 21148 5010 21188
rect 5050 21148 5092 21188
rect 5132 21148 5174 21188
rect 5214 21148 5256 21188
rect 5296 21148 5332 21188
rect 4892 19676 5332 21148
rect 4892 19636 4928 19676
rect 4968 19636 5010 19676
rect 5050 19636 5092 19676
rect 5132 19636 5174 19676
rect 5214 19636 5256 19676
rect 5296 19636 5332 19676
rect 4892 18164 5332 19636
rect 5452 68396 5492 68405
rect 5452 18416 5492 68356
rect 5548 66968 5588 69700
rect 5644 68312 5684 70456
rect 5644 68263 5684 68272
rect 5548 66919 5588 66928
rect 5452 18367 5492 18376
rect 5548 64784 5588 64793
rect 4892 18124 4928 18164
rect 4968 18124 5010 18164
rect 5050 18124 5092 18164
rect 5132 18124 5174 18164
rect 5214 18124 5256 18164
rect 5296 18124 5332 18164
rect 4780 16988 4820 16997
rect 4780 16316 4820 16948
rect 4780 16267 4820 16276
rect 4892 16652 5332 18124
rect 4892 16612 4928 16652
rect 4968 16612 5010 16652
rect 5050 16612 5092 16652
rect 5132 16612 5174 16652
rect 5214 16612 5256 16652
rect 5296 16612 5332 16652
rect 4684 5599 4724 5608
rect 4892 15140 5332 16612
rect 4892 15100 4928 15140
rect 4968 15100 5010 15140
rect 5050 15100 5092 15140
rect 5132 15100 5174 15140
rect 5214 15100 5256 15140
rect 5296 15100 5332 15140
rect 4892 13628 5332 15100
rect 4892 13588 4928 13628
rect 4968 13588 5010 13628
rect 5050 13588 5092 13628
rect 5132 13588 5174 13628
rect 5214 13588 5256 13628
rect 5296 13588 5332 13628
rect 4892 12116 5332 13588
rect 4892 12076 4928 12116
rect 4968 12076 5010 12116
rect 5050 12076 5092 12116
rect 5132 12076 5174 12116
rect 5214 12076 5256 12116
rect 5296 12076 5332 12116
rect 4892 10604 5332 12076
rect 4892 10564 4928 10604
rect 4968 10564 5010 10604
rect 5050 10564 5092 10604
rect 5132 10564 5174 10604
rect 5214 10564 5256 10604
rect 5296 10564 5332 10604
rect 4892 9092 5332 10564
rect 4892 9052 4928 9092
rect 4968 9052 5010 9092
rect 5050 9052 5092 9092
rect 5132 9052 5174 9092
rect 5214 9052 5256 9092
rect 5296 9052 5332 9092
rect 4892 7580 5332 9052
rect 4892 7540 4928 7580
rect 4968 7540 5010 7580
rect 5050 7540 5092 7580
rect 5132 7540 5174 7580
rect 5214 7540 5256 7580
rect 5296 7540 5332 7580
rect 4892 6068 5332 7540
rect 4892 6028 4928 6068
rect 4968 6028 5010 6068
rect 5050 6028 5092 6068
rect 5132 6028 5174 6068
rect 5214 6028 5256 6068
rect 5296 6028 5332 6068
rect 4588 2827 4628 2836
rect 4892 4556 5332 6028
rect 5548 5564 5588 64744
rect 5644 63692 5684 63701
rect 5644 63356 5684 63652
rect 5644 63307 5684 63316
rect 5644 58820 5684 58829
rect 5644 56972 5684 58780
rect 5644 56923 5684 56932
rect 5644 46052 5684 46061
rect 5644 45212 5684 46012
rect 5644 45163 5684 45172
rect 5644 44372 5684 44381
rect 5644 43700 5684 44332
rect 5644 43651 5684 43660
rect 5740 40340 5780 94144
rect 6124 94184 6164 94193
rect 5932 93932 5972 93941
rect 5836 84524 5876 84533
rect 5836 83264 5876 84484
rect 5836 83215 5876 83224
rect 5836 82256 5876 82265
rect 5836 81164 5876 82216
rect 5836 81115 5876 81124
rect 5836 70076 5876 70085
rect 5836 69320 5876 70036
rect 5836 69271 5876 69280
rect 5740 40291 5780 40300
rect 5836 64616 5876 64625
rect 5644 38492 5684 38501
rect 5644 28832 5684 38452
rect 5740 38156 5780 38165
rect 5740 31184 5780 38116
rect 5740 31135 5780 31144
rect 5644 28783 5684 28792
rect 5740 28748 5780 28757
rect 5644 27488 5684 27497
rect 5644 17156 5684 27448
rect 5740 25640 5780 28708
rect 5740 25591 5780 25600
rect 5740 22868 5780 22877
rect 5740 20852 5780 22828
rect 5740 20803 5780 20812
rect 5644 17107 5684 17116
rect 5548 5515 5588 5524
rect 4892 4516 4928 4556
rect 4968 4516 5010 4556
rect 5050 4516 5092 4556
rect 5132 4516 5174 4556
rect 5214 4516 5256 4556
rect 5296 4516 5332 4556
rect 4892 3044 5332 4516
rect 4892 3004 4928 3044
rect 4968 3004 5010 3044
rect 5050 3004 5092 3044
rect 5132 3004 5174 3044
rect 5214 3004 5256 3044
rect 5296 3004 5332 3044
rect 4492 2743 4532 2752
rect 3652 2248 3688 2288
rect 3728 2248 3770 2288
rect 3810 2248 3852 2288
rect 3892 2248 3934 2288
rect 3974 2248 4016 2288
rect 4056 2248 4092 2288
rect 2668 139 2708 148
rect 3652 0 4092 2248
rect 4892 1532 5332 3004
rect 5836 2120 5876 64576
rect 5932 54368 5972 93892
rect 6028 81500 6068 81509
rect 6028 79232 6068 81460
rect 6028 79183 6068 79192
rect 6028 76292 6068 76301
rect 6028 73520 6068 76252
rect 6028 73471 6068 73480
rect 6028 66968 6068 66977
rect 6028 61508 6068 66928
rect 6124 64784 6164 94144
rect 6220 74528 6260 74537
rect 6220 70580 6260 74488
rect 6220 70531 6260 70540
rect 6124 64735 6164 64744
rect 6028 61459 6068 61468
rect 6124 64532 6164 64541
rect 6124 63356 6164 64492
rect 6124 60752 6164 63316
rect 6124 60703 6164 60712
rect 5932 54319 5972 54328
rect 6220 55376 6260 55385
rect 6124 48740 6164 48749
rect 5932 44372 5972 44381
rect 5932 43280 5972 44332
rect 5932 43112 5972 43240
rect 5932 43063 5972 43072
rect 5932 42944 5972 42953
rect 5932 36980 5972 42904
rect 5932 34628 5972 36940
rect 5932 34579 5972 34588
rect 6028 41180 6068 41189
rect 5932 27404 5972 27413
rect 5932 20684 5972 27364
rect 6028 24548 6068 41140
rect 6124 41012 6164 48700
rect 6124 40963 6164 40972
rect 6028 24499 6068 24508
rect 6124 40844 6164 40853
rect 6124 40424 6164 40804
rect 6124 30344 6164 40384
rect 6124 23120 6164 30304
rect 6124 23071 6164 23080
rect 5932 20635 5972 20644
rect 6220 7160 6260 55336
rect 6316 28580 6356 94816
rect 6700 94856 6740 94865
rect 6604 92336 6644 92345
rect 6412 81080 6452 81089
rect 6412 58316 6452 81040
rect 6508 79316 6548 79325
rect 6508 70748 6548 79276
rect 6508 70699 6548 70708
rect 6412 58267 6452 58276
rect 6508 68480 6548 68489
rect 6316 28531 6356 28540
rect 6412 56384 6452 56393
rect 6220 7111 6260 7120
rect 5836 2071 5876 2080
rect 4892 1492 4928 1532
rect 4968 1492 5010 1532
rect 5050 1492 5092 1532
rect 5132 1492 5174 1532
rect 5214 1492 5256 1532
rect 5296 1492 5332 1532
rect 4892 0 5332 1492
rect 6412 272 6452 56344
rect 6508 44624 6548 68440
rect 6508 44575 6548 44584
rect 6508 44120 6548 44129
rect 6508 43448 6548 44080
rect 6508 43399 6548 43408
rect 6508 39668 6548 39677
rect 6508 1784 6548 39628
rect 6508 1735 6548 1744
rect 6604 1196 6644 92296
rect 6700 40172 6740 94816
rect 7084 94856 7124 94865
rect 6892 93848 6932 93857
rect 6796 75200 6836 75209
rect 6796 67640 6836 75160
rect 6796 67591 6836 67600
rect 6796 67472 6836 67481
rect 6796 63692 6836 67432
rect 6796 63643 6836 63652
rect 6700 40123 6740 40132
rect 6796 50420 6836 50429
rect 6700 39500 6740 39509
rect 6700 37704 6740 39460
rect 6796 38072 6836 50380
rect 6796 38023 6836 38032
rect 6700 37664 6836 37704
rect 6700 34544 6740 34553
rect 6700 14300 6740 34504
rect 6796 31940 6836 37664
rect 6796 31891 6836 31900
rect 6796 20096 6836 20105
rect 6796 18584 6836 20056
rect 6796 16232 6836 18544
rect 6796 15644 6836 16192
rect 6796 15595 6836 15604
rect 6700 14251 6740 14260
rect 6604 1147 6644 1156
rect 6892 356 6932 93808
rect 6988 75956 7028 75965
rect 6988 75116 7028 75916
rect 6988 75067 7028 75076
rect 6988 72764 7028 72773
rect 6988 70832 7028 72724
rect 6988 66128 7028 70792
rect 6988 66079 7028 66088
rect 7084 64112 7124 94816
rect 8812 94688 8852 94697
rect 8044 94184 8084 94193
rect 7756 93932 7796 93941
rect 7084 64063 7124 64072
rect 7180 93596 7220 93605
rect 7084 62852 7124 62861
rect 7084 61508 7124 62812
rect 7084 61459 7124 61468
rect 6988 59744 7028 59753
rect 6988 16484 7028 59704
rect 7084 40172 7124 40181
rect 7084 37148 7124 40132
rect 7084 37099 7124 37108
rect 7180 35468 7220 93556
rect 7660 88724 7700 88733
rect 7468 81836 7508 81845
rect 7372 80408 7412 80417
rect 7180 35419 7220 35428
rect 7276 75032 7316 75041
rect 7084 34712 7124 34721
rect 7084 32864 7124 34672
rect 7084 32815 7124 32824
rect 7180 25976 7220 25985
rect 7084 24968 7124 24977
rect 7084 20012 7124 24928
rect 7180 21608 7220 25936
rect 7180 21559 7220 21568
rect 7276 20180 7316 74992
rect 7372 70580 7412 80368
rect 7372 70531 7412 70540
rect 7372 67640 7412 67649
rect 7372 60752 7412 67600
rect 7372 60703 7412 60712
rect 7276 20131 7316 20140
rect 7372 48488 7412 48497
rect 7084 19963 7124 19972
rect 6988 16435 7028 16444
rect 7372 5732 7412 48448
rect 7468 34376 7508 81796
rect 7468 34327 7508 34336
rect 7564 69404 7604 69413
rect 7468 30176 7508 30185
rect 7468 24548 7508 30136
rect 7564 25892 7604 69364
rect 7660 68396 7700 88684
rect 7660 68347 7700 68356
rect 7660 38996 7700 39005
rect 7660 32696 7700 38956
rect 7660 27992 7700 32656
rect 7660 27943 7700 27952
rect 7564 25843 7604 25852
rect 7468 21608 7508 24508
rect 7660 25220 7700 25229
rect 7660 22952 7700 25180
rect 7660 22903 7700 22912
rect 7468 21559 7508 21568
rect 7372 5683 7412 5692
rect 7756 1448 7796 93892
rect 7948 86540 7988 86549
rect 7852 85112 7892 85121
rect 7852 18584 7892 85072
rect 7948 83264 7988 86500
rect 7948 83215 7988 83224
rect 7948 79904 7988 79913
rect 7948 77720 7988 79864
rect 7948 77671 7988 77680
rect 7948 76124 7988 76133
rect 7948 71504 7988 76084
rect 7948 71455 7988 71464
rect 7948 70244 7988 70253
rect 7948 68228 7988 70204
rect 7948 63104 7988 68188
rect 7948 63055 7988 63064
rect 7948 54284 7988 54293
rect 7948 30596 7988 54244
rect 8044 38828 8084 94144
rect 8332 91832 8372 91841
rect 8044 38779 8084 38788
rect 8140 91160 8180 91169
rect 7948 30547 7988 30556
rect 8044 32360 8084 32369
rect 7948 30092 7988 30101
rect 7948 24632 7988 30052
rect 7948 24583 7988 24592
rect 7852 18535 7892 18544
rect 8044 2456 8084 32320
rect 8044 2407 8084 2416
rect 7756 1399 7796 1408
rect 8140 1448 8180 91120
rect 8236 87968 8276 87977
rect 8236 73268 8276 87928
rect 8236 73219 8276 73228
rect 8236 68228 8276 68237
rect 8236 14300 8276 68188
rect 8236 14251 8276 14260
rect 8140 1399 8180 1408
rect 8332 1448 8372 91792
rect 8524 91160 8564 91169
rect 8428 84776 8468 84785
rect 8428 2876 8468 84736
rect 8428 2827 8468 2836
rect 8332 1399 8372 1408
rect 8524 1448 8564 91120
rect 8716 87548 8756 87557
rect 8620 76292 8660 76301
rect 8620 39920 8660 76252
rect 8716 60164 8756 87508
rect 8716 60115 8756 60124
rect 8812 56132 8852 94648
rect 9004 83432 9044 83441
rect 8908 78140 8948 78149
rect 8908 74612 8948 78100
rect 8908 74563 8948 74572
rect 9004 73520 9044 83392
rect 9004 73471 9044 73480
rect 8908 70580 8948 70589
rect 8908 64700 8948 70540
rect 8908 64651 8948 64660
rect 9004 68312 9044 68321
rect 8908 64028 8948 64037
rect 8908 63524 8948 63988
rect 8908 63475 8948 63484
rect 9004 63380 9044 68272
rect 8812 56083 8852 56092
rect 8908 63340 9044 63380
rect 8812 52856 8852 52865
rect 8620 39871 8660 39880
rect 8716 48404 8756 48413
rect 8620 32444 8660 32453
rect 8620 30428 8660 32404
rect 8620 24884 8660 30388
rect 8620 24835 8660 24844
rect 8620 23204 8660 23213
rect 8620 20852 8660 23164
rect 8620 20803 8660 20812
rect 8716 4304 8756 48364
rect 8716 4255 8756 4264
rect 8524 1399 8564 1408
rect 8812 1280 8852 52816
rect 8908 13712 8948 63340
rect 9004 62096 9044 62105
rect 9004 23204 9044 62056
rect 9004 23155 9044 23164
rect 9100 15056 9140 96580
rect 12556 95948 12596 95957
rect 9484 95696 9524 95705
rect 9388 94688 9428 94697
rect 9292 92672 9332 92681
rect 9196 77384 9236 77393
rect 9196 73352 9236 77344
rect 9196 73303 9236 73312
rect 9196 64952 9236 64961
rect 9196 62432 9236 64912
rect 9196 62383 9236 62392
rect 9196 62012 9236 62021
rect 9196 47984 9236 61972
rect 9292 56552 9332 92632
rect 9292 56503 9332 56512
rect 9388 48656 9428 94648
rect 9388 48607 9428 48616
rect 9196 47935 9236 47944
rect 9196 47228 9236 47237
rect 9196 45716 9236 47188
rect 9196 40928 9236 45676
rect 9196 40879 9236 40888
rect 9292 41516 9332 41525
rect 9196 39416 9236 39425
rect 9196 32108 9236 39376
rect 9196 32059 9236 32068
rect 9196 28580 9236 28589
rect 9196 23120 9236 28540
rect 9292 26312 9332 41476
rect 9292 26263 9332 26272
rect 9484 26228 9524 95656
rect 10636 94940 10676 94949
rect 9772 94688 9812 94697
rect 9676 88052 9716 88061
rect 9580 78308 9620 78317
rect 9580 70664 9620 78268
rect 9676 71504 9716 88012
rect 9676 71455 9716 71464
rect 9580 70615 9620 70624
rect 9676 70580 9716 70589
rect 9676 63188 9716 70540
rect 9676 63139 9716 63148
rect 9772 51932 9812 94648
rect 10540 94688 10580 94697
rect 9964 94016 10004 94025
rect 9868 78980 9908 78989
rect 9868 72176 9908 78940
rect 9868 72127 9908 72136
rect 9772 51883 9812 51892
rect 9868 54200 9908 54209
rect 9484 26179 9524 26188
rect 9580 49580 9620 49589
rect 9388 26144 9428 26153
rect 9388 25388 9428 26104
rect 9388 25339 9428 25348
rect 9196 23071 9236 23080
rect 9292 25304 9332 25313
rect 9100 15007 9140 15016
rect 8908 13663 8948 13672
rect 9292 1952 9332 25264
rect 9580 15812 9620 49540
rect 9580 15763 9620 15772
rect 9676 48824 9716 48833
rect 9580 14888 9620 14897
rect 9580 12452 9620 14848
rect 9580 12403 9620 12412
rect 9292 1903 9332 1912
rect 8812 1231 8852 1240
rect 9676 1196 9716 48784
rect 9676 1147 9716 1156
rect 9772 48740 9812 48749
rect 6892 307 6932 316
rect 9772 356 9812 48700
rect 9868 3128 9908 54160
rect 9964 53528 10004 93976
rect 10156 93932 10196 93941
rect 9964 53479 10004 53488
rect 10060 71588 10100 71597
rect 10060 48824 10100 71548
rect 10156 62012 10196 93892
rect 10252 86372 10292 86381
rect 10252 76964 10292 86332
rect 10444 85616 10484 85625
rect 10444 82844 10484 85576
rect 10444 82795 10484 82804
rect 10444 78812 10484 78821
rect 10252 76915 10292 76924
rect 10348 77468 10388 77477
rect 10348 76628 10388 77428
rect 10348 73688 10388 76588
rect 10348 73639 10388 73648
rect 10252 70076 10292 70085
rect 10252 67556 10292 70036
rect 10252 67507 10292 67516
rect 10348 69152 10388 69161
rect 10156 61963 10196 61972
rect 10348 50252 10388 69112
rect 10444 52520 10484 78772
rect 10444 52471 10484 52480
rect 10348 50203 10388 50212
rect 10060 48775 10100 48784
rect 10156 49580 10196 49589
rect 9964 44204 10004 44213
rect 9964 3212 10004 44164
rect 10060 26228 10100 26237
rect 10060 25304 10100 26188
rect 10060 25255 10100 25264
rect 10156 5984 10196 49540
rect 10540 48908 10580 94648
rect 10636 66212 10676 94900
rect 10636 66163 10676 66172
rect 10732 94772 10772 94781
rect 10540 48859 10580 48868
rect 10636 53444 10676 53453
rect 10156 5935 10196 5944
rect 10252 48068 10292 48077
rect 10252 3548 10292 48028
rect 10540 47900 10580 47909
rect 10540 47228 10580 47860
rect 10444 46556 10484 46565
rect 10348 40004 10388 40013
rect 10348 37316 10388 39964
rect 10444 39836 10484 46516
rect 10540 41012 10580 47188
rect 10540 40963 10580 40972
rect 10444 39787 10484 39796
rect 10540 40844 10580 40853
rect 10540 37568 10580 40804
rect 10540 37519 10580 37528
rect 10348 37267 10388 37276
rect 10444 32108 10484 32117
rect 10444 29924 10484 32068
rect 10444 29875 10484 29884
rect 10540 32024 10580 32033
rect 10348 29840 10388 29849
rect 10348 28664 10388 29800
rect 10540 28916 10580 31984
rect 10540 28867 10580 28876
rect 10348 28615 10388 28624
rect 10252 3499 10292 3508
rect 10348 19928 10388 19937
rect 9964 3163 10004 3172
rect 9868 3079 9908 3088
rect 10348 2624 10388 19888
rect 10636 9344 10676 53404
rect 10732 48908 10772 94732
rect 12364 94772 12404 94781
rect 11212 94688 11252 94697
rect 11020 94016 11060 94025
rect 10828 93932 10868 93941
rect 10828 50336 10868 93892
rect 10924 89900 10964 89909
rect 10924 79148 10964 89860
rect 10924 79099 10964 79108
rect 10828 49580 10868 50296
rect 10828 49531 10868 49540
rect 10924 76628 10964 76637
rect 10732 48859 10772 48868
rect 10828 42440 10868 42449
rect 10732 41096 10772 41105
rect 10732 34544 10772 41056
rect 10732 34495 10772 34504
rect 10732 32276 10772 32285
rect 10732 27572 10772 32236
rect 10828 30848 10868 42400
rect 10828 30799 10868 30808
rect 10732 27523 10772 27532
rect 10636 9295 10676 9304
rect 10732 23120 10772 23129
rect 10348 2575 10388 2584
rect 10732 2036 10772 23080
rect 10828 21524 10868 21533
rect 10828 2708 10868 21484
rect 10924 20180 10964 76588
rect 11020 50168 11060 93976
rect 11116 93932 11156 93941
rect 11116 62096 11156 93892
rect 11116 62047 11156 62056
rect 11020 50119 11060 50128
rect 11116 61844 11156 61853
rect 10924 20131 10964 20140
rect 11020 43532 11060 43541
rect 11020 8000 11060 43492
rect 11116 31604 11156 61804
rect 11212 51092 11252 94648
rect 11596 94688 11636 94697
rect 11404 69740 11444 69749
rect 11212 51043 11252 51052
rect 11308 65204 11348 65213
rect 11116 31555 11156 31564
rect 11212 50084 11252 50093
rect 11212 20348 11252 50044
rect 11308 40844 11348 65164
rect 11404 57644 11444 69700
rect 11404 57595 11444 57604
rect 11500 63692 11540 63701
rect 11308 40795 11348 40804
rect 11404 50336 11444 50345
rect 11308 38912 11348 38921
rect 11308 37568 11348 38872
rect 11308 33032 11348 37528
rect 11404 33284 11444 50296
rect 11404 33235 11444 33244
rect 11308 32983 11348 32992
rect 11212 20299 11252 20308
rect 11308 31436 11348 31445
rect 11308 17240 11348 31396
rect 11308 17191 11348 17200
rect 11404 22364 11444 22373
rect 11404 21944 11444 22324
rect 11404 16232 11444 21904
rect 11404 13964 11444 16192
rect 11404 13915 11444 13924
rect 11404 11024 11444 11033
rect 11404 10100 11444 10984
rect 11404 10051 11444 10060
rect 11020 7951 11060 7960
rect 10828 2659 10868 2668
rect 10732 1987 10772 1996
rect 11500 1952 11540 63652
rect 11596 60500 11636 94648
rect 12172 94688 12212 94697
rect 11884 93764 11924 93773
rect 11788 79736 11828 79745
rect 11596 60451 11636 60460
rect 11692 66968 11732 66977
rect 11692 66548 11732 66928
rect 11596 58568 11636 58577
rect 11596 57560 11636 58528
rect 11596 57511 11636 57520
rect 11596 33368 11636 33377
rect 11596 24968 11636 33328
rect 11596 24919 11636 24928
rect 11692 13460 11732 66508
rect 11788 27488 11828 79696
rect 11884 69152 11924 93724
rect 11884 69103 11924 69112
rect 11980 83012 12020 83021
rect 11884 62852 11924 62861
rect 11884 60248 11924 62812
rect 11884 60199 11924 60208
rect 11788 27439 11828 27448
rect 11884 59996 11924 60005
rect 11884 59240 11924 59956
rect 11692 13411 11732 13420
rect 11884 11864 11924 59200
rect 11980 32192 12020 82972
rect 11980 32143 12020 32152
rect 12076 80660 12116 80669
rect 11980 29252 12020 29261
rect 11980 25052 12020 29212
rect 11980 25003 12020 25012
rect 11884 11815 11924 11824
rect 12076 3380 12116 80620
rect 12172 60584 12212 94648
rect 12268 88892 12308 88901
rect 12268 62852 12308 88852
rect 12268 62803 12308 62812
rect 12172 60535 12212 60544
rect 12268 61172 12308 61181
rect 12172 59660 12212 59669
rect 12172 58232 12212 59620
rect 12172 58183 12212 58192
rect 12268 57980 12308 61132
rect 12268 57931 12308 57940
rect 12268 50336 12308 50345
rect 12172 47984 12212 47993
rect 12172 27404 12212 47944
rect 12268 30260 12308 50296
rect 12364 50252 12404 94732
rect 12460 94100 12500 94109
rect 12460 80072 12500 94060
rect 12460 80023 12500 80032
rect 12460 66380 12500 66389
rect 12460 63440 12500 66340
rect 12556 64196 12596 95908
rect 18220 94856 18260 94865
rect 13420 94772 13460 94781
rect 12748 94184 12788 94193
rect 12652 79988 12692 79997
rect 12652 74444 12692 79948
rect 12652 74395 12692 74404
rect 12556 64147 12596 64156
rect 12652 70496 12692 70505
rect 12460 63391 12500 63400
rect 12364 50203 12404 50212
rect 12460 60500 12500 60509
rect 12364 39752 12404 39761
rect 12364 36728 12404 39712
rect 12364 35720 12404 36688
rect 12364 35671 12404 35680
rect 12460 34544 12500 60460
rect 12652 60332 12692 70456
rect 12652 60283 12692 60292
rect 12652 50336 12692 50345
rect 12460 34495 12500 34504
rect 12556 46304 12596 46313
rect 12364 33368 12404 33377
rect 12364 33200 12404 33328
rect 12364 33151 12404 33160
rect 12268 30211 12308 30220
rect 12364 30344 12404 30353
rect 12172 27355 12212 27364
rect 12268 29084 12308 29093
rect 12268 26060 12308 29044
rect 12268 26011 12308 26020
rect 12364 12452 12404 30304
rect 12364 12403 12404 12412
rect 12460 30092 12500 30101
rect 12076 3331 12116 3340
rect 12460 2372 12500 30052
rect 12556 6068 12596 46264
rect 12556 6019 12596 6028
rect 12652 3800 12692 50296
rect 12748 48740 12788 94144
rect 13132 87968 13172 87977
rect 13036 86456 13076 86465
rect 12844 76460 12884 76469
rect 12844 73604 12884 76420
rect 12844 73555 12884 73564
rect 12844 73100 12884 73109
rect 12844 59912 12884 73060
rect 12844 59863 12884 59872
rect 12748 48691 12788 48700
rect 12940 43280 12980 43289
rect 12940 42720 12980 43240
rect 13036 42860 13076 86416
rect 13132 85028 13172 87928
rect 13132 84979 13172 84988
rect 13324 79820 13364 79829
rect 13324 75116 13364 79780
rect 13132 74528 13172 74537
rect 13132 67136 13172 74488
rect 13324 73352 13364 75076
rect 13324 73303 13364 73312
rect 13132 65120 13172 67096
rect 13132 65071 13172 65080
rect 13324 69152 13364 69161
rect 13228 65036 13268 65045
rect 13132 62516 13172 62525
rect 13132 58736 13172 62476
rect 13132 58687 13172 58696
rect 13036 42811 13076 42820
rect 13132 58568 13172 58577
rect 12940 42680 13076 42720
rect 12844 40340 12884 40349
rect 12748 37904 12788 37913
rect 12748 20852 12788 37864
rect 12748 20803 12788 20812
rect 12844 18668 12884 40300
rect 12940 39752 12980 39761
rect 12940 38996 12980 39712
rect 12940 38947 12980 38956
rect 13036 34056 13076 42680
rect 12940 34016 13076 34056
rect 12940 33116 12980 34016
rect 12940 33067 12980 33076
rect 13036 33872 13076 33881
rect 12940 29924 12980 29933
rect 12940 24380 12980 29884
rect 12940 24331 12980 24340
rect 12844 18619 12884 18628
rect 13036 16568 13076 33832
rect 13036 16519 13076 16528
rect 13036 14720 13076 14729
rect 13036 13124 13076 14680
rect 13036 13075 13076 13084
rect 12652 3751 12692 3760
rect 12460 2323 12500 2332
rect 11500 1903 11540 1912
rect 13132 1448 13172 58528
rect 13228 15392 13268 64996
rect 13324 63104 13364 69112
rect 13324 63055 13364 63064
rect 13228 15343 13268 15352
rect 13324 53360 13364 53369
rect 13132 1399 13172 1408
rect 13324 440 13364 53320
rect 13420 48740 13460 94732
rect 14380 94772 14420 94781
rect 13900 93932 13940 93941
rect 13804 89480 13844 89489
rect 13708 87968 13748 87977
rect 13612 82172 13652 82181
rect 13516 79904 13556 79913
rect 13516 78308 13556 79864
rect 13516 78259 13556 78268
rect 13516 64868 13556 64877
rect 13516 63272 13556 64828
rect 13516 63223 13556 63232
rect 13420 48691 13460 48700
rect 13516 46472 13556 46481
rect 13420 42860 13460 42869
rect 13420 40340 13460 42820
rect 13420 40291 13460 40300
rect 13420 39752 13460 39761
rect 13420 35300 13460 39712
rect 13516 36056 13556 46432
rect 13516 36007 13556 36016
rect 13420 35251 13460 35260
rect 13516 34628 13556 34637
rect 13420 33116 13460 33125
rect 13420 30092 13460 33076
rect 13420 30043 13460 30052
rect 13420 29756 13460 29765
rect 13420 23204 13460 29716
rect 13420 23155 13460 23164
rect 13420 20180 13460 20189
rect 13420 1952 13460 20140
rect 13516 17072 13556 34588
rect 13612 34460 13652 82132
rect 13708 42440 13748 87928
rect 13804 84104 13844 89440
rect 13804 82088 13844 84064
rect 13804 82039 13844 82048
rect 13708 42391 13748 42400
rect 13804 75620 13844 75629
rect 13708 42272 13748 42281
rect 13708 39416 13748 42232
rect 13708 39367 13748 39376
rect 13708 36644 13748 36653
rect 13708 35048 13748 36604
rect 13708 34999 13748 35008
rect 13804 34544 13844 75580
rect 13804 34495 13844 34504
rect 13612 34411 13652 34420
rect 13708 33284 13748 33293
rect 13612 32276 13652 32285
rect 13612 29084 13652 32236
rect 13612 29035 13652 29044
rect 13516 17023 13556 17032
rect 13612 21692 13652 21701
rect 13516 9596 13556 9605
rect 13516 8588 13556 9556
rect 13516 8539 13556 8548
rect 13612 2456 13652 21652
rect 13612 2407 13652 2416
rect 13420 1903 13460 1912
rect 13708 1364 13748 33244
rect 13804 31352 13844 31361
rect 13804 29420 13844 31312
rect 13804 26228 13844 29380
rect 13804 23288 13844 26188
rect 13804 23239 13844 23248
rect 13900 12452 13940 93892
rect 14284 93932 14324 93941
rect 14188 89060 14228 89069
rect 13996 85868 14036 85877
rect 13996 85028 14036 85828
rect 13996 75788 14036 84988
rect 14092 85196 14132 85205
rect 14092 83768 14132 85156
rect 14092 83719 14132 83728
rect 13996 75739 14036 75748
rect 14092 82760 14132 82769
rect 13996 68396 14036 68405
rect 13996 62936 14036 68356
rect 13996 62887 14036 62896
rect 13996 44960 14036 44969
rect 13996 40424 14036 44920
rect 13996 40375 14036 40384
rect 13996 38744 14036 38753
rect 13996 26312 14036 38704
rect 13996 26263 14036 26272
rect 14092 14804 14132 82720
rect 14188 31436 14228 89020
rect 14188 31387 14228 31396
rect 14092 14755 14132 14764
rect 14188 30260 14228 30269
rect 13900 11780 13940 12412
rect 13900 11731 13940 11740
rect 13708 1315 13748 1324
rect 14188 860 14228 30220
rect 14284 14552 14324 93892
rect 14380 16988 14420 94732
rect 16204 94184 16244 94193
rect 14668 93932 14708 93941
rect 14476 90740 14516 90749
rect 14476 84188 14516 90700
rect 14476 84139 14516 84148
rect 14476 76712 14516 76721
rect 14476 74444 14516 76672
rect 14476 74395 14516 74404
rect 14572 71252 14612 71261
rect 14476 69152 14516 69161
rect 14476 63692 14516 69112
rect 14476 63643 14516 63652
rect 14380 16939 14420 16948
rect 14476 60080 14516 60089
rect 14476 38240 14516 60040
rect 14284 14503 14324 14512
rect 14476 4136 14516 38200
rect 14572 21692 14612 71212
rect 14572 21643 14612 21652
rect 14572 20180 14612 20189
rect 14572 10100 14612 20140
rect 14668 13796 14708 93892
rect 15148 93932 15188 93941
rect 14860 89396 14900 89405
rect 14668 13747 14708 13756
rect 14764 83600 14804 83609
rect 14572 10051 14612 10060
rect 14476 4087 14516 4096
rect 14764 2624 14804 83560
rect 14860 33620 14900 89356
rect 14956 78140 14996 78149
rect 14956 35804 14996 78100
rect 15052 76376 15092 76385
rect 15052 73520 15092 76336
rect 15052 73471 15092 73480
rect 14956 35755 14996 35764
rect 15052 71252 15092 71261
rect 15052 70664 15092 71212
rect 14860 33571 14900 33580
rect 14956 34460 14996 34469
rect 14956 33368 14996 34420
rect 14860 33328 14996 33368
rect 14860 29756 14900 33328
rect 14860 29707 14900 29716
rect 14956 30008 14996 30017
rect 14860 29588 14900 29597
rect 14860 23792 14900 29548
rect 14956 29252 14996 29968
rect 14956 29203 14996 29212
rect 14860 23743 14900 23752
rect 15052 23120 15092 70624
rect 15052 23071 15092 23080
rect 15148 2876 15188 93892
rect 15340 87884 15380 87893
rect 15244 63608 15284 63617
rect 15244 62852 15284 63568
rect 15244 62803 15284 62812
rect 15244 62432 15284 62441
rect 15244 16484 15284 62392
rect 15340 51848 15380 87844
rect 15532 87884 15572 87893
rect 15436 66296 15476 66305
rect 15436 65288 15476 66256
rect 15436 65239 15476 65248
rect 15436 62684 15476 62693
rect 15436 59156 15476 62644
rect 15532 60500 15572 87844
rect 16108 82676 16148 82685
rect 16108 81584 16148 82636
rect 16108 81535 16148 81544
rect 15916 79316 15956 79325
rect 15820 76460 15860 76469
rect 15724 76292 15764 76301
rect 15628 71756 15668 71765
rect 15628 70580 15668 71716
rect 15628 70531 15668 70540
rect 15628 66212 15668 66221
rect 15628 61508 15668 66172
rect 15628 61459 15668 61468
rect 15532 60451 15572 60460
rect 15436 59107 15476 59116
rect 15340 51799 15380 51808
rect 15628 52184 15668 52193
rect 15436 40340 15476 40349
rect 15340 35384 15380 35393
rect 15340 20936 15380 35344
rect 15436 24632 15476 40300
rect 15532 38072 15572 38081
rect 15532 30932 15572 38032
rect 15532 30883 15572 30892
rect 15532 29840 15572 29849
rect 15532 27152 15572 29800
rect 15532 27103 15572 27112
rect 15436 24583 15476 24592
rect 15340 20887 15380 20896
rect 15340 20096 15380 20105
rect 15340 18500 15380 20056
rect 15340 18451 15380 18460
rect 15244 16435 15284 16444
rect 15628 9764 15668 52144
rect 15724 38408 15764 76252
rect 15820 71336 15860 76420
rect 15916 71588 15956 79276
rect 16012 73940 16052 73949
rect 16012 72932 16052 73900
rect 16012 72883 16052 72892
rect 15916 71539 15956 71548
rect 15820 71287 15860 71296
rect 15916 70580 15956 70589
rect 15916 48992 15956 70540
rect 16012 62432 16052 62441
rect 16012 61676 16052 62392
rect 16012 61627 16052 61636
rect 15916 48943 15956 48952
rect 16012 53360 16052 53369
rect 15724 38359 15764 38368
rect 15820 40004 15860 40013
rect 15820 32948 15860 39964
rect 15820 32899 15860 32908
rect 15916 36056 15956 36065
rect 15916 35552 15956 36016
rect 15820 32108 15860 32117
rect 15724 30008 15764 30017
rect 15724 29672 15764 29968
rect 15724 27152 15764 29632
rect 15724 27103 15764 27112
rect 15820 28832 15860 32068
rect 15916 30176 15956 35512
rect 15916 30127 15956 30136
rect 15820 20180 15860 28792
rect 15916 29420 15956 29429
rect 15916 23456 15956 29380
rect 15916 23407 15956 23416
rect 15820 20131 15860 20140
rect 16012 14972 16052 53320
rect 16108 49664 16148 49673
rect 16108 32108 16148 49624
rect 16108 32059 16148 32068
rect 16108 30260 16148 30269
rect 16108 26564 16148 30220
rect 16108 26515 16148 26524
rect 16108 23288 16148 23297
rect 16108 20684 16148 23248
rect 16108 20635 16148 20644
rect 16012 14923 16052 14932
rect 15628 9715 15668 9724
rect 15148 2827 15188 2836
rect 14764 2575 14804 2584
rect 14188 811 14228 820
rect 16204 524 16244 94144
rect 16972 94184 17012 94193
rect 16588 93932 16628 93941
rect 16492 89648 16532 89657
rect 16396 89060 16436 89069
rect 16300 77720 16340 77729
rect 16300 8168 16340 77680
rect 16396 60500 16436 89020
rect 16492 76292 16532 89608
rect 16492 76243 16532 76252
rect 16492 69320 16532 69329
rect 16492 65792 16532 69280
rect 16492 65743 16532 65752
rect 16396 60451 16436 60460
rect 16492 56132 16532 56141
rect 16300 8119 16340 8128
rect 16396 51932 16436 51941
rect 16396 1280 16436 51892
rect 16492 24044 16532 56092
rect 16588 27992 16628 93892
rect 16780 93680 16820 93689
rect 16684 86456 16724 86465
rect 16684 34544 16724 86416
rect 16684 34495 16724 34504
rect 16588 27943 16628 27952
rect 16492 23995 16532 24004
rect 16780 7160 16820 93640
rect 16876 84860 16916 84869
rect 16876 39752 16916 84820
rect 16876 39703 16916 39712
rect 16876 39164 16916 39173
rect 16876 30848 16916 39124
rect 16876 30799 16916 30808
rect 16780 7111 16820 7120
rect 16396 1231 16436 1240
rect 16972 1028 17012 94144
rect 18028 94184 18068 94193
rect 17740 93932 17780 93941
rect 17164 93344 17204 93353
rect 17068 78476 17108 78485
rect 17068 57644 17108 78436
rect 17068 57595 17108 57604
rect 17068 56216 17108 56225
rect 17068 31268 17108 56176
rect 17068 31219 17108 31228
rect 17164 1448 17204 93304
rect 17356 88136 17396 88145
rect 17260 85952 17300 85961
rect 17260 83852 17300 85912
rect 17260 83803 17300 83812
rect 17260 70076 17300 70085
rect 17260 62516 17300 70036
rect 17260 62467 17300 62476
rect 17260 60584 17300 60593
rect 17260 58568 17300 60544
rect 17260 58519 17300 58528
rect 17260 39668 17300 39677
rect 17260 32528 17300 39628
rect 17356 37400 17396 88096
rect 17644 87464 17684 87473
rect 17452 83600 17492 83609
rect 17452 83432 17492 83560
rect 17452 83383 17492 83392
rect 17452 80576 17492 80585
rect 17452 78140 17492 80536
rect 17452 74444 17492 78100
rect 17548 79820 17588 79829
rect 17548 77468 17588 79780
rect 17548 77419 17588 77428
rect 17452 70160 17492 74404
rect 17452 70111 17492 70120
rect 17548 75788 17588 75797
rect 17452 61508 17492 61517
rect 17452 57896 17492 61468
rect 17452 57847 17492 57856
rect 17356 37351 17396 37360
rect 17452 53360 17492 53369
rect 17260 32479 17300 32488
rect 17356 37232 17396 37241
rect 17356 12704 17396 37192
rect 17356 12655 17396 12664
rect 17452 4220 17492 53320
rect 17548 24464 17588 75748
rect 17644 56384 17684 87424
rect 17644 56335 17684 56344
rect 17548 24415 17588 24424
rect 17644 49328 17684 49337
rect 17452 4171 17492 4180
rect 17644 3464 17684 49288
rect 17644 3415 17684 3424
rect 17740 2792 17780 93892
rect 17932 86540 17972 86549
rect 17836 85784 17876 85793
rect 17836 59744 17876 85744
rect 17932 81836 17972 86500
rect 17932 81787 17972 81796
rect 17932 76796 17972 76805
rect 17932 71336 17972 76756
rect 17932 71287 17972 71296
rect 17932 70496 17972 70505
rect 17932 66296 17972 70456
rect 17932 63104 17972 66256
rect 17932 63055 17972 63064
rect 17836 59695 17876 59704
rect 17932 62852 17972 62861
rect 17932 62348 17972 62812
rect 17836 56216 17876 56225
rect 17836 37232 17876 56176
rect 17836 37183 17876 37192
rect 17836 34964 17876 34973
rect 17836 32864 17876 34924
rect 17836 32815 17876 32824
rect 17932 30344 17972 62308
rect 18028 51932 18068 94144
rect 18028 51883 18068 51892
rect 18124 93176 18164 93185
rect 18028 45212 18068 45221
rect 18028 38156 18068 45172
rect 18124 40424 18164 93136
rect 18220 64196 18260 94816
rect 18772 94520 19212 96768
rect 18772 94480 18808 94520
rect 18848 94480 18890 94520
rect 18930 94480 18972 94520
rect 19012 94480 19054 94520
rect 19094 94480 19136 94520
rect 19176 94480 19212 94520
rect 18772 93008 19212 94480
rect 20012 95276 20452 96768
rect 20012 95236 20048 95276
rect 20088 95236 20130 95276
rect 20170 95236 20212 95276
rect 20252 95236 20294 95276
rect 20334 95236 20376 95276
rect 20416 95236 20452 95276
rect 18772 92968 18808 93008
rect 18848 92968 18890 93008
rect 18930 92968 18972 93008
rect 19012 92968 19054 93008
rect 19094 92968 19136 93008
rect 19176 92968 19212 93008
rect 18772 91496 19212 92968
rect 18772 91456 18808 91496
rect 18848 91456 18890 91496
rect 18930 91456 18972 91496
rect 19012 91456 19054 91496
rect 19094 91456 19136 91496
rect 19176 91456 19212 91496
rect 18772 89984 19212 91456
rect 18772 89944 18808 89984
rect 18848 89944 18890 89984
rect 18930 89944 18972 89984
rect 19012 89944 19054 89984
rect 19094 89944 19136 89984
rect 19176 89944 19212 89984
rect 18604 88808 18644 88817
rect 18412 83600 18452 83609
rect 18316 83432 18356 83441
rect 18316 80744 18356 83392
rect 18316 80695 18356 80704
rect 18316 79148 18356 79157
rect 18316 76712 18356 79108
rect 18316 76663 18356 76672
rect 18316 76040 18356 76049
rect 18316 73772 18356 76000
rect 18316 73723 18356 73732
rect 18316 72428 18356 72437
rect 18316 68648 18356 72388
rect 18316 68599 18356 68608
rect 18220 64147 18260 64156
rect 18220 64028 18260 64037
rect 18220 63272 18260 63988
rect 18220 63223 18260 63232
rect 18316 63692 18356 63701
rect 18220 63104 18260 63113
rect 18220 61592 18260 63064
rect 18316 62852 18356 63652
rect 18316 62803 18356 62812
rect 18220 61543 18260 61552
rect 18316 59324 18356 59333
rect 18124 40375 18164 40384
rect 18220 58400 18260 58409
rect 18028 38107 18068 38116
rect 18124 39836 18164 39845
rect 18124 37704 18164 39796
rect 18028 37664 18164 37704
rect 18028 35216 18068 37664
rect 18028 35167 18068 35176
rect 18124 37568 18164 37577
rect 18124 34208 18164 37528
rect 18124 34159 18164 34168
rect 18124 33200 18164 33209
rect 17932 30295 17972 30304
rect 18028 33116 18068 33125
rect 18028 30092 18068 33076
rect 18124 32948 18164 33160
rect 18124 32899 18164 32908
rect 18124 32780 18164 32789
rect 18124 30428 18164 32740
rect 18124 30379 18164 30388
rect 17836 29756 17876 29765
rect 17836 26648 17876 29716
rect 17836 26599 17876 26608
rect 18028 29084 18068 30052
rect 18028 24716 18068 29044
rect 18124 30176 18164 30185
rect 18124 24800 18164 30136
rect 18124 24751 18164 24760
rect 18028 24667 18068 24676
rect 18124 24632 18164 24641
rect 18028 23624 18068 23633
rect 17836 22616 17876 22625
rect 17836 19928 17876 22576
rect 18028 21524 18068 23584
rect 18124 23372 18164 24592
rect 18124 23323 18164 23332
rect 18028 21475 18068 21484
rect 17836 19879 17876 19888
rect 17740 2743 17780 2752
rect 18220 1952 18260 58360
rect 18316 56384 18356 59284
rect 18316 54032 18356 56344
rect 18412 55544 18452 83560
rect 18412 55495 18452 55504
rect 18508 81500 18548 81509
rect 18316 53983 18356 53992
rect 18412 51932 18452 51941
rect 18316 38156 18356 38165
rect 18316 23792 18356 38116
rect 18316 23743 18356 23752
rect 18412 21692 18452 51892
rect 18508 30680 18548 81460
rect 18604 38996 18644 88768
rect 18604 38947 18644 38956
rect 18772 88472 19212 89944
rect 18772 88432 18808 88472
rect 18848 88432 18890 88472
rect 18930 88432 18972 88472
rect 19012 88432 19054 88472
rect 19094 88432 19136 88472
rect 19176 88432 19212 88472
rect 18772 86960 19212 88432
rect 18772 86920 18808 86960
rect 18848 86920 18890 86960
rect 18930 86920 18972 86960
rect 19012 86920 19054 86960
rect 19094 86920 19136 86960
rect 19176 86920 19212 86960
rect 18772 85448 19212 86920
rect 18772 85408 18808 85448
rect 18848 85408 18890 85448
rect 18930 85408 18972 85448
rect 19012 85408 19054 85448
rect 19094 85408 19136 85448
rect 19176 85408 19212 85448
rect 18772 83936 19212 85408
rect 19372 94184 19412 94193
rect 18772 83896 18808 83936
rect 18848 83896 18890 83936
rect 18930 83896 18972 83936
rect 19012 83896 19054 83936
rect 19094 83896 19136 83936
rect 19176 83896 19212 83936
rect 18772 82424 19212 83896
rect 18772 82384 18808 82424
rect 18848 82384 18890 82424
rect 18930 82384 18972 82424
rect 19012 82384 19054 82424
rect 19094 82384 19136 82424
rect 19176 82384 19212 82424
rect 18772 80912 19212 82384
rect 18772 80872 18808 80912
rect 18848 80872 18890 80912
rect 18930 80872 18972 80912
rect 19012 80872 19054 80912
rect 19094 80872 19136 80912
rect 19176 80872 19212 80912
rect 18772 79400 19212 80872
rect 18772 79360 18808 79400
rect 18848 79360 18890 79400
rect 18930 79360 18972 79400
rect 19012 79360 19054 79400
rect 19094 79360 19136 79400
rect 19176 79360 19212 79400
rect 18772 77888 19212 79360
rect 18772 77848 18808 77888
rect 18848 77848 18890 77888
rect 18930 77848 18972 77888
rect 19012 77848 19054 77888
rect 19094 77848 19136 77888
rect 19176 77848 19212 77888
rect 18772 76376 19212 77848
rect 18772 76336 18808 76376
rect 18848 76336 18890 76376
rect 18930 76336 18972 76376
rect 19012 76336 19054 76376
rect 19094 76336 19136 76376
rect 19176 76336 19212 76376
rect 18772 74864 19212 76336
rect 18772 74824 18808 74864
rect 18848 74824 18890 74864
rect 18930 74824 18972 74864
rect 19012 74824 19054 74864
rect 19094 74824 19136 74864
rect 19176 74824 19212 74864
rect 18772 73352 19212 74824
rect 18772 73312 18808 73352
rect 18848 73312 18890 73352
rect 18930 73312 18972 73352
rect 19012 73312 19054 73352
rect 19094 73312 19136 73352
rect 19176 73312 19212 73352
rect 18772 71840 19212 73312
rect 18772 71800 18808 71840
rect 18848 71800 18890 71840
rect 18930 71800 18972 71840
rect 19012 71800 19054 71840
rect 19094 71800 19136 71840
rect 19176 71800 19212 71840
rect 18772 70328 19212 71800
rect 18772 70288 18808 70328
rect 18848 70288 18890 70328
rect 18930 70288 18972 70328
rect 19012 70288 19054 70328
rect 19094 70288 19136 70328
rect 19176 70288 19212 70328
rect 18772 68816 19212 70288
rect 18772 68776 18808 68816
rect 18848 68776 18890 68816
rect 18930 68776 18972 68816
rect 19012 68776 19054 68816
rect 19094 68776 19136 68816
rect 19176 68776 19212 68816
rect 18772 67304 19212 68776
rect 18772 67264 18808 67304
rect 18848 67264 18890 67304
rect 18930 67264 18972 67304
rect 19012 67264 19054 67304
rect 19094 67264 19136 67304
rect 19176 67264 19212 67304
rect 18772 65792 19212 67264
rect 18772 65752 18808 65792
rect 18848 65752 18890 65792
rect 18930 65752 18972 65792
rect 19012 65752 19054 65792
rect 19094 65752 19136 65792
rect 19176 65752 19212 65792
rect 18772 64280 19212 65752
rect 18772 64240 18808 64280
rect 18848 64240 18890 64280
rect 18930 64240 18972 64280
rect 19012 64240 19054 64280
rect 19094 64240 19136 64280
rect 19176 64240 19212 64280
rect 18772 62768 19212 64240
rect 18772 62728 18808 62768
rect 18848 62728 18890 62768
rect 18930 62728 18972 62768
rect 19012 62728 19054 62768
rect 19094 62728 19136 62768
rect 19176 62728 19212 62768
rect 18772 61256 19212 62728
rect 18772 61216 18808 61256
rect 18848 61216 18890 61256
rect 18930 61216 18972 61256
rect 19012 61216 19054 61256
rect 19094 61216 19136 61256
rect 19176 61216 19212 61256
rect 18772 59744 19212 61216
rect 18772 59704 18808 59744
rect 18848 59704 18890 59744
rect 18930 59704 18972 59744
rect 19012 59704 19054 59744
rect 19094 59704 19136 59744
rect 19176 59704 19212 59744
rect 18772 58232 19212 59704
rect 18772 58192 18808 58232
rect 18848 58192 18890 58232
rect 18930 58192 18972 58232
rect 19012 58192 19054 58232
rect 19094 58192 19136 58232
rect 19176 58192 19212 58232
rect 18772 56720 19212 58192
rect 18772 56680 18808 56720
rect 18848 56680 18890 56720
rect 18930 56680 18972 56720
rect 19012 56680 19054 56720
rect 19094 56680 19136 56720
rect 19176 56680 19212 56720
rect 18772 55208 19212 56680
rect 18772 55168 18808 55208
rect 18848 55168 18890 55208
rect 18930 55168 18972 55208
rect 19012 55168 19054 55208
rect 19094 55168 19136 55208
rect 19176 55168 19212 55208
rect 18772 53696 19212 55168
rect 18772 53656 18808 53696
rect 18848 53656 18890 53696
rect 18930 53656 18972 53696
rect 19012 53656 19054 53696
rect 19094 53656 19136 53696
rect 19176 53656 19212 53696
rect 18772 52184 19212 53656
rect 18772 52144 18808 52184
rect 18848 52144 18890 52184
rect 18930 52144 18972 52184
rect 19012 52144 19054 52184
rect 19094 52144 19136 52184
rect 19176 52144 19212 52184
rect 18772 50672 19212 52144
rect 18772 50632 18808 50672
rect 18848 50632 18890 50672
rect 18930 50632 18972 50672
rect 19012 50632 19054 50672
rect 19094 50632 19136 50672
rect 19176 50632 19212 50672
rect 18772 49160 19212 50632
rect 18772 49120 18808 49160
rect 18848 49120 18890 49160
rect 18930 49120 18972 49160
rect 19012 49120 19054 49160
rect 19094 49120 19136 49160
rect 19176 49120 19212 49160
rect 18772 47648 19212 49120
rect 19276 84188 19316 84197
rect 19276 48236 19316 84148
rect 19276 48187 19316 48196
rect 18772 47608 18808 47648
rect 18848 47608 18890 47648
rect 18930 47608 18972 47648
rect 19012 47608 19054 47648
rect 19094 47608 19136 47648
rect 19176 47608 19212 47648
rect 18772 46136 19212 47608
rect 18772 46096 18808 46136
rect 18848 46096 18890 46136
rect 18930 46096 18972 46136
rect 19012 46096 19054 46136
rect 19094 46096 19136 46136
rect 19176 46096 19212 46136
rect 18772 44624 19212 46096
rect 18772 44584 18808 44624
rect 18848 44584 18890 44624
rect 18930 44584 18972 44624
rect 19012 44584 19054 44624
rect 19094 44584 19136 44624
rect 19176 44584 19212 44624
rect 18772 43112 19212 44584
rect 18772 43072 18808 43112
rect 18848 43072 18890 43112
rect 18930 43072 18972 43112
rect 19012 43072 19054 43112
rect 19094 43072 19136 43112
rect 19176 43072 19212 43112
rect 18772 41600 19212 43072
rect 18772 41560 18808 41600
rect 18848 41560 18890 41600
rect 18930 41560 18972 41600
rect 19012 41560 19054 41600
rect 19094 41560 19136 41600
rect 19176 41560 19212 41600
rect 18772 40088 19212 41560
rect 18772 40048 18808 40088
rect 18848 40048 18890 40088
rect 18930 40048 18972 40088
rect 19012 40048 19054 40088
rect 19094 40048 19136 40088
rect 19176 40048 19212 40088
rect 18604 38828 18644 38837
rect 18604 33284 18644 38788
rect 18604 33235 18644 33244
rect 18772 38576 19212 40048
rect 18772 38536 18808 38576
rect 18848 38536 18890 38576
rect 18930 38536 18972 38576
rect 19012 38536 19054 38576
rect 19094 38536 19136 38576
rect 19176 38536 19212 38576
rect 18772 37064 19212 38536
rect 19276 48068 19316 48077
rect 19276 38156 19316 48028
rect 19276 38107 19316 38116
rect 18772 37024 18808 37064
rect 18848 37024 18890 37064
rect 18930 37024 18972 37064
rect 19012 37024 19054 37064
rect 19094 37024 19136 37064
rect 19176 37024 19212 37064
rect 18772 35552 19212 37024
rect 18772 35512 18808 35552
rect 18848 35512 18890 35552
rect 18930 35512 18972 35552
rect 19012 35512 19054 35552
rect 19094 35512 19136 35552
rect 19176 35512 19212 35552
rect 18772 34040 19212 35512
rect 18772 34000 18808 34040
rect 18848 34000 18890 34040
rect 18930 34000 18972 34040
rect 19012 34000 19054 34040
rect 19094 34000 19136 34040
rect 19176 34000 19212 34040
rect 18508 30631 18548 30640
rect 18604 33116 18644 33125
rect 18508 30008 18548 30017
rect 18508 27824 18548 29968
rect 18508 27775 18548 27784
rect 18604 27672 18644 33076
rect 18508 27632 18644 27672
rect 18772 32528 19212 34000
rect 18772 32488 18808 32528
rect 18848 32488 18890 32528
rect 18930 32488 18972 32528
rect 19012 32488 19054 32528
rect 19094 32488 19136 32528
rect 19176 32488 19212 32528
rect 18772 31016 19212 32488
rect 18772 30976 18808 31016
rect 18848 30976 18890 31016
rect 18930 30976 18972 31016
rect 19012 30976 19054 31016
rect 19094 30976 19136 31016
rect 19176 30976 19212 31016
rect 18772 29504 19212 30976
rect 18772 29464 18808 29504
rect 18848 29464 18890 29504
rect 18930 29464 18972 29504
rect 19012 29464 19054 29504
rect 19094 29464 19136 29504
rect 19176 29464 19212 29504
rect 18772 27992 19212 29464
rect 18772 27952 18808 27992
rect 18848 27952 18890 27992
rect 18930 27952 18972 27992
rect 19012 27952 19054 27992
rect 19094 27952 19136 27992
rect 19176 27952 19212 27992
rect 18508 26312 18548 27632
rect 18508 26263 18548 26272
rect 18604 27404 18644 27413
rect 18604 23288 18644 27364
rect 18604 23239 18644 23248
rect 18772 26480 19212 27952
rect 18772 26440 18808 26480
rect 18848 26440 18890 26480
rect 18930 26440 18972 26480
rect 19012 26440 19054 26480
rect 19094 26440 19136 26480
rect 19176 26440 19212 26480
rect 18772 24968 19212 26440
rect 19276 37988 19316 37997
rect 19276 25388 19316 37948
rect 19276 25339 19316 25348
rect 18772 24928 18808 24968
rect 18848 24928 18890 24968
rect 18930 24928 18972 24968
rect 19012 24928 19054 24968
rect 19094 24928 19136 24968
rect 19176 24928 19212 24968
rect 18772 23456 19212 24928
rect 18772 23416 18808 23456
rect 18848 23416 18890 23456
rect 18930 23416 18972 23456
rect 19012 23416 19054 23456
rect 19094 23416 19136 23456
rect 19176 23416 19212 23456
rect 18412 21643 18452 21652
rect 18508 22448 18548 22457
rect 18508 21524 18548 22408
rect 18508 21104 18548 21484
rect 18508 21055 18548 21064
rect 18772 21944 19212 23416
rect 18772 21904 18808 21944
rect 18848 21904 18890 21944
rect 18930 21904 18972 21944
rect 19012 21904 19054 21944
rect 19094 21904 19136 21944
rect 19176 21904 19212 21944
rect 18772 20432 19212 21904
rect 18772 20392 18808 20432
rect 18848 20392 18890 20432
rect 18930 20392 18972 20432
rect 19012 20392 19054 20432
rect 19094 20392 19136 20432
rect 19176 20392 19212 20432
rect 18604 20096 18644 20105
rect 18508 19340 18548 19349
rect 18508 16316 18548 19300
rect 18508 16267 18548 16276
rect 18604 15476 18644 20056
rect 18604 15427 18644 15436
rect 18772 18920 19212 20392
rect 18772 18880 18808 18920
rect 18848 18880 18890 18920
rect 18930 18880 18972 18920
rect 19012 18880 19054 18920
rect 19094 18880 19136 18920
rect 19176 18880 19212 18920
rect 18772 17408 19212 18880
rect 18772 17368 18808 17408
rect 18848 17368 18890 17408
rect 18930 17368 18972 17408
rect 19012 17368 19054 17408
rect 19094 17368 19136 17408
rect 19176 17368 19212 17408
rect 18772 15896 19212 17368
rect 18772 15856 18808 15896
rect 18848 15856 18890 15896
rect 18930 15856 18972 15896
rect 19012 15856 19054 15896
rect 19094 15856 19136 15896
rect 19176 15856 19212 15896
rect 18772 14384 19212 15856
rect 18772 14344 18808 14384
rect 18848 14344 18890 14384
rect 18930 14344 18972 14384
rect 19012 14344 19054 14384
rect 19094 14344 19136 14384
rect 19176 14344 19212 14384
rect 18316 13040 18356 13049
rect 18316 12872 18356 13000
rect 18316 12823 18356 12832
rect 18772 12872 19212 14344
rect 18772 12832 18808 12872
rect 18848 12832 18890 12872
rect 18930 12832 18972 12872
rect 19012 12832 19054 12872
rect 19094 12832 19136 12872
rect 19176 12832 19212 12872
rect 18220 1903 18260 1912
rect 18772 11360 19212 12832
rect 18772 11320 18808 11360
rect 18848 11320 18890 11360
rect 18930 11320 18972 11360
rect 19012 11320 19054 11360
rect 19094 11320 19136 11360
rect 19176 11320 19212 11360
rect 18772 9848 19212 11320
rect 19276 25220 19316 25229
rect 19276 10184 19316 25180
rect 19276 10135 19316 10144
rect 18772 9808 18808 9848
rect 18848 9808 18890 9848
rect 18930 9808 18972 9848
rect 19012 9808 19054 9848
rect 19094 9808 19136 9848
rect 19176 9808 19212 9848
rect 18772 8336 19212 9808
rect 18772 8296 18808 8336
rect 18848 8296 18890 8336
rect 18930 8296 18972 8336
rect 19012 8296 19054 8336
rect 19094 8296 19136 8336
rect 19176 8296 19212 8336
rect 18772 6824 19212 8296
rect 18772 6784 18808 6824
rect 18848 6784 18890 6824
rect 18930 6784 18972 6824
rect 19012 6784 19054 6824
rect 19094 6784 19136 6824
rect 19176 6784 19212 6824
rect 18772 5312 19212 6784
rect 18772 5272 18808 5312
rect 18848 5272 18890 5312
rect 18930 5272 18972 5312
rect 19012 5272 19054 5312
rect 19094 5272 19136 5312
rect 19176 5272 19212 5312
rect 18772 3800 19212 5272
rect 18772 3760 18808 3800
rect 18848 3760 18890 3800
rect 18930 3760 18972 3800
rect 19012 3760 19054 3800
rect 19094 3760 19136 3800
rect 19176 3760 19212 3800
rect 18772 2288 19212 3760
rect 18772 2248 18808 2288
rect 18848 2248 18890 2288
rect 18930 2248 18972 2288
rect 19012 2248 19054 2288
rect 19094 2248 19136 2288
rect 19176 2248 19212 2288
rect 17164 1399 17204 1408
rect 16972 979 17012 988
rect 16204 475 16244 484
rect 13324 391 13364 400
rect 9772 307 9812 316
rect 6412 223 6452 232
rect 18772 0 19212 2248
rect 19372 188 19412 94144
rect 20012 93764 20452 95236
rect 20012 93724 20048 93764
rect 20088 93724 20130 93764
rect 20170 93724 20212 93764
rect 20252 93724 20294 93764
rect 20334 93724 20376 93764
rect 20416 93724 20452 93764
rect 19852 93344 19892 93353
rect 19468 92672 19508 92681
rect 19468 38324 19508 92632
rect 19660 92672 19700 92681
rect 19468 38275 19508 38284
rect 19564 91832 19604 91841
rect 19468 38156 19508 38165
rect 19468 25220 19508 38116
rect 19468 25171 19508 25180
rect 19468 25052 19508 25061
rect 19468 1448 19508 25012
rect 19564 9680 19604 91792
rect 19660 18096 19700 92632
rect 19756 87296 19796 87305
rect 19756 48404 19796 87256
rect 19756 48355 19796 48364
rect 19756 48236 19796 48245
rect 19756 18248 19796 48196
rect 19756 18199 19796 18208
rect 19660 18056 19796 18096
rect 19564 9631 19604 9640
rect 19660 17996 19700 18005
rect 19660 6320 19700 17956
rect 19756 10772 19796 18056
rect 19756 10723 19796 10732
rect 19660 6271 19700 6280
rect 19468 1399 19508 1408
rect 19852 608 19892 93304
rect 19852 559 19892 568
rect 20012 92252 20452 93724
rect 21484 94184 21524 94193
rect 20012 92212 20048 92252
rect 20088 92212 20130 92252
rect 20170 92212 20212 92252
rect 20252 92212 20294 92252
rect 20334 92212 20376 92252
rect 20416 92212 20452 92252
rect 20012 90740 20452 92212
rect 21388 93344 21428 93353
rect 20012 90700 20048 90740
rect 20088 90700 20130 90740
rect 20170 90700 20212 90740
rect 20252 90700 20294 90740
rect 20334 90700 20376 90740
rect 20416 90700 20452 90740
rect 20012 89228 20452 90700
rect 20908 91160 20948 91169
rect 20012 89188 20048 89228
rect 20088 89188 20130 89228
rect 20170 89188 20212 89228
rect 20252 89188 20294 89228
rect 20334 89188 20376 89228
rect 20416 89188 20452 89228
rect 20012 87716 20452 89188
rect 20812 89648 20852 89657
rect 20012 87676 20048 87716
rect 20088 87676 20130 87716
rect 20170 87676 20212 87716
rect 20252 87676 20294 87716
rect 20334 87676 20376 87716
rect 20416 87676 20452 87716
rect 20012 86204 20452 87676
rect 20012 86164 20048 86204
rect 20088 86164 20130 86204
rect 20170 86164 20212 86204
rect 20252 86164 20294 86204
rect 20334 86164 20376 86204
rect 20416 86164 20452 86204
rect 20012 84692 20452 86164
rect 20012 84652 20048 84692
rect 20088 84652 20130 84692
rect 20170 84652 20212 84692
rect 20252 84652 20294 84692
rect 20334 84652 20376 84692
rect 20416 84652 20452 84692
rect 20012 83180 20452 84652
rect 20524 88640 20564 88649
rect 20524 84608 20564 88600
rect 20524 84559 20564 84568
rect 20716 86624 20756 86633
rect 20012 83140 20048 83180
rect 20088 83140 20130 83180
rect 20170 83140 20212 83180
rect 20252 83140 20294 83180
rect 20334 83140 20376 83180
rect 20416 83140 20452 83180
rect 20012 81668 20452 83140
rect 20012 81628 20048 81668
rect 20088 81628 20130 81668
rect 20170 81628 20212 81668
rect 20252 81628 20294 81668
rect 20334 81628 20376 81668
rect 20416 81628 20452 81668
rect 20012 80156 20452 81628
rect 20012 80116 20048 80156
rect 20088 80116 20130 80156
rect 20170 80116 20212 80156
rect 20252 80116 20294 80156
rect 20334 80116 20376 80156
rect 20416 80116 20452 80156
rect 20012 78644 20452 80116
rect 20012 78604 20048 78644
rect 20088 78604 20130 78644
rect 20170 78604 20212 78644
rect 20252 78604 20294 78644
rect 20334 78604 20376 78644
rect 20416 78604 20452 78644
rect 20012 77132 20452 78604
rect 20012 77092 20048 77132
rect 20088 77092 20130 77132
rect 20170 77092 20212 77132
rect 20252 77092 20294 77132
rect 20334 77092 20376 77132
rect 20416 77092 20452 77132
rect 20012 75620 20452 77092
rect 20012 75580 20048 75620
rect 20088 75580 20130 75620
rect 20170 75580 20212 75620
rect 20252 75580 20294 75620
rect 20334 75580 20376 75620
rect 20416 75580 20452 75620
rect 20012 74108 20452 75580
rect 20012 74068 20048 74108
rect 20088 74068 20130 74108
rect 20170 74068 20212 74108
rect 20252 74068 20294 74108
rect 20334 74068 20376 74108
rect 20416 74068 20452 74108
rect 20012 72596 20452 74068
rect 20524 76628 20564 76637
rect 20524 72680 20564 76588
rect 20620 75956 20660 75965
rect 20620 73436 20660 75916
rect 20620 73387 20660 73396
rect 20524 72631 20564 72640
rect 20012 72556 20048 72596
rect 20088 72556 20130 72596
rect 20170 72556 20212 72596
rect 20252 72556 20294 72596
rect 20334 72556 20376 72596
rect 20416 72556 20452 72596
rect 20012 71084 20452 72556
rect 20012 71044 20048 71084
rect 20088 71044 20130 71084
rect 20170 71044 20212 71084
rect 20252 71044 20294 71084
rect 20334 71044 20376 71084
rect 20416 71044 20452 71084
rect 20012 69572 20452 71044
rect 20620 69824 20660 69833
rect 20012 69532 20048 69572
rect 20088 69532 20130 69572
rect 20170 69532 20212 69572
rect 20252 69532 20294 69572
rect 20334 69532 20376 69572
rect 20416 69532 20452 69572
rect 20012 68060 20452 69532
rect 20012 68020 20048 68060
rect 20088 68020 20130 68060
rect 20170 68020 20212 68060
rect 20252 68020 20294 68060
rect 20334 68020 20376 68060
rect 20416 68020 20452 68060
rect 20012 66548 20452 68020
rect 20524 69740 20564 69749
rect 20524 67892 20564 69700
rect 20620 69152 20660 69784
rect 20620 69103 20660 69112
rect 20524 67843 20564 67852
rect 20620 68984 20660 68993
rect 20620 67800 20660 68944
rect 20012 66508 20048 66548
rect 20088 66508 20130 66548
rect 20170 66508 20212 66548
rect 20252 66508 20294 66548
rect 20334 66508 20376 66548
rect 20416 66508 20452 66548
rect 20012 65036 20452 66508
rect 20012 64996 20048 65036
rect 20088 64996 20130 65036
rect 20170 64996 20212 65036
rect 20252 64996 20294 65036
rect 20334 64996 20376 65036
rect 20416 64996 20452 65036
rect 20012 63524 20452 64996
rect 20012 63484 20048 63524
rect 20088 63484 20130 63524
rect 20170 63484 20212 63524
rect 20252 63484 20294 63524
rect 20334 63484 20376 63524
rect 20416 63484 20452 63524
rect 20012 62012 20452 63484
rect 20012 61972 20048 62012
rect 20088 61972 20130 62012
rect 20170 61972 20212 62012
rect 20252 61972 20294 62012
rect 20334 61972 20376 62012
rect 20416 61972 20452 62012
rect 20012 60500 20452 61972
rect 20012 60460 20048 60500
rect 20088 60460 20130 60500
rect 20170 60460 20212 60500
rect 20252 60460 20294 60500
rect 20334 60460 20376 60500
rect 20416 60460 20452 60500
rect 20012 58988 20452 60460
rect 20012 58948 20048 58988
rect 20088 58948 20130 58988
rect 20170 58948 20212 58988
rect 20252 58948 20294 58988
rect 20334 58948 20376 58988
rect 20416 58948 20452 58988
rect 20012 57476 20452 58948
rect 20524 67760 20660 67800
rect 20524 58820 20564 67760
rect 20620 66716 20660 66725
rect 20620 63440 20660 66676
rect 20620 63391 20660 63400
rect 20524 58771 20564 58780
rect 20012 57436 20048 57476
rect 20088 57436 20130 57476
rect 20170 57436 20212 57476
rect 20252 57436 20294 57476
rect 20334 57436 20376 57476
rect 20416 57436 20452 57476
rect 20012 55964 20452 57436
rect 20012 55924 20048 55964
rect 20088 55924 20130 55964
rect 20170 55924 20212 55964
rect 20252 55924 20294 55964
rect 20334 55924 20376 55964
rect 20416 55924 20452 55964
rect 20012 54452 20452 55924
rect 20012 54412 20048 54452
rect 20088 54412 20130 54452
rect 20170 54412 20212 54452
rect 20252 54412 20294 54452
rect 20334 54412 20376 54452
rect 20416 54412 20452 54452
rect 20012 52940 20452 54412
rect 20012 52900 20048 52940
rect 20088 52900 20130 52940
rect 20170 52900 20212 52940
rect 20252 52900 20294 52940
rect 20334 52900 20376 52940
rect 20416 52900 20452 52940
rect 20012 51428 20452 52900
rect 20012 51388 20048 51428
rect 20088 51388 20130 51428
rect 20170 51388 20212 51428
rect 20252 51388 20294 51428
rect 20334 51388 20376 51428
rect 20416 51388 20452 51428
rect 20012 49916 20452 51388
rect 20012 49876 20048 49916
rect 20088 49876 20130 49916
rect 20170 49876 20212 49916
rect 20252 49876 20294 49916
rect 20334 49876 20376 49916
rect 20416 49876 20452 49916
rect 20012 48404 20452 49876
rect 20012 48364 20048 48404
rect 20088 48364 20130 48404
rect 20170 48364 20212 48404
rect 20252 48364 20294 48404
rect 20334 48364 20376 48404
rect 20416 48364 20452 48404
rect 20012 46892 20452 48364
rect 20012 46852 20048 46892
rect 20088 46852 20130 46892
rect 20170 46852 20212 46892
rect 20252 46852 20294 46892
rect 20334 46852 20376 46892
rect 20416 46852 20452 46892
rect 20012 45380 20452 46852
rect 20012 45340 20048 45380
rect 20088 45340 20130 45380
rect 20170 45340 20212 45380
rect 20252 45340 20294 45380
rect 20334 45340 20376 45380
rect 20416 45340 20452 45380
rect 20012 43868 20452 45340
rect 20012 43828 20048 43868
rect 20088 43828 20130 43868
rect 20170 43828 20212 43868
rect 20252 43828 20294 43868
rect 20334 43828 20376 43868
rect 20416 43828 20452 43868
rect 20012 42356 20452 43828
rect 20012 42316 20048 42356
rect 20088 42316 20130 42356
rect 20170 42316 20212 42356
rect 20252 42316 20294 42356
rect 20334 42316 20376 42356
rect 20416 42316 20452 42356
rect 20012 40844 20452 42316
rect 20012 40804 20048 40844
rect 20088 40804 20130 40844
rect 20170 40804 20212 40844
rect 20252 40804 20294 40844
rect 20334 40804 20376 40844
rect 20416 40804 20452 40844
rect 20012 39332 20452 40804
rect 20012 39292 20048 39332
rect 20088 39292 20130 39332
rect 20170 39292 20212 39332
rect 20252 39292 20294 39332
rect 20334 39292 20376 39332
rect 20416 39292 20452 39332
rect 20012 37820 20452 39292
rect 20012 37780 20048 37820
rect 20088 37780 20130 37820
rect 20170 37780 20212 37820
rect 20252 37780 20294 37820
rect 20334 37780 20376 37820
rect 20416 37780 20452 37820
rect 20012 36308 20452 37780
rect 20012 36268 20048 36308
rect 20088 36268 20130 36308
rect 20170 36268 20212 36308
rect 20252 36268 20294 36308
rect 20334 36268 20376 36308
rect 20416 36268 20452 36308
rect 20012 34796 20452 36268
rect 20012 34756 20048 34796
rect 20088 34756 20130 34796
rect 20170 34756 20212 34796
rect 20252 34756 20294 34796
rect 20334 34756 20376 34796
rect 20416 34756 20452 34796
rect 20012 33284 20452 34756
rect 20620 49496 20660 49505
rect 20012 33244 20048 33284
rect 20088 33244 20130 33284
rect 20170 33244 20212 33284
rect 20252 33244 20294 33284
rect 20334 33244 20376 33284
rect 20416 33244 20452 33284
rect 20012 31772 20452 33244
rect 20524 33368 20564 33377
rect 20524 33032 20564 33328
rect 20524 32983 20564 32992
rect 20012 31732 20048 31772
rect 20088 31732 20130 31772
rect 20170 31732 20212 31772
rect 20252 31732 20294 31772
rect 20334 31732 20376 31772
rect 20416 31732 20452 31772
rect 20012 30260 20452 31732
rect 20012 30220 20048 30260
rect 20088 30220 20130 30260
rect 20170 30220 20212 30260
rect 20252 30220 20294 30260
rect 20334 30220 20376 30260
rect 20416 30220 20452 30260
rect 20012 28748 20452 30220
rect 20012 28708 20048 28748
rect 20088 28708 20130 28748
rect 20170 28708 20212 28748
rect 20252 28708 20294 28748
rect 20334 28708 20376 28748
rect 20416 28708 20452 28748
rect 20012 27236 20452 28708
rect 20012 27196 20048 27236
rect 20088 27196 20130 27236
rect 20170 27196 20212 27236
rect 20252 27196 20294 27236
rect 20334 27196 20376 27236
rect 20416 27196 20452 27236
rect 20012 25724 20452 27196
rect 20012 25684 20048 25724
rect 20088 25684 20130 25724
rect 20170 25684 20212 25724
rect 20252 25684 20294 25724
rect 20334 25684 20376 25724
rect 20416 25684 20452 25724
rect 20012 24212 20452 25684
rect 20524 30344 20564 30353
rect 20524 25472 20564 30304
rect 20524 25423 20564 25432
rect 20012 24172 20048 24212
rect 20088 24172 20130 24212
rect 20170 24172 20212 24212
rect 20252 24172 20294 24212
rect 20334 24172 20376 24212
rect 20416 24172 20452 24212
rect 20012 22700 20452 24172
rect 20012 22660 20048 22700
rect 20088 22660 20130 22700
rect 20170 22660 20212 22700
rect 20252 22660 20294 22700
rect 20334 22660 20376 22700
rect 20416 22660 20452 22700
rect 20012 21188 20452 22660
rect 20012 21148 20048 21188
rect 20088 21148 20130 21188
rect 20170 21148 20212 21188
rect 20252 21148 20294 21188
rect 20334 21148 20376 21188
rect 20416 21148 20452 21188
rect 20012 19676 20452 21148
rect 20012 19636 20048 19676
rect 20088 19636 20130 19676
rect 20170 19636 20212 19676
rect 20252 19636 20294 19676
rect 20334 19636 20376 19676
rect 20416 19636 20452 19676
rect 20012 18164 20452 19636
rect 20524 24464 20564 24473
rect 20524 18584 20564 24424
rect 20620 19844 20660 49456
rect 20620 19795 20660 19804
rect 20524 18535 20564 18544
rect 20012 18124 20048 18164
rect 20088 18124 20130 18164
rect 20170 18124 20212 18164
rect 20252 18124 20294 18164
rect 20334 18124 20376 18164
rect 20416 18124 20452 18164
rect 20012 16652 20452 18124
rect 20012 16612 20048 16652
rect 20088 16612 20130 16652
rect 20170 16612 20212 16652
rect 20252 16612 20294 16652
rect 20334 16612 20376 16652
rect 20416 16612 20452 16652
rect 20012 15140 20452 16612
rect 20012 15100 20048 15140
rect 20088 15100 20130 15140
rect 20170 15100 20212 15140
rect 20252 15100 20294 15140
rect 20334 15100 20376 15140
rect 20416 15100 20452 15140
rect 20012 13628 20452 15100
rect 20012 13588 20048 13628
rect 20088 13588 20130 13628
rect 20170 13588 20212 13628
rect 20252 13588 20294 13628
rect 20334 13588 20376 13628
rect 20416 13588 20452 13628
rect 20012 12116 20452 13588
rect 20012 12076 20048 12116
rect 20088 12076 20130 12116
rect 20170 12076 20212 12116
rect 20252 12076 20294 12116
rect 20334 12076 20376 12116
rect 20416 12076 20452 12116
rect 20012 10604 20452 12076
rect 20012 10564 20048 10604
rect 20088 10564 20130 10604
rect 20170 10564 20212 10604
rect 20252 10564 20294 10604
rect 20334 10564 20376 10604
rect 20416 10564 20452 10604
rect 20012 9092 20452 10564
rect 20012 9052 20048 9092
rect 20088 9052 20130 9092
rect 20170 9052 20212 9092
rect 20252 9052 20294 9092
rect 20334 9052 20376 9092
rect 20416 9052 20452 9092
rect 20012 7580 20452 9052
rect 20012 7540 20048 7580
rect 20088 7540 20130 7580
rect 20170 7540 20212 7580
rect 20252 7540 20294 7580
rect 20334 7540 20376 7580
rect 20416 7540 20452 7580
rect 20012 6068 20452 7540
rect 20012 6028 20048 6068
rect 20088 6028 20130 6068
rect 20170 6028 20212 6068
rect 20252 6028 20294 6068
rect 20334 6028 20376 6068
rect 20416 6028 20452 6068
rect 20012 4556 20452 6028
rect 20716 5480 20756 86584
rect 20812 15308 20852 89608
rect 20908 22112 20948 91120
rect 21292 90320 21332 90329
rect 21196 87464 21236 87473
rect 21100 87296 21140 87305
rect 20908 22063 20948 22072
rect 21004 84272 21044 84281
rect 21004 17576 21044 84232
rect 21100 21440 21140 87256
rect 21196 85448 21236 87424
rect 21196 85399 21236 85408
rect 21292 85128 21332 90280
rect 21196 85088 21332 85128
rect 21196 34460 21236 85088
rect 21196 34411 21236 34420
rect 21292 83600 21332 83609
rect 21292 29168 21332 83560
rect 21388 45296 21428 93304
rect 21388 45247 21428 45256
rect 21292 29119 21332 29128
rect 21388 44960 21428 44969
rect 21100 21391 21140 21400
rect 21292 27320 21332 27329
rect 21004 17527 21044 17536
rect 20812 15259 20852 15268
rect 21292 8672 21332 27280
rect 21388 19508 21428 44920
rect 21388 19459 21428 19468
rect 21292 8623 21332 8632
rect 20716 5431 20756 5440
rect 20012 4516 20048 4556
rect 20088 4516 20130 4556
rect 20170 4516 20212 4556
rect 20252 4516 20294 4556
rect 20334 4516 20376 4556
rect 20416 4516 20452 4556
rect 20012 3044 20452 4516
rect 20012 3004 20048 3044
rect 20088 3004 20130 3044
rect 20170 3004 20212 3044
rect 20252 3004 20294 3044
rect 20334 3004 20376 3044
rect 20416 3004 20452 3044
rect 20012 1532 20452 3004
rect 20012 1492 20048 1532
rect 20088 1492 20130 1532
rect 20170 1492 20212 1532
rect 20252 1492 20294 1532
rect 20334 1492 20376 1532
rect 20416 1492 20452 1532
rect 19372 139 19412 148
rect 20012 0 20452 1492
rect 21484 1196 21524 94144
rect 21484 1147 21524 1156
use sg13g2_inv_1  _0297_
timestamp 1676382929
transform 1 0 4128 0 1 42336
box -48 -56 336 834
use sg13g2_inv_1  _0298_
timestamp 1676382929
transform -1 0 7200 0 1 40824
box -48 -56 336 834
use sg13g2_inv_1  _0299_
timestamp 1676382929
transform -1 0 7584 0 -1 46872
box -48 -56 336 834
use sg13g2_inv_1  _0300_
timestamp 1676382929
transform -1 0 20448 0 -1 74088
box -48 -56 336 834
use sg13g2_inv_1  _0301_
timestamp 1676382929
transform 1 0 12096 0 -1 78624
box -48 -56 336 834
use sg13g2_inv_1  _0302_
timestamp 1676382929
transform -1 0 5760 0 1 78624
box -48 -56 336 834
use sg13g2_inv_1  _0303_
timestamp 1676382929
transform -1 0 11520 0 -1 58968
box -48 -56 336 834
use sg13g2_inv_1  _0304_
timestamp 1676382929
transform 1 0 10368 0 1 46872
box -48 -56 336 834
use sg13g2_inv_1  _0305_
timestamp 1676382929
transform -1 0 14784 0 1 36288
box -48 -56 336 834
use sg13g2_inv_1  _0306_
timestamp 1676382929
transform 1 0 14112 0 -1 25704
box -48 -56 336 834
use sg13g2_inv_1  _0307_
timestamp 1676382929
transform 1 0 7104 0 1 34776
box -48 -56 336 834
use sg13g2_inv_1  _0308_
timestamp 1676382929
transform -1 0 9216 0 -1 65016
box -48 -56 336 834
use sg13g2_inv_1  _0309_
timestamp 1676382929
transform 1 0 19776 0 -1 77112
box -48 -56 336 834
use sg13g2_inv_1  _0310_
timestamp 1676382929
transform 1 0 13440 0 -1 86184
box -48 -56 336 834
use sg13g2_inv_1  _0311_
timestamp 1676382929
transform -1 0 9216 0 1 81648
box -48 -56 336 834
use sg13g2_inv_1  _0312_
timestamp 1676382929
transform -1 0 10848 0 1 52920
box -48 -56 336 834
use sg13g2_inv_1  _0313_
timestamp 1676382929
transform 1 0 16320 0 -1 60480
box -48 -56 336 834
use sg13g2_inv_1  _0314_
timestamp 1676382929
transform -1 0 16512 0 1 81648
box -48 -56 336 834
use sg13g2_inv_1  _0315_
timestamp 1676382929
transform 1 0 5664 0 1 83160
box -48 -56 336 834
use sg13g2_inv_1  _0316_
timestamp 1676382929
transform -1 0 5088 0 -1 33264
box -48 -56 336 834
use sg13g2_inv_1  _0317_
timestamp 1676382929
transform -1 0 5184 0 1 30240
box -48 -56 336 834
use sg13g2_inv_1  _0318_
timestamp 1676382929
transform 1 0 13440 0 1 19656
box -48 -56 336 834
use sg13g2_inv_1  _0319_
timestamp 1676382929
transform 1 0 13920 0 -1 19656
box -48 -56 336 834
use sg13g2_inv_1  _0320_
timestamp 1676382929
transform -1 0 18432 0 -1 36288
box -48 -56 336 834
use sg13g2_inv_1  _0321_
timestamp 1676382929
transform -1 0 18720 0 1 34776
box -48 -56 336 834
use sg13g2_inv_1  _0322_
timestamp 1676382929
transform 1 0 14112 0 -1 43848
box -48 -56 336 834
use sg13g2_inv_1  _0323_
timestamp 1676382929
transform 1 0 16032 0 1 40824
box -48 -56 336 834
use sg13g2_inv_1  _0324_
timestamp 1676382929
transform 1 0 2976 0 1 25704
box -48 -56 336 834
use sg13g2_inv_1  _0325_
timestamp 1676382929
transform 1 0 3168 0 1 27216
box -48 -56 336 834
use sg13g2_inv_1  _0326_
timestamp 1676382929
transform -1 0 18528 0 1 21168
box -48 -56 336 834
use sg13g2_inv_1  _0327_
timestamp 1676382929
transform -1 0 20448 0 1 19656
box -48 -56 336 834
use sg13g2_inv_1  _0328_
timestamp 1676382929
transform -1 0 14016 0 -1 31752
box -48 -56 336 834
use sg13g2_inv_1  _0329_
timestamp 1676382929
transform 1 0 12960 0 -1 30240
box -48 -56 336 834
use sg13g2_inv_1  _0330_
timestamp 1676382929
transform 1 0 12192 0 1 37800
box -48 -56 336 834
use sg13g2_inv_1  _0331_
timestamp 1676382929
transform 1 0 13440 0 -1 37800
box -48 -56 336 834
use sg13g2_inv_1  _0332_
timestamp 1676382929
transform -1 0 7104 0 1 43848
box -48 -56 336 834
use sg13g2_inv_1  _0333_
timestamp 1676382929
transform -1 0 6240 0 1 46872
box -48 -56 336 834
use sg13g2_inv_1  _0334_
timestamp 1676382929
transform 1 0 4512 0 1 39312
box -48 -56 336 834
use sg13g2_inv_1  _0335_
timestamp 1676382929
transform 1 0 5280 0 1 74088
box -48 -56 336 834
use sg13g2_inv_1  _0336_
timestamp 1676382929
transform 1 0 17472 0 1 74088
box -48 -56 336 834
use sg13g2_inv_1  _0337_
timestamp 1676382929
transform 1 0 12288 0 -1 86184
box -48 -56 336 834
use sg13g2_inv_1  _0338_
timestamp 1676382929
transform 1 0 3936 0 1 54432
box -48 -56 336 834
use sg13g2_inv_1  _0339_
timestamp 1676382929
transform 1 0 5280 0 -1 68040
box -48 -56 336 834
use sg13g2_mux4_1  _0340_
timestamp 1677257233
transform -1 0 9024 0 1 72576
box -48 -56 2064 834
use sg13g2_mux4_1  _0341_
timestamp 1677257233
transform 1 0 4032 0 -1 39312
box -48 -56 2064 834
use sg13g2_mux4_1  _0342_
timestamp 1677257233
transform 1 0 2496 0 -1 40824
box -48 -56 2064 834
use sg13g2_mux4_1  _0343_
timestamp 1677257233
transform 1 0 4896 0 1 48384
box -48 -56 2064 834
use sg13g2_o21ai_1  _0344_
timestamp 1685175443
transform -1 0 8064 0 1 45360
box -48 -56 538 834
use sg13g2_nor2_1  _0345_
timestamp 1676627187
transform -1 0 7488 0 1 43848
box -48 -56 432 834
use sg13g2_a22oi_1  _0346_
timestamp 1685173987
transform -1 0 7296 0 -1 45360
box -48 -56 624 834
use sg13g2_nand3_1  _0347_
timestamp 1683988354
transform 1 0 7104 0 1 45360
box -48 -56 528 834
use sg13g2_nand2_1  _0348_
timestamp 1676557249
transform -1 0 7296 0 -1 46872
box -48 -56 432 834
use sg13g2_o21ai_1  _0349_
timestamp 1685175443
transform -1 0 7104 0 1 45360
box -48 -56 538 834
use sg13g2_nand3b_1  _0350_
timestamp 1676573470
transform 1 0 7392 0 -1 45360
box -48 -56 720 834
use sg13g2_o21ai_1  _0351_
timestamp 1685175443
transform -1 0 9024 0 -1 45360
box -48 -56 538 834
use sg13g2_o21ai_1  _0352_
timestamp 1685175443
transform -1 0 8544 0 -1 45360
box -48 -56 538 834
use sg13g2_mux4_1  _0353_
timestamp 1677257233
transform 1 0 6336 0 -1 43848
box -48 -56 2064 834
use sg13g2_mux4_1  _0354_
timestamp 1677257233
transform 1 0 6144 0 1 42336
box -48 -56 2064 834
use sg13g2_mux2_1  _0355_
timestamp 1677247768
transform 1 0 8160 0 1 42336
box -48 -56 1008 834
use sg13g2_o21ai_1  _0356_
timestamp 1685175443
transform 1 0 9600 0 1 43848
box -48 -56 538 834
use sg13g2_a21oi_1  _0357_
timestamp 1683973020
transform -1 0 9600 0 1 43848
box -48 -56 528 834
use sg13g2_nand2b_1  _0358_
timestamp 1676567195
transform -1 0 17568 0 -1 72576
box -48 -56 528 834
use sg13g2_nor3_1  _0359_
timestamp 1676639442
transform 1 0 17568 0 -1 72576
box -48 -56 528 834
use sg13g2_a221oi_1  _0360_
timestamp 1685197497
transform 1 0 19200 0 1 72576
box -48 -56 816 834
use sg13g2_mux4_1  _0361_
timestamp 1677257233
transform 1 0 13344 0 -1 77112
box -48 -56 2064 834
use sg13g2_nand2b_1  _0362_
timestamp 1676567195
transform 1 0 14016 0 1 21168
box -48 -56 528 834
use sg13g2_nor3_1  _0363_
timestamp 1676639442
transform 1 0 13632 0 -1 22680
box -48 -56 528 834
use sg13g2_a221oi_1  _0364_
timestamp 1685197497
transform 1 0 14112 0 -1 22680
box -48 -56 816 834
use sg13g2_mux4_1  _0365_
timestamp 1677257233
transform 1 0 13824 0 -1 24192
box -48 -56 2064 834
use sg13g2_mux4_1  _0366_
timestamp 1677257233
transform 1 0 17472 0 1 69552
box -48 -56 2064 834
use sg13g2_mux4_1  _0367_
timestamp 1677257233
transform 1 0 14208 0 1 74088
box -48 -56 2064 834
use sg13g2_nand2b_1  _0368_
timestamp 1676567195
transform 1 0 12096 0 -1 80136
box -48 -56 528 834
use sg13g2_nor3_1  _0369_
timestamp 1676639442
transform -1 0 13056 0 -1 80136
box -48 -56 528 834
use sg13g2_a221oi_1  _0370_
timestamp 1685197497
transform 1 0 12672 0 1 78624
box -48 -56 816 834
use sg13g2_mux4_1  _0371_
timestamp 1677257233
transform -1 0 13920 0 1 75600
box -48 -56 2064 834
use sg13g2_nor3_1  _0372_
timestamp 1676639442
transform 1 0 11712 0 -1 36288
box -48 -56 528 834
use sg13g2_nand2b_1  _0373_
timestamp 1676567195
transform 1 0 13152 0 1 34776
box -48 -56 528 834
use sg13g2_a221oi_1  _0374_
timestamp 1685197497
transform 1 0 12192 0 -1 36288
box -48 -56 816 834
use sg13g2_mux4_1  _0375_
timestamp 1677257233
transform -1 0 14496 0 1 36288
box -48 -56 2064 834
use sg13g2_mux4_1  _0376_
timestamp 1677257233
transform 1 0 11040 0 1 81648
box -48 -56 2064 834
use sg13g2_mux4_1  _0377_
timestamp 1677257233
transform 1 0 13632 0 1 78624
box -48 -56 2064 834
use sg13g2_nand2b_1  _0378_
timestamp 1676567195
transform -1 0 3456 0 -1 78624
box -48 -56 528 834
use sg13g2_nor3_1  _0379_
timestamp 1676639442
transform -1 0 3648 0 1 78624
box -48 -56 528 834
use sg13g2_a221oi_1  _0380_
timestamp 1685197497
transform 1 0 3072 0 -1 80136
box -48 -56 816 834
use sg13g2_mux4_1  _0381_
timestamp 1677257233
transform 1 0 7584 0 -1 80136
box -48 -56 2064 834
use sg13g2_nor3_1  _0382_
timestamp 1676639442
transform 1 0 9504 0 -1 46872
box -48 -56 528 834
use sg13g2_nand2b_1  _0383_
timestamp 1676567195
transform 1 0 9984 0 -1 46872
box -48 -56 528 834
use sg13g2_a221oi_1  _0384_
timestamp 1685197497
transform 1 0 10752 0 -1 45360
box -48 -56 816 834
use sg13g2_mux4_1  _0385_
timestamp 1677257233
transform 1 0 7872 0 1 46872
box -48 -56 2064 834
use sg13g2_mux4_1  _0386_
timestamp 1677257233
transform 1 0 3264 0 1 74088
box -48 -56 2064 834
use sg13g2_mux4_1  _0387_
timestamp 1677257233
transform 1 0 7296 0 1 86184
box -48 -56 2064 834
use sg13g2_mux4_1  _0388_
timestamp 1677257233
transform -1 0 8736 0 -1 74088
box -48 -56 2064 834
use sg13g2_mux4_1  _0389_
timestamp 1677257233
transform 1 0 15072 0 -1 78624
box -48 -56 2064 834
use sg13g2_mux4_1  _0390_
timestamp 1677257233
transform 1 0 15744 0 1 49896
box -48 -56 2064 834
use sg13g2_mux4_1  _0391_
timestamp 1677257233
transform 1 0 13536 0 1 31752
box -48 -56 2064 834
use sg13g2_mux4_1  _0392_
timestamp 1677257233
transform 1 0 15552 0 -1 51408
box -48 -56 2064 834
use sg13g2_mux4_1  _0393_
timestamp 1677257233
transform 1 0 15360 0 1 77112
box -48 -56 2064 834
use sg13g2_mux4_1  _0394_
timestamp 1677257233
transform 1 0 11520 0 -1 71064
box -48 -56 2064 834
use sg13g2_mux4_1  _0395_
timestamp 1677257233
transform 1 0 10752 0 -1 43848
box -48 -56 2064 834
use sg13g2_mux4_1  _0396_
timestamp 1677257233
transform 1 0 10656 0 1 40824
box -48 -56 2064 834
use sg13g2_mux4_1  _0397_
timestamp 1677257233
transform 1 0 11520 0 1 48384
box -48 -56 2064 834
use sg13g2_mux4_1  _0398_
timestamp 1677257233
transform 1 0 11808 0 1 71064
box -48 -56 2064 834
use sg13g2_mux4_1  _0399_
timestamp 1677257233
transform -1 0 8928 0 1 69552
box -48 -56 2064 834
use sg13g2_mux4_1  _0400_
timestamp 1677257233
transform 1 0 5088 0 -1 42336
box -48 -56 2064 834
use sg13g2_mux4_1  _0401_
timestamp 1677257233
transform 1 0 2112 0 -1 36288
box -48 -56 2064 834
use sg13g2_mux4_1  _0402_
timestamp 1677257233
transform 1 0 4032 0 -1 48384
box -48 -56 2064 834
use sg13g2_mux4_1  _0403_
timestamp 1677257233
transform 1 0 6912 0 1 66528
box -48 -56 2064 834
use sg13g2_mux4_1  _0404_
timestamp 1677257233
transform -1 0 4800 0 1 51408
box -48 -56 2064 834
use sg13g2_mux4_1  _0405_
timestamp 1677257233
transform 1 0 2016 0 -1 48384
box -48 -56 2064 834
use sg13g2_mux4_1  _0406_
timestamp 1677257233
transform 1 0 2208 0 1 43848
box -48 -56 2064 834
use sg13g2_mux4_1  _0407_
timestamp 1677257233
transform 1 0 3168 0 1 46872
box -48 -56 2064 834
use sg13g2_mux4_1  _0408_
timestamp 1677257233
transform 1 0 2496 0 1 52920
box -48 -56 2064 834
use sg13g2_mux4_1  _0409_
timestamp 1677257233
transform 1 0 12576 0 -1 74088
box -48 -56 2064 834
use sg13g2_mux4_1  _0410_
timestamp 1677257233
transform 1 0 17952 0 1 48384
box -48 -56 2064 834
use sg13g2_mux4_1  _0411_
timestamp 1677257233
transform 1 0 17952 0 1 40824
box -48 -56 2064 834
use sg13g2_mux4_1  _0412_
timestamp 1677257233
transform -1 0 20448 0 1 49896
box -48 -56 2064 834
use sg13g2_mux4_1  _0413_
timestamp 1677257233
transform 1 0 12768 0 1 72576
box -48 -56 2064 834
use sg13g2_mux4_1  _0414_
timestamp 1677257233
transform 1 0 14784 0 -1 75600
box -48 -56 2064 834
use sg13g2_mux4_1  _0415_
timestamp 1677257233
transform 1 0 15552 0 -1 48384
box -48 -56 2064 834
use sg13g2_mux4_1  _0416_
timestamp 1677257233
transform 1 0 16320 0 1 30240
box -48 -56 2064 834
use sg13g2_mux4_1  _0417_
timestamp 1677257233
transform -1 0 17088 0 1 48384
box -48 -56 2064 834
use sg13g2_mux4_1  _0418_
timestamp 1677257233
transform 1 0 17760 0 1 74088
box -48 -56 2064 834
use sg13g2_mux4_1  _0419_
timestamp 1677257233
transform 1 0 7488 0 1 78624
box -48 -56 2064 834
use sg13g2_mux4_1  _0420_
timestamp 1677257233
transform 1 0 9504 0 -1 49896
box -48 -56 2064 834
use sg13g2_mux4_1  _0421_
timestamp 1677257233
transform 1 0 6912 0 -1 39312
box -48 -56 2064 834
use sg13g2_mux4_1  _0422_
timestamp 1677257233
transform 1 0 9024 0 1 49896
box -48 -56 2064 834
use sg13g2_mux4_1  _0423_
timestamp 1677257233
transform 1 0 8160 0 -1 77112
box -48 -56 2064 834
use sg13g2_nand2b_1  _0424_
timestamp 1676567195
transform 1 0 11904 0 1 57456
box -48 -56 528 834
use sg13g2_nor3_1  _0425_
timestamp 1676639442
transform -1 0 11904 0 1 57456
box -48 -56 528 834
use sg13g2_a221oi_1  _0426_
timestamp 1685197497
transform -1 0 11232 0 -1 58968
box -48 -56 816 834
use sg13g2_mux4_1  _0427_
timestamp 1677257233
transform 1 0 7872 0 1 60480
box -48 -56 2064 834
use sg13g2_nor3_1  _0428_
timestamp 1676639442
transform -1 0 8544 0 -1 33264
box -48 -56 528 834
use sg13g2_nand2b_1  _0429_
timestamp 1676567195
transform 1 0 7584 0 -1 33264
box -48 -56 528 834
use sg13g2_a221oi_1  _0430_
timestamp 1685197497
transform -1 0 8160 0 1 34776
box -48 -56 816 834
use sg13g2_mux4_1  _0431_
timestamp 1677257233
transform -1 0 10560 0 1 36288
box -48 -56 2064 834
use sg13g2_mux4_1  _0432_
timestamp 1677257233
transform 1 0 10560 0 1 58968
box -48 -56 2064 834
use sg13g2_mux4_1  _0433_
timestamp 1677257233
transform 1 0 17952 0 1 66528
box -48 -56 2064 834
use sg13g2_mux4_1  _0434_
timestamp 1677257233
transform 1 0 11040 0 1 66528
box -48 -56 2064 834
use sg13g2_mux4_1  _0435_
timestamp 1677257233
transform 1 0 2880 0 -1 74088
box -48 -56 2064 834
use sg13g2_mux4_1  _0436_
timestamp 1677257233
transform -1 0 4128 0 -1 65016
box -48 -56 2064 834
use sg13g2_mux4_1  _0437_
timestamp 1677257233
transform 1 0 15360 0 1 52920
box -48 -56 2064 834
use sg13g2_mux4_1  _0438_
timestamp 1677257233
transform 1 0 17952 0 -1 63504
box -48 -56 2064 834
use sg13g2_mux4_1  _0439_
timestamp 1677257233
transform 1 0 3360 0 1 55944
box -48 -56 2064 834
use sg13g2_mux4_1  _0440_
timestamp 1677257233
transform 1 0 2880 0 -1 68040
box -48 -56 2064 834
use sg13g2_mux4_1  _0441_
timestamp 1677257233
transform 1 0 13632 0 -1 63504
box -48 -56 2064 834
use sg13g2_mux4_1  _0442_
timestamp 1677257233
transform 1 0 18336 0 1 52920
box -48 -56 2064 834
use sg13g2_mux4_1  _0443_
timestamp 1677257233
transform 1 0 2016 0 -1 60480
box -48 -56 2064 834
use sg13g2_mux4_1  _0444_
timestamp 1677257233
transform 1 0 2496 0 -1 66528
box -48 -56 2064 834
use sg13g2_mux4_1  _0445_
timestamp 1677257233
transform 1 0 14976 0 -1 54432
box -48 -56 2064 834
use sg13g2_mux4_1  _0446_
timestamp 1677257233
transform 1 0 17952 0 1 63504
box -48 -56 2064 834
use sg13g2_mux4_1  _0447_
timestamp 1677257233
transform 1 0 3264 0 -1 61992
box -48 -56 2064 834
use sg13g2_mux4_1  _0448_
timestamp 1677257233
transform 1 0 2688 0 1 71064
box -48 -56 2064 834
use sg13g2_mux4_1  _0449_
timestamp 1677257233
transform 1 0 14592 0 1 61992
box -48 -56 2064 834
use sg13g2_mux4_1  _0450_
timestamp 1677257233
transform 1 0 18144 0 -1 54432
box -48 -56 2064 834
use sg13g2_mux4_1  _0451_
timestamp 1677257233
transform 1 0 2112 0 -1 58968
box -48 -56 2064 834
use sg13g2_mux4_1  _0452_
timestamp 1677257233
transform 1 0 2976 0 -1 69552
box -48 -56 2064 834
use sg13g2_mux4_1  _0453_
timestamp 1677257233
transform 1 0 14688 0 1 68040
box -48 -56 2064 834
use sg13g2_mux4_1  _0454_
timestamp 1677257233
transform 1 0 18144 0 1 57456
box -48 -56 2064 834
use sg13g2_mux4_1  _0455_
timestamp 1677257233
transform -1 0 10368 0 -1 58968
box -48 -56 2064 834
use sg13g2_mux4_1  _0456_
timestamp 1677257233
transform 1 0 4704 0 -1 57456
box -48 -56 2064 834
use sg13g2_mux4_1  _0457_
timestamp 1677257233
transform 1 0 2976 0 -1 77112
box -48 -56 2064 834
use sg13g2_mux4_1  _0458_
timestamp 1677257233
transform 1 0 3648 0 1 68040
box -48 -56 2064 834
use sg13g2_mux4_1  _0459_
timestamp 1677257233
transform 1 0 11232 0 -1 83160
box -48 -56 2064 834
use sg13g2_mux4_1  _0460_
timestamp 1677257233
transform 1 0 12480 0 1 65016
box -48 -56 2064 834
use sg13g2_mux4_1  _0461_
timestamp 1677257233
transform 1 0 17952 0 1 71064
box -48 -56 2064 834
use sg13g2_mux4_1  _0462_
timestamp 1677257233
transform 1 0 18240 0 1 58968
box -48 -56 2064 834
use sg13g2_mux4_1  _0463_
timestamp 1677257233
transform 1 0 9216 0 -1 54432
box -48 -56 2064 834
use sg13g2_mux4_1  _0464_
timestamp 1677257233
transform 1 0 3360 0 1 57456
box -48 -56 2064 834
use sg13g2_mux4_1  _0465_
timestamp 1677257233
transform 1 0 3456 0 -1 78624
box -48 -56 2064 834
use sg13g2_mux4_1  _0466_
timestamp 1677257233
transform 1 0 4224 0 -1 71064
box -48 -56 2064 834
use sg13g2_mux4_1  _0467_
timestamp 1677257233
transform 1 0 11136 0 -1 81648
box -48 -56 2064 834
use sg13g2_mux4_1  _0468_
timestamp 1677257233
transform 1 0 14976 0 1 65016
box -48 -56 2064 834
use sg13g2_mux4_1  _0469_
timestamp 1677257233
transform 1 0 18240 0 -1 72576
box -48 -56 2064 834
use sg13g2_mux4_1  _0470_
timestamp 1677257233
transform 1 0 18240 0 -1 61992
box -48 -56 2064 834
use sg13g2_mux4_1  _0471_
timestamp 1677257233
transform 1 0 8256 0 -1 55944
box -48 -56 2064 834
use sg13g2_mux4_1  _0472_
timestamp 1677257233
transform 1 0 3264 0 1 61992
box -48 -56 2064 834
use sg13g2_mux4_1  _0473_
timestamp 1677257233
transform 1 0 3264 0 1 75600
box -48 -56 2064 834
use sg13g2_mux4_1  _0474_
timestamp 1677257233
transform 1 0 2688 0 -1 72576
box -48 -56 2064 834
use sg13g2_mux4_1  _0475_
timestamp 1677257233
transform 1 0 11136 0 1 83160
box -48 -56 2064 834
use sg13g2_mux4_1  _0476_
timestamp 1677257233
transform 1 0 12096 0 1 68040
box -48 -56 2064 834
use sg13g2_mux4_1  _0477_
timestamp 1677257233
transform 1 0 18144 0 -1 69552
box -48 -56 2064 834
use sg13g2_mux4_1  _0478_
timestamp 1677257233
transform 1 0 18048 0 1 55944
box -48 -56 2064 834
use sg13g2_mux4_1  _0479_
timestamp 1677257233
transform 1 0 9408 0 1 54432
box -48 -56 2064 834
use sg13g2_mux4_1  _0480_
timestamp 1677257233
transform 1 0 5664 0 1 58968
box -48 -56 2064 834
use sg13g2_mux4_1  _0481_
timestamp 1677257233
transform 1 0 7680 0 1 68040
box -48 -56 2064 834
use sg13g2_mux4_1  _0482_
timestamp 1677257233
transform 1 0 14880 0 1 71064
box -48 -56 2064 834
use sg13g2_mux4_1  _0483_
timestamp 1677257233
transform 1 0 16512 0 1 80136
box -48 -56 2064 834
use sg13g2_mux4_1  _0484_
timestamp 1677257233
transform 1 0 4128 0 -1 65016
box -48 -56 2064 834
use sg13g2_mux4_1  _0485_
timestamp 1677257233
transform 1 0 5568 0 1 74088
box -48 -56 2064 834
use sg13g2_mux4_1  _0486_
timestamp 1677257233
transform 1 0 14688 0 -1 66528
box -48 -56 2064 834
use sg13g2_mux4_1  _0487_
timestamp 1677257233
transform 1 0 18048 0 -1 66528
box -48 -56 2064 834
use sg13g2_mux4_1  _0488_
timestamp 1677257233
transform 1 0 3456 0 1 60480
box -48 -56 2064 834
use sg13g2_mux4_1  _0489_
timestamp 1677257233
transform 1 0 6144 0 -1 72576
box -48 -56 2064 834
use sg13g2_mux4_1  _0490_
timestamp 1677257233
transform 1 0 14112 0 -1 69552
box -48 -56 2064 834
use sg13g2_mux4_1  _0491_
timestamp 1677257233
transform 1 0 16224 0 -1 61992
box -48 -56 2064 834
use sg13g2_mux4_1  _0492_
timestamp 1677257233
transform 1 0 5568 0 1 61992
box -48 -56 2064 834
use sg13g2_mux4_1  _0493_
timestamp 1677257233
transform 1 0 9792 0 1 61992
box -48 -56 2064 834
use sg13g2_mux4_1  _0494_
timestamp 1677257233
transform 1 0 18240 0 1 81648
box -48 -56 2064 834
use sg13g2_mux4_1  _0495_
timestamp 1677257233
transform 1 0 12864 0 1 87696
box -48 -56 2064 834
use sg13g2_mux4_1  _0496_
timestamp 1677257233
transform 1 0 2592 0 -1 84672
box -48 -56 2064 834
use sg13g2_mux4_1  _0497_
timestamp 1677257233
transform 1 0 6528 0 1 52920
box -48 -56 2064 834
use sg13g2_mux4_1  _0498_
timestamp 1677257233
transform 1 0 15168 0 -1 55944
box -48 -56 2064 834
use sg13g2_mux4_1  _0499_
timestamp 1677257233
transform 1 0 17664 0 1 83160
box -48 -56 2064 834
use sg13g2_mux4_1  _0500_
timestamp 1677257233
transform 1 0 4704 0 -1 87696
box -48 -56 2064 834
use sg13g2_mux4_1  _0501_
timestamp 1677257233
transform 1 0 9408 0 -1 65016
box -48 -56 2064 834
use sg13g2_mux4_1  _0502_
timestamp 1677257233
transform -1 0 19392 0 -1 87696
box -48 -56 2064 834
use sg13g2_mux4_1  _0503_
timestamp 1677257233
transform 1 0 14400 0 -1 89208
box -48 -56 2064 834
use sg13g2_mux4_1  _0504_
timestamp 1677257233
transform 1 0 3264 0 1 83160
box -48 -56 2064 834
use sg13g2_mux4_1  _0505_
timestamp 1677257233
transform 1 0 5760 0 1 51408
box -48 -56 2064 834
use sg13g2_mux4_1  _0506_
timestamp 1677257233
transform 1 0 13056 0 -1 57456
box -48 -56 2064 834
use sg13g2_mux4_1  _0507_
timestamp 1677257233
transform 1 0 14976 0 -1 84672
box -48 -56 2064 834
use sg13g2_mux4_1  _0508_
timestamp 1677257233
transform 1 0 6816 0 -1 87696
box -48 -56 2064 834
use sg13g2_mux4_1  _0509_
timestamp 1677257233
transform 1 0 9504 0 -1 61992
box -48 -56 2064 834
use sg13g2_mux4_1  _0510_
timestamp 1677257233
transform 1 0 18240 0 -1 81648
box -48 -56 2064 834
use sg13g2_mux4_1  _0511_
timestamp 1677257233
transform 1 0 12384 0 -1 89208
box -48 -56 2064 834
use sg13g2_mux4_1  _0512_
timestamp 1677257233
transform 1 0 3072 0 -1 83160
box -48 -56 2064 834
use sg13g2_mux4_1  _0513_
timestamp 1677257233
transform 1 0 6048 0 -1 54432
box -48 -56 2064 834
use sg13g2_mux4_1  _0514_
timestamp 1677257233
transform 1 0 15168 0 1 55944
box -48 -56 2064 834
use sg13g2_mux4_1  _0515_
timestamp 1677257233
transform 1 0 17664 0 -1 84672
box -48 -56 2064 834
use sg13g2_mux4_1  _0516_
timestamp 1677257233
transform 1 0 4704 0 1 87696
box -48 -56 2064 834
use sg13g2_mux4_1  _0517_
timestamp 1677257233
transform 1 0 9312 0 1 65016
box -48 -56 2064 834
use sg13g2_mux4_1  _0518_
timestamp 1677257233
transform 1 0 17376 0 1 86184
box -48 -56 2064 834
use sg13g2_mux4_1  _0519_
timestamp 1677257233
transform 1 0 12960 0 1 89208
box -48 -56 2064 834
use sg13g2_mux4_1  _0520_
timestamp 1677257233
transform 1 0 3072 0 1 81648
box -48 -56 2064 834
use sg13g2_mux4_1  _0521_
timestamp 1677257233
transform 1 0 5184 0 -1 52920
box -48 -56 2064 834
use sg13g2_mux4_1  _0522_
timestamp 1677257233
transform 1 0 13152 0 1 55944
box -48 -56 2064 834
use sg13g2_mux4_1  _0523_
timestamp 1677257233
transform 1 0 14976 0 1 84672
box -48 -56 2064 834
use sg13g2_mux4_1  _0524_
timestamp 1677257233
transform 1 0 4512 0 1 86184
box -48 -56 2064 834
use sg13g2_nor3_1  _0525_
timestamp 1676639442
transform 1 0 6048 0 -1 77112
box -48 -56 528 834
use sg13g2_nand2b_1  _0526_
timestamp 1676567195
transform 1 0 8640 0 -1 75600
box -48 -56 528 834
use sg13g2_a221oi_1  _0527_
timestamp 1685197497
transform 1 0 7872 0 -1 75600
box -48 -56 816 834
use sg13g2_nor3_1  _0528_
timestamp 1676639442
transform 1 0 16992 0 1 74088
box -48 -56 528 834
use sg13g2_nand2b_1  _0529_
timestamp 1676567195
transform -1 0 16992 0 1 74088
box -48 -56 528 834
use sg13g2_a221oi_1  _0530_
timestamp 1685197497
transform 1 0 17280 0 1 75600
box -48 -56 816 834
use sg13g2_nor3_1  _0531_
timestamp 1676639442
transform -1 0 13152 0 -1 87696
box -48 -56 528 834
use sg13g2_nand2b_1  _0532_
timestamp 1676567195
transform 1 0 13152 0 -1 87696
box -48 -56 528 834
use sg13g2_a221oi_1  _0533_
timestamp 1685197497
transform 1 0 12768 0 1 86184
box -48 -56 816 834
use sg13g2_nor3_1  _0534_
timestamp 1676639442
transform 1 0 3456 0 1 54432
box -48 -56 528 834
use sg13g2_nand2b_1  _0535_
timestamp 1676567195
transform 1 0 2976 0 1 54432
box -48 -56 528 834
use sg13g2_a221oi_1  _0536_
timestamp 1685197497
transform 1 0 3648 0 -1 54432
box -48 -56 816 834
use sg13g2_nor3_1  _0537_
timestamp 1676639442
transform 1 0 5376 0 -1 69552
box -48 -56 528 834
use sg13g2_nand2b_1  _0538_
timestamp 1676567195
transform 1 0 7104 0 -1 71064
box -48 -56 528 834
use sg13g2_a221oi_1  _0539_
timestamp 1685197497
transform 1 0 7488 0 -1 69552
box -48 -56 816 834
use sg13g2_mux2_1  _0540_
timestamp 1677247768
transform 1 0 7872 0 -1 63504
box -48 -56 1008 834
use sg13g2_nor2b_1  _0541_
timestamp 1685181386
transform 1 0 8448 0 -1 65016
box -54 -56 528 834
use sg13g2_o21ai_1  _0542_
timestamp 1685175443
transform 1 0 8928 0 1 63504
box -48 -56 538 834
use sg13g2_o21ai_1  _0543_
timestamp 1685175443
transform 1 0 8832 0 -1 63504
box -48 -56 538 834
use sg13g2_a21oi_1  _0544_
timestamp 1683973020
transform -1 0 8928 0 1 63504
box -48 -56 528 834
use sg13g2_mux4_1  _0545_
timestamp 1677257233
transform 1 0 7584 0 1 61992
box -48 -56 2064 834
use sg13g2_nor2_1  _0546_
timestamp 1676627187
transform -1 0 10080 0 -1 63504
box -48 -56 432 834
use sg13g2_nor2_1  _0547_
timestamp 1676627187
transform 1 0 9312 0 -1 63504
box -48 -56 432 834
use sg13g2_mux2_1  _0548_
timestamp 1677247768
transform 1 0 19008 0 1 77112
box -48 -56 1008 834
use sg13g2_nor2b_1  _0549_
timestamp 1685181386
transform -1 0 19968 0 -1 78624
box -54 -56 528 834
use sg13g2_o21ai_1  _0550_
timestamp 1685175443
transform 1 0 19968 0 -1 78624
box -48 -56 538 834
use sg13g2_o21ai_1  _0551_
timestamp 1685175443
transform 1 0 19680 0 1 78624
box -48 -56 538 834
use sg13g2_a21oi_1  _0552_
timestamp 1683973020
transform 1 0 19968 0 1 77112
box -48 -56 528 834
use sg13g2_mux4_1  _0553_
timestamp 1677257233
transform -1 0 19488 0 -1 78624
box -48 -56 2064 834
use sg13g2_nor2_1  _0554_
timestamp 1676627187
transform 1 0 14688 0 -1 78624
box -48 -56 432 834
use sg13g2_nor2_1  _0555_
timestamp 1676627187
transform -1 0 20064 0 1 83160
box -48 -56 432 834
use sg13g2_mux2_1  _0556_
timestamp 1677247768
transform 1 0 13152 0 -1 84672
box -48 -56 1008 834
use sg13g2_nor2b_1  _0557_
timestamp 1685181386
transform -1 0 14688 0 1 84672
box -54 -56 528 834
use sg13g2_o21ai_1  _0558_
timestamp 1685175443
transform -1 0 13440 0 -1 86184
box -48 -56 538 834
use sg13g2_o21ai_1  _0559_
timestamp 1685175443
transform -1 0 13152 0 -1 84672
box -48 -56 538 834
use sg13g2_a21oi_1  _0560_
timestamp 1683973020
transform 1 0 14112 0 -1 84672
box -48 -56 528 834
use sg13g2_mux4_1  _0561_
timestamp 1677257233
transform 1 0 12192 0 1 84672
box -48 -56 2064 834
use sg13g2_nor2_1  _0562_
timestamp 1676627187
transform -1 0 14976 0 -1 84672
box -48 -56 432 834
use sg13g2_nor2_1  _0563_
timestamp 1676627187
transform 1 0 12576 0 -1 86184
box -48 -56 432 834
use sg13g2_mux2_1  _0564_
timestamp 1677247768
transform 1 0 6720 0 -1 81648
box -48 -56 1008 834
use sg13g2_nor2b_1  _0565_
timestamp 1685181386
transform 1 0 6048 0 1 80136
box -54 -56 528 834
use sg13g2_o21ai_1  _0566_
timestamp 1685175443
transform 1 0 6720 0 1 81648
box -48 -56 538 834
use sg13g2_o21ai_1  _0567_
timestamp 1685175443
transform 1 0 6528 0 1 80136
box -48 -56 538 834
use sg13g2_a21oi_1  _0568_
timestamp 1683973020
transform -1 0 8160 0 -1 81648
box -48 -56 528 834
use sg13g2_mux4_1  _0569_
timestamp 1677257233
transform 1 0 4704 0 -1 81648
box -48 -56 2064 834
use sg13g2_nor2_1  _0570_
timestamp 1676627187
transform 1 0 7680 0 1 81648
box -48 -56 432 834
use sg13g2_nor2_1  _0571_
timestamp 1676627187
transform 1 0 8160 0 -1 81648
box -48 -56 432 834
use sg13g2_mux2_1  _0572_
timestamp 1677247768
transform 1 0 9216 0 1 52920
box -48 -56 1008 834
use sg13g2_nor2b_1  _0573_
timestamp 1685181386
transform -1 0 9120 0 1 52920
box -54 -56 528 834
use sg13g2_o21ai_1  _0574_
timestamp 1685175443
transform 1 0 9504 0 1 51408
box -48 -56 538 834
use sg13g2_o21ai_1  _0575_
timestamp 1685175443
transform 1 0 9984 0 -1 52920
box -48 -56 538 834
use sg13g2_a21oi_1  _0576_
timestamp 1683973020
transform -1 0 10464 0 1 51408
box -48 -56 528 834
use sg13g2_mux4_1  _0577_
timestamp 1677257233
transform 1 0 7968 0 -1 52920
box -48 -56 2064 834
use sg13g2_nor2_1  _0578_
timestamp 1676627187
transform -1 0 10848 0 1 51408
box -48 -56 432 834
use sg13g2_nor2_1  _0579_
timestamp 1676627187
transform 1 0 10464 0 -1 52920
box -48 -56 432 834
use sg13g2_mux2_1  _0580_
timestamp 1677247768
transform 1 0 16608 0 -1 60480
box -48 -56 1008 834
use sg13g2_nor2b_1  _0581_
timestamp 1685181386
transform -1 0 16320 0 -1 60480
box -54 -56 528 834
use sg13g2_o21ai_1  _0582_
timestamp 1685175443
transform -1 0 16224 0 1 57456
box -48 -56 538 834
use sg13g2_o21ai_1  _0583_
timestamp 1685175443
transform -1 0 15840 0 -1 60480
box -48 -56 538 834
use sg13g2_a21oi_1  _0584_
timestamp 1683973020
transform 1 0 17280 0 -1 58968
box -48 -56 528 834
use sg13g2_mux4_1  _0585_
timestamp 1677257233
transform 1 0 15264 0 -1 58968
box -48 -56 2064 834
use sg13g2_nor2_1  _0586_
timestamp 1676627187
transform -1 0 18144 0 -1 58968
box -48 -56 432 834
use sg13g2_nor2_1  _0587_
timestamp 1676627187
transform 1 0 17568 0 -1 60480
box -48 -56 432 834
use sg13g2_mux2_1  _0588_
timestamp 1677247768
transform -1 0 15840 0 -1 83160
box -48 -56 1008 834
use sg13g2_nor2b_1  _0589_
timestamp 1685181386
transform 1 0 15744 0 1 81648
box -54 -56 528 834
use sg13g2_o21ai_1  _0590_
timestamp 1685175443
transform -1 0 14880 0 -1 83160
box -48 -56 538 834
use sg13g2_o21ai_1  _0591_
timestamp 1685175443
transform 1 0 16704 0 -1 81648
box -48 -56 538 834
use sg13g2_a21oi_1  _0592_
timestamp 1683973020
transform -1 0 15360 0 1 83160
box -48 -56 528 834
use sg13g2_mux4_1  _0593_
timestamp 1677257233
transform 1 0 13728 0 1 81648
box -48 -56 2064 834
use sg13g2_nor2_1  _0594_
timestamp 1676627187
transform -1 0 16224 0 -1 83160
box -48 -56 432 834
use sg13g2_nor2_1  _0595_
timestamp 1676627187
transform -1 0 16608 0 -1 83160
box -48 -56 432 834
use sg13g2_mux2_1  _0596_
timestamp 1677247768
transform -1 0 8544 0 1 83160
box -48 -56 1008 834
use sg13g2_nor2b_1  _0597_
timestamp 1685181386
transform -1 0 7680 0 1 81648
box -54 -56 528 834
use sg13g2_o21ai_1  _0598_
timestamp 1685175443
transform 1 0 8544 0 1 83160
box -48 -56 538 834
use sg13g2_o21ai_1  _0599_
timestamp 1685175443
transform -1 0 8256 0 -1 84672
box -48 -56 538 834
use sg13g2_a21oi_1  _0600_
timestamp 1683973020
transform -1 0 7296 0 1 84672
box -48 -56 528 834
use sg13g2_mux4_1  _0601_
timestamp 1677257233
transform 1 0 5760 0 -1 84672
box -48 -56 2064 834
use sg13g2_nor2_1  _0602_
timestamp 1676627187
transform -1 0 8160 0 1 84672
box -48 -56 432 834
use sg13g2_nor2_1  _0603_
timestamp 1676627187
transform -1 0 8640 0 -1 84672
box -48 -56 432 834
use sg13g2_mux4_1  _0604_
timestamp 1677257233
transform 1 0 8544 0 1 22680
box -48 -56 2064 834
use sg13g2_mux4_1  _0605_
timestamp 1677257233
transform 1 0 13440 0 1 16632
box -48 -56 2064 834
use sg13g2_mux4_1  _0606_
timestamp 1677257233
transform 1 0 11712 0 1 12096
box -48 -56 2064 834
use sg13g2_mux4_1  _0607_
timestamp 1677257233
transform 1 0 9216 0 -1 34776
box -48 -56 2064 834
use sg13g2_mux4_1  _0608_
timestamp 1677257233
transform 1 0 7584 0 -1 57456
box -48 -56 2064 834
use sg13g2_mux4_1  _0609_
timestamp 1677257233
transform 1 0 5088 0 -1 33264
box -48 -56 2064 834
use sg13g2_mux4_1  _0610_
timestamp 1677257233
transform 1 0 13632 0 1 22680
box -48 -56 2064 834
use sg13g2_mux4_1  _0611_
timestamp 1677257233
transform 1 0 15360 0 1 36288
box -48 -56 2064 834
use sg13g2_mux4_1  _0612_
timestamp 1677257233
transform 1 0 10464 0 -1 46872
box -48 -56 2064 834
use sg13g2_mux4_1  _0613_
timestamp 1677257233
transform 1 0 2496 0 1 39312
box -48 -56 2064 834
use sg13g2_mux4_1  _0614_
timestamp 1677257233
transform 1 0 13536 0 -1 33264
box -48 -56 2064 834
use sg13g2_mux4_1  _0615_
timestamp 1677257233
transform 1 0 11328 0 -1 42336
box -48 -56 2064 834
use sg13g2_mux4_1  _0616_
timestamp 1677257233
transform 1 0 2112 0 1 36288
box -48 -56 2064 834
use sg13g2_mux4_1  _0617_
timestamp 1677257233
transform 1 0 2688 0 -1 34776
box -48 -56 2064 834
use sg13g2_mux4_1  _0618_
timestamp 1677257233
transform 1 0 18240 0 -1 27216
box -48 -56 2064 834
use sg13g2_mux4_1  _0619_
timestamp 1677257233
transform 1 0 16992 0 -1 30240
box -48 -56 2064 834
use sg13g2_mux4_1  _0620_
timestamp 1677257233
transform 1 0 6240 0 1 24192
box -48 -56 2064 834
use sg13g2_mux4_1  _0621_
timestamp 1677257233
transform 1 0 7392 0 1 18144
box -48 -56 2064 834
use sg13g2_mux4_1  _0622_
timestamp 1677257233
transform 1 0 12288 0 1 18144
box -48 -56 2064 834
use sg13g2_mux4_1  _0623_
timestamp 1677257233
transform 1 0 11328 0 1 10584
box -48 -56 2064 834
use sg13g2_mux4_1  _0624_
timestamp 1677257233
transform 1 0 9216 0 -1 21168
box -48 -56 2064 834
use sg13g2_mux4_1  _0625_
timestamp 1677257233
transform 1 0 5952 0 1 10584
box -48 -56 2064 834
use sg13g2_mux4_1  _0626_
timestamp 1677257233
transform 1 0 15264 0 1 6048
box -48 -56 2064 834
use sg13g2_mux4_1  _0627_
timestamp 1677257233
transform 1 0 8544 0 -1 12096
box -48 -56 2064 834
use sg13g2_mux4_1  _0628_
timestamp 1677257233
transform 1 0 2304 0 1 21168
box -48 -56 2064 834
use sg13g2_mux4_1  _0629_
timestamp 1677257233
transform 1 0 2304 0 1 12096
box -48 -56 2064 834
use sg13g2_mux4_1  _0630_
timestamp 1677257233
transform 1 0 8256 0 1 6048
box -48 -56 2064 834
use sg13g2_mux4_1  _0631_
timestamp 1677257233
transform 1 0 17760 0 1 9072
box -48 -56 2064 834
use sg13g2_mux4_1  _0632_
timestamp 1677257233
transform 1 0 3552 0 -1 16632
box -48 -56 2064 834
use sg13g2_mux4_1  _0633_
timestamp 1677257233
transform 1 0 6144 0 -1 9072
box -48 -56 2064 834
use sg13g2_mux4_1  _0634_
timestamp 1677257233
transform 1 0 13824 0 1 4536
box -48 -56 2064 834
use sg13g2_mux4_1  _0635_
timestamp 1677257233
transform 1 0 8256 0 -1 15120
box -48 -56 2064 834
use sg13g2_mux4_1  _0636_
timestamp 1677257233
transform 1 0 2304 0 1 18144
box -48 -56 2064 834
use sg13g2_mux4_1  _0637_
timestamp 1677257233
transform 1 0 2400 0 1 13608
box -48 -56 2064 834
use sg13g2_mux4_1  _0638_
timestamp 1677257233
transform 1 0 8544 0 -1 7560
box -48 -56 2064 834
use sg13g2_mux4_1  _0639_
timestamp 1677257233
transform -1 0 19872 0 -1 10584
box -48 -56 2064 834
use sg13g2_mux4_1  _0640_
timestamp 1677257233
transform 1 0 2880 0 1 16632
box -48 -56 2064 834
use sg13g2_mux4_1  _0641_
timestamp 1677257233
transform 1 0 7392 0 1 13608
box -48 -56 2064 834
use sg13g2_mux4_1  _0642_
timestamp 1677257233
transform 1 0 15648 0 -1 9072
box -48 -56 2064 834
use sg13g2_mux4_1  _0643_
timestamp 1677257233
transform 1 0 17760 0 1 12096
box -48 -56 2064 834
use sg13g2_mux4_1  _0644_
timestamp 1677257233
transform 1 0 3456 0 -1 22680
box -48 -56 2064 834
use sg13g2_mux4_1  _0645_
timestamp 1677257233
transform 1 0 9216 0 1 33264
box -48 -56 2064 834
use sg13g2_mux4_1  _0646_
timestamp 1677257233
transform 1 0 2688 0 -1 10584
box -48 -56 2064 834
use sg13g2_mux4_1  _0647_
timestamp 1677257233
transform 1 0 12096 0 -1 9072
box -48 -56 2064 834
use sg13g2_mux4_1  _0648_
timestamp 1677257233
transform 1 0 10752 0 -1 6048
box -48 -56 2064 834
use sg13g2_mux4_1  _0649_
timestamp 1677257233
transform 1 0 12672 0 -1 15120
box -48 -56 2064 834
use sg13g2_mux4_1  _0650_
timestamp 1677257233
transform 1 0 15264 0 1 10584
box -48 -56 2064 834
use sg13g2_mux4_1  _0651_
timestamp 1677257233
transform 1 0 8256 0 -1 18144
box -48 -56 2064 834
use sg13g2_mux4_1  _0652_
timestamp 1677257233
transform 1 0 3264 0 -1 18144
box -48 -56 2064 834
use sg13g2_mux4_1  _0653_
timestamp 1677257233
transform 1 0 9600 0 1 31752
box -48 -56 2064 834
use sg13g2_mux4_1  _0654_
timestamp 1677257233
transform 1 0 4128 0 -1 9072
box -48 -56 2064 834
use sg13g2_mux4_1  _0655_
timestamp 1677257233
transform 1 0 12288 0 -1 10584
box -48 -56 2064 834
use sg13g2_mux4_1  _0656_
timestamp 1677257233
transform 1 0 12768 0 -1 6048
box -48 -56 2064 834
use sg13g2_mux4_1  _0657_
timestamp 1677257233
transform 1 0 12960 0 1 13608
box -48 -56 2064 834
use sg13g2_mux4_1  _0658_
timestamp 1677257233
transform -1 0 18048 0 -1 15120
box -48 -56 2064 834
use sg13g2_mux4_1  _0659_
timestamp 1677257233
transform 1 0 7200 0 -1 21168
box -48 -56 2064 834
use sg13g2_mux4_1  _0660_
timestamp 1677257233
transform 1 0 2880 0 -1 19656
box -48 -56 2064 834
use sg13g2_mux4_1  _0661_
timestamp 1677257233
transform 1 0 9696 0 1 28728
box -48 -56 2064 834
use sg13g2_mux4_1  _0662_
timestamp 1677257233
transform 1 0 5376 0 1 13608
box -48 -56 2064 834
use sg13g2_mux4_1  _0663_
timestamp 1677257233
transform 1 0 12288 0 1 9072
box -48 -56 2064 834
use sg13g2_mux4_1  _0664_
timestamp 1677257233
transform 1 0 9120 0 1 9072
box -48 -56 2064 834
use sg13g2_mux4_1  _0665_
timestamp 1677257233
transform 1 0 13152 0 -1 16632
box -48 -56 2064 834
use sg13g2_mux4_1  _0666_
timestamp 1677257233
transform 1 0 17952 0 -1 13608
box -48 -56 2064 834
use sg13g2_mux4_1  _0667_
timestamp 1677257233
transform 1 0 6528 0 1 22680
box -48 -56 2064 834
use sg13g2_mux4_1  _0668_
timestamp 1677257233
transform 1 0 2880 0 -1 24192
box -48 -56 2064 834
use sg13g2_mux4_1  _0669_
timestamp 1677257233
transform 1 0 8832 0 1 16632
box -48 -56 2064 834
use sg13g2_mux4_1  _0670_
timestamp 1677257233
transform 1 0 14976 0 1 13608
box -48 -56 2064 834
use sg13g2_mux4_1  _0671_
timestamp 1677257233
transform 1 0 13248 0 -1 12096
box -48 -56 2064 834
use sg13g2_mux4_1  _0672_
timestamp 1677257233
transform 1 0 9504 0 -1 30240
box -48 -56 2064 834
use sg13g2_mux4_1  _0673_
timestamp 1677257233
transform 1 0 4032 0 1 9072
box -48 -56 2064 834
use sg13g2_mux4_1  _0674_
timestamp 1677257233
transform 1 0 10656 0 1 4536
box -48 -56 2064 834
use sg13g2_mux4_1  _0675_
timestamp 1677257233
transform 1 0 17376 0 -1 18144
box -48 -56 2064 834
use sg13g2_mux4_1  _0676_
timestamp 1677257233
transform 1 0 5472 0 -1 19656
box -48 -56 2064 834
use sg13g2_mux4_1  _0677_
timestamp 1677257233
transform 1 0 5184 0 1 12096
box -48 -56 2064 834
use sg13g2_mux4_1  _0678_
timestamp 1677257233
transform 1 0 10464 0 1 19656
box -48 -56 2064 834
use sg13g2_mux4_1  _0679_
timestamp 1677257233
transform 1 0 14976 0 -1 18144
box -48 -56 2064 834
use sg13g2_mux4_1  _0680_
timestamp 1677257233
transform 1 0 2880 0 1 24192
box -48 -56 2064 834
use sg13g2_nand3b_1  _0681_
timestamp 1676573470
transform 1 0 5856 0 -1 22680
box -48 -56 720 834
use sg13g2_nor2b_1  _0682_
timestamp 1685181386
transform 1 0 4896 0 1 21168
box -54 -56 528 834
use sg13g2_a21oi_1  _0683_
timestamp 1683973020
transform -1 0 8640 0 -1 22680
box -48 -56 528 834
use sg13g2_o21ai_1  _0684_
timestamp 1685175443
transform 1 0 8640 0 -1 22680
box -48 -56 538 834
use sg13g2_nand3b_1  _0685_
timestamp 1676573470
transform 1 0 15552 0 1 28728
box -48 -56 720 834
use sg13g2_nor2b_1  _0686_
timestamp 1685181386
transform 1 0 16320 0 -1 30240
box -54 -56 528 834
use sg13g2_a21oi_1  _0687_
timestamp 1683973020
transform 1 0 17856 0 1 28728
box -48 -56 528 834
use sg13g2_o21ai_1  _0688_
timestamp 1685175443
transform 1 0 16800 0 -1 27216
box -48 -56 538 834
use sg13g2_nand3b_1  _0689_
timestamp 1676573470
transform 1 0 19200 0 -1 28728
box -48 -56 720 834
use sg13g2_nor2b_1  _0690_
timestamp 1685181386
transform -1 0 20352 0 -1 28728
box -54 -56 528 834
use sg13g2_a21oi_1  _0691_
timestamp 1683973020
transform -1 0 19488 0 -1 30240
box -48 -56 528 834
use sg13g2_o21ai_1  _0692_
timestamp 1685175443
transform 1 0 19968 0 1 27216
box -48 -56 538 834
use sg13g2_nand3b_1  _0693_
timestamp 1676573470
transform 1 0 7200 0 -1 37800
box -48 -56 720 834
use sg13g2_nor2_1  _0694_
timestamp 1676627187
transform 1 0 6048 0 -1 36288
box -48 -56 432 834
use sg13g2_a21oi_1  _0695_
timestamp 1683973020
transform -1 0 8352 0 -1 37800
box -48 -56 528 834
use sg13g2_o21ai_1  _0696_
timestamp 1685175443
transform 1 0 8064 0 1 36288
box -48 -56 538 834
use sg13g2_nand3b_1  _0697_
timestamp 1676573470
transform -1 0 3456 0 1 33264
box -48 -56 720 834
use sg13g2_nor2b_1  _0698_
timestamp 1685181386
transform 1 0 2208 0 -1 34776
box -54 -56 528 834
use sg13g2_a21oi_1  _0699_
timestamp 1683973020
transform 1 0 3456 0 1 33264
box -48 -56 528 834
use sg13g2_o21ai_1  _0700_
timestamp 1685175443
transform -1 0 3264 0 1 31752
box -48 -56 538 834
use sg13g2_mux4_1  _0701_
timestamp 1677257233
transform 1 0 6528 0 -1 30240
box -48 -56 2064 834
use sg13g2_mux4_1  _0702_
timestamp 1677257233
transform 1 0 16896 0 1 24192
box -48 -56 2064 834
use sg13g2_mux4_1  _0703_
timestamp 1677257233
transform 1 0 18432 0 -1 40824
box -48 -56 2064 834
use sg13g2_mux4_1  _0704_
timestamp 1677257233
transform 1 0 17856 0 -1 45360
box -48 -56 2064 834
use sg13g2_mux4_1  _0705_
timestamp 1677257233
transform 1 0 8064 0 -1 27216
box -48 -56 2064 834
use sg13g2_mux4_1  _0706_
timestamp 1677257233
transform 1 0 18240 0 -1 16632
box -48 -56 2064 834
use sg13g2_mux4_1  _0707_
timestamp 1677257233
transform 1 0 18240 0 -1 33264
box -48 -56 2064 834
use sg13g2_mux4_1  _0708_
timestamp 1677257233
transform 1 0 14016 0 1 39312
box -48 -56 2064 834
use sg13g2_mux4_1  _0709_
timestamp 1677257233
transform 1 0 6816 0 1 30240
box -48 -56 2064 834
use sg13g2_mux4_1  _0710_
timestamp 1677257233
transform 1 0 15072 0 1 25704
box -48 -56 2064 834
use sg13g2_mux4_1  _0711_
timestamp 1677257233
transform 1 0 18336 0 -1 37800
box -48 -56 2064 834
use sg13g2_mux4_1  _0712_
timestamp 1677257233
transform 1 0 17856 0 1 42336
box -48 -56 2064 834
use sg13g2_mux4_1  _0713_
timestamp 1677257233
transform 1 0 9216 0 -1 25704
box -48 -56 2064 834
use sg13g2_mux4_1  _0714_
timestamp 1677257233
transform 1 0 18240 0 1 15120
box -48 -56 2064 834
use sg13g2_mux4_1  _0715_
timestamp 1677257233
transform 1 0 14112 0 -1 34776
box -48 -56 2064 834
use sg13g2_mux4_1  _0716_
timestamp 1677257233
transform 1 0 13248 0 -1 46872
box -48 -56 2064 834
use sg13g2_mux4_1  _0717_
timestamp 1677257233
transform 1 0 6912 0 -1 28728
box -48 -56 2064 834
use sg13g2_mux4_1  _0718_
timestamp 1677257233
transform 1 0 16032 0 -1 25704
box -48 -56 2064 834
use sg13g2_mux4_1  _0719_
timestamp 1677257233
transform 1 0 18432 0 -1 36288
box -48 -56 2064 834
use sg13g2_mux4_1  _0720_
timestamp 1677257233
transform 1 0 17664 0 1 45360
box -48 -56 2064 834
use sg13g2_mux4_1  _0721_
timestamp 1677257233
transform 1 0 7392 0 1 25704
box -48 -56 2064 834
use sg13g2_mux4_1  _0722_
timestamp 1677257233
transform 1 0 18240 0 -1 19656
box -48 -56 2064 834
use sg13g2_mux4_1  _0723_
timestamp 1677257233
transform 1 0 18240 0 1 31752
box -48 -56 2064 834
use sg13g2_mux4_1  _0724_
timestamp 1677257233
transform 1 0 14016 0 1 45360
box -48 -56 2064 834
use sg13g2_mux4_1  _0725_
timestamp 1677257233
transform 1 0 6624 0 1 28728
box -48 -56 2064 834
use sg13g2_mux4_1  _0726_
timestamp 1677257233
transform 1 0 15744 0 1 22680
box -48 -56 2064 834
use sg13g2_mux4_1  _0727_
timestamp 1677257233
transform 1 0 18336 0 1 37800
box -48 -56 2064 834
use sg13g2_mux4_1  _0728_
timestamp 1677257233
transform 1 0 17856 0 -1 43848
box -48 -56 2064 834
use sg13g2_mux4_1  _0729_
timestamp 1677257233
transform 1 0 9408 0 1 25704
box -48 -56 2064 834
use sg13g2_mux4_1  _0730_
timestamp 1677257233
transform 1 0 18144 0 1 19656
box -48 -56 2064 834
use sg13g2_mux4_1  _0731_
timestamp 1677257233
transform 1 0 13632 0 1 34776
box -48 -56 2064 834
use sg13g2_mux4_1  _0732_
timestamp 1677257233
transform 1 0 13344 0 -1 45360
box -48 -56 2064 834
use sg13g2_o21ai_1  _0733_
timestamp 1685175443
transform 1 0 3264 0 -1 28728
box -48 -56 538 834
use sg13g2_inv_1  _0734_
timestamp 1676382929
transform -1 0 4896 0 -1 30240
box -48 -56 336 834
use sg13g2_o21ai_1  _0735_
timestamp 1685175443
transform -1 0 4896 0 -1 28728
box -48 -56 538 834
use sg13g2_mux2_1  _0736_
timestamp 1677247768
transform -1 0 5568 0 -1 31752
box -48 -56 1008 834
use sg13g2_a21oi_1  _0737_
timestamp 1683973020
transform 1 0 4416 0 1 30240
box -48 -56 528 834
use sg13g2_nor2_1  _0738_
timestamp 1676627187
transform -1 0 9312 0 -1 30240
box -48 -56 432 834
use sg13g2_o21ai_1  _0739_
timestamp 1685175443
transform 1 0 6048 0 -1 31752
box -48 -56 538 834
use sg13g2_mux2_1  _0740_
timestamp 1677247768
transform 1 0 3456 0 1 28728
box -48 -56 1008 834
use sg13g2_o21ai_1  _0741_
timestamp 1685175443
transform -1 0 3456 0 1 28728
box -48 -56 538 834
use sg13g2_a21oi_1  _0742_
timestamp 1683973020
transform 1 0 3936 0 -1 28728
box -48 -56 528 834
use sg13g2_a21oi_1  _0743_
timestamp 1683973020
transform 1 0 5568 0 -1 31752
box -48 -56 528 834
use sg13g2_o21ai_1  _0744_
timestamp 1685175443
transform -1 0 14976 0 1 21168
box -48 -56 538 834
use sg13g2_inv_1  _0745_
timestamp 1676382929
transform -1 0 14496 0 -1 19656
box -48 -56 336 834
use sg13g2_o21ai_1  _0746_
timestamp 1685175443
transform 1 0 14112 0 1 19656
box -48 -56 538 834
use sg13g2_mux2_1  _0747_
timestamp 1677247768
transform -1 0 16224 0 -1 21168
box -48 -56 1008 834
use sg13g2_a21oi_1  _0748_
timestamp 1683973020
transform -1 0 15456 0 -1 19656
box -48 -56 528 834
use sg13g2_nor2_1  _0749_
timestamp 1676627187
transform 1 0 14496 0 -1 19656
box -48 -56 432 834
use sg13g2_o21ai_1  _0750_
timestamp 1685175443
transform 1 0 14976 0 1 21168
box -48 -56 538 834
use sg13g2_mux2_1  _0751_
timestamp 1677247768
transform 1 0 14592 0 1 19656
box -48 -56 1008 834
use sg13g2_o21ai_1  _0752_
timestamp 1685175443
transform 1 0 15456 0 1 21168
box -48 -56 538 834
use sg13g2_a21oi_1  _0753_
timestamp 1683973020
transform 1 0 15936 0 1 21168
box -48 -56 528 834
use sg13g2_a21oi_1  _0754_
timestamp 1683973020
transform -1 0 16032 0 1 19656
box -48 -56 528 834
use sg13g2_o21ai_1  _0755_
timestamp 1685175443
transform 1 0 17376 0 1 36288
box -48 -56 538 834
use sg13g2_inv_1  _0756_
timestamp 1676382929
transform -1 0 18624 0 1 36288
box -48 -56 336 834
use sg13g2_o21ai_1  _0757_
timestamp 1685175443
transform -1 0 16032 0 -1 36288
box -48 -56 538 834
use sg13g2_mux2_1  _0758_
timestamp 1677247768
transform 1 0 17088 0 1 34776
box -48 -56 1008 834
use sg13g2_a21oi_1  _0759_
timestamp 1683973020
transform 1 0 17856 0 1 36288
box -48 -56 528 834
use sg13g2_nor2_1  _0760_
timestamp 1676627187
transform -1 0 16128 0 1 34776
box -48 -56 432 834
use sg13g2_o21ai_1  _0761_
timestamp 1685175443
transform 1 0 16128 0 1 34776
box -48 -56 538 834
use sg13g2_mux2_1  _0762_
timestamp 1677247768
transform 1 0 16032 0 1 33264
box -48 -56 1008 834
use sg13g2_o21ai_1  _0763_
timestamp 1685175443
transform 1 0 16608 0 1 34776
box -48 -56 538 834
use sg13g2_a21oi_1  _0764_
timestamp 1683973020
transform -1 0 17568 0 -1 34776
box -48 -56 528 834
use sg13g2_a21oi_1  _0765_
timestamp 1683973020
transform 1 0 17664 0 -1 36288
box -48 -56 528 834
use sg13g2_o21ai_1  _0766_
timestamp 1685175443
transform -1 0 15936 0 -1 42336
box -48 -56 538 834
use sg13g2_inv_1  _0767_
timestamp 1676382929
transform -1 0 15552 0 1 40824
box -48 -56 336 834
use sg13g2_o21ai_1  _0768_
timestamp 1685175443
transform -1 0 14880 0 -1 43848
box -48 -56 538 834
use sg13g2_mux2_1  _0769_
timestamp 1677247768
transform 1 0 15168 0 1 43848
box -48 -56 1008 834
use sg13g2_a21oi_1  _0770_
timestamp 1683973020
transform 1 0 15552 0 1 40824
box -48 -56 528 834
use sg13g2_nor2_1  _0771_
timestamp 1676627187
transform -1 0 16224 0 1 42336
box -48 -56 432 834
use sg13g2_o21ai_1  _0772_
timestamp 1685175443
transform 1 0 15360 0 1 42336
box -48 -56 538 834
use sg13g2_mux2_1  _0773_
timestamp 1677247768
transform 1 0 14880 0 -1 43848
box -48 -56 1008 834
use sg13g2_o21ai_1  _0774_
timestamp 1685175443
transform -1 0 15456 0 -1 42336
box -48 -56 538 834
use sg13g2_a21oi_1  _0775_
timestamp 1683973020
transform 1 0 15936 0 -1 42336
box -48 -56 528 834
use sg13g2_a21oi_1  _0776_
timestamp 1683973020
transform -1 0 13728 0 1 42336
box -48 -56 528 834
use sg13g2_o21ai_1  _0777_
timestamp 1685175443
transform -1 0 2976 0 1 28728
box -48 -56 538 834
use sg13g2_inv_1  _0778_
timestamp 1676382929
transform 1 0 3072 0 -1 27216
box -48 -56 336 834
use sg13g2_o21ai_1  _0779_
timestamp 1685175443
transform 1 0 3264 0 1 25704
box -48 -56 538 834
use sg13g2_mux2_1  _0780_
timestamp 1677247768
transform 1 0 3360 0 -1 27216
box -48 -56 1008 834
use sg13g2_a21oi_1  _0781_
timestamp 1683973020
transform 1 0 3744 0 1 25704
box -48 -56 528 834
use sg13g2_nor2_1  _0782_
timestamp 1676627187
transform 1 0 3456 0 1 22680
box -48 -56 432 834
use sg13g2_o21ai_1  _0783_
timestamp 1685175443
transform 1 0 4896 0 1 27216
box -48 -56 538 834
use sg13g2_mux2_1  _0784_
timestamp 1677247768
transform 1 0 3456 0 1 27216
box -48 -56 1008 834
use sg13g2_o21ai_1  _0785_
timestamp 1685175443
transform 1 0 5376 0 1 27216
box -48 -56 538 834
use sg13g2_a21oi_1  _0786_
timestamp 1683973020
transform -1 0 4896 0 1 27216
box -48 -56 528 834
use sg13g2_a21oi_1  _0787_
timestamp 1683973020
transform -1 0 4704 0 1 25704
box -48 -56 528 834
use sg13g2_o21ai_1  _0788_
timestamp 1685175443
transform 1 0 19392 0 -1 22680
box -48 -56 538 834
use sg13g2_inv_1  _0789_
timestamp 1676382929
transform -1 0 20448 0 1 22680
box -48 -56 336 834
use sg13g2_o21ai_1  _0790_
timestamp 1685175443
transform 1 0 18912 0 -1 22680
box -48 -56 538 834
use sg13g2_mux2_1  _0791_
timestamp 1677247768
transform 1 0 19488 0 1 21168
box -48 -56 1008 834
use sg13g2_a21oi_1  _0792_
timestamp 1683973020
transform 1 0 19872 0 -1 24192
box -48 -56 528 834
use sg13g2_nor2_1  _0793_
timestamp 1676627187
transform -1 0 18432 0 1 18144
box -48 -56 432 834
use sg13g2_o21ai_1  _0794_
timestamp 1685175443
transform 1 0 18432 0 -1 22680
box -48 -56 538 834
use sg13g2_mux2_1  _0795_
timestamp 1677247768
transform 1 0 18528 0 1 21168
box -48 -56 1008 834
use sg13g2_o21ai_1  _0796_
timestamp 1685175443
transform 1 0 18912 0 -1 24192
box -48 -56 538 834
use sg13g2_a21oi_1  _0797_
timestamp 1683973020
transform -1 0 19872 0 -1 24192
box -48 -56 528 834
use sg13g2_a21oi_1  _0798_
timestamp 1683973020
transform 1 0 19872 0 -1 22680
box -48 -56 528 834
use sg13g2_o21ai_1  _0799_
timestamp 1685175443
transform -1 0 13728 0 1 30240
box -48 -56 538 834
use sg13g2_inv_1  _0800_
timestamp 1676382929
transform 1 0 12960 0 1 30240
box -48 -56 336 834
use sg13g2_o21ai_1  _0801_
timestamp 1685175443
transform 1 0 14112 0 -1 30240
box -48 -56 538 834
use sg13g2_mux2_1  _0802_
timestamp 1677247768
transform 1 0 14016 0 -1 31752
box -48 -56 1008 834
use sg13g2_a21oi_1  _0803_
timestamp 1683973020
transform 1 0 15072 0 -1 30240
box -48 -56 528 834
use sg13g2_nor2_1  _0804_
timestamp 1676627187
transform 1 0 13248 0 -1 30240
box -48 -56 432 834
use sg13g2_o21ai_1  _0805_
timestamp 1685175443
transform 1 0 13632 0 -1 30240
box -48 -56 538 834
use sg13g2_mux2_1  _0806_
timestamp 1677247768
transform 1 0 13728 0 1 30240
box -48 -56 1008 834
use sg13g2_o21ai_1  _0807_
timestamp 1685175443
transform 1 0 14592 0 -1 30240
box -48 -56 538 834
use sg13g2_a21oi_1  _0808_
timestamp 1683973020
transform 1 0 14976 0 -1 31752
box -48 -56 528 834
use sg13g2_a21oi_1  _0809_
timestamp 1683973020
transform -1 0 14592 0 1 28728
box -48 -56 528 834
use sg13g2_o21ai_1  _0810_
timestamp 1685175443
transform -1 0 12576 0 1 39312
box -48 -56 538 834
use sg13g2_inv_1  _0811_
timestamp 1676382929
transform 1 0 11808 0 1 39312
box -48 -56 336 834
use sg13g2_o21ai_1  _0812_
timestamp 1685175443
transform 1 0 13536 0 1 39312
box -48 -56 538 834
use sg13g2_mux2_1  _0813_
timestamp 1677247768
transform 1 0 13056 0 -1 39312
box -48 -56 1008 834
use sg13g2_a21oi_1  _0814_
timestamp 1683973020
transform 1 0 13824 0 -1 40824
box -48 -56 528 834
use sg13g2_nor2_1  _0815_
timestamp 1676627187
transform -1 0 13056 0 -1 39312
box -48 -56 432 834
use sg13g2_o21ai_1  _0816_
timestamp 1685175443
transform 1 0 12480 0 1 37800
box -48 -56 538 834
use sg13g2_mux2_1  _0817_
timestamp 1677247768
transform 1 0 12576 0 1 39312
box -48 -56 1008 834
use sg13g2_o21ai_1  _0818_
timestamp 1685175443
transform 1 0 12576 0 -1 37800
box -48 -56 538 834
use sg13g2_a21oi_1  _0819_
timestamp 1683973020
transform 1 0 13344 0 -1 40824
box -48 -56 528 834
use sg13g2_a21oi_1  _0820_
timestamp 1683973020
transform 1 0 12864 0 -1 40824
box -48 -56 528 834
use sg13g2_nor2b_1  _0821_
timestamp 1685181386
transform 1 0 4800 0 -1 43848
box -54 -56 528 834
use sg13g2_nand2b_1  _0822_
timestamp 1676567195
transform 1 0 3840 0 1 45360
box -48 -56 528 834
use sg13g2_nand2_1  _0823_
timestamp 1676557249
transform 1 0 5760 0 1 42336
box -48 -56 432 834
use sg13g2_or2_1  _0824_
timestamp 1684236171
transform 1 0 4320 0 1 43848
box -48 -56 528 834
use sg13g2_a21oi_1  _0825_
timestamp 1683973020
transform 1 0 6048 0 -1 45360
box -48 -56 528 834
use sg13g2_nand2_1  _0826_
timestamp 1676557249
transform -1 0 6816 0 1 43848
box -48 -56 432 834
use sg13g2_nand2_1  _0827_
timestamp 1676557249
transform 1 0 4416 0 1 42336
box -48 -56 432 834
use sg13g2_nand4_1  _0828_
timestamp 1685201930
transform 1 0 5280 0 1 43848
box -48 -56 624 834
use sg13g2_a21oi_1  _0829_
timestamp 1683973020
transform 1 0 5280 0 1 42336
box -48 -56 528 834
use sg13g2_o21ai_1  _0830_
timestamp 1685175443
transform 1 0 4320 0 -1 43848
box -48 -56 538 834
use sg13g2_and2_1  _0831_
timestamp 1676901763
transform 1 0 4800 0 1 42336
box -48 -56 528 834
use sg13g2_a21oi_1  _0832_
timestamp 1683973020
transform 1 0 5760 0 -1 43848
box -48 -56 528 834
use sg13g2_a22oi_1  _0833_
timestamp 1685173987
transform 1 0 5856 0 1 43848
box -48 -56 624 834
use sg13g2_nand3_1  _0834_
timestamp 1683988354
transform -1 0 5760 0 -1 43848
box -48 -56 528 834
use sg13g2_nand2b_1  _0835_
timestamp 1676567195
transform 1 0 4800 0 1 43848
box -48 -56 528 834
use sg13g2_or3_1  _0836_
timestamp 1677141922
transform 1 0 4320 0 -1 45360
box -48 -56 720 834
use sg13g2_or2_1  _0837_
timestamp 1684236171
transform 1 0 4800 0 -1 46872
box -48 -56 528 834
use sg13g2_nand4_1  _0838_
timestamp 1685201930
transform 1 0 4992 0 -1 45360
box -48 -56 624 834
use sg13g2_nand2b_1  _0839_
timestamp 1676567195
transform 1 0 6144 0 1 45360
box -48 -56 528 834
use sg13g2_nor3_1  _0840_
timestamp 1676639442
transform 1 0 4320 0 1 45360
box -48 -56 528 834
use sg13g2_a221oi_1  _0841_
timestamp 1685197497
transform 1 0 5376 0 1 45360
box -48 -56 816 834
use sg13g2_a21oi_1  _0842_
timestamp 1683973020
transform 1 0 5568 0 -1 45360
box -48 -56 528 834
use sg13g2_a22oi_1  _0843_
timestamp 1685173987
transform 1 0 4800 0 1 45360
box -48 -56 624 834
use sg13g2_mux4_1  _0844_
timestamp 1677257233
transform 1 0 4896 0 -1 40824
box -48 -56 2064 834
use sg13g2_nand2_1  _0845_
timestamp 1676557249
transform 1 0 5088 0 1 40824
box -48 -56 432 834
use sg13g2_nor2b_1  _0846_
timestamp 1685181386
transform 1 0 5952 0 1 40824
box -54 -56 528 834
use sg13g2_nor3_1  _0847_
timestamp 1676639442
transform -1 0 7392 0 -1 40824
box -48 -56 528 834
use sg13g2_nand2_1  _0848_
timestamp 1676557249
transform -1 0 6912 0 -1 39312
box -48 -56 432 834
use sg13g2_nand2b_1  _0849_
timestamp 1676567195
transform 1 0 5472 0 1 40824
box -48 -56 528 834
use sg13g2_a21oi_1  _0850_
timestamp 1683973020
transform 1 0 6816 0 1 39312
box -48 -56 528 834
use sg13g2_a22oi_1  _0851_
timestamp 1685173987
transform 1 0 5760 0 1 39312
box -48 -56 624 834
use sg13g2_o21ai_1  _0852_
timestamp 1685175443
transform 1 0 7392 0 -1 40824
box -48 -56 538 834
use sg13g2_nor3_1  _0853_
timestamp 1676639442
transform 1 0 4800 0 1 39312
box -48 -56 528 834
use sg13g2_nor3_1  _0854_
timestamp 1676639442
transform -1 0 7392 0 1 37800
box -48 -56 528 834
use sg13g2_o21ai_1  _0855_
timestamp 1685175443
transform 1 0 5280 0 1 39312
box -48 -56 538 834
use sg13g2_nor3_1  _0856_
timestamp 1676639442
transform 1 0 5472 0 1 37800
box -48 -56 528 834
use sg13g2_a21oi_1  _0857_
timestamp 1683973020
transform 1 0 6336 0 1 39312
box -48 -56 528 834
use sg13g2_a21oi_1  _0858_
timestamp 1683973020
transform 1 0 6432 0 1 40824
box -48 -56 528 834
use sg13g2_nor3_1  _0859_
timestamp 1676639442
transform -1 0 6432 0 1 37800
box -48 -56 528 834
use sg13g2_nor3_1  _0860_
timestamp 1676639442
transform -1 0 6528 0 -1 39312
box -48 -56 528 834
use sg13g2_o21ai_1  _0861_
timestamp 1685175443
transform -1 0 5472 0 1 37800
box -48 -56 538 834
use sg13g2_o21ai_1  _0862_
timestamp 1685175443
transform 1 0 6432 0 1 37800
box -48 -56 538 834
use sg13g2_dlhq_1  _0863_
timestamp 1678805552
transform 1 0 1536 0 -1 81648
box -50 -56 1692 834
use sg13g2_dlhq_1  _0864_
timestamp 1678805552
transform -1 0 7104 0 -1 78624
box -50 -56 1692 834
use sg13g2_dlhq_1  _0865_
timestamp 1678805552
transform 1 0 11040 0 1 78624
box -50 -56 1692 834
use sg13g2_dlhq_1  _0866_
timestamp 1678805552
transform 1 0 10464 0 -1 78624
box -50 -56 1692 834
use sg13g2_dlhq_1  _0867_
timestamp 1678805552
transform 1 0 17568 0 1 72576
box -50 -56 1692 834
use sg13g2_dlhq_1  _0868_
timestamp 1678805552
transform 1 0 15936 0 1 72576
box -50 -56 1692 834
use sg13g2_dlhq_1  _0869_
timestamp 1678805552
transform 1 0 9792 0 -1 57456
box -50 -56 1692 834
use sg13g2_dlhq_1  _0870_
timestamp 1678805552
transform 1 0 9792 0 1 57456
box -50 -56 1692 834
use sg13g2_dlhq_1  _0871_
timestamp 1678805552
transform 1 0 7680 0 -1 49896
box -50 -56 1692 834
use sg13g2_dlhq_1  _0872_
timestamp 1678805552
transform 1 0 8832 0 -1 51408
box -50 -56 1692 834
use sg13g2_dlhq_1  _0873_
timestamp 1678805552
transform 1 0 14112 0 1 49896
box -50 -56 1692 834
use sg13g2_dlhq_1  _0874_
timestamp 1678805552
transform 1 0 12480 0 1 49896
box -50 -56 1692 834
use sg13g2_dlhq_1  _0875_
timestamp 1678805552
transform 1 0 17568 0 -1 51408
box -50 -56 1692 834
use sg13g2_dlhq_1  _0876_
timestamp 1678805552
transform 1 0 18144 0 1 51408
box -50 -56 1692 834
use sg13g2_dlhq_1  _0877_
timestamp 1678805552
transform 1 0 2016 0 1 49896
box -50 -56 1692 834
use sg13g2_dlhq_1  _0878_
timestamp 1678805552
transform -1 0 5568 0 -1 49896
box -50 -56 1692 834
use sg13g2_dlhq_1  _0879_
timestamp 1678805552
transform 1 0 3936 0 1 49896
box -50 -56 1692 834
use sg13g2_dlhq_1  _0880_
timestamp 1678805552
transform 1 0 1920 0 -1 49896
box -50 -56 1692 834
use sg13g2_dlhq_1  _0881_
timestamp 1678805552
transform 1 0 11904 0 -1 49896
box -50 -56 1692 834
use sg13g2_dlhq_1  _0882_
timestamp 1678805552
transform 1 0 10464 0 -1 51408
box -50 -56 1692 834
use sg13g2_dlhq_1  _0883_
timestamp 1678805552
transform 1 0 14784 0 1 51408
box -50 -56 1692 834
use sg13g2_dlhq_1  _0884_
timestamp 1678805552
transform -1 0 18048 0 1 51408
box -50 -56 1692 834
use sg13g2_dlhq_1  _0885_
timestamp 1678805552
transform -1 0 8544 0 1 48384
box -50 -56 1692 834
use sg13g2_dlhq_1  _0886_
timestamp 1678805552
transform -1 0 7680 0 -1 49896
box -50 -56 1692 834
use sg13g2_dlhq_1  _0887_
timestamp 1678805552
transform 1 0 8544 0 1 74088
box -50 -56 1692 834
use sg13g2_dlhq_1  _0888_
timestamp 1678805552
transform 1 0 1344 0 -1 77112
box -50 -56 1692 834
use sg13g2_dlhq_1  _0889_
timestamp 1678805552
transform 1 0 8544 0 -1 83160
box -50 -56 1692 834
use sg13g2_dlhq_1  _0890_
timestamp 1678805552
transform 1 0 9216 0 1 81648
box -50 -56 1692 834
use sg13g2_dlhq_1  _0891_
timestamp 1678805552
transform 1 0 17472 0 1 68040
box -50 -56 1692 834
use sg13g2_dlhq_1  _0892_
timestamp 1678805552
transform 1 0 16032 0 -1 71064
box -50 -56 1692 834
use sg13g2_dlhq_1  _0893_
timestamp 1678805552
transform -1 0 10368 0 1 58968
box -50 -56 1692 834
use sg13g2_dlhq_1  _0894_
timestamp 1678805552
transform 1 0 6720 0 -1 58968
box -50 -56 1692 834
use sg13g2_dlhq_1  _0895_
timestamp 1678805552
transform 1 0 1632 0 1 80136
box -50 -56 1692 834
use sg13g2_dlhq_1  _0896_
timestamp 1678805552
transform 1 0 1440 0 -1 80136
box -50 -56 1692 834
use sg13g2_dlhq_1  _0897_
timestamp 1678805552
transform 1 0 8736 0 -1 86184
box -50 -56 1692 834
use sg13g2_dlhq_1  _0898_
timestamp 1678805552
transform 1 0 8928 0 1 84672
box -50 -56 1692 834
use sg13g2_dlhq_1  _0899_
timestamp 1678805552
transform 1 0 18528 0 -1 74088
box -50 -56 1692 834
use sg13g2_dlhq_1  _0900_
timestamp 1678805552
transform 1 0 16320 0 -1 74088
box -50 -56 1692 834
use sg13g2_dlhq_1  _0901_
timestamp 1678805552
transform -1 0 12192 0 -1 55944
box -50 -56 1692 834
use sg13g2_dlhq_1  _0902_
timestamp 1678805552
transform 1 0 7776 0 1 54432
box -50 -56 1692 834
use sg13g2_dlhq_1  _0903_
timestamp 1678805552
transform 1 0 3840 0 1 78624
box -50 -56 1692 834
use sg13g2_dlhq_1  _0904_
timestamp 1678805552
transform 1 0 1440 0 1 81648
box -50 -56 1692 834
use sg13g2_dlhq_1  _0905_
timestamp 1678805552
transform 1 0 5088 0 1 81648
box -50 -56 1692 834
use sg13g2_dlhq_1  _0906_
timestamp 1678805552
transform 1 0 9024 0 -1 81648
box -50 -56 1692 834
use sg13g2_dlhq_1  _0907_
timestamp 1678805552
transform 1 0 18816 0 -1 75600
box -50 -56 1692 834
use sg13g2_dlhq_1  _0908_
timestamp 1678805552
transform 1 0 18144 0 -1 77112
box -50 -56 1692 834
use sg13g2_dlhq_1  _0909_
timestamp 1678805552
transform 1 0 8448 0 1 55944
box -50 -56 1692 834
use sg13g2_dlhq_1  _0910_
timestamp 1678805552
transform 1 0 6528 0 -1 55944
box -50 -56 1692 834
use sg13g2_dlhq_1  _0911_
timestamp 1678805552
transform 1 0 3744 0 1 77112
box -50 -56 1692 834
use sg13g2_dlhq_1  _0912_
timestamp 1678805552
transform 1 0 1536 0 1 78624
box -50 -56 1692 834
use sg13g2_dlhq_1  _0913_
timestamp 1678805552
transform 1 0 9504 0 1 83160
box -50 -56 1692 834
use sg13g2_dlhq_1  _0914_
timestamp 1678805552
transform 1 0 9216 0 -1 84672
box -50 -56 1692 834
use sg13g2_dlhq_1  _0915_
timestamp 1678805552
transform 1 0 18720 0 -1 71064
box -50 -56 1692 834
use sg13g2_dlhq_1  _0916_
timestamp 1678805552
transform 1 0 16512 0 -1 69552
box -50 -56 1692 834
use sg13g2_dlhq_1  _0917_
timestamp 1678805552
transform -1 0 12864 0 -1 54432
box -50 -56 1692 834
use sg13g2_dlhq_1  _0918_
timestamp 1678805552
transform 1 0 7392 0 1 49896
box -50 -56 1692 834
use sg13g2_dlhq_1  _0919_
timestamp 1678805552
transform 1 0 5856 0 -1 69552
box -50 -56 1692 834
use sg13g2_dlhq_1  _0920_
timestamp 1678805552
transform 1 0 5280 0 1 69552
box -50 -56 1692 834
use sg13g2_dlhq_1  _0921_
timestamp 1678805552
transform 1 0 1344 0 1 54432
box -50 -56 1692 834
use sg13g2_dlhq_1  _0922_
timestamp 1678805552
transform 1 0 1344 0 -1 55944
box -50 -56 1692 834
use sg13g2_dlhq_1  _0923_
timestamp 1678805552
transform 1 0 11040 0 -1 87696
box -50 -56 1692 834
use sg13g2_dlhq_1  _0924_
timestamp 1678805552
transform 1 0 10752 0 1 86184
box -50 -56 1692 834
use sg13g2_dlhq_1  _0925_
timestamp 1678805552
transform 1 0 16128 0 -1 77112
box -50 -56 1692 834
use sg13g2_dlhq_1  _0926_
timestamp 1678805552
transform 1 0 15648 0 1 75600
box -50 -56 1692 834
use sg13g2_dlhq_1  _0927_
timestamp 1678805552
transform 1 0 6528 0 -1 77112
box -50 -56 1692 834
use sg13g2_dlhq_1  _0928_
timestamp 1678805552
transform -1 0 8928 0 1 77112
box -50 -56 1692 834
use sg13g2_dlhq_1  _0929_
timestamp 1678805552
transform 1 0 4320 0 -1 86184
box -50 -56 1692 834
use sg13g2_dlhq_1  _0930_
timestamp 1678805552
transform 1 0 2880 0 1 86184
box -50 -56 1692 834
use sg13g2_dlhq_1  _0931_
timestamp 1678805552
transform 1 0 15360 0 -1 86184
box -50 -56 1692 834
use sg13g2_dlhq_1  _0932_
timestamp 1678805552
transform 1 0 13728 0 -1 86184
box -50 -56 1692 834
use sg13g2_dlhq_1  _0933_
timestamp 1678805552
transform 1 0 12384 0 1 57456
box -50 -56 1692 834
use sg13g2_dlhq_1  _0934_
timestamp 1678805552
transform 1 0 11904 0 1 54432
box -50 -56 1692 834
use sg13g2_dlhq_1  _0935_
timestamp 1678805552
transform 1 0 4800 0 1 52920
box -50 -56 1692 834
use sg13g2_dlhq_1  _0936_
timestamp 1678805552
transform 1 0 3552 0 -1 52920
box -50 -56 1692 834
use sg13g2_dlhq_1  _0937_
timestamp 1678805552
transform 1 0 1440 0 -1 83160
box -50 -56 1692 834
use sg13g2_dlhq_1  _0938_
timestamp 1678805552
transform 1 0 1440 0 1 83160
box -50 -56 1692 834
use sg13g2_dlhq_1  _0939_
timestamp 1678805552
transform -1 0 16608 0 1 89208
box -50 -56 1692 834
use sg13g2_dlhq_1  _0940_
timestamp 1678805552
transform 1 0 11328 0 -1 90720
box -50 -56 1692 834
use sg13g2_dlhq_1  _0941_
timestamp 1678805552
transform 1 0 16800 0 -1 89208
box -50 -56 1692 834
use sg13g2_dlhq_1  _0942_
timestamp 1678805552
transform 1 0 15648 0 -1 87696
box -50 -56 1692 834
use sg13g2_dlhq_1  _0943_
timestamp 1678805552
transform 1 0 9792 0 -1 66528
box -50 -56 1692 834
use sg13g2_dlhq_1  _0944_
timestamp 1678805552
transform 1 0 7872 0 -1 66528
box -50 -56 1692 834
use sg13g2_dlhq_1  _0945_
timestamp 1678805552
transform 1 0 4416 0 -1 89208
box -50 -56 1692 834
use sg13g2_dlhq_1  _0946_
timestamp 1678805552
transform 1 0 2688 0 1 87696
box -50 -56 1692 834
use sg13g2_dlhq_1  _0947_
timestamp 1678805552
transform 1 0 18528 0 -1 86184
box -50 -56 1692 834
use sg13g2_dlhq_1  _0948_
timestamp 1678805552
transform 1 0 16992 0 1 84672
box -50 -56 1692 834
use sg13g2_dlhq_1  _0949_
timestamp 1678805552
transform 1 0 15264 0 1 54432
box -50 -56 1692 834
use sg13g2_dlhq_1  _0950_
timestamp 1678805552
transform 1 0 13536 0 1 54432
box -50 -56 1692 834
use sg13g2_dlhq_1  _0951_
timestamp 1678805552
transform 1 0 6144 0 1 54432
box -50 -56 1692 834
use sg13g2_dlhq_1  _0952_
timestamp 1678805552
transform 1 0 4224 0 1 54432
box -50 -56 1692 834
use sg13g2_dlhq_1  _0953_
timestamp 1678805552
transform -1 0 6720 0 -1 83160
box -50 -56 1692 834
use sg13g2_dlhq_1  _0954_
timestamp 1678805552
transform 1 0 1344 0 1 84672
box -50 -56 1692 834
use sg13g2_dlhq_1  _0955_
timestamp 1678805552
transform 1 0 10752 0 -1 89208
box -50 -56 1692 834
use sg13g2_dlhq_1  _0956_
timestamp 1678805552
transform 1 0 10656 0 1 87696
box -50 -56 1692 834
use sg13g2_dlhq_1  _0957_
timestamp 1678805552
transform 1 0 18624 0 1 84672
box -50 -56 1692 834
use sg13g2_dlhq_1  _0958_
timestamp 1678805552
transform -1 0 20064 0 -1 83160
box -50 -56 1692 834
use sg13g2_dlhq_1  _0959_
timestamp 1678805552
transform 1 0 9984 0 1 60480
box -50 -56 1692 834
use sg13g2_dlhq_1  _0960_
timestamp 1678805552
transform 1 0 7872 0 -1 61992
box -50 -56 1692 834
use sg13g2_dlhq_1  _0961_
timestamp 1678805552
transform -1 0 10464 0 -1 87696
box -50 -56 1692 834
use sg13g2_dlhq_1  _0962_
timestamp 1678805552
transform -1 0 8640 0 -1 89208
box -50 -56 1692 834
use sg13g2_dlhq_1  _0963_
timestamp 1678805552
transform 1 0 15456 0 1 86184
box -50 -56 1692 834
use sg13g2_dlhq_1  _0964_
timestamp 1678805552
transform 1 0 13824 0 1 86184
box -50 -56 1692 834
use sg13g2_dlhq_1  _0965_
timestamp 1678805552
transform 1 0 11520 0 1 55944
box -50 -56 1692 834
use sg13g2_dlhq_1  _0966_
timestamp 1678805552
transform 1 0 11424 0 -1 57456
box -50 -56 1692 834
use sg13g2_dlhq_1  _0967_
timestamp 1678805552
transform 1 0 6048 0 -1 51408
box -50 -56 1692 834
use sg13g2_dlhq_1  _0968_
timestamp 1678805552
transform 1 0 4416 0 -1 51408
box -50 -56 1692 834
use sg13g2_dlhq_1  _0969_
timestamp 1678805552
transform 1 0 3360 0 1 84672
box -50 -56 1692 834
use sg13g2_dlhq_1  _0970_
timestamp 1678805552
transform 1 0 1536 0 -1 87696
box -50 -56 1692 834
use sg13g2_dlhq_1  _0971_
timestamp 1678805552
transform 1 0 14304 0 -1 90720
box -50 -56 1692 834
use sg13g2_dlhq_1  _0972_
timestamp 1678805552
transform 1 0 11328 0 1 89208
box -50 -56 1692 834
use sg13g2_dlhq_1  _0973_
timestamp 1678805552
transform 1 0 16800 0 1 89208
box -50 -56 1692 834
use sg13g2_dlhq_1  _0974_
timestamp 1678805552
transform 1 0 16512 0 1 87696
box -50 -56 1692 834
use sg13g2_dlhq_1  _0975_
timestamp 1678805552
transform 1 0 9408 0 1 66528
box -50 -56 1692 834
use sg13g2_dlhq_1  _0976_
timestamp 1678805552
transform 1 0 7680 0 1 65016
box -50 -56 1692 834
use sg13g2_dlhq_1  _0977_
timestamp 1678805552
transform 1 0 4608 0 1 89208
box -50 -56 1692 834
use sg13g2_dlhq_1  _0978_
timestamp 1678805552
transform 1 0 2688 0 -1 89208
box -50 -56 1692 834
use sg13g2_dlhq_1  _0979_
timestamp 1678805552
transform 1 0 18528 0 1 87696
box -50 -56 1692 834
use sg13g2_dlhq_1  _0980_
timestamp 1678805552
transform 1 0 16032 0 1 83160
box -50 -56 1692 834
use sg13g2_dlhq_1  _0981_
timestamp 1678805552
transform 1 0 15264 0 -1 57456
box -50 -56 1692 834
use sg13g2_dlhq_1  _0982_
timestamp 1678805552
transform 1 0 13536 0 -1 55944
box -50 -56 1692 834
use sg13g2_dlhq_1  _0983_
timestamp 1678805552
transform -1 0 9408 0 1 51408
box -50 -56 1692 834
use sg13g2_dlhq_1  _0984_
timestamp 1678805552
transform 1 0 4416 0 -1 54432
box -50 -56 1692 834
use sg13g2_dlhq_1  _0985_
timestamp 1678805552
transform 1 0 1632 0 -1 86184
box -50 -56 1692 834
use sg13g2_dlhq_1  _0986_
timestamp 1678805552
transform 1 0 1248 0 1 86184
box -50 -56 1692 834
use sg13g2_dlhq_1  _0987_
timestamp 1678805552
transform -1 0 16512 0 1 87696
box -50 -56 1692 834
use sg13g2_dlhq_1  _0988_
timestamp 1678805552
transform -1 0 10656 0 1 87696
box -50 -56 1692 834
use sg13g2_dlhq_1  _0989_
timestamp 1678805552
transform 1 0 16416 0 1 78624
box -50 -56 1692 834
use sg13g2_dlhq_1  _0990_
timestamp 1678805552
transform 1 0 16800 0 -1 83160
box -50 -56 1692 834
use sg13g2_dlhq_1  _0991_
timestamp 1678805552
transform 1 0 10272 0 -1 63504
box -50 -56 1692 834
use sg13g2_dlhq_1  _0992_
timestamp 1678805552
transform 1 0 9984 0 1 63504
box -50 -56 1692 834
use sg13g2_dlhq_1  _0993_
timestamp 1678805552
transform 1 0 4416 0 1 65016
box -50 -56 1692 834
use sg13g2_dlhq_1  _0994_
timestamp 1678805552
transform 1 0 5856 0 -1 61992
box -50 -56 1692 834
use sg13g2_dlhq_1  _0995_
timestamp 1678805552
transform 1 0 14976 0 1 60480
box -50 -56 1692 834
use sg13g2_dlhq_1  _0996_
timestamp 1678805552
transform 1 0 16608 0 1 60480
box -50 -56 1692 834
use sg13g2_dlhq_1  _0997_
timestamp 1678805552
transform 1 0 12672 0 1 69552
box -50 -56 1692 834
use sg13g2_dlhq_1  _0998_
timestamp 1678805552
transform 1 0 14400 0 1 69552
box -50 -56 1692 834
use sg13g2_dlhq_1  _0999_
timestamp 1678805552
transform 1 0 4896 0 1 72576
box -50 -56 1692 834
use sg13g2_dlhq_1  _1000_
timestamp 1678805552
transform 1 0 6624 0 1 71064
box -50 -56 1692 834
use sg13g2_dlhq_1  _1001_
timestamp 1678805552
transform 1 0 4032 0 -1 60480
box -50 -56 1692 834
use sg13g2_dlhq_1  _1002_
timestamp 1678805552
transform 1 0 1632 0 -1 63504
box -50 -56 1692 834
use sg13g2_dlhq_1  _1003_
timestamp 1678805552
transform 1 0 18624 0 1 65016
box -50 -56 1692 834
use sg13g2_dlhq_1  _1004_
timestamp 1678805552
transform 1 0 16320 0 1 66528
box -50 -56 1692 834
use sg13g2_dlhq_1  _1005_
timestamp 1678805552
transform 1 0 12960 0 -1 66528
box -50 -56 1692 834
use sg13g2_dlhq_1  _1006_
timestamp 1678805552
transform -1 0 18624 0 1 65016
box -50 -56 1692 834
use sg13g2_dlhq_1  _1007_
timestamp 1678805552
transform 1 0 4608 0 -1 75600
box -50 -56 1692 834
use sg13g2_dlhq_1  _1008_
timestamp 1678805552
transform 1 0 5088 0 -1 74088
box -50 -56 1692 834
use sg13g2_dlhq_1  _1009_
timestamp 1678805552
transform 1 0 4704 0 -1 66528
box -50 -56 1692 834
use sg13g2_dlhq_1  _1010_
timestamp 1678805552
transform 1 0 1248 0 -1 68040
box -50 -56 1692 834
use sg13g2_dlhq_1  _1011_
timestamp 1678805552
transform 1 0 16512 0 1 81648
box -50 -56 1692 834
use sg13g2_dlhq_1  _1012_
timestamp 1678805552
transform 1 0 14880 0 1 80136
box -50 -56 1692 834
use sg13g2_dlhq_1  _1013_
timestamp 1678805552
transform 1 0 15168 0 -1 72576
box -50 -56 1692 834
use sg13g2_dlhq_1  _1014_
timestamp 1678805552
transform 1 0 13728 0 -1 71064
box -50 -56 1692 834
use sg13g2_dlhq_1  _1015_
timestamp 1678805552
transform 1 0 8352 0 -1 69552
box -50 -56 1692 834
use sg13g2_dlhq_1  _1016_
timestamp 1678805552
transform 1 0 5280 0 1 66528
box -50 -56 1692 834
use sg13g2_dlhq_1  _1017_
timestamp 1678805552
transform 1 0 5760 0 -1 60480
box -50 -56 1692 834
use sg13g2_dlhq_1  _1018_
timestamp 1678805552
transform 1 0 4032 0 1 58968
box -50 -56 1692 834
use sg13g2_dlhq_1  _1019_
timestamp 1678805552
transform 1 0 18528 0 -1 57456
box -50 -56 1692 834
use sg13g2_dlhq_1  _1020_
timestamp 1678805552
transform 1 0 16896 0 -1 57456
box -50 -56 1692 834
use sg13g2_dlhq_1  _1021_
timestamp 1678805552
transform 1 0 11424 0 -1 69552
box -50 -56 1692 834
use sg13g2_dlhq_1  _1022_
timestamp 1678805552
transform 1 0 10368 0 1 68040
box -50 -56 1692 834
use sg13g2_dlhq_1  _1023_
timestamp 1678805552
transform 1 0 1248 0 -1 74088
box -50 -56 1692 834
use sg13g2_dlhq_1  _1024_
timestamp 1678805552
transform 1 0 1152 0 1 74088
box -50 -56 1692 834
use sg13g2_dlhq_1  _1025_
timestamp 1678805552
transform 1 0 3840 0 1 63504
box -50 -56 1692 834
use sg13g2_dlhq_1  _1026_
timestamp 1678805552
transform 1 0 1440 0 1 65016
box -50 -56 1692 834
use sg13g2_dlhq_1  _1027_
timestamp 1678805552
transform 1 0 18528 0 1 60480
box -50 -56 1692 834
use sg13g2_dlhq_1  _1028_
timestamp 1678805552
transform 1 0 16608 0 1 61992
box -50 -56 1692 834
use sg13g2_dlhq_1  _1029_
timestamp 1678805552
transform 1 0 14592 0 -1 65016
box -50 -56 1692 834
use sg13g2_dlhq_1  _1030_
timestamp 1678805552
transform 1 0 13536 0 1 66528
box -50 -56 1692 834
use sg13g2_dlhq_1  _1031_
timestamp 1678805552
transform 1 0 4704 0 1 71064
box -50 -56 1692 834
use sg13g2_dlhq_1  _1032_
timestamp 1678805552
transform 1 0 2880 0 1 72576
box -50 -56 1692 834
use sg13g2_dlhq_1  _1033_
timestamp 1678805552
transform 1 0 4128 0 -1 58968
box -50 -56 1692 834
use sg13g2_dlhq_1  _1034_
timestamp 1678805552
transform 1 0 1440 0 1 57456
box -50 -56 1692 834
use sg13g2_dlhq_1  _1035_
timestamp 1678805552
transform 1 0 18624 0 -1 60480
box -50 -56 1692 834
use sg13g2_dlhq_1  _1036_
timestamp 1678805552
transform 1 0 16608 0 1 58968
box -50 -56 1692 834
use sg13g2_dlhq_1  _1037_
timestamp 1678805552
transform 1 0 12576 0 -1 65016
box -50 -56 1692 834
use sg13g2_dlhq_1  _1038_
timestamp 1678805552
transform 1 0 12000 0 1 61992
box -50 -56 1692 834
use sg13g2_dlhq_1  _1039_
timestamp 1678805552
transform -1 0 7296 0 1 68040
box -50 -56 1692 834
use sg13g2_dlhq_1  _1040_
timestamp 1678805552
transform 1 0 1440 0 1 69552
box -50 -56 1692 834
use sg13g2_dlhq_1  _1041_
timestamp 1678805552
transform -1 0 7008 0 1 57456
box -50 -56 1692 834
use sg13g2_dlhq_1  _1042_
timestamp 1678805552
transform 1 0 2688 0 -1 57456
box -50 -56 1692 834
use sg13g2_dlhq_1  _1043_
timestamp 1678805552
transform 1 0 18624 0 -1 58968
box -50 -56 1692 834
use sg13g2_dlhq_1  _1044_
timestamp 1678805552
transform 1 0 16512 0 1 57456
box -50 -56 1692 834
use sg13g2_dlhq_1  _1045_
timestamp 1678805552
transform 1 0 14688 0 -1 68040
box -50 -56 1692 834
use sg13g2_dlhq_1  _1046_
timestamp 1678805552
transform 1 0 12672 0 -1 68040
box -50 -56 1692 834
use sg13g2_dlhq_1  _1047_
timestamp 1678805552
transform 1 0 1920 0 -1 71064
box -50 -56 1692 834
use sg13g2_dlhq_1  _1048_
timestamp 1678805552
transform 1 0 1248 0 1 72576
box -50 -56 1692 834
use sg13g2_dlhq_1  _1049_
timestamp 1678805552
transform 1 0 1536 0 1 58968
box -50 -56 1692 834
use sg13g2_dlhq_1  _1050_
timestamp 1678805552
transform 1 0 1152 0 1 60480
box -50 -56 1692 834
use sg13g2_dlhq_1  _1051_
timestamp 1678805552
transform 1 0 17952 0 -1 55944
box -50 -56 1692 834
use sg13g2_dlhq_1  _1052_
timestamp 1678805552
transform 1 0 16992 0 1 54432
box -50 -56 1692 834
use sg13g2_dlhq_1  _1053_
timestamp 1678805552
transform -1 0 17280 0 -1 63504
box -50 -56 1692 834
use sg13g2_dlhq_1  _1054_
timestamp 1678805552
transform 1 0 13728 0 -1 61992
box -50 -56 1692 834
use sg13g2_dlhq_1  _1055_
timestamp 1678805552
transform 1 0 2592 0 -1 75600
box -50 -56 1692 834
use sg13g2_dlhq_1  _1056_
timestamp 1678805552
transform 1 0 1152 0 1 75600
box -50 -56 1692 834
use sg13g2_dlhq_1  _1057_
timestamp 1678805552
transform 1 0 3840 0 -1 63504
box -50 -56 1692 834
use sg13g2_dlhq_1  _1058_
timestamp 1678805552
transform 1 0 1440 0 1 63504
box -50 -56 1692 834
use sg13g2_dlhq_1  _1059_
timestamp 1678805552
transform 1 0 18240 0 -1 65016
box -50 -56 1692 834
use sg13g2_dlhq_1  _1060_
timestamp 1678805552
transform 1 0 16320 0 1 63504
box -50 -56 1692 834
use sg13g2_dlhq_1  _1061_
timestamp 1678805552
transform 1 0 13728 0 1 52920
box -50 -56 1692 834
use sg13g2_dlhq_1  _1062_
timestamp 1678805552
transform 1 0 13344 0 -1 54432
box -50 -56 1692 834
use sg13g2_dlhq_1  _1063_
timestamp 1678805552
transform -1 0 4896 0 1 66528
box -50 -56 1692 834
use sg13g2_dlhq_1  _1064_
timestamp 1678805552
transform 1 0 1152 0 1 68040
box -50 -56 1692 834
use sg13g2_dlhq_1  _1065_
timestamp 1678805552
transform 1 0 1632 0 -1 61992
box -50 -56 1692 834
use sg13g2_dlhq_1  _1066_
timestamp 1678805552
transform 1 0 1152 0 1 61992
box -50 -56 1692 834
use sg13g2_dlhq_1  _1067_
timestamp 1678805552
transform 1 0 18816 0 1 54432
box -50 -56 1692 834
use sg13g2_dlhq_1  _1068_
timestamp 1678805552
transform 1 0 17376 0 -1 52920
box -50 -56 1692 834
use sg13g2_dlhq_1  _1069_
timestamp 1678805552
transform 1 0 12672 0 1 63504
box -50 -56 1692 834
use sg13g2_dlhq_1  _1070_
timestamp 1678805552
transform 1 0 12096 0 -1 61992
box -50 -56 1692 834
use sg13g2_dlhq_1  _1071_
timestamp 1678805552
transform -1 0 5280 0 1 69552
box -50 -56 1692 834
use sg13g2_dlhq_1  _1072_
timestamp 1678805552
transform 1 0 1344 0 -1 69552
box -50 -56 1692 834
use sg13g2_dlhq_1  _1073_
timestamp 1678805552
transform 1 0 3840 0 -1 55944
box -50 -56 1692 834
use sg13g2_dlhq_1  _1074_
timestamp 1678805552
transform 1 0 1632 0 1 55944
box -50 -56 1692 834
use sg13g2_dlhq_1  _1075_
timestamp 1678805552
transform 1 0 18336 0 1 61992
box -50 -56 1692 834
use sg13g2_dlhq_1  _1076_
timestamp 1678805552
transform 1 0 16512 0 -1 65016
box -50 -56 1692 834
use sg13g2_dlhq_1  _1077_
timestamp 1678805552
transform 1 0 15744 0 -1 52920
box -50 -56 1692 834
use sg13g2_dlhq_1  _1078_
timestamp 1678805552
transform 1 0 14112 0 -1 52920
box -50 -56 1692 834
use sg13g2_dlhq_1  _1079_
timestamp 1678805552
transform 1 0 1632 0 1 66528
box -50 -56 1692 834
use sg13g2_dlhq_1  _1080_
timestamp 1678805552
transform -1 0 7104 0 -1 63504
box -50 -56 1692 834
use sg13g2_dlhq_1  _1081_
timestamp 1678805552
transform 1 0 1152 0 -1 78624
box -50 -56 1692 834
use sg13g2_dlhq_1  _1082_
timestamp 1678805552
transform 1 0 2112 0 1 77112
box -50 -56 1692 834
use sg13g2_dlhq_1  _1083_
timestamp 1678805552
transform 1 0 9408 0 -1 68040
box -50 -56 1692 834
use sg13g2_dlhq_1  _1084_
timestamp 1678805552
transform 1 0 11040 0 -1 68040
box -50 -56 1692 834
use sg13g2_dlhq_1  _1085_
timestamp 1678805552
transform 1 0 16896 0 -1 68040
box -50 -56 1692 834
use sg13g2_dlhq_1  _1086_
timestamp 1678805552
transform 1 0 18528 0 -1 68040
box -50 -56 1692 834
use sg13g2_dlhq_1  _1087_
timestamp 1678805552
transform 1 0 9024 0 -1 60480
box -50 -56 1692 834
use sg13g2_dlhq_1  _1088_
timestamp 1678805552
transform 1 0 10656 0 -1 60480
box -50 -56 1692 834
use sg13g2_dlhq_1  _1089_
timestamp 1678805552
transform 1 0 5952 0 1 83160
box -50 -56 1692 834
use sg13g2_dlhq_1  _1090_
timestamp 1678805552
transform 1 0 5184 0 1 84672
box -50 -56 1692 834
use sg13g2_dlhq_1  _1091_
timestamp 1678805552
transform 1 0 6912 0 -1 83160
box -50 -56 1692 834
use sg13g2_dlhq_1  _1092_
timestamp 1678805552
transform 1 0 13440 0 -1 81648
box -50 -56 1692 834
use sg13g2_dlhq_1  _1093_
timestamp 1678805552
transform 1 0 10656 0 1 80136
box -50 -56 1692 834
use sg13g2_dlhq_1  _1094_
timestamp 1678805552
transform 1 0 13152 0 1 80136
box -50 -56 1692 834
use sg13g2_dlhq_1  _1095_
timestamp 1678805552
transform 1 0 14784 0 1 58968
box -50 -56 1692 834
use sg13g2_dlhq_1  _1096_
timestamp 1678805552
transform 1 0 13152 0 1 58968
box -50 -56 1692 834
use sg13g2_dlhq_1  _1097_
timestamp 1678805552
transform 1 0 13536 0 -1 58968
box -50 -56 1692 834
use sg13g2_dlhq_1  _1098_
timestamp 1678805552
transform -1 0 12480 0 1 51408
box -50 -56 1692 834
use sg13g2_dlhq_1  _1099_
timestamp 1678805552
transform -1 0 14112 0 -1 52920
box -50 -56 1692 834
use sg13g2_dlhq_1  _1100_
timestamp 1678805552
transform -1 0 12480 0 -1 52920
box -50 -56 1692 834
use sg13g2_dlhq_1  _1101_
timestamp 1678805552
transform 1 0 7200 0 -1 78624
box -50 -56 1692 834
use sg13g2_dlhq_1  _1102_
timestamp 1678805552
transform 1 0 5760 0 1 78624
box -50 -56 1692 834
use sg13g2_dlhq_1  _1103_
timestamp 1678805552
transform 1 0 10176 0 1 74088
box -50 -56 1692 834
use sg13g2_dlhq_1  _1104_
timestamp 1678805552
transform 1 0 9216 0 -1 75600
box -50 -56 1692 834
use sg13g2_dlhq_1  _1105_
timestamp 1678805552
transform 1 0 11904 0 1 74088
box -50 -56 1692 834
use sg13g2_dlhq_1  _1106_
timestamp 1678805552
transform 1 0 10560 0 -1 74088
box -50 -56 1692 834
use sg13g2_dlhq_1  _1107_
timestamp 1678805552
transform -1 0 14784 0 1 51408
box -50 -56 1692 834
use sg13g2_dlhq_1  _1108_
timestamp 1678805552
transform -1 0 14880 0 -1 51408
box -50 -56 1692 834
use sg13g2_dlhq_1  _1109_
timestamp 1678805552
transform -1 0 9216 0 -1 71064
box -50 -56 1692 834
use sg13g2_dlhq_1  _1110_
timestamp 1678805552
transform -1 0 11136 0 1 69552
box -50 -56 1692 834
use sg13g2_dlhq_1  _1111_
timestamp 1678805552
transform 1 0 8544 0 1 71064
box -50 -56 1692 834
use sg13g2_dlhq_1  _1112_
timestamp 1678805552
transform 1 0 9408 0 -1 71064
box -50 -56 1692 834
use sg13g2_dlhq_1  _1113_
timestamp 1678805552
transform 1 0 9024 0 1 77112
box -50 -56 1692 834
use sg13g2_dlhq_1  _1114_
timestamp 1678805552
transform 1 0 8832 0 -1 78624
box -50 -56 1692 834
use sg13g2_dlhq_1  _1115_
timestamp 1678805552
transform -1 0 10944 0 1 72576
box -50 -56 1692 834
use sg13g2_dlhq_1  _1116_
timestamp 1678805552
transform -1 0 10368 0 -1 74088
box -50 -56 1692 834
use sg13g2_dlhq_1  _1117_
timestamp 1678805552
transform -1 0 10272 0 1 80136
box -50 -56 1692 834
use sg13g2_dlhq_1  _1118_
timestamp 1678805552
transform 1 0 7008 0 1 80136
box -50 -56 1692 834
use sg13g2_dlhq_1  _1119_
timestamp 1678805552
transform 1 0 10656 0 1 77112
box -50 -56 1692 834
use sg13g2_dlhq_1  _1120_
timestamp 1678805552
transform 1 0 10176 0 1 75600
box -50 -56 1692 834
use sg13g2_dlhq_1  _1121_
timestamp 1678805552
transform 1 0 13056 0 1 77112
box -50 -56 1692 834
use sg13g2_dlhq_1  _1122_
timestamp 1678805552
transform 1 0 11520 0 -1 77112
box -50 -56 1692 834
use sg13g2_dlhq_1  _1123_
timestamp 1678805552
transform 1 0 6240 0 1 60480
box -50 -56 1692 834
use sg13g2_dlhq_1  _1124_
timestamp 1678805552
transform -1 0 14112 0 1 60480
box -50 -56 1692 834
use sg13g2_dlhq_1  _1125_
timestamp 1678805552
transform 1 0 5952 0 -1 80136
box -50 -56 1692 834
use sg13g2_dlhq_1  _1126_
timestamp 1678805552
transform 1 0 4320 0 -1 80136
box -50 -56 1692 834
use sg13g2_dlhq_1  _1127_
timestamp 1678805552
transform 1 0 4416 0 1 80136
box -50 -56 1692 834
use sg13g2_dlhq_1  _1128_
timestamp 1678805552
transform 1 0 10368 0 -1 86184
box -50 -56 1692 834
use sg13g2_dlhq_1  _1129_
timestamp 1678805552
transform 1 0 10848 0 -1 84672
box -50 -56 1692 834
use sg13g2_dlhq_1  _1130_
timestamp 1678805552
transform 1 0 10560 0 1 84672
box -50 -56 1692 834
use sg13g2_dlhq_1  _1131_
timestamp 1678805552
transform 1 0 18528 0 1 80136
box -50 -56 1692 834
use sg13g2_dlhq_1  _1132_
timestamp 1678805552
transform 1 0 18048 0 1 78624
box -50 -56 1692 834
use sg13g2_dlhq_1  _1133_
timestamp 1678805552
transform 1 0 17376 0 -1 80136
box -50 -56 1692 834
use sg13g2_dlhq_1  _1134_
timestamp 1678805552
transform 1 0 6816 0 1 63504
box -50 -56 1692 834
use sg13g2_dlhq_1  _1135_
timestamp 1678805552
transform 1 0 6816 0 -1 65016
box -50 -56 1692 834
use sg13g2_dlhq_1  _1136_
timestamp 1678805552
transform 1 0 6048 0 1 65016
box -50 -56 1692 834
use sg13g2_dlhq_1  _1137_
timestamp 1678805552
transform 1 0 8448 0 1 75600
box -50 -56 1692 834
use sg13g2_dlhq_1  _1138_
timestamp 1678805552
transform 1 0 6816 0 1 75600
box -50 -56 1692 834
use sg13g2_dlhq_1  _1139_
timestamp 1678805552
transform 1 0 18432 0 1 75600
box -50 -56 1692 834
use sg13g2_dlhq_1  _1140_
timestamp 1678805552
transform 1 0 16800 0 -1 75600
box -50 -56 1692 834
use sg13g2_dlhq_1  _1141_
timestamp 1678805552
transform 1 0 13536 0 -1 72576
box -50 -56 1692 834
use sg13g2_dlhq_1  _1142_
timestamp 1678805552
transform 1 0 10944 0 1 72576
box -50 -56 1692 834
use sg13g2_dlhq_1  _1143_
timestamp 1678805552
transform 1 0 2016 0 -1 54432
box -50 -56 1692 834
use sg13g2_dlhq_1  _1144_
timestamp 1678805552
transform 1 0 1152 0 -1 52920
box -50 -56 1692 834
use sg13g2_dlhq_1  _1145_
timestamp 1678805552
transform 1 0 7296 0 -1 68040
box -50 -56 1692 834
use sg13g2_dlhq_1  _1146_
timestamp 1678805552
transform 1 0 5568 0 -1 68040
box -50 -56 1692 834
use sg13g2_dlhq_1  _1147_
timestamp 1678805552
transform 1 0 11904 0 -1 72576
box -50 -56 1692 834
use sg13g2_dlhq_1  _1148_
timestamp 1678805552
transform 1 0 10176 0 1 71064
box -50 -56 1692 834
use sg13g2_dlhq_1  _1149_
timestamp 1678805552
transform -1 0 19008 0 1 77112
box -50 -56 1692 834
use sg13g2_dlhq_1  _1150_
timestamp 1678805552
transform 1 0 14688 0 -1 80136
box -50 -56 1692 834
use sg13g2_dlhq_1  _1151_
timestamp 1678805552
transform 1 0 5664 0 1 77112
box -50 -56 1692 834
use sg13g2_dlhq_1  _1152_
timestamp 1678805552
transform 1 0 6240 0 -1 75600
box -50 -56 1692 834
use sg13g2_dlhq_1  _1153_
timestamp 1678805552
transform 1 0 7104 0 -1 86184
box -50 -56 1692 834
use sg13g2_dlhq_1  _1154_
timestamp 1678805552
transform -1 0 8352 0 1 87696
box -50 -56 1692 834
use sg13g2_dlhq_1  _1155_
timestamp 1678805552
transform -1 0 16704 0 -1 81648
box -50 -56 1692 834
use sg13g2_dlhq_1  _1156_
timestamp 1678805552
transform 1 0 12384 0 -1 78624
box -50 -56 1692 834
use sg13g2_dlhq_1  _1157_
timestamp 1678805552
transform 1 0 14016 0 1 75600
box -50 -56 1692 834
use sg13g2_dlhq_1  _1158_
timestamp 1678805552
transform 1 0 13056 0 -1 80136
box -50 -56 1692 834
use sg13g2_dlhq_1  _1159_
timestamp 1678805552
transform 1 0 6528 0 1 55944
box -50 -56 1692 834
use sg13g2_dlhq_1  _1160_
timestamp 1678805552
transform 1 0 7392 0 1 57456
box -50 -56 1692 834
use sg13g2_dlhq_1  _1161_
timestamp 1678805552
transform 1 0 9120 0 -1 45360
box -50 -56 1692 834
use sg13g2_dlhq_1  _1162_
timestamp 1678805552
transform 1 0 8256 0 1 45360
box -50 -56 1692 834
use sg13g2_dlhq_1  _1163_
timestamp 1678805552
transform 1 0 8160 0 1 34776
box -50 -56 1692 834
use sg13g2_dlhq_1  _1164_
timestamp 1678805552
transform 1 0 6816 0 -1 36288
box -50 -56 1692 834
use sg13g2_dlhq_1  _1165_
timestamp 1678805552
transform 1 0 12000 0 1 22680
box -50 -56 1692 834
use sg13g2_dlhq_1  _1166_
timestamp 1678805552
transform 1 0 11616 0 -1 22680
box -50 -56 1692 834
use sg13g2_dlhq_1  _1167_
timestamp 1678805552
transform 1 0 5952 0 1 33264
box -50 -56 1692 834
use sg13g2_dlhq_1  _1168_
timestamp 1678805552
transform 1 0 5952 0 -1 34776
box -50 -56 1692 834
use sg13g2_dlhq_1  _1169_
timestamp 1678805552
transform 1 0 9888 0 1 48384
box -50 -56 1692 834
use sg13g2_dlhq_1  _1170_
timestamp 1678805552
transform 1 0 9024 0 1 40824
box -50 -56 1692 834
use sg13g2_dlhq_1  _1171_
timestamp 1678805552
transform 1 0 15936 0 1 46872
box -50 -56 1692 834
use sg13g2_dlhq_1  _1172_
timestamp 1678805552
transform 1 0 14304 0 1 46872
box -50 -56 1692 834
use sg13g2_dlhq_1  _1173_
timestamp 1678805552
transform 1 0 17952 0 1 46872
box -50 -56 1692 834
use sg13g2_dlhq_1  _1174_
timestamp 1678805552
transform 1 0 17568 0 -1 48384
box -50 -56 1692 834
use sg13g2_dlhq_1  _1175_
timestamp 1678805552
transform 1 0 1536 0 1 46872
box -50 -56 1692 834
use sg13g2_dlhq_1  _1176_
timestamp 1678805552
transform 1 0 1248 0 -1 46872
box -50 -56 1692 834
use sg13g2_dlhq_1  _1177_
timestamp 1678805552
transform 1 0 3456 0 -1 42336
box -50 -56 1692 834
use sg13g2_dlhq_1  _1178_
timestamp 1678805552
transform 1 0 6432 0 1 36288
box -50 -56 1692 834
use sg13g2_dlhq_1  _1179_
timestamp 1678805552
transform 1 0 9216 0 -1 42336
box -50 -56 1692 834
use sg13g2_dlhq_1  _1180_
timestamp 1678805552
transform 1 0 9888 0 1 34776
box -50 -56 1692 834
use sg13g2_dlhq_1  _1181_
timestamp 1678805552
transform 1 0 15936 0 -1 49896
box -50 -56 1692 834
use sg13g2_dlhq_1  _1182_
timestamp 1678805552
transform 1 0 14304 0 -1 49896
box -50 -56 1692 834
use sg13g2_dlhq_1  _1183_
timestamp 1678805552
transform 1 0 4416 0 -1 36288
box -50 -56 1692 834
use sg13g2_dlhq_1  _1184_
timestamp 1678805552
transform 1 0 3840 0 1 34776
box -50 -56 1692 834
use sg13g2_dlhq_1  _1185_
timestamp 1678805552
transform 1 0 8448 0 -1 36288
box -50 -56 1692 834
use sg13g2_dlhq_1  _1186_
timestamp 1678805552
transform 1 0 7584 0 1 33264
box -50 -56 1692 834
use sg13g2_dlhq_1  _1187_
timestamp 1678805552
transform 1 0 11136 0 -1 13608
box -50 -56 1692 834
use sg13g2_dlhq_1  _1188_
timestamp 1678805552
transform 1 0 9504 0 -1 13608
box -50 -56 1692 834
use sg13g2_dlhq_1  _1189_
timestamp 1678805552
transform -1 0 16800 0 -1 16632
box -50 -56 1692 834
use sg13g2_dlhq_1  _1190_
timestamp 1678805552
transform 1 0 11424 0 1 16632
box -50 -56 1692 834
use sg13g2_dlhq_1  _1191_
timestamp 1678805552
transform 1 0 9312 0 -1 22680
box -50 -56 1692 834
use sg13g2_dlhq_1  _1192_
timestamp 1678805552
transform -1 0 10560 0 1 21168
box -50 -56 1692 834
use sg13g2_dlhq_1  _1193_
timestamp 1678805552
transform 1 0 8640 0 -1 33264
box -50 -56 1692 834
use sg13g2_dlhq_1  _1194_
timestamp 1678805552
transform 1 0 7584 0 -1 34776
box -50 -56 1692 834
use sg13g2_dlhq_1  _1195_
timestamp 1678805552
transform 1 0 12288 0 1 7560
box -50 -56 1692 834
use sg13g2_dlhq_1  _1196_
timestamp 1678805552
transform 1 0 10272 0 1 7560
box -50 -56 1692 834
use sg13g2_dlhq_1  _1197_
timestamp 1678805552
transform 1 0 10944 0 1 15120
box -50 -56 1692 834
use sg13g2_dlhq_1  _1198_
timestamp 1678805552
transform 1 0 10848 0 1 13608
box -50 -56 1692 834
use sg13g2_dlhq_1  _1199_
timestamp 1678805552
transform 1 0 9120 0 -1 16632
box -50 -56 1692 834
use sg13g2_dlhq_1  _1200_
timestamp 1678805552
transform 1 0 6624 0 1 16632
box -50 -56 1692 834
use sg13g2_dlhq_1  _1201_
timestamp 1678805552
transform 1 0 10080 0 -1 31752
box -50 -56 1692 834
use sg13g2_dlhq_1  _1202_
timestamp 1678805552
transform 1 0 8448 0 -1 31752
box -50 -56 1692 834
use sg13g2_dlhq_1  _1203_
timestamp 1678805552
transform -1 0 15552 0 1 7560
box -50 -56 1692 834
use sg13g2_dlhq_1  _1204_
timestamp 1678805552
transform 1 0 10560 0 -1 7560
box -50 -56 1692 834
use sg13g2_dlhq_1  _1205_
timestamp 1678805552
transform 1 0 12864 0 -1 13608
box -50 -56 1692 834
use sg13g2_dlhq_1  _1206_
timestamp 1678805552
transform 1 0 10944 0 -1 15120
box -50 -56 1692 834
use sg13g2_dlhq_1  _1207_
timestamp 1678805552
transform 1 0 7200 0 1 19656
box -50 -56 1692 834
use sg13g2_dlhq_1  _1208_
timestamp 1678805552
transform 1 0 5568 0 -1 21168
box -50 -56 1692 834
use sg13g2_dlhq_1  _1209_
timestamp 1678805552
transform -1 0 12096 0 -1 28728
box -50 -56 1692 834
use sg13g2_dlhq_1  _1210_
timestamp 1678805552
transform -1 0 12768 0 1 27216
box -50 -56 1692 834
use sg13g2_dlhq_1  _1211_
timestamp 1678805552
transform 1 0 12768 0 -1 7560
box -50 -56 1692 834
use sg13g2_dlhq_1  _1212_
timestamp 1678805552
transform 1 0 10368 0 -1 9072
box -50 -56 1692 834
use sg13g2_dlhq_1  _1213_
timestamp 1678805552
transform 1 0 13056 0 1 15120
box -50 -56 1692 834
use sg13g2_dlhq_1  _1214_
timestamp 1678805552
transform 1 0 11136 0 -1 16632
box -50 -56 1692 834
use sg13g2_dlhq_1  _1215_
timestamp 1678805552
transform 1 0 6528 0 -1 22680
box -50 -56 1692 834
use sg13g2_dlhq_1  _1216_
timestamp 1678805552
transform 1 0 4608 0 1 22680
box -50 -56 1692 834
use sg13g2_dlhq_1  _1217_
timestamp 1678805552
transform 1 0 3936 0 -1 37800
box -50 -56 1692 834
use sg13g2_dlhq_1  _1218_
timestamp 1678805552
transform 1 0 4320 0 1 33264
box -50 -56 1692 834
use sg13g2_dlhq_1  _1219_
timestamp 1678805552
transform 1 0 4800 0 1 28728
box -50 -56 1692 834
use sg13g2_dlhq_1  _1220_
timestamp 1678805552
transform 1 0 5472 0 1 34776
box -50 -56 1692 834
use sg13g2_dlhq_1  _1221_
timestamp 1678805552
transform -1 0 6912 0 -1 46872
box -50 -56 1692 834
use sg13g2_dlhq_1  _1222_
timestamp 1678805552
transform 1 0 2688 0 -1 45360
box -50 -56 1692 834
use sg13g2_dlhq_1  _1223_
timestamp 1678805552
transform 1 0 2400 0 -1 43848
box -50 -56 1692 834
use sg13g2_dlhq_1  _1224_
timestamp 1678805552
transform 1 0 2496 0 1 42336
box -50 -56 1692 834
use sg13g2_dlhq_1  _1225_
timestamp 1678805552
transform 1 0 8832 0 -1 43848
box -50 -56 1692 834
use sg13g2_dlhq_1  _1226_
timestamp 1678805552
transform 1 0 7488 0 1 43848
box -50 -56 1692 834
use sg13g2_dlhq_1  _1227_
timestamp 1678805552
transform 1 0 7584 0 -1 42336
box -50 -56 1692 834
use sg13g2_dlhq_1  _1228_
timestamp 1678805552
transform 1 0 7392 0 1 40824
box -50 -56 1692 834
use sg13g2_dlhq_1  _1229_
timestamp 1678805552
transform 1 0 13536 0 1 43848
box -50 -56 1692 834
use sg13g2_dlhq_1  _1230_
timestamp 1678805552
transform 1 0 11904 0 1 43848
box -50 -56 1692 834
use sg13g2_dlhq_1  _1231_
timestamp 1678805552
transform 1 0 12960 0 -1 36288
box -50 -56 1692 834
use sg13g2_dlhq_1  _1232_
timestamp 1678805552
transform 1 0 11520 0 1 34776
box -50 -56 1692 834
use sg13g2_dlhq_1  _1233_
timestamp 1678805552
transform 1 0 18432 0 -1 21168
box -50 -56 1692 834
use sg13g2_dlhq_1  _1234_
timestamp 1678805552
transform 1 0 16512 0 1 19656
box -50 -56 1692 834
use sg13g2_dlhq_1  _1235_
timestamp 1678805552
transform -1 0 13632 0 1 25704
box -50 -56 1692 834
use sg13g2_dlhq_1  _1236_
timestamp 1678805552
transform -1 0 12960 0 -1 27216
box -50 -56 1692 834
use sg13g2_dlhq_1  _1237_
timestamp 1678805552
transform 1 0 18144 0 -1 42336
box -50 -56 1692 834
use sg13g2_dlhq_1  _1238_
timestamp 1678805552
transform 1 0 16224 0 -1 43848
box -50 -56 1692 834
use sg13g2_dlhq_1  _1239_
timestamp 1678805552
transform 1 0 18624 0 1 36288
box -50 -56 1692 834
use sg13g2_dlhq_1  _1240_
timestamp 1678805552
transform 1 0 16896 0 -1 39312
box -50 -56 1692 834
use sg13g2_dlhq_1  _1241_
timestamp 1678805552
transform 1 0 16608 0 -1 22680
box -50 -56 1692 834
use sg13g2_dlhq_1  _1242_
timestamp 1678805552
transform 1 0 14976 0 -1 22680
box -50 -56 1692 834
use sg13g2_dlhq_1  _1243_
timestamp 1678805552
transform -1 0 9312 0 1 27216
box -50 -56 1692 834
use sg13g2_dlhq_1  _1244_
timestamp 1678805552
transform 1 0 5280 0 -1 28728
box -50 -56 1692 834
use sg13g2_dlhq_1  _1245_
timestamp 1678805552
transform -1 0 16896 0 -1 46872
box -50 -56 1692 834
use sg13g2_dlhq_1  _1246_
timestamp 1678805552
transform 1 0 12672 0 1 46872
box -50 -56 1692 834
use sg13g2_dlhq_1  _1247_
timestamp 1678805552
transform 1 0 18720 0 -1 31752
box -50 -56 1692 834
use sg13g2_dlhq_1  _1248_
timestamp 1678805552
transform 1 0 16992 0 -1 31752
box -50 -56 1692 834
use sg13g2_dlhq_1  _1249_
timestamp 1678805552
transform 1 0 18432 0 1 18144
box -50 -56 1692 834
use sg13g2_dlhq_1  _1250_
timestamp 1678805552
transform 1 0 16416 0 -1 19656
box -50 -56 1692 834
use sg13g2_dlhq_1  _1251_
timestamp 1678805552
transform -1 0 12960 0 -1 25704
box -50 -56 1692 834
use sg13g2_dlhq_1  _1252_
timestamp 1678805552
transform 1 0 4320 0 -1 27216
box -50 -56 1692 834
use sg13g2_dlhq_1  _1253_
timestamp 1678805552
transform 1 0 17760 0 -1 46872
box -50 -56 1692 834
use sg13g2_dlhq_1  _1254_
timestamp 1678805552
transform 1 0 15936 0 -1 45360
box -50 -56 1692 834
use sg13g2_dlhq_1  _1255_
timestamp 1678805552
transform 1 0 18720 0 1 34776
box -50 -56 1692 834
use sg13g2_dlhq_1  _1256_
timestamp 1678805552
transform 1 0 17568 0 -1 34776
box -50 -56 1692 834
use sg13g2_dlhq_1  _1257_
timestamp 1678805552
transform -1 0 18720 0 1 25704
box -50 -56 1692 834
use sg13g2_dlhq_1  _1258_
timestamp 1678805552
transform 1 0 14400 0 -1 25704
box -50 -56 1692 834
use sg13g2_dlhq_1  _1259_
timestamp 1678805552
transform 1 0 6048 0 1 27216
box -50 -56 1692 834
use sg13g2_dlhq_1  _1260_
timestamp 1678805552
transform 1 0 5952 0 -1 27216
box -50 -56 1692 834
use sg13g2_dlhq_1  _1261_
timestamp 1678805552
transform 1 0 12864 0 -1 48384
box -50 -56 1692 834
use sg13g2_dlhq_1  _1262_
timestamp 1678805552
transform 1 0 11904 0 1 45360
box -50 -56 1692 834
use sg13g2_dlhq_1  _1263_
timestamp 1678805552
transform 1 0 14112 0 1 33264
box -50 -56 1692 834
use sg13g2_dlhq_1  _1264_
timestamp 1678805552
transform 1 0 12384 0 -1 34776
box -50 -56 1692 834
use sg13g2_dlhq_1  _1265_
timestamp 1678805552
transform 1 0 18720 0 1 13608
box -50 -56 1692 834
use sg13g2_dlhq_1  _1266_
timestamp 1678805552
transform 1 0 16992 0 1 13608
box -50 -56 1692 834
use sg13g2_dlhq_1  _1267_
timestamp 1678805552
transform 1 0 9792 0 1 24192
box -50 -56 1692 834
use sg13g2_dlhq_1  _1268_
timestamp 1678805552
transform 1 0 7776 0 -1 24192
box -50 -56 1692 834
use sg13g2_dlhq_1  _1269_
timestamp 1678805552
transform 1 0 16512 0 -1 42336
box -50 -56 1692 834
use sg13g2_dlhq_1  _1270_
timestamp 1678805552
transform 1 0 16224 0 1 42336
box -50 -56 1692 834
use sg13g2_dlhq_1  _1271_
timestamp 1678805552
transform 1 0 18624 0 -1 39312
box -50 -56 1692 834
use sg13g2_dlhq_1  _1272_
timestamp 1678805552
transform 1 0 16704 0 1 37800
box -50 -56 1692 834
use sg13g2_dlhq_1  _1273_
timestamp 1678805552
transform 1 0 15168 0 -1 27216
box -50 -56 1692 834
use sg13g2_dlhq_1  _1274_
timestamp 1678805552
transform 1 0 13536 0 -1 27216
box -50 -56 1692 834
use sg13g2_dlhq_1  _1275_
timestamp 1678805552
transform -1 0 10464 0 1 30240
box -50 -56 1692 834
use sg13g2_dlhq_1  _1276_
timestamp 1678805552
transform 1 0 5184 0 1 30240
box -50 -56 1692 834
use sg13g2_dlhq_1  _1277_
timestamp 1678805552
transform 1 0 14400 0 -1 39312
box -50 -56 1692 834
use sg13g2_dlhq_1  _1278_
timestamp 1678805552
transform 1 0 13152 0 1 37800
box -50 -56 1692 834
use sg13g2_dlhq_1  _1279_
timestamp 1678805552
transform 1 0 18624 0 1 33264
box -50 -56 1692 834
use sg13g2_dlhq_1  _1280_
timestamp 1678805552
transform 1 0 16992 0 1 33264
box -50 -56 1692 834
use sg13g2_dlhq_1  _1281_
timestamp 1678805552
transform 1 0 18624 0 -1 15120
box -50 -56 1692 834
use sg13g2_dlhq_1  _1282_
timestamp 1678805552
transform 1 0 16608 0 1 15120
box -50 -56 1692 834
use sg13g2_dlhq_1  _1283_
timestamp 1678805552
transform 1 0 7584 0 -1 25704
box -50 -56 1692 834
use sg13g2_dlhq_1  _1284_
timestamp 1678805552
transform 1 0 5760 0 1 25704
box -50 -56 1692 834
use sg13g2_dlhq_1  _1285_
timestamp 1678805552
transform 1 0 18624 0 1 43848
box -50 -56 1692 834
use sg13g2_dlhq_1  _1286_
timestamp 1678805552
transform 1 0 16128 0 1 43848
box -50 -56 1692 834
use sg13g2_dlhq_1  _1287_
timestamp 1678805552
transform 1 0 18816 0 1 39312
box -50 -56 1692 834
use sg13g2_dlhq_1  _1288_
timestamp 1678805552
transform 1 0 16320 0 1 40824
box -50 -56 1692 834
use sg13g2_dlhq_1  _1289_
timestamp 1678805552
transform 1 0 18048 0 -1 25704
box -50 -56 1692 834
use sg13g2_dlhq_1  _1290_
timestamp 1678805552
transform 1 0 15264 0 1 24192
box -50 -56 1692 834
use sg13g2_dlhq_1  _1291_
timestamp 1678805552
transform 1 0 6720 0 -1 31752
box -50 -56 1692 834
use sg13g2_dlhq_1  _1292_
timestamp 1678805552
transform 1 0 4896 0 -1 30240
box -50 -56 1692 834
use sg13g2_dlhq_1  _1293_
timestamp 1678805552
transform -1 0 4608 0 -1 31752
box -50 -56 1692 834
use sg13g2_dlhq_1  _1294_
timestamp 1678805552
transform 1 0 1152 0 1 30240
box -50 -56 1692 834
use sg13g2_dlhq_1  _1295_
timestamp 1678805552
transform 1 0 4800 0 1 36288
box -50 -56 1692 834
use sg13g2_dlhq_1  _1296_
timestamp 1678805552
transform 1 0 5568 0 -1 37800
box -50 -56 1692 834
use sg13g2_dlhq_1  _1297_
timestamp 1678805552
transform 1 0 18336 0 1 27216
box -50 -56 1692 834
use sg13g2_dlhq_1  _1298_
timestamp 1678805552
transform 1 0 17568 0 -1 28728
box -50 -56 1692 834
use sg13g2_dlhq_1  _1299_
timestamp 1678805552
transform 1 0 14976 0 1 27216
box -50 -56 1692 834
use sg13g2_dlhq_1  _1300_
timestamp 1678805552
transform 1 0 14304 0 -1 28728
box -50 -56 1692 834
use sg13g2_dlhq_1  _1301_
timestamp 1678805552
transform 1 0 5376 0 1 21168
box -50 -56 1692 834
use sg13g2_dlhq_1  _1302_
timestamp 1678805552
transform 1 0 5088 0 1 19656
box -50 -56 1692 834
use sg13g2_dlhq_1  _1303_
timestamp 1678805552
transform 1 0 1344 0 1 25704
box -50 -56 1692 834
use sg13g2_dlhq_1  _1304_
timestamp 1678805552
transform 1 0 1824 0 -1 25704
box -50 -56 1692 834
use sg13g2_dlhq_1  _1305_
timestamp 1678805552
transform 1 0 14304 0 1 18144
box -50 -56 1692 834
use sg13g2_dlhq_1  _1306_
timestamp 1678805552
transform 1 0 15456 0 1 16632
box -50 -56 1692 834
use sg13g2_dlhq_1  _1307_
timestamp 1678805552
transform 1 0 8832 0 1 19656
box -50 -56 1692 834
use sg13g2_dlhq_1  _1308_
timestamp 1678805552
transform 1 0 10752 0 -1 19656
box -50 -56 1692 834
use sg13g2_dlhq_1  _1309_
timestamp 1678805552
transform 1 0 4032 0 -1 13608
box -50 -56 1692 834
use sg13g2_dlhq_1  _1310_
timestamp 1678805552
transform 1 0 4992 0 -1 12096
box -50 -56 1692 834
use sg13g2_dlhq_1  _1311_
timestamp 1678805552
transform 1 0 5664 0 1 18144
box -50 -56 1692 834
use sg13g2_dlhq_1  _1312_
timestamp 1678805552
transform 1 0 3456 0 1 19656
box -50 -56 1692 834
use sg13g2_dlhq_1  _1313_
timestamp 1678805552
transform 1 0 17664 0 1 16632
box -50 -56 1692 834
use sg13g2_dlhq_1  _1314_
timestamp 1678805552
transform 1 0 15936 0 1 18144
box -50 -56 1692 834
use sg13g2_dlhq_1  _1315_
timestamp 1678805552
transform 1 0 6432 0 1 6048
box -50 -56 1692 834
use sg13g2_dlhq_1  _1316_
timestamp 1678805552
transform 1 0 5184 0 -1 6048
box -50 -56 1692 834
use sg13g2_dlhq_1  _1317_
timestamp 1678805552
transform 1 0 2976 0 1 7560
box -50 -56 1692 834
use sg13g2_dlhq_1  _1318_
timestamp 1678805552
transform 1 0 4704 0 -1 10584
box -50 -56 1692 834
use sg13g2_dlhq_1  _1319_
timestamp 1678805552
transform 1 0 9504 0 1 27216
box -50 -56 1692 834
use sg13g2_dlhq_1  _1320_
timestamp 1678805552
transform -1 0 11904 0 -1 33264
box -50 -56 1692 834
use sg13g2_dlhq_1  _1321_
timestamp 1678805552
transform 1 0 13536 0 1 10584
box -50 -56 1692 834
use sg13g2_dlhq_1  _1322_
timestamp 1678805552
transform 1 0 11616 0 -1 12096
box -50 -56 1692 834
use sg13g2_dlhq_1  _1323_
timestamp 1678805552
transform 1 0 15360 0 1 12096
box -50 -56 1692 834
use sg13g2_dlhq_1  _1324_
timestamp 1678805552
transform 1 0 13728 0 1 12096
box -50 -56 1692 834
use sg13g2_dlhq_1  _1325_
timestamp 1678805552
transform 1 0 9216 0 1 15120
box -50 -56 1692 834
use sg13g2_dlhq_1  _1326_
timestamp 1678805552
transform 1 0 7392 0 -1 16632
box -50 -56 1692 834
use sg13g2_dlhq_1  _1327_
timestamp 1678805552
transform 1 0 1248 0 1 24192
box -50 -56 1692 834
use sg13g2_dlhq_1  _1328_
timestamp 1678805552
transform 1 0 1248 0 -1 24192
box -50 -56 1692 834
use sg13g2_dlhq_1  _1329_
timestamp 1678805552
transform 1 0 18432 0 -1 12096
box -50 -56 1692 834
use sg13g2_dlhq_1  _1330_
timestamp 1678805552
transform 1 0 16800 0 -1 12096
box -50 -56 1692 834
use sg13g2_dlhq_1  _1331_
timestamp 1678805552
transform 1 0 8544 0 -1 9072
box -50 -56 1692 834
use sg13g2_dlhq_1  _1332_
timestamp 1678805552
transform 1 0 7488 0 1 9072
box -50 -56 1692 834
use sg13g2_dlhq_1  _1333_
timestamp 1678805552
transform 1 0 4608 0 -1 15120
box -50 -56 1692 834
use sg13g2_dlhq_1  _1334_
timestamp 1678805552
transform 1 0 2976 0 -1 15120
box -50 -56 1692 834
use sg13g2_dlhq_1  _1335_
timestamp 1678805552
transform 1 0 1248 0 -1 19656
box -50 -56 1692 834
use sg13g2_dlhq_1  _1336_
timestamp 1678805552
transform 1 0 1152 0 1 19656
box -50 -56 1692 834
use sg13g2_dlhq_1  _1337_
timestamp 1678805552
transform 1 0 15840 0 -1 13608
box -50 -56 1692 834
use sg13g2_dlhq_1  _1338_
timestamp 1678805552
transform 1 0 14976 0 1 15120
box -50 -56 1692 834
use sg13g2_dlhq_1  _1339_
timestamp 1678805552
transform 1 0 13152 0 1 6048
box -50 -56 1692 834
use sg13g2_dlhq_1  _1340_
timestamp 1678805552
transform 1 0 11040 0 1 6048
box -50 -56 1692 834
use sg13g2_dlhq_1  _1341_
timestamp 1678805552
transform 1 0 4704 0 1 7560
box -50 -56 1692 834
use sg13g2_dlhq_1  _1342_
timestamp 1678805552
transform -1 0 5472 0 1 6048
box -50 -56 1692 834
use sg13g2_dlhq_1  _1343_
timestamp 1678805552
transform -1 0 6240 0 1 15120
box -50 -56 1692 834
use sg13g2_dlhq_1  _1344_
timestamp 1678805552
transform 1 0 1536 0 -1 13608
box -50 -56 1692 834
use sg13g2_dlhq_1  _1345_
timestamp 1678805552
transform 1 0 15360 0 1 9072
box -50 -56 1692 834
use sg13g2_dlhq_1  _1346_
timestamp 1678805552
transform 1 0 14304 0 -1 10584
box -50 -56 1692 834
use sg13g2_dlhq_1  _1347_
timestamp 1678805552
transform 1 0 10848 0 -1 4536
box -50 -56 1692 834
use sg13g2_dlhq_1  _1348_
timestamp 1678805552
transform 1 0 9024 0 1 4536
box -50 -56 1692 834
use sg13g2_dlhq_1  _1349_
timestamp 1678805552
transform 1 0 2304 0 -1 7560
box -50 -56 1692 834
use sg13g2_dlhq_1  _1350_
timestamp 1678805552
transform 1 0 1344 0 1 7560
box -50 -56 1692 834
use sg13g2_dlhq_1  _1351_
timestamp 1678805552
transform 1 0 3840 0 -1 21168
box -50 -56 1692 834
use sg13g2_dlhq_1  _1352_
timestamp 1678805552
transform 1 0 1824 0 -1 22680
box -50 -56 1692 834
use sg13g2_dlhq_1  _1353_
timestamp 1678805552
transform 1 0 17856 0 1 10584
box -50 -56 1692 834
use sg13g2_dlhq_1  _1354_
timestamp 1678805552
transform 1 0 16128 0 -1 10584
box -50 -56 1692 834
use sg13g2_dlhq_1  _1355_
timestamp 1678805552
transform -1 0 19296 0 -1 7560
box -50 -56 1692 834
use sg13g2_dlhq_1  _1356_
timestamp 1678805552
transform -1 0 17664 0 -1 7560
box -50 -56 1692 834
use sg13g2_dlhq_1  _1357_
timestamp 1678805552
transform 1 0 6912 0 -1 12096
box -50 -56 1692 834
use sg13g2_dlhq_1  _1358_
timestamp 1678805552
transform 1 0 5760 0 -1 13608
box -50 -56 1692 834
use sg13g2_dlhq_1  _1359_
timestamp 1678805552
transform 1 0 1632 0 -1 16632
box -50 -56 1692 834
use sg13g2_dlhq_1  _1360_
timestamp 1678805552
transform 1 0 1248 0 1 15120
box -50 -56 1692 834
use sg13g2_dlhq_1  _1361_
timestamp 1678805552
transform 1 0 18432 0 1 7560
box -50 -56 1692 834
use sg13g2_dlhq_1  _1362_
timestamp 1678805552
transform 1 0 17664 0 -1 9072
box -50 -56 1692 834
use sg13g2_dlhq_1  _1363_
timestamp 1678805552
transform 1 0 8544 0 1 7560
box -50 -56 1692 834
use sg13g2_dlhq_1  _1364_
timestamp 1678805552
transform 1 0 6912 0 -1 7560
box -50 -56 1692 834
use sg13g2_dlhq_1  _1365_
timestamp 1678805552
transform 1 0 2112 0 -1 12096
box -50 -56 1692 834
use sg13g2_dlhq_1  _1366_
timestamp 1678805552
transform 1 0 1152 0 1 10584
box -50 -56 1692 834
use sg13g2_dlhq_1  _1367_
timestamp 1678805552
transform 1 0 1536 0 -1 18144
box -50 -56 1692 834
use sg13g2_dlhq_1  _1368_
timestamp 1678805552
transform 1 0 1152 0 1 16632
box -50 -56 1692 834
use sg13g2_dlhq_1  _1369_
timestamp 1678805552
transform 1 0 7584 0 1 15120
box -50 -56 1692 834
use sg13g2_dlhq_1  _1370_
timestamp 1678805552
transform 1 0 6240 0 -1 15120
box -50 -56 1692 834
use sg13g2_dlhq_1  _1371_
timestamp 1678805552
transform 1 0 14784 0 -1 6048
box -50 -56 1692 834
use sg13g2_dlhq_1  _1372_
timestamp 1678805552
transform 1 0 8448 0 -1 6048
box -50 -56 1692 834
use sg13g2_dlhq_1  _1373_
timestamp 1678805552
transform 1 0 6432 0 1 7560
box -50 -56 1692 834
use sg13g2_dlhq_1  _1374_
timestamp 1678805552
transform 1 0 5184 0 -1 7560
box -50 -56 1692 834
use sg13g2_dlhq_1  _1375_
timestamp 1678805552
transform 1 0 2976 0 1 15120
box -50 -56 1692 834
use sg13g2_dlhq_1  _1376_
timestamp 1678805552
transform 1 0 1344 0 -1 15120
box -50 -56 1692 834
use sg13g2_dlhq_1  _1377_
timestamp 1678805552
transform 1 0 18240 0 1 6048
box -50 -56 1692 834
use sg13g2_dlhq_1  _1378_
timestamp 1678805552
transform 1 0 16224 0 1 7560
box -50 -56 1692 834
use sg13g2_dlhq_1  _1379_
timestamp 1678805552
transform 1 0 6816 0 -1 6048
box -50 -56 1692 834
use sg13g2_dlhq_1  _1380_
timestamp 1678805552
transform 1 0 6528 0 1 4536
box -50 -56 1692 834
use sg13g2_dlhq_1  _1381_
timestamp 1678805552
transform 1 0 1824 0 1 9072
box -50 -56 1692 834
use sg13g2_dlhq_1  _1382_
timestamp 1678805552
transform 1 0 1152 0 -1 9072
box -50 -56 1692 834
use sg13g2_dlhq_1  _1383_
timestamp 1678805552
transform 1 0 1824 0 1 22680
box -50 -56 1692 834
use sg13g2_dlhq_1  _1384_
timestamp 1678805552
transform 1 0 1152 0 -1 21168
box -50 -56 1692 834
use sg13g2_dlhq_1  _1385_
timestamp 1678805552
transform 1 0 8544 0 1 12096
box -50 -56 1692 834
use sg13g2_dlhq_1  _1386_
timestamp 1678805552
transform -1 0 9600 0 1 10584
box -50 -56 1692 834
use sg13g2_dlhq_1  _1387_
timestamp 1678805552
transform -1 0 18048 0 -1 6048
box -50 -56 1692 834
use sg13g2_dlhq_1  _1388_
timestamp 1678805552
transform -1 0 16032 0 -1 7560
box -50 -56 1692 834
use sg13g2_dlhq_1  _1389_
timestamp 1678805552
transform 1 0 6432 0 -1 10584
box -50 -56 1692 834
use sg13g2_dlhq_1  _1390_
timestamp 1678805552
transform 1 0 4320 0 1 10584
box -50 -56 1692 834
use sg13g2_dlhq_1  _1391_
timestamp 1678805552
transform 1 0 7296 0 1 21168
box -50 -56 1692 834
use sg13g2_dlhq_1  _1392_
timestamp 1678805552
transform -1 0 12192 0 1 21168
box -50 -56 1692 834
use sg13g2_dlhq_1  _1393_
timestamp 1678805552
transform 1 0 9696 0 1 10584
box -50 -56 1692 834
use sg13g2_dlhq_1  _1394_
timestamp 1678805552
transform 1 0 10656 0 -1 10584
box -50 -56 1692 834
use sg13g2_dlhq_1  _1395_
timestamp 1678805552
transform 1 0 10656 0 1 18144
box -50 -56 1692 834
use sg13g2_dlhq_1  _1396_
timestamp 1678805552
transform 1 0 11808 0 -1 18144
box -50 -56 1692 834
use sg13g2_dlhq_1  _1397_
timestamp 1678805552
transform 1 0 4992 0 1 16632
box -50 -56 1692 834
use sg13g2_dlhq_1  _1398_
timestamp 1678805552
transform 1 0 6624 0 -1 18144
box -50 -56 1692 834
use sg13g2_dlhq_1  _1399_
timestamp 1678805552
transform 1 0 11040 0 -1 39312
box -50 -56 1692 834
use sg13g2_dlhq_1  _1400_
timestamp 1678805552
transform 1 0 10560 0 1 37800
box -50 -56 1692 834
use sg13g2_dlhq_1  _1401_
timestamp 1678805552
transform 1 0 10656 0 -1 37800
box -50 -56 1692 834
use sg13g2_dlhq_1  _1402_
timestamp 1678805552
transform 1 0 12480 0 -1 28728
box -50 -56 1692 834
use sg13g2_dlhq_1  _1403_
timestamp 1678805552
transform 1 0 11232 0 1 30240
box -50 -56 1692 834
use sg13g2_dlhq_1  _1404_
timestamp 1678805552
transform 1 0 11904 0 -1 31752
box -50 -56 1692 834
use sg13g2_dlhq_1  _1405_
timestamp 1678805552
transform 1 0 16608 0 1 21168
box -50 -56 1692 834
use sg13g2_dlhq_1  _1406_
timestamp 1678805552
transform 1 0 16608 0 -1 21168
box -50 -56 1692 834
use sg13g2_dlhq_1  _1407_
timestamp 1678805552
transform 1 0 18528 0 1 22680
box -50 -56 1692 834
use sg13g2_dlhq_1  _1408_
timestamp 1678805552
transform 1 0 1440 0 -1 27216
box -50 -56 1692 834
use sg13g2_dlhq_1  _1409_
timestamp 1678805552
transform 1 0 1536 0 1 27216
box -50 -56 1692 834
use sg13g2_dlhq_1  _1410_
timestamp 1678805552
transform 1 0 1440 0 -1 28728
box -50 -56 1692 834
use sg13g2_dlhq_1  _1411_
timestamp 1678805552
transform 1 0 5280 0 -1 25704
box -50 -56 1692 834
use sg13g2_dlhq_1  _1412_
timestamp 1678805552
transform 1 0 5952 0 -1 24192
box -50 -56 1692 834
use sg13g2_dlhq_1  _1413_
timestamp 1678805552
transform 1 0 18336 0 1 28728
box -50 -56 1692 834
use sg13g2_dlhq_1  _1414_
timestamp 1678805552
transform 1 0 15936 0 -1 28728
box -50 -56 1692 834
use sg13g2_dlhq_1  _1415_
timestamp 1678805552
transform 1 0 18720 0 1 25704
box -50 -56 1692 834
use sg13g2_dlhq_1  _1416_
timestamp 1678805552
transform 1 0 16704 0 1 27216
box -50 -56 1692 834
use sg13g2_dlhq_1  _1417_
timestamp 1678805552
transform 1 0 1344 0 -1 31752
box -50 -56 1692 834
use sg13g2_dlhq_1  _1418_
timestamp 1678805552
transform 1 0 3168 0 -1 33264
box -50 -56 1692 834
use sg13g2_dlhq_1  _1419_
timestamp 1678805552
transform 1 0 1152 0 1 33264
box -50 -56 1692 834
use sg13g2_dlhq_1  _1420_
timestamp 1678805552
transform 1 0 2016 0 1 34776
box -50 -56 1692 834
use sg13g2_dlhq_1  _1421_
timestamp 1678805552
transform 1 0 9600 0 1 42336
box -50 -56 1692 834
use sg13g2_dlhq_1  _1422_
timestamp 1678805552
transform 1 0 11232 0 1 42336
box -50 -56 1692 834
use sg13g2_dlhq_1  _1423_
timestamp 1678805552
transform 1 0 12480 0 1 33264
box -50 -56 1692 834
use sg13g2_dlhq_1  _1424_
timestamp 1678805552
transform 1 0 11904 0 -1 33264
box -50 -56 1692 834
use sg13g2_dlhq_1  _1425_
timestamp 1678805552
transform 1 0 2400 0 -1 39312
box -50 -56 1692 834
use sg13g2_dlhq_1  _1426_
timestamp 1678805552
transform 1 0 1152 0 -1 37800
box -50 -56 1692 834
use sg13g2_dlhq_1  _1427_
timestamp 1678805552
transform 1 0 10752 0 1 46872
box -50 -56 1692 834
use sg13g2_dlhq_1  _1428_
timestamp 1678805552
transform 1 0 9888 0 1 45360
box -50 -56 1692 834
use sg13g2_dlhq_1  _1429_
timestamp 1678805552
transform 1 0 16032 0 -1 36288
box -50 -56 1692 834
use sg13g2_dlhq_1  _1430_
timestamp 1678805552
transform -1 0 16992 0 -1 37800
box -50 -56 1692 834
use sg13g2_dlhq_1  _1431_
timestamp 1678805552
transform 1 0 13248 0 1 24192
box -50 -56 1692 834
use sg13g2_dlhq_1  _1432_
timestamp 1678805552
transform 1 0 12096 0 -1 24192
box -50 -56 1692 834
use sg13g2_dlhq_1  _1433_
timestamp 1678805552
transform 1 0 4896 0 1 31752
box -50 -56 1692 834
use sg13g2_dlhq_1  _1434_
timestamp 1678805552
transform 1 0 3264 0 1 31752
box -50 -56 1692 834
use sg13g2_dlhq_1  _1435_
timestamp 1678805552
transform 1 0 13728 0 1 42336
box -50 -56 1692 834
use sg13g2_dlhq_1  _1436_
timestamp 1678805552
transform 1 0 13344 0 -1 42336
box -50 -56 1692 834
use sg13g2_dlhq_1  _1437_
timestamp 1678805552
transform 1 0 13632 0 1 40824
box -50 -56 1692 834
use sg13g2_dlhq_1  _1438_
timestamp 1678805552
transform 1 0 13728 0 -1 37800
box -50 -56 1692 834
use sg13g2_dlhq_1  _1439_
timestamp 1678805552
transform 1 0 15552 0 1 31752
box -50 -56 1692 834
use sg13g2_dlhq_1  _1440_
timestamp 1678805552
transform 1 0 15648 0 -1 33264
box -50 -56 1692 834
use sg13g2_dlhq_1  _1441_
timestamp 1678805552
transform 1 0 13632 0 -1 21168
box -50 -56 1692 834
use sg13g2_dlhq_1  _1442_
timestamp 1678805552
transform 1 0 12384 0 1 21168
box -50 -56 1692 834
use sg13g2_dlhq_1  _1443_
timestamp 1678805552
transform 1 0 12000 0 -1 21168
box -50 -56 1692 834
use sg13g2_dlhq_1  _1444_
timestamp 1678805552
transform -1 0 4608 0 -1 30240
box -50 -56 1692 834
use sg13g2_dlhq_1  _1445_
timestamp 1678805552
transform 1 0 1344 0 -1 30240
box -50 -56 1692 834
use sg13g2_dlhq_1  _1446_
timestamp 1678805552
transform 1 0 2784 0 1 30240
box -50 -56 1692 834
use sg13g2_dlhq_1  _1447_
timestamp 1678805552
transform 1 0 7488 0 1 39312
box -50 -56 1692 834
use sg13g2_dlhq_1  _1448_
timestamp 1678805552
transform 1 0 2784 0 1 37800
box -50 -56 1692 834
use sg13g2_dlhq_1  _1449_
timestamp 1678805552
transform 1 0 14688 0 1 30240
box -50 -56 1692 834
use sg13g2_dlhq_1  _1450_
timestamp 1678805552
transform 1 0 16224 0 1 28728
box -50 -56 1692 834
use sg13g2_dlhq_1  _1451_
timestamp 1678805552
transform 1 0 16224 0 1 39312
box -50 -56 1692 834
use sg13g2_dlhq_1  _1452_
timestamp 1678805552
transform 1 0 16128 0 -1 40824
box -50 -56 1692 834
use sg13g2_dlhq_1  _1453_
timestamp 1678805552
transform 1 0 1344 0 -1 42336
box -50 -56 1692 834
use sg13g2_dlhq_1  _1454_
timestamp 1678805552
transform 1 0 1152 0 1 40824
box -50 -56 1692 834
use sg13g2_dlhq_1  _1455_
timestamp 1678805552
transform 1 0 1152 0 1 31752
box -50 -56 1692 834
use sg13g2_dlhq_1  _1456_
timestamp 1678805552
transform 1 0 1536 0 -1 33264
box -50 -56 1692 834
use sg13g2_dlhq_1  _1457_
timestamp 1678805552
transform 1 0 9120 0 1 39312
box -50 -56 1692 834
use sg13g2_dlhq_1  _1458_
timestamp 1678805552
transform 1 0 9696 0 -1 40824
box -50 -56 1692 834
use sg13g2_dlhq_1  _1459_
timestamp 1678805552
transform 1 0 13056 0 1 27216
box -50 -56 1692 834
use sg13g2_dlhq_1  _1460_
timestamp 1678805552
transform 1 0 12000 0 1 28728
box -50 -56 1692 834
use sg13g2_dlhq_1  _1461_
timestamp 1678805552
transform 1 0 2784 0 1 40824
box -50 -56 1692 834
use sg13g2_dlhq_1  _1462_
timestamp 1678805552
transform 1 0 1152 0 1 37800
box -50 -56 1692 834
use sg13g2_dlhq_1  _1463_
timestamp 1678805552
transform 1 0 6240 0 1 46872
box -50 -56 1692 834
use sg13g2_dlhq_1  _1464_
timestamp 1678805552
transform 1 0 7872 0 -1 46872
box -50 -56 1692 834
use sg13g2_dlhq_1  _1465_
timestamp 1678805552
transform 1 0 10848 0 1 36288
box -50 -56 1692 834
use sg13g2_dlhq_1  _1466_
timestamp 1678805552
transform 1 0 10080 0 -1 36288
box -50 -56 1692 834
use sg13g2_dlhq_1  _1467_
timestamp 1678805552
transform 1 0 10464 0 -1 24192
box -50 -56 1692 834
use sg13g2_dlhq_1  _1468_
timestamp 1678805552
transform 1 0 11424 0 1 24192
box -50 -56 1692 834
use sg13g2_dlhq_1  _1469_
timestamp 1678805552
transform 1 0 8928 0 -1 39312
box -50 -56 1692 834
use sg13g2_dlhq_1  _1470_
timestamp 1678805552
transform -1 0 10656 0 -1 37800
box -50 -56 1692 834
use sg13g2_buf_1  _1473_
timestamp 1676381911
transform -1 0 19680 0 -1 93744
box -48 -56 432 834
use sg13g2_buf_1  _1474_
timestamp 1676381911
transform 1 0 16512 0 -1 68040
box -48 -56 432 834
use sg13g2_buf_1  _1475_
timestamp 1676381911
transform 1 0 14592 0 1 57456
box -48 -56 432 834
use sg13g2_buf_1  _1476_
timestamp 1676381911
transform -1 0 17568 0 -1 55944
box -48 -56 432 834
use sg13g2_buf_1  _1477_
timestamp 1676381911
transform 1 0 11136 0 1 69552
box -48 -56 432 834
use sg13g2_buf_1  _1478_
timestamp 1676381911
transform 1 0 1920 0 -1 57456
box -48 -56 432 834
use sg13g2_buf_1  _1479_
timestamp 1676381911
transform 1 0 2976 0 -1 55944
box -48 -56 432 834
use sg13g2_buf_1  _1480_
timestamp 1676381911
transform 1 0 1632 0 -1 54432
box -48 -56 432 834
use sg13g2_buf_1  _1481_
timestamp 1676381911
transform 1 0 1824 0 1 52920
box -48 -56 432 834
use sg13g2_buf_1  _1482_
timestamp 1676381911
transform 1 0 9312 0 -1 72576
box -48 -56 432 834
use sg13g2_buf_1  _1483_
timestamp 1676381911
transform 1 0 15168 0 1 66528
box -48 -56 432 834
use sg13g2_buf_1  _1484_
timestamp 1676381911
transform 1 0 16992 0 -1 84672
box -48 -56 432 834
use sg13g2_buf_1  _1485_
timestamp 1676381911
transform 1 0 13536 0 1 83160
box -48 -56 432 834
use sg13g2_buf_1  _1486_
timestamp 1676381911
transform 1 0 1824 0 1 87696
box -48 -56 432 834
use sg13g2_buf_1  _1487_
timestamp 1676381911
transform 1 0 4320 0 1 87696
box -48 -56 432 834
use sg13g2_buf_1  _1488_
timestamp 1676381911
transform 1 0 1824 0 1 71064
box -48 -56 432 834
use sg13g2_buf_1  _1489_
timestamp 1676381911
transform 1 0 9696 0 1 68040
box -48 -56 432 834
use sg13g2_buf_1  _1490_
timestamp 1676381911
transform 1 0 14016 0 1 57456
box -48 -56 432 834
use sg13g2_buf_1  _1491_
timestamp 1676381911
transform 1 0 12288 0 1 69552
box -48 -56 432 834
use sg13g2_buf_1  _1492_
timestamp 1676381911
transform 1 0 13344 0 -1 83160
box -48 -56 432 834
use sg13g2_buf_1  _1493_
timestamp 1676381911
transform 1 0 15072 0 -1 74088
box -48 -56 432 834
use sg13g2_buf_1  _1494_
timestamp 1676381911
transform 1 0 2208 0 1 87696
box -48 -56 432 834
use sg13g2_buf_1  _1495_
timestamp 1676381911
transform 1 0 8544 0 1 81648
box -48 -56 432 834
use sg13g2_buf_1  _1496_
timestamp 1676381911
transform 1 0 2304 0 1 89208
box -48 -56 432 834
use sg13g2_buf_1  _1497_
timestamp 1676381911
transform 1 0 9888 0 1 78624
box -48 -56 432 834
use sg13g2_buf_1  _1498_
timestamp 1676381911
transform 1 0 12768 0 1 80136
box -48 -56 432 834
use sg13g2_buf_1  _1499_
timestamp 1676381911
transform 1 0 9600 0 -1 80136
box -48 -56 432 834
use sg13g2_buf_1  _1500_
timestamp 1676381911
transform 1 0 14016 0 1 61992
box -48 -56 432 834
use sg13g2_buf_1  _1501_
timestamp 1676381911
transform -1 0 14496 0 1 60480
box -48 -56 432 834
use sg13g2_buf_1  _1502_
timestamp 1676381911
transform 1 0 2304 0 -1 90720
box -48 -56 432 834
use sg13g2_buf_1  _1503_
timestamp 1676381911
transform 1 0 9984 0 1 86184
box -48 -56 432 834
use sg13g2_buf_1  _1504_
timestamp 1676381911
transform 1 0 2976 0 1 84672
box -48 -56 432 834
use sg13g2_buf_1  _1505_
timestamp 1676381911
transform 1 0 7584 0 -1 60480
box -48 -56 432 834
use sg13g2_buf_1  _1506_
timestamp 1676381911
transform 1 0 10848 0 -1 75600
box -48 -56 432 834
use sg13g2_buf_1  _1507_
timestamp 1676381911
transform 1 0 3264 0 -1 86184
box -48 -56 432 834
use sg13g2_buf_1  _1508_
timestamp 1676381911
transform -1 0 17376 0 -1 90720
box -48 -56 432 834
use sg13g2_buf_1  _1509_
timestamp 1676381911
transform 1 0 9120 0 -1 89208
box -48 -56 432 834
use sg13g2_buf_1  _1510_
timestamp 1676381911
transform 1 0 17088 0 1 69552
box -48 -56 432 834
use sg13g2_buf_1  _1511_
timestamp 1676381911
transform -1 0 20352 0 1 63504
box -48 -56 432 834
use sg13g2_buf_1  _1512_
timestamp 1676381911
transform 1 0 12672 0 -1 58968
box -48 -56 432 834
use sg13g2_buf_1  _1513_
timestamp 1676381911
transform 1 0 12288 0 -1 60480
box -48 -56 432 834
use sg13g2_buf_1  _1514_
timestamp 1676381911
transform 1 0 6624 0 1 72576
box -48 -56 432 834
use sg13g2_buf_1  _1515_
timestamp 1676381911
transform 1 0 10368 0 1 86184
box -48 -56 432 834
use sg13g2_buf_1  _1516_
timestamp 1676381911
transform 1 0 2496 0 -1 3024
box -48 -56 432 834
use sg13g2_buf_1  _1517_
timestamp 1676381911
transform 1 0 16896 0 1 93744
box -48 -56 432 834
use sg13g2_buf_1  _1518_
timestamp 1676381911
transform 1 0 17280 0 1 93744
box -48 -56 432 834
use sg13g2_buf_1  _1519_
timestamp 1676381911
transform 1 0 16128 0 1 93744
box -48 -56 432 834
use sg13g2_buf_1  _1520_
timestamp 1676381911
transform 1 0 18048 0 1 93744
box -48 -56 432 834
use sg13g2_buf_1  _1521_
timestamp 1676381911
transform -1 0 20352 0 1 93744
box -48 -56 432 834
use sg13g2_buf_1  _1522_
timestamp 1676381911
transform 1 0 8160 0 -1 3024
box -48 -56 432 834
use sg13g2_buf_1  _1523_
timestamp 1676381911
transform -1 0 19968 0 1 93744
box -48 -56 432 834
use sg13g2_buf_1  _1524_
timestamp 1676381911
transform 1 0 18912 0 -1 93744
box -48 -56 432 834
use sg13g2_buf_1  _1525_
timestamp 1676381911
transform -1 0 19680 0 1 92232
box -48 -56 432 834
use sg13g2_buf_1  _1526_
timestamp 1676381911
transform -1 0 10464 0 1 55944
box -48 -56 432 834
use sg13g2_buf_1  _1527_
timestamp 1676381911
transform -1 0 15840 0 -1 74088
box -48 -56 432 834
use sg13g2_buf_1  _1528_
timestamp 1676381911
transform -1 0 16032 0 1 78624
box -48 -56 432 834
use sg13g2_buf_1  _1529_
timestamp 1676381911
transform -1 0 9024 0 1 87696
box -48 -56 432 834
use sg13g2_buf_1  _1530_
timestamp 1676381911
transform -1 0 8544 0 1 74088
box -48 -56 432 834
use sg13g2_buf_1  _1531_
timestamp 1676381911
transform -1 0 17376 0 -1 80136
box -48 -56 432 834
use sg13g2_buf_1  _1532_
timestamp 1676381911
transform -1 0 14208 0 1 71064
box -48 -56 432 834
use sg13g2_buf_1  _1533_
timestamp 1676381911
transform -1 0 9312 0 1 66528
box -48 -56 432 834
use sg13g2_buf_1  _1534_
timestamp 1676381911
transform -1 0 5184 0 1 51408
box -48 -56 432 834
use sg13g2_buf_1  _1535_
timestamp 1676381911
transform -1 0 14976 0 -1 74088
box -48 -56 432 834
use sg13g2_buf_1  _1536_
timestamp 1676381911
transform -1 0 14400 0 -1 75600
box -48 -56 432 834
use sg13g2_buf_1  _1537_
timestamp 1676381911
transform -1 0 10560 0 -1 77112
box -48 -56 432 834
use sg13g2_buf_1  _1538_
timestamp 1676381911
transform -1 0 4896 0 1 40824
box -48 -56 432 834
use sg13g2_buf_1  _1539_
timestamp 1676381911
transform -1 0 15072 0 1 48384
box -48 -56 432 834
use sg13g2_buf_1  _1540_
timestamp 1676381911
transform -1 0 13248 0 1 42336
box -48 -56 432 834
use sg13g2_buf_1  _1541_
timestamp 1676381911
transform 1 0 4032 0 -1 46872
box -48 -56 432 834
use sg13g2_buf_1  _1542_
timestamp 1676381911
transform 1 0 3552 0 -1 46872
box -48 -56 432 834
use sg13g2_buf_1  _1543_
timestamp 1676381911
transform -1 0 20352 0 1 48384
box -48 -56 432 834
use sg13g2_buf_1  _1544_
timestamp 1676381911
transform -1 0 16992 0 -1 31752
box -48 -56 432 834
use sg13g2_buf_1  _1545_
timestamp 1676381911
transform -1 0 9312 0 -1 40824
box -48 -56 432 834
use sg13g2_buf_1  _1546_
timestamp 1676381911
transform 1 0 2688 0 1 93744
box -48 -56 432 834
use sg13g2_buf_1  _1547_
timestamp 1676381911
transform 1 0 2688 0 -1 6048
box -48 -56 432 834
use sg13g2_buf_1  _1548_
timestamp 1676381911
transform 1 0 3072 0 1 93744
box -48 -56 432 834
use sg13g2_buf_1  _1549_
timestamp 1676381911
transform -1 0 8544 0 1 93744
box -48 -56 432 834
use sg13g2_buf_1  _1550_
timestamp 1676381911
transform 1 0 4608 0 -1 6048
box -48 -56 432 834
use sg13g2_buf_1  _1551_
timestamp 1676381911
transform -1 0 8064 0 1 90720
box -48 -56 432 834
use sg13g2_buf_1  _1552_
timestamp 1676381911
transform -1 0 8160 0 -1 92232
box -48 -56 432 834
use sg13g2_buf_1  _1553_
timestamp 1676381911
transform -1 0 8448 0 1 90720
box -48 -56 432 834
use sg13g2_buf_1  _1554_
timestamp 1676381911
transform 1 0 4896 0 -1 28728
box -48 -56 432 834
use sg13g2_buf_1  _1555_
timestamp 1676381911
transform -1 0 16608 0 -1 21168
box -48 -56 432 834
use sg13g2_buf_1  _1556_
timestamp 1676381911
transform -1 0 17760 0 -1 37800
box -48 -56 432 834
use sg13g2_buf_1  _1557_
timestamp 1676381911
transform -1 0 15552 0 -1 36288
box -48 -56 432 834
use sg13g2_buf_1  _1558_
timestamp 1676381911
transform -1 0 9792 0 1 63504
box -48 -56 432 834
use sg13g2_buf_1  _1559_
timestamp 1676381911
transform -1 0 17856 0 -1 81648
box -48 -56 432 834
use sg13g2_buf_1  _1560_
timestamp 1676381911
transform -1 0 14304 0 1 83160
box -48 -56 432 834
use sg13g2_buf_1  _1561_
timestamp 1676381911
transform 1 0 8544 0 -1 81648
box -48 -56 432 834
use sg13g2_buf_1  _1562_
timestamp 1676381911
transform -1 0 20064 0 -1 93744
box -48 -56 432 834
use sg13g2_buf_1  _1563_
timestamp 1676381911
transform -1 0 12960 0 1 58968
box -48 -56 432 834
use sg13g2_buf_1  _1564_
timestamp 1676381911
transform -1 0 17088 0 1 69552
box -48 -56 432 834
use sg13g2_buf_1  _1565_
timestamp 1676381911
transform -1 0 12960 0 -1 66528
box -48 -56 432 834
use sg13g2_buf_1  _1566_
timestamp 1676381911
transform -1 0 5664 0 1 75600
box -48 -56 432 834
use sg13g2_buf_1  _1567_
timestamp 1676381911
transform -1 0 4416 0 1 65016
box -48 -56 432 834
use sg13g2_buf_1  _1568_
timestamp 1676381911
transform -1 0 18144 0 1 52920
box -48 -56 432 834
use sg13g2_buf_1  _1569_
timestamp 1676381911
transform -1 0 14688 0 1 63504
box -48 -56 432 834
use sg13g2_buf_1  _1570_
timestamp 1676381911
transform -1 0 5760 0 1 55944
box -48 -56 432 834
use sg13g2_buf_1  _1571_
timestamp 1676381911
transform -1 0 3648 0 1 69552
box -48 -56 432 834
use sg13g2_buf_1  _1572_
timestamp 1676381911
transform -1 0 15840 0 1 63504
box -48 -56 432 834
use sg13g2_buf_1  _1573_
timestamp 1676381911
transform -1 0 19776 0 -1 52920
box -48 -56 432 834
use sg13g2_buf_1  _1574_
timestamp 1676381911
transform -1 0 3648 0 1 58968
box -48 -56 432 834
use sg13g2_buf_1  _1575_
timestamp 1676381911
transform -1 0 5280 0 -1 68040
box -48 -56 432 834
use sg13g2_buf_1  _1576_
timestamp 1676381911
transform -1 0 17376 0 -1 54432
box -48 -56 432 834
use sg13g2_buf_1  _1577_
timestamp 1676381911
transform -1 0 19776 0 1 68040
box -48 -56 432 834
use sg13g2_buf_1  _1578_
timestamp 1676381911
transform -1 0 6240 0 1 60480
box -48 -56 432 834
use sg13g2_buf_1  _1579_
timestamp 1676381911
transform -1 0 5856 0 -1 72576
box -48 -56 432 834
use sg13g2_buf_1  _1580_
timestamp 1676381911
transform -1 0 15840 0 -1 61992
box -48 -56 432 834
use sg13g2_buf_1  _1581_
timestamp 1676381911
transform -1 0 18144 0 -1 54432
box -48 -56 432 834
use sg13g2_buf_1  _1582_
timestamp 1676381911
transform -1 0 4032 0 1 58968
box -48 -56 432 834
use sg13g2_buf_1  _1583_
timestamp 1676381911
transform -1 0 10368 0 -1 69552
box -48 -56 432 834
use sg13g2_buf_1  _1584_
timestamp 1676381911
transform -1 0 16032 0 -1 71064
box -48 -56 432 834
use sg13g2_buf_1  _1585_
timestamp 1676381911
transform -1 0 18528 0 -1 86184
box -48 -56 432 834
use sg13g2_buf_1  _1586_
timestamp 1676381911
transform -1 0 6528 0 -1 65016
box -48 -56 432 834
use sg13g2_buf_1  _1587_
timestamp 1676381911
transform 1 0 6432 0 1 75600
box -48 -56 432 834
use sg13g2_buf_1  _1588_
timestamp 1676381911
transform -1 0 17088 0 -1 66528
box -48 -56 432 834
use sg13g2_buf_1  _1589_
timestamp 1676381911
transform -1 0 18720 0 -1 71064
box -48 -56 432 834
use sg13g2_buf_1  _1590_
timestamp 1676381911
transform -1 0 5856 0 1 60480
box -48 -56 432 834
use sg13g2_buf_1  _1591_
timestamp 1676381911
transform -1 0 8544 0 -1 72576
box -48 -56 432 834
use sg13g2_buf_1  _1592_
timestamp 1676381911
transform -1 0 16416 0 1 69552
box -48 -56 432 834
use sg13g2_buf_1  _1593_
timestamp 1676381911
transform -1 0 16320 0 1 63504
box -48 -56 432 834
use sg13g2_buf_1  _1594_
timestamp 1676381911
transform -1 0 7872 0 -1 61992
box -48 -56 432 834
use sg13g2_buf_1  _1595_
timestamp 1676381911
transform 1 0 6240 0 -1 71064
box -48 -56 432 834
use sg13g2_buf_1  _1596_
timestamp 1676381911
transform -1 0 16512 0 -1 69552
box -48 -56 432 834
use sg13g2_buf_1  _1597_
timestamp 1676381911
transform -1 0 15360 0 1 57456
box -48 -56 432 834
use sg13g2_buf_1  _1598_
timestamp 1676381911
transform -1 0 7104 0 -1 57456
box -48 -56 432 834
use sg13g2_buf_1  _1599_
timestamp 1676381911
transform -1 0 5376 0 -1 69552
box -48 -56 432 834
use sg13g2_buf_1  _1600_
timestamp 1676381911
transform -1 0 14880 0 1 65016
box -48 -56 432 834
use sg13g2_buf_1  _1601_
timestamp 1676381911
transform -1 0 16224 0 -1 61992
box -48 -56 432 834
use sg13g2_buf_1  _1602_
timestamp 1676381911
transform -1 0 6144 0 -1 58968
box -48 -56 432 834
use sg13g2_buf_1  _1603_
timestamp 1676381911
transform -1 0 7008 0 -1 71064
box -48 -56 432 834
use sg13g2_buf_1  _1604_
timestamp 1676381911
transform -1 0 17472 0 -1 66528
box -48 -56 432 834
use sg13g2_buf_1  _1605_
timestamp 1676381911
transform -1 0 20352 0 1 66528
box -48 -56 432 834
use sg13g2_buf_1  _1606_
timestamp 1676381911
transform -1 0 5664 0 -1 61992
box -48 -56 432 834
use sg13g2_buf_1  _1607_
timestamp 1676381911
transform -1 0 5472 0 -1 72576
box -48 -56 432 834
use sg13g2_buf_1  _1608_
timestamp 1676381911
transform -1 0 14496 0 1 68040
box -48 -56 432 834
use sg13g2_buf_1  _1609_
timestamp 1676381911
transform -1 0 17664 0 1 55944
box -48 -56 432 834
use sg13g2_buf_1  _1610_
timestamp 1676381911
transform -1 0 8544 0 1 58968
box -48 -56 432 834
use sg13g2_buf_1  _1611_
timestamp 1676381911
transform 1 0 2976 0 -1 42336
box -48 -56 432 834
use sg13g2_buf_1  _1612_
timestamp 1676381911
transform 1 0 8928 0 1 28728
box -48 -56 432 834
use sg13g2_buf_1  _1613_
timestamp 1676381911
transform 1 0 6048 0 -1 18144
box -48 -56 432 834
use sg13g2_buf_1  _1614_
timestamp 1676381911
transform 1 0 1920 0 1 6048
box -48 -56 432 834
use sg13g2_buf_1  _1615_
timestamp 1676381911
transform 1 0 4224 0 -1 6048
box -48 -56 432 834
use sg13g2_buf_1  _1616_
timestamp 1676381911
transform 1 0 7584 0 -1 27216
box -48 -56 432 834
use sg13g2_buf_1  _1617_
timestamp 1676381911
transform 1 0 10080 0 -1 28728
box -48 -56 432 834
use sg13g2_buf_1  _1618_
timestamp 1676381911
transform 1 0 1920 0 1 21168
box -48 -56 432 834
use sg13g2_buf_1  _1619_
timestamp 1676381911
transform 1 0 1824 0 -1 10584
box -48 -56 432 834
use sg13g2_buf_1  _1620_
timestamp 1676381911
transform 1 0 6816 0 -1 16632
box -48 -56 432 834
use sg13g2_buf_1  _1621_
timestamp 1676381911
transform 1 0 15840 0 1 7560
box -48 -56 432 834
use sg13g2_buf_1  _1622_
timestamp 1676381911
transform -1 0 15648 0 -1 9072
box -48 -56 432 834
use sg13g2_buf_1  _1623_
timestamp 1676381911
transform 1 0 12000 0 -1 34776
box -48 -56 432 834
use sg13g2_buf_1  _1624_
timestamp 1676381911
transform 1 0 10464 0 1 30240
box -48 -56 432 834
use sg13g2_buf_1  _1625_
timestamp 1676381911
transform 1 0 7104 0 1 15120
box -48 -56 432 834
use sg13g2_buf_1  _1626_
timestamp 1676381911
transform 1 0 4704 0 1 18144
box -48 -56 432 834
use sg13g2_buf_1  _1627_
timestamp 1676381911
transform 1 0 16992 0 -1 37800
box -48 -56 432 834
use sg13g2_buf_1  _1628_
timestamp 1676381911
transform 1 0 15360 0 1 37800
box -48 -56 432 834
use sg13g2_buf_1  _1629_
timestamp 1676381911
transform 1 0 3168 0 1 10584
box -48 -56 432 834
use sg13g2_buf_1  _1630_
timestamp 1676381911
transform 1 0 16704 0 -1 34776
box -48 -56 432 834
use sg13g2_buf_1  _1631_
timestamp 1676381911
transform 1 0 10944 0 -1 27216
box -48 -56 432 834
use sg13g2_buf_1  _1632_
timestamp 1676381911
transform 1 0 13632 0 1 25704
box -48 -56 432 834
use sg13g2_buf_1  _1633_
timestamp 1676381911
transform 1 0 1920 0 1 39312
box -48 -56 432 834
use sg13g2_buf_1  _1634_
timestamp 1676381911
transform 1 0 8160 0 -1 40824
box -48 -56 432 834
use sg13g2_buf_1  _1635_
timestamp 1676381911
transform 1 0 10944 0 -1 22680
box -48 -56 432 834
use sg13g2_buf_1  _1636_
timestamp 1676381911
transform 1 0 9024 0 1 24192
box -48 -56 432 834
use sg13g2_buf_1  _1637_
timestamp 1676381911
transform 1 0 11616 0 -1 45360
box -48 -56 432 834
use sg13g2_buf_1  _1638_
timestamp 1676381911
transform 1 0 11520 0 1 45360
box -48 -56 432 834
use sg13g2_buf_1  _1639_
timestamp 1676381911
transform 1 0 14976 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  _1640_
timestamp 1676381911
transform 1 0 15744 0 -1 40824
box -48 -56 432 834
use sg13g2_buf_1  _1641_
timestamp 1676381911
transform 1 0 3936 0 1 10584
box -48 -56 432 834
use sg13g2_buf_1  _1642_
timestamp 1676381911
transform 1 0 3168 0 -1 9072
box -48 -56 432 834
use sg13g2_buf_1  _1643_
timestamp 1676381911
transform 1 0 6912 0 1 31752
box -48 -56 432 834
use sg13g2_buf_1  _1644_
timestamp 1676381911
transform -1 0 16224 0 -1 24192
box -48 -56 432 834
use sg13g2_buf_1  _1645_
timestamp 1676381911
transform -1 0 18432 0 1 34776
box -48 -56 432 834
use sg13g2_buf_1  _1646_
timestamp 1676381911
transform -1 0 12864 0 -1 46872
box -48 -56 432 834
use sg13g2_buf_1  _1647_
timestamp 1676381911
transform 1 0 2016 0 -1 43848
box -48 -56 432 834
use sg13g2_buf_1  _1648_
timestamp 1676381911
transform -1 0 17664 0 -1 33264
box -48 -56 432 834
use sg13g2_buf_1  _1649_
timestamp 1676381911
transform -1 0 13536 0 -1 43848
box -48 -56 432 834
use sg13g2_buf_1  _1650_
timestamp 1676381911
transform 1 0 7296 0 1 31752
box -48 -56 432 834
use sg13g2_buf_1  _1651_
timestamp 1676381911
transform 1 0 4704 0 -1 34776
box -48 -56 432 834
use sg13g2_buf_1  _1652_
timestamp 1676381911
transform -1 0 17952 0 -1 24192
box -48 -56 432 834
use sg13g2_buf_1  _1653_
timestamp 1676381911
transform -1 0 18240 0 -1 27216
box -48 -56 432 834
use sg13g2_buf_1  _1654_
timestamp 1676381911
transform 1 0 8256 0 1 24192
box -48 -56 432 834
use sg13g2_buf_1  _1655_
timestamp 1676381911
transform 1 0 5856 0 -1 55944
box -48 -56 432 834
use sg13g2_buf_1  _1656_
timestamp 1676381911
transform -1 0 17760 0 1 52920
box -48 -56 432 834
use sg13g2_buf_1  _1657_
timestamp 1676381911
transform -1 0 12672 0 1 63504
box -48 -56 432 834
use sg13g2_buf_1  _1658_
timestamp 1676381911
transform 1 0 7296 0 1 68040
box -48 -56 432 834
use sg13g2_buf_1  _1659_
timestamp 1676381911
transform 1 0 3744 0 1 48384
box -48 -56 432 834
use sg13g2_buf_1  _1660_
timestamp 1676381911
transform -1 0 14880 0 1 71064
box -48 -56 432 834
use sg13g2_buf_1  _1661_
timestamp 1676381911
transform -1 0 17952 0 -1 49896
box -48 -56 432 834
use sg13g2_buf_1  _1662_
timestamp 1676381911
transform 1 0 10560 0 -1 77112
box -48 -56 432 834
use sg13g2_buf_1  _1663_
timestamp 1676381911
transform -1 0 14688 0 1 93744
box -48 -56 432 834
use sg13g2_buf_1  _1664_
timestamp 1676381911
transform 1 0 2016 0 -1 3024
box -48 -56 432 834
use sg13g2_buf_1  _1665_
timestamp 1676381911
transform -1 0 15072 0 1 93744
box -48 -56 432 834
use sg13g2_buf_1  _1666_
timestamp 1676381911
transform 1 0 1632 0 -1 3024
box -48 -56 432 834
use sg13g2_buf_1  _1667_
timestamp 1676381911
transform -1 0 18048 0 1 93744
box -48 -56 432 834
use sg13g2_buf_1  _1668_
timestamp 1676381911
transform -1 0 16896 0 1 93744
box -48 -56 432 834
use sg13g2_buf_1  _1669_
timestamp 1676381911
transform -1 0 15456 0 1 93744
box -48 -56 432 834
use sg13g2_buf_1  _1670_
timestamp 1676381911
transform 1 0 2304 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  _1671_
timestamp 1676381911
transform 1 0 10176 0 1 52920
box -48 -56 432 834
use sg13g2_buf_1  _1672_
timestamp 1676381911
transform -1 0 18528 0 -1 58968
box -48 -56 432 834
use sg13g2_buf_1  _1673_
timestamp 1676381911
transform -1 0 16032 0 1 83160
box -48 -56 432 834
use sg13g2_buf_1  _1674_
timestamp 1676381911
transform 1 0 7392 0 1 84672
box -48 -56 432 834
use sg13g2_buf_1  _1675_
timestamp 1676381911
transform 1 0 4416 0 1 13608
box -48 -56 432 834
use sg13g2_buf_1  _1676_
timestamp 1676381911
transform -1 0 19776 0 -1 18144
box -48 -56 432 834
use sg13g2_buf_1  _1677_
timestamp 1676381911
transform 1 0 14592 0 1 28728
box -48 -56 432 834
use sg13g2_buf_1  _1678_
timestamp 1676381911
transform 1 0 12480 0 -1 40824
box -48 -56 432 834
use sg13g2_buf_1  _1679_
timestamp 1676381911
transform -1 0 9792 0 1 18144
box -48 -56 432 834
use sg13g2_buf_1  _1680_
timestamp 1676381911
transform -1 0 14496 0 -1 18144
box -48 -56 432 834
use sg13g2_buf_1  _1681_
timestamp 1676381911
transform -1 0 14688 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  _1682_
timestamp 1676381911
transform -1 0 11616 0 -1 21168
box -48 -56 432 834
use sg13g2_buf_1  _1683_
timestamp 1676381911
transform -1 0 8448 0 -1 10584
box -48 -56 432 834
use sg13g2_buf_1  _1684_
timestamp 1676381911
transform -1 0 17664 0 1 6048
box -48 -56 432 834
use sg13g2_buf_1  _1685_
timestamp 1676381911
transform -1 0 10944 0 -1 12096
box -48 -56 432 834
use sg13g2_buf_1  _1686_
timestamp 1676381911
transform -1 0 4704 0 1 18144
box -48 -56 432 834
use sg13g2_buf_1  _1687_
timestamp 1676381911
transform -1 0 4992 0 -1 12096
box -48 -56 432 834
use sg13g2_buf_1  _1688_
timestamp 1676381911
transform -1 0 10464 0 -1 6048
box -48 -56 432 834
use sg13g2_buf_1  _1689_
timestamp 1676381911
transform -1 0 19776 0 -1 7560
box -48 -56 432 834
use sg13g2_buf_1  _1690_
timestamp 1676381911
transform -1 0 6624 0 1 15120
box -48 -56 432 834
use sg13g2_buf_1  _1691_
timestamp 1676381911
transform -1 0 8544 0 -1 9072
box -48 -56 432 834
use sg13g2_buf_1  _1692_
timestamp 1676381911
transform -1 0 16224 0 1 4536
box -48 -56 432 834
use sg13g2_buf_1  _1693_
timestamp 1676381911
transform -1 0 10368 0 1 13608
box -48 -56 432 834
use sg13g2_buf_1  _1694_
timestamp 1676381911
transform -1 0 8640 0 -1 19656
box -48 -56 432 834
use sg13g2_buf_1  _1695_
timestamp 1676381911
transform -1 0 4608 0 -1 12096
box -48 -56 432 834
use sg13g2_buf_1  _1696_
timestamp 1676381911
transform -1 0 10656 0 1 6048
box -48 -56 432 834
use sg13g2_buf_1  _1697_
timestamp 1676381911
transform -1 0 17760 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  _1698_
timestamp 1676381911
transform -1 0 6336 0 -1 16632
box -48 -56 432 834
use sg13g2_buf_1  _1699_
timestamp 1676381911
transform -1 0 11232 0 1 16632
box -48 -56 432 834
use sg13g2_buf_1  _1700_
timestamp 1676381911
transform -1 0 17856 0 -1 13608
box -48 -56 432 834
use sg13g2_buf_1  _1701_
timestamp 1676381911
transform -1 0 15648 0 -1 12096
box -48 -56 432 834
use sg13g2_buf_1  _1702_
timestamp 1676381911
transform -1 0 11904 0 -1 30240
box -48 -56 432 834
use sg13g2_buf_1  _1703_
timestamp 1676381911
transform -1 0 6432 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  _1704_
timestamp 1676381911
transform -1 0 13056 0 1 4536
box -48 -56 432 834
use sg13g2_buf_1  _1705_
timestamp 1676381911
transform -1 0 14976 0 -1 18144
box -48 -56 432 834
use sg13g2_buf_1  _1706_
timestamp 1676381911
transform -1 0 8256 0 -1 19656
box -48 -56 432 834
use sg13g2_buf_1  _1707_
timestamp 1676381911
transform -1 0 7584 0 1 12096
box -48 -56 432 834
use sg13g2_buf_1  _1708_
timestamp 1676381911
transform -1 0 12864 0 1 19656
box -48 -56 432 834
use sg13g2_buf_1  _1709_
timestamp 1676381911
transform -1 0 17376 0 -1 18144
box -48 -56 432 834
use sg13g2_buf_1  _1710_
timestamp 1676381911
transform 1 0 4224 0 1 22680
box -48 -56 432 834
use sg13g2_buf_1  _1711_
timestamp 1676381911
transform -1 0 9792 0 1 13608
box -48 -56 432 834
use sg13g2_buf_1  _1712_
timestamp 1676381911
transform -1 0 18240 0 1 7560
box -48 -56 432 834
use sg13g2_buf_1  _1713_
timestamp 1676381911
transform -1 0 16800 0 -1 12096
box -48 -56 432 834
use sg13g2_buf_1  _1714_
timestamp 1676381911
transform -1 0 7104 0 1 19656
box -48 -56 432 834
use sg13g2_buf_1  _1715_
timestamp 1676381911
transform -1 0 4128 0 -1 9072
box -48 -56 432 834
use sg13g2_buf_1  _1716_
timestamp 1676381911
transform -1 0 13440 0 1 4536
box -48 -56 432 834
use sg13g2_buf_1  _1717_
timestamp 1676381911
transform -1 0 17664 0 1 10584
box -48 -56 432 834
use sg13g2_buf_1  _1718_
timestamp 1676381911
transform -1 0 5952 0 -1 16632
box -48 -56 432 834
use sg13g2_buf_1  _1719_
timestamp 1676381911
transform -1 0 7008 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  _1720_
timestamp 1676381911
transform -1 0 15168 0 1 6048
box -48 -56 432 834
use sg13g2_buf_1  _1721_
timestamp 1676381911
transform -1 0 16032 0 -1 15120
box -48 -56 432 834
use sg13g2_buf_1  _1722_
timestamp 1676381911
transform 1 0 5280 0 -1 18144
box -48 -56 432 834
use sg13g2_buf_1  _1723_
timestamp 1676381911
transform -1 0 8064 0 -1 13608
box -48 -56 432 834
use sg13g2_buf_1  _1724_
timestamp 1676381911
transform -1 0 11520 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  _1725_
timestamp 1676381911
transform -1 0 17376 0 1 12096
box -48 -56 432 834
use sg13g2_buf_1  _1726_
timestamp 1676381911
transform -1 0 7296 0 -1 25704
box -48 -56 432 834
use sg13g2_buf_1  fanout623
timestamp 1676381911
transform 1 0 8928 0 -1 68040
box -48 -56 432 834
use sg13g2_buf_1  fanout624
timestamp 1676381911
transform -1 0 17184 0 1 68040
box -48 -56 432 834
use sg13g2_buf_1  fanout625
timestamp 1676381911
transform 1 0 14976 0 -1 60480
box -48 -56 432 834
use sg13g2_buf_1  fanout626
timestamp 1676381911
transform 1 0 4896 0 1 66528
box -48 -56 432 834
use sg13g2_buf_1  fanout627
timestamp 1676381911
transform -1 0 4896 0 1 48384
box -48 -56 432 834
use sg13g2_buf_1  fanout628
timestamp 1676381911
transform -1 0 5856 0 -1 55944
box -48 -56 432 834
use sg13g2_buf_1  fanout629
timestamp 1676381911
transform 1 0 13248 0 -1 69552
box -48 -56 432 834
use sg13g2_buf_1  fanout630
timestamp 1676381911
transform -1 0 19392 0 -1 52920
box -48 -56 432 834
use sg13g2_buf_1  fanout631
timestamp 1676381911
transform 1 0 8544 0 -1 72576
box -48 -56 432 834
use sg13g2_buf_1  fanout632
timestamp 1676381911
transform -1 0 8544 0 1 37800
box -48 -56 432 834
use sg13g2_buf_1  fanout633
timestamp 1676381911
transform -1 0 16320 0 -1 30240
box -48 -56 432 834
use sg13g2_buf_1  fanout634
timestamp 1676381911
transform -1 0 18144 0 1 22680
box -48 -56 432 834
use sg13g2_buf_1  fanout635
timestamp 1676381911
transform 1 0 4896 0 -1 19656
box -48 -56 432 834
use sg13g2_buf_1  fanout636
timestamp 1676381911
transform 1 0 4416 0 -1 46872
box -48 -56 432 834
use sg13g2_buf_1  fanout637
timestamp 1676381911
transform 1 0 4128 0 1 36288
box -48 -56 432 834
use sg13g2_buf_1  fanout638
timestamp 1676381911
transform -1 0 15552 0 1 28728
box -48 -56 432 834
use sg13g2_buf_1  fanout639
timestamp 1676381911
transform -1 0 16416 0 -1 19656
box -48 -56 432 834
use sg13g2_buf_1  fanout640
timestamp 1676381911
transform 1 0 5664 0 1 24192
box -48 -56 432 834
use sg13g2_buf_1  fanout641
timestamp 1676381911
transform 1 0 11712 0 1 31752
box -48 -56 432 834
use sg13g2_buf_1  fanout642
timestamp 1676381911
transform -1 0 10656 0 1 43848
box -48 -56 432 834
use sg13g2_buf_1  fanout643
timestamp 1676381911
transform 1 0 9600 0 -1 48384
box -48 -56 432 834
use sg13g2_buf_1  fanout644
timestamp 1676381911
transform 1 0 8544 0 1 84672
box -48 -56 432 834
use sg13g2_buf_1  fanout645
timestamp 1676381911
transform -1 0 8928 0 1 48384
box -48 -56 432 834
use sg13g2_buf_1  fanout646
timestamp 1676381911
transform -1 0 9312 0 1 48384
box -48 -56 432 834
use sg13g2_buf_1  fanout647
timestamp 1676381911
transform 1 0 13056 0 -1 37800
box -48 -56 432 834
use sg13g2_buf_1  fanout648
timestamp 1676381911
transform -1 0 13920 0 -1 25704
box -48 -56 432 834
use sg13g2_buf_1  fanout649
timestamp 1676381911
transform -1 0 4800 0 1 28728
box -48 -56 432 834
use sg13g2_buf_1  fanout650
timestamp 1676381911
transform 1 0 14784 0 1 36288
box -48 -56 432 834
use sg13g2_buf_1  fanout651
timestamp 1676381911
transform -1 0 15168 0 1 37800
box -48 -56 432 834
use sg13g2_buf_1  fanout652
timestamp 1676381911
transform -1 0 12864 0 -1 75600
box -48 -56 432 834
use sg13g2_buf_1  fanout653
timestamp 1676381911
transform 1 0 12672 0 1 77112
box -48 -56 432 834
use sg13g2_buf_1  fanout654
timestamp 1676381911
transform 1 0 13248 0 -1 75600
box -48 -56 432 834
use sg13g2_buf_1  fanout655
timestamp 1676381911
transform -1 0 12672 0 1 77112
box -48 -56 432 834
use sg13g2_buf_1  fanout656
timestamp 1676381911
transform 1 0 12864 0 -1 75600
box -48 -56 432 834
use sg13g2_buf_1  fanout657
timestamp 1676381911
transform -1 0 14496 0 -1 60480
box -48 -56 432 834
use sg13g2_buf_1  fanout658
timestamp 1676381911
transform 1 0 14784 0 -1 9072
box -48 -56 432 834
use sg13g2_buf_1  fanout659
timestamp 1676381911
transform -1 0 16512 0 1 19656
box -48 -56 432 834
use sg13g2_buf_1  fanout660
timestamp 1676381911
transform 1 0 16800 0 -1 24192
box -48 -56 432 834
use sg13g2_buf_1  fanout661
timestamp 1676381911
transform -1 0 12000 0 1 22680
box -48 -56 432 834
use sg13g2_buf_1  fanout662
timestamp 1676381911
transform 1 0 12192 0 -1 30240
box -48 -56 432 834
use sg13g2_buf_1  fanout663
timestamp 1676381911
transform 1 0 12096 0 1 52920
box -48 -56 432 834
use sg13g2_buf_1  fanout664
timestamp 1676381911
transform 1 0 11040 0 -1 80136
box -48 -56 432 834
use sg13g2_buf_1  fanout665
timestamp 1676381911
transform -1 0 11616 0 -1 72576
box -48 -56 432 834
use sg13g2_buf_1  fanout666
timestamp 1676381911
transform -1 0 11424 0 -1 71064
box -48 -56 432 834
use sg13g2_buf_1  fanout667
timestamp 1676381911
transform -1 0 12480 0 -1 51408
box -48 -56 432 834
use sg13g2_buf_1  fanout668
timestamp 1676381911
transform -1 0 12384 0 1 49896
box -48 -56 432 834
use sg13g2_buf_1  fanout669
timestamp 1676381911
transform -1 0 8544 0 1 12096
box -48 -56 432 834
use sg13g2_buf_1  fanout670
timestamp 1676381911
transform 1 0 4800 0 1 12096
box -48 -56 432 834
use sg13g2_buf_1  fanout671
timestamp 1676381911
transform 1 0 16032 0 -1 12096
box -48 -56 432 834
use sg13g2_buf_1  fanout672
timestamp 1676381911
transform 1 0 4320 0 1 12096
box -48 -56 432 834
use sg13g2_buf_1  fanout673
timestamp 1676381911
transform 1 0 3168 0 -1 13608
box -48 -56 432 834
use sg13g2_buf_1  fanout674
timestamp 1676381911
transform -1 0 2880 0 -1 51408
box -48 -56 432 834
use sg13g2_buf_1  fanout675
timestamp 1676381911
transform 1 0 13536 0 1 74088
box -48 -56 432 834
use sg13g2_buf_1  fanout676
timestamp 1676381911
transform -1 0 3456 0 1 65016
box -48 -56 432 834
use sg13g2_buf_1  fanout677
timestamp 1676381911
transform 1 0 13056 0 1 66528
box -48 -56 432 834
use sg13g2_buf_1  fanout678
timestamp 1676381911
transform 1 0 2016 0 1 51408
box -48 -56 432 834
use sg13g2_buf_1  fanout679
timestamp 1676381911
transform 1 0 2400 0 1 51408
box -48 -56 432 834
use sg13g2_buf_1  fanout680
timestamp 1676381911
transform -1 0 3168 0 1 6048
box -48 -56 432 834
use sg13g2_buf_1  fanout681
timestamp 1676381911
transform 1 0 6336 0 -1 16632
box -48 -56 432 834
use sg13g2_buf_1  fanout682
timestamp 1676381911
transform 1 0 10464 0 1 13608
box -48 -56 432 834
use sg13g2_buf_1  fanout683
timestamp 1676381911
transform 1 0 10560 0 -1 15120
box -48 -56 432 834
use sg13g2_buf_1  fanout684
timestamp 1676381911
transform -1 0 10752 0 -1 18144
box -48 -56 432 834
use sg13g2_buf_1  fanout685
timestamp 1676381911
transform -1 0 6432 0 1 63504
box -48 -56 432 834
use sg13g2_buf_1  fanout686
timestamp 1676381911
transform -1 0 6048 0 1 63504
box -48 -56 432 834
use sg13g2_buf_1  fanout687
timestamp 1676381911
transform 1 0 13632 0 1 61992
box -48 -56 432 834
use sg13g2_buf_1  fanout688
timestamp 1676381911
transform 1 0 13248 0 -1 63504
box -48 -56 432 834
use sg13g2_buf_1  fanout689
timestamp 1676381911
transform -1 0 12096 0 -1 61992
box -48 -56 432 834
use sg13g2_buf_1  fanout690
timestamp 1676381911
transform 1 0 12480 0 1 51408
box -48 -56 432 834
use sg13g2_buf_1  fanout691
timestamp 1676381911
transform -1 0 11520 0 1 49896
box -48 -56 432 834
use sg13g2_buf_1  fanout692
timestamp 1676381911
transform -1 0 7872 0 -1 19656
box -48 -56 432 834
use sg13g2_buf_1  fanout693
timestamp 1676381911
transform 1 0 12864 0 1 19656
box -48 -56 432 834
use sg13g2_buf_1  fanout694
timestamp 1676381911
transform -1 0 18336 0 -1 24192
box -48 -56 432 834
use sg13g2_buf_1  fanout695
timestamp 1676381911
transform -1 0 12480 0 -1 28728
box -48 -56 432 834
use sg13g2_buf_1  fanout696
timestamp 1676381911
transform -1 0 12864 0 1 52920
box -48 -56 432 834
use sg13g2_buf_1  fanout697
timestamp 1676381911
transform 1 0 6528 0 -1 66528
box -48 -56 432 834
use sg13g2_buf_1  fanout698
timestamp 1676381911
transform 1 0 11712 0 1 65016
box -48 -56 432 834
use sg13g2_buf_1  fanout699
timestamp 1676381911
transform -1 0 12480 0 1 65016
box -48 -56 432 834
use sg13g2_buf_1  fanout700
timestamp 1676381911
transform 1 0 15840 0 -1 74088
box -48 -56 432 834
use sg13g2_buf_1  fanout701
timestamp 1676381911
transform 1 0 15552 0 1 66528
box -48 -56 432 834
use sg13g2_buf_1  fanout702
timestamp 1676381911
transform -1 0 13248 0 -1 54432
box -48 -56 432 834
use sg13g2_buf_1  fanout703
timestamp 1676381911
transform 1 0 17184 0 1 31752
box -48 -56 432 834
use sg13g2_buf_1  fanout704
timestamp 1676381911
transform 1 0 15744 0 1 37800
box -48 -56 432 834
use sg13g2_buf_1  fanout705
timestamp 1676381911
transform -1 0 16416 0 -1 39312
box -48 -56 432 834
use sg13g2_buf_1  fanout706
timestamp 1676381911
transform 1 0 15360 0 -1 40824
box -48 -56 432 834
use sg13g2_buf_1  fanout707
timestamp 1676381911
transform 1 0 16416 0 -1 39312
box -48 -56 432 834
use sg13g2_buf_1  fanout708
timestamp 1676381911
transform 1 0 13056 0 -1 58968
box -48 -56 432 834
use sg13g2_buf_1  fanout709
timestamp 1676381911
transform -1 0 13536 0 -1 60480
box -48 -56 432 834
use sg13g2_buf_1  fanout710
timestamp 1676381911
transform -1 0 9888 0 -1 89208
box -48 -56 432 834
use sg13g2_buf_1  fanout711
timestamp 1676381911
transform 1 0 12480 0 1 87696
box -48 -56 432 834
use sg13g2_buf_1  fanout712
timestamp 1676381911
transform -1 0 10272 0 -1 89208
box -48 -56 432 834
use sg13g2_buf_1  fanout713
timestamp 1676381911
transform -1 0 13152 0 -1 60480
box -48 -56 432 834
use sg13g2_buf_1  fanout714
timestamp 1676381911
transform -1 0 17856 0 -1 27216
box -48 -56 432 834
use sg13g2_buf_1  fanout715
timestamp 1676381911
transform -1 0 15936 0 -1 30240
box -48 -56 432 834
use sg13g2_buf_1  fanout716
timestamp 1676381911
transform 1 0 17760 0 1 43848
box -48 -56 432 834
use sg13g2_buf_1  fanout717
timestamp 1676381911
transform 1 0 12768 0 -1 43848
box -48 -56 432 834
use sg13g2_buf_1  fanout718
timestamp 1676381911
transform -1 0 12768 0 -1 45360
box -48 -56 432 834
use sg13g2_buf_1  fanout719
timestamp 1676381911
transform 1 0 12192 0 -1 55944
box -48 -56 432 834
use sg13g2_buf_1  fanout720
timestamp 1676381911
transform -1 0 6432 0 -1 86184
box -48 -56 432 834
use sg13g2_buf_1  fanout721
timestamp 1676381911
transform 1 0 12384 0 1 86184
box -48 -56 432 834
use sg13g2_buf_1  fanout722
timestamp 1676381911
transform 1 0 8832 0 -1 84672
box -48 -56 432 834
use sg13g2_buf_1  fanout723
timestamp 1676381911
transform 1 0 11616 0 1 63504
box -48 -56 432 834
use sg13g2_buf_1  fanout724
timestamp 1676381911
transform -1 0 6528 0 1 55944
box -48 -56 432 834
use sg13g2_buf_1  fanout725
timestamp 1676381911
transform 1 0 10752 0 -1 16632
box -48 -56 432 834
use sg13g2_buf_1  fanout726
timestamp 1676381911
transform 1 0 12576 0 1 15120
box -48 -56 432 834
use sg13g2_buf_1  fanout727
timestamp 1676381911
transform 1 0 9408 0 -1 24192
box -48 -56 432 834
use sg13g2_buf_1  fanout728
timestamp 1676381911
transform 1 0 8928 0 -1 28728
box -48 -56 432 834
use sg13g2_buf_1  fanout729
timestamp 1676381911
transform -1 0 5664 0 1 25704
box -48 -56 432 834
use sg13g2_buf_1  fanout730
timestamp 1676381911
transform 1 0 8640 0 1 24192
box -48 -56 432 834
use sg13g2_buf_1  fanout731
timestamp 1676381911
transform 1 0 7872 0 -1 48384
box -48 -56 432 834
use sg13g2_buf_1  fanout732
timestamp 1676381911
transform 1 0 7776 0 1 74088
box -48 -56 432 834
use sg13g2_buf_1  fanout733
timestamp 1676381911
transform 1 0 10272 0 1 80136
box -48 -56 432 834
use sg13g2_buf_1  fanout734
timestamp 1676381911
transform -1 0 5664 0 1 83160
box -48 -56 432 834
use sg13g2_buf_1  fanout735
timestamp 1676381911
transform 1 0 10656 0 -1 81648
box -48 -56 432 834
use sg13g2_buf_1  fanout736
timestamp 1676381911
transform -1 0 8160 0 1 58968
box -48 -56 432 834
use sg13g2_buf_1  fanout737
timestamp 1676381911
transform 1 0 7008 0 1 57456
box -48 -56 432 834
use sg13g2_buf_1  fanout738
timestamp 1676381911
transform 1 0 10272 0 -1 48384
box -48 -56 432 834
use sg13g2_buf_1  fanout739
timestamp 1676381911
transform -1 0 11040 0 -1 48384
box -48 -56 432 834
use sg13g2_buf_1  fanout740
timestamp 1676381911
transform 1 0 8640 0 -1 37800
box -48 -56 432 834
use sg13g2_buf_1  fanout741
timestamp 1676381911
transform -1 0 8928 0 1 37800
box -48 -56 432 834
use sg13g2_buf_1  fanout742
timestamp 1676381911
transform -1 0 9408 0 -1 48384
box -48 -56 432 834
use sg13g2_buf_1  fanout743
timestamp 1676381911
transform 1 0 11616 0 1 49896
box -48 -56 432 834
use sg13g2_buf_1  fanout744
timestamp 1676381911
transform 1 0 15936 0 1 66528
box -48 -56 432 834
use sg13g2_buf_1  fanout745
timestamp 1676381911
transform -1 0 15744 0 1 57456
box -48 -56 432 834
use sg13g2_buf_1  fanout746
timestamp 1676381911
transform -1 0 12576 0 -1 74088
box -48 -56 432 834
use sg13g2_buf_1  fanout747
timestamp 1676381911
transform 1 0 11712 0 -1 58968
box -48 -56 432 834
use sg13g2_buf_1  fanout748
timestamp 1676381911
transform 1 0 11520 0 -1 49896
box -48 -56 432 834
use sg13g2_buf_1  fanout749
timestamp 1676381911
transform -1 0 9792 0 1 48384
box -48 -56 432 834
use sg13g2_buf_1  fanout750
timestamp 1676381911
transform 1 0 5280 0 -1 24192
box -48 -56 432 834
use sg13g2_buf_1  fanout751
timestamp 1676381911
transform -1 0 4704 0 1 21168
box -48 -56 432 834
use sg13g2_buf_1  fanout752
timestamp 1676381911
transform 1 0 3840 0 1 22680
box -48 -56 432 834
use sg13g2_buf_1  fanout753
timestamp 1676381911
transform -1 0 5664 0 1 24192
box -48 -56 432 834
use sg13g2_buf_1  fanout754
timestamp 1676381911
transform 1 0 4896 0 -1 25704
box -48 -56 432 834
use sg13g2_buf_1  fanout755
timestamp 1676381911
transform -1 0 4704 0 -1 25704
box -48 -56 432 834
use sg13g2_buf_1  fanout756
timestamp 1676381911
transform -1 0 17664 0 1 45360
box -48 -56 432 834
use sg13g2_buf_1  fanout757
timestamp 1676381911
transform 1 0 9120 0 1 31752
box -48 -56 432 834
use sg13g2_buf_1  fanout758
timestamp 1676381911
transform -1 0 8256 0 1 31752
box -48 -56 432 834
use sg13g2_buf_1  fanout759
timestamp 1676381911
transform -1 0 15840 0 -1 45360
box -48 -56 432 834
use sg13g2_buf_1  fanout760
timestamp 1676381911
transform 1 0 7200 0 -1 33264
box -48 -56 432 834
use sg13g2_buf_1  fanout761
timestamp 1676381911
transform 1 0 6528 0 1 31752
box -48 -56 432 834
use sg13g2_buf_1  fanout762
timestamp 1676381911
transform -1 0 11904 0 1 43848
box -48 -56 432 834
use sg13g2_buf_1  fanout763
timestamp 1676381911
transform -1 0 11520 0 1 43848
box -48 -56 432 834
use sg13g2_buf_1  fanout764
timestamp 1676381911
transform -1 0 6816 0 -1 36288
box -48 -56 432 834
use sg13g2_buf_1  fanout765
timestamp 1676381911
transform -1 0 5952 0 -1 34776
box -48 -56 432 834
use sg13g2_buf_1  fanout766
timestamp 1676381911
transform 1 0 9312 0 -1 40824
box -48 -56 432 834
use sg13g2_buf_1  fanout767
timestamp 1676381911
transform 1 0 10752 0 1 39312
box -48 -56 432 834
use sg13g2_buf_1  fanout768
timestamp 1676381911
transform 1 0 11616 0 1 25704
box -48 -56 432 834
use sg13g2_buf_1  fanout769
timestamp 1676381911
transform 1 0 12960 0 -1 27216
box -48 -56 432 834
use sg13g2_buf_1  fanout770
timestamp 1676381911
transform 1 0 9312 0 1 28728
box -48 -56 432 834
use sg13g2_buf_1  fanout771
timestamp 1676381911
transform -1 0 18528 0 1 43848
box -48 -56 432 834
use sg13g2_buf_1  fanout772
timestamp 1676381911
transform 1 0 15840 0 -1 43848
box -48 -56 432 834
use sg13g2_buf_1  fanout773
timestamp 1676381911
transform -1 0 18240 0 -1 37800
box -48 -56 432 834
use sg13g2_buf_1  fanout774
timestamp 1676381911
transform -1 0 16608 0 1 37800
box -48 -56 432 834
use sg13g2_buf_1  fanout775
timestamp 1676381911
transform -1 0 14400 0 1 25704
box -48 -56 432 834
use sg13g2_buf_1  fanout776
timestamp 1676381911
transform -1 0 10944 0 -1 27216
box -48 -56 432 834
use sg13g2_buf_1  fanout777
timestamp 1676381911
transform 1 0 8544 0 -1 30240
box -48 -56 432 834
use sg13g2_buf_1  fanout778
timestamp 1676381911
transform -1 0 12480 0 1 31752
box -48 -56 432 834
use sg13g2_buf_1  fanout779
timestamp 1676381911
transform 1 0 8544 0 -1 40824
box -48 -56 432 834
use sg13g2_buf_1  fanout780
timestamp 1676381911
transform -1 0 9792 0 1 37800
box -48 -56 432 834
use sg13g2_buf_1  fanout781
timestamp 1676381911
transform -1 0 18048 0 -1 33264
box -48 -56 432 834
use sg13g2_buf_1  fanout782
timestamp 1676381911
transform 1 0 14304 0 -1 68040
box -48 -56 432 834
use sg13g2_buf_1  fanout783
timestamp 1676381911
transform 1 0 10368 0 -1 69552
box -48 -56 432 834
use sg13g2_buf_1  fanout784
timestamp 1676381911
transform -1 0 9312 0 1 69552
box -48 -56 432 834
use sg13g2_buf_1  fanout785
timestamp 1676381911
transform -1 0 4608 0 -1 75600
box -48 -56 432 834
use sg13g2_buf_1  fanout786
timestamp 1676381911
transform -1 0 8544 0 1 81648
box -48 -56 432 834
use sg13g2_buf_1  fanout787
timestamp 1676381911
transform -1 0 4704 0 -1 87696
box -48 -56 432 834
use sg13g2_buf_1  fanout788
timestamp 1676381911
transform 1 0 10656 0 -1 87696
box -48 -56 432 834
use sg13g2_buf_1  fanout789
timestamp 1676381911
transform -1 0 4320 0 -1 81648
box -48 -56 432 834
use sg13g2_buf_1  fanout790
timestamp 1676381911
transform 1 0 4320 0 -1 81648
box -48 -56 432 834
use sg13g2_buf_1  fanout791
timestamp 1676381911
transform -1 0 10752 0 -1 89208
box -48 -56 432 834
use sg13g2_buf_1  fanout792
timestamp 1676381911
transform 1 0 6912 0 1 86184
box -48 -56 432 834
use sg13g2_buf_1  fanout793
timestamp 1676381911
transform 1 0 9312 0 1 86184
box -48 -56 432 834
use sg13g2_buf_1  fanout794
timestamp 1676381911
transform 1 0 13344 0 1 81648
box -48 -56 432 834
use sg13g2_buf_1  fanout795
timestamp 1676381911
transform 1 0 12384 0 1 80136
box -48 -56 432 834
use sg13g2_buf_1  fanout796
timestamp 1676381911
transform -1 0 10848 0 1 78624
box -48 -56 432 834
use sg13g2_buf_1  fanout797
timestamp 1676381911
transform 1 0 14016 0 -1 78624
box -48 -56 432 834
use sg13g2_buf_1  fanout798
timestamp 1676381911
transform -1 0 9888 0 1 78624
box -48 -56 432 834
use sg13g2_buf_1  fanout799
timestamp 1676381911
transform -1 0 10080 0 -1 72576
box -48 -56 432 834
use sg13g2_buf_1  fanout800
timestamp 1676381911
transform -1 0 3552 0 -1 87696
box -48 -56 432 834
use sg13g2_buf_1  fanout801
timestamp 1676381911
transform 1 0 3552 0 -1 87696
box -48 -56 432 834
use sg13g2_buf_1  fanout802
timestamp 1676381911
transform -1 0 16128 0 -1 77112
box -48 -56 432 834
use sg13g2_buf_1  fanout803
timestamp 1676381911
transform 1 0 18048 0 1 75600
box -48 -56 432 834
use sg13g2_buf_1  fanout804
timestamp 1676381911
transform 1 0 17088 0 -1 78624
box -48 -56 432 834
use sg13g2_buf_1  fanout805
timestamp 1676381911
transform 1 0 12192 0 -1 65016
box -48 -56 432 834
use sg13g2_buf_1  fanout806
timestamp 1676381911
transform 1 0 12096 0 -1 63504
box -48 -56 432 834
use sg13g2_buf_1  fanout807
timestamp 1676381911
transform 1 0 6912 0 -1 66528
box -48 -56 432 834
use sg13g2_buf_1  fanout808
timestamp 1676381911
transform 1 0 2208 0 1 71064
box -48 -56 432 834
use sg13g2_buf_1  fanout809
timestamp 1676381911
transform 1 0 6048 0 -1 89208
box -48 -56 432 834
use sg13g2_buf_1  fanout810
timestamp 1676381911
transform 1 0 3072 0 1 89208
box -48 -56 432 834
use sg13g2_buf_1  fanout811
timestamp 1676381911
transform -1 0 17376 0 -1 86184
box -48 -56 432 834
use sg13g2_buf_1  fanout812
timestamp 1676381911
transform 1 0 14496 0 1 83160
box -48 -56 432 834
use sg13g2_buf_1  fanout813
timestamp 1676381911
transform 1 0 15360 0 -1 77112
box -48 -56 432 834
use sg13g2_fill_1  FILLER_0_0
timestamp 1677579658
transform 1 0 1152 0 1 1512
box -48 -56 144 834
use sg13g2_decap_4  FILLER_0_69
timestamp 1679577901
transform 1 0 7776 0 1 1512
box -48 -56 432 834
use sg13g2_decap_8  FILLER_0_161
timestamp 1679581782
transform 1 0 16608 0 1 1512
box -48 -56 720 834
use sg13g2_fill_1  FILLER_0_168
timestamp 1677579658
transform 1 0 17280 0 1 1512
box -48 -56 144 834
use sg13g2_decap_8  FILLER_0_173
timestamp 1679581782
transform 1 0 17760 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_180
timestamp 1679581782
transform 1 0 18432 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_187
timestamp 1679581782
transform 1 0 19104 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_194
timestamp 1679581782
transform 1 0 19776 0 1 1512
box -48 -56 720 834
use sg13g2_fill_1  FILLER_1_4
timestamp 1677579658
transform 1 0 1536 0 -1 3024
box -48 -56 144 834
use sg13g2_fill_1  FILLER_1_13
timestamp 1677579658
transform 1 0 2400 0 -1 3024
box -48 -56 144 834
use sg13g2_fill_2  FILLER_1_18
timestamp 1677580104
transform 1 0 2880 0 -1 3024
box -48 -56 240 834
use sg13g2_fill_1  FILLER_1_20
timestamp 1677579658
transform 1 0 3072 0 -1 3024
box -48 -56 144 834
use sg13g2_decap_8  FILLER_1_53
timestamp 1679581782
transform 1 0 6240 0 -1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_60
timestamp 1679581782
transform 1 0 6912 0 -1 3024
box -48 -56 720 834
use sg13g2_decap_4  FILLER_1_67
timestamp 1679577901
transform 1 0 7584 0 -1 3024
box -48 -56 432 834
use sg13g2_fill_2  FILLER_1_71
timestamp 1677580104
transform 1 0 7968 0 -1 3024
box -48 -56 240 834
use sg13g2_decap_4  FILLER_1_77
timestamp 1679577901
transform 1 0 8544 0 -1 3024
box -48 -56 432 834
use sg13g2_decap_8  FILLER_1_105
timestamp 1679581782
transform 1 0 11232 0 -1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_112
timestamp 1679581782
transform 1 0 11904 0 -1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_151
timestamp 1679581782
transform 1 0 15648 0 -1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_158
timestamp 1679581782
transform 1 0 16320 0 -1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_165
timestamp 1679581782
transform 1 0 16992 0 -1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_172
timestamp 1679581782
transform 1 0 17664 0 -1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_179
timestamp 1679581782
transform 1 0 18336 0 -1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_186
timestamp 1679581782
transform 1 0 19008 0 -1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_193
timestamp 1679581782
transform 1 0 19680 0 -1 3024
box -48 -56 720 834
use sg13g2_fill_1  FILLER_1_200
timestamp 1677579658
transform 1 0 20352 0 -1 3024
box -48 -56 144 834
use sg13g2_decap_8  FILLER_2_28
timestamp 1679581782
transform 1 0 3840 0 1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_35
timestamp 1679581782
transform 1 0 4512 0 1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_42
timestamp 1679581782
transform 1 0 5184 0 1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_49
timestamp 1679581782
transform 1 0 5856 0 1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_56
timestamp 1679581782
transform 1 0 6528 0 1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_63
timestamp 1679581782
transform 1 0 7200 0 1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_70
timestamp 1679581782
transform 1 0 7872 0 1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_77
timestamp 1679581782
transform 1 0 8544 0 1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_84
timestamp 1679581782
transform 1 0 9216 0 1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_91
timestamp 1679581782
transform 1 0 9888 0 1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_98
timestamp 1679581782
transform 1 0 10560 0 1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_105
timestamp 1679581782
transform 1 0 11232 0 1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_112
timestamp 1679581782
transform 1 0 11904 0 1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_119
timestamp 1679581782
transform 1 0 12576 0 1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_126
timestamp 1679581782
transform 1 0 13248 0 1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_133
timestamp 1679581782
transform 1 0 13920 0 1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_140
timestamp 1679581782
transform 1 0 14592 0 1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_147
timestamp 1679581782
transform 1 0 15264 0 1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_154
timestamp 1679581782
transform 1 0 15936 0 1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_161
timestamp 1679581782
transform 1 0 16608 0 1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_168
timestamp 1679581782
transform 1 0 17280 0 1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_175
timestamp 1679581782
transform 1 0 17952 0 1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_182
timestamp 1679581782
transform 1 0 18624 0 1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_189
timestamp 1679581782
transform 1 0 19296 0 1 3024
box -48 -56 720 834
use sg13g2_fill_1  FILLER_2_196
timestamp 1677579658
transform 1 0 19968 0 1 3024
box -48 -56 144 834
use sg13g2_decap_8  FILLER_3_20
timestamp 1679581782
transform 1 0 3072 0 -1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_27
timestamp 1679581782
transform 1 0 3744 0 -1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_34
timestamp 1679581782
transform 1 0 4416 0 -1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_41
timestamp 1679581782
transform 1 0 5088 0 -1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_48
timestamp 1679581782
transform 1 0 5760 0 -1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_55
timestamp 1679581782
transform 1 0 6432 0 -1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_62
timestamp 1679581782
transform 1 0 7104 0 -1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_69
timestamp 1679581782
transform 1 0 7776 0 -1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_76
timestamp 1679581782
transform 1 0 8448 0 -1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_83
timestamp 1679581782
transform 1 0 9120 0 -1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_90
timestamp 1679581782
transform 1 0 9792 0 -1 4536
box -48 -56 720 834
use sg13g2_decap_4  FILLER_3_97
timestamp 1679577901
transform 1 0 10464 0 -1 4536
box -48 -56 432 834
use sg13g2_decap_8  FILLER_3_118
timestamp 1679581782
transform 1 0 12480 0 -1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_125
timestamp 1679581782
transform 1 0 13152 0 -1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_132
timestamp 1679581782
transform 1 0 13824 0 -1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_139
timestamp 1679581782
transform 1 0 14496 0 -1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_146
timestamp 1679581782
transform 1 0 15168 0 -1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_153
timestamp 1679581782
transform 1 0 15840 0 -1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_160
timestamp 1679581782
transform 1 0 16512 0 -1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_167
timestamp 1679581782
transform 1 0 17184 0 -1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_174
timestamp 1679581782
transform 1 0 17856 0 -1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_181
timestamp 1679581782
transform 1 0 18528 0 -1 4536
box -48 -56 720 834
use sg13g2_decap_4  FILLER_3_188
timestamp 1679577901
transform 1 0 19200 0 -1 4536
box -48 -56 432 834
use sg13g2_fill_1  FILLER_3_192
timestamp 1677579658
transform 1 0 19584 0 -1 4536
box -48 -56 144 834
use sg13g2_decap_8  FILLER_4_20
timestamp 1679581782
transform 1 0 3072 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_27
timestamp 1679581782
transform 1 0 3744 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_34
timestamp 1679581782
transform 1 0 4416 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_41
timestamp 1679581782
transform 1 0 5088 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_48
timestamp 1679581782
transform 1 0 5760 0 1 4536
box -48 -56 720 834
use sg13g2_fill_1  FILLER_4_55
timestamp 1677579658
transform 1 0 6432 0 1 4536
box -48 -56 144 834
use sg13g2_decap_8  FILLER_4_73
timestamp 1679581782
transform 1 0 8160 0 1 4536
box -48 -56 720 834
use sg13g2_fill_2  FILLER_4_80
timestamp 1677580104
transform 1 0 8832 0 1 4536
box -48 -56 240 834
use sg13g2_decap_4  FILLER_4_128
timestamp 1679577901
transform 1 0 13440 0 1 4536
box -48 -56 432 834
use sg13g2_decap_8  FILLER_4_157
timestamp 1679581782
transform 1 0 16224 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_164
timestamp 1679581782
transform 1 0 16896 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_171
timestamp 1679581782
transform 1 0 17568 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_178
timestamp 1679581782
transform 1 0 18240 0 1 4536
box -48 -56 720 834
use sg13g2_decap_4  FILLER_4_185
timestamp 1679577901
transform 1 0 18912 0 1 4536
box -48 -56 432 834
use sg13g2_decap_8  FILLER_5_24
timestamp 1679581782
transform 1 0 3456 0 -1 6048
box -48 -56 720 834
use sg13g2_fill_1  FILLER_5_31
timestamp 1677579658
transform 1 0 4128 0 -1 6048
box -48 -56 144 834
use sg13g2_fill_2  FILLER_5_40
timestamp 1677580104
transform 1 0 4992 0 -1 6048
box -48 -56 240 834
use sg13g2_fill_2  FILLER_5_97
timestamp 1677580104
transform 1 0 10464 0 -1 6048
box -48 -56 240 834
use sg13g2_fill_1  FILLER_5_99
timestamp 1677579658
transform 1 0 10656 0 -1 6048
box -48 -56 144 834
use sg13g2_decap_8  FILLER_5_176
timestamp 1679581782
transform 1 0 18048 0 -1 6048
box -48 -56 720 834
use sg13g2_fill_2  FILLER_5_183
timestamp 1677580104
transform 1 0 18720 0 -1 6048
box -48 -56 240 834
use sg13g2_fill_1  FILLER_6_16
timestamp 1677579658
transform 1 0 2688 0 1 6048
box -48 -56 144 834
use sg13g2_fill_2  FILLER_6_25
timestamp 1677580104
transform 1 0 3552 0 1 6048
box -48 -56 240 834
use sg13g2_fill_1  FILLER_6_27
timestamp 1677579658
transform 1 0 3744 0 1 6048
box -48 -56 144 834
use sg13g2_decap_8  FILLER_6_45
timestamp 1679581782
transform 1 0 5472 0 1 6048
box -48 -56 720 834
use sg13g2_fill_2  FILLER_6_52
timestamp 1677580104
transform 1 0 6144 0 1 6048
box -48 -56 240 834
use sg13g2_fill_1  FILLER_6_54
timestamp 1677579658
transform 1 0 6336 0 1 6048
box -48 -56 144 834
use sg13g2_fill_2  FILLER_6_72
timestamp 1677580104
transform 1 0 8064 0 1 6048
box -48 -56 240 834
use sg13g2_decap_4  FILLER_6_99
timestamp 1679577901
transform 1 0 10656 0 1 6048
box -48 -56 432 834
use sg13g2_decap_4  FILLER_6_120
timestamp 1679577901
transform 1 0 12672 0 1 6048
box -48 -56 432 834
use sg13g2_fill_1  FILLER_6_124
timestamp 1677579658
transform 1 0 13056 0 1 6048
box -48 -56 144 834
use sg13g2_fill_1  FILLER_6_146
timestamp 1677579658
transform 1 0 15168 0 1 6048
box -48 -56 144 834
use sg13g2_decap_4  FILLER_6_172
timestamp 1679577901
transform 1 0 17664 0 1 6048
box -48 -56 432 834
use sg13g2_fill_2  FILLER_6_176
timestamp 1677580104
transform 1 0 18048 0 1 6048
box -48 -56 240 834
use sg13g2_fill_2  FILLER_6_195
timestamp 1677580104
transform 1 0 19872 0 1 6048
box -48 -56 240 834
use sg13g2_fill_1  FILLER_7_41
timestamp 1677579658
transform 1 0 5088 0 -1 7560
box -48 -56 144 834
use sg13g2_fill_1  FILLER_7_59
timestamp 1677579658
transform 1 0 6816 0 -1 7560
box -48 -56 144 834
use sg13g2_decap_4  FILLER_7_115
timestamp 1679577901
transform 1 0 12192 0 -1 7560
box -48 -56 432 834
use sg13g2_fill_2  FILLER_7_119
timestamp 1677580104
transform 1 0 12576 0 -1 7560
box -48 -56 240 834
use sg13g2_fill_1  FILLER_7_189
timestamp 1677579658
transform 1 0 19296 0 -1 7560
box -48 -56 144 834
use sg13g2_fill_2  FILLER_7_194
timestamp 1677580104
transform 1 0 19776 0 -1 7560
box -48 -56 240 834
use sg13g2_fill_1  FILLER_7_196
timestamp 1677579658
transform 1 0 19968 0 -1 7560
box -48 -56 144 834
use sg13g2_fill_2  FILLER_8_0
timestamp 1677580104
transform 1 0 1152 0 1 7560
box -48 -56 240 834
use sg13g2_fill_1  FILLER_8_36
timestamp 1677579658
transform 1 0 4608 0 1 7560
box -48 -56 144 834
use sg13g2_fill_1  FILLER_8_54
timestamp 1677579658
transform 1 0 6336 0 1 7560
box -48 -56 144 834
use sg13g2_decap_4  FILLER_8_72
timestamp 1679577901
transform 1 0 8064 0 1 7560
box -48 -56 432 834
use sg13g2_fill_1  FILLER_8_76
timestamp 1677579658
transform 1 0 8448 0 1 7560
box -48 -56 144 834
use sg13g2_fill_1  FILLER_8_94
timestamp 1677579658
transform 1 0 10176 0 1 7560
box -48 -56 144 834
use sg13g2_decap_4  FILLER_8_112
timestamp 1679577901
transform 1 0 11904 0 1 7560
box -48 -56 432 834
use sg13g2_fill_2  FILLER_8_150
timestamp 1677580104
transform 1 0 15552 0 1 7560
box -48 -56 240 834
use sg13g2_fill_1  FILLER_8_152
timestamp 1677579658
transform 1 0 15744 0 1 7560
box -48 -56 144 834
use sg13g2_fill_2  FILLER_8_178
timestamp 1677580104
transform 1 0 18240 0 1 7560
box -48 -56 240 834
use sg13g2_fill_2  FILLER_9_25
timestamp 1677580104
transform 1 0 3552 0 -1 9072
box -48 -56 240 834
use sg13g2_fill_2  FILLER_9_94
timestamp 1677580104
transform 1 0 10176 0 -1 9072
box -48 -56 240 834
use sg13g2_fill_1  FILLER_9_113
timestamp 1677579658
transform 1 0 12000 0 -1 9072
box -48 -56 144 834
use sg13g2_decap_8  FILLER_9_135
timestamp 1679581782
transform 1 0 14112 0 -1 9072
box -48 -56 720 834
use sg13g2_fill_1  FILLER_9_146
timestamp 1677579658
transform 1 0 15168 0 -1 9072
box -48 -56 144 834
use sg13g2_fill_2  FILLER_10_4
timestamp 1677580104
transform 1 0 1536 0 1 9072
box -48 -56 240 834
use sg13g2_fill_1  FILLER_10_6
timestamp 1677579658
transform 1 0 1728 0 1 9072
box -48 -56 144 834
use sg13g2_fill_2  FILLER_10_28
timestamp 1677580104
transform 1 0 3840 0 1 9072
box -48 -56 240 834
use sg13g2_fill_2  FILLER_10_55
timestamp 1677580104
transform 1 0 6432 0 1 9072
box -48 -56 240 834
use sg13g2_decap_4  FILLER_10_61
timestamp 1679577901
transform 1 0 7008 0 1 9072
box -48 -56 432 834
use sg13g2_fill_1  FILLER_10_65
timestamp 1677579658
transform 1 0 7392 0 1 9072
box -48 -56 144 834
use sg13g2_decap_8  FILLER_10_108
timestamp 1679581782
transform 1 0 11520 0 1 9072
box -48 -56 720 834
use sg13g2_fill_1  FILLER_10_115
timestamp 1677579658
transform 1 0 12192 0 1 9072
box -48 -56 144 834
use sg13g2_fill_2  FILLER_10_141
timestamp 1677580104
transform 1 0 14688 0 1 9072
box -48 -56 240 834
use sg13g2_fill_1  FILLER_10_143
timestamp 1677579658
transform 1 0 14880 0 1 9072
box -48 -56 144 834
use sg13g2_fill_2  FILLER_10_194
timestamp 1677580104
transform 1 0 19776 0 1 9072
box -48 -56 240 834
use sg13g2_fill_1  FILLER_10_196
timestamp 1677579658
transform 1 0 19968 0 1 9072
box -48 -56 144 834
use sg13g2_fill_2  FILLER_11_4
timestamp 1677580104
transform 1 0 1536 0 -1 10584
box -48 -56 240 834
use sg13g2_fill_1  FILLER_11_6
timestamp 1677579658
transform 1 0 1728 0 -1 10584
box -48 -56 144 834
use sg13g2_fill_1  FILLER_11_15
timestamp 1677579658
transform 1 0 2592 0 -1 10584
box -48 -56 144 834
use sg13g2_fill_1  FILLER_11_54
timestamp 1677579658
transform 1 0 6336 0 -1 10584
box -48 -56 144 834
use sg13g2_decap_8  FILLER_11_76
timestamp 1679581782
transform 1 0 8448 0 -1 10584
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_83
timestamp 1679581782
transform 1 0 9120 0 -1 10584
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_90
timestamp 1679581782
transform 1 0 9792 0 -1 10584
box -48 -56 720 834
use sg13g2_fill_2  FILLER_11_97
timestamp 1677580104
transform 1 0 10464 0 -1 10584
box -48 -56 240 834
use sg13g2_fill_2  FILLER_11_154
timestamp 1677580104
transform 1 0 15936 0 -1 10584
box -48 -56 240 834
use sg13g2_fill_1  FILLER_11_173
timestamp 1677579658
transform 1 0 17760 0 -1 10584
box -48 -56 144 834
use sg13g2_fill_2  FILLER_11_195
timestamp 1677580104
transform 1 0 19872 0 -1 10584
box -48 -56 240 834
use sg13g2_fill_1  FILLER_12_88
timestamp 1677579658
transform 1 0 9600 0 1 10584
box -48 -56 144 834
use sg13g2_fill_2  FILLER_12_127
timestamp 1677580104
transform 1 0 13344 0 1 10584
box -48 -56 240 834
use sg13g2_fill_1  FILLER_12_146
timestamp 1677579658
transform 1 0 15168 0 1 10584
box -48 -56 144 834
use sg13g2_fill_2  FILLER_12_172
timestamp 1677580104
transform 1 0 17664 0 1 10584
box -48 -56 240 834
use sg13g2_fill_2  FILLER_12_191
timestamp 1677580104
transform 1 0 19488 0 1 10584
box -48 -56 240 834
use sg13g2_fill_2  FILLER_13_8
timestamp 1677580104
transform 1 0 1920 0 -1 12096
box -48 -56 240 834
use sg13g2_fill_1  FILLER_13_31
timestamp 1677579658
transform 1 0 4128 0 -1 12096
box -48 -56 144 834
use sg13g2_fill_2  FILLER_13_57
timestamp 1677580104
transform 1 0 6624 0 -1 12096
box -48 -56 240 834
use sg13g2_fill_1  FILLER_13_59
timestamp 1677579658
transform 1 0 6816 0 -1 12096
box -48 -56 144 834
use sg13g2_decap_8  FILLER_13_102
timestamp 1679581782
transform 1 0 10944 0 -1 12096
box -48 -56 720 834
use sg13g2_decap_4  FILLER_13_151
timestamp 1679577901
transform 1 0 15648 0 -1 12096
box -48 -56 432 834
use sg13g2_fill_1  FILLER_14_37
timestamp 1677579658
transform 1 0 4704 0 1 12096
box -48 -56 144 834
use sg13g2_fill_2  FILLER_14_71
timestamp 1677580104
transform 1 0 7968 0 1 12096
box -48 -56 240 834
use sg13g2_decap_8  FILLER_14_94
timestamp 1679581782
transform 1 0 10176 0 1 12096
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_101
timestamp 1679581782
transform 1 0 10848 0 1 12096
box -48 -56 720 834
use sg13g2_fill_2  FILLER_14_108
timestamp 1677580104
transform 1 0 11520 0 1 12096
box -48 -56 240 834
use sg13g2_fill_2  FILLER_14_194
timestamp 1677580104
transform 1 0 19776 0 1 12096
box -48 -56 240 834
use sg13g2_fill_1  FILLER_14_196
timestamp 1677579658
transform 1 0 19968 0 1 12096
box -48 -56 144 834
use sg13g2_fill_1  FILLER_15_29
timestamp 1677579658
transform 1 0 3936 0 -1 13608
box -48 -56 144 834
use sg13g2_fill_1  FILLER_15_47
timestamp 1677579658
transform 1 0 5664 0 -1 13608
box -48 -56 144 834
use sg13g2_fill_2  FILLER_15_65
timestamp 1677580104
transform 1 0 7392 0 -1 13608
box -48 -56 240 834
use sg13g2_fill_1  FILLER_15_67
timestamp 1677579658
transform 1 0 7584 0 -1 13608
box -48 -56 144 834
use sg13g2_decap_8  FILLER_15_80
timestamp 1679581782
transform 1 0 8832 0 -1 13608
box -48 -56 720 834
use sg13g2_fill_1  FILLER_15_121
timestamp 1677579658
transform 1 0 12768 0 -1 13608
box -48 -56 144 834
use sg13g2_decap_8  FILLER_15_139
timestamp 1679581782
transform 1 0 14496 0 -1 13608
box -48 -56 720 834
use sg13g2_fill_2  FILLER_15_146
timestamp 1677580104
transform 1 0 15168 0 -1 13608
box -48 -56 240 834
use sg13g2_fill_1  FILLER_15_148
timestamp 1677579658
transform 1 0 15360 0 -1 13608
box -48 -56 144 834
use sg13g2_fill_1  FILLER_15_174
timestamp 1677579658
transform 1 0 17856 0 -1 13608
box -48 -56 144 834
use sg13g2_fill_1  FILLER_15_196
timestamp 1677579658
transform 1 0 19968 0 -1 13608
box -48 -56 144 834
use sg13g2_fill_1  FILLER_16_12
timestamp 1677579658
transform 1 0 2304 0 1 13608
box -48 -56 144 834
use sg13g2_fill_2  FILLER_16_42
timestamp 1677580104
transform 1 0 5184 0 1 13608
box -48 -56 240 834
use sg13g2_fill_2  FILLER_16_90
timestamp 1677580104
transform 1 0 9792 0 1 13608
box -48 -56 240 834
use sg13g2_fill_1  FILLER_16_96
timestamp 1677579658
transform 1 0 10368 0 1 13608
box -48 -56 144 834
use sg13g2_decap_4  FILLER_16_118
timestamp 1679577901
transform 1 0 12480 0 1 13608
box -48 -56 432 834
use sg13g2_fill_1  FILLER_16_122
timestamp 1677579658
transform 1 0 12864 0 1 13608
box -48 -56 144 834
use sg13g2_fill_1  FILLER_16_182
timestamp 1677579658
transform 1 0 18624 0 1 13608
box -48 -56 144 834
use sg13g2_fill_1  FILLER_16_200
timestamp 1677579658
transform 1 0 20352 0 1 13608
box -48 -56 144 834
use sg13g2_fill_2  FILLER_17_0
timestamp 1677580104
transform 1 0 1152 0 -1 15120
box -48 -56 240 834
use sg13g2_fill_2  FILLER_17_95
timestamp 1677580104
transform 1 0 10272 0 -1 15120
box -48 -56 240 834
use sg13g2_fill_1  FILLER_17_97
timestamp 1677579658
transform 1 0 10464 0 -1 15120
box -48 -56 144 834
use sg13g2_fill_1  FILLER_17_119
timestamp 1677579658
transform 1 0 12576 0 -1 15120
box -48 -56 144 834
use sg13g2_decap_4  FILLER_17_141
timestamp 1679577901
transform 1 0 14688 0 -1 15120
box -48 -56 432 834
use sg13g2_fill_2  FILLER_17_145
timestamp 1677580104
transform 1 0 15072 0 -1 15120
box -48 -56 240 834
use sg13g2_fill_2  FILLER_17_176
timestamp 1677580104
transform 1 0 18048 0 -1 15120
box -48 -56 240 834
use sg13g2_fill_2  FILLER_17_199
timestamp 1677580104
transform 1 0 20256 0 -1 15120
box -48 -56 240 834
use sg13g2_fill_1  FILLER_18_0
timestamp 1677579658
transform 1 0 1152 0 1 15120
box -48 -56 144 834
use sg13g2_fill_1  FILLER_18_18
timestamp 1677579658
transform 1 0 2880 0 1 15120
box -48 -56 144 834
use sg13g2_fill_1  FILLER_18_61
timestamp 1677579658
transform 1 0 7008 0 1 15120
box -48 -56 144 834
use sg13g2_fill_1  FILLER_18_66
timestamp 1677579658
transform 1 0 7488 0 1 15120
box -48 -56 144 834
use sg13g2_fill_1  FILLER_18_101
timestamp 1677579658
transform 1 0 10848 0 1 15120
box -48 -56 144 834
use sg13g2_fill_1  FILLER_18_123
timestamp 1677579658
transform 1 0 12960 0 1 15120
box -48 -56 144 834
use sg13g2_fill_2  FILLER_18_141
timestamp 1677580104
transform 1 0 14688 0 1 15120
box -48 -56 240 834
use sg13g2_fill_1  FILLER_18_143
timestamp 1677579658
transform 1 0 14880 0 1 15120
box -48 -56 144 834
use sg13g2_fill_2  FILLER_18_199
timestamp 1677580104
transform 1 0 20256 0 1 15120
box -48 -56 240 834
use sg13g2_fill_1  FILLER_19_4
timestamp 1677579658
transform 1 0 1536 0 -1 16632
box -48 -56 144 834
use sg13g2_fill_2  FILLER_19_22
timestamp 1677580104
transform 1 0 3264 0 -1 16632
box -48 -56 240 834
use sg13g2_fill_1  FILLER_19_24
timestamp 1677579658
transform 1 0 3456 0 -1 16632
box -48 -56 144 834
use sg13g2_fill_1  FILLER_19_58
timestamp 1677579658
transform 1 0 6720 0 -1 16632
box -48 -56 144 834
use sg13g2_fill_2  FILLER_19_63
timestamp 1677580104
transform 1 0 7200 0 -1 16632
box -48 -56 240 834
use sg13g2_fill_1  FILLER_19_82
timestamp 1677579658
transform 1 0 9024 0 -1 16632
box -48 -56 144 834
use sg13g2_decap_4  FILLER_19_121
timestamp 1679577901
transform 1 0 12768 0 -1 16632
box -48 -56 432 834
use sg13g2_fill_2  FILLER_19_163
timestamp 1677580104
transform 1 0 16800 0 -1 16632
box -48 -56 240 834
use sg13g2_fill_1  FILLER_19_165
timestamp 1677579658
transform 1 0 16992 0 -1 16632
box -48 -56 144 834
use sg13g2_fill_2  FILLER_19_199
timestamp 1677580104
transform 1 0 20256 0 -1 16632
box -48 -56 240 834
use sg13g2_fill_1  FILLER_20_17
timestamp 1677579658
transform 1 0 2784 0 1 16632
box -48 -56 144 834
use sg13g2_fill_1  FILLER_20_39
timestamp 1677579658
transform 1 0 4896 0 1 16632
box -48 -56 144 834
use sg13g2_fill_2  FILLER_20_78
timestamp 1677580104
transform 1 0 8640 0 1 16632
box -48 -56 240 834
use sg13g2_fill_2  FILLER_20_105
timestamp 1677580104
transform 1 0 11232 0 1 16632
box -48 -56 240 834
use sg13g2_decap_4  FILLER_20_124
timestamp 1679577901
transform 1 0 13056 0 1 16632
box -48 -56 432 834
use sg13g2_fill_2  FILLER_20_166
timestamp 1677580104
transform 1 0 17088 0 1 16632
box -48 -56 240 834
use sg13g2_fill_1  FILLER_21_21
timestamp 1677579658
transform 1 0 3168 0 -1 18144
box -48 -56 144 834
use sg13g2_fill_2  FILLER_21_55
timestamp 1677580104
transform 1 0 6432 0 -1 18144
box -48 -56 240 834
use sg13g2_fill_1  FILLER_21_95
timestamp 1677579658
transform 1 0 10272 0 -1 18144
box -48 -56 144 834
use sg13g2_decap_8  FILLER_21_100
timestamp 1679581782
transform 1 0 10752 0 -1 18144
box -48 -56 720 834
use sg13g2_decap_4  FILLER_21_107
timestamp 1679577901
transform 1 0 11424 0 -1 18144
box -48 -56 432 834
use sg13g2_decap_8  FILLER_21_128
timestamp 1679581782
transform 1 0 13440 0 -1 18144
box -48 -56 720 834
use sg13g2_fill_1  FILLER_21_139
timestamp 1677579658
transform 1 0 14496 0 -1 18144
box -48 -56 144 834
use sg13g2_fill_2  FILLER_21_194
timestamp 1677580104
transform 1 0 19776 0 -1 18144
box -48 -56 240 834
use sg13g2_fill_1  FILLER_21_196
timestamp 1677579658
transform 1 0 19968 0 -1 18144
box -48 -56 144 834
use sg13g2_fill_2  FILLER_22_45
timestamp 1677580104
transform 1 0 5472 0 1 18144
box -48 -56 240 834
use sg13g2_fill_1  FILLER_22_64
timestamp 1677579658
transform 1 0 7296 0 1 18144
box -48 -56 144 834
use sg13g2_decap_8  FILLER_22_90
timestamp 1679581782
transform 1 0 9792 0 1 18144
box -48 -56 720 834
use sg13g2_fill_2  FILLER_22_97
timestamp 1677580104
transform 1 0 10464 0 1 18144
box -48 -56 240 834
use sg13g2_fill_1  FILLER_22_171
timestamp 1677579658
transform 1 0 17568 0 1 18144
box -48 -56 144 834
use sg13g2_fill_1  FILLER_23_0
timestamp 1677579658
transform 1 0 1152 0 -1 19656
box -48 -56 144 834
use sg13g2_fill_2  FILLER_23_43
timestamp 1677580104
transform 1 0 5280 0 -1 19656
box -48 -56 240 834
use sg13g2_fill_2  FILLER_23_98
timestamp 1677580104
transform 1 0 10560 0 -1 19656
box -48 -56 240 834
use sg13g2_decap_8  FILLER_23_117
timestamp 1679581782
transform 1 0 12384 0 -1 19656
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_124
timestamp 1679581782
transform 1 0 13056 0 -1 19656
box -48 -56 720 834
use sg13g2_fill_2  FILLER_23_131
timestamp 1677580104
transform 1 0 13728 0 -1 19656
box -48 -56 240 834
use sg13g2_fill_1  FILLER_23_143
timestamp 1677579658
transform 1 0 14880 0 -1 19656
box -48 -56 144 834
use sg13g2_fill_2  FILLER_23_149
timestamp 1677580104
transform 1 0 15456 0 -1 19656
box -48 -56 240 834
use sg13g2_fill_2  FILLER_23_176
timestamp 1677580104
transform 1 0 18048 0 -1 19656
box -48 -56 240 834
use sg13g2_fill_2  FILLER_23_199
timestamp 1677580104
transform 1 0 20256 0 -1 19656
box -48 -56 240 834
use sg13g2_fill_2  FILLER_24_21
timestamp 1677580104
transform 1 0 3168 0 1 19656
box -48 -56 240 834
use sg13g2_fill_1  FILLER_24_23
timestamp 1677579658
transform 1 0 3360 0 1 19656
box -48 -56 144 834
use sg13g2_fill_1  FILLER_24_62
timestamp 1677579658
transform 1 0 7104 0 1 19656
box -48 -56 144 834
use sg13g2_fill_2  FILLER_24_126
timestamp 1677580104
transform 1 0 13248 0 1 19656
box -48 -56 240 834
use sg13g2_fill_1  FILLER_24_155
timestamp 1677579658
transform 1 0 16032 0 1 19656
box -48 -56 144 834
use sg13g2_fill_2  FILLER_25_25
timestamp 1677580104
transform 1 0 3552 0 -1 21168
box -48 -56 240 834
use sg13g2_fill_1  FILLER_25_27
timestamp 1677579658
transform 1 0 3744 0 -1 21168
box -48 -56 144 834
use sg13g2_fill_1  FILLER_25_45
timestamp 1677579658
transform 1 0 5472 0 -1 21168
box -48 -56 144 834
use sg13g2_decap_4  FILLER_25_109
timestamp 1679577901
transform 1 0 11616 0 -1 21168
box -48 -56 432 834
use sg13g2_fill_2  FILLER_25_178
timestamp 1677580104
transform 1 0 18240 0 -1 21168
box -48 -56 240 834
use sg13g2_fill_2  FILLER_26_37
timestamp 1677580104
transform 1 0 4704 0 1 21168
box -48 -56 240 834
use sg13g2_fill_2  FILLER_26_61
timestamp 1677580104
transform 1 0 7008 0 1 21168
box -48 -56 240 834
use sg13g2_fill_1  FILLER_26_63
timestamp 1677579658
transform 1 0 7200 0 1 21168
box -48 -56 144 834
use sg13g2_fill_2  FILLER_26_115
timestamp 1677580104
transform 1 0 12192 0 1 21168
box -48 -56 240 834
use sg13g2_fill_2  FILLER_26_159
timestamp 1677580104
transform 1 0 16416 0 1 21168
box -48 -56 240 834
use sg13g2_fill_2  FILLER_27_4
timestamp 1677580104
transform 1 0 1536 0 -1 22680
box -48 -56 240 834
use sg13g2_fill_1  FILLER_27_6
timestamp 1677579658
transform 1 0 1728 0 -1 22680
box -48 -56 144 834
use sg13g2_fill_2  FILLER_27_83
timestamp 1677580104
transform 1 0 9120 0 -1 22680
box -48 -56 240 834
use sg13g2_fill_2  FILLER_27_106
timestamp 1677580104
transform 1 0 11328 0 -1 22680
box -48 -56 240 834
use sg13g2_fill_1  FILLER_27_108
timestamp 1677579658
transform 1 0 11520 0 -1 22680
box -48 -56 144 834
use sg13g2_decap_4  FILLER_27_126
timestamp 1679577901
transform 1 0 13248 0 -1 22680
box -48 -56 432 834
use sg13g2_fill_1  FILLER_27_143
timestamp 1677579658
transform 1 0 14880 0 -1 22680
box -48 -56 144 834
use sg13g2_fill_2  FILLER_27_178
timestamp 1677580104
transform 1 0 18240 0 -1 22680
box -48 -56 240 834
use sg13g2_fill_1  FILLER_27_200
timestamp 1677579658
transform 1 0 20352 0 -1 22680
box -48 -56 144 834
use sg13g2_fill_2  FILLER_28_4
timestamp 1677580104
transform 1 0 1536 0 1 22680
box -48 -56 240 834
use sg13g2_fill_1  FILLER_28_6
timestamp 1677579658
transform 1 0 1728 0 1 22680
box -48 -56 144 834
use sg13g2_fill_2  FILLER_28_53
timestamp 1677580104
transform 1 0 6240 0 1 22680
box -48 -56 240 834
use sg13g2_fill_1  FILLER_28_55
timestamp 1677579658
transform 1 0 6432 0 1 22680
box -48 -56 144 834
use sg13g2_fill_2  FILLER_28_106
timestamp 1677580104
transform 1 0 11328 0 1 22680
box -48 -56 240 834
use sg13g2_fill_1  FILLER_28_108
timestamp 1677579658
transform 1 0 11520 0 1 22680
box -48 -56 144 834
use sg13g2_fill_1  FILLER_28_151
timestamp 1677579658
transform 1 0 15648 0 1 22680
box -48 -56 144 834
use sg13g2_fill_1  FILLER_29_0
timestamp 1677579658
transform 1 0 1152 0 -1 24192
box -48 -56 144 834
use sg13g2_fill_2  FILLER_29_47
timestamp 1677580104
transform 1 0 5664 0 -1 24192
box -48 -56 240 834
use sg13g2_fill_1  FILLER_29_49
timestamp 1677579658
transform 1 0 5856 0 -1 24192
box -48 -56 144 834
use sg13g2_fill_2  FILLER_29_67
timestamp 1677580104
transform 1 0 7584 0 -1 24192
box -48 -56 240 834
use sg13g2_fill_2  FILLER_29_94
timestamp 1677580104
transform 1 0 10176 0 -1 24192
box -48 -56 240 834
use sg13g2_fill_1  FILLER_29_96
timestamp 1677579658
transform 1 0 10368 0 -1 24192
box -48 -56 144 834
use sg13g2_fill_1  FILLER_29_131
timestamp 1677579658
transform 1 0 13728 0 -1 24192
box -48 -56 144 834
use sg13g2_fill_2  FILLER_29_157
timestamp 1677580104
transform 1 0 16224 0 -1 24192
box -48 -56 240 834
use sg13g2_fill_2  FILLER_29_179
timestamp 1677580104
transform 1 0 18336 0 -1 24192
box -48 -56 240 834
use sg13g2_fill_1  FILLER_29_200
timestamp 1677579658
transform 1 0 20352 0 -1 24192
box -48 -56 144 834
use sg13g2_fill_1  FILLER_30_0
timestamp 1677579658
transform 1 0 1152 0 1 24192
box -48 -56 144 834
use sg13g2_fill_2  FILLER_30_51
timestamp 1677580104
transform 1 0 6048 0 1 24192
box -48 -56 240 834
use sg13g2_fill_2  FILLER_30_124
timestamp 1677580104
transform 1 0 13056 0 1 24192
box -48 -56 240 834
use sg13g2_fill_2  FILLER_31_4
timestamp 1677580104
transform 1 0 1536 0 -1 25704
box -48 -56 240 834
use sg13g2_fill_1  FILLER_31_6
timestamp 1677579658
transform 1 0 1728 0 -1 25704
box -48 -56 144 834
use sg13g2_fill_1  FILLER_31_32
timestamp 1677579658
transform 1 0 4224 0 -1 25704
box -48 -56 144 834
use sg13g2_fill_2  FILLER_31_37
timestamp 1677580104
transform 1 0 4704 0 -1 25704
box -48 -56 240 834
use sg13g2_fill_2  FILLER_31_64
timestamp 1677580104
transform 1 0 7296 0 -1 25704
box -48 -56 240 834
use sg13g2_fill_1  FILLER_31_66
timestamp 1677579658
transform 1 0 7488 0 -1 25704
box -48 -56 144 834
use sg13g2_fill_1  FILLER_31_105
timestamp 1677579658
transform 1 0 11232 0 -1 25704
box -48 -56 144 834
use sg13g2_decap_4  FILLER_31_123
timestamp 1679577901
transform 1 0 12960 0 -1 25704
box -48 -56 432 834
use sg13g2_fill_2  FILLER_31_127
timestamp 1677580104
transform 1 0 13344 0 -1 25704
box -48 -56 240 834
use sg13g2_fill_2  FILLER_31_133
timestamp 1677580104
transform 1 0 13920 0 -1 25704
box -48 -56 240 834
use sg13g2_fill_2  FILLER_32_0
timestamp 1677580104
transform 1 0 1152 0 1 25704
box -48 -56 240 834
use sg13g2_fill_2  FILLER_32_41
timestamp 1677580104
transform 1 0 5088 0 1 25704
box -48 -56 240 834
use sg13g2_fill_1  FILLER_32_47
timestamp 1677579658
transform 1 0 5664 0 1 25704
box -48 -56 144 834
use sg13g2_fill_2  FILLER_32_107
timestamp 1677580104
transform 1 0 11424 0 1 25704
box -48 -56 240 834
use sg13g2_fill_2  FILLER_32_138
timestamp 1677580104
transform 1 0 14400 0 1 25704
box -48 -56 240 834
use sg13g2_fill_1  FILLER_32_140
timestamp 1677579658
transform 1 0 14592 0 1 25704
box -48 -56 144 834
use sg13g2_fill_1  FILLER_32_200
timestamp 1677579658
transform 1 0 20352 0 1 25704
box -48 -56 144 834
use sg13g2_fill_2  FILLER_33_0
timestamp 1677580104
transform 1 0 1152 0 -1 27216
box -48 -56 240 834
use sg13g2_fill_1  FILLER_33_2
timestamp 1677579658
transform 1 0 1344 0 -1 27216
box -48 -56 144 834
use sg13g2_fill_1  FILLER_33_71
timestamp 1677579658
transform 1 0 7968 0 -1 27216
box -48 -56 144 834
use sg13g2_fill_1  FILLER_33_97
timestamp 1677579658
transform 1 0 10464 0 -1 27216
box -48 -56 144 834
use sg13g2_fill_2  FILLER_33_127
timestamp 1677580104
transform 1 0 13344 0 -1 27216
box -48 -56 240 834
use sg13g2_fill_2  FILLER_33_168
timestamp 1677580104
transform 1 0 17280 0 -1 27216
box -48 -56 240 834
use sg13g2_fill_2  FILLER_33_199
timestamp 1677580104
transform 1 0 20256 0 -1 27216
box -48 -56 240 834
use sg13g2_fill_2  FILLER_34_49
timestamp 1677580104
transform 1 0 5856 0 1 27216
box -48 -56 240 834
use sg13g2_fill_2  FILLER_34_85
timestamp 1677580104
transform 1 0 9312 0 1 27216
box -48 -56 240 834
use sg13g2_fill_2  FILLER_34_121
timestamp 1677580104
transform 1 0 12768 0 1 27216
box -48 -56 240 834
use sg13g2_fill_1  FILLER_34_123
timestamp 1677579658
transform 1 0 12960 0 1 27216
box -48 -56 144 834
use sg13g2_fill_2  FILLER_34_141
timestamp 1677580104
transform 1 0 14688 0 1 27216
box -48 -56 240 834
use sg13g2_fill_1  FILLER_34_143
timestamp 1677579658
transform 1 0 14880 0 1 27216
box -48 -56 144 834
use sg13g2_fill_1  FILLER_34_161
timestamp 1677579658
transform 1 0 16608 0 1 27216
box -48 -56 144 834
use sg13g2_fill_2  FILLER_35_0
timestamp 1677580104
transform 1 0 1152 0 -1 28728
box -48 -56 240 834
use sg13g2_fill_1  FILLER_35_2
timestamp 1677579658
transform 1 0 1344 0 -1 28728
box -48 -56 144 834
use sg13g2_fill_2  FILLER_35_20
timestamp 1677580104
transform 1 0 3072 0 -1 28728
box -48 -56 240 834
use sg13g2_fill_2  FILLER_35_27
timestamp 1677580104
transform 1 0 3744 0 -1 28728
box -48 -56 240 834
use sg13g2_fill_2  FILLER_35_135
timestamp 1677580104
transform 1 0 14112 0 -1 28728
box -48 -56 240 834
use sg13g2_fill_1  FILLER_35_200
timestamp 1677579658
transform 1 0 20352 0 -1 28728
box -48 -56 144 834
use sg13g2_fill_2  FILLER_36_12
timestamp 1677580104
transform 1 0 2304 0 1 28728
box -48 -56 240 834
use sg13g2_fill_2  FILLER_36_55
timestamp 1677580104
transform 1 0 6432 0 1 28728
box -48 -56 240 834
use sg13g2_fill_2  FILLER_36_78
timestamp 1677580104
transform 1 0 8640 0 1 28728
box -48 -56 240 834
use sg13g2_fill_1  FILLER_36_80
timestamp 1677579658
transform 1 0 8832 0 1 28728
box -48 -56 144 834
use sg13g2_fill_2  FILLER_36_110
timestamp 1677580104
transform 1 0 11712 0 1 28728
box -48 -56 240 834
use sg13g2_fill_1  FILLER_36_112
timestamp 1677579658
transform 1 0 11904 0 1 28728
box -48 -56 144 834
use sg13g2_decap_4  FILLER_36_130
timestamp 1679577901
transform 1 0 13632 0 1 28728
box -48 -56 432 834
use sg13g2_fill_1  FILLER_36_134
timestamp 1677579658
transform 1 0 14016 0 1 28728
box -48 -56 144 834
use sg13g2_fill_2  FILLER_36_144
timestamp 1677580104
transform 1 0 14976 0 1 28728
box -48 -56 240 834
use sg13g2_fill_1  FILLER_36_196
timestamp 1677579658
transform 1 0 19968 0 1 28728
box -48 -56 144 834
use sg13g2_fill_2  FILLER_37_0
timestamp 1677580104
transform 1 0 1152 0 -1 30240
box -48 -56 240 834
use sg13g2_fill_2  FILLER_37_85
timestamp 1677580104
transform 1 0 9312 0 -1 30240
box -48 -56 240 834
use sg13g2_fill_2  FILLER_37_112
timestamp 1677580104
transform 1 0 11904 0 -1 30240
box -48 -56 240 834
use sg13g2_fill_1  FILLER_37_114
timestamp 1677579658
transform 1 0 12096 0 -1 30240
box -48 -56 144 834
use sg13g2_decap_4  FILLER_37_119
timestamp 1679577901
transform 1 0 12576 0 -1 30240
box -48 -56 432 834
use sg13g2_fill_2  FILLER_37_163
timestamp 1677580104
transform 1 0 16800 0 -1 30240
box -48 -56 240 834
use sg13g2_fill_2  FILLER_37_191
timestamp 1677580104
transform 1 0 19488 0 -1 30240
box -48 -56 240 834
use sg13g2_fill_1  FILLER_38_122
timestamp 1677579658
transform 1 0 12864 0 1 30240
box -48 -56 144 834
use sg13g2_fill_2  FILLER_38_179
timestamp 1677580104
transform 1 0 18336 0 1 30240
box -48 -56 240 834
use sg13g2_fill_2  FILLER_39_0
timestamp 1677580104
transform 1 0 1152 0 -1 31752
box -48 -56 240 834
use sg13g2_fill_2  FILLER_39_56
timestamp 1677580104
transform 1 0 6528 0 -1 31752
box -48 -56 240 834
use sg13g2_fill_1  FILLER_39_75
timestamp 1677579658
transform 1 0 8352 0 -1 31752
box -48 -56 144 834
use sg13g2_fill_2  FILLER_39_110
timestamp 1677580104
transform 1 0 11712 0 -1 31752
box -48 -56 240 834
use sg13g2_fill_2  FILLER_39_129
timestamp 1677580104
transform 1 0 13536 0 -1 31752
box -48 -56 240 834
use sg13g2_fill_1  FILLER_39_182
timestamp 1677579658
transform 1 0 18624 0 -1 31752
box -48 -56 144 834
use sg13g2_fill_1  FILLER_39_200
timestamp 1677579658
transform 1 0 20352 0 -1 31752
box -48 -56 144 834
use sg13g2_fill_2  FILLER_40_68
timestamp 1677580104
transform 1 0 7680 0 1 31752
box -48 -56 240 834
use sg13g2_fill_1  FILLER_40_82
timestamp 1677579658
transform 1 0 9024 0 1 31752
box -48 -56 144 834
use sg13g2_fill_1  FILLER_40_87
timestamp 1677579658
transform 1 0 9504 0 1 31752
box -48 -56 144 834
use sg13g2_fill_1  FILLER_40_109
timestamp 1677579658
transform 1 0 11616 0 1 31752
box -48 -56 144 834
use sg13g2_decap_8  FILLER_40_118
timestamp 1679581782
transform 1 0 12480 0 1 31752
box -48 -56 720 834
use sg13g2_decap_4  FILLER_40_125
timestamp 1679577901
transform 1 0 13152 0 1 31752
box -48 -56 432 834
use sg13g2_fill_2  FILLER_40_171
timestamp 1677580104
transform 1 0 17568 0 1 31752
box -48 -56 240 834
use sg13g2_fill_1  FILLER_40_173
timestamp 1677579658
transform 1 0 17760 0 1 31752
box -48 -56 144 834
use sg13g2_fill_2  FILLER_40_199
timestamp 1677580104
transform 1 0 20256 0 1 31752
box -48 -56 240 834
use sg13g2_fill_1  FILLER_41_62
timestamp 1677579658
transform 1 0 7104 0 -1 33264
box -48 -56 144 834
use sg13g2_fill_1  FILLER_41_77
timestamp 1677579658
transform 1 0 8544 0 -1 33264
box -48 -56 144 834
use sg13g2_fill_1  FILLER_41_150
timestamp 1677579658
transform 1 0 15552 0 -1 33264
box -48 -56 144 834
use sg13g2_fill_2  FILLER_41_176
timestamp 1677580104
transform 1 0 18048 0 -1 33264
box -48 -56 240 834
use sg13g2_fill_2  FILLER_41_199
timestamp 1677580104
transform 1 0 20256 0 -1 33264
box -48 -56 240 834
use sg13g2_decap_8  FILLER_42_105
timestamp 1679581782
transform 1 0 11232 0 1 33264
box -48 -56 720 834
use sg13g2_decap_4  FILLER_42_112
timestamp 1679577901
transform 1 0 11904 0 1 33264
box -48 -56 432 834
use sg13g2_fill_2  FILLER_42_116
timestamp 1677580104
transform 1 0 12288 0 1 33264
box -48 -56 240 834
use sg13g2_fill_2  FILLER_42_152
timestamp 1677580104
transform 1 0 15744 0 1 33264
box -48 -56 240 834
use sg13g2_fill_1  FILLER_42_154
timestamp 1677579658
transform 1 0 15936 0 1 33264
box -48 -56 144 834
use sg13g2_fill_2  FILLER_42_199
timestamp 1677580104
transform 1 0 20256 0 1 33264
box -48 -56 240 834
use sg13g2_fill_2  FILLER_43_8
timestamp 1677580104
transform 1 0 1920 0 -1 34776
box -48 -56 240 834
use sg13g2_fill_1  FILLER_43_10
timestamp 1677579658
transform 1 0 2112 0 -1 34776
box -48 -56 144 834
use sg13g2_fill_1  FILLER_43_45
timestamp 1677579658
transform 1 0 5472 0 -1 34776
box -48 -56 144 834
use sg13g2_decap_8  FILLER_43_105
timestamp 1679581782
transform 1 0 11232 0 -1 34776
box -48 -56 720 834
use sg13g2_fill_1  FILLER_43_112
timestamp 1677579658
transform 1 0 11904 0 -1 34776
box -48 -56 144 834
use sg13g2_fill_1  FILLER_43_134
timestamp 1677579658
transform 1 0 14016 0 -1 34776
box -48 -56 144 834
use sg13g2_fill_2  FILLER_43_156
timestamp 1677580104
transform 1 0 16128 0 -1 34776
box -48 -56 240 834
use sg13g2_fill_1  FILLER_43_188
timestamp 1677579658
transform 1 0 19200 0 -1 34776
box -48 -56 144 834
use sg13g2_fill_1  FILLER_44_8
timestamp 1677579658
transform 1 0 1920 0 1 34776
box -48 -56 144 834
use sg13g2_fill_2  FILLER_44_26
timestamp 1677580104
transform 1 0 3648 0 1 34776
box -48 -56 240 834
use sg13g2_fill_1  FILLER_44_90
timestamp 1677579658
transform 1 0 9792 0 1 34776
box -48 -56 144 834
use sg13g2_fill_1  FILLER_44_151
timestamp 1677579658
transform 1 0 15648 0 1 34776
box -48 -56 144 834
use sg13g2_fill_1  FILLER_44_200
timestamp 1677579658
transform 1 0 20352 0 1 34776
box -48 -56 144 834
use sg13g2_fill_2  FILLER_45_8
timestamp 1677580104
transform 1 0 1920 0 -1 36288
box -48 -56 240 834
use sg13g2_fill_2  FILLER_45_31
timestamp 1677580104
transform 1 0 4128 0 -1 36288
box -48 -56 240 834
use sg13g2_fill_1  FILLER_45_33
timestamp 1677579658
transform 1 0 4320 0 -1 36288
box -48 -56 144 834
use sg13g2_fill_2  FILLER_45_140
timestamp 1677580104
transform 1 0 14592 0 -1 36288
box -48 -56 240 834
use sg13g2_fill_2  FILLER_46_8
timestamp 1677580104
transform 1 0 1920 0 1 36288
box -48 -56 240 834
use sg13g2_fill_2  FILLER_46_35
timestamp 1677580104
transform 1 0 4512 0 1 36288
box -48 -56 240 834
use sg13g2_fill_1  FILLER_46_37
timestamp 1677579658
transform 1 0 4704 0 1 36288
box -48 -56 144 834
use sg13g2_fill_2  FILLER_46_98
timestamp 1677580104
transform 1 0 10560 0 1 36288
box -48 -56 240 834
use sg13g2_fill_1  FILLER_46_100
timestamp 1677579658
transform 1 0 10752 0 1 36288
box -48 -56 144 834
use sg13g2_fill_2  FILLER_46_146
timestamp 1677580104
transform 1 0 15168 0 1 36288
box -48 -56 240 834
use sg13g2_fill_2  FILLER_46_199
timestamp 1677580104
transform 1 0 20256 0 1 36288
box -48 -56 240 834
use sg13g2_fill_2  FILLER_47_75
timestamp 1677580104
transform 1 0 8352 0 -1 37800
box -48 -56 240 834
use sg13g2_fill_1  FILLER_47_77
timestamp 1677579658
transform 1 0 8544 0 -1 37800
box -48 -56 144 834
use sg13g2_fill_2  FILLER_47_116
timestamp 1677580104
transform 1 0 12288 0 -1 37800
box -48 -56 240 834
use sg13g2_fill_1  FILLER_47_118
timestamp 1677579658
transform 1 0 12480 0 -1 37800
box -48 -56 144 834
use sg13g2_fill_1  FILLER_47_173
timestamp 1677579658
transform 1 0 17760 0 -1 37800
box -48 -56 144 834
use sg13g2_fill_1  FILLER_47_178
timestamp 1677579658
transform 1 0 18240 0 -1 37800
box -48 -56 144 834
use sg13g2_fill_1  FILLER_47_200
timestamp 1677579658
transform 1 0 20352 0 -1 37800
box -48 -56 144 834
use sg13g2_fill_2  FILLER_48_38
timestamp 1677580104
transform 1 0 4800 0 1 37800
box -48 -56 240 834
use sg13g2_decap_8  FILLER_48_65
timestamp 1679581782
transform 1 0 7392 0 1 37800
box -48 -56 720 834
use sg13g2_fill_1  FILLER_48_72
timestamp 1677579658
transform 1 0 8064 0 1 37800
box -48 -56 144 834
use sg13g2_decap_4  FILLER_48_81
timestamp 1679577901
transform 1 0 8928 0 1 37800
box -48 -56 432 834
use sg13g2_fill_1  FILLER_48_85
timestamp 1677579658
transform 1 0 9312 0 1 37800
box -48 -56 144 834
use sg13g2_decap_8  FILLER_48_90
timestamp 1679581782
transform 1 0 9792 0 1 37800
box -48 -56 720 834
use sg13g2_fill_1  FILLER_48_97
timestamp 1677579658
transform 1 0 10464 0 1 37800
box -48 -56 144 834
use sg13g2_fill_2  FILLER_48_123
timestamp 1677580104
transform 1 0 12960 0 1 37800
box -48 -56 240 834
use sg13g2_fill_2  FILLER_48_146
timestamp 1677580104
transform 1 0 15168 0 1 37800
box -48 -56 240 834
use sg13g2_fill_1  FILLER_48_156
timestamp 1677579658
transform 1 0 16128 0 1 37800
box -48 -56 144 834
use sg13g2_fill_1  FILLER_48_161
timestamp 1677579658
transform 1 0 16608 0 1 37800
box -48 -56 144 834
use sg13g2_fill_1  FILLER_48_200
timestamp 1677579658
transform 1 0 20352 0 1 37800
box -48 -56 144 834
use sg13g2_fill_1  FILLER_49_12
timestamp 1677579658
transform 1 0 2304 0 -1 39312
box -48 -56 144 834
use sg13g2_decap_4  FILLER_49_98
timestamp 1679577901
transform 1 0 10560 0 -1 39312
box -48 -56 432 834
use sg13g2_fill_1  FILLER_49_102
timestamp 1677579658
transform 1 0 10944 0 -1 39312
box -48 -56 144 834
use sg13g2_fill_1  FILLER_49_163
timestamp 1677579658
transform 1 0 16800 0 -1 39312
box -48 -56 144 834
use sg13g2_fill_1  FILLER_49_181
timestamp 1677579658
transform 1 0 18528 0 -1 39312
box -48 -56 144 834
use sg13g2_fill_2  FILLER_49_199
timestamp 1677580104
transform 1 0 20256 0 -1 39312
box -48 -56 240 834
use sg13g2_fill_2  FILLER_50_12
timestamp 1677580104
transform 1 0 2304 0 1 39312
box -48 -56 240 834
use sg13g2_fill_2  FILLER_50_64
timestamp 1677580104
transform 1 0 7296 0 1 39312
box -48 -56 240 834
use sg13g2_decap_8  FILLER_50_104
timestamp 1679581782
transform 1 0 11136 0 1 39312
box -48 -56 720 834
use sg13g2_fill_2  FILLER_50_155
timestamp 1677580104
transform 1 0 16032 0 1 39312
box -48 -56 240 834
use sg13g2_fill_2  FILLER_50_174
timestamp 1677580104
transform 1 0 17856 0 1 39312
box -48 -56 240 834
use sg13g2_fill_2  FILLER_51_12
timestamp 1677580104
transform 1 0 2304 0 -1 40824
box -48 -56 240 834
use sg13g2_decap_4  FILLER_51_35
timestamp 1679577901
transform 1 0 4512 0 -1 40824
box -48 -56 432 834
use sg13g2_fill_2  FILLER_51_70
timestamp 1677580104
transform 1 0 7872 0 -1 40824
box -48 -56 240 834
use sg13g2_fill_1  FILLER_51_72
timestamp 1677579658
transform 1 0 8064 0 -1 40824
box -48 -56 144 834
use sg13g2_decap_8  FILLER_51_106
timestamp 1679581782
transform 1 0 11328 0 -1 40824
box -48 -56 720 834
use sg13g2_decap_4  FILLER_51_113
timestamp 1679577901
transform 1 0 12000 0 -1 40824
box -48 -56 432 834
use sg13g2_fill_1  FILLER_51_117
timestamp 1677579658
transform 1 0 12384 0 -1 40824
box -48 -56 144 834
use sg13g2_fill_2  FILLER_51_137
timestamp 1677580104
transform 1 0 14304 0 -1 40824
box -48 -56 240 834
use sg13g2_fill_1  FILLER_51_139
timestamp 1677579658
transform 1 0 14496 0 -1 40824
box -48 -56 144 834
use sg13g2_fill_2  FILLER_51_173
timestamp 1677580104
transform 1 0 17760 0 -1 40824
box -48 -56 240 834
use sg13g2_fill_1  FILLER_51_175
timestamp 1677579658
transform 1 0 17952 0 -1 40824
box -48 -56 144 834
use sg13g2_fill_1  FILLER_52_34
timestamp 1677579658
transform 1 0 4416 0 1 40824
box -48 -56 144 834
use sg13g2_fill_2  FILLER_52_39
timestamp 1677580104
transform 1 0 4896 0 1 40824
box -48 -56 240 834
use sg13g2_fill_2  FILLER_52_63
timestamp 1677580104
transform 1 0 7200 0 1 40824
box -48 -56 240 834
use sg13g2_decap_8  FILLER_52_120
timestamp 1679581782
transform 1 0 12672 0 1 40824
box -48 -56 720 834
use sg13g2_fill_2  FILLER_52_127
timestamp 1677580104
transform 1 0 13344 0 1 40824
box -48 -56 240 834
use sg13g2_fill_1  FILLER_52_129
timestamp 1677579658
transform 1 0 13536 0 1 40824
box -48 -56 144 834
use sg13g2_fill_1  FILLER_52_196
timestamp 1677579658
transform 1 0 19968 0 1 40824
box -48 -56 144 834
use sg13g2_fill_2  FILLER_53_0
timestamp 1677580104
transform 1 0 1152 0 -1 42336
box -48 -56 240 834
use sg13g2_fill_1  FILLER_53_23
timestamp 1677579658
transform 1 0 3360 0 -1 42336
box -48 -56 144 834
use sg13g2_decap_4  FILLER_53_62
timestamp 1679577901
transform 1 0 7104 0 -1 42336
box -48 -56 432 834
use sg13g2_fill_1  FILLER_53_66
timestamp 1677579658
transform 1 0 7488 0 -1 42336
box -48 -56 144 834
use sg13g2_decap_4  FILLER_53_101
timestamp 1679577901
transform 1 0 10848 0 -1 42336
box -48 -56 432 834
use sg13g2_fill_1  FILLER_53_105
timestamp 1677579658
transform 1 0 11232 0 -1 42336
box -48 -56 144 834
use sg13g2_fill_1  FILLER_53_159
timestamp 1677579658
transform 1 0 16416 0 -1 42336
box -48 -56 144 834
use sg13g2_fill_2  FILLER_53_194
timestamp 1677580104
transform 1 0 19776 0 -1 42336
box -48 -56 240 834
use sg13g2_fill_1  FILLER_53_196
timestamp 1677579658
transform 1 0 19968 0 -1 42336
box -48 -56 144 834
use sg13g2_fill_2  FILLER_54_12
timestamp 1677580104
transform 1 0 2304 0 1 42336
box -48 -56 240 834
use sg13g2_decap_4  FILLER_54_83
timestamp 1679577901
transform 1 0 9120 0 1 42336
box -48 -56 432 834
use sg13g2_fill_1  FILLER_54_87
timestamp 1677579658
transform 1 0 9504 0 1 42336
box -48 -56 144 834
use sg13g2_fill_2  FILLER_54_195
timestamp 1677580104
transform 1 0 19872 0 1 42336
box -48 -56 240 834
use sg13g2_fill_1  FILLER_55_8
timestamp 1677579658
transform 1 0 1920 0 -1 43848
box -48 -56 144 834
use sg13g2_fill_2  FILLER_55_30
timestamp 1677580104
transform 1 0 4032 0 -1 43848
box -48 -56 240 834
use sg13g2_fill_1  FILLER_55_32
timestamp 1677579658
transform 1 0 4224 0 -1 43848
box -48 -56 144 834
use sg13g2_fill_1  FILLER_55_53
timestamp 1677579658
transform 1 0 6240 0 -1 43848
box -48 -56 144 834
use sg13g2_decap_4  FILLER_55_75
timestamp 1679577901
transform 1 0 8352 0 -1 43848
box -48 -56 432 834
use sg13g2_fill_1  FILLER_55_79
timestamp 1677579658
transform 1 0 8736 0 -1 43848
box -48 -56 144 834
use sg13g2_fill_2  FILLER_55_97
timestamp 1677580104
transform 1 0 10464 0 -1 43848
box -48 -56 240 834
use sg13g2_fill_1  FILLER_55_99
timestamp 1677579658
transform 1 0 10656 0 -1 43848
box -48 -56 144 834
use sg13g2_decap_4  FILLER_55_129
timestamp 1679577901
transform 1 0 13536 0 -1 43848
box -48 -56 432 834
use sg13g2_fill_2  FILLER_55_133
timestamp 1677580104
transform 1 0 13920 0 -1 43848
box -48 -56 240 834
use sg13g2_fill_2  FILLER_55_195
timestamp 1677580104
transform 1 0 19872 0 -1 43848
box -48 -56 240 834
use sg13g2_fill_2  FILLER_56_8
timestamp 1677580104
transform 1 0 1920 0 1 43848
box -48 -56 240 834
use sg13g2_fill_1  FILLER_56_10
timestamp 1677579658
transform 1 0 2112 0 1 43848
box -48 -56 144 834
use sg13g2_fill_1  FILLER_56_32
timestamp 1677579658
transform 1 0 4224 0 1 43848
box -48 -56 144 834
use sg13g2_fill_2  FILLER_56_93
timestamp 1677580104
transform 1 0 10080 0 1 43848
box -48 -56 240 834
use sg13g2_decap_4  FILLER_56_99
timestamp 1679577901
transform 1 0 10656 0 1 43848
box -48 -56 432 834
use sg13g2_fill_1  FILLER_56_103
timestamp 1677579658
transform 1 0 11040 0 1 43848
box -48 -56 144 834
use sg13g2_fill_1  FILLER_56_181
timestamp 1677579658
transform 1 0 18528 0 1 43848
box -48 -56 144 834
use sg13g2_fill_2  FILLER_56_199
timestamp 1677580104
transform 1 0 20256 0 1 43848
box -48 -56 240 834
use sg13g2_decap_8  FILLER_57_8
timestamp 1679581782
transform 1 0 1920 0 -1 45360
box -48 -56 720 834
use sg13g2_fill_1  FILLER_57_15
timestamp 1677579658
transform 1 0 2592 0 -1 45360
box -48 -56 144 834
use sg13g2_fill_2  FILLER_57_56
timestamp 1677580104
transform 1 0 6528 0 -1 45360
box -48 -56 240 834
use sg13g2_fill_1  FILLER_57_64
timestamp 1677579658
transform 1 0 7296 0 -1 45360
box -48 -56 144 834
use sg13g2_fill_1  FILLER_57_82
timestamp 1677579658
transform 1 0 9024 0 -1 45360
box -48 -56 144 834
use sg13g2_fill_1  FILLER_57_108
timestamp 1677579658
transform 1 0 11520 0 -1 45360
box -48 -56 144 834
use sg13g2_decap_4  FILLER_57_113
timestamp 1679577901
transform 1 0 12000 0 -1 45360
box -48 -56 432 834
use sg13g2_decap_4  FILLER_57_121
timestamp 1679577901
transform 1 0 12768 0 -1 45360
box -48 -56 432 834
use sg13g2_fill_2  FILLER_57_125
timestamp 1677580104
transform 1 0 13152 0 -1 45360
box -48 -56 240 834
use sg13g2_fill_1  FILLER_57_148
timestamp 1677579658
transform 1 0 15360 0 -1 45360
box -48 -56 144 834
use sg13g2_fill_1  FILLER_57_153
timestamp 1677579658
transform 1 0 15840 0 -1 45360
box -48 -56 144 834
use sg13g2_fill_2  FILLER_57_171
timestamp 1677580104
transform 1 0 17568 0 -1 45360
box -48 -56 240 834
use sg13g2_fill_1  FILLER_57_173
timestamp 1677579658
transform 1 0 17760 0 -1 45360
box -48 -56 144 834
use sg13g2_fill_2  FILLER_57_195
timestamp 1677580104
transform 1 0 19872 0 -1 45360
box -48 -56 240 834
use sg13g2_decap_8  FILLER_58_8
timestamp 1679581782
transform 1 0 1920 0 1 45360
box -48 -56 720 834
use sg13g2_decap_8  FILLER_58_15
timestamp 1679581782
transform 1 0 2592 0 1 45360
box -48 -56 720 834
use sg13g2_decap_4  FILLER_58_22
timestamp 1679577901
transform 1 0 3264 0 1 45360
box -48 -56 432 834
use sg13g2_fill_2  FILLER_58_26
timestamp 1677580104
transform 1 0 3648 0 1 45360
box -48 -56 240 834
use sg13g2_fill_2  FILLER_58_72
timestamp 1677580104
transform 1 0 8064 0 1 45360
box -48 -56 240 834
use sg13g2_decap_4  FILLER_58_129
timestamp 1679577901
transform 1 0 13536 0 1 45360
box -48 -56 432 834
use sg13g2_fill_1  FILLER_58_133
timestamp 1677579658
transform 1 0 13920 0 1 45360
box -48 -56 144 834
use sg13g2_decap_8  FILLER_58_155
timestamp 1679581782
transform 1 0 16032 0 1 45360
box -48 -56 720 834
use sg13g2_decap_4  FILLER_58_162
timestamp 1679577901
transform 1 0 16704 0 1 45360
box -48 -56 432 834
use sg13g2_fill_2  FILLER_58_166
timestamp 1677580104
transform 1 0 17088 0 1 45360
box -48 -56 240 834
use sg13g2_fill_1  FILLER_59_0
timestamp 1677579658
transform 1 0 1152 0 -1 46872
box -48 -56 144 834
use sg13g2_decap_8  FILLER_59_18
timestamp 1679581782
transform 1 0 2880 0 -1 46872
box -48 -56 720 834
use sg13g2_fill_1  FILLER_59_29
timestamp 1677579658
transform 1 0 3936 0 -1 46872
box -48 -56 144 834
use sg13g2_fill_2  FILLER_59_67
timestamp 1677580104
transform 1 0 7584 0 -1 46872
box -48 -56 240 834
use sg13g2_fill_1  FILLER_59_69
timestamp 1677579658
transform 1 0 7776 0 -1 46872
box -48 -56 144 834
use sg13g2_decap_4  FILLER_59_122
timestamp 1679577901
transform 1 0 12864 0 -1 46872
box -48 -56 432 834
use sg13g2_decap_8  FILLER_59_164
timestamp 1679581782
transform 1 0 16896 0 -1 46872
box -48 -56 720 834
use sg13g2_fill_2  FILLER_59_171
timestamp 1677580104
transform 1 0 17568 0 -1 46872
box -48 -56 240 834
use sg13g2_fill_2  FILLER_59_190
timestamp 1677580104
transform 1 0 19392 0 -1 46872
box -48 -56 240 834
use sg13g2_fill_1  FILLER_59_192
timestamp 1677579658
transform 1 0 19584 0 -1 46872
box -48 -56 144 834
use sg13g2_decap_4  FILLER_60_0
timestamp 1679577901
transform 1 0 1152 0 1 46872
box -48 -56 432 834
use sg13g2_decap_8  FILLER_60_42
timestamp 1679581782
transform 1 0 5184 0 1 46872
box -48 -56 720 834
use sg13g2_fill_1  FILLER_60_49
timestamp 1677579658
transform 1 0 5856 0 1 46872
box -48 -56 144 834
use sg13g2_decap_4  FILLER_60_91
timestamp 1679577901
transform 1 0 9888 0 1 46872
box -48 -56 432 834
use sg13g2_fill_1  FILLER_60_95
timestamp 1677579658
transform 1 0 10272 0 1 46872
box -48 -56 144 834
use sg13g2_fill_1  FILLER_60_99
timestamp 1677579658
transform 1 0 10656 0 1 46872
box -48 -56 144 834
use sg13g2_fill_2  FILLER_60_117
timestamp 1677580104
transform 1 0 12384 0 1 46872
box -48 -56 240 834
use sg13g2_fill_1  FILLER_60_119
timestamp 1677579658
transform 1 0 12576 0 1 46872
box -48 -56 144 834
use sg13g2_decap_4  FILLER_60_171
timestamp 1679577901
transform 1 0 17568 0 1 46872
box -48 -56 432 834
use sg13g2_fill_1  FILLER_60_192
timestamp 1677579658
transform 1 0 19584 0 1 46872
box -48 -56 144 834
use sg13g2_decap_8  FILLER_61_0
timestamp 1679581782
transform 1 0 1152 0 -1 48384
box -48 -56 720 834
use sg13g2_fill_2  FILLER_61_7
timestamp 1677580104
transform 1 0 1824 0 -1 48384
box -48 -56 240 834
use sg13g2_decap_8  FILLER_61_51
timestamp 1679581782
transform 1 0 6048 0 -1 48384
box -48 -56 720 834
use sg13g2_decap_8  FILLER_61_58
timestamp 1679581782
transform 1 0 6720 0 -1 48384
box -48 -56 720 834
use sg13g2_decap_4  FILLER_61_65
timestamp 1679577901
transform 1 0 7392 0 -1 48384
box -48 -56 432 834
use sg13g2_fill_1  FILLER_61_69
timestamp 1677579658
transform 1 0 7776 0 -1 48384
box -48 -56 144 834
use sg13g2_decap_8  FILLER_61_74
timestamp 1679581782
transform 1 0 8256 0 -1 48384
box -48 -56 720 834
use sg13g2_fill_1  FILLER_61_81
timestamp 1677579658
transform 1 0 8928 0 -1 48384
box -48 -56 144 834
use sg13g2_fill_2  FILLER_61_86
timestamp 1677580104
transform 1 0 9408 0 -1 48384
box -48 -56 240 834
use sg13g2_fill_2  FILLER_61_92
timestamp 1677580104
transform 1 0 9984 0 -1 48384
box -48 -56 240 834
use sg13g2_fill_1  FILLER_61_94
timestamp 1677579658
transform 1 0 10176 0 -1 48384
box -48 -56 144 834
use sg13g2_decap_8  FILLER_61_103
timestamp 1679581782
transform 1 0 11040 0 -1 48384
box -48 -56 720 834
use sg13g2_decap_8  FILLER_61_110
timestamp 1679581782
transform 1 0 11712 0 -1 48384
box -48 -56 720 834
use sg13g2_decap_4  FILLER_61_117
timestamp 1679577901
transform 1 0 12384 0 -1 48384
box -48 -56 432 834
use sg13g2_fill_1  FILLER_61_121
timestamp 1677579658
transform 1 0 12768 0 -1 48384
box -48 -56 144 834
use sg13g2_decap_8  FILLER_61_139
timestamp 1679581782
transform 1 0 14496 0 -1 48384
box -48 -56 720 834
use sg13g2_decap_4  FILLER_61_146
timestamp 1679577901
transform 1 0 15168 0 -1 48384
box -48 -56 432 834
use sg13g2_decap_4  FILLER_61_188
timestamp 1679577901
transform 1 0 19200 0 -1 48384
box -48 -56 432 834
use sg13g2_fill_1  FILLER_61_192
timestamp 1677579658
transform 1 0 19584 0 -1 48384
box -48 -56 144 834
use sg13g2_decap_8  FILLER_62_0
timestamp 1679581782
transform 1 0 1152 0 1 48384
box -48 -56 720 834
use sg13g2_decap_8  FILLER_62_7
timestamp 1679581782
transform 1 0 1824 0 1 48384
box -48 -56 720 834
use sg13g2_decap_8  FILLER_62_14
timestamp 1679581782
transform 1 0 2496 0 1 48384
box -48 -56 720 834
use sg13g2_decap_4  FILLER_62_21
timestamp 1679577901
transform 1 0 3168 0 1 48384
box -48 -56 432 834
use sg13g2_fill_2  FILLER_62_25
timestamp 1677580104
transform 1 0 3552 0 1 48384
box -48 -56 240 834
use sg13g2_decap_4  FILLER_62_31
timestamp 1679577901
transform 1 0 4128 0 1 48384
box -48 -56 432 834
use sg13g2_fill_1  FILLER_62_85
timestamp 1677579658
transform 1 0 9312 0 1 48384
box -48 -56 144 834
use sg13g2_fill_1  FILLER_62_90
timestamp 1677579658
transform 1 0 9792 0 1 48384
box -48 -56 144 834
use sg13g2_decap_8  FILLER_62_129
timestamp 1679581782
transform 1 0 13536 0 1 48384
box -48 -56 720 834
use sg13g2_decap_4  FILLER_62_136
timestamp 1679577901
transform 1 0 14208 0 1 48384
box -48 -56 432 834
use sg13g2_fill_1  FILLER_62_140
timestamp 1677579658
transform 1 0 14592 0 1 48384
box -48 -56 144 834
use sg13g2_decap_8  FILLER_62_166
timestamp 1679581782
transform 1 0 17088 0 1 48384
box -48 -56 720 834
use sg13g2_fill_2  FILLER_62_173
timestamp 1677580104
transform 1 0 17760 0 1 48384
box -48 -56 240 834
use sg13g2_fill_1  FILLER_62_200
timestamp 1677579658
transform 1 0 20352 0 1 48384
box -48 -56 144 834
use sg13g2_decap_8  FILLER_63_0
timestamp 1679581782
transform 1 0 1152 0 -1 49896
box -48 -56 720 834
use sg13g2_fill_1  FILLER_63_7
timestamp 1677579658
transform 1 0 1824 0 -1 49896
box -48 -56 144 834
use sg13g2_decap_4  FILLER_63_25
timestamp 1679577901
transform 1 0 3552 0 -1 49896
box -48 -56 432 834
use sg13g2_decap_4  FILLER_63_46
timestamp 1679577901
transform 1 0 5568 0 -1 49896
box -48 -56 432 834
use sg13g2_fill_1  FILLER_63_50
timestamp 1677579658
transform 1 0 5952 0 -1 49896
box -48 -56 144 834
use sg13g2_fill_2  FILLER_63_85
timestamp 1677580104
transform 1 0 9312 0 -1 49896
box -48 -56 240 834
use sg13g2_decap_8  FILLER_63_129
timestamp 1679581782
transform 1 0 13536 0 -1 49896
box -48 -56 720 834
use sg13g2_fill_1  FILLER_63_136
timestamp 1677579658
transform 1 0 14208 0 -1 49896
box -48 -56 144 834
use sg13g2_decap_8  FILLER_63_175
timestamp 1679581782
transform 1 0 17952 0 -1 49896
box -48 -56 720 834
use sg13g2_decap_8  FILLER_63_182
timestamp 1679581782
transform 1 0 18624 0 -1 49896
box -48 -56 720 834
use sg13g2_decap_8  FILLER_64_0
timestamp 1679581782
transform 1 0 1152 0 1 49896
box -48 -56 720 834
use sg13g2_fill_2  FILLER_64_7
timestamp 1677580104
transform 1 0 1824 0 1 49896
box -48 -56 240 834
use sg13g2_fill_2  FILLER_64_26
timestamp 1677580104
transform 1 0 3648 0 1 49896
box -48 -56 240 834
use sg13g2_fill_1  FILLER_64_28
timestamp 1677579658
transform 1 0 3840 0 1 49896
box -48 -56 144 834
use sg13g2_decap_8  FILLER_64_46
timestamp 1679581782
transform 1 0 5568 0 1 49896
box -48 -56 720 834
use sg13g2_decap_8  FILLER_64_53
timestamp 1679581782
transform 1 0 6240 0 1 49896
box -48 -56 720 834
use sg13g2_decap_4  FILLER_64_60
timestamp 1679577901
transform 1 0 6912 0 1 49896
box -48 -56 432 834
use sg13g2_fill_1  FILLER_64_64
timestamp 1677579658
transform 1 0 7296 0 1 49896
box -48 -56 144 834
use sg13g2_fill_1  FILLER_64_103
timestamp 1677579658
transform 1 0 11040 0 1 49896
box -48 -56 144 834
use sg13g2_fill_1  FILLER_64_108
timestamp 1677579658
transform 1 0 11520 0 1 49896
box -48 -56 144 834
use sg13g2_fill_1  FILLER_64_117
timestamp 1677579658
transform 1 0 12384 0 1 49896
box -48 -56 144 834
use sg13g2_decap_8  FILLER_64_173
timestamp 1679581782
transform 1 0 17760 0 1 49896
box -48 -56 720 834
use sg13g2_decap_4  FILLER_65_8
timestamp 1679577901
transform 1 0 1920 0 -1 51408
box -48 -56 432 834
use sg13g2_fill_2  FILLER_65_12
timestamp 1677580104
transform 1 0 2304 0 -1 51408
box -48 -56 240 834
use sg13g2_decap_8  FILLER_65_18
timestamp 1679581782
transform 1 0 2880 0 -1 51408
box -48 -56 720 834
use sg13g2_decap_8  FILLER_65_25
timestamp 1679581782
transform 1 0 3552 0 -1 51408
box -48 -56 720 834
use sg13g2_fill_2  FILLER_65_32
timestamp 1677580104
transform 1 0 4224 0 -1 51408
box -48 -56 240 834
use sg13g2_decap_8  FILLER_65_68
timestamp 1679581782
transform 1 0 7680 0 -1 51408
box -48 -56 720 834
use sg13g2_decap_4  FILLER_65_75
timestamp 1679577901
transform 1 0 8352 0 -1 51408
box -48 -56 432 834
use sg13g2_fill_1  FILLER_65_79
timestamp 1677579658
transform 1 0 8736 0 -1 51408
box -48 -56 144 834
use sg13g2_decap_8  FILLER_65_118
timestamp 1679581782
transform 1 0 12480 0 -1 51408
box -48 -56 720 834
use sg13g2_fill_1  FILLER_65_125
timestamp 1677579658
transform 1 0 13152 0 -1 51408
box -48 -56 144 834
use sg13g2_decap_8  FILLER_65_143
timestamp 1679581782
transform 1 0 14880 0 -1 51408
box -48 -56 720 834
use sg13g2_fill_1  FILLER_65_188
timestamp 1677579658
transform 1 0 19200 0 -1 51408
box -48 -56 144 834
use sg13g2_fill_1  FILLER_66_8
timestamp 1677579658
transform 1 0 1920 0 1 51408
box -48 -56 144 834
use sg13g2_decap_4  FILLER_66_42
timestamp 1679577901
transform 1 0 5184 0 1 51408
box -48 -56 432 834
use sg13g2_fill_2  FILLER_66_46
timestamp 1677580104
transform 1 0 5568 0 1 51408
box -48 -56 240 834
use sg13g2_fill_1  FILLER_66_86
timestamp 1677579658
transform 1 0 9408 0 1 51408
box -48 -56 144 834
use sg13g2_fill_2  FILLER_66_122
timestamp 1677580104
transform 1 0 12864 0 1 51408
box -48 -56 240 834
use sg13g2_fill_1  FILLER_66_124
timestamp 1677579658
transform 1 0 13056 0 1 51408
box -48 -56 144 834
use sg13g2_fill_1  FILLER_66_176
timestamp 1677579658
transform 1 0 18048 0 1 51408
box -48 -56 144 834
use sg13g2_fill_2  FILLER_66_194
timestamp 1677580104
transform 1 0 19776 0 1 51408
box -48 -56 240 834
use sg13g2_fill_1  FILLER_66_196
timestamp 1677579658
transform 1 0 19968 0 1 51408
box -48 -56 144 834
use sg13g2_decap_4  FILLER_67_21
timestamp 1679577901
transform 1 0 3168 0 -1 52920
box -48 -56 432 834
use sg13g2_decap_8  FILLER_67_63
timestamp 1679581782
transform 1 0 7200 0 -1 52920
box -48 -56 720 834
use sg13g2_fill_1  FILLER_67_70
timestamp 1677579658
transform 1 0 7872 0 -1 52920
box -48 -56 144 834
use sg13g2_fill_2  FILLER_67_194
timestamp 1677580104
transform 1 0 19776 0 -1 52920
box -48 -56 240 834
use sg13g2_fill_1  FILLER_67_196
timestamp 1677579658
transform 1 0 19968 0 -1 52920
box -48 -56 144 834
use sg13g2_fill_2  FILLER_68_4
timestamp 1677580104
transform 1 0 1536 0 1 52920
box -48 -56 240 834
use sg13g2_fill_1  FILLER_68_6
timestamp 1677579658
transform 1 0 1728 0 1 52920
box -48 -56 144 834
use sg13g2_fill_2  FILLER_68_11
timestamp 1677580104
transform 1 0 2208 0 1 52920
box -48 -56 240 834
use sg13g2_fill_1  FILLER_68_13
timestamp 1677579658
transform 1 0 2400 0 1 52920
box -48 -56 144 834
use sg13g2_fill_2  FILLER_68_35
timestamp 1677580104
transform 1 0 4512 0 1 52920
box -48 -56 240 834
use sg13g2_fill_1  FILLER_68_37
timestamp 1677579658
transform 1 0 4704 0 1 52920
box -48 -56 144 834
use sg13g2_fill_1  FILLER_68_55
timestamp 1677579658
transform 1 0 6432 0 1 52920
box -48 -56 144 834
use sg13g2_fill_1  FILLER_68_77
timestamp 1677579658
transform 1 0 8544 0 1 52920
box -48 -56 144 834
use sg13g2_fill_1  FILLER_68_83
timestamp 1677579658
transform 1 0 9120 0 1 52920
box -48 -56 144 834
use sg13g2_decap_8  FILLER_68_101
timestamp 1679581782
transform 1 0 10848 0 1 52920
box -48 -56 720 834
use sg13g2_decap_4  FILLER_68_108
timestamp 1679577901
transform 1 0 11520 0 1 52920
box -48 -56 432 834
use sg13g2_fill_2  FILLER_68_112
timestamp 1677580104
transform 1 0 11904 0 1 52920
box -48 -56 240 834
use sg13g2_decap_8  FILLER_68_122
timestamp 1679581782
transform 1 0 12864 0 1 52920
box -48 -56 720 834
use sg13g2_fill_2  FILLER_68_129
timestamp 1677580104
transform 1 0 13536 0 1 52920
box -48 -56 240 834
use sg13g2_fill_2  FILLER_68_177
timestamp 1677580104
transform 1 0 18144 0 1 52920
box -48 -56 240 834
use sg13g2_fill_1  FILLER_68_200
timestamp 1677579658
transform 1 0 20352 0 1 52920
box -48 -56 144 834
use sg13g2_fill_1  FILLER_69_4
timestamp 1677579658
transform 1 0 1536 0 -1 54432
box -48 -56 144 834
use sg13g2_decap_8  FILLER_69_72
timestamp 1679581782
transform 1 0 8064 0 -1 54432
box -48 -56 720 834
use sg13g2_decap_4  FILLER_69_79
timestamp 1679577901
transform 1 0 8736 0 -1 54432
box -48 -56 432 834
use sg13g2_fill_1  FILLER_69_83
timestamp 1677579658
transform 1 0 9120 0 -1 54432
box -48 -56 144 834
use sg13g2_fill_1  FILLER_69_126
timestamp 1677579658
transform 1 0 13248 0 -1 54432
box -48 -56 144 834
use sg13g2_fill_2  FILLER_69_198
timestamp 1677580104
transform 1 0 20160 0 -1 54432
box -48 -56 240 834
use sg13g2_fill_1  FILLER_69_200
timestamp 1677579658
transform 1 0 20352 0 -1 54432
box -48 -56 144 834
use sg13g2_fill_2  FILLER_70_0
timestamp 1677580104
transform 1 0 1152 0 1 54432
box -48 -56 240 834
use sg13g2_fill_2  FILLER_70_49
timestamp 1677580104
transform 1 0 5856 0 1 54432
box -48 -56 240 834
use sg13g2_fill_1  FILLER_70_51
timestamp 1677579658
transform 1 0 6048 0 1 54432
box -48 -56 144 834
use sg13g2_decap_4  FILLER_70_107
timestamp 1679577901
transform 1 0 11424 0 1 54432
box -48 -56 432 834
use sg13g2_fill_1  FILLER_70_111
timestamp 1677579658
transform 1 0 11808 0 1 54432
box -48 -56 144 834
use sg13g2_fill_1  FILLER_70_146
timestamp 1677579658
transform 1 0 15168 0 1 54432
box -48 -56 144 834
use sg13g2_fill_1  FILLER_70_164
timestamp 1677579658
transform 1 0 16896 0 1 54432
box -48 -56 144 834
use sg13g2_fill_2  FILLER_70_182
timestamp 1677580104
transform 1 0 18624 0 1 54432
box -48 -56 240 834
use sg13g2_fill_2  FILLER_71_0
timestamp 1677580104
transform 1 0 1152 0 -1 55944
box -48 -56 240 834
use sg13g2_fill_1  FILLER_71_27
timestamp 1677579658
transform 1 0 3744 0 -1 55944
box -48 -56 144 834
use sg13g2_fill_2  FILLER_71_53
timestamp 1677580104
transform 1 0 6240 0 -1 55944
box -48 -56 240 834
use sg13g2_fill_1  FILLER_71_55
timestamp 1677579658
transform 1 0 6432 0 -1 55944
box -48 -56 144 834
use sg13g2_fill_1  FILLER_71_73
timestamp 1677579658
transform 1 0 8160 0 -1 55944
box -48 -56 144 834
use sg13g2_fill_2  FILLER_71_95
timestamp 1677580104
transform 1 0 10272 0 -1 55944
box -48 -56 240 834
use sg13g2_fill_1  FILLER_71_97
timestamp 1677579658
transform 1 0 10464 0 -1 55944
box -48 -56 144 834
use sg13g2_decap_8  FILLER_71_119
timestamp 1679581782
transform 1 0 12576 0 -1 55944
box -48 -56 720 834
use sg13g2_fill_2  FILLER_71_126
timestamp 1677580104
transform 1 0 13248 0 -1 55944
box -48 -56 240 834
use sg13g2_fill_1  FILLER_71_128
timestamp 1677579658
transform 1 0 13440 0 -1 55944
box -48 -56 144 834
use sg13g2_fill_1  FILLER_71_192
timestamp 1677579658
transform 1 0 19584 0 -1 55944
box -48 -56 144 834
use sg13g2_fill_1  FILLER_72_4
timestamp 1677579658
transform 1 0 1536 0 1 55944
box -48 -56 144 834
use sg13g2_fill_1  FILLER_72_22
timestamp 1677579658
transform 1 0 3264 0 1 55944
box -48 -56 144 834
use sg13g2_decap_4  FILLER_72_48
timestamp 1679577901
transform 1 0 5760 0 1 55944
box -48 -56 432 834
use sg13g2_fill_2  FILLER_72_73
timestamp 1677580104
transform 1 0 8160 0 1 55944
box -48 -56 240 834
use sg13g2_fill_1  FILLER_72_75
timestamp 1677579658
transform 1 0 8352 0 1 55944
box -48 -56 144 834
use sg13g2_decap_8  FILLER_72_97
timestamp 1679581782
transform 1 0 10464 0 1 55944
box -48 -56 720 834
use sg13g2_decap_4  FILLER_72_104
timestamp 1679577901
transform 1 0 11136 0 1 55944
box -48 -56 432 834
use sg13g2_fill_1  FILLER_72_167
timestamp 1677579658
transform 1 0 17184 0 1 55944
box -48 -56 144 834
use sg13g2_decap_4  FILLER_73_62
timestamp 1679577901
transform 1 0 7104 0 -1 57456
box -48 -56 432 834
use sg13g2_fill_1  FILLER_73_66
timestamp 1677579658
transform 1 0 7488 0 -1 57456
box -48 -56 144 834
use sg13g2_fill_2  FILLER_73_88
timestamp 1677580104
transform 1 0 9600 0 -1 57456
box -48 -56 240 834
use sg13g2_fill_2  FILLER_73_145
timestamp 1677580104
transform 1 0 15072 0 -1 57456
box -48 -56 240 834
use sg13g2_fill_2  FILLER_73_198
timestamp 1677580104
transform 1 0 20160 0 -1 57456
box -48 -56 240 834
use sg13g2_fill_1  FILLER_73_200
timestamp 1677579658
transform 1 0 20352 0 -1 57456
box -48 -56 144 834
use sg13g2_fill_2  FILLER_74_0
timestamp 1677580104
transform 1 0 1152 0 1 57456
box -48 -56 240 834
use sg13g2_fill_1  FILLER_74_2
timestamp 1677579658
transform 1 0 1344 0 1 57456
box -48 -56 144 834
use sg13g2_fill_2  FILLER_74_20
timestamp 1677580104
transform 1 0 3072 0 1 57456
box -48 -56 240 834
use sg13g2_fill_1  FILLER_74_22
timestamp 1677579658
transform 1 0 3264 0 1 57456
box -48 -56 144 834
use sg13g2_decap_8  FILLER_74_82
timestamp 1679581782
transform 1 0 9024 0 1 57456
box -48 -56 720 834
use sg13g2_fill_1  FILLER_74_89
timestamp 1677579658
transform 1 0 9696 0 1 57456
box -48 -56 144 834
use sg13g2_fill_2  FILLER_74_138
timestamp 1677580104
transform 1 0 14400 0 1 57456
box -48 -56 240 834
use sg13g2_fill_2  FILLER_74_157
timestamp 1677580104
transform 1 0 16224 0 1 57456
box -48 -56 240 834
use sg13g2_fill_1  FILLER_74_159
timestamp 1677579658
transform 1 0 16416 0 1 57456
box -48 -56 144 834
use sg13g2_fill_2  FILLER_74_198
timestamp 1677580104
transform 1 0 20160 0 1 57456
box -48 -56 240 834
use sg13g2_fill_1  FILLER_74_200
timestamp 1677579658
transform 1 0 20352 0 1 57456
box -48 -56 144 834
use sg13g2_fill_2  FILLER_75_8
timestamp 1677580104
transform 1 0 1920 0 -1 58968
box -48 -56 240 834
use sg13g2_fill_2  FILLER_75_56
timestamp 1677580104
transform 1 0 6528 0 -1 58968
box -48 -56 240 834
use sg13g2_fill_1  FILLER_75_96
timestamp 1677579658
transform 1 0 10368 0 -1 58968
box -48 -56 144 834
use sg13g2_fill_2  FILLER_75_108
timestamp 1677580104
transform 1 0 11520 0 -1 58968
box -48 -56 240 834
use sg13g2_decap_4  FILLER_75_114
timestamp 1679577901
transform 1 0 12096 0 -1 58968
box -48 -56 432 834
use sg13g2_fill_2  FILLER_75_118
timestamp 1677580104
transform 1 0 12480 0 -1 58968
box -48 -56 240 834
use sg13g2_fill_1  FILLER_75_128
timestamp 1677579658
transform 1 0 13440 0 -1 58968
box -48 -56 144 834
use sg13g2_fill_1  FILLER_75_146
timestamp 1677579658
transform 1 0 15168 0 -1 58968
box -48 -56 144 834
use sg13g2_fill_1  FILLER_75_181
timestamp 1677579658
transform 1 0 18528 0 -1 58968
box -48 -56 144 834
use sg13g2_fill_2  FILLER_75_199
timestamp 1677580104
transform 1 0 20256 0 -1 58968
box -48 -56 240 834
use sg13g2_fill_1  FILLER_76_21
timestamp 1677579658
transform 1 0 3168 0 1 58968
box -48 -56 144 834
use sg13g2_fill_1  FILLER_76_68
timestamp 1677579658
transform 1 0 7680 0 1 58968
box -48 -56 144 834
use sg13g2_fill_2  FILLER_76_77
timestamp 1677580104
transform 1 0 8544 0 1 58968
box -48 -56 240 834
use sg13g2_fill_2  FILLER_76_96
timestamp 1677580104
transform 1 0 10368 0 1 58968
box -48 -56 240 834
use sg13g2_fill_2  FILLER_76_123
timestamp 1677580104
transform 1 0 12960 0 1 58968
box -48 -56 240 834
use sg13g2_fill_2  FILLER_76_159
timestamp 1677580104
transform 1 0 16416 0 1 58968
box -48 -56 240 834
use sg13g2_fill_2  FILLER_76_199
timestamp 1677580104
transform 1 0 20256 0 1 58968
box -48 -56 240 834
use sg13g2_fill_1  FILLER_77_8
timestamp 1677579658
transform 1 0 1920 0 -1 60480
box -48 -56 144 834
use sg13g2_fill_1  FILLER_77_47
timestamp 1677579658
transform 1 0 5664 0 -1 60480
box -48 -56 144 834
use sg13g2_fill_2  FILLER_77_65
timestamp 1677580104
transform 1 0 7392 0 -1 60480
box -48 -56 240 834
use sg13g2_decap_8  FILLER_77_71
timestamp 1679581782
transform 1 0 7968 0 -1 60480
box -48 -56 720 834
use sg13g2_decap_4  FILLER_77_78
timestamp 1679577901
transform 1 0 8640 0 -1 60480
box -48 -56 432 834
use sg13g2_fill_1  FILLER_77_120
timestamp 1677579658
transform 1 0 12672 0 -1 60480
box -48 -56 144 834
use sg13g2_fill_2  FILLER_77_129
timestamp 1677580104
transform 1 0 13536 0 -1 60480
box -48 -56 240 834
use sg13g2_fill_1  FILLER_77_139
timestamp 1677579658
transform 1 0 14496 0 -1 60480
box -48 -56 144 834
use sg13g2_fill_2  FILLER_77_175
timestamp 1677580104
transform 1 0 17952 0 -1 60480
box -48 -56 240 834
use sg13g2_fill_1  FILLER_77_177
timestamp 1677579658
transform 1 0 18144 0 -1 60480
box -48 -56 144 834
use sg13g2_fill_2  FILLER_77_199
timestamp 1677580104
transform 1 0 20256 0 -1 60480
box -48 -56 240 834
use sg13g2_fill_2  FILLER_78_21
timestamp 1677580104
transform 1 0 3168 0 1 60480
box -48 -56 240 834
use sg13g2_fill_1  FILLER_78_23
timestamp 1677579658
transform 1 0 3360 0 1 60480
box -48 -56 144 834
use sg13g2_fill_1  FILLER_78_91
timestamp 1677579658
transform 1 0 9888 0 1 60480
box -48 -56 144 834
use sg13g2_decap_4  FILLER_78_109
timestamp 1679577901
transform 1 0 11616 0 1 60480
box -48 -56 432 834
use sg13g2_fill_1  FILLER_78_113
timestamp 1677579658
transform 1 0 12000 0 1 60480
box -48 -56 144 834
use sg13g2_fill_1  FILLER_78_139
timestamp 1677579658
transform 1 0 14496 0 1 60480
box -48 -56 144 834
use sg13g2_fill_2  FILLER_78_178
timestamp 1677580104
transform 1 0 18240 0 1 60480
box -48 -56 240 834
use sg13g2_fill_1  FILLER_78_180
timestamp 1677579658
transform 1 0 18432 0 1 60480
box -48 -56 144 834
use sg13g2_fill_2  FILLER_78_198
timestamp 1677580104
transform 1 0 20160 0 1 60480
box -48 -56 240 834
use sg13g2_fill_1  FILLER_78_200
timestamp 1677579658
transform 1 0 20352 0 1 60480
box -48 -56 144 834
use sg13g2_fill_1  FILLER_79_4
timestamp 1677579658
transform 1 0 1536 0 -1 61992
box -48 -56 144 834
use sg13g2_fill_2  FILLER_79_47
timestamp 1677580104
transform 1 0 5664 0 -1 61992
box -48 -56 240 834
use sg13g2_fill_2  FILLER_79_108
timestamp 1677580104
transform 1 0 11520 0 -1 61992
box -48 -56 240 834
use sg13g2_fill_1  FILLER_79_148
timestamp 1677579658
transform 1 0 15360 0 -1 61992
box -48 -56 144 834
use sg13g2_fill_2  FILLER_79_199
timestamp 1677580104
transform 1 0 20256 0 -1 61992
box -48 -56 240 834
use sg13g2_fill_1  FILLER_80_21
timestamp 1677579658
transform 1 0 3168 0 1 61992
box -48 -56 144 834
use sg13g2_fill_2  FILLER_80_43
timestamp 1677580104
transform 1 0 5280 0 1 61992
box -48 -56 240 834
use sg13g2_fill_1  FILLER_80_45
timestamp 1677579658
transform 1 0 5472 0 1 61992
box -48 -56 144 834
use sg13g2_fill_2  FILLER_80_88
timestamp 1677580104
transform 1 0 9600 0 1 61992
box -48 -56 240 834
use sg13g2_fill_2  FILLER_80_111
timestamp 1677580104
transform 1 0 11808 0 1 61992
box -48 -56 240 834
use sg13g2_fill_2  FILLER_80_138
timestamp 1677580104
transform 1 0 14400 0 1 61992
box -48 -56 240 834
use sg13g2_fill_1  FILLER_80_178
timestamp 1677579658
transform 1 0 18240 0 1 61992
box -48 -56 144 834
use sg13g2_fill_1  FILLER_80_196
timestamp 1677579658
transform 1 0 19968 0 1 61992
box -48 -56 144 834
use sg13g2_fill_1  FILLER_81_4
timestamp 1677579658
transform 1 0 1536 0 -1 63504
box -48 -56 144 834
use sg13g2_fill_2  FILLER_81_26
timestamp 1677580104
transform 1 0 3648 0 -1 63504
box -48 -56 240 834
use sg13g2_fill_2  FILLER_81_93
timestamp 1677580104
transform 1 0 10080 0 -1 63504
box -48 -56 240 834
use sg13g2_fill_2  FILLER_81_112
timestamp 1677580104
transform 1 0 11904 0 -1 63504
box -48 -56 240 834
use sg13g2_decap_4  FILLER_81_118
timestamp 1679577901
transform 1 0 12480 0 -1 63504
box -48 -56 432 834
use sg13g2_fill_2  FILLER_81_168
timestamp 1677580104
transform 1 0 17280 0 -1 63504
box -48 -56 240 834
use sg13g2_fill_1  FILLER_81_170
timestamp 1677579658
transform 1 0 17472 0 -1 63504
box -48 -56 144 834
use sg13g2_fill_1  FILLER_81_196
timestamp 1677579658
transform 1 0 19968 0 -1 63504
box -48 -56 144 834
use sg13g2_fill_2  FILLER_82_0
timestamp 1677580104
transform 1 0 1152 0 1 63504
box -48 -56 240 834
use sg13g2_fill_1  FILLER_82_2
timestamp 1677579658
transform 1 0 1344 0 1 63504
box -48 -56 144 834
use sg13g2_fill_2  FILLER_82_45
timestamp 1677580104
transform 1 0 5472 0 1 63504
box -48 -56 240 834
use sg13g2_fill_2  FILLER_82_90
timestamp 1677580104
transform 1 0 9792 0 1 63504
box -48 -56 240 834
use sg13g2_fill_2  FILLER_82_113
timestamp 1677580104
transform 1 0 12000 0 1 63504
box -48 -56 240 834
use sg13g2_fill_1  FILLER_82_115
timestamp 1677579658
transform 1 0 12192 0 1 63504
box -48 -56 144 834
use sg13g2_fill_1  FILLER_82_153
timestamp 1677579658
transform 1 0 15840 0 1 63504
box -48 -56 144 834
use sg13g2_fill_1  FILLER_82_200
timestamp 1677579658
transform 1 0 20352 0 1 63504
box -48 -56 144 834
use sg13g2_fill_2  FILLER_83_8
timestamp 1677580104
transform 1 0 1920 0 -1 65016
box -48 -56 240 834
use sg13g2_fill_2  FILLER_83_56
timestamp 1677580104
transform 1 0 6528 0 -1 65016
box -48 -56 240 834
use sg13g2_fill_1  FILLER_83_58
timestamp 1677579658
transform 1 0 6720 0 -1 65016
box -48 -56 144 834
use sg13g2_fill_2  FILLER_83_84
timestamp 1677580104
transform 1 0 9216 0 -1 65016
box -48 -56 240 834
use sg13g2_decap_8  FILLER_83_107
timestamp 1679581782
transform 1 0 11424 0 -1 65016
box -48 -56 720 834
use sg13g2_fill_1  FILLER_83_114
timestamp 1677579658
transform 1 0 12096 0 -1 65016
box -48 -56 144 834
use sg13g2_fill_2  FILLER_83_157
timestamp 1677580104
transform 1 0 16224 0 -1 65016
box -48 -56 240 834
use sg13g2_fill_1  FILLER_83_159
timestamp 1677579658
transform 1 0 16416 0 -1 65016
box -48 -56 144 834
use sg13g2_fill_1  FILLER_83_177
timestamp 1677579658
transform 1 0 18144 0 -1 65016
box -48 -56 144 834
use sg13g2_fill_2  FILLER_83_195
timestamp 1677580104
transform 1 0 19872 0 -1 65016
box -48 -56 240 834
use sg13g2_fill_2  FILLER_84_0
timestamp 1677580104
transform 1 0 1152 0 1 65016
box -48 -56 240 834
use sg13g2_fill_1  FILLER_84_2
timestamp 1677579658
transform 1 0 1344 0 1 65016
box -48 -56 144 834
use sg13g2_fill_2  FILLER_84_28
timestamp 1677580104
transform 1 0 3840 0 1 65016
box -48 -56 240 834
use sg13g2_decap_4  FILLER_84_106
timestamp 1679577901
transform 1 0 11328 0 1 65016
box -48 -56 432 834
use sg13g2_fill_1  FILLER_84_143
timestamp 1677579658
transform 1 0 14880 0 1 65016
box -48 -56 144 834
use sg13g2_fill_2  FILLER_84_199
timestamp 1677580104
transform 1 0 20256 0 1 65016
box -48 -56 240 834
use sg13g2_fill_2  FILLER_85_12
timestamp 1677580104
transform 1 0 2304 0 -1 66528
box -48 -56 240 834
use sg13g2_fill_2  FILLER_85_35
timestamp 1677580104
transform 1 0 4512 0 -1 66528
box -48 -56 240 834
use sg13g2_fill_2  FILLER_85_54
timestamp 1677580104
transform 1 0 6336 0 -1 66528
box -48 -56 240 834
use sg13g2_fill_2  FILLER_85_68
timestamp 1677580104
transform 1 0 7680 0 -1 66528
box -48 -56 240 834
use sg13g2_fill_2  FILLER_85_87
timestamp 1677580104
transform 1 0 9504 0 -1 66528
box -48 -56 240 834
use sg13g2_fill_1  FILLER_85_89
timestamp 1677579658
transform 1 0 9696 0 -1 66528
box -48 -56 144 834
use sg13g2_decap_8  FILLER_85_107
timestamp 1679581782
transform 1 0 11424 0 -1 66528
box -48 -56 720 834
use sg13g2_decap_4  FILLER_85_114
timestamp 1679577901
transform 1 0 12096 0 -1 66528
box -48 -56 432 834
use sg13g2_fill_1  FILLER_85_118
timestamp 1677579658
transform 1 0 12480 0 -1 66528
box -48 -56 144 834
use sg13g2_fill_1  FILLER_85_140
timestamp 1677579658
transform 1 0 14592 0 -1 66528
box -48 -56 144 834
use sg13g2_fill_2  FILLER_85_170
timestamp 1677580104
transform 1 0 17472 0 -1 66528
box -48 -56 240 834
use sg13g2_fill_1  FILLER_86_4
timestamp 1677579658
transform 1 0 1536 0 1 66528
box -48 -56 144 834
use sg13g2_fill_1  FILLER_86_85
timestamp 1677579658
transform 1 0 9312 0 1 66528
box -48 -56 144 834
use sg13g2_fill_1  FILLER_86_128
timestamp 1677579658
transform 1 0 13440 0 1 66528
box -48 -56 144 834
use sg13g2_fill_1  FILLER_86_200
timestamp 1677579658
transform 1 0 20352 0 1 66528
box -48 -56 144 834
use sg13g2_fill_1  FILLER_87_0
timestamp 1677579658
transform 1 0 1152 0 -1 68040
box -48 -56 144 834
use sg13g2_fill_1  FILLER_87_63
timestamp 1677579658
transform 1 0 7200 0 -1 68040
box -48 -56 144 834
use sg13g2_fill_1  FILLER_87_85
timestamp 1677579658
transform 1 0 9312 0 -1 68040
box -48 -56 144 834
use sg13g2_fill_2  FILLER_87_158
timestamp 1677580104
transform 1 0 16320 0 -1 68040
box -48 -56 240 834
use sg13g2_fill_2  FILLER_87_198
timestamp 1677580104
transform 1 0 20160 0 -1 68040
box -48 -56 240 834
use sg13g2_fill_1  FILLER_87_200
timestamp 1677579658
transform 1 0 20352 0 -1 68040
box -48 -56 144 834
use sg13g2_fill_1  FILLER_88_25
timestamp 1677579658
transform 1 0 3552 0 1 68040
box -48 -56 144 834
use sg13g2_fill_2  FILLER_88_93
timestamp 1677580104
transform 1 0 10080 0 1 68040
box -48 -56 240 834
use sg13g2_fill_1  FILLER_88_95
timestamp 1677579658
transform 1 0 10272 0 1 68040
box -48 -56 144 834
use sg13g2_fill_1  FILLER_88_113
timestamp 1677579658
transform 1 0 12000 0 1 68040
box -48 -56 144 834
use sg13g2_fill_2  FILLER_88_139
timestamp 1677580104
transform 1 0 14496 0 1 68040
box -48 -56 240 834
use sg13g2_fill_1  FILLER_88_162
timestamp 1677579658
transform 1 0 16704 0 1 68040
box -48 -56 144 834
use sg13g2_fill_2  FILLER_88_167
timestamp 1677580104
transform 1 0 17184 0 1 68040
box -48 -56 240 834
use sg13g2_fill_1  FILLER_88_169
timestamp 1677579658
transform 1 0 17376 0 1 68040
box -48 -56 144 834
use sg13g2_fill_2  FILLER_88_187
timestamp 1677580104
transform 1 0 19104 0 1 68040
box -48 -56 240 834
use sg13g2_fill_1  FILLER_88_189
timestamp 1677579658
transform 1 0 19296 0 1 68040
box -48 -56 144 834
use sg13g2_fill_2  FILLER_88_194
timestamp 1677580104
transform 1 0 19776 0 1 68040
box -48 -56 240 834
use sg13g2_fill_1  FILLER_88_196
timestamp 1677579658
transform 1 0 19968 0 1 68040
box -48 -56 144 834
use sg13g2_fill_2  FILLER_89_0
timestamp 1677580104
transform 1 0 1152 0 -1 69552
box -48 -56 240 834
use sg13g2_fill_1  FILLER_89_74
timestamp 1677579658
transform 1 0 8256 0 -1 69552
box -48 -56 144 834
use sg13g2_decap_8  FILLER_89_100
timestamp 1679581782
transform 1 0 10752 0 -1 69552
box -48 -56 720 834
use sg13g2_fill_2  FILLER_89_124
timestamp 1677580104
transform 1 0 13056 0 -1 69552
box -48 -56 240 834
use sg13g2_fill_1  FILLER_89_130
timestamp 1677579658
transform 1 0 13632 0 -1 69552
box -48 -56 144 834
use sg13g2_fill_2  FILLER_89_198
timestamp 1677580104
transform 1 0 20160 0 -1 69552
box -48 -56 240 834
use sg13g2_fill_1  FILLER_89_200
timestamp 1677579658
transform 1 0 20352 0 -1 69552
box -48 -56 144 834
use sg13g2_fill_2  FILLER_90_0
timestamp 1677580104
transform 1 0 1152 0 1 69552
box -48 -56 240 834
use sg13g2_fill_1  FILLER_90_2
timestamp 1677579658
transform 1 0 1344 0 1 69552
box -48 -56 144 834
use sg13g2_fill_2  FILLER_90_20
timestamp 1677580104
transform 1 0 3072 0 1 69552
box -48 -56 240 834
use sg13g2_fill_2  FILLER_90_85
timestamp 1677580104
transform 1 0 9312 0 1 69552
box -48 -56 240 834
use sg13g2_decap_8  FILLER_90_108
timestamp 1679581782
transform 1 0 11520 0 1 69552
box -48 -56 720 834
use sg13g2_fill_1  FILLER_90_115
timestamp 1677579658
transform 1 0 12192 0 1 69552
box -48 -56 144 834
use sg13g2_fill_1  FILLER_90_137
timestamp 1677579658
transform 1 0 14304 0 1 69552
box -48 -56 144 834
use sg13g2_fill_2  FILLER_90_159
timestamp 1677580104
transform 1 0 16416 0 1 69552
box -48 -56 240 834
use sg13g2_fill_1  FILLER_90_161
timestamp 1677579658
transform 1 0 16608 0 1 69552
box -48 -56 144 834
use sg13g2_fill_2  FILLER_90_191
timestamp 1677580104
transform 1 0 19488 0 1 69552
box -48 -56 240 834
use sg13g2_fill_2  FILLER_91_29
timestamp 1677580104
transform 1 0 3936 0 -1 71064
box -48 -56 240 834
use sg13g2_fill_1  FILLER_91_31
timestamp 1677579658
transform 1 0 4128 0 -1 71064
box -48 -56 144 834
use sg13g2_fill_1  FILLER_91_61
timestamp 1677579658
transform 1 0 7008 0 -1 71064
box -48 -56 144 834
use sg13g2_fill_2  FILLER_91_84
timestamp 1677580104
transform 1 0 9216 0 -1 71064
box -48 -56 240 834
use sg13g2_fill_1  FILLER_91_107
timestamp 1677579658
transform 1 0 11424 0 -1 71064
box -48 -56 144 834
use sg13g2_fill_2  FILLER_91_129
timestamp 1677580104
transform 1 0 13536 0 -1 71064
box -48 -56 240 834
use sg13g2_fill_2  FILLER_91_148
timestamp 1677580104
transform 1 0 15360 0 -1 71064
box -48 -56 240 834
use sg13g2_fill_1  FILLER_91_150
timestamp 1677579658
transform 1 0 15552 0 -1 71064
box -48 -56 144 834
use sg13g2_fill_2  FILLER_91_172
timestamp 1677580104
transform 1 0 17664 0 -1 71064
box -48 -56 240 834
use sg13g2_fill_1  FILLER_91_174
timestamp 1677579658
transform 1 0 17856 0 -1 71064
box -48 -56 144 834
use sg13g2_fill_1  FILLER_91_200
timestamp 1677579658
transform 1 0 20352 0 -1 71064
box -48 -56 144 834
use sg13g2_fill_2  FILLER_92_4
timestamp 1677580104
transform 1 0 1536 0 1 71064
box -48 -56 240 834
use sg13g2_fill_1  FILLER_92_6
timestamp 1677579658
transform 1 0 1728 0 1 71064
box -48 -56 144 834
use sg13g2_fill_1  FILLER_92_15
timestamp 1677579658
transform 1 0 2592 0 1 71064
box -48 -56 144 834
use sg13g2_fill_2  FILLER_92_54
timestamp 1677580104
transform 1 0 6336 0 1 71064
box -48 -56 240 834
use sg13g2_fill_1  FILLER_92_56
timestamp 1677579658
transform 1 0 6528 0 1 71064
box -48 -56 144 834
use sg13g2_fill_2  FILLER_92_74
timestamp 1677580104
transform 1 0 8256 0 1 71064
box -48 -56 240 834
use sg13g2_fill_1  FILLER_92_76
timestamp 1677579658
transform 1 0 8448 0 1 71064
box -48 -56 144 834
use sg13g2_fill_2  FILLER_92_136
timestamp 1677580104
transform 1 0 14208 0 1 71064
box -48 -56 240 834
use sg13g2_fill_1  FILLER_92_138
timestamp 1677579658
transform 1 0 14400 0 1 71064
box -48 -56 144 834
use sg13g2_fill_2  FILLER_92_164
timestamp 1677580104
transform 1 0 16896 0 1 71064
box -48 -56 240 834
use sg13g2_fill_1  FILLER_92_166
timestamp 1677579658
transform 1 0 17088 0 1 71064
box -48 -56 144 834
use sg13g2_fill_1  FILLER_92_196
timestamp 1677579658
transform 1 0 19968 0 1 71064
box -48 -56 144 834
use sg13g2_fill_2  FILLER_93_49
timestamp 1677580104
transform 1 0 5856 0 -1 72576
box -48 -56 240 834
use sg13g2_fill_1  FILLER_93_51
timestamp 1677579658
transform 1 0 6048 0 -1 72576
box -48 -56 144 834
use sg13g2_decap_4  FILLER_93_101
timestamp 1679577901
transform 1 0 10848 0 -1 72576
box -48 -56 432 834
use sg13g2_fill_2  FILLER_93_109
timestamp 1677580104
transform 1 0 11616 0 -1 72576
box -48 -56 240 834
use sg13g2_fill_1  FILLER_93_111
timestamp 1677579658
transform 1 0 11808 0 -1 72576
box -48 -56 144 834
use sg13g2_fill_2  FILLER_93_163
timestamp 1677580104
transform 1 0 16800 0 -1 72576
box -48 -56 240 834
use sg13g2_fill_1  FILLER_93_165
timestamp 1677579658
transform 1 0 16992 0 -1 72576
box -48 -56 144 834
use sg13g2_fill_2  FILLER_93_176
timestamp 1677580104
transform 1 0 18048 0 -1 72576
box -48 -56 240 834
use sg13g2_fill_2  FILLER_93_199
timestamp 1677580104
transform 1 0 20256 0 -1 72576
box -48 -56 240 834
use sg13g2_fill_1  FILLER_94_0
timestamp 1677579658
transform 1 0 1152 0 1 72576
box -48 -56 144 834
use sg13g2_fill_1  FILLER_94_56
timestamp 1677579658
transform 1 0 6528 0 1 72576
box -48 -56 144 834
use sg13g2_fill_2  FILLER_94_82
timestamp 1677580104
transform 1 0 9024 0 1 72576
box -48 -56 240 834
use sg13g2_fill_1  FILLER_94_84
timestamp 1677579658
transform 1 0 9216 0 1 72576
box -48 -56 144 834
use sg13g2_fill_2  FILLER_94_119
timestamp 1677580104
transform 1 0 12576 0 1 72576
box -48 -56 240 834
use sg13g2_fill_1  FILLER_94_196
timestamp 1677579658
transform 1 0 19968 0 1 72576
box -48 -56 144 834
use sg13g2_fill_1  FILLER_95_0
timestamp 1677579658
transform 1 0 1152 0 -1 74088
box -48 -56 144 834
use sg13g2_fill_2  FILLER_95_39
timestamp 1677580104
transform 1 0 4896 0 -1 74088
box -48 -56 240 834
use sg13g2_fill_2  FILLER_95_96
timestamp 1677580104
transform 1 0 10368 0 -1 74088
box -48 -56 240 834
use sg13g2_fill_1  FILLER_95_144
timestamp 1677579658
transform 1 0 14976 0 -1 74088
box -48 -56 144 834
use sg13g2_fill_1  FILLER_95_157
timestamp 1677579658
transform 1 0 16224 0 -1 74088
box -48 -56 144 834
use sg13g2_fill_2  FILLER_95_175
timestamp 1677580104
transform 1 0 17952 0 -1 74088
box -48 -56 240 834
use sg13g2_fill_1  FILLER_96_21
timestamp 1677579658
transform 1 0 3168 0 1 74088
box -48 -56 144 834
use sg13g2_fill_2  FILLER_96_67
timestamp 1677580104
transform 1 0 7584 0 1 74088
box -48 -56 240 834
use sg13g2_fill_1  FILLER_96_111
timestamp 1677579658
transform 1 0 11808 0 1 74088
box -48 -56 144 834
use sg13g2_fill_2  FILLER_96_133
timestamp 1677580104
transform 1 0 13920 0 1 74088
box -48 -56 240 834
use sg13g2_fill_1  FILLER_96_135
timestamp 1677579658
transform 1 0 14112 0 1 74088
box -48 -56 144 834
use sg13g2_fill_2  FILLER_96_157
timestamp 1677580104
transform 1 0 16224 0 1 74088
box -48 -56 240 834
use sg13g2_fill_1  FILLER_96_159
timestamp 1677579658
transform 1 0 16416 0 1 74088
box -48 -56 144 834
use sg13g2_fill_2  FILLER_96_194
timestamp 1677580104
transform 1 0 19776 0 1 74088
box -48 -56 240 834
use sg13g2_fill_1  FILLER_96_196
timestamp 1677579658
transform 1 0 19968 0 1 74088
box -48 -56 144 834
use sg13g2_fill_2  FILLER_97_12
timestamp 1677580104
transform 1 0 2304 0 -1 75600
box -48 -56 240 834
use sg13g2_fill_1  FILLER_97_14
timestamp 1677579658
transform 1 0 2496 0 -1 75600
box -48 -56 144 834
use sg13g2_fill_1  FILLER_97_83
timestamp 1677579658
transform 1 0 9120 0 -1 75600
box -48 -56 144 834
use sg13g2_decap_8  FILLER_97_105
timestamp 1679581782
transform 1 0 11232 0 -1 75600
box -48 -56 720 834
use sg13g2_decap_4  FILLER_97_112
timestamp 1679577901
transform 1 0 11904 0 -1 75600
box -48 -56 432 834
use sg13g2_fill_2  FILLER_97_116
timestamp 1677580104
transform 1 0 12288 0 -1 75600
box -48 -56 240 834
use sg13g2_fill_1  FILLER_98_21
timestamp 1677579658
transform 1 0 3168 0 1 75600
box -48 -56 144 834
use sg13g2_fill_1  FILLER_98_93
timestamp 1677579658
transform 1 0 10080 0 1 75600
box -48 -56 144 834
use sg13g2_fill_1  FILLER_98_111
timestamp 1677579658
transform 1 0 11808 0 1 75600
box -48 -56 144 834
use sg13g2_fill_1  FILLER_98_133
timestamp 1677579658
transform 1 0 13920 0 1 75600
box -48 -56 144 834
use sg13g2_fill_2  FILLER_99_0
timestamp 1677580104
transform 1 0 1152 0 -1 77112
box -48 -56 240 834
use sg13g2_fill_2  FILLER_99_48
timestamp 1677580104
transform 1 0 5760 0 -1 77112
box -48 -56 240 834
use sg13g2_fill_1  FILLER_99_50
timestamp 1677579658
transform 1 0 5952 0 -1 77112
box -48 -56 144 834
use sg13g2_fill_2  FILLER_99_106
timestamp 1677580104
transform 1 0 11328 0 -1 77112
box -48 -56 240 834
use sg13g2_fill_2  FILLER_99_125
timestamp 1677580104
transform 1 0 13152 0 -1 77112
box -48 -56 240 834
use sg13g2_fill_2  FILLER_100_8
timestamp 1677580104
transform 1 0 1920 0 1 77112
box -48 -56 240 834
use sg13g2_fill_2  FILLER_100_44
timestamp 1677580104
transform 1 0 5376 0 1 77112
box -48 -56 240 834
use sg13g2_fill_1  FILLER_100_46
timestamp 1677579658
transform 1 0 5568 0 1 77112
box -48 -56 144 834
use sg13g2_fill_1  FILLER_100_81
timestamp 1677579658
transform 1 0 8928 0 1 77112
box -48 -56 144 834
use sg13g2_fill_2  FILLER_100_141
timestamp 1677580104
transform 1 0 14688 0 1 77112
box -48 -56 240 834
use sg13g2_fill_1  FILLER_100_143
timestamp 1677579658
transform 1 0 14880 0 1 77112
box -48 -56 144 834
use sg13g2_fill_2  FILLER_101_17
timestamp 1677580104
transform 1 0 2784 0 -1 78624
box -48 -56 240 834
use sg13g2_fill_1  FILLER_101_62
timestamp 1677579658
transform 1 0 7104 0 -1 78624
box -48 -56 144 834
use sg13g2_fill_2  FILLER_101_138
timestamp 1677580104
transform 1 0 14400 0 -1 78624
box -48 -56 240 834
use sg13g2_fill_1  FILLER_101_140
timestamp 1677579658
transform 1 0 14592 0 -1 78624
box -48 -56 144 834
use sg13g2_fill_2  FILLER_102_26
timestamp 1677580104
transform 1 0 3648 0 1 78624
box -48 -56 240 834
use sg13g2_fill_1  FILLER_102_65
timestamp 1677579658
transform 1 0 7392 0 1 78624
box -48 -56 144 834
use sg13g2_fill_2  FILLER_102_95
timestamp 1677580104
transform 1 0 10272 0 1 78624
box -48 -56 240 834
use sg13g2_fill_2  FILLER_102_101
timestamp 1677580104
transform 1 0 10848 0 1 78624
box -48 -56 240 834
use sg13g2_fill_2  FILLER_102_128
timestamp 1677580104
transform 1 0 13440 0 1 78624
box -48 -56 240 834
use sg13g2_fill_2  FILLER_102_198
timestamp 1677580104
transform 1 0 20160 0 1 78624
box -48 -56 240 834
use sg13g2_fill_1  FILLER_102_200
timestamp 1677579658
transform 1 0 20352 0 1 78624
box -48 -56 144 834
use sg13g2_fill_2  FILLER_103_0
timestamp 1677580104
transform 1 0 1152 0 -1 80136
box -48 -56 240 834
use sg13g2_fill_1  FILLER_103_2
timestamp 1677579658
transform 1 0 1344 0 -1 80136
box -48 -56 144 834
use sg13g2_fill_1  FILLER_103_32
timestamp 1677579658
transform 1 0 4224 0 -1 80136
box -48 -56 144 834
use sg13g2_fill_2  FILLER_103_100
timestamp 1677580104
transform 1 0 10752 0 -1 80136
box -48 -56 240 834
use sg13g2_fill_1  FILLER_103_102
timestamp 1677579658
transform 1 0 10944 0 -1 80136
box -48 -56 144 834
use sg13g2_fill_2  FILLER_103_107
timestamp 1677580104
transform 1 0 11424 0 -1 80136
box -48 -56 240 834
use sg13g2_fill_1  FILLER_103_109
timestamp 1677579658
transform 1 0 11616 0 -1 80136
box -48 -56 144 834
use sg13g2_fill_2  FILLER_103_158
timestamp 1677580104
transform 1 0 16320 0 -1 80136
box -48 -56 240 834
use sg13g2_fill_1  FILLER_103_160
timestamp 1677579658
transform 1 0 16512 0 -1 80136
box -48 -56 144 834
use sg13g2_fill_2  FILLER_103_186
timestamp 1677580104
transform 1 0 19008 0 -1 80136
box -48 -56 240 834
use sg13g2_fill_1  FILLER_103_188
timestamp 1677579658
transform 1 0 19200 0 -1 80136
box -48 -56 144 834
use sg13g2_fill_1  FILLER_104_4
timestamp 1677579658
transform 1 0 1536 0 1 80136
box -48 -56 144 834
use sg13g2_fill_1  FILLER_104_116
timestamp 1677579658
transform 1 0 12288 0 1 80136
box -48 -56 144 834
use sg13g2_fill_1  FILLER_104_142
timestamp 1677579658
transform 1 0 14784 0 1 80136
box -48 -56 144 834
use sg13g2_fill_2  FILLER_104_198
timestamp 1677580104
transform 1 0 20160 0 1 80136
box -48 -56 240 834
use sg13g2_fill_1  FILLER_104_200
timestamp 1677579658
transform 1 0 20352 0 1 80136
box -48 -56 144 834
use sg13g2_fill_1  FILLER_105_81
timestamp 1677579658
transform 1 0 8928 0 -1 81648
box -48 -56 144 834
use sg13g2_fill_1  FILLER_105_103
timestamp 1677579658
transform 1 0 11040 0 -1 81648
box -48 -56 144 834
use sg13g2_fill_2  FILLER_105_125
timestamp 1677580104
transform 1 0 13152 0 -1 81648
box -48 -56 240 834
use sg13g2_fill_1  FILLER_105_127
timestamp 1677579658
transform 1 0 13344 0 -1 81648
box -48 -56 144 834
use sg13g2_fill_2  FILLER_105_167
timestamp 1677580104
transform 1 0 17184 0 -1 81648
box -48 -56 240 834
use sg13g2_fill_1  FILLER_105_169
timestamp 1677579658
transform 1 0 17376 0 -1 81648
box -48 -56 144 834
use sg13g2_fill_2  FILLER_105_199
timestamp 1677580104
transform 1 0 20256 0 -1 81648
box -48 -56 240 834
use sg13g2_fill_2  FILLER_106_0
timestamp 1677580104
transform 1 0 1152 0 1 81648
box -48 -56 240 834
use sg13g2_fill_1  FILLER_106_2
timestamp 1677579658
transform 1 0 1344 0 1 81648
box -48 -56 144 834
use sg13g2_fill_1  FILLER_106_72
timestamp 1677579658
transform 1 0 8064 0 1 81648
box -48 -56 144 834
use sg13g2_fill_2  FILLER_106_101
timestamp 1677580104
transform 1 0 10848 0 1 81648
box -48 -56 240 834
use sg13g2_fill_2  FILLER_106_124
timestamp 1677580104
transform 1 0 13056 0 1 81648
box -48 -56 240 834
use sg13g2_fill_1  FILLER_106_126
timestamp 1677579658
transform 1 0 13248 0 1 81648
box -48 -56 144 834
use sg13g2_fill_1  FILLER_106_177
timestamp 1677579658
transform 1 0 18144 0 1 81648
box -48 -56 144 834
use sg13g2_fill_2  FILLER_106_199
timestamp 1677580104
transform 1 0 20256 0 1 81648
box -48 -56 240 834
use sg13g2_fill_2  FILLER_107_0
timestamp 1677580104
transform 1 0 1152 0 -1 83160
box -48 -56 240 834
use sg13g2_fill_1  FILLER_107_2
timestamp 1677579658
transform 1 0 1344 0 -1 83160
box -48 -56 144 834
use sg13g2_fill_2  FILLER_107_58
timestamp 1677580104
transform 1 0 6720 0 -1 83160
box -48 -56 240 834
use sg13g2_decap_8  FILLER_107_94
timestamp 1679581782
transform 1 0 10176 0 -1 83160
box -48 -56 720 834
use sg13g2_decap_4  FILLER_107_101
timestamp 1679577901
transform 1 0 10848 0 -1 83160
box -48 -56 432 834
use sg13g2_fill_1  FILLER_107_126
timestamp 1677579658
transform 1 0 13248 0 -1 83160
box -48 -56 144 834
use sg13g2_fill_2  FILLER_107_131
timestamp 1677580104
transform 1 0 13728 0 -1 83160
box -48 -56 240 834
use sg13g2_fill_1  FILLER_107_133
timestamp 1677579658
transform 1 0 13920 0 -1 83160
box -48 -56 144 834
use sg13g2_fill_2  FILLER_107_161
timestamp 1677580104
transform 1 0 16608 0 -1 83160
box -48 -56 240 834
use sg13g2_fill_2  FILLER_108_0
timestamp 1677580104
transform 1 0 1152 0 1 83160
box -48 -56 240 834
use sg13g2_fill_1  FILLER_108_2
timestamp 1677579658
transform 1 0 1344 0 1 83160
box -48 -56 144 834
use sg13g2_fill_2  FILLER_108_20
timestamp 1677580104
transform 1 0 3072 0 1 83160
box -48 -56 240 834
use sg13g2_fill_1  FILLER_108_86
timestamp 1677579658
transform 1 0 9408 0 1 83160
box -48 -56 144 834
use sg13g2_decap_4  FILLER_108_125
timestamp 1679577901
transform 1 0 13152 0 1 83160
box -48 -56 432 834
use sg13g2_fill_2  FILLER_108_137
timestamp 1677580104
transform 1 0 14304 0 1 83160
box -48 -56 240 834
use sg13g2_fill_2  FILLER_108_148
timestamp 1677580104
transform 1 0 15360 0 1 83160
box -48 -56 240 834
use sg13g2_fill_1  FILLER_108_150
timestamp 1677579658
transform 1 0 15552 0 1 83160
box -48 -56 144 834
use sg13g2_fill_2  FILLER_109_12
timestamp 1677580104
transform 1 0 2304 0 -1 84672
box -48 -56 240 834
use sg13g2_fill_1  FILLER_109_14
timestamp 1677579658
transform 1 0 2496 0 -1 84672
box -48 -56 144 834
use sg13g2_fill_2  FILLER_109_78
timestamp 1677580104
transform 1 0 8640 0 -1 84672
box -48 -56 240 834
use sg13g2_fill_2  FILLER_109_118
timestamp 1677580104
transform 1 0 12480 0 -1 84672
box -48 -56 240 834
use sg13g2_fill_2  FILLER_109_169
timestamp 1677580104
transform 1 0 17376 0 -1 84672
box -48 -56 240 834
use sg13g2_fill_1  FILLER_109_171
timestamp 1677579658
transform 1 0 17568 0 -1 84672
box -48 -56 144 834
use sg13g2_fill_2  FILLER_110_0
timestamp 1677580104
transform 1 0 1152 0 1 84672
box -48 -56 240 834
use sg13g2_fill_2  FILLER_110_40
timestamp 1677580104
transform 1 0 4992 0 1 84672
box -48 -56 240 834
use sg13g2_fill_1  FILLER_110_64
timestamp 1677579658
transform 1 0 7296 0 1 84672
box -48 -56 144 834
use sg13g2_fill_2  FILLER_110_141
timestamp 1677580104
transform 1 0 14688 0 1 84672
box -48 -56 240 834
use sg13g2_fill_1  FILLER_110_143
timestamp 1677579658
transform 1 0 14880 0 1 84672
box -48 -56 144 834
use sg13g2_fill_2  FILLER_110_199
timestamp 1677580104
transform 1 0 20256 0 1 84672
box -48 -56 240 834
use sg13g2_fill_1  FILLER_111_4
timestamp 1677579658
transform 1 0 1536 0 -1 86184
box -48 -56 144 834
use sg13g2_fill_2  FILLER_111_30
timestamp 1677580104
transform 1 0 4032 0 -1 86184
box -48 -56 240 834
use sg13g2_fill_1  FILLER_111_32
timestamp 1677579658
transform 1 0 4224 0 -1 86184
box -48 -56 144 834
use sg13g2_fill_1  FILLER_111_50
timestamp 1677579658
transform 1 0 5952 0 -1 86184
box -48 -56 144 834
use sg13g2_fill_2  FILLER_111_59
timestamp 1677580104
transform 1 0 6816 0 -1 86184
box -48 -56 240 834
use sg13g2_fill_1  FILLER_111_61
timestamp 1677579658
transform 1 0 7008 0 -1 86184
box -48 -56 144 834
use sg13g2_fill_2  FILLER_111_113
timestamp 1677580104
transform 1 0 12000 0 -1 86184
box -48 -56 240 834
use sg13g2_fill_1  FILLER_111_115
timestamp 1677579658
transform 1 0 12192 0 -1 86184
box -48 -56 144 834
use sg13g2_fill_2  FILLER_111_198
timestamp 1677580104
transform 1 0 20160 0 -1 86184
box -48 -56 240 834
use sg13g2_fill_1  FILLER_111_200
timestamp 1677579658
transform 1 0 20352 0 -1 86184
box -48 -56 144 834
use sg13g2_fill_1  FILLER_112_0
timestamp 1677579658
transform 1 0 1152 0 1 86184
box -48 -56 144 834
use sg13g2_fill_2  FILLER_112_89
timestamp 1677580104
transform 1 0 9696 0 1 86184
box -48 -56 240 834
use sg13g2_fill_1  FILLER_112_91
timestamp 1677579658
transform 1 0 9888 0 1 86184
box -48 -56 144 834
use sg13g2_fill_2  FILLER_112_129
timestamp 1677580104
transform 1 0 13536 0 1 86184
box -48 -56 240 834
use sg13g2_fill_1  FILLER_112_131
timestamp 1677579658
transform 1 0 13728 0 1 86184
box -48 -56 144 834
use sg13g2_fill_2  FILLER_112_166
timestamp 1677580104
transform 1 0 17088 0 1 86184
box -48 -56 240 834
use sg13g2_fill_1  FILLER_112_168
timestamp 1677579658
transform 1 0 17280 0 1 86184
box -48 -56 144 834
use sg13g2_fill_2  FILLER_112_190
timestamp 1677580104
transform 1 0 19392 0 1 86184
box -48 -56 240 834
use sg13g2_fill_1  FILLER_112_192
timestamp 1677579658
transform 1 0 19584 0 1 86184
box -48 -56 144 834
use sg13g2_fill_1  FILLER_113_58
timestamp 1677579658
transform 1 0 6720 0 -1 87696
box -48 -56 144 834
use sg13g2_fill_2  FILLER_113_97
timestamp 1677580104
transform 1 0 10464 0 -1 87696
box -48 -56 240 834
use sg13g2_decap_8  FILLER_113_130
timestamp 1679581782
transform 1 0 13632 0 -1 87696
box -48 -56 720 834
use sg13g2_decap_8  FILLER_113_137
timestamp 1679581782
transform 1 0 14304 0 -1 87696
box -48 -56 720 834
use sg13g2_decap_8  FILLER_113_144
timestamp 1679581782
transform 1 0 14976 0 -1 87696
box -48 -56 720 834
use sg13g2_fill_1  FILLER_113_168
timestamp 1677579658
transform 1 0 17280 0 -1 87696
box -48 -56 144 834
use sg13g2_fill_2  FILLER_113_190
timestamp 1677580104
transform 1 0 19392 0 -1 87696
box -48 -56 240 834
use sg13g2_fill_1  FILLER_113_192
timestamp 1677579658
transform 1 0 19584 0 -1 87696
box -48 -56 144 834
use sg13g2_fill_2  FILLER_114_4
timestamp 1677580104
transform 1 0 1536 0 1 87696
box -48 -56 240 834
use sg13g2_fill_1  FILLER_114_6
timestamp 1677579658
transform 1 0 1728 0 1 87696
box -48 -56 144 834
use sg13g2_fill_1  FILLER_114_15
timestamp 1677579658
transform 1 0 2592 0 1 87696
box -48 -56 144 834
use sg13g2_fill_2  FILLER_114_75
timestamp 1677580104
transform 1 0 8352 0 1 87696
box -48 -56 240 834
use sg13g2_fill_1  FILLER_114_77
timestamp 1677579658
transform 1 0 8544 0 1 87696
box -48 -56 144 834
use sg13g2_fill_2  FILLER_114_116
timestamp 1677580104
transform 1 0 12288 0 1 87696
box -48 -56 240 834
use sg13g2_fill_2  FILLER_114_198
timestamp 1677580104
transform 1 0 20160 0 1 87696
box -48 -56 240 834
use sg13g2_fill_1  FILLER_114_200
timestamp 1677579658
transform 1 0 20352 0 1 87696
box -48 -56 144 834
use sg13g2_fill_1  FILLER_115_33
timestamp 1677579658
transform 1 0 4320 0 -1 89208
box -48 -56 144 834
use sg13g2_decap_4  FILLER_115_55
timestamp 1679577901
transform 1 0 6432 0 -1 89208
box -48 -56 432 834
use sg13g2_fill_2  FILLER_115_59
timestamp 1677580104
transform 1 0 6816 0 -1 89208
box -48 -56 240 834
use sg13g2_decap_4  FILLER_115_78
timestamp 1679577901
transform 1 0 8640 0 -1 89208
box -48 -56 432 834
use sg13g2_fill_1  FILLER_115_82
timestamp 1677579658
transform 1 0 9024 0 -1 89208
box -48 -56 144 834
use sg13g2_fill_1  FILLER_115_95
timestamp 1677579658
transform 1 0 10272 0 -1 89208
box -48 -56 144 834
use sg13g2_decap_4  FILLER_115_159
timestamp 1679577901
transform 1 0 16416 0 -1 89208
box -48 -56 432 834
use sg13g2_fill_1  FILLER_115_180
timestamp 1677579658
transform 1 0 18432 0 -1 89208
box -48 -56 144 834
use sg13g2_decap_8  FILLER_116_53
timestamp 1679581782
transform 1 0 6240 0 1 89208
box -48 -56 720 834
use sg13g2_decap_8  FILLER_116_60
timestamp 1679581782
transform 1 0 6912 0 1 89208
box -48 -56 720 834
use sg13g2_decap_8  FILLER_116_67
timestamp 1679581782
transform 1 0 7584 0 1 89208
box -48 -56 720 834
use sg13g2_decap_8  FILLER_116_74
timestamp 1679581782
transform 1 0 8256 0 1 89208
box -48 -56 720 834
use sg13g2_decap_8  FILLER_116_81
timestamp 1679581782
transform 1 0 8928 0 1 89208
box -48 -56 720 834
use sg13g2_decap_8  FILLER_116_88
timestamp 1679581782
transform 1 0 9600 0 1 89208
box -48 -56 720 834
use sg13g2_decap_8  FILLER_116_95
timestamp 1679581782
transform 1 0 10272 0 1 89208
box -48 -56 720 834
use sg13g2_decap_4  FILLER_116_102
timestamp 1679577901
transform 1 0 10944 0 1 89208
box -48 -56 432 834
use sg13g2_fill_2  FILLER_116_161
timestamp 1677580104
transform 1 0 16608 0 1 89208
box -48 -56 240 834
use sg13g2_decap_4  FILLER_116_180
timestamp 1679577901
transform 1 0 18432 0 1 89208
box -48 -56 432 834
use sg13g2_fill_1  FILLER_116_184
timestamp 1677579658
transform 1 0 18816 0 1 89208
box -48 -56 144 834
use sg13g2_decap_8  FILLER_117_32
timestamp 1679581782
transform 1 0 4224 0 -1 90720
box -48 -56 720 834
use sg13g2_decap_8  FILLER_117_39
timestamp 1679581782
transform 1 0 4896 0 -1 90720
box -48 -56 720 834
use sg13g2_decap_8  FILLER_117_46
timestamp 1679581782
transform 1 0 5568 0 -1 90720
box -48 -56 720 834
use sg13g2_decap_8  FILLER_117_53
timestamp 1679581782
transform 1 0 6240 0 -1 90720
box -48 -56 720 834
use sg13g2_decap_8  FILLER_117_60
timestamp 1679581782
transform 1 0 6912 0 -1 90720
box -48 -56 720 834
use sg13g2_decap_8  FILLER_117_67
timestamp 1679581782
transform 1 0 7584 0 -1 90720
box -48 -56 720 834
use sg13g2_decap_8  FILLER_117_74
timestamp 1679581782
transform 1 0 8256 0 -1 90720
box -48 -56 720 834
use sg13g2_decap_8  FILLER_117_81
timestamp 1679581782
transform 1 0 8928 0 -1 90720
box -48 -56 720 834
use sg13g2_decap_8  FILLER_117_88
timestamp 1679581782
transform 1 0 9600 0 -1 90720
box -48 -56 720 834
use sg13g2_decap_8  FILLER_117_95
timestamp 1679581782
transform 1 0 10272 0 -1 90720
box -48 -56 720 834
use sg13g2_decap_4  FILLER_117_102
timestamp 1679577901
transform 1 0 10944 0 -1 90720
box -48 -56 432 834
use sg13g2_decap_8  FILLER_117_123
timestamp 1679581782
transform 1 0 12960 0 -1 90720
box -48 -56 720 834
use sg13g2_decap_8  FILLER_117_130
timestamp 1679581782
transform 1 0 13632 0 -1 90720
box -48 -56 720 834
use sg13g2_decap_8  FILLER_117_154
timestamp 1679581782
transform 1 0 15936 0 -1 90720
box -48 -56 720 834
use sg13g2_decap_4  FILLER_117_161
timestamp 1679577901
transform 1 0 16608 0 -1 90720
box -48 -56 432 834
use sg13g2_decap_8  FILLER_117_169
timestamp 1679581782
transform 1 0 17376 0 -1 90720
box -48 -56 720 834
use sg13g2_decap_8  FILLER_117_176
timestamp 1679581782
transform 1 0 18048 0 -1 90720
box -48 -56 720 834
use sg13g2_decap_4  FILLER_117_183
timestamp 1679577901
transform 1 0 18720 0 -1 90720
box -48 -56 432 834
use sg13g2_fill_2  FILLER_117_187
timestamp 1677580104
transform 1 0 19104 0 -1 90720
box -48 -56 240 834
use sg13g2_decap_8  FILLER_118_20
timestamp 1679581782
transform 1 0 3072 0 1 90720
box -48 -56 720 834
use sg13g2_decap_8  FILLER_118_27
timestamp 1679581782
transform 1 0 3744 0 1 90720
box -48 -56 720 834
use sg13g2_decap_8  FILLER_118_34
timestamp 1679581782
transform 1 0 4416 0 1 90720
box -48 -56 720 834
use sg13g2_decap_8  FILLER_118_41
timestamp 1679581782
transform 1 0 5088 0 1 90720
box -48 -56 720 834
use sg13g2_decap_8  FILLER_118_48
timestamp 1679581782
transform 1 0 5760 0 1 90720
box -48 -56 720 834
use sg13g2_decap_8  FILLER_118_55
timestamp 1679581782
transform 1 0 6432 0 1 90720
box -48 -56 720 834
use sg13g2_decap_4  FILLER_118_62
timestamp 1679577901
transform 1 0 7104 0 1 90720
box -48 -56 432 834
use sg13g2_fill_2  FILLER_118_66
timestamp 1677580104
transform 1 0 7488 0 1 90720
box -48 -56 240 834
use sg13g2_decap_8  FILLER_118_76
timestamp 1679581782
transform 1 0 8448 0 1 90720
box -48 -56 720 834
use sg13g2_decap_8  FILLER_118_83
timestamp 1679581782
transform 1 0 9120 0 1 90720
box -48 -56 720 834
use sg13g2_decap_8  FILLER_118_90
timestamp 1679581782
transform 1 0 9792 0 1 90720
box -48 -56 720 834
use sg13g2_decap_8  FILLER_118_97
timestamp 1679581782
transform 1 0 10464 0 1 90720
box -48 -56 720 834
use sg13g2_decap_8  FILLER_118_104
timestamp 1679581782
transform 1 0 11136 0 1 90720
box -48 -56 720 834
use sg13g2_decap_8  FILLER_118_111
timestamp 1679581782
transform 1 0 11808 0 1 90720
box -48 -56 720 834
use sg13g2_decap_8  FILLER_118_118
timestamp 1679581782
transform 1 0 12480 0 1 90720
box -48 -56 720 834
use sg13g2_decap_8  FILLER_118_125
timestamp 1679581782
transform 1 0 13152 0 1 90720
box -48 -56 720 834
use sg13g2_decap_8  FILLER_118_132
timestamp 1679581782
transform 1 0 13824 0 1 90720
box -48 -56 720 834
use sg13g2_decap_8  FILLER_118_139
timestamp 1679581782
transform 1 0 14496 0 1 90720
box -48 -56 720 834
use sg13g2_decap_8  FILLER_118_146
timestamp 1679581782
transform 1 0 15168 0 1 90720
box -48 -56 720 834
use sg13g2_decap_8  FILLER_118_153
timestamp 1679581782
transform 1 0 15840 0 1 90720
box -48 -56 720 834
use sg13g2_decap_8  FILLER_118_160
timestamp 1679581782
transform 1 0 16512 0 1 90720
box -48 -56 720 834
use sg13g2_decap_8  FILLER_118_167
timestamp 1679581782
transform 1 0 17184 0 1 90720
box -48 -56 720 834
use sg13g2_decap_8  FILLER_118_174
timestamp 1679581782
transform 1 0 17856 0 1 90720
box -48 -56 720 834
use sg13g2_decap_8  FILLER_118_181
timestamp 1679581782
transform 1 0 18528 0 1 90720
box -48 -56 720 834
use sg13g2_decap_4  FILLER_118_188
timestamp 1679577901
transform 1 0 19200 0 1 90720
box -48 -56 432 834
use sg13g2_fill_1  FILLER_118_192
timestamp 1677579658
transform 1 0 19584 0 1 90720
box -48 -56 144 834
use sg13g2_decap_8  FILLER_119_20
timestamp 1679581782
transform 1 0 3072 0 -1 92232
box -48 -56 720 834
use sg13g2_decap_8  FILLER_119_27
timestamp 1679581782
transform 1 0 3744 0 -1 92232
box -48 -56 720 834
use sg13g2_decap_8  FILLER_119_34
timestamp 1679581782
transform 1 0 4416 0 -1 92232
box -48 -56 720 834
use sg13g2_decap_8  FILLER_119_41
timestamp 1679581782
transform 1 0 5088 0 -1 92232
box -48 -56 720 834
use sg13g2_decap_8  FILLER_119_48
timestamp 1679581782
transform 1 0 5760 0 -1 92232
box -48 -56 720 834
use sg13g2_decap_8  FILLER_119_55
timestamp 1679581782
transform 1 0 6432 0 -1 92232
box -48 -56 720 834
use sg13g2_decap_8  FILLER_119_62
timestamp 1679581782
transform 1 0 7104 0 -1 92232
box -48 -56 720 834
use sg13g2_decap_8  FILLER_119_73
timestamp 1679581782
transform 1 0 8160 0 -1 92232
box -48 -56 720 834
use sg13g2_decap_8  FILLER_119_80
timestamp 1679581782
transform 1 0 8832 0 -1 92232
box -48 -56 720 834
use sg13g2_decap_8  FILLER_119_87
timestamp 1679581782
transform 1 0 9504 0 -1 92232
box -48 -56 720 834
use sg13g2_decap_8  FILLER_119_94
timestamp 1679581782
transform 1 0 10176 0 -1 92232
box -48 -56 720 834
use sg13g2_decap_8  FILLER_119_101
timestamp 1679581782
transform 1 0 10848 0 -1 92232
box -48 -56 720 834
use sg13g2_decap_8  FILLER_119_108
timestamp 1679581782
transform 1 0 11520 0 -1 92232
box -48 -56 720 834
use sg13g2_decap_8  FILLER_119_115
timestamp 1679581782
transform 1 0 12192 0 -1 92232
box -48 -56 720 834
use sg13g2_decap_8  FILLER_119_122
timestamp 1679581782
transform 1 0 12864 0 -1 92232
box -48 -56 720 834
use sg13g2_decap_8  FILLER_119_129
timestamp 1679581782
transform 1 0 13536 0 -1 92232
box -48 -56 720 834
use sg13g2_decap_8  FILLER_119_136
timestamp 1679581782
transform 1 0 14208 0 -1 92232
box -48 -56 720 834
use sg13g2_decap_8  FILLER_119_143
timestamp 1679581782
transform 1 0 14880 0 -1 92232
box -48 -56 720 834
use sg13g2_decap_8  FILLER_119_150
timestamp 1679581782
transform 1 0 15552 0 -1 92232
box -48 -56 720 834
use sg13g2_decap_8  FILLER_119_157
timestamp 1679581782
transform 1 0 16224 0 -1 92232
box -48 -56 720 834
use sg13g2_decap_8  FILLER_119_164
timestamp 1679581782
transform 1 0 16896 0 -1 92232
box -48 -56 720 834
use sg13g2_decap_8  FILLER_119_171
timestamp 1679581782
transform 1 0 17568 0 -1 92232
box -48 -56 720 834
use sg13g2_decap_8  FILLER_119_178
timestamp 1679581782
transform 1 0 18240 0 -1 92232
box -48 -56 720 834
use sg13g2_decap_4  FILLER_119_185
timestamp 1679577901
transform 1 0 18912 0 -1 92232
box -48 -56 432 834
use sg13g2_decap_8  FILLER_120_20
timestamp 1679581782
transform 1 0 3072 0 1 92232
box -48 -56 720 834
use sg13g2_decap_8  FILLER_120_27
timestamp 1679581782
transform 1 0 3744 0 1 92232
box -48 -56 720 834
use sg13g2_decap_8  FILLER_120_34
timestamp 1679581782
transform 1 0 4416 0 1 92232
box -48 -56 720 834
use sg13g2_decap_8  FILLER_120_41
timestamp 1679581782
transform 1 0 5088 0 1 92232
box -48 -56 720 834
use sg13g2_decap_8  FILLER_120_48
timestamp 1679581782
transform 1 0 5760 0 1 92232
box -48 -56 720 834
use sg13g2_decap_8  FILLER_120_55
timestamp 1679581782
transform 1 0 6432 0 1 92232
box -48 -56 720 834
use sg13g2_decap_8  FILLER_120_62
timestamp 1679581782
transform 1 0 7104 0 1 92232
box -48 -56 720 834
use sg13g2_decap_8  FILLER_120_69
timestamp 1679581782
transform 1 0 7776 0 1 92232
box -48 -56 720 834
use sg13g2_decap_8  FILLER_120_76
timestamp 1679581782
transform 1 0 8448 0 1 92232
box -48 -56 720 834
use sg13g2_decap_8  FILLER_120_83
timestamp 1679581782
transform 1 0 9120 0 1 92232
box -48 -56 720 834
use sg13g2_decap_8  FILLER_120_90
timestamp 1679581782
transform 1 0 9792 0 1 92232
box -48 -56 720 834
use sg13g2_decap_8  FILLER_120_97
timestamp 1679581782
transform 1 0 10464 0 1 92232
box -48 -56 720 834
use sg13g2_decap_8  FILLER_120_104
timestamp 1679581782
transform 1 0 11136 0 1 92232
box -48 -56 720 834
use sg13g2_decap_8  FILLER_120_111
timestamp 1679581782
transform 1 0 11808 0 1 92232
box -48 -56 720 834
use sg13g2_decap_8  FILLER_120_118
timestamp 1679581782
transform 1 0 12480 0 1 92232
box -48 -56 720 834
use sg13g2_decap_8  FILLER_120_125
timestamp 1679581782
transform 1 0 13152 0 1 92232
box -48 -56 720 834
use sg13g2_decap_8  FILLER_120_132
timestamp 1679581782
transform 1 0 13824 0 1 92232
box -48 -56 720 834
use sg13g2_decap_8  FILLER_120_139
timestamp 1679581782
transform 1 0 14496 0 1 92232
box -48 -56 720 834
use sg13g2_decap_8  FILLER_120_146
timestamp 1679581782
transform 1 0 15168 0 1 92232
box -48 -56 720 834
use sg13g2_decap_8  FILLER_120_153
timestamp 1679581782
transform 1 0 15840 0 1 92232
box -48 -56 720 834
use sg13g2_decap_8  FILLER_120_160
timestamp 1679581782
transform 1 0 16512 0 1 92232
box -48 -56 720 834
use sg13g2_decap_8  FILLER_120_167
timestamp 1679581782
transform 1 0 17184 0 1 92232
box -48 -56 720 834
use sg13g2_decap_8  FILLER_120_174
timestamp 1679581782
transform 1 0 17856 0 1 92232
box -48 -56 720 834
use sg13g2_decap_8  FILLER_121_24
timestamp 1679581782
transform 1 0 3456 0 -1 93744
box -48 -56 720 834
use sg13g2_decap_8  FILLER_121_31
timestamp 1679581782
transform 1 0 4128 0 -1 93744
box -48 -56 720 834
use sg13g2_decap_8  FILLER_121_38
timestamp 1679581782
transform 1 0 4800 0 -1 93744
box -48 -56 720 834
use sg13g2_decap_8  FILLER_121_45
timestamp 1679581782
transform 1 0 5472 0 -1 93744
box -48 -56 720 834
use sg13g2_decap_8  FILLER_121_52
timestamp 1679581782
transform 1 0 6144 0 -1 93744
box -48 -56 720 834
use sg13g2_decap_8  FILLER_121_59
timestamp 1679581782
transform 1 0 6816 0 -1 93744
box -48 -56 720 834
use sg13g2_decap_8  FILLER_121_66
timestamp 1679581782
transform 1 0 7488 0 -1 93744
box -48 -56 720 834
use sg13g2_decap_8  FILLER_121_73
timestamp 1679581782
transform 1 0 8160 0 -1 93744
box -48 -56 720 834
use sg13g2_decap_8  FILLER_121_80
timestamp 1679581782
transform 1 0 8832 0 -1 93744
box -48 -56 720 834
use sg13g2_decap_8  FILLER_121_87
timestamp 1679581782
transform 1 0 9504 0 -1 93744
box -48 -56 720 834
use sg13g2_decap_8  FILLER_121_94
timestamp 1679581782
transform 1 0 10176 0 -1 93744
box -48 -56 720 834
use sg13g2_decap_8  FILLER_121_101
timestamp 1679581782
transform 1 0 10848 0 -1 93744
box -48 -56 720 834
use sg13g2_decap_8  FILLER_121_108
timestamp 1679581782
transform 1 0 11520 0 -1 93744
box -48 -56 720 834
use sg13g2_decap_8  FILLER_121_115
timestamp 1679581782
transform 1 0 12192 0 -1 93744
box -48 -56 720 834
use sg13g2_decap_8  FILLER_121_122
timestamp 1679581782
transform 1 0 12864 0 -1 93744
box -48 -56 720 834
use sg13g2_decap_8  FILLER_121_129
timestamp 1679581782
transform 1 0 13536 0 -1 93744
box -48 -56 720 834
use sg13g2_decap_8  FILLER_121_136
timestamp 1679581782
transform 1 0 14208 0 -1 93744
box -48 -56 720 834
use sg13g2_decap_8  FILLER_121_143
timestamp 1679581782
transform 1 0 14880 0 -1 93744
box -48 -56 720 834
use sg13g2_decap_8  FILLER_121_150
timestamp 1679581782
transform 1 0 15552 0 -1 93744
box -48 -56 720 834
use sg13g2_decap_8  FILLER_121_157
timestamp 1679581782
transform 1 0 16224 0 -1 93744
box -48 -56 720 834
use sg13g2_decap_8  FILLER_121_164
timestamp 1679581782
transform 1 0 16896 0 -1 93744
box -48 -56 720 834
use sg13g2_fill_2  FILLER_121_171
timestamp 1677580104
transform 1 0 17568 0 -1 93744
box -48 -56 240 834
use sg13g2_fill_1  FILLER_122_24
timestamp 1677579658
transform 1 0 3456 0 1 93744
box -48 -56 144 834
use sg13g2_decap_8  FILLER_122_105
timestamp 1679581782
transform 1 0 11232 0 1 93744
box -48 -56 720 834
use sg13g2_decap_8  FILLER_122_112
timestamp 1679581782
transform 1 0 11904 0 1 93744
box -48 -56 720 834
use sg13g2_fill_2  FILLER_122_135
timestamp 1677580104
transform 1 0 14112 0 1 93744
box -48 -56 240 834
use sg13g2_decap_8  FILLER_122_149
timestamp 1679581782
transform 1 0 15456 0 1 93744
box -48 -56 720 834
use sg13g2_fill_1  FILLER_122_200
timestamp 1677579658
transform 1 0 20352 0 1 93744
box -48 -56 144 834
use sg13g2_fill_1  FILLER_123_0
timestamp 1677579658
transform 1 0 1152 0 -1 95256
box -48 -56 144 834
use sg13g2_decap_4  FILLER_123_145
timestamp 1679577901
transform 1 0 15072 0 -1 95256
box -48 -56 432 834
use sg13g2_fill_2  FILLER_123_149
timestamp 1677580104
transform 1 0 15456 0 -1 95256
box -48 -56 240 834
use sg13g2_fill_2  FILLER_123_199
timestamp 1677580104
transform 1 0 20256 0 -1 95256
box -48 -56 240 834
use sg13g2_tielo  IHP_SRAM_582
timestamp 1680000637
transform 1 0 20064 0 -1 66528
box -48 -56 432 834
use sg13g2_tiehi  IHP_SRAM_583
timestamp 1680000651
transform 1 0 13728 0 -1 60480
box -48 -56 432 834
use sg13g2_buf_1  input1
timestamp 1676381911
transform -1 0 20448 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  input2
timestamp 1676381911
transform -1 0 20064 0 -1 4536
box -48 -56 432 834
use sg13g2_buf_1  input3
timestamp 1676381911
transform -1 0 19680 0 1 4536
box -48 -56 432 834
use sg13g2_buf_1  input4
timestamp 1676381911
transform -1 0 20448 0 1 6048
box -48 -56 432 834
use sg13g2_buf_1  input5
timestamp 1676381911
transform -1 0 20448 0 -1 7560
box -48 -56 432 834
use sg13g2_buf_1  input6
timestamp 1676381911
transform -1 0 19680 0 -1 9072
box -48 -56 432 834
use sg13g2_buf_1  input7
timestamp 1676381911
transform -1 0 20448 0 1 7560
box -48 -56 432 834
use sg13g2_buf_1  input8
timestamp 1676381911
transform -1 0 20064 0 -1 9072
box -48 -56 432 834
use sg13g2_buf_1  input9
timestamp 1676381911
transform -1 0 20448 0 -1 9072
box -48 -56 432 834
use sg13g2_buf_1  input10
timestamp 1676381911
transform -1 0 15840 0 -1 13608
box -48 -56 432 834
use sg13g2_buf_1  input11
timestamp 1676381911
transform -1 0 20448 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  input12
timestamp 1676381911
transform -1 0 17760 0 1 12096
box -48 -56 432 834
use sg13g2_buf_1  input13
timestamp 1676381911
transform -1 0 20448 0 -1 10584
box -48 -56 432 834
use sg13g2_buf_1  input14
timestamp 1676381911
transform -1 0 20448 0 -1 4536
box -48 -56 432 834
use sg13g2_buf_1  input15
timestamp 1676381911
transform -1 0 20064 0 1 10584
box -48 -56 432 834
use sg13g2_buf_1  input16
timestamp 1676381911
transform -1 0 15648 0 -1 15120
box -48 -56 432 834
use sg13g2_buf_1  input17
timestamp 1676381911
transform -1 0 20448 0 1 10584
box -48 -56 432 834
use sg13g2_buf_1  input18
timestamp 1676381911
transform -1 0 20448 0 -1 12096
box -48 -56 432 834
use sg13g2_buf_1  input19
timestamp 1676381911
transform -1 0 20448 0 1 12096
box -48 -56 432 834
use sg13g2_buf_1  input20
timestamp 1676381911
transform -1 0 18624 0 -1 15120
box -48 -56 432 834
use sg13g2_buf_1  input21
timestamp 1676381911
transform -1 0 20448 0 -1 13608
box -48 -56 432 834
use sg13g2_buf_1  input22
timestamp 1676381911
transform -1 0 17472 0 -1 16632
box -48 -56 432 834
use sg13g2_buf_1  input23
timestamp 1676381911
transform -1 0 17856 0 -1 16632
box -48 -56 432 834
use sg13g2_buf_1  input24
timestamp 1676381911
transform -1 0 18240 0 -1 16632
box -48 -56 432 834
use sg13g2_buf_1  input25
timestamp 1676381911
transform -1 0 19296 0 -1 6048
box -48 -56 432 834
use sg13g2_buf_1  input26
timestamp 1676381911
transform 1 0 13728 0 1 19656
box -48 -56 432 834
use sg13g2_buf_1  input27
timestamp 1676381911
transform -1 0 17664 0 1 16632
box -48 -56 432 834
use sg13g2_buf_1  input28
timestamp 1676381911
transform -1 0 20064 0 1 4536
box -48 -56 432 834
use sg13g2_buf_1  input29
timestamp 1676381911
transform -1 0 19680 0 -1 6048
box -48 -56 432 834
use sg13g2_buf_1  input30
timestamp 1676381911
transform -1 0 20448 0 1 4536
box -48 -56 432 834
use sg13g2_buf_1  input31
timestamp 1676381911
transform -1 0 20064 0 -1 6048
box -48 -56 432 834
use sg13g2_buf_1  input32
timestamp 1676381911
transform -1 0 20448 0 -1 6048
box -48 -56 432 834
use sg13g2_buf_1  input33
timestamp 1676381911
transform -1 0 17376 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  input34
timestamp 1676381911
transform 1 0 1152 0 -1 75600
box -48 -56 432 834
use sg13g2_buf_1  input35
timestamp 1676381911
transform 1 0 1536 0 -1 75600
box -48 -56 432 834
use sg13g2_buf_1  input36
timestamp 1676381911
transform 1 0 1920 0 -1 75600
box -48 -56 432 834
use sg13g2_buf_1  input37
timestamp 1676381911
transform 1 0 2784 0 1 74088
box -48 -56 432 834
use sg13g2_buf_1  input38
timestamp 1676381911
transform -1 0 10848 0 -1 72576
box -48 -56 432 834
use sg13g2_buf_1  input39
timestamp 1676381911
transform 1 0 4992 0 -1 77112
box -48 -56 432 834
use sg13g2_buf_1  input40
timestamp 1676381911
transform 1 0 6048 0 1 75600
box -48 -56 432 834
use sg13g2_buf_1  input41
timestamp 1676381911
transform -1 0 5760 0 -1 77112
box -48 -56 432 834
use sg13g2_buf_1  input42
timestamp 1676381911
transform 1 0 1152 0 1 80136
box -48 -56 432 834
use sg13g2_buf_1  input43
timestamp 1676381911
transform 1 0 1152 0 -1 81648
box -48 -56 432 834
use sg13g2_buf_1  input44
timestamp 1676381911
transform 1 0 3840 0 -1 80136
box -48 -56 432 834
use sg13g2_buf_1  input45
timestamp 1676381911
transform 1 0 3264 0 1 80136
box -48 -56 432 834
use sg13g2_buf_1  input46
timestamp 1676381911
transform 1 0 4512 0 1 72576
box -48 -56 432 834
use sg13g2_buf_1  input47
timestamp 1676381911
transform 1 0 2784 0 1 75600
box -48 -56 432 834
use sg13g2_buf_1  input48
timestamp 1676381911
transform 1 0 1152 0 1 77112
box -48 -56 432 834
use sg13g2_buf_1  input49
timestamp 1676381911
transform 1 0 1536 0 1 77112
box -48 -56 432 834
use sg13g2_buf_1  input50
timestamp 1676381911
transform -1 0 9312 0 -1 72576
box -48 -56 432 834
use sg13g2_buf_1  input51
timestamp 1676381911
transform 1 0 1152 0 1 78624
box -48 -56 432 834
use sg13g2_buf_1  input52
timestamp 1676381911
transform 1 0 5664 0 1 75600
box -48 -56 432 834
use sg13g2_buf_1  input53
timestamp 1676381911
transform -1 0 10464 0 -1 72576
box -48 -56 432 834
use sg13g2_buf_1  input54
timestamp 1676381911
transform 1 0 1152 0 1 87696
box -48 -56 432 834
use sg13g2_buf_1  input55
timestamp 1676381911
transform 1 0 9024 0 1 83160
box -48 -56 432 834
use sg13g2_buf_1  input56
timestamp 1676381911
transform 1 0 1152 0 -1 90720
box -48 -56 432 834
use sg13g2_buf_1  input57
timestamp 1676381911
transform 1 0 1152 0 -1 89208
box -48 -56 432 834
use sg13g2_buf_1  input58
timestamp 1676381911
transform 1 0 1536 0 -1 89208
box -48 -56 432 834
use sg13g2_buf_1  input59
timestamp 1676381911
transform 1 0 1920 0 -1 89208
box -48 -56 432 834
use sg13g2_buf_1  input60
timestamp 1676381911
transform 1 0 3936 0 -1 87696
box -48 -56 432 834
use sg13g2_buf_1  input61
timestamp 1676381911
transform 1 0 1152 0 1 89208
box -48 -56 432 834
use sg13g2_buf_1  input62
timestamp 1676381911
transform 1 0 1536 0 1 89208
box -48 -56 432 834
use sg13g2_buf_1  input63
timestamp 1676381911
transform 1 0 2304 0 -1 89208
box -48 -56 432 834
use sg13g2_buf_1  input64
timestamp 1676381911
transform 1 0 1920 0 1 89208
box -48 -56 432 834
use sg13g2_buf_1  input65
timestamp 1676381911
transform 1 0 6432 0 -1 86184
box -48 -56 432 834
use sg13g2_buf_1  input66
timestamp 1676381911
transform 1 0 3648 0 1 80136
box -48 -56 432 834
use sg13g2_buf_1  input67
timestamp 1676381911
transform 1 0 9984 0 -1 80136
box -48 -56 432 834
use sg13g2_buf_1  input68
timestamp 1676381911
transform -1 0 10752 0 -1 80136
box -48 -56 432 834
use sg13g2_buf_1  input69
timestamp 1676381911
transform 1 0 1152 0 -1 87696
box -48 -56 432 834
use sg13g2_buf_1  input70
timestamp 1676381911
transform 1 0 4992 0 -1 84672
box -48 -56 432 834
use sg13g2_buf_1  input71
timestamp 1676381911
transform 1 0 3648 0 -1 86184
box -48 -56 432 834
use sg13g2_buf_1  input72
timestamp 1676381911
transform 1 0 5376 0 -1 84672
box -48 -56 432 834
use sg13g2_buf_1  input73
timestamp 1676381911
transform 1 0 3168 0 -1 81648
box -48 -56 432 834
use sg13g2_buf_1  input74
timestamp 1676381911
transform 1 0 4032 0 1 80136
box -48 -56 432 834
use sg13g2_buf_1  input75
timestamp 1676381911
transform 1 0 3552 0 -1 81648
box -48 -56 432 834
use sg13g2_buf_1  input76
timestamp 1676381911
transform 1 0 1152 0 -1 84672
box -48 -56 432 834
use sg13g2_buf_1  input77
timestamp 1676381911
transform 1 0 1536 0 -1 84672
box -48 -56 432 834
use sg13g2_buf_1  input78
timestamp 1676381911
transform 1 0 1920 0 -1 84672
box -48 -56 432 834
use sg13g2_buf_1  input79
timestamp 1676381911
transform -1 0 11328 0 -1 77112
box -48 -56 432 834
use sg13g2_buf_1  input80
timestamp 1676381911
transform 1 0 1152 0 -1 86184
box -48 -56 432 834
use sg13g2_buf_1  input81
timestamp 1676381911
transform 1 0 4608 0 -1 84672
box -48 -56 432 834
use sg13g2_buf_1  input82
timestamp 1676381911
transform 1 0 1536 0 -1 90720
box -48 -56 432 834
use sg13g2_buf_1  input83
timestamp 1676381911
transform 1 0 3840 0 1 89208
box -48 -56 432 834
use sg13g2_buf_1  input84
timestamp 1676381911
transform 1 0 1152 0 -1 92232
box -48 -56 432 834
use sg13g2_buf_1  input85
timestamp 1676381911
transform 1 0 1536 0 -1 92232
box -48 -56 432 834
use sg13g2_buf_1  input86
timestamp 1676381911
transform 1 0 2304 0 1 90720
box -48 -56 432 834
use sg13g2_buf_1  input87
timestamp 1676381911
transform -1 0 3456 0 -1 90720
box -48 -56 432 834
use sg13g2_buf_1  input88
timestamp 1676381911
transform 1 0 1920 0 -1 92232
box -48 -56 432 834
use sg13g2_buf_1  input89
timestamp 1676381911
transform 1 0 2688 0 1 90720
box -48 -56 432 834
use sg13g2_buf_1  input90
timestamp 1676381911
transform 1 0 3456 0 -1 90720
box -48 -56 432 834
use sg13g2_buf_1  input91
timestamp 1676381911
transform 1 0 4224 0 1 89208
box -48 -56 432 834
use sg13g2_buf_1  input92
timestamp 1676381911
transform 1 0 3840 0 -1 90720
box -48 -56 432 834
use sg13g2_buf_1  input93
timestamp 1676381911
transform 1 0 1920 0 -1 90720
box -48 -56 432 834
use sg13g2_buf_1  input94
timestamp 1676381911
transform 1 0 1152 0 1 92232
box -48 -56 432 834
use sg13g2_buf_1  input95
timestamp 1676381911
transform 1 0 1536 0 1 92232
box -48 -56 432 834
use sg13g2_buf_1  input96
timestamp 1676381911
transform 1 0 2304 0 -1 92232
box -48 -56 432 834
use sg13g2_buf_1  input97
timestamp 1676381911
transform 1 0 1920 0 1 92232
box -48 -56 432 834
use sg13g2_buf_1  input98
timestamp 1676381911
transform 1 0 2688 0 -1 92232
box -48 -56 432 834
use sg13g2_buf_1  input99
timestamp 1676381911
transform 1 0 1152 0 -1 93744
box -48 -56 432 834
use sg13g2_buf_1  input100
timestamp 1676381911
transform 1 0 1536 0 -1 93744
box -48 -56 432 834
use sg13g2_buf_1  input101
timestamp 1676381911
transform 1 0 2304 0 1 92232
box -48 -56 432 834
use sg13g2_buf_1  input102
timestamp 1676381911
transform 1 0 1920 0 -1 93744
box -48 -56 432 834
use sg13g2_buf_1  input103
timestamp 1676381911
transform 1 0 1152 0 1 93744
box -48 -56 432 834
use sg13g2_buf_1  input104
timestamp 1676381911
transform 1 0 2688 0 1 89208
box -48 -56 432 834
use sg13g2_buf_1  input105
timestamp 1676381911
transform 1 0 2304 0 -1 93744
box -48 -56 432 834
use sg13g2_buf_1  input106
timestamp 1676381911
transform 1 0 3072 0 -1 93744
box -48 -56 432 834
use sg13g2_buf_1  input107
timestamp 1676381911
transform 1 0 6528 0 1 86184
box -48 -56 432 834
use sg13g2_buf_1  input108
timestamp 1676381911
transform -1 0 8544 0 1 84672
box -48 -56 432 834
use sg13g2_buf_1  input109
timestamp 1676381911
transform 1 0 1152 0 1 90720
box -48 -56 432 834
use sg13g2_buf_1  input110
timestamp 1676381911
transform 1 0 1536 0 1 90720
box -48 -56 432 834
use sg13g2_buf_1  input111
timestamp 1676381911
transform 1 0 1920 0 1 90720
box -48 -56 432 834
use sg13g2_buf_1  input112
timestamp 1676381911
transform 1 0 2688 0 -1 90720
box -48 -56 432 834
use sg13g2_buf_1  input113
timestamp 1676381911
transform 1 0 3456 0 1 89208
box -48 -56 432 834
use sg13g2_buf_1  input114
timestamp 1676381911
transform 1 0 8160 0 -1 95256
box -48 -56 432 834
use sg13g2_buf_1  input115
timestamp 1676381911
transform 1 0 8928 0 1 93744
box -48 -56 432 834
use sg13g2_buf_1  input116
timestamp 1676381911
transform 1 0 8544 0 -1 95256
box -48 -56 432 834
use sg13g2_buf_1  input117
timestamp 1676381911
transform -1 0 9696 0 1 93744
box -48 -56 432 834
use sg13g2_buf_1  input118
timestamp 1676381911
transform -1 0 10848 0 -1 95256
box -48 -56 432 834
use sg13g2_buf_1  input119
timestamp 1676381911
transform 1 0 10848 0 -1 95256
box -48 -56 432 834
use sg13g2_buf_1  input120
timestamp 1676381911
transform 1 0 11232 0 -1 95256
box -48 -56 432 834
use sg13g2_buf_1  input121
timestamp 1676381911
transform -1 0 12000 0 -1 95256
box -48 -56 432 834
use sg13g2_buf_1  input122
timestamp 1676381911
transform -1 0 12768 0 -1 95256
box -48 -56 432 834
use sg13g2_buf_1  input123
timestamp 1676381911
transform 1 0 12000 0 -1 95256
box -48 -56 432 834
use sg13g2_buf_1  input124
timestamp 1676381911
transform 1 0 12768 0 -1 95256
box -48 -56 432 834
use sg13g2_buf_1  input125
timestamp 1676381911
transform -1 0 13536 0 -1 95256
box -48 -56 432 834
use sg13g2_buf_1  input126
timestamp 1676381911
transform -1 0 9312 0 -1 95256
box -48 -56 432 834
use sg13g2_buf_1  input127
timestamp 1676381911
transform 1 0 9696 0 1 93744
box -48 -56 432 834
use sg13g2_buf_1  input128
timestamp 1676381911
transform -1 0 9696 0 -1 95256
box -48 -56 432 834
use sg13g2_buf_1  input129
timestamp 1676381911
transform -1 0 10464 0 1 93744
box -48 -56 432 834
use sg13g2_buf_1  input130
timestamp 1676381911
transform -1 0 10080 0 -1 95256
box -48 -56 432 834
use sg13g2_buf_1  input131
timestamp 1676381911
transform 1 0 10464 0 1 93744
box -48 -56 432 834
use sg13g2_buf_1  input132
timestamp 1676381911
transform 1 0 10080 0 -1 95256
box -48 -56 432 834
use sg13g2_buf_1  input133
timestamp 1676381911
transform -1 0 11232 0 1 93744
box -48 -56 432 834
use sg13g2_buf_1  input134
timestamp 1676381911
transform -1 0 12960 0 1 93744
box -48 -56 432 834
use sg13g2_buf_1  input135
timestamp 1676381911
transform 1 0 13536 0 -1 95256
box -48 -56 432 834
use sg13g2_buf_1  input136
timestamp 1676381911
transform 1 0 12960 0 1 93744
box -48 -56 432 834
use sg13g2_buf_1  input137
timestamp 1676381911
transform -1 0 14304 0 -1 95256
box -48 -56 432 834
use sg13g2_buf_1  input138
timestamp 1676381911
transform -1 0 13728 0 1 93744
box -48 -56 432 834
use sg13g2_buf_1  input139
timestamp 1676381911
transform 1 0 14304 0 -1 95256
box -48 -56 432 834
use sg13g2_buf_1  input140
timestamp 1676381911
transform 1 0 13728 0 1 93744
box -48 -56 432 834
use sg13g2_buf_1  input141
timestamp 1676381911
transform -1 0 15072 0 -1 95256
box -48 -56 432 834
use sg13g2_buf_1  input142
timestamp 1676381911
transform 1 0 9792 0 -1 19656
box -48 -56 432 834
use sg13g2_buf_1  input143
timestamp 1676381911
transform 1 0 1920 0 1 12096
box -48 -56 432 834
use sg13g2_buf_1  input144
timestamp 1676381911
transform 1 0 1536 0 1 12096
box -48 -56 432 834
use sg13g2_buf_1  input145
timestamp 1676381911
transform 1 0 1152 0 1 12096
box -48 -56 432 834
use sg13g2_buf_1  input146
timestamp 1676381911
transform -1 0 11328 0 1 22680
box -48 -56 432 834
use sg13g2_buf_1  input147
timestamp 1676381911
transform 1 0 5088 0 1 18144
box -48 -56 432 834
use sg13g2_buf_1  input148
timestamp 1676381911
transform 1 0 10560 0 1 22680
box -48 -56 432 834
use sg13g2_buf_1  input149
timestamp 1676381911
transform 1 0 1152 0 -1 16632
box -48 -56 432 834
use sg13g2_buf_1  input150
timestamp 1676381911
transform -1 0 10176 0 -1 24192
box -48 -56 432 834
use sg13g2_buf_1  input151
timestamp 1676381911
transform 1 0 1152 0 -1 18144
box -48 -56 432 834
use sg13g2_buf_1  input152
timestamp 1676381911
transform 1 0 9408 0 1 24192
box -48 -56 432 834
use sg13g2_buf_1  input153
timestamp 1676381911
transform 1 0 1920 0 1 18144
box -48 -56 432 834
use sg13g2_buf_1  input154
timestamp 1676381911
transform -1 0 9792 0 -1 19656
box -48 -56 432 834
use sg13g2_buf_1  input155
timestamp 1676381911
transform 1 0 9024 0 -1 19656
box -48 -56 432 834
use sg13g2_buf_1  input156
timestamp 1676381911
transform 1 0 1152 0 -1 13608
box -48 -56 432 834
use sg13g2_buf_1  input157
timestamp 1676381911
transform -1 0 9024 0 -1 19656
box -48 -56 432 834
use sg13g2_buf_1  input158
timestamp 1676381911
transform 1 0 1920 0 1 13608
box -48 -56 432 834
use sg13g2_buf_1  input159
timestamp 1676381911
transform 1 0 1536 0 1 13608
box -48 -56 432 834
use sg13g2_buf_1  input160
timestamp 1676381911
transform 1 0 1152 0 1 13608
box -48 -56 432 834
use sg13g2_buf_1  input161
timestamp 1676381911
transform -1 0 6048 0 -1 18144
box -48 -56 432 834
use sg13g2_buf_1  input162
timestamp 1676381911
transform 1 0 4704 0 1 25704
box -48 -56 432 834
use sg13g2_buf_1  input163
timestamp 1676381911
transform 1 0 1152 0 1 28728
box -48 -56 432 834
use sg13g2_buf_1  input164
timestamp 1676381911
transform 1 0 5088 0 -1 34776
box -48 -56 432 834
use sg13g2_buf_1  input165
timestamp 1676381911
transform 1 0 3840 0 -1 25704
box -48 -56 432 834
use sg13g2_buf_1  input166
timestamp 1676381911
transform 1 0 3456 0 -1 25704
box -48 -56 432 834
use sg13g2_buf_1  input167
timestamp 1676381911
transform 1 0 1152 0 -1 25704
box -48 -56 432 834
use sg13g2_buf_1  input168
timestamp 1676381911
transform 1 0 8640 0 1 31752
box -48 -56 432 834
use sg13g2_buf_1  input169
timestamp 1676381911
transform 1 0 8256 0 1 31752
box -48 -56 432 834
use sg13g2_buf_1  input170
timestamp 1676381911
transform 1 0 4416 0 1 37800
box -48 -56 432 834
use sg13g2_buf_1  input171
timestamp 1676381911
transform 1 0 1152 0 1 27216
box -48 -56 432 834
use sg13g2_buf_1  input172
timestamp 1676381911
transform 1 0 1920 0 1 28728
box -48 -56 432 834
use sg13g2_buf_1  input173
timestamp 1676381911
transform 1 0 1536 0 1 28728
box -48 -56 432 834
use sg13g2_buf_1  input174
timestamp 1676381911
transform 1 0 1536 0 1 18144
box -48 -56 432 834
use sg13g2_buf_1  input175
timestamp 1676381911
transform 1 0 9696 0 -1 28728
box -48 -56 432 834
use sg13g2_buf_1  input176
timestamp 1676381911
transform 1 0 9312 0 -1 28728
box -48 -56 432 834
use sg13g2_buf_1  input177
timestamp 1676381911
transform 1 0 4896 0 1 24192
box -48 -56 432 834
use sg13g2_buf_1  input178
timestamp 1676381911
transform 1 0 1152 0 -1 22680
box -48 -56 432 834
use sg13g2_buf_1  input179
timestamp 1676381911
transform 1 0 10848 0 1 30240
box -48 -56 432 834
use sg13g2_buf_1  input180
timestamp 1676381911
transform 1 0 1152 0 1 22680
box -48 -56 432 834
use sg13g2_buf_1  input181
timestamp 1676381911
transform 1 0 1152 0 1 18144
box -48 -56 432 834
use sg13g2_buf_1  input182
timestamp 1676381911
transform 1 0 5472 0 -1 22680
box -48 -56 432 834
use sg13g2_buf_1  input183
timestamp 1676381911
transform 1 0 2784 0 1 19656
box -48 -56 432 834
use sg13g2_buf_1  input184
timestamp 1676381911
transform 1 0 3168 0 -1 21168
box -48 -56 432 834
use sg13g2_buf_1  input185
timestamp 1676381911
transform 1 0 10080 0 -1 27216
box -48 -56 432 834
use sg13g2_buf_1  input186
timestamp 1676381911
transform 1 0 2784 0 -1 21168
box -48 -56 432 834
use sg13g2_buf_1  input187
timestamp 1676381911
transform 1 0 4896 0 -1 24192
box -48 -56 432 834
use sg13g2_buf_1  input188
timestamp 1676381911
transform 1 0 1536 0 1 21168
box -48 -56 432 834
use sg13g2_buf_1  input189
timestamp 1676381911
transform 1 0 1152 0 1 21168
box -48 -56 432 834
use sg13g2_buf_1  input190
timestamp 1676381911
transform 1 0 3936 0 1 33264
box -48 -56 432 834
use sg13g2_buf_1  input191
timestamp 1676381911
transform 1 0 2784 0 -1 37800
box -48 -56 432 834
use sg13g2_buf_1  input192
timestamp 1676381911
transform 1 0 1536 0 1 36288
box -48 -56 432 834
use sg13g2_buf_1  input193
timestamp 1676381911
transform 1 0 1152 0 1 36288
box -48 -56 432 834
use sg13g2_buf_1  input194
timestamp 1676381911
transform 1 0 1920 0 -1 39312
box -48 -56 432 834
use sg13g2_buf_1  input195
timestamp 1676381911
transform 1 0 1536 0 -1 39312
box -48 -56 432 834
use sg13g2_buf_1  input196
timestamp 1676381911
transform 1 0 1152 0 -1 39312
box -48 -56 432 834
use sg13g2_buf_1  input197
timestamp 1676381911
transform 1 0 1536 0 1 39312
box -48 -56 432 834
use sg13g2_buf_1  input198
timestamp 1676381911
transform 1 0 1152 0 1 39312
box -48 -56 432 834
use sg13g2_buf_1  input199
timestamp 1676381911
transform 1 0 1920 0 -1 40824
box -48 -56 432 834
use sg13g2_buf_1  input200
timestamp 1676381911
transform 1 0 1536 0 -1 40824
box -48 -56 432 834
use sg13g2_buf_1  input201
timestamp 1676381911
transform 1 0 1152 0 -1 33264
box -48 -56 432 834
use sg13g2_buf_1  input202
timestamp 1676381911
transform 1 0 1152 0 -1 40824
box -48 -56 432 834
use sg13g2_buf_1  input203
timestamp 1676381911
transform 1 0 1920 0 1 42336
box -48 -56 432 834
use sg13g2_buf_1  input204
timestamp 1676381911
transform 1 0 1536 0 1 42336
box -48 -56 432 834
use sg13g2_buf_1  input205
timestamp 1676381911
transform 1 0 1152 0 1 42336
box -48 -56 432 834
use sg13g2_buf_1  input206
timestamp 1676381911
transform 1 0 1536 0 -1 43848
box -48 -56 432 834
use sg13g2_buf_1  input207
timestamp 1676381911
transform 1 0 1152 0 -1 43848
box -48 -56 432 834
use sg13g2_buf_1  input208
timestamp 1676381911
transform 1 0 1536 0 1 43848
box -48 -56 432 834
use sg13g2_buf_1  input209
timestamp 1676381911
transform 1 0 1152 0 1 43848
box -48 -56 432 834
use sg13g2_buf_1  input210
timestamp 1676381911
transform 1 0 1536 0 -1 45360
box -48 -56 432 834
use sg13g2_buf_1  input211
timestamp 1676381911
transform 1 0 1152 0 -1 45360
box -48 -56 432 834
use sg13g2_buf_1  input212
timestamp 1676381911
transform 1 0 1536 0 -1 34776
box -48 -56 432 834
use sg13g2_buf_1  input213
timestamp 1676381911
transform 1 0 1536 0 1 45360
box -48 -56 432 834
use sg13g2_buf_1  input214
timestamp 1676381911
transform 1 0 1152 0 1 45360
box -48 -56 432 834
use sg13g2_buf_1  input215
timestamp 1676381911
transform 1 0 1152 0 -1 34776
box -48 -56 432 834
use sg13g2_buf_1  input216
timestamp 1676381911
transform 1 0 1536 0 1 34776
box -48 -56 432 834
use sg13g2_buf_1  input217
timestamp 1676381911
transform 1 0 1152 0 1 34776
box -48 -56 432 834
use sg13g2_buf_1  input218
timestamp 1676381911
transform 1 0 3552 0 -1 37800
box -48 -56 432 834
use sg13g2_buf_1  input219
timestamp 1676381911
transform 1 0 3168 0 -1 37800
box -48 -56 432 834
use sg13g2_buf_1  input220
timestamp 1676381911
transform 1 0 1536 0 -1 36288
box -48 -56 432 834
use sg13g2_buf_1  input221
timestamp 1676381911
transform 1 0 1152 0 -1 36288
box -48 -56 432 834
use sg13g2_buf_1  input222
timestamp 1676381911
transform -1 0 17760 0 1 1512
box -48 -56 432 834
use sg13g2_buf_1  input223
timestamp 1676381911
transform 1 0 3456 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  input224
timestamp 1676381911
transform 1 0 2688 0 -1 4536
box -48 -56 432 834
use sg13g2_buf_1  input225
timestamp 1676381911
transform 1 0 3072 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  input226
timestamp 1676381911
transform 1 0 1248 0 1 1512
box -48 -56 432 834
use sg13g2_buf_1  input227
timestamp 1676381911
transform 1 0 3552 0 1 1512
box -48 -56 432 834
use sg13g2_buf_1  input228
timestamp 1676381911
transform 1 0 4320 0 -1 3024
box -48 -56 432 834
use sg13g2_buf_1  input229
timestamp 1676381911
transform 1 0 3936 0 1 1512
box -48 -56 432 834
use sg13g2_buf_1  input230
timestamp 1676381911
transform 1 0 4704 0 -1 3024
box -48 -56 432 834
use sg13g2_buf_1  input231
timestamp 1676381911
transform -1 0 4704 0 1 1512
box -48 -56 432 834
use sg13g2_buf_1  input232
timestamp 1676381911
transform 1 0 5088 0 -1 3024
box -48 -56 432 834
use sg13g2_buf_1  input233
timestamp 1676381911
transform 1 0 4704 0 1 1512
box -48 -56 432 834
use sg13g2_buf_1  input234
timestamp 1676381911
transform 1 0 5472 0 -1 3024
box -48 -56 432 834
use sg13g2_buf_1  input235
timestamp 1676381911
transform 1 0 1632 0 1 1512
box -48 -56 432 834
use sg13g2_buf_1  input236
timestamp 1676381911
transform 1 0 2016 0 1 1512
box -48 -56 432 834
use sg13g2_buf_1  input237
timestamp 1676381911
transform 1 0 2400 0 1 1512
box -48 -56 432 834
use sg13g2_buf_1  input238
timestamp 1676381911
transform 1 0 3168 0 -1 3024
box -48 -56 432 834
use sg13g2_buf_1  input239
timestamp 1676381911
transform -1 0 3168 0 1 1512
box -48 -56 432 834
use sg13g2_buf_1  input240
timestamp 1676381911
transform 1 0 3552 0 -1 3024
box -48 -56 432 834
use sg13g2_buf_1  input241
timestamp 1676381911
transform 1 0 3168 0 1 1512
box -48 -56 432 834
use sg13g2_buf_1  input242
timestamp 1676381911
transform 1 0 3936 0 -1 3024
box -48 -56 432 834
use sg13g2_buf_1  input243
timestamp 1676381911
transform 1 0 5088 0 1 1512
box -48 -56 432 834
use sg13g2_buf_1  input244
timestamp 1676381911
transform 1 0 5856 0 -1 3024
box -48 -56 432 834
use sg13g2_buf_1  input245
timestamp 1676381911
transform 1 0 5472 0 1 1512
box -48 -56 432 834
use sg13g2_buf_1  input246
timestamp 1676381911
transform 1 0 5856 0 1 1512
box -48 -56 432 834
use sg13g2_buf_1  input247
timestamp 1676381911
transform 1 0 6240 0 1 1512
box -48 -56 432 834
use sg13g2_buf_1  input248
timestamp 1676381911
transform 1 0 6624 0 1 1512
box -48 -56 432 834
use sg13g2_buf_1  input249
timestamp 1676381911
transform 1 0 7392 0 1 1512
box -48 -56 432 834
use sg13g2_buf_1  input250
timestamp 1676381911
transform -1 0 7392 0 1 1512
box -48 -56 432 834
use sg13g2_buf_1  output251
timestamp 1676381911
transform 1 0 15648 0 -1 19656
box -48 -56 432 834
use sg13g2_buf_1  output252
timestamp 1676381911
transform 1 0 17664 0 1 18144
box -48 -56 432 834
use sg13g2_buf_1  output253
timestamp 1676381911
transform 1 0 19296 0 1 16632
box -48 -56 432 834
use sg13g2_buf_1  output254
timestamp 1676381911
transform 1 0 19680 0 1 16632
box -48 -56 432 834
use sg13g2_buf_1  output255
timestamp 1676381911
transform 1 0 20064 0 1 16632
box -48 -56 432 834
use sg13g2_buf_1  output256
timestamp 1676381911
transform 1 0 20064 0 -1 18144
box -48 -56 432 834
use sg13g2_buf_1  output257
timestamp 1676381911
transform 1 0 20064 0 1 18144
box -48 -56 432 834
use sg13g2_buf_1  output258
timestamp 1676381911
transform 1 0 14880 0 1 24192
box -48 -56 432 834
use sg13g2_buf_1  output259
timestamp 1676381911
transform 1 0 16416 0 -1 24192
box -48 -56 432 834
use sg13g2_buf_1  output260
timestamp 1676381911
transform 1 0 20064 0 -1 21168
box -48 -56 432 834
use sg13g2_buf_1  output261
timestamp 1676381911
transform 1 0 14688 0 1 25704
box -48 -56 432 834
use sg13g2_buf_1  output262
timestamp 1676381911
transform 1 0 17184 0 -1 24192
box -48 -56 432 834
use sg13g2_buf_1  output263
timestamp 1676381911
transform 1 0 15456 0 -1 31752
box -48 -56 432 834
use sg13g2_buf_1  output264
timestamp 1676381911
transform 1 0 15840 0 -1 31752
box -48 -56 432 834
use sg13g2_buf_1  output265
timestamp 1676381911
transform 1 0 16224 0 -1 31752
box -48 -56 432 834
use sg13g2_buf_1  output266
timestamp 1676381911
transform 1 0 18528 0 1 30240
box -48 -56 432 834
use sg13g2_buf_1  output267
timestamp 1676381911
transform 1 0 20064 0 1 28728
box -48 -56 432 834
use sg13g2_buf_1  output268
timestamp 1676381911
transform 1 0 18912 0 1 30240
box -48 -56 432 834
use sg13g2_buf_1  output269
timestamp 1676381911
transform 1 0 19680 0 -1 30240
box -48 -56 432 834
use sg13g2_buf_1  output270
timestamp 1676381911
transform 1 0 19296 0 1 30240
box -48 -56 432 834
use sg13g2_buf_1  output271
timestamp 1676381911
transform 1 0 20064 0 -1 30240
box -48 -56 432 834
use sg13g2_buf_1  output272
timestamp 1676381911
transform 1 0 17856 0 1 31752
box -48 -56 432 834
use sg13g2_buf_1  output273
timestamp 1676381911
transform 1 0 18144 0 1 22680
box -48 -56 432 834
use sg13g2_buf_1  output274
timestamp 1676381911
transform 1 0 19680 0 1 30240
box -48 -56 432 834
use sg13g2_buf_1  output275
timestamp 1676381911
transform 1 0 20064 0 1 30240
box -48 -56 432 834
use sg13g2_buf_1  output276
timestamp 1676381911
transform 1 0 14784 0 -1 36288
box -48 -56 432 834
use sg13g2_buf_1  output277
timestamp 1676381911
transform 1 0 16320 0 -1 34776
box -48 -56 432 834
use sg13g2_buf_1  output278
timestamp 1676381911
transform 1 0 14016 0 -1 39312
box -48 -56 432 834
use sg13g2_buf_1  output279
timestamp 1676381911
transform 1 0 19296 0 -1 34776
box -48 -56 432 834
use sg13g2_buf_1  output280
timestamp 1676381911
transform 1 0 19680 0 -1 34776
box -48 -56 432 834
use sg13g2_buf_1  output281
timestamp 1676381911
transform 1 0 20064 0 -1 34776
box -48 -56 432 834
use sg13g2_buf_1  output282
timestamp 1676381911
transform 1 0 14592 0 -1 40824
box -48 -56 432 834
use sg13g2_buf_1  output283
timestamp 1676381911
transform 1 0 14976 0 -1 40824
box -48 -56 432 834
use sg13g2_buf_1  output284
timestamp 1676381911
transform 1 0 18528 0 -1 24192
box -48 -56 432 834
use sg13g2_buf_1  output285
timestamp 1676381911
transform 1 0 18048 0 1 39312
box -48 -56 432 834
use sg13g2_buf_1  output286
timestamp 1676381911
transform 1 0 18432 0 1 39312
box -48 -56 432 834
use sg13g2_buf_1  output287
timestamp 1676381911
transform 1 0 18912 0 1 24192
box -48 -56 432 834
use sg13g2_buf_1  output288
timestamp 1676381911
transform 1 0 19296 0 1 24192
box -48 -56 432 834
use sg13g2_buf_1  output289
timestamp 1676381911
transform 1 0 19680 0 1 24192
box -48 -56 432 834
use sg13g2_buf_1  output290
timestamp 1676381911
transform 1 0 20064 0 1 24192
box -48 -56 432 834
use sg13g2_buf_1  output291
timestamp 1676381911
transform 1 0 19680 0 -1 25704
box -48 -56 432 834
use sg13g2_buf_1  output292
timestamp 1676381911
transform 1 0 20064 0 -1 25704
box -48 -56 432 834
use sg13g2_buf_1  output293
timestamp 1676381911
transform 1 0 18048 0 -1 40824
box -48 -56 432 834
use sg13g2_buf_1  output294
timestamp 1676381911
transform 1 0 20064 0 1 40824
box -48 -56 432 834
use sg13g2_buf_1  output295
timestamp 1676381911
transform 1 0 20064 0 -1 42336
box -48 -56 432 834
use sg13g2_buf_1  output296
timestamp 1676381911
transform 1 0 20064 0 1 46872
box -48 -56 432 834
use sg13g2_buf_1  output297
timestamp 1676381911
transform 1 0 19680 0 -1 48384
box -48 -56 432 834
use sg13g2_buf_1  output298
timestamp 1676381911
transform 1 0 20064 0 -1 48384
box -48 -56 432 834
use sg13g2_buf_1  output299
timestamp 1676381911
transform 1 0 19296 0 -1 49896
box -48 -56 432 834
use sg13g2_buf_1  output300
timestamp 1676381911
transform 1 0 19680 0 -1 49896
box -48 -56 432 834
use sg13g2_buf_1  output301
timestamp 1676381911
transform 1 0 20064 0 -1 49896
box -48 -56 432 834
use sg13g2_buf_1  output302
timestamp 1676381911
transform 1 0 20064 0 -1 51408
box -48 -56 432 834
use sg13g2_buf_1  output303
timestamp 1676381911
transform 1 0 19680 0 -1 51408
box -48 -56 432 834
use sg13g2_buf_1  output304
timestamp 1676381911
transform 1 0 20064 0 1 51408
box -48 -56 432 834
use sg13g2_buf_1  output305
timestamp 1676381911
transform 1 0 20064 0 -1 52920
box -48 -56 432 834
use sg13g2_buf_1  output306
timestamp 1676381911
transform 1 0 20064 0 1 42336
box -48 -56 432 834
use sg13g2_buf_1  output307
timestamp 1676381911
transform 1 0 19296 0 -1 51408
box -48 -56 432 834
use sg13g2_buf_1  output308
timestamp 1676381911
transform 1 0 20064 0 -1 55944
box -48 -56 432 834
use sg13g2_buf_1  output309
timestamp 1676381911
transform 1 0 19680 0 -1 55944
box -48 -56 432 834
use sg13g2_buf_1  output310
timestamp 1676381911
transform 1 0 20064 0 1 55944
box -48 -56 432 834
use sg13g2_buf_1  output311
timestamp 1676381911
transform 1 0 17568 0 -1 55944
box -48 -56 432 834
use sg13g2_buf_1  output312
timestamp 1676381911
transform 1 0 17664 0 1 55944
box -48 -56 432 834
use sg13g2_buf_1  output313
timestamp 1676381911
transform 1 0 17376 0 -1 54432
box -48 -56 432 834
use sg13g2_buf_1  output314
timestamp 1676381911
transform 1 0 18240 0 -1 60480
box -48 -56 432 834
use sg13g2_buf_1  output315
timestamp 1676381911
transform 1 0 20064 0 1 61992
box -48 -56 432 834
use sg13g2_buf_1  output316
timestamp 1676381911
transform 1 0 20064 0 -1 63504
box -48 -56 432 834
use sg13g2_buf_1  output317
timestamp 1676381911
transform 1 0 20064 0 -1 43848
box -48 -56 432 834
use sg13g2_buf_1  output318
timestamp 1676381911
transform 1 0 20064 0 -1 65016
box -48 -56 432 834
use sg13g2_buf_1  output319
timestamp 1676381911
transform 1 0 14592 0 -1 60480
box -48 -56 432 834
use sg13g2_buf_1  output320
timestamp 1676381911
transform 1 0 19680 0 1 45360
box -48 -56 432 834
use sg13g2_buf_1  output321
timestamp 1676381911
transform 1 0 20064 0 -1 45360
box -48 -56 432 834
use sg13g2_buf_1  output322
timestamp 1676381911
transform 1 0 20064 0 1 45360
box -48 -56 432 834
use sg13g2_buf_1  output323
timestamp 1676381911
transform 1 0 19680 0 -1 46872
box -48 -56 432 834
use sg13g2_buf_1  output324
timestamp 1676381911
transform 1 0 20064 0 -1 46872
box -48 -56 432 834
use sg13g2_buf_1  output325
timestamp 1676381911
transform 1 0 19680 0 1 46872
box -48 -56 432 834
use sg13g2_buf_1  output326
timestamp 1676381911
transform 1 0 17568 0 -1 63504
box -48 -56 432 834
use sg13g2_buf_1  output327
timestamp 1676381911
transform 1 0 14592 0 1 60480
box -48 -56 432 834
use sg13g2_buf_1  output328
timestamp 1676381911
transform 1 0 20064 0 1 68040
box -48 -56 432 834
use sg13g2_buf_1  output329
timestamp 1676381911
transform 1 0 20064 0 1 72576
box -48 -56 432 834
use sg13g2_buf_1  output330
timestamp 1676381911
transform 1 0 17568 0 1 71064
box -48 -56 432 834
use sg13g2_buf_1  output331
timestamp 1676381911
transform 1 0 17184 0 1 71064
box -48 -56 432 834
use sg13g2_buf_1  output332
timestamp 1676381911
transform 1 0 20064 0 1 74088
box -48 -56 432 834
use sg13g2_buf_1  output333
timestamp 1676381911
transform 1 0 13728 0 -1 69552
box -48 -56 432 834
use sg13g2_buf_1  output334
timestamp 1676381911
transform 1 0 18144 0 -1 74088
box -48 -56 432 834
use sg13g2_buf_1  output335
timestamp 1676381911
transform 1 0 20064 0 1 75600
box -48 -56 432 834
use sg13g2_buf_1  output336
timestamp 1676381911
transform 1 0 20064 0 -1 77112
box -48 -56 432 834
use sg13g2_buf_1  output337
timestamp 1676381911
transform 1 0 18432 0 -1 75600
box -48 -56 432 834
use sg13g2_buf_1  output338
timestamp 1676381911
transform 1 0 15552 0 1 72576
box -48 -56 432 834
use sg13g2_buf_1  output339
timestamp 1676381911
transform 1 0 17664 0 -1 66528
box -48 -56 432 834
use sg13g2_buf_1  output340
timestamp 1676381911
transform 1 0 15168 0 1 72576
box -48 -56 432 834
use sg13g2_buf_1  output341
timestamp 1676381911
transform 1 0 14784 0 1 72576
box -48 -56 432 834
use sg13g2_buf_1  output342
timestamp 1676381911
transform 1 0 17760 0 -1 77112
box -48 -56 432 834
use sg13g2_buf_1  output343
timestamp 1676381911
transform 1 0 20064 0 -1 80136
box -48 -56 432 834
use sg13g2_buf_1  output344
timestamp 1676381911
transform 1 0 14400 0 -1 75600
box -48 -56 432 834
use sg13g2_buf_1  output345
timestamp 1676381911
transform 1 0 19680 0 -1 80136
box -48 -56 432 834
use sg13g2_buf_1  output346
timestamp 1676381911
transform 1 0 19296 0 -1 80136
box -48 -56 432 834
use sg13g2_buf_1  output347
timestamp 1676381911
transform 1 0 13632 0 -1 75600
box -48 -56 432 834
use sg13g2_buf_1  output348
timestamp 1676381911
transform 1 0 14976 0 1 77112
box -48 -56 432 834
use sg13g2_buf_1  output349
timestamp 1676381911
transform 1 0 20064 0 -1 83160
box -48 -56 432 834
use sg13g2_buf_1  output350
timestamp 1676381911
transform 1 0 15072 0 1 63504
box -48 -56 432 834
use sg13g2_buf_1  output351
timestamp 1676381911
transform 1 0 16032 0 1 78624
box -48 -56 432 834
use sg13g2_buf_1  output352
timestamp 1676381911
transform 1 0 16608 0 -1 80136
box -48 -56 432 834
use sg13g2_buf_1  output353
timestamp 1676381911
transform 1 0 14688 0 1 63504
box -48 -56 432 834
use sg13g2_buf_1  output354
timestamp 1676381911
transform 1 0 12864 0 -1 63504
box -48 -56 432 834
use sg13g2_buf_1  output355
timestamp 1676381911
transform 1 0 20064 0 1 69552
box -48 -56 432 834
use sg13g2_buf_1  output356
timestamp 1676381911
transform 1 0 14208 0 -1 65016
box -48 -56 432 834
use sg13g2_buf_1  output357
timestamp 1676381911
transform 1 0 19680 0 1 69552
box -48 -56 432 834
use sg13g2_buf_1  output358
timestamp 1676381911
transform 1 0 20064 0 1 71064
box -48 -56 432 834
use sg13g2_buf_1  output359
timestamp 1676381911
transform 1 0 17952 0 -1 71064
box -48 -56 432 834
use sg13g2_buf_1  output360
timestamp 1676381911
transform -1 0 16416 0 -1 95256
box -48 -56 432 834
use sg13g2_buf_1  output361
timestamp 1676381911
transform -1 0 19872 0 -1 95256
box -48 -56 432 834
use sg13g2_buf_1  output362
timestamp 1676381911
transform -1 0 19200 0 1 93744
box -48 -56 432 834
use sg13g2_buf_1  output363
timestamp 1676381911
transform -1 0 20256 0 -1 95256
box -48 -56 432 834
use sg13g2_buf_1  output364
timestamp 1676381911
transform -1 0 19584 0 1 93744
box -48 -56 432 834
use sg13g2_buf_1  output365
timestamp 1676381911
transform -1 0 18912 0 -1 93744
box -48 -56 432 834
use sg13g2_buf_1  output366
timestamp 1676381911
transform 1 0 18144 0 -1 93744
box -48 -56 432 834
use sg13g2_buf_1  output367
timestamp 1676381911
transform -1 0 19296 0 1 92232
box -48 -56 432 834
use sg13g2_buf_1  output368
timestamp 1676381911
transform 1 0 18528 0 1 92232
box -48 -56 432 834
use sg13g2_buf_1  output369
timestamp 1676381911
transform -1 0 19680 0 -1 92232
box -48 -56 432 834
use sg13g2_buf_1  output370
timestamp 1676381911
transform 1 0 17760 0 -1 93744
box -48 -56 432 834
use sg13g2_buf_1  output371
timestamp 1676381911
transform -1 0 16800 0 -1 95256
box -48 -56 432 834
use sg13g2_buf_1  output372
timestamp 1676381911
transform -1 0 17184 0 -1 95256
box -48 -56 432 834
use sg13g2_buf_1  output373
timestamp 1676381911
transform -1 0 17568 0 -1 95256
box -48 -56 432 834
use sg13g2_buf_1  output374
timestamp 1676381911
transform -1 0 17952 0 -1 95256
box -48 -56 432 834
use sg13g2_buf_1  output375
timestamp 1676381911
transform -1 0 18336 0 -1 95256
box -48 -56 432 834
use sg13g2_buf_1  output376
timestamp 1676381911
transform -1 0 18720 0 -1 95256
box -48 -56 432 834
use sg13g2_buf_1  output377
timestamp 1676381911
transform -1 0 19104 0 -1 95256
box -48 -56 432 834
use sg13g2_buf_1  output378
timestamp 1676381911
transform -1 0 19488 0 -1 95256
box -48 -56 432 834
use sg13g2_buf_1  output379
timestamp 1676381911
transform -1 0 18816 0 1 93744
box -48 -56 432 834
use sg13g2_buf_1  output380
timestamp 1676381911
transform -1 0 3072 0 1 92232
box -48 -56 432 834
use sg13g2_buf_1  output381
timestamp 1676381911
transform -1 0 3072 0 -1 93744
box -48 -56 432 834
use sg13g2_buf_1  output382
timestamp 1676381911
transform 1 0 1536 0 1 93744
box -48 -56 432 834
use sg13g2_buf_1  output383
timestamp 1676381911
transform 1 0 1920 0 1 93744
box -48 -56 432 834
use sg13g2_buf_1  output384
timestamp 1676381911
transform 1 0 1248 0 -1 95256
box -48 -56 432 834
use sg13g2_buf_1  output385
timestamp 1676381911
transform 1 0 2304 0 1 93744
box -48 -56 432 834
use sg13g2_buf_1  output386
timestamp 1676381911
transform 1 0 1632 0 -1 95256
box -48 -56 432 834
use sg13g2_buf_1  output387
timestamp 1676381911
transform 1 0 2016 0 -1 95256
box -48 -56 432 834
use sg13g2_buf_1  output388
timestamp 1676381911
transform 1 0 2400 0 -1 95256
box -48 -56 432 834
use sg13g2_buf_1  output389
timestamp 1676381911
transform -1 0 3936 0 1 93744
box -48 -56 432 834
use sg13g2_buf_1  output390
timestamp 1676381911
transform 1 0 2784 0 -1 95256
box -48 -56 432 834
use sg13g2_buf_1  output391
timestamp 1676381911
transform -1 0 4320 0 1 93744
box -48 -56 432 834
use sg13g2_buf_1  output392
timestamp 1676381911
transform 1 0 3168 0 -1 95256
box -48 -56 432 834
use sg13g2_buf_1  output393
timestamp 1676381911
transform -1 0 4704 0 1 93744
box -48 -56 432 834
use sg13g2_buf_1  output394
timestamp 1676381911
transform 1 0 3552 0 -1 95256
box -48 -56 432 834
use sg13g2_buf_1  output395
timestamp 1676381911
transform -1 0 5088 0 1 93744
box -48 -56 432 834
use sg13g2_buf_1  output396
timestamp 1676381911
transform 1 0 3936 0 -1 95256
box -48 -56 432 834
use sg13g2_buf_1  output397
timestamp 1676381911
transform -1 0 5472 0 1 93744
box -48 -56 432 834
use sg13g2_buf_1  output398
timestamp 1676381911
transform 1 0 4320 0 -1 95256
box -48 -56 432 834
use sg13g2_buf_1  output399
timestamp 1676381911
transform -1 0 5856 0 1 93744
box -48 -56 432 834
use sg13g2_buf_1  output400
timestamp 1676381911
transform 1 0 4704 0 -1 95256
box -48 -56 432 834
use sg13g2_buf_1  output401
timestamp 1676381911
transform 1 0 6624 0 -1 95256
box -48 -56 432 834
use sg13g2_buf_1  output402
timestamp 1676381911
transform -1 0 8160 0 1 93744
box -48 -56 432 834
use sg13g2_buf_1  output403
timestamp 1676381911
transform 1 0 7008 0 -1 95256
box -48 -56 432 834
use sg13g2_buf_1  output404
timestamp 1676381911
transform 1 0 7392 0 -1 95256
box -48 -56 432 834
use sg13g2_buf_1  output405
timestamp 1676381911
transform 1 0 7776 0 -1 95256
box -48 -56 432 834
use sg13g2_buf_1  output406
timestamp 1676381911
transform -1 0 8928 0 1 93744
box -48 -56 432 834
use sg13g2_buf_1  output407
timestamp 1676381911
transform -1 0 6240 0 1 93744
box -48 -56 432 834
use sg13g2_buf_1  output408
timestamp 1676381911
transform 1 0 5088 0 -1 95256
box -48 -56 432 834
use sg13g2_buf_1  output409
timestamp 1676381911
transform -1 0 6624 0 1 93744
box -48 -56 432 834
use sg13g2_buf_1  output410
timestamp 1676381911
transform 1 0 5472 0 -1 95256
box -48 -56 432 834
use sg13g2_buf_1  output411
timestamp 1676381911
transform -1 0 7008 0 1 93744
box -48 -56 432 834
use sg13g2_buf_1  output412
timestamp 1676381911
transform 1 0 5856 0 -1 95256
box -48 -56 432 834
use sg13g2_buf_1  output413
timestamp 1676381911
transform -1 0 7392 0 1 93744
box -48 -56 432 834
use sg13g2_buf_1  output414
timestamp 1676381911
transform 1 0 6240 0 -1 95256
box -48 -56 432 834
use sg13g2_buf_1  output415
timestamp 1676381911
transform -1 0 7776 0 1 93744
box -48 -56 432 834
use sg13g2_buf_1  output416
timestamp 1676381911
transform -1 0 16032 0 -1 95256
box -48 -56 432 834
use sg13g2_buf_1  output417
timestamp 1676381911
transform -1 0 1536 0 1 51408
box -48 -56 432 834
use sg13g2_buf_1  output418
timestamp 1676381911
transform -1 0 1920 0 1 51408
box -48 -56 432 834
use sg13g2_buf_1  output419
timestamp 1676381911
transform -1 0 1536 0 1 52920
box -48 -56 432 834
use sg13g2_buf_1  output420
timestamp 1676381911
transform -1 0 3168 0 -1 52920
box -48 -56 432 834
use sg13g2_buf_1  output421
timestamp 1676381911
transform -1 0 1536 0 -1 51408
box -48 -56 432 834
use sg13g2_buf_1  output422
timestamp 1676381911
transform -1 0 1536 0 -1 54432
box -48 -56 432 834
use sg13g2_buf_1  output423
timestamp 1676381911
transform -1 0 1920 0 -1 51408
box -48 -56 432 834
use sg13g2_buf_1  output424
timestamp 1676381911
transform -1 0 1536 0 1 55944
box -48 -56 432 834
use sg13g2_buf_1  output425
timestamp 1676381911
transform -1 0 1536 0 -1 57456
box -48 -56 432 834
use sg13g2_buf_1  output426
timestamp 1676381911
transform -1 0 1920 0 -1 57456
box -48 -56 432 834
use sg13g2_buf_1  output427
timestamp 1676381911
transform -1 0 3744 0 -1 55944
box -48 -56 432 834
use sg13g2_buf_1  output428
timestamp 1676381911
transform -1 0 2688 0 -1 57456
box -48 -56 432 834
use sg13g2_buf_1  output429
timestamp 1676381911
transform -1 0 1536 0 -1 58968
box -48 -56 432 834
use sg13g2_buf_1  output430
timestamp 1676381911
transform -1 0 1920 0 -1 58968
box -48 -56 432 834
use sg13g2_buf_1  output431
timestamp 1676381911
transform -1 0 1536 0 1 58968
box -48 -56 432 834
use sg13g2_buf_1  output432
timestamp 1676381911
transform -1 0 4704 0 -1 57456
box -48 -56 432 834
use sg13g2_buf_1  output433
timestamp 1676381911
transform -1 0 1536 0 -1 60480
box -48 -56 432 834
use sg13g2_buf_1  output434
timestamp 1676381911
transform -1 0 1920 0 -1 60480
box -48 -56 432 834
use sg13g2_buf_1  output435
timestamp 1676381911
transform -1 0 1536 0 -1 61992
box -48 -56 432 834
use sg13g2_buf_1  output436
timestamp 1676381911
transform -1 0 3168 0 1 60480
box -48 -56 432 834
use sg13g2_buf_1  output437
timestamp 1676381911
transform -1 0 3168 0 1 68040
box -48 -56 432 834
use sg13g2_buf_1  output438
timestamp 1676381911
transform -1 0 2688 0 -1 72576
box -48 -56 432 834
use sg13g2_buf_1  output439
timestamp 1676381911
transform -1 0 5088 0 -1 72576
box -48 -56 432 834
use sg13g2_buf_1  output440
timestamp 1676381911
transform -1 0 3552 0 1 68040
box -48 -56 432 834
use sg13g2_buf_1  output441
timestamp 1676381911
transform -1 0 1536 0 -1 71064
box -48 -56 432 834
use sg13g2_buf_1  output442
timestamp 1676381911
transform -1 0 1920 0 -1 71064
box -48 -56 432 834
use sg13g2_buf_1  output443
timestamp 1676381911
transform -1 0 7680 0 -1 66528
box -48 -56 432 834
use sg13g2_buf_1  output444
timestamp 1676381911
transform -1 0 1536 0 1 71064
box -48 -56 432 834
use sg13g2_buf_1  output445
timestamp 1676381911
transform -1 0 1536 0 -1 72576
box -48 -56 432 834
use sg13g2_buf_1  output446
timestamp 1676381911
transform -1 0 1920 0 -1 72576
box -48 -56 432 834
use sg13g2_buf_1  output447
timestamp 1676381911
transform -1 0 2304 0 -1 72576
box -48 -56 432 834
use sg13g2_buf_1  output448
timestamp 1676381911
transform -1 0 3936 0 -1 71064
box -48 -56 432 834
use sg13g2_buf_1  output449
timestamp 1676381911
transform -1 0 6528 0 -1 58968
box -48 -56 432 834
use sg13g2_buf_1  output450
timestamp 1676381911
transform -1 0 2304 0 -1 66528
box -48 -56 432 834
use sg13g2_buf_1  output451
timestamp 1676381911
transform -1 0 1536 0 1 66528
box -48 -56 432 834
use sg13g2_buf_1  output452
timestamp 1676381911
transform -1 0 3840 0 1 65016
box -48 -56 432 834
use sg13g2_buf_1  output453
timestamp 1676381911
transform -1 0 7488 0 -1 63504
box -48 -56 432 834
use sg13g2_buf_1  output454
timestamp 1676381911
transform -1 0 6816 0 1 63504
box -48 -56 432 834
use sg13g2_buf_1  output455
timestamp 1676381911
transform -1 0 7872 0 -1 63504
box -48 -56 432 834
use sg13g2_buf_1  output456
timestamp 1676381911
transform -1 0 1536 0 -1 63504
box -48 -56 432 834
use sg13g2_buf_1  output457
timestamp 1676381911
transform -1 0 3168 0 1 61992
box -48 -56 432 834
use sg13g2_buf_1  output458
timestamp 1676381911
transform -1 0 1536 0 -1 65016
box -48 -56 432 834
use sg13g2_buf_1  output459
timestamp 1676381911
transform -1 0 1920 0 -1 65016
box -48 -56 432 834
use sg13g2_buf_1  output460
timestamp 1676381911
transform -1 0 3648 0 -1 63504
box -48 -56 432 834
use sg13g2_buf_1  output461
timestamp 1676381911
transform -1 0 3456 0 1 63504
box -48 -56 432 834
use sg13g2_buf_1  output462
timestamp 1676381911
transform -1 0 3840 0 1 63504
box -48 -56 432 834
use sg13g2_buf_1  output463
timestamp 1676381911
transform -1 0 1536 0 -1 66528
box -48 -56 432 834
use sg13g2_buf_1  output464
timestamp 1676381911
transform -1 0 1920 0 -1 66528
box -48 -56 432 834
use sg13g2_buf_1  output465
timestamp 1676381911
transform 1 0 17856 0 -1 81648
box -48 -56 432 834
use sg13g2_buf_1  output466
timestamp 1676381911
transform 1 0 17376 0 -1 86184
box -48 -56 432 834
use sg13g2_buf_1  output467
timestamp 1676381911
transform 1 0 14016 0 -1 83160
box -48 -56 432 834
use sg13g2_buf_1  output468
timestamp 1676381911
transform 1 0 20064 0 -1 89208
box -48 -56 432 834
use sg13g2_buf_1  output469
timestamp 1676381911
transform 1 0 19680 0 -1 89208
box -48 -56 432 834
use sg13g2_buf_1  output470
timestamp 1676381911
transform 1 0 20064 0 1 89208
box -48 -56 432 834
use sg13g2_buf_1  output471
timestamp 1676381911
transform 1 0 19296 0 -1 89208
box -48 -56 432 834
use sg13g2_buf_1  output472
timestamp 1676381911
transform 1 0 18144 0 1 87696
box -48 -56 432 834
use sg13g2_buf_1  output473
timestamp 1676381911
transform 1 0 19680 0 1 89208
box -48 -56 432 834
use sg13g2_buf_1  output474
timestamp 1676381911
transform 1 0 18912 0 -1 89208
box -48 -56 432 834
use sg13g2_buf_1  output475
timestamp 1676381911
transform 1 0 20064 0 -1 90720
box -48 -56 432 834
use sg13g2_buf_1  output476
timestamp 1676381911
transform 1 0 20064 0 1 83160
box -48 -56 432 834
use sg13g2_buf_1  output477
timestamp 1676381911
transform 1 0 19296 0 1 89208
box -48 -56 432 834
use sg13g2_buf_1  output478
timestamp 1676381911
transform 1 0 18528 0 -1 89208
box -48 -56 432 834
use sg13g2_buf_1  output479
timestamp 1676381911
transform 1 0 19680 0 -1 90720
box -48 -56 432 834
use sg13g2_buf_1  output480
timestamp 1676381911
transform 1 0 18912 0 1 89208
box -48 -56 432 834
use sg13g2_buf_1  output481
timestamp 1676381911
transform 1 0 20064 0 1 90720
box -48 -56 432 834
use sg13g2_buf_1  output482
timestamp 1676381911
transform 1 0 19296 0 -1 90720
box -48 -56 432 834
use sg13g2_buf_1  output483
timestamp 1676381911
transform 1 0 19680 0 1 90720
box -48 -56 432 834
use sg13g2_buf_1  output484
timestamp 1676381911
transform 1 0 20064 0 -1 92232
box -48 -56 432 834
use sg13g2_buf_1  output485
timestamp 1676381911
transform 1 0 19680 0 -1 92232
box -48 -56 432 834
use sg13g2_buf_1  output486
timestamp 1676381911
transform 1 0 20064 0 1 92232
box -48 -56 432 834
use sg13g2_buf_1  output487
timestamp 1676381911
transform 1 0 20064 0 -1 84672
box -48 -56 432 834
use sg13g2_buf_1  output488
timestamp 1676381911
transform 1 0 19680 0 1 92232
box -48 -56 432 834
use sg13g2_buf_1  output489
timestamp 1676381911
transform 1 0 20064 0 -1 93744
box -48 -56 432 834
use sg13g2_buf_1  output490
timestamp 1676381911
transform 1 0 19680 0 -1 84672
box -48 -56 432 834
use sg13g2_buf_1  output491
timestamp 1676381911
transform 1 0 20064 0 1 86184
box -48 -56 432 834
use sg13g2_buf_1  output492
timestamp 1676381911
transform 1 0 11712 0 -1 80136
box -48 -56 432 834
use sg13g2_buf_1  output493
timestamp 1676381911
transform 1 0 19680 0 1 86184
box -48 -56 432 834
use sg13g2_buf_1  output494
timestamp 1676381911
transform 1 0 20064 0 -1 87696
box -48 -56 432 834
use sg13g2_buf_1  output495
timestamp 1676381911
transform 1 0 19680 0 -1 87696
box -48 -56 432 834
use sg13g2_buf_1  output496
timestamp 1676381911
transform 1 0 17760 0 -1 86184
box -48 -56 432 834
use sg13g2_buf_1  output497
timestamp 1676381911
transform 1 0 8160 0 1 1512
box -48 -56 432 834
use sg13g2_buf_1  output498
timestamp 1676381911
transform -1 0 9312 0 -1 3024
box -48 -56 432 834
use sg13g2_buf_1  output499
timestamp 1676381911
transform 1 0 8544 0 1 1512
box -48 -56 432 834
use sg13g2_buf_1  output500
timestamp 1676381911
transform -1 0 9696 0 -1 3024
box -48 -56 432 834
use sg13g2_buf_1  output501
timestamp 1676381911
transform 1 0 8928 0 1 1512
box -48 -56 432 834
use sg13g2_buf_1  output502
timestamp 1676381911
transform -1 0 10080 0 -1 3024
box -48 -56 432 834
use sg13g2_buf_1  output503
timestamp 1676381911
transform 1 0 9312 0 1 1512
box -48 -56 432 834
use sg13g2_buf_1  output504
timestamp 1676381911
transform -1 0 10464 0 -1 3024
box -48 -56 432 834
use sg13g2_buf_1  output505
timestamp 1676381911
transform 1 0 9696 0 1 1512
box -48 -56 432 834
use sg13g2_buf_1  output506
timestamp 1676381911
transform -1 0 10848 0 -1 3024
box -48 -56 432 834
use sg13g2_buf_1  output507
timestamp 1676381911
transform 1 0 10080 0 1 1512
box -48 -56 432 834
use sg13g2_buf_1  output508
timestamp 1676381911
transform -1 0 11232 0 -1 3024
box -48 -56 432 834
use sg13g2_buf_1  output509
timestamp 1676381911
transform 1 0 10464 0 1 1512
box -48 -56 432 834
use sg13g2_buf_1  output510
timestamp 1676381911
transform 1 0 10848 0 1 1512
box -48 -56 432 834
use sg13g2_buf_1  output511
timestamp 1676381911
transform -1 0 11616 0 1 1512
box -48 -56 432 834
use sg13g2_buf_1  output512
timestamp 1676381911
transform -1 0 12000 0 1 1512
box -48 -56 432 834
use sg13g2_buf_1  output513
timestamp 1676381911
transform -1 0 12768 0 1 1512
box -48 -56 432 834
use sg13g2_buf_1  output514
timestamp 1676381911
transform -1 0 12384 0 1 1512
box -48 -56 432 834
use sg13g2_buf_1  output515
timestamp 1676381911
transform -1 0 13152 0 1 1512
box -48 -56 432 834
use sg13g2_buf_1  output516
timestamp 1676381911
transform -1 0 13536 0 1 1512
box -48 -56 432 834
use sg13g2_buf_1  output517
timestamp 1676381911
transform -1 0 12960 0 -1 3024
box -48 -56 432 834
use sg13g2_buf_1  output518
timestamp 1676381911
transform -1 0 14880 0 -1 3024
box -48 -56 432 834
use sg13g2_buf_1  output519
timestamp 1676381911
transform -1 0 15840 0 1 1512
box -48 -56 432 834
use sg13g2_buf_1  output520
timestamp 1676381911
transform -1 0 15264 0 -1 3024
box -48 -56 432 834
use sg13g2_buf_1  output521
timestamp 1676381911
transform -1 0 16224 0 1 1512
box -48 -56 432 834
use sg13g2_buf_1  output522
timestamp 1676381911
transform -1 0 15648 0 -1 3024
box -48 -56 432 834
use sg13g2_buf_1  output523
timestamp 1676381911
transform -1 0 16608 0 1 1512
box -48 -56 432 834
use sg13g2_buf_1  output524
timestamp 1676381911
transform -1 0 13920 0 1 1512
box -48 -56 432 834
use sg13g2_buf_1  output525
timestamp 1676381911
transform -1 0 13344 0 -1 3024
box -48 -56 432 834
use sg13g2_buf_1  output526
timestamp 1676381911
transform -1 0 14304 0 1 1512
box -48 -56 432 834
use sg13g2_buf_1  output527
timestamp 1676381911
transform -1 0 13728 0 -1 3024
box -48 -56 432 834
use sg13g2_buf_1  output528
timestamp 1676381911
transform -1 0 14688 0 1 1512
box -48 -56 432 834
use sg13g2_buf_1  output529
timestamp 1676381911
transform -1 0 14112 0 -1 3024
box -48 -56 432 834
use sg13g2_buf_1  output530
timestamp 1676381911
transform -1 0 15072 0 1 1512
box -48 -56 432 834
use sg13g2_buf_1  output531
timestamp 1676381911
transform -1 0 14496 0 -1 3024
box -48 -56 432 834
use sg13g2_buf_1  output532
timestamp 1676381911
transform -1 0 15456 0 1 1512
box -48 -56 432 834
use sg13g2_buf_1  output533
timestamp 1676381911
transform -1 0 3072 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  output534
timestamp 1676381911
transform -1 0 1536 0 -1 3024
box -48 -56 432 834
use sg13g2_buf_1  output535
timestamp 1676381911
transform -1 0 2304 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  output536
timestamp 1676381911
transform -1 0 2688 0 -1 4536
box -48 -56 432 834
use sg13g2_buf_1  output537
timestamp 1676381911
transform -1 0 1920 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  output538
timestamp 1676381911
transform -1 0 1536 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  output539
timestamp 1676381911
transform -1 0 3072 0 1 4536
box -48 -56 432 834
use sg13g2_buf_1  output540
timestamp 1676381911
transform -1 0 2304 0 -1 4536
box -48 -56 432 834
use sg13g2_buf_1  output541
timestamp 1676381911
transform -1 0 3456 0 -1 6048
box -48 -56 432 834
use sg13g2_buf_1  output542
timestamp 1676381911
transform -1 0 2688 0 1 4536
box -48 -56 432 834
use sg13g2_buf_1  output543
timestamp 1676381911
transform -1 0 1920 0 -1 4536
box -48 -56 432 834
use sg13g2_buf_1  output544
timestamp 1676381911
transform -1 0 1536 0 -1 4536
box -48 -56 432 834
use sg13g2_buf_1  output545
timestamp 1676381911
transform -1 0 5088 0 -1 7560
box -48 -56 432 834
use sg13g2_buf_1  output546
timestamp 1676381911
transform -1 0 4704 0 -1 7560
box -48 -56 432 834
use sg13g2_buf_1  output547
timestamp 1676381911
transform -1 0 2304 0 1 4536
box -48 -56 432 834
use sg13g2_buf_1  output548
timestamp 1676381911
transform -1 0 3552 0 1 6048
box -48 -56 432 834
use sg13g2_buf_1  output549
timestamp 1676381911
transform -1 0 2688 0 -1 6048
box -48 -56 432 834
use sg13g2_buf_1  output550
timestamp 1676381911
transform -1 0 1920 0 1 4536
box -48 -56 432 834
use sg13g2_buf_1  output551
timestamp 1676381911
transform -1 0 1536 0 1 4536
box -48 -56 432 834
use sg13g2_buf_1  output552
timestamp 1676381911
transform -1 0 4320 0 -1 7560
box -48 -56 432 834
use sg13g2_buf_1  output553
timestamp 1676381911
transform -1 0 2592 0 -1 10584
box -48 -56 432 834
use sg13g2_buf_1  output554
timestamp 1676381911
transform -1 0 1536 0 -1 12096
box -48 -56 432 834
use sg13g2_buf_1  output555
timestamp 1676381911
transform -1 0 10560 0 -1 19656
box -48 -56 432 834
use sg13g2_buf_1  output556
timestamp 1676381911
transform -1 0 1536 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  output557
timestamp 1676381911
transform -1 0 4128 0 -1 12096
box -48 -56 432 834
use sg13g2_buf_1  output558
timestamp 1676381911
transform -1 0 3168 0 1 10584
box -48 -56 432 834
use sg13g2_buf_1  output559
timestamp 1676381911
transform -1 0 1536 0 -1 10584
box -48 -56 432 834
use sg13g2_buf_1  output560
timestamp 1676381911
transform -1 0 8640 0 1 16632
box -48 -56 432 834
use sg13g2_buf_1  output561
timestamp 1676381911
transform -1 0 7008 0 1 15120
box -48 -56 432 834
use sg13g2_buf_1  output562
timestamp 1676381911
transform -1 0 5184 0 1 13608
box -48 -56 432 834
use sg13g2_buf_1  output563
timestamp 1676381911
transform -1 0 3936 0 -1 13608
box -48 -56 432 834
use sg13g2_buf_1  output564
timestamp 1676381911
transform -1 0 1920 0 -1 12096
box -48 -56 432 834
use sg13g2_buf_1  output565
timestamp 1676381911
transform -1 0 2304 0 -1 6048
box -48 -56 432 834
use sg13g2_buf_1  output566
timestamp 1676381911
transform -1 0 7968 0 1 12096
box -48 -56 432 834
use sg13g2_buf_1  output567
timestamp 1676381911
transform -1 0 8448 0 -1 13608
box -48 -56 432 834
use sg13g2_buf_1  output568
timestamp 1676381911
transform -1 0 3168 0 -1 9072
box -48 -56 432 834
use sg13g2_buf_1  output569
timestamp 1676381911
transform -1 0 3840 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  output570
timestamp 1676381911
transform -1 0 8256 0 -1 15120
box -48 -56 432 834
use sg13g2_buf_1  output571
timestamp 1676381911
transform -1 0 3936 0 1 10584
box -48 -56 432 834
use sg13g2_buf_1  output572
timestamp 1676381911
transform -1 0 2688 0 1 6048
box -48 -56 432 834
use sg13g2_buf_1  output573
timestamp 1676381911
transform -1 0 1920 0 -1 6048
box -48 -56 432 834
use sg13g2_buf_1  output574
timestamp 1676381911
transform -1 0 1536 0 -1 6048
box -48 -56 432 834
use sg13g2_buf_1  output575
timestamp 1676381911
transform -1 0 1920 0 1 6048
box -48 -56 432 834
use sg13g2_buf_1  output576
timestamp 1676381911
transform -1 0 1536 0 1 6048
box -48 -56 432 834
use sg13g2_buf_1  output577
timestamp 1676381911
transform -1 0 2304 0 -1 7560
box -48 -56 432 834
use sg13g2_buf_1  output578
timestamp 1676381911
transform -1 0 1920 0 -1 7560
box -48 -56 432 834
use sg13g2_buf_1  output579
timestamp 1676381911
transform -1 0 1536 0 -1 7560
box -48 -56 432 834
use sg13g2_buf_1  output580
timestamp 1676381911
transform -1 0 8832 0 -1 13608
box -48 -56 432 834
use sg13g2_buf_1  output581
timestamp 1676381911
transform 1 0 12096 0 1 60480
box -48 -56 432 834
<< labels >>
flabel metal2 s 21510 20540 21600 20620 0 FreeSans 320 0 0 0 ADDR_SRAM0
port 0 nsew signal output
flabel metal2 s 21510 21044 21600 21124 0 FreeSans 320 0 0 0 ADDR_SRAM1
port 1 nsew signal output
flabel metal2 s 21510 21548 21600 21628 0 FreeSans 320 0 0 0 ADDR_SRAM2
port 2 nsew signal output
flabel metal2 s 21510 22052 21600 22132 0 FreeSans 320 0 0 0 ADDR_SRAM3
port 3 nsew signal output
flabel metal2 s 21510 22556 21600 22636 0 FreeSans 320 0 0 0 ADDR_SRAM4
port 4 nsew signal output
flabel metal2 s 21510 23060 21600 23140 0 FreeSans 320 0 0 0 ADDR_SRAM5
port 5 nsew signal output
flabel metal2 s 21510 23564 21600 23644 0 FreeSans 320 0 0 0 ADDR_SRAM6
port 6 nsew signal output
flabel metal2 s 21510 24068 21600 24148 0 FreeSans 320 0 0 0 ADDR_SRAM7
port 7 nsew signal output
flabel metal2 s 21510 24572 21600 24652 0 FreeSans 320 0 0 0 ADDR_SRAM8
port 8 nsew signal output
flabel metal2 s 21510 25076 21600 25156 0 FreeSans 320 0 0 0 ADDR_SRAM9
port 9 nsew signal output
flabel metal2 s 21510 25580 21600 25660 0 FreeSans 320 0 0 0 BM_SRAM0
port 10 nsew signal output
flabel metal2 s 21510 26084 21600 26164 0 FreeSans 320 0 0 0 BM_SRAM1
port 11 nsew signal output
flabel metal2 s 21510 30620 21600 30700 0 FreeSans 320 0 0 0 BM_SRAM10
port 12 nsew signal output
flabel metal2 s 21510 31124 21600 31204 0 FreeSans 320 0 0 0 BM_SRAM11
port 13 nsew signal output
flabel metal2 s 21510 31628 21600 31708 0 FreeSans 320 0 0 0 BM_SRAM12
port 14 nsew signal output
flabel metal2 s 21510 32132 21600 32212 0 FreeSans 320 0 0 0 BM_SRAM13
port 15 nsew signal output
flabel metal2 s 21510 32636 21600 32716 0 FreeSans 320 0 0 0 BM_SRAM14
port 16 nsew signal output
flabel metal2 s 21510 33140 21600 33220 0 FreeSans 320 0 0 0 BM_SRAM15
port 17 nsew signal output
flabel metal2 s 21510 33644 21600 33724 0 FreeSans 320 0 0 0 BM_SRAM16
port 18 nsew signal output
flabel metal2 s 21510 34148 21600 34228 0 FreeSans 320 0 0 0 BM_SRAM17
port 19 nsew signal output
flabel metal2 s 21510 34652 21600 34732 0 FreeSans 320 0 0 0 BM_SRAM18
port 20 nsew signal output
flabel metal2 s 21510 35156 21600 35236 0 FreeSans 320 0 0 0 BM_SRAM19
port 21 nsew signal output
flabel metal2 s 21510 26588 21600 26668 0 FreeSans 320 0 0 0 BM_SRAM2
port 22 nsew signal output
flabel metal2 s 21510 35660 21600 35740 0 FreeSans 320 0 0 0 BM_SRAM20
port 23 nsew signal output
flabel metal2 s 21510 36164 21600 36244 0 FreeSans 320 0 0 0 BM_SRAM21
port 24 nsew signal output
flabel metal2 s 21510 36668 21600 36748 0 FreeSans 320 0 0 0 BM_SRAM22
port 25 nsew signal output
flabel metal2 s 21510 37172 21600 37252 0 FreeSans 320 0 0 0 BM_SRAM23
port 26 nsew signal output
flabel metal2 s 21510 37676 21600 37756 0 FreeSans 320 0 0 0 BM_SRAM24
port 27 nsew signal output
flabel metal2 s 21510 38180 21600 38260 0 FreeSans 320 0 0 0 BM_SRAM25
port 28 nsew signal output
flabel metal2 s 21510 38684 21600 38764 0 FreeSans 320 0 0 0 BM_SRAM26
port 29 nsew signal output
flabel metal2 s 21510 39188 21600 39268 0 FreeSans 320 0 0 0 BM_SRAM27
port 30 nsew signal output
flabel metal2 s 21510 39692 21600 39772 0 FreeSans 320 0 0 0 BM_SRAM28
port 31 nsew signal output
flabel metal2 s 21510 40196 21600 40276 0 FreeSans 320 0 0 0 BM_SRAM29
port 32 nsew signal output
flabel metal2 s 21510 27092 21600 27172 0 FreeSans 320 0 0 0 BM_SRAM3
port 33 nsew signal output
flabel metal2 s 21510 40700 21600 40780 0 FreeSans 320 0 0 0 BM_SRAM30
port 34 nsew signal output
flabel metal2 s 21510 41204 21600 41284 0 FreeSans 320 0 0 0 BM_SRAM31
port 35 nsew signal output
flabel metal2 s 21510 27596 21600 27676 0 FreeSans 320 0 0 0 BM_SRAM4
port 36 nsew signal output
flabel metal2 s 21510 28100 21600 28180 0 FreeSans 320 0 0 0 BM_SRAM5
port 37 nsew signal output
flabel metal2 s 21510 28604 21600 28684 0 FreeSans 320 0 0 0 BM_SRAM6
port 38 nsew signal output
flabel metal2 s 21510 29108 21600 29188 0 FreeSans 320 0 0 0 BM_SRAM7
port 39 nsew signal output
flabel metal2 s 21510 29612 21600 29692 0 FreeSans 320 0 0 0 BM_SRAM8
port 40 nsew signal output
flabel metal2 s 21510 30116 21600 30196 0 FreeSans 320 0 0 0 BM_SRAM9
port 41 nsew signal output
flabel metal2 s 21510 41708 21600 41788 0 FreeSans 320 0 0 0 CLK_SRAM
port 42 nsew signal output
flabel metal2 s 21510 3908 21600 3988 0 FreeSans 320 0 0 0 CONFIGURED_top
port 43 nsew signal input
flabel metal2 s 21510 42212 21600 42292 0 FreeSans 320 0 0 0 DIN_SRAM0
port 44 nsew signal output
flabel metal2 s 21510 42716 21600 42796 0 FreeSans 320 0 0 0 DIN_SRAM1
port 45 nsew signal output
flabel metal2 s 21510 47252 21600 47332 0 FreeSans 320 0 0 0 DIN_SRAM10
port 46 nsew signal output
flabel metal2 s 21510 47756 21600 47836 0 FreeSans 320 0 0 0 DIN_SRAM11
port 47 nsew signal output
flabel metal2 s 21510 48260 21600 48340 0 FreeSans 320 0 0 0 DIN_SRAM12
port 48 nsew signal output
flabel metal2 s 21510 48764 21600 48844 0 FreeSans 320 0 0 0 DIN_SRAM13
port 49 nsew signal output
flabel metal2 s 21510 49268 21600 49348 0 FreeSans 320 0 0 0 DIN_SRAM14
port 50 nsew signal output
flabel metal2 s 21510 49772 21600 49852 0 FreeSans 320 0 0 0 DIN_SRAM15
port 51 nsew signal output
flabel metal2 s 21510 50276 21600 50356 0 FreeSans 320 0 0 0 DIN_SRAM16
port 52 nsew signal output
flabel metal2 s 21510 50780 21600 50860 0 FreeSans 320 0 0 0 DIN_SRAM17
port 53 nsew signal output
flabel metal2 s 21510 51284 21600 51364 0 FreeSans 320 0 0 0 DIN_SRAM18
port 54 nsew signal output
flabel metal2 s 21510 51788 21600 51868 0 FreeSans 320 0 0 0 DIN_SRAM19
port 55 nsew signal output
flabel metal2 s 21510 43220 21600 43300 0 FreeSans 320 0 0 0 DIN_SRAM2
port 56 nsew signal output
flabel metal2 s 21510 52292 21600 52372 0 FreeSans 320 0 0 0 DIN_SRAM20
port 57 nsew signal output
flabel metal2 s 21510 52796 21600 52876 0 FreeSans 320 0 0 0 DIN_SRAM21
port 58 nsew signal output
flabel metal2 s 21510 53300 21600 53380 0 FreeSans 320 0 0 0 DIN_SRAM22
port 59 nsew signal output
flabel metal2 s 21510 53804 21600 53884 0 FreeSans 320 0 0 0 DIN_SRAM23
port 60 nsew signal output
flabel metal2 s 21510 54308 21600 54388 0 FreeSans 320 0 0 0 DIN_SRAM24
port 61 nsew signal output
flabel metal2 s 21510 54812 21600 54892 0 FreeSans 320 0 0 0 DIN_SRAM25
port 62 nsew signal output
flabel metal2 s 21510 55316 21600 55396 0 FreeSans 320 0 0 0 DIN_SRAM26
port 63 nsew signal output
flabel metal2 s 21510 55820 21600 55900 0 FreeSans 320 0 0 0 DIN_SRAM27
port 64 nsew signal output
flabel metal2 s 21510 56324 21600 56404 0 FreeSans 320 0 0 0 DIN_SRAM28
port 65 nsew signal output
flabel metal2 s 21510 56828 21600 56908 0 FreeSans 320 0 0 0 DIN_SRAM29
port 66 nsew signal output
flabel metal2 s 21510 43724 21600 43804 0 FreeSans 320 0 0 0 DIN_SRAM3
port 67 nsew signal output
flabel metal2 s 21510 57332 21600 57412 0 FreeSans 320 0 0 0 DIN_SRAM30
port 68 nsew signal output
flabel metal2 s 21510 57836 21600 57916 0 FreeSans 320 0 0 0 DIN_SRAM31
port 69 nsew signal output
flabel metal2 s 21510 44228 21600 44308 0 FreeSans 320 0 0 0 DIN_SRAM4
port 70 nsew signal output
flabel metal2 s 21510 44732 21600 44812 0 FreeSans 320 0 0 0 DIN_SRAM5
port 71 nsew signal output
flabel metal2 s 21510 45236 21600 45316 0 FreeSans 320 0 0 0 DIN_SRAM6
port 72 nsew signal output
flabel metal2 s 21510 45740 21600 45820 0 FreeSans 320 0 0 0 DIN_SRAM7
port 73 nsew signal output
flabel metal2 s 21510 46244 21600 46324 0 FreeSans 320 0 0 0 DIN_SRAM8
port 74 nsew signal output
flabel metal2 s 21510 46748 21600 46828 0 FreeSans 320 0 0 0 DIN_SRAM9
port 75 nsew signal output
flabel metal2 s 21510 4412 21600 4492 0 FreeSans 320 0 0 0 DOUT_SRAM0
port 76 nsew signal input
flabel metal2 s 21510 4916 21600 4996 0 FreeSans 320 0 0 0 DOUT_SRAM1
port 77 nsew signal input
flabel metal2 s 21510 9452 21600 9532 0 FreeSans 320 0 0 0 DOUT_SRAM10
port 78 nsew signal input
flabel metal2 s 21510 9956 21600 10036 0 FreeSans 320 0 0 0 DOUT_SRAM11
port 79 nsew signal input
flabel metal2 s 21510 10460 21600 10540 0 FreeSans 320 0 0 0 DOUT_SRAM12
port 80 nsew signal input
flabel metal2 s 21510 10964 21600 11044 0 FreeSans 320 0 0 0 DOUT_SRAM13
port 81 nsew signal input
flabel metal2 s 21510 11468 21600 11548 0 FreeSans 320 0 0 0 DOUT_SRAM14
port 82 nsew signal input
flabel metal2 s 21510 11972 21600 12052 0 FreeSans 320 0 0 0 DOUT_SRAM15
port 83 nsew signal input
flabel metal2 s 21510 12476 21600 12556 0 FreeSans 320 0 0 0 DOUT_SRAM16
port 84 nsew signal input
flabel metal2 s 21510 12980 21600 13060 0 FreeSans 320 0 0 0 DOUT_SRAM17
port 85 nsew signal input
flabel metal2 s 21510 13484 21600 13564 0 FreeSans 320 0 0 0 DOUT_SRAM18
port 86 nsew signal input
flabel metal2 s 21510 13988 21600 14068 0 FreeSans 320 0 0 0 DOUT_SRAM19
port 87 nsew signal input
flabel metal2 s 21510 5420 21600 5500 0 FreeSans 320 0 0 0 DOUT_SRAM2
port 88 nsew signal input
flabel metal2 s 21510 14492 21600 14572 0 FreeSans 320 0 0 0 DOUT_SRAM20
port 89 nsew signal input
flabel metal2 s 21510 14996 21600 15076 0 FreeSans 320 0 0 0 DOUT_SRAM21
port 90 nsew signal input
flabel metal2 s 21510 15500 21600 15580 0 FreeSans 320 0 0 0 DOUT_SRAM22
port 91 nsew signal input
flabel metal2 s 21510 16004 21600 16084 0 FreeSans 320 0 0 0 DOUT_SRAM23
port 92 nsew signal input
flabel metal2 s 21510 16508 21600 16588 0 FreeSans 320 0 0 0 DOUT_SRAM24
port 93 nsew signal input
flabel metal2 s 21510 17012 21600 17092 0 FreeSans 320 0 0 0 DOUT_SRAM25
port 94 nsew signal input
flabel metal2 s 21510 17516 21600 17596 0 FreeSans 320 0 0 0 DOUT_SRAM26
port 95 nsew signal input
flabel metal2 s 21510 18020 21600 18100 0 FreeSans 320 0 0 0 DOUT_SRAM27
port 96 nsew signal input
flabel metal2 s 21510 18524 21600 18604 0 FreeSans 320 0 0 0 DOUT_SRAM28
port 97 nsew signal input
flabel metal2 s 21510 19028 21600 19108 0 FreeSans 320 0 0 0 DOUT_SRAM29
port 98 nsew signal input
flabel metal2 s 21510 5924 21600 6004 0 FreeSans 320 0 0 0 DOUT_SRAM3
port 99 nsew signal input
flabel metal2 s 21510 19532 21600 19612 0 FreeSans 320 0 0 0 DOUT_SRAM30
port 100 nsew signal input
flabel metal2 s 21510 20036 21600 20116 0 FreeSans 320 0 0 0 DOUT_SRAM31
port 101 nsew signal input
flabel metal2 s 21510 6428 21600 6508 0 FreeSans 320 0 0 0 DOUT_SRAM4
port 102 nsew signal input
flabel metal2 s 21510 6932 21600 7012 0 FreeSans 320 0 0 0 DOUT_SRAM5
port 103 nsew signal input
flabel metal2 s 21510 7436 21600 7516 0 FreeSans 320 0 0 0 DOUT_SRAM6
port 104 nsew signal input
flabel metal2 s 21510 7940 21600 8020 0 FreeSans 320 0 0 0 DOUT_SRAM7
port 105 nsew signal input
flabel metal2 s 21510 8444 21600 8524 0 FreeSans 320 0 0 0 DOUT_SRAM8
port 106 nsew signal input
flabel metal2 s 21510 8948 21600 9028 0 FreeSans 320 0 0 0 DOUT_SRAM9
port 107 nsew signal input
flabel metal2 s 21510 58340 21600 58420 0 FreeSans 320 0 0 0 MEN_SRAM
port 108 nsew signal output
flabel metal2 s 21510 58844 21600 58924 0 FreeSans 320 0 0 0 REN_SRAM
port 109 nsew signal output
flabel metal2 s 21510 59348 21600 59428 0 FreeSans 320 0 0 0 TIE_HIGH_SRAM
port 110 nsew signal output
flabel metal2 s 21510 59852 21600 59932 0 FreeSans 320 0 0 0 TIE_LOW_SRAM
port 111 nsew signal output
flabel metal2 s 0 67244 90 67324 0 FreeSans 320 0 0 0 Tile_X0Y0_E1END[0]
port 112 nsew signal input
flabel metal2 s 0 67580 90 67660 0 FreeSans 320 0 0 0 Tile_X0Y0_E1END[1]
port 113 nsew signal input
flabel metal2 s 0 67916 90 67996 0 FreeSans 320 0 0 0 Tile_X0Y0_E1END[2]
port 114 nsew signal input
flabel metal2 s 0 68252 90 68332 0 FreeSans 320 0 0 0 Tile_X0Y0_E1END[3]
port 115 nsew signal input
flabel metal2 s 0 71276 90 71356 0 FreeSans 320 0 0 0 Tile_X0Y0_E2END[0]
port 116 nsew signal input
flabel metal2 s 0 71612 90 71692 0 FreeSans 320 0 0 0 Tile_X0Y0_E2END[1]
port 117 nsew signal input
flabel metal2 s 0 71948 90 72028 0 FreeSans 320 0 0 0 Tile_X0Y0_E2END[2]
port 118 nsew signal input
flabel metal2 s 0 72284 90 72364 0 FreeSans 320 0 0 0 Tile_X0Y0_E2END[3]
port 119 nsew signal input
flabel metal2 s 0 72620 90 72700 0 FreeSans 320 0 0 0 Tile_X0Y0_E2END[4]
port 120 nsew signal input
flabel metal2 s 0 72956 90 73036 0 FreeSans 320 0 0 0 Tile_X0Y0_E2END[5]
port 121 nsew signal input
flabel metal2 s 0 73292 90 73372 0 FreeSans 320 0 0 0 Tile_X0Y0_E2END[6]
port 122 nsew signal input
flabel metal2 s 0 73628 90 73708 0 FreeSans 320 0 0 0 Tile_X0Y0_E2END[7]
port 123 nsew signal input
flabel metal2 s 0 68588 90 68668 0 FreeSans 320 0 0 0 Tile_X0Y0_E2MID[0]
port 124 nsew signal input
flabel metal2 s 0 68924 90 69004 0 FreeSans 320 0 0 0 Tile_X0Y0_E2MID[1]
port 125 nsew signal input
flabel metal2 s 0 69260 90 69340 0 FreeSans 320 0 0 0 Tile_X0Y0_E2MID[2]
port 126 nsew signal input
flabel metal2 s 0 69596 90 69676 0 FreeSans 320 0 0 0 Tile_X0Y0_E2MID[3]
port 127 nsew signal input
flabel metal2 s 0 69932 90 70012 0 FreeSans 320 0 0 0 Tile_X0Y0_E2MID[4]
port 128 nsew signal input
flabel metal2 s 0 70268 90 70348 0 FreeSans 320 0 0 0 Tile_X0Y0_E2MID[5]
port 129 nsew signal input
flabel metal2 s 0 70604 90 70684 0 FreeSans 320 0 0 0 Tile_X0Y0_E2MID[6]
port 130 nsew signal input
flabel metal2 s 0 70940 90 71020 0 FreeSans 320 0 0 0 Tile_X0Y0_E2MID[7]
port 131 nsew signal input
flabel metal2 s 0 79340 90 79420 0 FreeSans 320 0 0 0 Tile_X0Y0_E6END[0]
port 132 nsew signal input
flabel metal2 s 0 82700 90 82780 0 FreeSans 320 0 0 0 Tile_X0Y0_E6END[10]
port 133 nsew signal input
flabel metal2 s 0 83036 90 83116 0 FreeSans 320 0 0 0 Tile_X0Y0_E6END[11]
port 134 nsew signal input
flabel metal2 s 0 79676 90 79756 0 FreeSans 320 0 0 0 Tile_X0Y0_E6END[1]
port 135 nsew signal input
flabel metal2 s 0 80012 90 80092 0 FreeSans 320 0 0 0 Tile_X0Y0_E6END[2]
port 136 nsew signal input
flabel metal2 s 0 80348 90 80428 0 FreeSans 320 0 0 0 Tile_X0Y0_E6END[3]
port 137 nsew signal input
flabel metal2 s 0 80684 90 80764 0 FreeSans 320 0 0 0 Tile_X0Y0_E6END[4]
port 138 nsew signal input
flabel metal2 s 0 81020 90 81100 0 FreeSans 320 0 0 0 Tile_X0Y0_E6END[5]
port 139 nsew signal input
flabel metal2 s 0 81356 90 81436 0 FreeSans 320 0 0 0 Tile_X0Y0_E6END[6]
port 140 nsew signal input
flabel metal2 s 0 81692 90 81772 0 FreeSans 320 0 0 0 Tile_X0Y0_E6END[7]
port 141 nsew signal input
flabel metal2 s 0 82028 90 82108 0 FreeSans 320 0 0 0 Tile_X0Y0_E6END[8]
port 142 nsew signal input
flabel metal2 s 0 82364 90 82444 0 FreeSans 320 0 0 0 Tile_X0Y0_E6END[9]
port 143 nsew signal input
flabel metal2 s 0 73964 90 74044 0 FreeSans 320 0 0 0 Tile_X0Y0_EE4END[0]
port 144 nsew signal input
flabel metal2 s 0 77324 90 77404 0 FreeSans 320 0 0 0 Tile_X0Y0_EE4END[10]
port 145 nsew signal input
flabel metal2 s 0 77660 90 77740 0 FreeSans 320 0 0 0 Tile_X0Y0_EE4END[11]
port 146 nsew signal input
flabel metal2 s 0 77996 90 78076 0 FreeSans 320 0 0 0 Tile_X0Y0_EE4END[12]
port 147 nsew signal input
flabel metal2 s 0 78332 90 78412 0 FreeSans 320 0 0 0 Tile_X0Y0_EE4END[13]
port 148 nsew signal input
flabel metal2 s 0 78668 90 78748 0 FreeSans 320 0 0 0 Tile_X0Y0_EE4END[14]
port 149 nsew signal input
flabel metal2 s 0 79004 90 79084 0 FreeSans 320 0 0 0 Tile_X0Y0_EE4END[15]
port 150 nsew signal input
flabel metal2 s 0 74300 90 74380 0 FreeSans 320 0 0 0 Tile_X0Y0_EE4END[1]
port 151 nsew signal input
flabel metal2 s 0 74636 90 74716 0 FreeSans 320 0 0 0 Tile_X0Y0_EE4END[2]
port 152 nsew signal input
flabel metal2 s 0 74972 90 75052 0 FreeSans 320 0 0 0 Tile_X0Y0_EE4END[3]
port 153 nsew signal input
flabel metal2 s 0 75308 90 75388 0 FreeSans 320 0 0 0 Tile_X0Y0_EE4END[4]
port 154 nsew signal input
flabel metal2 s 0 75644 90 75724 0 FreeSans 320 0 0 0 Tile_X0Y0_EE4END[5]
port 155 nsew signal input
flabel metal2 s 0 75980 90 76060 0 FreeSans 320 0 0 0 Tile_X0Y0_EE4END[6]
port 156 nsew signal input
flabel metal2 s 0 76316 90 76396 0 FreeSans 320 0 0 0 Tile_X0Y0_EE4END[7]
port 157 nsew signal input
flabel metal2 s 0 76652 90 76732 0 FreeSans 320 0 0 0 Tile_X0Y0_EE4END[8]
port 158 nsew signal input
flabel metal2 s 0 76988 90 77068 0 FreeSans 320 0 0 0 Tile_X0Y0_EE4END[9]
port 159 nsew signal input
flabel metal2 s 0 83372 90 83452 0 FreeSans 320 0 0 0 Tile_X0Y0_FrameData[0]
port 160 nsew signal input
flabel metal2 s 0 86732 90 86812 0 FreeSans 320 0 0 0 Tile_X0Y0_FrameData[10]
port 161 nsew signal input
flabel metal2 s 0 87068 90 87148 0 FreeSans 320 0 0 0 Tile_X0Y0_FrameData[11]
port 162 nsew signal input
flabel metal2 s 0 87404 90 87484 0 FreeSans 320 0 0 0 Tile_X0Y0_FrameData[12]
port 163 nsew signal input
flabel metal2 s 0 87740 90 87820 0 FreeSans 320 0 0 0 Tile_X0Y0_FrameData[13]
port 164 nsew signal input
flabel metal2 s 0 88076 90 88156 0 FreeSans 320 0 0 0 Tile_X0Y0_FrameData[14]
port 165 nsew signal input
flabel metal2 s 0 88412 90 88492 0 FreeSans 320 0 0 0 Tile_X0Y0_FrameData[15]
port 166 nsew signal input
flabel metal2 s 0 88748 90 88828 0 FreeSans 320 0 0 0 Tile_X0Y0_FrameData[16]
port 167 nsew signal input
flabel metal2 s 0 89084 90 89164 0 FreeSans 320 0 0 0 Tile_X0Y0_FrameData[17]
port 168 nsew signal input
flabel metal2 s 0 89420 90 89500 0 FreeSans 320 0 0 0 Tile_X0Y0_FrameData[18]
port 169 nsew signal input
flabel metal2 s 0 89756 90 89836 0 FreeSans 320 0 0 0 Tile_X0Y0_FrameData[19]
port 170 nsew signal input
flabel metal2 s 0 83708 90 83788 0 FreeSans 320 0 0 0 Tile_X0Y0_FrameData[1]
port 171 nsew signal input
flabel metal2 s 0 90092 90 90172 0 FreeSans 320 0 0 0 Tile_X0Y0_FrameData[20]
port 172 nsew signal input
flabel metal2 s 0 90428 90 90508 0 FreeSans 320 0 0 0 Tile_X0Y0_FrameData[21]
port 173 nsew signal input
flabel metal2 s 0 90764 90 90844 0 FreeSans 320 0 0 0 Tile_X0Y0_FrameData[22]
port 174 nsew signal input
flabel metal2 s 0 91100 90 91180 0 FreeSans 320 0 0 0 Tile_X0Y0_FrameData[23]
port 175 nsew signal input
flabel metal2 s 0 91436 90 91516 0 FreeSans 320 0 0 0 Tile_X0Y0_FrameData[24]
port 176 nsew signal input
flabel metal2 s 0 91772 90 91852 0 FreeSans 320 0 0 0 Tile_X0Y0_FrameData[25]
port 177 nsew signal input
flabel metal2 s 0 92108 90 92188 0 FreeSans 320 0 0 0 Tile_X0Y0_FrameData[26]
port 178 nsew signal input
flabel metal2 s 0 92444 90 92524 0 FreeSans 320 0 0 0 Tile_X0Y0_FrameData[27]
port 179 nsew signal input
flabel metal2 s 0 92780 90 92860 0 FreeSans 320 0 0 0 Tile_X0Y0_FrameData[28]
port 180 nsew signal input
flabel metal2 s 0 93116 90 93196 0 FreeSans 320 0 0 0 Tile_X0Y0_FrameData[29]
port 181 nsew signal input
flabel metal2 s 0 84044 90 84124 0 FreeSans 320 0 0 0 Tile_X0Y0_FrameData[2]
port 182 nsew signal input
flabel metal2 s 0 93452 90 93532 0 FreeSans 320 0 0 0 Tile_X0Y0_FrameData[30]
port 183 nsew signal input
flabel metal2 s 0 93788 90 93868 0 FreeSans 320 0 0 0 Tile_X0Y0_FrameData[31]
port 184 nsew signal input
flabel metal2 s 0 84380 90 84460 0 FreeSans 320 0 0 0 Tile_X0Y0_FrameData[3]
port 185 nsew signal input
flabel metal2 s 0 84716 90 84796 0 FreeSans 320 0 0 0 Tile_X0Y0_FrameData[4]
port 186 nsew signal input
flabel metal2 s 0 85052 90 85132 0 FreeSans 320 0 0 0 Tile_X0Y0_FrameData[5]
port 187 nsew signal input
flabel metal2 s 0 85388 90 85468 0 FreeSans 320 0 0 0 Tile_X0Y0_FrameData[6]
port 188 nsew signal input
flabel metal2 s 0 85724 90 85804 0 FreeSans 320 0 0 0 Tile_X0Y0_FrameData[7]
port 189 nsew signal input
flabel metal2 s 0 86060 90 86140 0 FreeSans 320 0 0 0 Tile_X0Y0_FrameData[8]
port 190 nsew signal input
flabel metal2 s 0 86396 90 86476 0 FreeSans 320 0 0 0 Tile_X0Y0_FrameData[9]
port 191 nsew signal input
flabel metal2 s 21510 60860 21600 60940 0 FreeSans 320 0 0 0 Tile_X0Y0_FrameData_O[0]
port 192 nsew signal output
flabel metal2 s 21510 65900 21600 65980 0 FreeSans 320 0 0 0 Tile_X0Y0_FrameData_O[10]
port 193 nsew signal output
flabel metal2 s 21510 66404 21600 66484 0 FreeSans 320 0 0 0 Tile_X0Y0_FrameData_O[11]
port 194 nsew signal output
flabel metal2 s 21510 66908 21600 66988 0 FreeSans 320 0 0 0 Tile_X0Y0_FrameData_O[12]
port 195 nsew signal output
flabel metal2 s 21510 67412 21600 67492 0 FreeSans 320 0 0 0 Tile_X0Y0_FrameData_O[13]
port 196 nsew signal output
flabel metal2 s 21510 67916 21600 67996 0 FreeSans 320 0 0 0 Tile_X0Y0_FrameData_O[14]
port 197 nsew signal output
flabel metal2 s 21510 68420 21600 68500 0 FreeSans 320 0 0 0 Tile_X0Y0_FrameData_O[15]
port 198 nsew signal output
flabel metal2 s 21510 68924 21600 69004 0 FreeSans 320 0 0 0 Tile_X0Y0_FrameData_O[16]
port 199 nsew signal output
flabel metal2 s 21510 69428 21600 69508 0 FreeSans 320 0 0 0 Tile_X0Y0_FrameData_O[17]
port 200 nsew signal output
flabel metal2 s 21510 69932 21600 70012 0 FreeSans 320 0 0 0 Tile_X0Y0_FrameData_O[18]
port 201 nsew signal output
flabel metal2 s 21510 70436 21600 70516 0 FreeSans 320 0 0 0 Tile_X0Y0_FrameData_O[19]
port 202 nsew signal output
flabel metal2 s 21510 61364 21600 61444 0 FreeSans 320 0 0 0 Tile_X0Y0_FrameData_O[1]
port 203 nsew signal output
flabel metal2 s 21510 70940 21600 71020 0 FreeSans 320 0 0 0 Tile_X0Y0_FrameData_O[20]
port 204 nsew signal output
flabel metal2 s 21510 71444 21600 71524 0 FreeSans 320 0 0 0 Tile_X0Y0_FrameData_O[21]
port 205 nsew signal output
flabel metal2 s 21510 71948 21600 72028 0 FreeSans 320 0 0 0 Tile_X0Y0_FrameData_O[22]
port 206 nsew signal output
flabel metal2 s 21510 72452 21600 72532 0 FreeSans 320 0 0 0 Tile_X0Y0_FrameData_O[23]
port 207 nsew signal output
flabel metal2 s 21510 72956 21600 73036 0 FreeSans 320 0 0 0 Tile_X0Y0_FrameData_O[24]
port 208 nsew signal output
flabel metal2 s 21510 73460 21600 73540 0 FreeSans 320 0 0 0 Tile_X0Y0_FrameData_O[25]
port 209 nsew signal output
flabel metal2 s 21510 73964 21600 74044 0 FreeSans 320 0 0 0 Tile_X0Y0_FrameData_O[26]
port 210 nsew signal output
flabel metal2 s 21510 74468 21600 74548 0 FreeSans 320 0 0 0 Tile_X0Y0_FrameData_O[27]
port 211 nsew signal output
flabel metal2 s 21510 74972 21600 75052 0 FreeSans 320 0 0 0 Tile_X0Y0_FrameData_O[28]
port 212 nsew signal output
flabel metal2 s 21510 75476 21600 75556 0 FreeSans 320 0 0 0 Tile_X0Y0_FrameData_O[29]
port 213 nsew signal output
flabel metal2 s 21510 61868 21600 61948 0 FreeSans 320 0 0 0 Tile_X0Y0_FrameData_O[2]
port 214 nsew signal output
flabel metal2 s 21510 75980 21600 76060 0 FreeSans 320 0 0 0 Tile_X0Y0_FrameData_O[30]
port 215 nsew signal output
flabel metal2 s 21510 76484 21600 76564 0 FreeSans 320 0 0 0 Tile_X0Y0_FrameData_O[31]
port 216 nsew signal output
flabel metal2 s 21510 62372 21600 62452 0 FreeSans 320 0 0 0 Tile_X0Y0_FrameData_O[3]
port 217 nsew signal output
flabel metal2 s 21510 62876 21600 62956 0 FreeSans 320 0 0 0 Tile_X0Y0_FrameData_O[4]
port 218 nsew signal output
flabel metal2 s 21510 63380 21600 63460 0 FreeSans 320 0 0 0 Tile_X0Y0_FrameData_O[5]
port 219 nsew signal output
flabel metal2 s 21510 63884 21600 63964 0 FreeSans 320 0 0 0 Tile_X0Y0_FrameData_O[6]
port 220 nsew signal output
flabel metal2 s 21510 64388 21600 64468 0 FreeSans 320 0 0 0 Tile_X0Y0_FrameData_O[7]
port 221 nsew signal output
flabel metal2 s 21510 64892 21600 64972 0 FreeSans 320 0 0 0 Tile_X0Y0_FrameData_O[8]
port 222 nsew signal output
flabel metal2 s 21510 65396 21600 65476 0 FreeSans 320 0 0 0 Tile_X0Y0_FrameData_O[9]
port 223 nsew signal output
flabel metal3 s 15800 96688 15880 96768 0 FreeSans 320 0 0 0 Tile_X0Y0_FrameStrobe_O[0]
port 224 nsew signal output
flabel metal3 s 17720 96688 17800 96768 0 FreeSans 320 0 0 0 Tile_X0Y0_FrameStrobe_O[10]
port 225 nsew signal output
flabel metal3 s 17912 96688 17992 96768 0 FreeSans 320 0 0 0 Tile_X0Y0_FrameStrobe_O[11]
port 226 nsew signal output
flabel metal3 s 18104 96688 18184 96768 0 FreeSans 320 0 0 0 Tile_X0Y0_FrameStrobe_O[12]
port 227 nsew signal output
flabel metal3 s 18296 96688 18376 96768 0 FreeSans 320 0 0 0 Tile_X0Y0_FrameStrobe_O[13]
port 228 nsew signal output
flabel metal3 s 18488 96688 18568 96768 0 FreeSans 320 0 0 0 Tile_X0Y0_FrameStrobe_O[14]
port 229 nsew signal output
flabel metal3 s 18680 96688 18760 96768 0 FreeSans 320 0 0 0 Tile_X0Y0_FrameStrobe_O[15]
port 230 nsew signal output
flabel metal3 s 18872 96688 18952 96768 0 FreeSans 320 0 0 0 Tile_X0Y0_FrameStrobe_O[16]
port 231 nsew signal output
flabel metal3 s 19064 96688 19144 96768 0 FreeSans 320 0 0 0 Tile_X0Y0_FrameStrobe_O[17]
port 232 nsew signal output
flabel metal3 s 19256 96688 19336 96768 0 FreeSans 320 0 0 0 Tile_X0Y0_FrameStrobe_O[18]
port 233 nsew signal output
flabel metal3 s 19448 96688 19528 96768 0 FreeSans 320 0 0 0 Tile_X0Y0_FrameStrobe_O[19]
port 234 nsew signal output
flabel metal3 s 15992 96688 16072 96768 0 FreeSans 320 0 0 0 Tile_X0Y0_FrameStrobe_O[1]
port 235 nsew signal output
flabel metal3 s 16184 96688 16264 96768 0 FreeSans 320 0 0 0 Tile_X0Y0_FrameStrobe_O[2]
port 236 nsew signal output
flabel metal3 s 16376 96688 16456 96768 0 FreeSans 320 0 0 0 Tile_X0Y0_FrameStrobe_O[3]
port 237 nsew signal output
flabel metal3 s 16568 96688 16648 96768 0 FreeSans 320 0 0 0 Tile_X0Y0_FrameStrobe_O[4]
port 238 nsew signal output
flabel metal3 s 16760 96688 16840 96768 0 FreeSans 320 0 0 0 Tile_X0Y0_FrameStrobe_O[5]
port 239 nsew signal output
flabel metal3 s 16952 96688 17032 96768 0 FreeSans 320 0 0 0 Tile_X0Y0_FrameStrobe_O[6]
port 240 nsew signal output
flabel metal3 s 17144 96688 17224 96768 0 FreeSans 320 0 0 0 Tile_X0Y0_FrameStrobe_O[7]
port 241 nsew signal output
flabel metal3 s 17336 96688 17416 96768 0 FreeSans 320 0 0 0 Tile_X0Y0_FrameStrobe_O[8]
port 242 nsew signal output
flabel metal3 s 17528 96688 17608 96768 0 FreeSans 320 0 0 0 Tile_X0Y0_FrameStrobe_O[9]
port 243 nsew signal output
flabel metal3 s 1784 96688 1864 96768 0 FreeSans 320 0 0 0 Tile_X0Y0_N1BEG[0]
port 244 nsew signal output
flabel metal3 s 1976 96688 2056 96768 0 FreeSans 320 0 0 0 Tile_X0Y0_N1BEG[1]
port 245 nsew signal output
flabel metal3 s 2168 96688 2248 96768 0 FreeSans 320 0 0 0 Tile_X0Y0_N1BEG[2]
port 246 nsew signal output
flabel metal3 s 2360 96688 2440 96768 0 FreeSans 320 0 0 0 Tile_X0Y0_N1BEG[3]
port 247 nsew signal output
flabel metal3 s 2552 96688 2632 96768 0 FreeSans 320 0 0 0 Tile_X0Y0_N2BEG[0]
port 248 nsew signal output
flabel metal3 s 2744 96688 2824 96768 0 FreeSans 320 0 0 0 Tile_X0Y0_N2BEG[1]
port 249 nsew signal output
flabel metal3 s 2936 96688 3016 96768 0 FreeSans 320 0 0 0 Tile_X0Y0_N2BEG[2]
port 250 nsew signal output
flabel metal3 s 3128 96688 3208 96768 0 FreeSans 320 0 0 0 Tile_X0Y0_N2BEG[3]
port 251 nsew signal output
flabel metal3 s 3320 96688 3400 96768 0 FreeSans 320 0 0 0 Tile_X0Y0_N2BEG[4]
port 252 nsew signal output
flabel metal3 s 3512 96688 3592 96768 0 FreeSans 320 0 0 0 Tile_X0Y0_N2BEG[5]
port 253 nsew signal output
flabel metal3 s 3704 96688 3784 96768 0 FreeSans 320 0 0 0 Tile_X0Y0_N2BEG[6]
port 254 nsew signal output
flabel metal3 s 3896 96688 3976 96768 0 FreeSans 320 0 0 0 Tile_X0Y0_N2BEG[7]
port 255 nsew signal output
flabel metal3 s 4088 96688 4168 96768 0 FreeSans 320 0 0 0 Tile_X0Y0_N2BEGb[0]
port 256 nsew signal output
flabel metal3 s 4280 96688 4360 96768 0 FreeSans 320 0 0 0 Tile_X0Y0_N2BEGb[1]
port 257 nsew signal output
flabel metal3 s 4472 96688 4552 96768 0 FreeSans 320 0 0 0 Tile_X0Y0_N2BEGb[2]
port 258 nsew signal output
flabel metal3 s 4664 96688 4744 96768 0 FreeSans 320 0 0 0 Tile_X0Y0_N2BEGb[3]
port 259 nsew signal output
flabel metal3 s 4856 96688 4936 96768 0 FreeSans 320 0 0 0 Tile_X0Y0_N2BEGb[4]
port 260 nsew signal output
flabel metal3 s 5048 96688 5128 96768 0 FreeSans 320 0 0 0 Tile_X0Y0_N2BEGb[5]
port 261 nsew signal output
flabel metal3 s 5240 96688 5320 96768 0 FreeSans 320 0 0 0 Tile_X0Y0_N2BEGb[6]
port 262 nsew signal output
flabel metal3 s 5432 96688 5512 96768 0 FreeSans 320 0 0 0 Tile_X0Y0_N2BEGb[7]
port 263 nsew signal output
flabel metal3 s 5624 96688 5704 96768 0 FreeSans 320 0 0 0 Tile_X0Y0_N4BEG[0]
port 264 nsew signal output
flabel metal3 s 7544 96688 7624 96768 0 FreeSans 320 0 0 0 Tile_X0Y0_N4BEG[10]
port 265 nsew signal output
flabel metal3 s 7736 96688 7816 96768 0 FreeSans 320 0 0 0 Tile_X0Y0_N4BEG[11]
port 266 nsew signal output
flabel metal3 s 7928 96688 8008 96768 0 FreeSans 320 0 0 0 Tile_X0Y0_N4BEG[12]
port 267 nsew signal output
flabel metal3 s 8120 96688 8200 96768 0 FreeSans 320 0 0 0 Tile_X0Y0_N4BEG[13]
port 268 nsew signal output
flabel metal3 s 8312 96688 8392 96768 0 FreeSans 320 0 0 0 Tile_X0Y0_N4BEG[14]
port 269 nsew signal output
flabel metal3 s 8504 96688 8584 96768 0 FreeSans 320 0 0 0 Tile_X0Y0_N4BEG[15]
port 270 nsew signal output
flabel metal3 s 5816 96688 5896 96768 0 FreeSans 320 0 0 0 Tile_X0Y0_N4BEG[1]
port 271 nsew signal output
flabel metal3 s 6008 96688 6088 96768 0 FreeSans 320 0 0 0 Tile_X0Y0_N4BEG[2]
port 272 nsew signal output
flabel metal3 s 6200 96688 6280 96768 0 FreeSans 320 0 0 0 Tile_X0Y0_N4BEG[3]
port 273 nsew signal output
flabel metal3 s 6392 96688 6472 96768 0 FreeSans 320 0 0 0 Tile_X0Y0_N4BEG[4]
port 274 nsew signal output
flabel metal3 s 6584 96688 6664 96768 0 FreeSans 320 0 0 0 Tile_X0Y0_N4BEG[5]
port 275 nsew signal output
flabel metal3 s 6776 96688 6856 96768 0 FreeSans 320 0 0 0 Tile_X0Y0_N4BEG[6]
port 276 nsew signal output
flabel metal3 s 6968 96688 7048 96768 0 FreeSans 320 0 0 0 Tile_X0Y0_N4BEG[7]
port 277 nsew signal output
flabel metal3 s 7160 96688 7240 96768 0 FreeSans 320 0 0 0 Tile_X0Y0_N4BEG[8]
port 278 nsew signal output
flabel metal3 s 7352 96688 7432 96768 0 FreeSans 320 0 0 0 Tile_X0Y0_N4BEG[9]
port 279 nsew signal output
flabel metal3 s 8696 96688 8776 96768 0 FreeSans 320 0 0 0 Tile_X0Y0_S1END[0]
port 280 nsew signal input
flabel metal3 s 8888 96688 8968 96768 0 FreeSans 320 0 0 0 Tile_X0Y0_S1END[1]
port 281 nsew signal input
flabel metal3 s 9080 96688 9160 96768 0 FreeSans 320 0 0 0 Tile_X0Y0_S1END[2]
port 282 nsew signal input
flabel metal3 s 9272 96688 9352 96768 0 FreeSans 320 0 0 0 Tile_X0Y0_S1END[3]
port 283 nsew signal input
flabel metal3 s 11000 96688 11080 96768 0 FreeSans 320 0 0 0 Tile_X0Y0_S2END[0]
port 284 nsew signal input
flabel metal3 s 11192 96688 11272 96768 0 FreeSans 320 0 0 0 Tile_X0Y0_S2END[1]
port 285 nsew signal input
flabel metal3 s 11384 96688 11464 96768 0 FreeSans 320 0 0 0 Tile_X0Y0_S2END[2]
port 286 nsew signal input
flabel metal3 s 11576 96688 11656 96768 0 FreeSans 320 0 0 0 Tile_X0Y0_S2END[3]
port 287 nsew signal input
flabel metal3 s 11768 96688 11848 96768 0 FreeSans 320 0 0 0 Tile_X0Y0_S2END[4]
port 288 nsew signal input
flabel metal3 s 11960 96688 12040 96768 0 FreeSans 320 0 0 0 Tile_X0Y0_S2END[5]
port 289 nsew signal input
flabel metal3 s 12152 96688 12232 96768 0 FreeSans 320 0 0 0 Tile_X0Y0_S2END[6]
port 290 nsew signal input
flabel metal3 s 12344 96688 12424 96768 0 FreeSans 320 0 0 0 Tile_X0Y0_S2END[7]
port 291 nsew signal input
flabel metal3 s 9464 96688 9544 96768 0 FreeSans 320 0 0 0 Tile_X0Y0_S2MID[0]
port 292 nsew signal input
flabel metal3 s 9656 96688 9736 96768 0 FreeSans 320 0 0 0 Tile_X0Y0_S2MID[1]
port 293 nsew signal input
flabel metal3 s 9848 96688 9928 96768 0 FreeSans 320 0 0 0 Tile_X0Y0_S2MID[2]
port 294 nsew signal input
flabel metal3 s 10040 96688 10120 96768 0 FreeSans 320 0 0 0 Tile_X0Y0_S2MID[3]
port 295 nsew signal input
flabel metal3 s 10232 96688 10312 96768 0 FreeSans 320 0 0 0 Tile_X0Y0_S2MID[4]
port 296 nsew signal input
flabel metal3 s 10424 96688 10504 96768 0 FreeSans 320 0 0 0 Tile_X0Y0_S2MID[5]
port 297 nsew signal input
flabel metal3 s 10616 96688 10696 96768 0 FreeSans 320 0 0 0 Tile_X0Y0_S2MID[6]
port 298 nsew signal input
flabel metal3 s 10808 96688 10888 96768 0 FreeSans 320 0 0 0 Tile_X0Y0_S2MID[7]
port 299 nsew signal input
flabel metal3 s 12536 96688 12616 96768 0 FreeSans 320 0 0 0 Tile_X0Y0_S4END[0]
port 300 nsew signal input
flabel metal3 s 14456 96688 14536 96768 0 FreeSans 320 0 0 0 Tile_X0Y0_S4END[10]
port 301 nsew signal input
flabel metal3 s 14648 96688 14728 96768 0 FreeSans 320 0 0 0 Tile_X0Y0_S4END[11]
port 302 nsew signal input
flabel metal3 s 14840 96688 14920 96768 0 FreeSans 320 0 0 0 Tile_X0Y0_S4END[12]
port 303 nsew signal input
flabel metal3 s 15032 96688 15112 96768 0 FreeSans 320 0 0 0 Tile_X0Y0_S4END[13]
port 304 nsew signal input
flabel metal3 s 15224 96688 15304 96768 0 FreeSans 320 0 0 0 Tile_X0Y0_S4END[14]
port 305 nsew signal input
flabel metal3 s 15416 96688 15496 96768 0 FreeSans 320 0 0 0 Tile_X0Y0_S4END[15]
port 306 nsew signal input
flabel metal3 s 12728 96688 12808 96768 0 FreeSans 320 0 0 0 Tile_X0Y0_S4END[1]
port 307 nsew signal input
flabel metal3 s 12920 96688 13000 96768 0 FreeSans 320 0 0 0 Tile_X0Y0_S4END[2]
port 308 nsew signal input
flabel metal3 s 13112 96688 13192 96768 0 FreeSans 320 0 0 0 Tile_X0Y0_S4END[3]
port 309 nsew signal input
flabel metal3 s 13304 96688 13384 96768 0 FreeSans 320 0 0 0 Tile_X0Y0_S4END[4]
port 310 nsew signal input
flabel metal3 s 13496 96688 13576 96768 0 FreeSans 320 0 0 0 Tile_X0Y0_S4END[5]
port 311 nsew signal input
flabel metal3 s 13688 96688 13768 96768 0 FreeSans 320 0 0 0 Tile_X0Y0_S4END[6]
port 312 nsew signal input
flabel metal3 s 13880 96688 13960 96768 0 FreeSans 320 0 0 0 Tile_X0Y0_S4END[7]
port 313 nsew signal input
flabel metal3 s 14072 96688 14152 96768 0 FreeSans 320 0 0 0 Tile_X0Y0_S4END[8]
port 314 nsew signal input
flabel metal3 s 14264 96688 14344 96768 0 FreeSans 320 0 0 0 Tile_X0Y0_S4END[9]
port 315 nsew signal input
flabel metal3 s 15608 96688 15688 96768 0 FreeSans 320 0 0 0 Tile_X0Y0_UserCLKo
port 316 nsew signal output
flabel metal2 s 0 51116 90 51196 0 FreeSans 320 0 0 0 Tile_X0Y0_W1BEG[0]
port 317 nsew signal output
flabel metal2 s 0 51452 90 51532 0 FreeSans 320 0 0 0 Tile_X0Y0_W1BEG[1]
port 318 nsew signal output
flabel metal2 s 0 51788 90 51868 0 FreeSans 320 0 0 0 Tile_X0Y0_W1BEG[2]
port 319 nsew signal output
flabel metal2 s 0 52124 90 52204 0 FreeSans 320 0 0 0 Tile_X0Y0_W1BEG[3]
port 320 nsew signal output
flabel metal2 s 0 52460 90 52540 0 FreeSans 320 0 0 0 Tile_X0Y0_W2BEG[0]
port 321 nsew signal output
flabel metal2 s 0 52796 90 52876 0 FreeSans 320 0 0 0 Tile_X0Y0_W2BEG[1]
port 322 nsew signal output
flabel metal2 s 0 53132 90 53212 0 FreeSans 320 0 0 0 Tile_X0Y0_W2BEG[2]
port 323 nsew signal output
flabel metal2 s 0 53468 90 53548 0 FreeSans 320 0 0 0 Tile_X0Y0_W2BEG[3]
port 324 nsew signal output
flabel metal2 s 0 53804 90 53884 0 FreeSans 320 0 0 0 Tile_X0Y0_W2BEG[4]
port 325 nsew signal output
flabel metal2 s 0 54140 90 54220 0 FreeSans 320 0 0 0 Tile_X0Y0_W2BEG[5]
port 326 nsew signal output
flabel metal2 s 0 54476 90 54556 0 FreeSans 320 0 0 0 Tile_X0Y0_W2BEG[6]
port 327 nsew signal output
flabel metal2 s 0 54812 90 54892 0 FreeSans 320 0 0 0 Tile_X0Y0_W2BEG[7]
port 328 nsew signal output
flabel metal2 s 0 55148 90 55228 0 FreeSans 320 0 0 0 Tile_X0Y0_W2BEGb[0]
port 329 nsew signal output
flabel metal2 s 0 55484 90 55564 0 FreeSans 320 0 0 0 Tile_X0Y0_W2BEGb[1]
port 330 nsew signal output
flabel metal2 s 0 55820 90 55900 0 FreeSans 320 0 0 0 Tile_X0Y0_W2BEGb[2]
port 331 nsew signal output
flabel metal2 s 0 56156 90 56236 0 FreeSans 320 0 0 0 Tile_X0Y0_W2BEGb[3]
port 332 nsew signal output
flabel metal2 s 0 56492 90 56572 0 FreeSans 320 0 0 0 Tile_X0Y0_W2BEGb[4]
port 333 nsew signal output
flabel metal2 s 0 56828 90 56908 0 FreeSans 320 0 0 0 Tile_X0Y0_W2BEGb[5]
port 334 nsew signal output
flabel metal2 s 0 57164 90 57244 0 FreeSans 320 0 0 0 Tile_X0Y0_W2BEGb[6]
port 335 nsew signal output
flabel metal2 s 0 57500 90 57580 0 FreeSans 320 0 0 0 Tile_X0Y0_W2BEGb[7]
port 336 nsew signal output
flabel metal2 s 0 63212 90 63292 0 FreeSans 320 0 0 0 Tile_X0Y0_W6BEG[0]
port 337 nsew signal output
flabel metal2 s 0 66572 90 66652 0 FreeSans 320 0 0 0 Tile_X0Y0_W6BEG[10]
port 338 nsew signal output
flabel metal2 s 0 66908 90 66988 0 FreeSans 320 0 0 0 Tile_X0Y0_W6BEG[11]
port 339 nsew signal output
flabel metal2 s 0 63548 90 63628 0 FreeSans 320 0 0 0 Tile_X0Y0_W6BEG[1]
port 340 nsew signal output
flabel metal2 s 0 63884 90 63964 0 FreeSans 320 0 0 0 Tile_X0Y0_W6BEG[2]
port 341 nsew signal output
flabel metal2 s 0 64220 90 64300 0 FreeSans 320 0 0 0 Tile_X0Y0_W6BEG[3]
port 342 nsew signal output
flabel metal2 s 0 64556 90 64636 0 FreeSans 320 0 0 0 Tile_X0Y0_W6BEG[4]
port 343 nsew signal output
flabel metal2 s 0 64892 90 64972 0 FreeSans 320 0 0 0 Tile_X0Y0_W6BEG[5]
port 344 nsew signal output
flabel metal2 s 0 65228 90 65308 0 FreeSans 320 0 0 0 Tile_X0Y0_W6BEG[6]
port 345 nsew signal output
flabel metal2 s 0 65564 90 65644 0 FreeSans 320 0 0 0 Tile_X0Y0_W6BEG[7]
port 346 nsew signal output
flabel metal2 s 0 65900 90 65980 0 FreeSans 320 0 0 0 Tile_X0Y0_W6BEG[8]
port 347 nsew signal output
flabel metal2 s 0 66236 90 66316 0 FreeSans 320 0 0 0 Tile_X0Y0_W6BEG[9]
port 348 nsew signal output
flabel metal2 s 0 57836 90 57916 0 FreeSans 320 0 0 0 Tile_X0Y0_WW4BEG[0]
port 349 nsew signal output
flabel metal2 s 0 61196 90 61276 0 FreeSans 320 0 0 0 Tile_X0Y0_WW4BEG[10]
port 350 nsew signal output
flabel metal2 s 0 61532 90 61612 0 FreeSans 320 0 0 0 Tile_X0Y0_WW4BEG[11]
port 351 nsew signal output
flabel metal2 s 0 61868 90 61948 0 FreeSans 320 0 0 0 Tile_X0Y0_WW4BEG[12]
port 352 nsew signal output
flabel metal2 s 0 62204 90 62284 0 FreeSans 320 0 0 0 Tile_X0Y0_WW4BEG[13]
port 353 nsew signal output
flabel metal2 s 0 62540 90 62620 0 FreeSans 320 0 0 0 Tile_X0Y0_WW4BEG[14]
port 354 nsew signal output
flabel metal2 s 0 62876 90 62956 0 FreeSans 320 0 0 0 Tile_X0Y0_WW4BEG[15]
port 355 nsew signal output
flabel metal2 s 0 58172 90 58252 0 FreeSans 320 0 0 0 Tile_X0Y0_WW4BEG[1]
port 356 nsew signal output
flabel metal2 s 0 58508 90 58588 0 FreeSans 320 0 0 0 Tile_X0Y0_WW4BEG[2]
port 357 nsew signal output
flabel metal2 s 0 58844 90 58924 0 FreeSans 320 0 0 0 Tile_X0Y0_WW4BEG[3]
port 358 nsew signal output
flabel metal2 s 0 59180 90 59260 0 FreeSans 320 0 0 0 Tile_X0Y0_WW4BEG[4]
port 359 nsew signal output
flabel metal2 s 0 59516 90 59596 0 FreeSans 320 0 0 0 Tile_X0Y0_WW4BEG[5]
port 360 nsew signal output
flabel metal2 s 0 59852 90 59932 0 FreeSans 320 0 0 0 Tile_X0Y0_WW4BEG[6]
port 361 nsew signal output
flabel metal2 s 0 60188 90 60268 0 FreeSans 320 0 0 0 Tile_X0Y0_WW4BEG[7]
port 362 nsew signal output
flabel metal2 s 0 60524 90 60604 0 FreeSans 320 0 0 0 Tile_X0Y0_WW4BEG[8]
port 363 nsew signal output
flabel metal2 s 0 60860 90 60940 0 FreeSans 320 0 0 0 Tile_X0Y0_WW4BEG[9]
port 364 nsew signal output
flabel metal2 s 0 18860 90 18940 0 FreeSans 320 0 0 0 Tile_X0Y1_E1END[0]
port 365 nsew signal input
flabel metal2 s 0 19196 90 19276 0 FreeSans 320 0 0 0 Tile_X0Y1_E1END[1]
port 366 nsew signal input
flabel metal2 s 0 19532 90 19612 0 FreeSans 320 0 0 0 Tile_X0Y1_E1END[2]
port 367 nsew signal input
flabel metal2 s 0 19868 90 19948 0 FreeSans 320 0 0 0 Tile_X0Y1_E1END[3]
port 368 nsew signal input
flabel metal2 s 0 22892 90 22972 0 FreeSans 320 0 0 0 Tile_X0Y1_E2END[0]
port 369 nsew signal input
flabel metal2 s 0 23228 90 23308 0 FreeSans 320 0 0 0 Tile_X0Y1_E2END[1]
port 370 nsew signal input
flabel metal2 s 0 23564 90 23644 0 FreeSans 320 0 0 0 Tile_X0Y1_E2END[2]
port 371 nsew signal input
flabel metal2 s 0 23900 90 23980 0 FreeSans 320 0 0 0 Tile_X0Y1_E2END[3]
port 372 nsew signal input
flabel metal2 s 0 24236 90 24316 0 FreeSans 320 0 0 0 Tile_X0Y1_E2END[4]
port 373 nsew signal input
flabel metal2 s 0 24572 90 24652 0 FreeSans 320 0 0 0 Tile_X0Y1_E2END[5]
port 374 nsew signal input
flabel metal2 s 0 24908 90 24988 0 FreeSans 320 0 0 0 Tile_X0Y1_E2END[6]
port 375 nsew signal input
flabel metal2 s 0 25244 90 25324 0 FreeSans 320 0 0 0 Tile_X0Y1_E2END[7]
port 376 nsew signal input
flabel metal2 s 0 20204 90 20284 0 FreeSans 320 0 0 0 Tile_X0Y1_E2MID[0]
port 377 nsew signal input
flabel metal2 s 0 20540 90 20620 0 FreeSans 320 0 0 0 Tile_X0Y1_E2MID[1]
port 378 nsew signal input
flabel metal2 s 0 20876 90 20956 0 FreeSans 320 0 0 0 Tile_X0Y1_E2MID[2]
port 379 nsew signal input
flabel metal2 s 0 21212 90 21292 0 FreeSans 320 0 0 0 Tile_X0Y1_E2MID[3]
port 380 nsew signal input
flabel metal2 s 0 21548 90 21628 0 FreeSans 320 0 0 0 Tile_X0Y1_E2MID[4]
port 381 nsew signal input
flabel metal2 s 0 21884 90 21964 0 FreeSans 320 0 0 0 Tile_X0Y1_E2MID[5]
port 382 nsew signal input
flabel metal2 s 0 22220 90 22300 0 FreeSans 320 0 0 0 Tile_X0Y1_E2MID[6]
port 383 nsew signal input
flabel metal2 s 0 22556 90 22636 0 FreeSans 320 0 0 0 Tile_X0Y1_E2MID[7]
port 384 nsew signal input
flabel metal2 s 0 30956 90 31036 0 FreeSans 320 0 0 0 Tile_X0Y1_E6END[0]
port 385 nsew signal input
flabel metal2 s 0 34316 90 34396 0 FreeSans 320 0 0 0 Tile_X0Y1_E6END[10]
port 386 nsew signal input
flabel metal2 s 0 34652 90 34732 0 FreeSans 320 0 0 0 Tile_X0Y1_E6END[11]
port 387 nsew signal input
flabel metal2 s 0 31292 90 31372 0 FreeSans 320 0 0 0 Tile_X0Y1_E6END[1]
port 388 nsew signal input
flabel metal2 s 0 31628 90 31708 0 FreeSans 320 0 0 0 Tile_X0Y1_E6END[2]
port 389 nsew signal input
flabel metal2 s 0 31964 90 32044 0 FreeSans 320 0 0 0 Tile_X0Y1_E6END[3]
port 390 nsew signal input
flabel metal2 s 0 32300 90 32380 0 FreeSans 320 0 0 0 Tile_X0Y1_E6END[4]
port 391 nsew signal input
flabel metal2 s 0 32636 90 32716 0 FreeSans 320 0 0 0 Tile_X0Y1_E6END[5]
port 392 nsew signal input
flabel metal2 s 0 32972 90 33052 0 FreeSans 320 0 0 0 Tile_X0Y1_E6END[6]
port 393 nsew signal input
flabel metal2 s 0 33308 90 33388 0 FreeSans 320 0 0 0 Tile_X0Y1_E6END[7]
port 394 nsew signal input
flabel metal2 s 0 33644 90 33724 0 FreeSans 320 0 0 0 Tile_X0Y1_E6END[8]
port 395 nsew signal input
flabel metal2 s 0 33980 90 34060 0 FreeSans 320 0 0 0 Tile_X0Y1_E6END[9]
port 396 nsew signal input
flabel metal2 s 0 25580 90 25660 0 FreeSans 320 0 0 0 Tile_X0Y1_EE4END[0]
port 397 nsew signal input
flabel metal2 s 0 28940 90 29020 0 FreeSans 320 0 0 0 Tile_X0Y1_EE4END[10]
port 398 nsew signal input
flabel metal2 s 0 29276 90 29356 0 FreeSans 320 0 0 0 Tile_X0Y1_EE4END[11]
port 399 nsew signal input
flabel metal2 s 0 29612 90 29692 0 FreeSans 320 0 0 0 Tile_X0Y1_EE4END[12]
port 400 nsew signal input
flabel metal2 s 0 29948 90 30028 0 FreeSans 320 0 0 0 Tile_X0Y1_EE4END[13]
port 401 nsew signal input
flabel metal2 s 0 30284 90 30364 0 FreeSans 320 0 0 0 Tile_X0Y1_EE4END[14]
port 402 nsew signal input
flabel metal2 s 0 30620 90 30700 0 FreeSans 320 0 0 0 Tile_X0Y1_EE4END[15]
port 403 nsew signal input
flabel metal2 s 0 25916 90 25996 0 FreeSans 320 0 0 0 Tile_X0Y1_EE4END[1]
port 404 nsew signal input
flabel metal2 s 0 26252 90 26332 0 FreeSans 320 0 0 0 Tile_X0Y1_EE4END[2]
port 405 nsew signal input
flabel metal2 s 0 26588 90 26668 0 FreeSans 320 0 0 0 Tile_X0Y1_EE4END[3]
port 406 nsew signal input
flabel metal2 s 0 26924 90 27004 0 FreeSans 320 0 0 0 Tile_X0Y1_EE4END[4]
port 407 nsew signal input
flabel metal2 s 0 27260 90 27340 0 FreeSans 320 0 0 0 Tile_X0Y1_EE4END[5]
port 408 nsew signal input
flabel metal2 s 0 27596 90 27676 0 FreeSans 320 0 0 0 Tile_X0Y1_EE4END[6]
port 409 nsew signal input
flabel metal2 s 0 27932 90 28012 0 FreeSans 320 0 0 0 Tile_X0Y1_EE4END[7]
port 410 nsew signal input
flabel metal2 s 0 28268 90 28348 0 FreeSans 320 0 0 0 Tile_X0Y1_EE4END[8]
port 411 nsew signal input
flabel metal2 s 0 28604 90 28684 0 FreeSans 320 0 0 0 Tile_X0Y1_EE4END[9]
port 412 nsew signal input
flabel metal2 s 0 34988 90 35068 0 FreeSans 320 0 0 0 Tile_X0Y1_FrameData[0]
port 413 nsew signal input
flabel metal2 s 0 38348 90 38428 0 FreeSans 320 0 0 0 Tile_X0Y1_FrameData[10]
port 414 nsew signal input
flabel metal2 s 0 38684 90 38764 0 FreeSans 320 0 0 0 Tile_X0Y1_FrameData[11]
port 415 nsew signal input
flabel metal2 s 0 39020 90 39100 0 FreeSans 320 0 0 0 Tile_X0Y1_FrameData[12]
port 416 nsew signal input
flabel metal2 s 0 39356 90 39436 0 FreeSans 320 0 0 0 Tile_X0Y1_FrameData[13]
port 417 nsew signal input
flabel metal2 s 0 39692 90 39772 0 FreeSans 320 0 0 0 Tile_X0Y1_FrameData[14]
port 418 nsew signal input
flabel metal2 s 0 40028 90 40108 0 FreeSans 320 0 0 0 Tile_X0Y1_FrameData[15]
port 419 nsew signal input
flabel metal2 s 0 40364 90 40444 0 FreeSans 320 0 0 0 Tile_X0Y1_FrameData[16]
port 420 nsew signal input
flabel metal2 s 0 40700 90 40780 0 FreeSans 320 0 0 0 Tile_X0Y1_FrameData[17]
port 421 nsew signal input
flabel metal2 s 0 41036 90 41116 0 FreeSans 320 0 0 0 Tile_X0Y1_FrameData[18]
port 422 nsew signal input
flabel metal2 s 0 41372 90 41452 0 FreeSans 320 0 0 0 Tile_X0Y1_FrameData[19]
port 423 nsew signal input
flabel metal2 s 0 35324 90 35404 0 FreeSans 320 0 0 0 Tile_X0Y1_FrameData[1]
port 424 nsew signal input
flabel metal2 s 0 41708 90 41788 0 FreeSans 320 0 0 0 Tile_X0Y1_FrameData[20]
port 425 nsew signal input
flabel metal2 s 0 42044 90 42124 0 FreeSans 320 0 0 0 Tile_X0Y1_FrameData[21]
port 426 nsew signal input
flabel metal2 s 0 42380 90 42460 0 FreeSans 320 0 0 0 Tile_X0Y1_FrameData[22]
port 427 nsew signal input
flabel metal2 s 0 42716 90 42796 0 FreeSans 320 0 0 0 Tile_X0Y1_FrameData[23]
port 428 nsew signal input
flabel metal2 s 0 43052 90 43132 0 FreeSans 320 0 0 0 Tile_X0Y1_FrameData[24]
port 429 nsew signal input
flabel metal2 s 0 43388 90 43468 0 FreeSans 320 0 0 0 Tile_X0Y1_FrameData[25]
port 430 nsew signal input
flabel metal2 s 0 43724 90 43804 0 FreeSans 320 0 0 0 Tile_X0Y1_FrameData[26]
port 431 nsew signal input
flabel metal2 s 0 44060 90 44140 0 FreeSans 320 0 0 0 Tile_X0Y1_FrameData[27]
port 432 nsew signal input
flabel metal2 s 0 44396 90 44476 0 FreeSans 320 0 0 0 Tile_X0Y1_FrameData[28]
port 433 nsew signal input
flabel metal2 s 0 44732 90 44812 0 FreeSans 320 0 0 0 Tile_X0Y1_FrameData[29]
port 434 nsew signal input
flabel metal2 s 0 35660 90 35740 0 FreeSans 320 0 0 0 Tile_X0Y1_FrameData[2]
port 435 nsew signal input
flabel metal2 s 0 45068 90 45148 0 FreeSans 320 0 0 0 Tile_X0Y1_FrameData[30]
port 436 nsew signal input
flabel metal2 s 0 45404 90 45484 0 FreeSans 320 0 0 0 Tile_X0Y1_FrameData[31]
port 437 nsew signal input
flabel metal2 s 0 35996 90 36076 0 FreeSans 320 0 0 0 Tile_X0Y1_FrameData[3]
port 438 nsew signal input
flabel metal2 s 0 36332 90 36412 0 FreeSans 320 0 0 0 Tile_X0Y1_FrameData[4]
port 439 nsew signal input
flabel metal2 s 0 36668 90 36748 0 FreeSans 320 0 0 0 Tile_X0Y1_FrameData[5]
port 440 nsew signal input
flabel metal2 s 0 37004 90 37084 0 FreeSans 320 0 0 0 Tile_X0Y1_FrameData[6]
port 441 nsew signal input
flabel metal2 s 0 37340 90 37420 0 FreeSans 320 0 0 0 Tile_X0Y1_FrameData[7]
port 442 nsew signal input
flabel metal2 s 0 37676 90 37756 0 FreeSans 320 0 0 0 Tile_X0Y1_FrameData[8]
port 443 nsew signal input
flabel metal2 s 0 38012 90 38092 0 FreeSans 320 0 0 0 Tile_X0Y1_FrameData[9]
port 444 nsew signal input
flabel metal2 s 21510 76988 21600 77068 0 FreeSans 320 0 0 0 Tile_X0Y1_FrameData_O[0]
port 445 nsew signal output
flabel metal2 s 21510 82028 21600 82108 0 FreeSans 320 0 0 0 Tile_X0Y1_FrameData_O[10]
port 446 nsew signal output
flabel metal2 s 21510 82532 21600 82612 0 FreeSans 320 0 0 0 Tile_X0Y1_FrameData_O[11]
port 447 nsew signal output
flabel metal2 s 21510 83036 21600 83116 0 FreeSans 320 0 0 0 Tile_X0Y1_FrameData_O[12]
port 448 nsew signal output
flabel metal2 s 21510 83540 21600 83620 0 FreeSans 320 0 0 0 Tile_X0Y1_FrameData_O[13]
port 449 nsew signal output
flabel metal2 s 21510 84044 21600 84124 0 FreeSans 320 0 0 0 Tile_X0Y1_FrameData_O[14]
port 450 nsew signal output
flabel metal2 s 21510 84548 21600 84628 0 FreeSans 320 0 0 0 Tile_X0Y1_FrameData_O[15]
port 451 nsew signal output
flabel metal2 s 21510 85052 21600 85132 0 FreeSans 320 0 0 0 Tile_X0Y1_FrameData_O[16]
port 452 nsew signal output
flabel metal2 s 21510 85556 21600 85636 0 FreeSans 320 0 0 0 Tile_X0Y1_FrameData_O[17]
port 453 nsew signal output
flabel metal2 s 21510 86060 21600 86140 0 FreeSans 320 0 0 0 Tile_X0Y1_FrameData_O[18]
port 454 nsew signal output
flabel metal2 s 21510 86564 21600 86644 0 FreeSans 320 0 0 0 Tile_X0Y1_FrameData_O[19]
port 455 nsew signal output
flabel metal2 s 21510 77492 21600 77572 0 FreeSans 320 0 0 0 Tile_X0Y1_FrameData_O[1]
port 456 nsew signal output
flabel metal2 s 21510 87068 21600 87148 0 FreeSans 320 0 0 0 Tile_X0Y1_FrameData_O[20]
port 457 nsew signal output
flabel metal2 s 21510 87572 21600 87652 0 FreeSans 320 0 0 0 Tile_X0Y1_FrameData_O[21]
port 458 nsew signal output
flabel metal2 s 21510 88076 21600 88156 0 FreeSans 320 0 0 0 Tile_X0Y1_FrameData_O[22]
port 459 nsew signal output
flabel metal2 s 21510 88580 21600 88660 0 FreeSans 320 0 0 0 Tile_X0Y1_FrameData_O[23]
port 460 nsew signal output
flabel metal2 s 21510 89084 21600 89164 0 FreeSans 320 0 0 0 Tile_X0Y1_FrameData_O[24]
port 461 nsew signal output
flabel metal2 s 21510 89588 21600 89668 0 FreeSans 320 0 0 0 Tile_X0Y1_FrameData_O[25]
port 462 nsew signal output
flabel metal2 s 21510 90092 21600 90172 0 FreeSans 320 0 0 0 Tile_X0Y1_FrameData_O[26]
port 463 nsew signal output
flabel metal2 s 21510 90596 21600 90676 0 FreeSans 320 0 0 0 Tile_X0Y1_FrameData_O[27]
port 464 nsew signal output
flabel metal2 s 21510 91100 21600 91180 0 FreeSans 320 0 0 0 Tile_X0Y1_FrameData_O[28]
port 465 nsew signal output
flabel metal2 s 21510 91604 21600 91684 0 FreeSans 320 0 0 0 Tile_X0Y1_FrameData_O[29]
port 466 nsew signal output
flabel metal2 s 21510 77996 21600 78076 0 FreeSans 320 0 0 0 Tile_X0Y1_FrameData_O[2]
port 467 nsew signal output
flabel metal2 s 21510 92108 21600 92188 0 FreeSans 320 0 0 0 Tile_X0Y1_FrameData_O[30]
port 468 nsew signal output
flabel metal2 s 21510 92612 21600 92692 0 FreeSans 320 0 0 0 Tile_X0Y1_FrameData_O[31]
port 469 nsew signal output
flabel metal2 s 21510 78500 21600 78580 0 FreeSans 320 0 0 0 Tile_X0Y1_FrameData_O[3]
port 470 nsew signal output
flabel metal2 s 21510 79004 21600 79084 0 FreeSans 320 0 0 0 Tile_X0Y1_FrameData_O[4]
port 471 nsew signal output
flabel metal2 s 21510 79508 21600 79588 0 FreeSans 320 0 0 0 Tile_X0Y1_FrameData_O[5]
port 472 nsew signal output
flabel metal2 s 21510 80012 21600 80092 0 FreeSans 320 0 0 0 Tile_X0Y1_FrameData_O[6]
port 473 nsew signal output
flabel metal2 s 21510 80516 21600 80596 0 FreeSans 320 0 0 0 Tile_X0Y1_FrameData_O[7]
port 474 nsew signal output
flabel metal2 s 21510 81020 21600 81100 0 FreeSans 320 0 0 0 Tile_X0Y1_FrameData_O[8]
port 475 nsew signal output
flabel metal2 s 21510 81524 21600 81604 0 FreeSans 320 0 0 0 Tile_X0Y1_FrameData_O[9]
port 476 nsew signal output
flabel metal3 s 15800 0 15880 80 0 FreeSans 320 0 0 0 Tile_X0Y1_FrameStrobe[0]
port 477 nsew signal input
flabel metal3 s 17720 0 17800 80 0 FreeSans 320 0 0 0 Tile_X0Y1_FrameStrobe[10]
port 478 nsew signal input
flabel metal3 s 17912 0 17992 80 0 FreeSans 320 0 0 0 Tile_X0Y1_FrameStrobe[11]
port 479 nsew signal input
flabel metal3 s 18104 0 18184 80 0 FreeSans 320 0 0 0 Tile_X0Y1_FrameStrobe[12]
port 480 nsew signal input
flabel metal3 s 18296 0 18376 80 0 FreeSans 320 0 0 0 Tile_X0Y1_FrameStrobe[13]
port 481 nsew signal input
flabel metal3 s 18488 0 18568 80 0 FreeSans 320 0 0 0 Tile_X0Y1_FrameStrobe[14]
port 482 nsew signal input
flabel metal3 s 18680 0 18760 80 0 FreeSans 320 0 0 0 Tile_X0Y1_FrameStrobe[15]
port 483 nsew signal input
flabel metal3 s 18872 0 18952 80 0 FreeSans 320 0 0 0 Tile_X0Y1_FrameStrobe[16]
port 484 nsew signal input
flabel metal3 s 19064 0 19144 80 0 FreeSans 320 0 0 0 Tile_X0Y1_FrameStrobe[17]
port 485 nsew signal input
flabel metal3 s 19256 0 19336 80 0 FreeSans 320 0 0 0 Tile_X0Y1_FrameStrobe[18]
port 486 nsew signal input
flabel metal3 s 19448 0 19528 80 0 FreeSans 320 0 0 0 Tile_X0Y1_FrameStrobe[19]
port 487 nsew signal input
flabel metal3 s 15992 0 16072 80 0 FreeSans 320 0 0 0 Tile_X0Y1_FrameStrobe[1]
port 488 nsew signal input
flabel metal3 s 16184 0 16264 80 0 FreeSans 320 0 0 0 Tile_X0Y1_FrameStrobe[2]
port 489 nsew signal input
flabel metal3 s 16376 0 16456 80 0 FreeSans 320 0 0 0 Tile_X0Y1_FrameStrobe[3]
port 490 nsew signal input
flabel metal3 s 16568 0 16648 80 0 FreeSans 320 0 0 0 Tile_X0Y1_FrameStrobe[4]
port 491 nsew signal input
flabel metal3 s 16760 0 16840 80 0 FreeSans 320 0 0 0 Tile_X0Y1_FrameStrobe[5]
port 492 nsew signal input
flabel metal3 s 16952 0 17032 80 0 FreeSans 320 0 0 0 Tile_X0Y1_FrameStrobe[6]
port 493 nsew signal input
flabel metal3 s 17144 0 17224 80 0 FreeSans 320 0 0 0 Tile_X0Y1_FrameStrobe[7]
port 494 nsew signal input
flabel metal3 s 17336 0 17416 80 0 FreeSans 320 0 0 0 Tile_X0Y1_FrameStrobe[8]
port 495 nsew signal input
flabel metal3 s 17528 0 17608 80 0 FreeSans 320 0 0 0 Tile_X0Y1_FrameStrobe[9]
port 496 nsew signal input
flabel metal3 s 1784 0 1864 80 0 FreeSans 320 0 0 0 Tile_X0Y1_N1END[0]
port 497 nsew signal input
flabel metal3 s 1976 0 2056 80 0 FreeSans 320 0 0 0 Tile_X0Y1_N1END[1]
port 498 nsew signal input
flabel metal3 s 2168 0 2248 80 0 FreeSans 320 0 0 0 Tile_X0Y1_N1END[2]
port 499 nsew signal input
flabel metal3 s 2360 0 2440 80 0 FreeSans 320 0 0 0 Tile_X0Y1_N1END[3]
port 500 nsew signal input
flabel metal3 s 4088 0 4168 80 0 FreeSans 320 0 0 0 Tile_X0Y1_N2END[0]
port 501 nsew signal input
flabel metal3 s 4280 0 4360 80 0 FreeSans 320 0 0 0 Tile_X0Y1_N2END[1]
port 502 nsew signal input
flabel metal3 s 4472 0 4552 80 0 FreeSans 320 0 0 0 Tile_X0Y1_N2END[2]
port 503 nsew signal input
flabel metal3 s 4664 0 4744 80 0 FreeSans 320 0 0 0 Tile_X0Y1_N2END[3]
port 504 nsew signal input
flabel metal3 s 4856 0 4936 80 0 FreeSans 320 0 0 0 Tile_X0Y1_N2END[4]
port 505 nsew signal input
flabel metal3 s 5048 0 5128 80 0 FreeSans 320 0 0 0 Tile_X0Y1_N2END[5]
port 506 nsew signal input
flabel metal3 s 5240 0 5320 80 0 FreeSans 320 0 0 0 Tile_X0Y1_N2END[6]
port 507 nsew signal input
flabel metal3 s 5432 0 5512 80 0 FreeSans 320 0 0 0 Tile_X0Y1_N2END[7]
port 508 nsew signal input
flabel metal3 s 2552 0 2632 80 0 FreeSans 320 0 0 0 Tile_X0Y1_N2MID[0]
port 509 nsew signal input
flabel metal3 s 2744 0 2824 80 0 FreeSans 320 0 0 0 Tile_X0Y1_N2MID[1]
port 510 nsew signal input
flabel metal3 s 2936 0 3016 80 0 FreeSans 320 0 0 0 Tile_X0Y1_N2MID[2]
port 511 nsew signal input
flabel metal3 s 3128 0 3208 80 0 FreeSans 320 0 0 0 Tile_X0Y1_N2MID[3]
port 512 nsew signal input
flabel metal3 s 3320 0 3400 80 0 FreeSans 320 0 0 0 Tile_X0Y1_N2MID[4]
port 513 nsew signal input
flabel metal3 s 3512 0 3592 80 0 FreeSans 320 0 0 0 Tile_X0Y1_N2MID[5]
port 514 nsew signal input
flabel metal3 s 3704 0 3784 80 0 FreeSans 320 0 0 0 Tile_X0Y1_N2MID[6]
port 515 nsew signal input
flabel metal3 s 3896 0 3976 80 0 FreeSans 320 0 0 0 Tile_X0Y1_N2MID[7]
port 516 nsew signal input
flabel metal3 s 5624 0 5704 80 0 FreeSans 320 0 0 0 Tile_X0Y1_N4END[0]
port 517 nsew signal input
flabel metal3 s 7544 0 7624 80 0 FreeSans 320 0 0 0 Tile_X0Y1_N4END[10]
port 518 nsew signal input
flabel metal3 s 7736 0 7816 80 0 FreeSans 320 0 0 0 Tile_X0Y1_N4END[11]
port 519 nsew signal input
flabel metal3 s 7928 0 8008 80 0 FreeSans 320 0 0 0 Tile_X0Y1_N4END[12]
port 520 nsew signal input
flabel metal3 s 8120 0 8200 80 0 FreeSans 320 0 0 0 Tile_X0Y1_N4END[13]
port 521 nsew signal input
flabel metal3 s 8312 0 8392 80 0 FreeSans 320 0 0 0 Tile_X0Y1_N4END[14]
port 522 nsew signal input
flabel metal3 s 8504 0 8584 80 0 FreeSans 320 0 0 0 Tile_X0Y1_N4END[15]
port 523 nsew signal input
flabel metal3 s 5816 0 5896 80 0 FreeSans 320 0 0 0 Tile_X0Y1_N4END[1]
port 524 nsew signal input
flabel metal3 s 6008 0 6088 80 0 FreeSans 320 0 0 0 Tile_X0Y1_N4END[2]
port 525 nsew signal input
flabel metal3 s 6200 0 6280 80 0 FreeSans 320 0 0 0 Tile_X0Y1_N4END[3]
port 526 nsew signal input
flabel metal3 s 6392 0 6472 80 0 FreeSans 320 0 0 0 Tile_X0Y1_N4END[4]
port 527 nsew signal input
flabel metal3 s 6584 0 6664 80 0 FreeSans 320 0 0 0 Tile_X0Y1_N4END[5]
port 528 nsew signal input
flabel metal3 s 6776 0 6856 80 0 FreeSans 320 0 0 0 Tile_X0Y1_N4END[6]
port 529 nsew signal input
flabel metal3 s 6968 0 7048 80 0 FreeSans 320 0 0 0 Tile_X0Y1_N4END[7]
port 530 nsew signal input
flabel metal3 s 7160 0 7240 80 0 FreeSans 320 0 0 0 Tile_X0Y1_N4END[8]
port 531 nsew signal input
flabel metal3 s 7352 0 7432 80 0 FreeSans 320 0 0 0 Tile_X0Y1_N4END[9]
port 532 nsew signal input
flabel metal3 s 8696 0 8776 80 0 FreeSans 320 0 0 0 Tile_X0Y1_S1BEG[0]
port 533 nsew signal output
flabel metal3 s 8888 0 8968 80 0 FreeSans 320 0 0 0 Tile_X0Y1_S1BEG[1]
port 534 nsew signal output
flabel metal3 s 9080 0 9160 80 0 FreeSans 320 0 0 0 Tile_X0Y1_S1BEG[2]
port 535 nsew signal output
flabel metal3 s 9272 0 9352 80 0 FreeSans 320 0 0 0 Tile_X0Y1_S1BEG[3]
port 536 nsew signal output
flabel metal3 s 9464 0 9544 80 0 FreeSans 320 0 0 0 Tile_X0Y1_S2BEG[0]
port 537 nsew signal output
flabel metal3 s 9656 0 9736 80 0 FreeSans 320 0 0 0 Tile_X0Y1_S2BEG[1]
port 538 nsew signal output
flabel metal3 s 9848 0 9928 80 0 FreeSans 320 0 0 0 Tile_X0Y1_S2BEG[2]
port 539 nsew signal output
flabel metal3 s 10040 0 10120 80 0 FreeSans 320 0 0 0 Tile_X0Y1_S2BEG[3]
port 540 nsew signal output
flabel metal3 s 10232 0 10312 80 0 FreeSans 320 0 0 0 Tile_X0Y1_S2BEG[4]
port 541 nsew signal output
flabel metal3 s 10424 0 10504 80 0 FreeSans 320 0 0 0 Tile_X0Y1_S2BEG[5]
port 542 nsew signal output
flabel metal3 s 10616 0 10696 80 0 FreeSans 320 0 0 0 Tile_X0Y1_S2BEG[6]
port 543 nsew signal output
flabel metal3 s 10808 0 10888 80 0 FreeSans 320 0 0 0 Tile_X0Y1_S2BEG[7]
port 544 nsew signal output
flabel metal3 s 11000 0 11080 80 0 FreeSans 320 0 0 0 Tile_X0Y1_S2BEGb[0]
port 545 nsew signal output
flabel metal3 s 11192 0 11272 80 0 FreeSans 320 0 0 0 Tile_X0Y1_S2BEGb[1]
port 546 nsew signal output
flabel metal3 s 11384 0 11464 80 0 FreeSans 320 0 0 0 Tile_X0Y1_S2BEGb[2]
port 547 nsew signal output
flabel metal3 s 11576 0 11656 80 0 FreeSans 320 0 0 0 Tile_X0Y1_S2BEGb[3]
port 548 nsew signal output
flabel metal3 s 11768 0 11848 80 0 FreeSans 320 0 0 0 Tile_X0Y1_S2BEGb[4]
port 549 nsew signal output
flabel metal3 s 11960 0 12040 80 0 FreeSans 320 0 0 0 Tile_X0Y1_S2BEGb[5]
port 550 nsew signal output
flabel metal3 s 12152 0 12232 80 0 FreeSans 320 0 0 0 Tile_X0Y1_S2BEGb[6]
port 551 nsew signal output
flabel metal3 s 12344 0 12424 80 0 FreeSans 320 0 0 0 Tile_X0Y1_S2BEGb[7]
port 552 nsew signal output
flabel metal3 s 12536 0 12616 80 0 FreeSans 320 0 0 0 Tile_X0Y1_S4BEG[0]
port 553 nsew signal output
flabel metal3 s 14456 0 14536 80 0 FreeSans 320 0 0 0 Tile_X0Y1_S4BEG[10]
port 554 nsew signal output
flabel metal3 s 14648 0 14728 80 0 FreeSans 320 0 0 0 Tile_X0Y1_S4BEG[11]
port 555 nsew signal output
flabel metal3 s 14840 0 14920 80 0 FreeSans 320 0 0 0 Tile_X0Y1_S4BEG[12]
port 556 nsew signal output
flabel metal3 s 15032 0 15112 80 0 FreeSans 320 0 0 0 Tile_X0Y1_S4BEG[13]
port 557 nsew signal output
flabel metal3 s 15224 0 15304 80 0 FreeSans 320 0 0 0 Tile_X0Y1_S4BEG[14]
port 558 nsew signal output
flabel metal3 s 15416 0 15496 80 0 FreeSans 320 0 0 0 Tile_X0Y1_S4BEG[15]
port 559 nsew signal output
flabel metal3 s 12728 0 12808 80 0 FreeSans 320 0 0 0 Tile_X0Y1_S4BEG[1]
port 560 nsew signal output
flabel metal3 s 12920 0 13000 80 0 FreeSans 320 0 0 0 Tile_X0Y1_S4BEG[2]
port 561 nsew signal output
flabel metal3 s 13112 0 13192 80 0 FreeSans 320 0 0 0 Tile_X0Y1_S4BEG[3]
port 562 nsew signal output
flabel metal3 s 13304 0 13384 80 0 FreeSans 320 0 0 0 Tile_X0Y1_S4BEG[4]
port 563 nsew signal output
flabel metal3 s 13496 0 13576 80 0 FreeSans 320 0 0 0 Tile_X0Y1_S4BEG[5]
port 564 nsew signal output
flabel metal3 s 13688 0 13768 80 0 FreeSans 320 0 0 0 Tile_X0Y1_S4BEG[6]
port 565 nsew signal output
flabel metal3 s 13880 0 13960 80 0 FreeSans 320 0 0 0 Tile_X0Y1_S4BEG[7]
port 566 nsew signal output
flabel metal3 s 14072 0 14152 80 0 FreeSans 320 0 0 0 Tile_X0Y1_S4BEG[8]
port 567 nsew signal output
flabel metal3 s 14264 0 14344 80 0 FreeSans 320 0 0 0 Tile_X0Y1_S4BEG[9]
port 568 nsew signal output
flabel metal3 s 15608 0 15688 80 0 FreeSans 320 0 0 0 Tile_X0Y1_UserCLK
port 569 nsew signal input
flabel metal2 s 0 2732 90 2812 0 FreeSans 320 0 0 0 Tile_X0Y1_W1BEG[0]
port 570 nsew signal output
flabel metal2 s 0 3068 90 3148 0 FreeSans 320 0 0 0 Tile_X0Y1_W1BEG[1]
port 571 nsew signal output
flabel metal2 s 0 3404 90 3484 0 FreeSans 320 0 0 0 Tile_X0Y1_W1BEG[2]
port 572 nsew signal output
flabel metal2 s 0 3740 90 3820 0 FreeSans 320 0 0 0 Tile_X0Y1_W1BEG[3]
port 573 nsew signal output
flabel metal2 s 0 4076 90 4156 0 FreeSans 320 0 0 0 Tile_X0Y1_W2BEG[0]
port 574 nsew signal output
flabel metal2 s 0 4412 90 4492 0 FreeSans 320 0 0 0 Tile_X0Y1_W2BEG[1]
port 575 nsew signal output
flabel metal2 s 0 4748 90 4828 0 FreeSans 320 0 0 0 Tile_X0Y1_W2BEG[2]
port 576 nsew signal output
flabel metal2 s 0 5084 90 5164 0 FreeSans 320 0 0 0 Tile_X0Y1_W2BEG[3]
port 577 nsew signal output
flabel metal2 s 0 5420 90 5500 0 FreeSans 320 0 0 0 Tile_X0Y1_W2BEG[4]
port 578 nsew signal output
flabel metal2 s 0 5756 90 5836 0 FreeSans 320 0 0 0 Tile_X0Y1_W2BEG[5]
port 579 nsew signal output
flabel metal2 s 0 6092 90 6172 0 FreeSans 320 0 0 0 Tile_X0Y1_W2BEG[6]
port 580 nsew signal output
flabel metal2 s 0 6428 90 6508 0 FreeSans 320 0 0 0 Tile_X0Y1_W2BEG[7]
port 581 nsew signal output
flabel metal2 s 0 6764 90 6844 0 FreeSans 320 0 0 0 Tile_X0Y1_W2BEGb[0]
port 582 nsew signal output
flabel metal2 s 0 7100 90 7180 0 FreeSans 320 0 0 0 Tile_X0Y1_W2BEGb[1]
port 583 nsew signal output
flabel metal2 s 0 7436 90 7516 0 FreeSans 320 0 0 0 Tile_X0Y1_W2BEGb[2]
port 584 nsew signal output
flabel metal2 s 0 7772 90 7852 0 FreeSans 320 0 0 0 Tile_X0Y1_W2BEGb[3]
port 585 nsew signal output
flabel metal2 s 0 8108 90 8188 0 FreeSans 320 0 0 0 Tile_X0Y1_W2BEGb[4]
port 586 nsew signal output
flabel metal2 s 0 8444 90 8524 0 FreeSans 320 0 0 0 Tile_X0Y1_W2BEGb[5]
port 587 nsew signal output
flabel metal2 s 0 8780 90 8860 0 FreeSans 320 0 0 0 Tile_X0Y1_W2BEGb[6]
port 588 nsew signal output
flabel metal2 s 0 9116 90 9196 0 FreeSans 320 0 0 0 Tile_X0Y1_W2BEGb[7]
port 589 nsew signal output
flabel metal2 s 0 14828 90 14908 0 FreeSans 320 0 0 0 Tile_X0Y1_W6BEG[0]
port 590 nsew signal output
flabel metal2 s 0 18188 90 18268 0 FreeSans 320 0 0 0 Tile_X0Y1_W6BEG[10]
port 591 nsew signal output
flabel metal2 s 0 18524 90 18604 0 FreeSans 320 0 0 0 Tile_X0Y1_W6BEG[11]
port 592 nsew signal output
flabel metal2 s 0 15164 90 15244 0 FreeSans 320 0 0 0 Tile_X0Y1_W6BEG[1]
port 593 nsew signal output
flabel metal2 s 0 15500 90 15580 0 FreeSans 320 0 0 0 Tile_X0Y1_W6BEG[2]
port 594 nsew signal output
flabel metal2 s 0 15836 90 15916 0 FreeSans 320 0 0 0 Tile_X0Y1_W6BEG[3]
port 595 nsew signal output
flabel metal2 s 0 16172 90 16252 0 FreeSans 320 0 0 0 Tile_X0Y1_W6BEG[4]
port 596 nsew signal output
flabel metal2 s 0 16508 90 16588 0 FreeSans 320 0 0 0 Tile_X0Y1_W6BEG[5]
port 597 nsew signal output
flabel metal2 s 0 16844 90 16924 0 FreeSans 320 0 0 0 Tile_X0Y1_W6BEG[6]
port 598 nsew signal output
flabel metal2 s 0 17180 90 17260 0 FreeSans 320 0 0 0 Tile_X0Y1_W6BEG[7]
port 599 nsew signal output
flabel metal2 s 0 17516 90 17596 0 FreeSans 320 0 0 0 Tile_X0Y1_W6BEG[8]
port 600 nsew signal output
flabel metal2 s 0 17852 90 17932 0 FreeSans 320 0 0 0 Tile_X0Y1_W6BEG[9]
port 601 nsew signal output
flabel metal2 s 0 9452 90 9532 0 FreeSans 320 0 0 0 Tile_X0Y1_WW4BEG[0]
port 602 nsew signal output
flabel metal2 s 0 12812 90 12892 0 FreeSans 320 0 0 0 Tile_X0Y1_WW4BEG[10]
port 603 nsew signal output
flabel metal2 s 0 13148 90 13228 0 FreeSans 320 0 0 0 Tile_X0Y1_WW4BEG[11]
port 604 nsew signal output
flabel metal2 s 0 13484 90 13564 0 FreeSans 320 0 0 0 Tile_X0Y1_WW4BEG[12]
port 605 nsew signal output
flabel metal2 s 0 13820 90 13900 0 FreeSans 320 0 0 0 Tile_X0Y1_WW4BEG[13]
port 606 nsew signal output
flabel metal2 s 0 14156 90 14236 0 FreeSans 320 0 0 0 Tile_X0Y1_WW4BEG[14]
port 607 nsew signal output
flabel metal2 s 0 14492 90 14572 0 FreeSans 320 0 0 0 Tile_X0Y1_WW4BEG[15]
port 608 nsew signal output
flabel metal2 s 0 9788 90 9868 0 FreeSans 320 0 0 0 Tile_X0Y1_WW4BEG[1]
port 609 nsew signal output
flabel metal2 s 0 10124 90 10204 0 FreeSans 320 0 0 0 Tile_X0Y1_WW4BEG[2]
port 610 nsew signal output
flabel metal2 s 0 10460 90 10540 0 FreeSans 320 0 0 0 Tile_X0Y1_WW4BEG[3]
port 611 nsew signal output
flabel metal2 s 0 10796 90 10876 0 FreeSans 320 0 0 0 Tile_X0Y1_WW4BEG[4]
port 612 nsew signal output
flabel metal2 s 0 11132 90 11212 0 FreeSans 320 0 0 0 Tile_X0Y1_WW4BEG[5]
port 613 nsew signal output
flabel metal2 s 0 11468 90 11548 0 FreeSans 320 0 0 0 Tile_X0Y1_WW4BEG[6]
port 614 nsew signal output
flabel metal2 s 0 11804 90 11884 0 FreeSans 320 0 0 0 Tile_X0Y1_WW4BEG[7]
port 615 nsew signal output
flabel metal2 s 0 12140 90 12220 0 FreeSans 320 0 0 0 Tile_X0Y1_WW4BEG[8]
port 616 nsew signal output
flabel metal2 s 0 12476 90 12556 0 FreeSans 320 0 0 0 Tile_X0Y1_WW4BEG[9]
port 617 nsew signal output
flabel metal5 s 4892 0 5332 96768 0 FreeSans 2560 90 0 0 VGND
port 618 nsew ground bidirectional
flabel metal5 s 4892 0 5332 40 0 FreeSans 320 0 0 0 VGND
port 618 nsew ground bidirectional
flabel metal5 s 4892 96728 5332 96768 0 FreeSans 320 0 0 0 VGND
port 618 nsew ground bidirectional
flabel metal5 s 20012 0 20452 96768 0 FreeSans 2560 90 0 0 VGND
port 618 nsew ground bidirectional
flabel metal5 s 20012 0 20452 40 0 FreeSans 320 0 0 0 VGND
port 618 nsew ground bidirectional
flabel metal5 s 20012 96728 20452 96768 0 FreeSans 320 0 0 0 VGND
port 618 nsew ground bidirectional
flabel metal5 s 3652 0 4092 96768 0 FreeSans 2560 90 0 0 VPWR
port 619 nsew power bidirectional
flabel metal5 s 3652 0 4092 40 0 FreeSans 320 0 0 0 VPWR
port 619 nsew power bidirectional
flabel metal5 s 3652 96728 4092 96768 0 FreeSans 320 0 0 0 VPWR
port 619 nsew power bidirectional
flabel metal5 s 18772 0 19212 96768 0 FreeSans 2560 90 0 0 VPWR
port 619 nsew power bidirectional
flabel metal5 s 18772 0 19212 40 0 FreeSans 320 0 0 0 VPWR
port 619 nsew power bidirectional
flabel metal5 s 18772 96728 19212 96768 0 FreeSans 320 0 0 0 VPWR
port 619 nsew power bidirectional
flabel metal2 s 21510 60356 21600 60436 0 FreeSans 320 0 0 0 WEN_SRAM
port 620 nsew signal output
rlabel metal1 10802 95256 10802 95256 0 VGND
rlabel metal1 10800 94500 10800 94500 0 VPWR
rlabel metal2 17400 19488 17400 19488 0 ADDR_SRAM0
rlabel metal2 18120 18312 18120 18312 0 ADDR_SRAM1
rlabel metal2 19704 17220 19704 17220 0 ADDR_SRAM2
rlabel metal2 20664 17136 20664 17136 0 ADDR_SRAM3
rlabel metal2 20712 17220 20712 17220 0 ADDR_SRAM4
rlabel metal2 20760 17976 20760 17976 0 ADDR_SRAM5
rlabel metal2 20616 18648 20616 18648 0 ADDR_SRAM6
rlabel metal2 19695 24108 19695 24108 0 ADDR_SRAM7
rlabel metal3 21120 24738 21120 24738 0 ADDR_SRAM8
rlabel metal2 20568 21000 20568 21000 0 ADDR_SRAM9
rlabel metal2 21039 25620 21039 25620 0 BM_SRAM0
rlabel metal2 20847 26124 20847 26124 0 BM_SRAM1
rlabel metal2 21216 30786 21216 30786 0 BM_SRAM10
rlabel metal2 20223 31164 20223 31164 0 BM_SRAM11
rlabel metal2 20832 31584 20832 31584 0 BM_SRAM12
rlabel metal2 19224 30828 19224 30828 0 BM_SRAM13
rlabel metal2 20520 29316 20520 29316 0 BM_SRAM14
rlabel metal2 21087 33180 21087 33180 0 BM_SRAM15
rlabel metal2 19944 30072 19944 30072 0 BM_SRAM16
rlabel metal2 21327 34188 21327 34188 0 BM_SRAM17
rlabel metal2 21279 34692 21279 34692 0 BM_SRAM18
rlabel metal2 21039 35196 21039 35196 0 BM_SRAM19
rlabel metal2 19032 23268 19032 23268 0 BM_SRAM2
rlabel metal2 19680 33180 19680 33180 0 BM_SRAM20
rlabel metal2 21231 36204 21231 36204 0 BM_SRAM21
rlabel metal2 15144 35868 15144 35868 0 BM_SRAM22
rlabel metal2 16968 34524 16968 34524 0 BM_SRAM23
rlabel metal2 21279 37716 21279 37716 0 BM_SRAM24
rlabel metal2 19656 34524 19656 34524 0 BM_SRAM25
rlabel metal2 19944 34524 19944 34524 0 BM_SRAM26
rlabel metal2 20520 34524 20520 34524 0 BM_SRAM27
rlabel metal2 19392 40152 19392 40152 0 BM_SRAM28
rlabel metal2 20511 40236 20511 40236 0 BM_SRAM29
rlabel metal2 18936 23940 18936 23940 0 BM_SRAM3
rlabel metal2 19224 39816 19224 39816 0 BM_SRAM30
rlabel metal2 19368 39900 19368 39900 0 BM_SRAM31
rlabel metal2 19272 24780 19272 24780 0 BM_SRAM4
rlabel metal2 19656 24612 19656 24612 0 BM_SRAM5
rlabel metal2 19944 24780 19944 24780 0 BM_SRAM6
rlabel metal2 20712 24780 20712 24780 0 BM_SRAM7
rlabel metal2 20616 25452 20616 25452 0 BM_SRAM8
rlabel metal2 20760 25536 20760 25536 0 BM_SRAM9
rlabel metal2 18408 40656 18408 40656 0 CLK_SRAM
rlabel metal2 20943 3948 20943 3948 0 CONFIGURED_top
rlabel metal2 20520 41328 20520 41328 0 DIN_SRAM0
rlabel metal2 20472 42168 20472 42168 0 DIN_SRAM1
rlabel metal2 20967 47292 20967 47292 0 DIN_SRAM10
rlabel metal2 21183 47796 21183 47796 0 DIN_SRAM11
rlabel metal2 20400 48258 20400 48258 0 DIN_SRAM12
rlabel metal2 21375 48804 21375 48804 0 DIN_SRAM13
rlabel metal2 21183 49308 21183 49308 0 DIN_SRAM14
rlabel metal2 20400 49770 20400 49770 0 DIN_SRAM15
rlabel metal2 21135 50316 21135 50316 0 DIN_SRAM16
rlabel metal2 21183 50820 21183 50820 0 DIN_SRAM17
rlabel metal2 21279 51324 21279 51324 0 DIN_SRAM18
rlabel metal2 20991 51828 20991 51828 0 DIN_SRAM19
rlabel metal2 20904 42924 20904 42924 0 DIN_SRAM2
rlabel metal2 19704 51240 19704 51240 0 DIN_SRAM20
rlabel metal2 20664 55356 20664 55356 0 DIN_SRAM21
rlabel metal2 21183 53340 21183 53340 0 DIN_SRAM22
rlabel metal2 21279 53844 21279 53844 0 DIN_SRAM23
rlabel metal2 21087 54348 21087 54348 0 DIN_SRAM24
rlabel metal2 21135 54852 21135 54852 0 DIN_SRAM25
rlabel metal2 17832 54264 17832 54264 0 DIN_SRAM26
rlabel metal2 20607 55860 20607 55860 0 DIN_SRAM27
rlabel metal2 21231 56364 21231 56364 0 DIN_SRAM28
rlabel metal2 21183 56868 21183 56868 0 DIN_SRAM29
rlabel metal2 20400 43722 20400 43722 0 DIN_SRAM3
rlabel metal4 20784 62328 20784 62328 0 DIN_SRAM30
rlabel metal2 21135 57876 21135 57876 0 DIN_SRAM31
rlabel metal2 21279 44268 21279 44268 0 DIN_SRAM4
rlabel metal2 20967 44772 20967 44772 0 DIN_SRAM5
rlabel metal2 21231 45276 21231 45276 0 DIN_SRAM6
rlabel metal2 21087 45780 21087 45780 0 DIN_SRAM7
rlabel metal2 20967 46284 20967 46284 0 DIN_SRAM8
rlabel metal2 21135 46788 21135 46788 0 DIN_SRAM9
rlabel metal2 20751 4452 20751 4452 0 DOUT_SRAM0
rlabel metal2 21087 4956 21087 4956 0 DOUT_SRAM1
rlabel metal2 21375 9492 21375 9492 0 DOUT_SRAM10
rlabel metal2 21327 9996 21327 9996 0 DOUT_SRAM11
rlabel metal2 20559 10500 20559 10500 0 DOUT_SRAM12
rlabel metal2 21471 11004 21471 11004 0 DOUT_SRAM13
rlabel metal2 21135 11508 21135 11508 0 DOUT_SRAM14
rlabel metal2 21279 12012 21279 12012 0 DOUT_SRAM15
rlabel metal2 17856 13524 17856 13524 0 DOUT_SRAM16
rlabel metal2 21231 13020 21231 13020 0 DOUT_SRAM17
rlabel metal2 20415 13524 20415 13524 0 DOUT_SRAM18
rlabel metal2 21183 14028 21183 14028 0 DOUT_SRAM19
rlabel metal2 21423 5460 21423 5460 0 DOUT_SRAM2
rlabel metal2 20655 14532 20655 14532 0 DOUT_SRAM20
rlabel metal2 19680 14574 19680 14574 0 DOUT_SRAM21
rlabel metal2 21375 15540 21375 15540 0 DOUT_SRAM22
rlabel metal2 21471 16044 21471 16044 0 DOUT_SRAM23
rlabel metal2 21279 16548 21279 16548 0 DOUT_SRAM24
rlabel metal3 19872 15708 19872 15708 0 DOUT_SRAM25
rlabel metal2 21231 17556 21231 17556 0 DOUT_SRAM26
rlabel metal2 20463 18060 20463 18060 0 DOUT_SRAM27
rlabel metal2 20895 18564 20895 18564 0 DOUT_SRAM28
rlabel metal2 21135 19068 21135 19068 0 DOUT_SRAM29
rlabel metal2 20367 5964 20367 5964 0 DOUT_SRAM3
rlabel metal2 20928 19656 20928 19656 0 DOUT_SRAM30
rlabel metal2 21375 20076 21375 20076 0 DOUT_SRAM31
rlabel metal2 21135 6468 21135 6468 0 DOUT_SRAM4
rlabel metal2 20559 6972 20559 6972 0 DOUT_SRAM5
rlabel metal2 21039 7476 21039 7476 0 DOUT_SRAM6
rlabel metal2 21519 7980 21519 7980 0 DOUT_SRAM7
rlabel metal2 21231 8484 21231 8484 0 DOUT_SRAM8
rlabel metal2 20511 8988 20511 8988 0 DOUT_SRAM9
rlabel metal2 21327 58380 21327 58380 0 MEN_SRAM
rlabel metal2 19887 58884 19887 58884 0 REN_SRAM
rlabel metal2 960 75180 960 75180 0 Tile_X0Y0_E1END[0]
rlabel metal3 1440 74760 1440 74760 0 Tile_X0Y0_E1END[1]
rlabel metal2 1440 75096 1440 75096 0 Tile_X0Y0_E1END[2]
rlabel metal2 560 68292 560 68292 0 Tile_X0Y0_E1END[3]
rlabel metal2 1184 71316 1184 71316 0 Tile_X0Y0_E2END[0]
rlabel metal2 656 71652 656 71652 0 Tile_X0Y0_E2END[1]
rlabel metal2 320 71988 320 71988 0 Tile_X0Y0_E2END[2]
rlabel metal2 80 72324 80 72324 0 Tile_X0Y0_E2END[3]
rlabel metal2 1008 80556 1008 80556 0 Tile_X0Y0_E2END[4]
rlabel metal2 672 81228 672 81228 0 Tile_X0Y0_E2END[5]
rlabel metal5 384 74676 384 74676 0 Tile_X0Y0_E2END[6]
rlabel metal2 176 73668 176 73668 0 Tile_X0Y0_E2END[7]
rlabel via2 80 68628 80 68628 0 Tile_X0Y0_E2MID[0]
rlabel metal2 656 68964 656 68964 0 Tile_X0Y0_E2MID[1]
rlabel metal2 864 77532 864 77532 0 Tile_X0Y0_E2MID[2]
rlabel metal2 1344 77490 1344 77490 0 Tile_X0Y0_E2MID[3]
rlabel metal2 80 69972 80 69972 0 Tile_X0Y0_E2MID[4]
rlabel metal2 720 79044 720 79044 0 Tile_X0Y0_E2MID[5]
rlabel metal2 416 70644 416 70644 0 Tile_X0Y0_E2MID[6]
rlabel metal2 10368 72198 10368 72198 0 Tile_X0Y0_E2MID[7]
rlabel metal2 320 79380 320 79380 0 Tile_X0Y0_E6END[0]
rlabel metal2 80 82740 80 82740 0 Tile_X0Y0_E6END[10]
rlabel metal2 80 83076 80 83076 0 Tile_X0Y0_E6END[11]
rlabel metal2 224 79716 224 79716 0 Tile_X0Y0_E6END[1]
rlabel metal2 272 80052 272 80052 0 Tile_X0Y0_E6END[2]
rlabel metal2 368 80388 368 80388 0 Tile_X0Y0_E6END[3]
rlabel metal2 608 80724 608 80724 0 Tile_X0Y0_E6END[4]
rlabel metal2 512 81060 512 81060 0 Tile_X0Y0_E6END[5]
rlabel metal2 128 81396 128 81396 0 Tile_X0Y0_E6END[6]
rlabel via2 80 81732 80 81732 0 Tile_X0Y0_E6END[7]
rlabel metal2 752 82068 752 82068 0 Tile_X0Y0_E6END[8]
rlabel metal2 1472 82404 1472 82404 0 Tile_X0Y0_E6END[9]
rlabel metal2 224 74004 224 74004 0 Tile_X0Y0_EE4END[0]
rlabel metal2 1616 77364 1616 77364 0 Tile_X0Y0_EE4END[10]
rlabel metal2 10656 79590 10656 79590 0 Tile_X0Y0_EE4END[11]
rlabel metal2 704 78036 704 78036 0 Tile_X0Y0_EE4END[12]
rlabel metal2 464 78372 464 78372 0 Tile_X0Y0_EE4END[13]
rlabel metal2 992 78708 992 78708 0 Tile_X0Y0_EE4END[14]
rlabel metal2 80 79044 80 79044 0 Tile_X0Y0_EE4END[15]
rlabel metal2 944 74340 944 74340 0 Tile_X0Y0_EE4END[1]
rlabel metal2 320 74676 320 74676 0 Tile_X0Y0_EE4END[2]
rlabel metal2 320 75012 320 75012 0 Tile_X0Y0_EE4END[3]
rlabel metal2 176 75348 176 75348 0 Tile_X0Y0_EE4END[4]
rlabel metal2 512 75684 512 75684 0 Tile_X0Y0_EE4END[5]
rlabel metal2 752 76020 752 76020 0 Tile_X0Y0_EE4END[6]
rlabel metal2 1472 76356 1472 76356 0 Tile_X0Y0_EE4END[7]
rlabel metal2 656 76692 656 76692 0 Tile_X0Y0_EE4END[8]
rlabel metal2 2288 77028 2288 77028 0 Tile_X0Y0_EE4END[9]
rlabel metal2 560 83412 560 83412 0 Tile_X0Y0_FrameData[0]
rlabel metal2 752 86772 752 86772 0 Tile_X0Y0_FrameData[10]
rlabel metal2 416 87108 416 87108 0 Tile_X0Y0_FrameData[11]
rlabel metal2 800 87444 800 87444 0 Tile_X0Y0_FrameData[12]
rlabel metal2 1328 87780 1328 87780 0 Tile_X0Y0_FrameData[13]
rlabel metal2 608 88116 608 88116 0 Tile_X0Y0_FrameData[14]
rlabel metal2 608 88452 608 88452 0 Tile_X0Y0_FrameData[15]
rlabel via2 80 88788 80 88788 0 Tile_X0Y0_FrameData[16]
rlabel metal3 3552 89712 3552 89712 0 Tile_X0Y0_FrameData[17]
rlabel metal2 752 89460 752 89460 0 Tile_X0Y0_FrameData[18]
rlabel metal2 128 89796 128 89796 0 Tile_X0Y0_FrameData[19]
rlabel metal2 1424 83748 1424 83748 0 Tile_X0Y0_FrameData[1]
rlabel metal2 656 90132 656 90132 0 Tile_X0Y0_FrameData[20]
rlabel metal2 752 90468 752 90468 0 Tile_X0Y0_FrameData[21]
rlabel metal2 704 90804 704 90804 0 Tile_X0Y0_FrameData[22]
rlabel metal2 416 91140 416 91140 0 Tile_X0Y0_FrameData[23]
rlabel metal2 128 91476 128 91476 0 Tile_X0Y0_FrameData[24]
rlabel metal2 272 91812 272 91812 0 Tile_X0Y0_FrameData[25]
rlabel metal2 848 92148 848 92148 0 Tile_X0Y0_FrameData[26]
rlabel metal2 1232 92484 1232 92484 0 Tile_X0Y0_FrameData[27]
rlabel metal2 704 92820 704 92820 0 Tile_X0Y0_FrameData[28]
rlabel metal2 656 93156 656 93156 0 Tile_X0Y0_FrameData[29]
rlabel metal2 704 84084 704 84084 0 Tile_X0Y0_FrameData[2]
rlabel metal2 1232 93492 1232 93492 0 Tile_X0Y0_FrameData[30]
rlabel via2 80 93828 80 93828 0 Tile_X0Y0_FrameData[31]
rlabel metal2 128 84420 128 84420 0 Tile_X0Y0_FrameData[3]
rlabel metal2 752 84756 752 84756 0 Tile_X0Y0_FrameData[4]
rlabel metal2 464 85092 464 85092 0 Tile_X0Y0_FrameData[5]
rlabel metal2 176 85428 176 85428 0 Tile_X0Y0_FrameData[6]
rlabel metal2 512 85764 512 85764 0 Tile_X0Y0_FrameData[7]
rlabel metal2 608 86100 608 86100 0 Tile_X0Y0_FrameData[8]
rlabel metal2 128 86436 128 86436 0 Tile_X0Y0_FrameData[9]
rlabel via2 21519 60900 21519 60900 0 Tile_X0Y0_FrameData_O[0]
rlabel via2 21519 65940 21519 65940 0 Tile_X0Y0_FrameData_O[10]
rlabel metal4 20496 69720 20496 69720 0 Tile_X0Y0_FrameData_O[11]
rlabel metal4 20496 69804 20496 69804 0 Tile_X0Y0_FrameData_O[12]
rlabel metal2 20856 74256 20856 74256 0 Tile_X0Y0_FrameData_O[13]
rlabel metal3 20256 68754 20256 68754 0 Tile_X0Y0_FrameData_O[14]
rlabel metal2 19080 73500 19080 73500 0 Tile_X0Y0_FrameData_O[15]
rlabel metal2 20664 75768 20664 75768 0 Tile_X0Y0_FrameData_O[16]
rlabel metal2 21471 69468 21471 69468 0 Tile_X0Y0_FrameData_O[17]
rlabel metal3 19200 73878 19200 73878 0 Tile_X0Y0_FrameData_O[18]
rlabel metal2 20127 70476 20127 70476 0 Tile_X0Y0_FrameData_O[19]
rlabel metal2 21471 61404 21471 61404 0 Tile_X0Y0_FrameData_O[1]
rlabel metal2 20415 70980 20415 70980 0 Tile_X0Y0_FrameData_O[20]
rlabel metal2 20943 71484 20943 71484 0 Tile_X0Y0_FrameData_O[21]
rlabel metal3 20448 76188 20448 76188 0 Tile_X0Y0_FrameData_O[22]
rlabel metal2 20712 79632 20712 79632 0 Tile_X0Y0_FrameData_O[23]
rlabel metal2 21327 72996 21327 72996 0 Tile_X0Y0_FrameData_O[24]
rlabel metal2 21375 73500 21375 73500 0 Tile_X0Y0_FrameData_O[25]
rlabel metal2 21375 74004 21375 74004 0 Tile_X0Y0_FrameData_O[26]
rlabel metal2 20943 74508 20943 74508 0 Tile_X0Y0_FrameData_O[27]
rlabel metal2 21423 75012 21423 75012 0 Tile_X0Y0_FrameData_O[28]
rlabel metal2 21327 75516 21327 75516 0 Tile_X0Y0_FrameData_O[29]
rlabel metal4 20976 63084 20976 63084 0 Tile_X0Y0_FrameData_O[2]
rlabel metal2 20895 76020 20895 76020 0 Tile_X0Y0_FrameData_O[30]
rlabel metal2 19968 76314 19968 76314 0 Tile_X0Y0_FrameData_O[31]
rlabel metal2 19440 62496 19440 62496 0 Tile_X0Y0_FrameData_O[3]
rlabel metal2 20928 63084 20928 63084 0 Tile_X0Y0_FrameData_O[4]
rlabel metal2 21375 63420 21375 63420 0 Tile_X0Y0_FrameData_O[5]
rlabel metal3 21120 64344 21120 64344 0 Tile_X0Y0_FrameData_O[6]
rlabel metal3 21024 69090 21024 69090 0 Tile_X0Y0_FrameData_O[7]
rlabel metal2 21327 64932 21327 64932 0 Tile_X0Y0_FrameData_O[8]
rlabel metal2 20799 65436 20799 65436 0 Tile_X0Y0_FrameData_O[9]
rlabel metal2 16008 95004 16008 95004 0 Tile_X0Y0_FrameStrobe_O[0]
rlabel metal2 19416 94668 19416 94668 0 Tile_X0Y0_FrameStrobe_O[10]
rlabel metal2 18888 94164 18888 94164 0 Tile_X0Y0_FrameStrobe_O[11]
rlabel metal2 19464 95004 19464 95004 0 Tile_X0Y0_FrameStrobe_O[12]
rlabel metal2 19080 93912 19080 93912 0 Tile_X0Y0_FrameStrobe_O[13]
rlabel metal2 18552 93576 18552 93576 0 Tile_X0Y0_FrameStrobe_O[14]
rlabel metal2 18600 93492 18600 93492 0 Tile_X0Y0_FrameStrobe_O[15]
rlabel metal3 19104 94668 19104 94668 0 Tile_X0Y0_FrameStrobe_O[16]
rlabel metal4 19296 94836 19296 94836 0 Tile_X0Y0_FrameStrobe_O[17]
rlabel metal3 19344 94752 19344 94752 0 Tile_X0Y0_FrameStrobe_O[18]
rlabel metal4 19344 94248 19344 94248 0 Tile_X0Y0_FrameStrobe_O[19]
rlabel metal2 16248 94668 16248 94668 0 Tile_X0Y0_FrameStrobe_O[1]
rlabel metal2 16536 95004 16536 95004 0 Tile_X0Y0_FrameStrobe_O[2]
rlabel metal2 17112 95004 17112 95004 0 Tile_X0Y0_FrameStrobe_O[3]
rlabel metal3 16608 95688 16608 95688 0 Tile_X0Y0_FrameStrobe_O[4]
rlabel metal2 17760 94626 17760 94626 0 Tile_X0Y0_FrameStrobe_O[5]
rlabel metal2 17856 94962 17856 94962 0 Tile_X0Y0_FrameStrobe_O[6]
rlabel metal2 18648 95004 18648 95004 0 Tile_X0Y0_FrameStrobe_O[7]
rlabel metal2 18648 94668 18648 94668 0 Tile_X0Y0_FrameStrobe_O[8]
rlabel metal2 18264 93912 18264 93912 0 Tile_X0Y0_FrameStrobe_O[9]
rlabel via1 10184 58652 10184 58652 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame0_bit0.Q
rlabel metal3 8640 58884 8640 58884 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame0_bit1.Q
rlabel metal2 17280 51114 17280 51114 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame0_bit10.Q
rlabel metal2 15744 51114 15744 51114 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame0_bit11.Q
rlabel metal2 11712 48762 11712 48762 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame0_bit12.Q
rlabel metal2 13368 48720 13368 48720 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame0_bit13.Q
rlabel metal2 4161 48048 4161 48048 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame0_bit14.Q
rlabel metal3 5760 49056 5760 49056 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame0_bit15.Q
rlabel metal2 4808 47208 4808 47208 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame0_bit16.Q
rlabel metal2 3360 47250 3360 47250 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame0_bit17.Q
rlabel metal2 18912 50232 18912 50232 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame0_bit18.Q
rlabel via1 20258 50232 20258 50232 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame0_bit19.Q
rlabel metal2 17601 69888 17601 69888 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame0_bit2.Q
rlabel metal3 15360 49392 15360 49392 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame0_bit20.Q
rlabel via1 16904 48739 16904 48739 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame0_bit21.Q
rlabel metal2 10568 50232 10568 50232 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame0_bit22.Q
rlabel metal2 9216 49980 9216 49980 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame0_bit23.Q
rlabel metal2 10944 58044 10944 58044 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame0_bit24.Q
rlabel metal2 11088 57288 11088 57288 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame0_bit25.Q
rlabel metal2 17472 73206 17472 73206 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame0_bit26.Q
rlabel metal4 18336 72744 18336 72744 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame0_bit27.Q
rlabel metal3 13248 79338 13248 79338 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame0_bit28.Q
rlabel metal2 12552 78876 12552 78876 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame0_bit29.Q
rlabel metal2 19272 69888 19272 69888 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame0_bit3.Q
rlabel metal2 3360 78330 3360 78330 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame0_bit30.Q
rlabel metal2 3264 79884 3264 79884 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame0_bit31.Q
rlabel metal2 10992 81984 10992 81984 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame0_bit4.Q
rlabel metal2 12680 81984 12680 81984 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame0_bit5.Q
rlabel metal3 2688 75474 2688 75474 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame0_bit6.Q
rlabel metal2 5064 74424 5064 74424 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame0_bit7.Q
rlabel via2 6632 48720 6632 48720 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame0_bit8.Q
rlabel metal2 5088 48762 5088 48762 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame0_bit9.Q
rlabel metal2 17232 75768 17232 75768 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame1_bit0.Q
rlabel metal2 17760 75978 17760 75978 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame1_bit1.Q
rlabel metal2 18336 69258 18336 69258 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame1_bit10.Q
rlabel metal3 19872 69888 19872 69888 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame1_bit11.Q
rlabel metal2 11265 83496 11265 83496 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame1_bit12.Q
rlabel metal2 12680 83496 12680 83496 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame1_bit13.Q
rlabel metal2 3393 75936 3393 75936 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame1_bit14.Q
rlabel metal2 5064 75936 5064 75936 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame1_bit15.Q
rlabel metal2 8256 55608 8256 55608 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame1_bit16.Q
rlabel metal3 9984 55860 9984 55860 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame1_bit17.Q
rlabel metal2 18369 72240 18369 72240 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame1_bit18.Q
rlabel metal3 20016 74256 20016 74256 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame1_bit19.Q
rlabel via1 12971 86520 12971 86520 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame1_bit2.Q
rlabel metal2 11328 81354 11328 81354 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame1_bit20.Q
rlabel metal2 12672 81312 12672 81312 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame1_bit21.Q
rlabel metal2 3216 81816 3216 81816 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame1_bit22.Q
rlabel metal2 5040 78288 5040 78288 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame1_bit23.Q
rlabel metal2 9360 54096 9360 54096 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame1_bit24.Q
rlabel metal3 10944 54726 10944 54726 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame1_bit25.Q
rlabel metal2 18000 71400 18000 71400 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame1_bit26.Q
rlabel metal2 19920 73500 19920 73500 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame1_bit27.Q
rlabel metal2 10944 82824 10944 82824 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame1_bit28.Q
rlabel metal2 12864 82824 12864 82824 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame1_bit29.Q
rlabel metal2 12768 87276 12768 87276 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame1_bit3.Q
rlabel metal2 3168 76734 3168 76734 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame1_bit30.Q
rlabel metal3 4704 78498 4704 78498 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame1_bit31.Q
rlabel via2 3744 54852 3744 54852 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame1_bit4.Q
rlabel metal2 3840 54726 3840 54726 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame1_bit5.Q
rlabel metal2 6339 69720 6339 69720 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame1_bit6.Q
rlabel metal2 7200 70686 7200 70686 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame1_bit7.Q
rlabel metal2 9408 54768 9408 54768 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame1_bit8.Q
rlabel metal3 11328 54516 11328 54516 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame1_bit9.Q
rlabel metal2 18432 81354 18432 81354 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame2_bit0.Q
rlabel metal2 20352 81312 20352 81312 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame2_bit1.Q
rlabel metal2 17856 84378 17856 84378 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame2_bit10.Q
rlabel metal3 19392 84966 19392 84966 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame2_bit11.Q
rlabel metal2 4560 88032 4560 88032 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame2_bit12.Q
rlabel metal2 6344 88032 6344 88032 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame2_bit13.Q
rlabel metal2 9504 65394 9504 65394 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame2_bit14.Q
rlabel via2 11048 65352 11048 65352 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame2_bit15.Q
rlabel metal2 17376 86520 17376 86520 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame2_bit16.Q
rlabel metal2 18920 86520 18920 86520 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame2_bit17.Q
rlabel metal3 13056 89880 13056 89880 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame2_bit18.Q
rlabel metal2 14736 89586 14736 89586 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame2_bit19.Q
rlabel metal3 12192 88578 12192 88578 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame2_bit2.Q
rlabel metal2 3120 81984 3120 81984 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame2_bit20.Q
rlabel metal2 4616 81984 4616 81984 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame2_bit21.Q
rlabel metal2 5232 52584 5232 52584 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame2_bit22.Q
rlabel metal3 6912 52668 6912 52668 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame2_bit23.Q
rlabel metal3 13440 55608 13440 55608 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame2_bit24.Q
rlabel via2 14888 56280 14888 56280 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame2_bit25.Q
rlabel metal2 15168 85050 15168 85050 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame2_bit26.Q
rlabel metal2 16824 85008 16824 85008 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame2_bit27.Q
rlabel metal2 4560 86520 4560 86520 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame2_bit28.Q
rlabel metal2 6056 86520 6056 86520 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame2_bit29.Q
rlabel metal2 14112 88914 14112 88914 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame2_bit3.Q
rlabel metal2 7728 77280 7728 77280 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame2_bit30.Q
rlabel metal2 7248 76608 7248 76608 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame2_bit31.Q
rlabel metal2 3072 82824 3072 82824 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame2_bit4.Q
rlabel metal2 4800 82866 4800 82866 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame2_bit5.Q
rlabel metal2 6240 54138 6240 54138 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame2_bit6.Q
rlabel metal3 7776 54348 7776 54348 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame2_bit7.Q
rlabel metal3 15072 55650 15072 55650 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame2_bit8.Q
rlabel metal2 16856 56280 16856 56280 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame2_bit9.Q
rlabel metal2 18369 81984 18369 81984 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame3_bit0.Q
rlabel metal2 19832 81984 19832 81984 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame3_bit1.Q
rlabel metal2 17568 83454 17568 83454 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame3_bit10.Q
rlabel metal2 19560 83496 19560 83496 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame3_bit11.Q
rlabel metal2 4833 87360 4833 87360 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame3_bit12.Q
rlabel metal3 6432 88368 6432 88368 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame3_bit13.Q
rlabel metal2 9552 64680 9552 64680 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame3_bit14.Q
rlabel metal3 11136 65688 11136 65688 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame3_bit15.Q
rlabel metal2 19263 87360 19263 87360 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame3_bit16.Q
rlabel metal3 17664 88368 17664 88368 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame3_bit17.Q
rlabel metal2 14496 88872 14496 88872 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame3_bit18.Q
rlabel metal3 16128 89502 16128 89502 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame3_bit19.Q
rlabel metal2 13008 88032 13008 88032 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame3_bit2.Q
rlabel metal2 3360 83496 3360 83496 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame3_bit20.Q
rlabel metal2 4904 83496 4904 83496 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame3_bit21.Q
rlabel metal2 5952 51492 5952 51492 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame3_bit22.Q
rlabel metal2 7544 51240 7544 51240 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame3_bit23.Q
rlabel metal2 13248 57162 13248 57162 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame3_bit24.Q
rlabel metal2 13920 56532 13920 56532 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame3_bit25.Q
rlabel metal2 15168 84378 15168 84378 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame3_bit26.Q
rlabel metal2 16848 84336 16848 84336 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame3_bit27.Q
rlabel metal2 7008 87402 7008 87402 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame3_bit28.Q
rlabel metal2 8736 87360 8736 87360 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame3_bit29.Q
rlabel metal2 14808 88032 14808 88032 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame3_bit3.Q
rlabel metal2 9552 61656 9552 61656 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame3_bit30.Q
rlabel metal2 11232 61614 11232 61614 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame3_bit31.Q
rlabel metal2 2784 84378 2784 84378 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame3_bit4.Q
rlabel metal3 4320 84924 4320 84924 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame3_bit5.Q
rlabel metal2 6657 53256 6657 53256 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame3_bit6.Q
rlabel via2 8264 53256 8264 53256 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame3_bit7.Q
rlabel metal2 15360 55650 15360 55650 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame3_bit8.Q
rlabel metal3 16896 56238 16896 56238 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame3_bit9.Q
rlabel metal2 12288 68334 12288 68334 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame4_bit0.Q
rlabel via2 13832 68376 13832 68376 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame4_bit1.Q
rlabel metal2 16560 80472 16560 80472 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame4_bit10.Q
rlabel metal2 18152 80472 18152 80472 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame4_bit11.Q
rlabel metal2 4320 64638 4320 64638 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame4_bit12.Q
rlabel metal3 5856 65310 5856 65310 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame4_bit13.Q
rlabel metal2 7256 74424 7256 74424 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame4_bit14.Q
rlabel metal2 5760 74466 5760 74466 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame4_bit15.Q
rlabel metal3 16416 65856 16416 65856 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame4_bit16.Q
rlabel metal2 14688 66192 14688 66192 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame4_bit17.Q
rlabel metal2 18048 66192 18048 66192 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame4_bit18.Q
rlabel metal2 19968 66192 19968 66192 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame4_bit19.Q
rlabel via1 18216 56280 18216 56280 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame4_bit2.Q
rlabel metal2 3408 60816 3408 60816 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame4_bit20.Q
rlabel metal3 5568 60564 5568 60564 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame4_bit21.Q
rlabel metal3 7872 71946 7872 71946 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame4_bit22.Q
rlabel metal2 6225 72240 6225 72240 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame4_bit23.Q
rlabel metal2 15696 69216 15696 69216 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame4_bit24.Q
rlabel metal2 14256 69216 14256 69216 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame4_bit25.Q
rlabel metal2 17952 61572 17952 61572 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame4_bit26.Q
rlabel metal2 16464 61068 16464 61068 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame4_bit27.Q
rlabel metal3 7392 62076 7392 62076 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame4_bit28.Q
rlabel via1 5758 62328 5758 62328 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame4_bit29.Q
rlabel metal2 19776 56385 19776 56385 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame4_bit3.Q
rlabel metal2 10032 62412 10032 62412 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame4_bit30.Q
rlabel metal2 11640 62328 11640 62328 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame4_bit31.Q
rlabel metal2 5856 59262 5856 59262 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame4_bit4.Q
rlabel metal2 7352 59304 7352 59304 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame4_bit5.Q
rlabel metal2 7104 66780 7104 66780 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame4_bit6.Q
rlabel metal2 9672 68376 9672 68376 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame4_bit7.Q
rlabel metal2 15288 70896 15288 70896 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame4_bit8.Q
rlabel metal2 16680 71400 16680 71400 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame4_bit9.Q
rlabel metal2 14880 61824 14880 61824 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame5_bit0.Q
rlabel metal2 16184 62328 16184 62328 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame5_bit1.Q
rlabel metal2 18336 57750 18336 57750 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame5_bit10.Q
rlabel metal2 20040 57792 20040 57792 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame5_bit11.Q
rlabel metal2 4560 57120 4560 57120 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame5_bit12.Q
rlabel metal3 6432 57372 6432 57372 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame5_bit13.Q
rlabel metal2 3408 68376 3408 68376 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame5_bit14.Q
rlabel metal2 5592 68376 5592 68376 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame5_bit15.Q
rlabel metal3 13536 63924 13536 63924 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame5_bit16.Q
rlabel metal2 14168 65352 14168 65352 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame5_bit17.Q
rlabel metal2 18432 59262 18432 59262 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame5_bit18.Q
rlabel metal2 20088 59304 20088 59304 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame5_bit19.Q
rlabel metal2 18336 54138 18336 54138 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame5_bit2.Q
rlabel metal2 3552 57750 3552 57750 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame5_bit20.Q
rlabel metal2 5088 57897 5088 57897 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame5_bit21.Q
rlabel metal2 4416 70770 4416 70770 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame5_bit22.Q
rlabel metal2 6000 70728 6000 70728 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame5_bit23.Q
rlabel metal2 15105 65352 15105 65352 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame5_bit24.Q
rlabel via2 16712 65352 16712 65352 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame5_bit25.Q
rlabel metal2 18288 61656 18288 61656 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame5_bit26.Q
rlabel metal2 20016 61656 20016 61656 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame5_bit27.Q
rlabel metal2 3216 62328 3216 62328 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame5_bit28.Q
rlabel metal2 5208 62328 5208 62328 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame5_bit29.Q
rlabel metal3 19872 54726 19872 54726 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame5_bit3.Q
rlabel metal3 2688 73248 2688 73248 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame5_bit30.Q
rlabel metal2 3552 73500 3552 73500 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame5_bit31.Q
rlabel metal2 2304 58674 2304 58674 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame5_bit4.Q
rlabel metal3 3840 58926 3840 58926 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame5_bit5.Q
rlabel metal2 2928 72744 2928 72744 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame5_bit6.Q
rlabel metal2 4512 69216 4512 69216 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame5_bit7.Q
rlabel metal2 14304 67536 14304 67536 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame5_bit8.Q
rlabel metal2 16328 68376 16328 68376 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame5_bit9.Q
rlabel metal2 19896 66864 19896 66864 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame6_bit0.Q
rlabel metal2 18144 66906 18144 66906 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame6_bit1.Q
rlabel metal2 18081 63168 18081 63168 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame6_bit10.Q
rlabel metal2 19968 63168 19968 63168 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame6_bit11.Q
rlabel metal2 3552 56238 3552 56238 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame6_bit12.Q
rlabel metal3 5376 56028 5376 56028 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame6_bit13.Q
rlabel metal3 2784 68334 2784 68334 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame6_bit14.Q
rlabel metal3 4608 68712 4608 68712 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame6_bit15.Q
rlabel metal3 13632 62496 13632 62496 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame6_bit16.Q
rlabel metal2 15360 63126 15360 63126 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame6_bit17.Q
rlabel metal2 18720 52752 18720 52752 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame6_bit18.Q
rlabel metal2 20160 54936 20160 54936 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame6_bit19.Q
rlabel metal2 12680 66864 12680 66864 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame6_bit2.Q
rlabel metal2 2208 60186 2208 60186 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame6_bit20.Q
rlabel metal2 3648 60144 3648 60144 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame6_bit21.Q
rlabel metal2 2625 66192 2625 66192 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame6_bit22.Q
rlabel metal3 4224 66444 4224 66444 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame6_bit23.Q
rlabel metal2 15168 54138 15168 54138 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame6_bit24.Q
rlabel metal2 15984 53508 15984 53508 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame6_bit25.Q
rlabel metal2 18000 63840 18000 63840 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame6_bit26.Q
rlabel metal2 19738 63840 19738 63840 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame6_bit27.Q
rlabel metal2 3393 61656 3393 61656 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame6_bit28.Q
rlabel metal2 5232 61656 5232 61656 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame6_bit29.Q
rlabel metal2 11088 66864 11088 66864 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame6_bit3.Q
rlabel metal2 2817 71400 2817 71400 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame6_bit30.Q
rlabel metal2 4280 71400 4280 71400 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame6_bit31.Q
rlabel metal3 4608 75516 4608 75516 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame6_bit4.Q
rlabel metal2 3072 73794 3072 73794 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame6_bit5.Q
rlabel metal2 5568 63378 5568 63378 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame6_bit6.Q
rlabel metal3 2688 65688 2688 65688 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame6_bit7.Q
rlabel metal2 15600 52752 15600 52752 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame6_bit8.Q
rlabel metal2 17232 52752 17232 52752 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame6_bit9.Q
rlabel metal2 7776 79842 7776 79842 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit0.Q
rlabel metal2 9312 79842 9312 79842 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit1.Q
rlabel metal2 9024 51030 9024 51030 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit10.Q
rlabel metal2 13248 51450 13248 51450 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit11.Q
rlabel metal2 12768 73794 12768 73794 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit12.Q
rlabel metal2 14256 73752 14256 73752 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit13.Q
rlabel metal2 14976 75306 14976 75306 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit14.Q
rlabel metal2 12240 74676 12240 74676 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit15.Q
rlabel metal2 7488 78960 7488 78960 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit16.Q
rlabel via1 9224 78960 9224 78960 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit17.Q
rlabel metal2 9525 51744 9525 51744 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit18.Q
rlabel metal2 11664 53256 11664 53256 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit19.Q
rlabel metal2 8880 73500 8880 73500 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit2.Q
rlabel metal3 10944 52206 10944 52206 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit20.Q
rlabel metal2 16203 57792 16203 57792 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit21.Q
rlabel metal2 15552 59556 15552 59556 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit22.Q
rlabel metal2 17184 59136 17184 59136 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit23.Q
rlabel metal2 15416 81984 15416 81984 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit24.Q
rlabel metal2 13488 81984 13488 81984 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit25.Q
rlabel metal2 16992 81354 16992 81354 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit26.Q
rlabel metal3 8352 83664 8352 83664 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit27.Q
rlabel via2 5856 83496 5856 83496 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit28.Q
rlabel metal3 8064 84336 8064 84336 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit29.Q
rlabel metal2 7296 72828 7296 72828 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit3.Q
rlabel metal2 12336 59346 12336 59346 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit30.Q
rlabel metal2 10752 59346 10752 59346 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit31.Q
rlabel metal2 15264 78204 15264 78204 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit4.Q
rlabel metal2 12096 77700 12096 77700 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit5.Q
rlabel metal2 11712 70770 11712 70770 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit6.Q
rlabel metal2 13248 70686 13248 70686 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit7.Q
rlabel metal2 9183 69888 9183 69888 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit8.Q
rlabel metal3 7200 70182 7200 70182 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit9.Q
rlabel metal2 15552 77490 15552 77490 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit0.Q
rlabel metal2 17136 77406 17136 77406 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit1.Q
rlabel metal2 17952 74466 17952 74466 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit10.Q
rlabel metal2 19752 74424 19752 74424 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit11.Q
rlabel metal3 8352 76440 8352 76440 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit12.Q
rlabel metal3 9888 76482 9888 76482 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit13.Q
rlabel metal3 8544 64932 8544 64932 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit14.Q
rlabel metal2 9432 62328 9432 62328 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit15.Q
rlabel metal2 9120 63210 9120 63210 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit16.Q
rlabel metal2 19872 78330 19872 78330 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit17.Q
rlabel metal2 20208 78288 20208 78288 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit18.Q
rlabel metal2 19968 79086 19968 79086 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit19.Q
rlabel metal2 11856 71400 11856 71400 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit2.Q
rlabel metal2 13344 84378 13344 84378 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit20.Q
rlabel metal2 13536 85890 13536 85890 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit21.Q
rlabel metal2 12720 84336 12720 84336 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit22.Q
rlabel metal2 6816 81312 6816 81312 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit23.Q
rlabel metal2 7008 82026 7008 82026 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit24.Q
rlabel metal3 7488 80808 7488 80808 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit25.Q
rlabel metal2 9816 60816 9816 60816 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit26.Q
rlabel metal2 8064 60774 8064 60774 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit27.Q
rlabel metal2 13296 76776 13296 76776 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit28.Q
rlabel metal2 14952 76776 14952 76776 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit29.Q
rlabel metal2 13496 71400 13496 71400 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit3.Q
rlabel metal2 13745 75978 13745 75978 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit30.Q
rlabel metal3 12192 76608 12192 76608 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit31.Q
rlabel metal2 7104 67158 7104 67158 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit4.Q
rlabel metal2 8760 66864 8760 66864 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit5.Q
rlabel metal2 2688 53004 2688 53004 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit6.Q
rlabel metal2 3888 53928 3888 53928 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit7.Q
rlabel metal2 12720 72912 12720 72912 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit8.Q
rlabel metal2 14880 72408 14880 72408 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit9.Q
rlabel metal3 9312 57372 9312 57372 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame9_bit22.Q
rlabel metal2 7968 56532 7968 56532 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame9_bit23.Q
rlabel metal2 14400 74466 14400 74466 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame9_bit24.Q
rlabel metal2 15752 74424 15752 74424 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame9_bit25.Q
rlabel metal2 13824 78456 13824 78456 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame9_bit26.Q
rlabel metal2 15272 78960 15272 78960 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame9_bit27.Q
rlabel metal2 7425 86520 7425 86520 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame9_bit28.Q
rlabel metal2 8840 86520 8840 86520 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame9_bit29.Q
rlabel via1 8546 73752 8546 73752 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame9_bit30.Q
rlabel metal2 7104 73752 7104 73752 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame9_bit31.Q
rlabel metal3 6912 70056 6912 70056 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS2_BEG0
rlabel metal4 17616 60060 17616 60060 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS2_BEG1
rlabel metal3 13440 58296 13440 58296 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS2_BEG2
rlabel metal2 5808 55524 5808 55524 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS2_BEG3
rlabel metal2 4944 47040 4944 47040 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS2_BEG4
rlabel metal2 15264 60060 15264 60060 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS2_BEG5
rlabel metal2 16464 60480 16464 60480 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS2_BEG6
rlabel metal3 9024 62916 9024 62916 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS2_BEG7
rlabel metal2 11064 54852 11064 54852 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG0
rlabel metal2 16704 58632 16704 58632 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG1
rlabel metal2 15264 82782 15264 82782 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG10
rlabel metal2 4320 68376 4320 68376 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG11
rlabel metal4 8496 63252 8496 63252 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG12
rlabel metal2 19392 69678 19392 69678 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG13
rlabel via2 14699 82740 14699 82740 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG14
rlabel metal2 3936 69132 3936 69132 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG15
rlabel metal2 14496 81900 14496 81900 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG2
rlabel metal3 4320 82950 4320 82950 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG3
rlabel metal2 6240 62496 6240 62496 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG4
rlabel metal2 16416 56322 16416 56322 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG5
rlabel metal2 13968 81480 13968 81480 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG6
rlabel metal2 5904 87360 5904 87360 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG7
rlabel metal2 10320 53424 10320 53424 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG8
rlabel metal2 19056 59304 19056 59304 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG9
rlabel metal2 9768 56868 9768 56868 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.N1BEG0
rlabel metal2 15792 73668 15792 73668 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.N1BEG1
rlabel metal2 15768 79044 15768 79044 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.N1BEG2
rlabel metal2 9096 86772 9096 86772 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.N1BEG3
rlabel metal2 8880 36540 8880 36540 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.N1END0
rlabel metal4 17424 56112 17424 56112 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.N1END1
rlabel metal2 12336 36456 12336 36456 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.N1END2
rlabel metal3 9360 61740 9360 61740 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.N1END3
rlabel metal2 8448 74466 8448 74466 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.N2BEG0
rlabel metal3 17280 78498 17280 78498 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.N2BEG1
rlabel metal2 13944 71484 13944 71484 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.N2BEG2
rlabel metal2 9216 66864 9216 66864 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.N2BEG3
rlabel metal2 4752 51828 4752 51828 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.N2BEG4
rlabel metal2 14784 73668 14784 73668 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.N2BEG5
rlabel metal2 19392 74256 19392 74256 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.N2BEG6
rlabel metal2 10296 76692 10296 76692 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.N2BEG7
rlabel metal2 4656 41244 4656 41244 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.N2BEGb0
rlabel metal2 15504 31920 15504 31920 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.N2BEGb1
rlabel metal3 12672 41874 12672 41874 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.N2BEGb2
rlabel metal2 4128 46410 4128 46410 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.N2BEGb3
rlabel metal2 3552 46452 3552 46452 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.N2BEGb4
rlabel metal2 19872 41244 19872 41244 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.N2BEGb5
rlabel metal2 16944 31332 16944 31332 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.N2BEGb6
rlabel metal2 9120 40404 9120 40404 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.N2BEGb7
rlabel metal2 9600 63336 9600 63336 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.N4BEG0
rlabel metal4 19488 82404 19488 82404 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.N4BEG1
rlabel metal2 14208 83622 14208 83622 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.N4BEG2
rlabel metal2 8544 81228 8544 81228 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.N4BEG3
rlabel metal4 4368 43092 4368 43092 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.S2BEG0
rlabel metal4 17040 57624 17040 57624 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.S2BEG1
rlabel metal3 11280 58296 11280 58296 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.S2BEG2
rlabel metal2 6000 42000 6000 42000 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.S2BEG3
rlabel metal3 2784 50190 2784 50190 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.S2BEG4
rlabel metal3 17616 56112 17616 56112 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.S2BEG5
rlabel metal2 16656 75432 16656 75432 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.S2BEG6
rlabel metal2 9408 78708 9408 78708 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.S2BEG7
rlabel metal2 10704 52752 10704 52752 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.S4BEG0
rlabel metal3 18432 59220 18432 59220 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.S4BEG1
rlabel metal2 16176 82656 16176 82656 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.S4BEG2
rlabel metal2 8448 84546 8448 84546 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.S4BEG3
rlabel metal2 12696 59388 12696 59388 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.W1BEG0
rlabel metal2 19824 66696 19824 66696 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.W1BEG1
rlabel metal3 13056 66402 13056 66402 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.W1BEG2
rlabel metal3 5568 74970 5568 74970 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.W1BEG3
rlabel metal2 3840 64806 3840 64806 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.W2BEG0
rlabel metal2 18048 53382 18048 53382 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.W2BEG1
rlabel metal2 19344 63336 19344 63336 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.W2BEG2
rlabel metal2 5496 56364 5496 56364 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.W2BEG3
rlabel metal2 3552 70014 3552 70014 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.W2BEG4
rlabel metal2 15648 63336 15648 63336 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.W2BEG5
rlabel metal3 19680 52794 19680 52794 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.W2BEG6
rlabel metal2 3768 59892 3768 59892 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.W2BEG7
rlabel metal2 4992 67620 4992 67620 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.W2BEGb0
rlabel metal2 17112 54012 17112 54012 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.W2BEGb1
rlabel metal3 19872 66066 19872 66066 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.W2BEGb2
rlabel via1 5208 61404 5208 61404 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.W2BEGb3
rlabel metal2 5184 71232 5184 71232 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.W2BEGb4
rlabel metal2 15792 61572 15792 61572 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.W2BEGb5
rlabel metal2 18048 54138 18048 54138 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.W2BEGb6
rlabel metal3 3936 59094 3936 59094 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.W2BEGb7
rlabel metal2 9600 68250 9600 68250 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.W6BEG0
rlabel metal2 16560 70644 16560 70644 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.W6BEG1
rlabel metal2 17760 61824 17760 61824 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.W6BEG10
rlabel metal3 7776 61866 7776 61866 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.W6BEG11
rlabel metal3 18432 83034 18432 83034 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.W6BEG2
rlabel metal2 6264 64596 6264 64596 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.W6BEG3
rlabel metal3 7488 75138 7488 75138 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.W6BEG4
rlabel metal2 16824 66108 16824 66108 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.W6BEG5
rlabel metal3 18624 68334 18624 68334 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.W6BEG6
rlabel metal2 5592 60900 5592 60900 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.W6BEG7
rlabel metal2 8280 72156 8280 72156 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.W6BEG8
rlabel metal2 16248 69972 16248 69972 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.W6BEG9
rlabel metal2 6192 70644 6192 70644 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.WW4BEG0
rlabel metal3 16608 68670 16608 68670 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.WW4BEG1
rlabel metal2 20448 61824 20448 61824 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.WW4BEG10
rlabel metal3 5568 61866 5568 61866 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.WW4BEG11
rlabel metal2 5376 72198 5376 72198 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.WW4BEG12
rlabel metal2 14232 68460 14232 68460 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.WW4BEG13
rlabel metal2 17568 56238 17568 56238 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.WW4BEG14
rlabel metal2 8448 59346 8448 59346 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.WW4BEG15
rlabel metal2 15408 57876 15408 57876 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.WW4BEG2
rlabel metal2 6840 57036 6840 57036 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.WW4BEG3
rlabel metal3 5568 68670 5568 68670 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.WW4BEG4
rlabel metal2 14616 65436 14616 65436 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.WW4BEG5
rlabel metal2 20160 59094 20160 59094 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.WW4BEG6
rlabel metal2 5448 58044 5448 58044 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.WW4BEG7
rlabel metal2 6720 70644 6720 70644 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.WW4BEG8
rlabel metal2 17160 65604 17160 65604 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.WW4BEG9
rlabel metal2 17760 36120 17760 36120 0 Tile_X0Y0_IHP_SRAM_top.N4BEG_outbuf_10.A
rlabel metal2 15456 35700 15456 35700 0 Tile_X0Y0_IHP_SRAM_top.N4BEG_outbuf_11.A
rlabel metal2 5328 28308 5328 28308 0 Tile_X0Y0_IHP_SRAM_top.N4BEG_outbuf_8.A
rlabel metal2 16224 20244 16224 20244 0 Tile_X0Y0_IHP_SRAM_top.N4BEG_outbuf_9.A
rlabel metal3 1824 95154 1824 95154 0 Tile_X0Y0_N1BEG[0]
rlabel metal2 2376 93576 2376 93576 0 Tile_X0Y0_N1BEG[1]
rlabel metal2 2040 94248 2040 94248 0 Tile_X0Y0_N1BEG[2]
rlabel metal2 2328 94332 2328 94332 0 Tile_X0Y0_N1BEG[3]
rlabel metal2 2088 95004 2088 95004 0 Tile_X0Y0_N2BEG[0]
rlabel metal2 2712 94332 2712 94332 0 Tile_X0Y0_N2BEG[1]
rlabel metal3 2976 95730 2976 95730 0 Tile_X0Y0_N2BEG[2]
rlabel metal2 2616 94668 2616 94668 0 Tile_X0Y0_N2BEG[3]
rlabel metal3 3360 95856 3360 95856 0 Tile_X0Y0_N2BEG[4]
rlabel metal2 3576 94332 3576 94332 0 Tile_X0Y0_N2BEG[5]
rlabel metal2 3432 94752 3432 94752 0 Tile_X0Y0_N2BEG[6]
rlabel metal2 4056 94332 4056 94332 0 Tile_X0Y0_N2BEG[7]
rlabel metal2 3864 95004 3864 95004 0 Tile_X0Y0_N2BEGb[0]
rlabel metal2 4344 94332 4344 94332 0 Tile_X0Y0_N2BEGb[1]
rlabel metal2 4200 94752 4200 94752 0 Tile_X0Y0_N2BEGb[2]
rlabel metal2 4728 94332 4728 94332 0 Tile_X0Y0_N2BEGb[3]
rlabel metal2 4392 94668 4392 94668 0 Tile_X0Y0_N2BEGb[4]
rlabel metal2 5256 94332 5256 94332 0 Tile_X0Y0_N2BEGb[5]
rlabel metal2 4632 95004 4632 95004 0 Tile_X0Y0_N2BEGb[6]
rlabel metal2 5496 94248 5496 94248 0 Tile_X0Y0_N2BEGb[7]
rlabel metal2 5352 95004 5352 95004 0 Tile_X0Y0_N4BEG[0]
rlabel metal2 7272 95004 7272 95004 0 Tile_X0Y0_N4BEG[10]
rlabel metal2 7800 94332 7800 94332 0 Tile_X0Y0_N4BEG[11]
rlabel metal2 7512 95088 7512 95088 0 Tile_X0Y0_N4BEG[12]
rlabel metal2 7944 94752 7944 94752 0 Tile_X0Y0_N4BEG[13]
rlabel metal2 8232 95004 8232 95004 0 Tile_X0Y0_N4BEG[14]
rlabel metal2 8568 94332 8568 94332 0 Tile_X0Y0_N4BEG[15]
rlabel metal2 5880 94332 5880 94332 0 Tile_X0Y0_N4BEG[1]
rlabel metal2 5736 94752 5736 94752 0 Tile_X0Y0_N4BEG[2]
rlabel metal2 6264 94332 6264 94332 0 Tile_X0Y0_N4BEG[3]
rlabel metal2 6120 95004 6120 95004 0 Tile_X0Y0_N4BEG[4]
rlabel metal2 6648 94332 6648 94332 0 Tile_X0Y0_N4BEG[5]
rlabel metal2 6504 94752 6504 94752 0 Tile_X0Y0_N4BEG[6]
rlabel metal2 7032 94332 7032 94332 0 Tile_X0Y0_N4BEG[7]
rlabel metal2 6888 94668 6888 94668 0 Tile_X0Y0_N4BEG[8]
rlabel metal2 7416 94332 7416 94332 0 Tile_X0Y0_N4BEG[9]
rlabel metal3 8736 95814 8736 95814 0 Tile_X0Y0_S1END[0]
rlabel metal3 8928 95478 8928 95478 0 Tile_X0Y0_S1END[1]
rlabel metal3 9120 95814 9120 95814 0 Tile_X0Y0_S1END[2]
rlabel metal3 9312 95436 9312 95436 0 Tile_X0Y0_S1END[3]
rlabel metal3 11040 95814 11040 95814 0 Tile_X0Y0_S2END[0]
rlabel metal3 11232 95814 11232 95814 0 Tile_X0Y0_S2END[1]
rlabel metal3 11424 95772 11424 95772 0 Tile_X0Y0_S2END[2]
rlabel metal3 11616 95772 11616 95772 0 Tile_X0Y0_S2END[3]
rlabel metal3 11808 95730 11808 95730 0 Tile_X0Y0_S2END[4]
rlabel metal3 12000 95814 12000 95814 0 Tile_X0Y0_S2END[5]
rlabel metal3 12192 95814 12192 95814 0 Tile_X0Y0_S2END[6]
rlabel metal2 13440 94710 13440 94710 0 Tile_X0Y0_S2END[7]
rlabel metal3 9504 95814 9504 95814 0 Tile_X0Y0_S2MID[0]
rlabel metal3 9696 95478 9696 95478 0 Tile_X0Y0_S2MID[1]
rlabel metal3 9888 95814 9888 95814 0 Tile_X0Y0_S2MID[2]
rlabel metal3 10080 95436 10080 95436 0 Tile_X0Y0_S2MID[3]
rlabel metal3 10272 95814 10272 95814 0 Tile_X0Y0_S2MID[4]
rlabel metal3 10464 95478 10464 95478 0 Tile_X0Y0_S2MID[5]
rlabel metal3 10656 95814 10656 95814 0 Tile_X0Y0_S2MID[6]
rlabel metal3 10848 95436 10848 95436 0 Tile_X0Y0_S2MID[7]
rlabel metal3 12576 95436 12576 95436 0 Tile_X0Y0_S4END[0]
rlabel metal3 14496 95478 14496 95478 0 Tile_X0Y0_S4END[10]
rlabel metal3 14688 96654 14688 96654 0 Tile_X0Y0_S4END[11]
rlabel metal2 17952 94122 17952 94122 0 Tile_X0Y0_S4END[12]
rlabel metal3 15072 95478 15072 95478 0 Tile_X0Y0_S4END[13]
rlabel metal3 15264 95436 15264 95436 0 Tile_X0Y0_S4END[14]
rlabel metal3 15456 96192 15456 96192 0 Tile_X0Y0_S4END[15]
rlabel metal2 13632 94920 13632 94920 0 Tile_X0Y0_S4END[1]
rlabel metal2 13008 94164 13008 94164 0 Tile_X0Y0_S4END[2]
rlabel metal3 13152 95814 13152 95814 0 Tile_X0Y0_S4END[3]
rlabel metal3 13344 95436 13344 95436 0 Tile_X0Y0_S4END[4]
rlabel metal3 13536 95898 13536 95898 0 Tile_X0Y0_S4END[5]
rlabel metal3 13728 95478 13728 95478 0 Tile_X0Y0_S4END[6]
rlabel metal3 13920 95646 13920 95646 0 Tile_X0Y0_S4END[7]
rlabel metal3 14112 95436 14112 95436 0 Tile_X0Y0_S4END[8]
rlabel metal3 14304 96318 14304 96318 0 Tile_X0Y0_S4END[9]
rlabel metal2 15672 95004 15672 95004 0 Tile_X0Y0_UserCLKo
rlabel metal2 320 51156 320 51156 0 Tile_X0Y0_W1BEG[0]
rlabel metal2 704 51492 704 51492 0 Tile_X0Y0_W1BEG[1]
rlabel metal2 888 53340 888 53340 0 Tile_X0Y0_W1BEG[2]
rlabel metal2 128 52164 128 52164 0 Tile_X0Y0_W1BEG[3]
rlabel metal2 368 52500 368 52500 0 Tile_X0Y0_W2BEG[0]
rlabel metal2 936 53844 936 53844 0 Tile_X0Y0_W2BEG[1]
rlabel metal2 704 53172 704 53172 0 Tile_X0Y0_W2BEG[2]
rlabel metal2 320 53508 320 53508 0 Tile_X0Y0_W2BEG[3]
rlabel metal2 272 53844 272 53844 0 Tile_X0Y0_W2BEG[4]
rlabel metal2 704 54180 704 54180 0 Tile_X0Y0_W2BEG[5]
rlabel metal2 1424 54516 1424 54516 0 Tile_X0Y0_W2BEG[6]
rlabel metal2 944 54852 944 54852 0 Tile_X0Y0_W2BEG[7]
rlabel metal2 368 55188 368 55188 0 Tile_X0Y0_W2BEGb[0]
rlabel metal2 752 55524 752 55524 0 Tile_X0Y0_W2BEGb[1]
rlabel metal2 416 55860 416 55860 0 Tile_X0Y0_W2BEGb[2]
rlabel metal2 128 56196 128 56196 0 Tile_X0Y0_W2BEGb[3]
rlabel via2 80 56532 80 56532 0 Tile_X0Y0_W2BEGb[4]
rlabel metal2 176 56868 176 56868 0 Tile_X0Y0_W2BEGb[5]
rlabel metal2 128 57204 128 57204 0 Tile_X0Y0_W2BEGb[6]
rlabel metal2 800 57540 800 57540 0 Tile_X0Y0_W2BEGb[7]
rlabel metal2 656 63252 656 63252 0 Tile_X0Y0_W6BEG[0]
rlabel metal2 512 66612 512 66612 0 Tile_X0Y0_W6BEG[10]
rlabel metal2 128 66948 128 66948 0 Tile_X0Y0_W6BEG[11]
rlabel metal2 656 63588 656 63588 0 Tile_X0Y0_W6BEG[1]
rlabel metal2 416 63924 416 63924 0 Tile_X0Y0_W6BEG[2]
rlabel metal2 608 64260 608 64260 0 Tile_X0Y0_W6BEG[3]
rlabel metal2 656 64596 656 64596 0 Tile_X0Y0_W6BEG[4]
rlabel metal2 320 64932 320 64932 0 Tile_X0Y0_W6BEG[5]
rlabel metal2 224 65268 224 65268 0 Tile_X0Y0_W6BEG[6]
rlabel metal2 176 65604 176 65604 0 Tile_X0Y0_W6BEG[7]
rlabel metal2 272 65940 272 65940 0 Tile_X0Y0_W6BEG[8]
rlabel metal2 656 66276 656 66276 0 Tile_X0Y0_W6BEG[9]
rlabel metal2 752 57876 752 57876 0 Tile_X0Y0_WW4BEG[0]
rlabel metal2 1040 61236 1040 61236 0 Tile_X0Y0_WW4BEG[10]
rlabel metal2 368 61572 368 61572 0 Tile_X0Y0_WW4BEG[11]
rlabel metal2 560 61908 560 61908 0 Tile_X0Y0_WW4BEG[12]
rlabel metal2 848 62244 848 62244 0 Tile_X0Y0_WW4BEG[13]
rlabel metal2 752 62580 752 62580 0 Tile_X0Y0_WW4BEG[14]
rlabel metal2 224 62916 224 62916 0 Tile_X0Y0_WW4BEG[15]
rlabel metal2 272 58212 272 58212 0 Tile_X0Y0_WW4BEG[1]
rlabel metal2 704 58548 704 58548 0 Tile_X0Y0_WW4BEG[2]
rlabel metal2 320 58884 320 58884 0 Tile_X0Y0_WW4BEG[3]
rlabel metal2 944 59220 944 59220 0 Tile_X0Y0_WW4BEG[4]
rlabel metal2 992 59556 992 59556 0 Tile_X0Y0_WW4BEG[5]
rlabel metal2 128 59892 128 59892 0 Tile_X0Y0_WW4BEG[6]
rlabel metal2 704 60228 704 60228 0 Tile_X0Y0_WW4BEG[7]
rlabel metal2 512 60564 512 60564 0 Tile_X0Y0_WW4BEG[8]
rlabel metal2 848 60900 848 60900 0 Tile_X0Y0_WW4BEG[9]
rlabel metal2 1808 18900 1808 18900 0 Tile_X0Y1_E1END[0]
rlabel metal2 416 19236 416 19236 0 Tile_X0Y1_E1END[1]
rlabel metal2 272 19572 272 19572 0 Tile_X0Y1_E1END[2]
rlabel metal2 464 19908 464 19908 0 Tile_X0Y1_E1END[3]
rlabel metal2 11232 22974 11232 22974 0 Tile_X0Y1_E2END[0]
rlabel metal2 80 23268 80 23268 0 Tile_X0Y1_E2END[1]
rlabel metal2 10656 23226 10656 23226 0 Tile_X0Y1_E2END[2]
rlabel metal2 1152 16212 1152 16212 0 Tile_X0Y1_E2END[3]
rlabel metal2 10080 24024 10080 24024 0 Tile_X0Y1_E2END[4]
rlabel metal2 960 17724 960 17724 0 Tile_X0Y1_E2END[5]
rlabel metal2 1808 24948 1808 24948 0 Tile_X0Y1_E2END[6]
rlabel metal2 912 18396 912 18396 0 Tile_X0Y1_E2END[7]
rlabel metal2 1472 20244 1472 20244 0 Tile_X0Y1_E2MID[0]
rlabel metal2 1472 20580 1472 20580 0 Tile_X0Y1_E2MID[1]
rlabel metal2 512 20916 512 20916 0 Tile_X0Y1_E2MID[2]
rlabel metal2 80 21252 80 21252 0 Tile_X0Y1_E2MID[3]
rlabel metal2 512 21588 512 21588 0 Tile_X0Y1_E2MID[4]
rlabel metal2 752 21924 752 21924 0 Tile_X0Y1_E2MID[5]
rlabel metal2 128 22260 128 22260 0 Tile_X0Y1_E2MID[6]
rlabel metal3 5856 20496 5856 20496 0 Tile_X0Y1_E2MID[7]
rlabel metal2 1136 30996 1136 30996 0 Tile_X0Y1_E6END[0]
rlabel metal2 272 34356 272 34356 0 Tile_X0Y1_E6END[10]
rlabel metal2 848 34692 848 34692 0 Tile_X0Y1_E6END[11]
rlabel metal2 368 31332 368 31332 0 Tile_X0Y1_E6END[1]
rlabel metal2 128 31668 128 31668 0 Tile_X0Y1_E6END[2]
rlabel metal2 656 32004 656 32004 0 Tile_X0Y1_E6END[3]
rlabel metal2 1808 32340 1808 32340 0 Tile_X0Y1_E6END[4]
rlabel via2 80 32676 80 32676 0 Tile_X0Y1_E6END[5]
rlabel via2 80 33012 80 33012 0 Tile_X0Y1_E6END[6]
rlabel metal2 176 33348 176 33348 0 Tile_X0Y1_E6END[7]
rlabel metal2 1040 33684 1040 33684 0 Tile_X0Y1_E6END[8]
rlabel metal2 848 34020 848 34020 0 Tile_X0Y1_E6END[9]
rlabel metal2 1104 18480 1104 18480 0 Tile_X0Y1_EE4END[0]
rlabel metal2 2976 28896 2976 28896 0 Tile_X0Y1_EE4END[10]
rlabel metal2 704 29316 704 29316 0 Tile_X0Y1_EE4END[11]
rlabel via2 80 29652 80 29652 0 Tile_X0Y1_EE4END[12]
rlabel metal2 1056 22260 1056 22260 0 Tile_X0Y1_EE4END[13]
rlabel metal2 11424 30534 11424 30534 0 Tile_X0Y1_EE4END[14]
rlabel metal2 416 30660 416 30660 0 Tile_X0Y1_EE4END[15]
rlabel metal2 1296 18564 1296 18564 0 Tile_X0Y1_EE4END[1]
rlabel metal2 3600 22512 3600 22512 0 Tile_X0Y1_EE4END[2]
rlabel metal2 176 26628 176 26628 0 Tile_X0Y1_EE4END[3]
rlabel metal2 272 26964 272 26964 0 Tile_X0Y1_EE4END[4]
rlabel metal3 6528 27132 6528 27132 0 Tile_X0Y1_EE4END[5]
rlabel metal2 128 27636 128 27636 0 Tile_X0Y1_EE4END[6]
rlabel metal2 1040 27972 1040 27972 0 Tile_X0Y1_EE4END[7]
rlabel metal2 272 28308 272 28308 0 Tile_X0Y1_EE4END[8]
rlabel metal3 1248 22314 1248 22314 0 Tile_X0Y1_EE4END[9]
rlabel metal2 704 35028 704 35028 0 Tile_X0Y1_FrameData[0]
rlabel metal2 752 38388 752 38388 0 Tile_X0Y1_FrameData[10]
rlabel metal2 848 38724 848 38724 0 Tile_X0Y1_FrameData[11]
rlabel metal2 656 39060 656 39060 0 Tile_X0Y1_FrameData[12]
rlabel metal2 704 39396 704 39396 0 Tile_X0Y1_FrameData[13]
rlabel metal2 464 39732 464 39732 0 Tile_X0Y1_FrameData[14]
rlabel metal2 224 40068 224 40068 0 Tile_X0Y1_FrameData[15]
rlabel metal2 80 40404 80 40404 0 Tile_X0Y1_FrameData[16]
rlabel metal2 656 40740 656 40740 0 Tile_X0Y1_FrameData[17]
rlabel via2 80 41076 80 41076 0 Tile_X0Y1_FrameData[18]
rlabel metal2 848 41412 848 41412 0 Tile_X0Y1_FrameData[19]
rlabel metal2 128 35364 128 35364 0 Tile_X0Y1_FrameData[1]
rlabel metal2 128 41748 128 41748 0 Tile_X0Y1_FrameData[20]
rlabel metal2 128 42084 128 42084 0 Tile_X0Y1_FrameData[21]
rlabel metal2 128 42420 128 42420 0 Tile_X0Y1_FrameData[22]
rlabel metal2 656 42756 656 42756 0 Tile_X0Y1_FrameData[23]
rlabel metal2 848 43092 848 43092 0 Tile_X0Y1_FrameData[24]
rlabel metal2 656 43428 656 43428 0 Tile_X0Y1_FrameData[25]
rlabel metal2 128 43764 128 43764 0 Tile_X0Y1_FrameData[26]
rlabel via2 80 44100 80 44100 0 Tile_X0Y1_FrameData[27]
rlabel metal2 848 44436 848 44436 0 Tile_X0Y1_FrameData[28]
rlabel via2 80 44772 80 44772 0 Tile_X0Y1_FrameData[29]
rlabel metal2 464 35700 464 35700 0 Tile_X0Y1_FrameData[2]
rlabel metal2 848 45108 848 45108 0 Tile_X0Y1_FrameData[30]
rlabel via2 80 45444 80 45444 0 Tile_X0Y1_FrameData[31]
rlabel metal2 656 36036 656 36036 0 Tile_X0Y1_FrameData[3]
rlabel metal2 752 36372 752 36372 0 Tile_X0Y1_FrameData[4]
rlabel metal2 368 36708 368 36708 0 Tile_X0Y1_FrameData[5]
rlabel metal2 1472 37044 1472 37044 0 Tile_X0Y1_FrameData[6]
rlabel metal2 128 37380 128 37380 0 Tile_X0Y1_FrameData[7]
rlabel metal2 464 37716 464 37716 0 Tile_X0Y1_FrameData[8]
rlabel metal2 416 38052 416 38052 0 Tile_X0Y1_FrameData[9]
rlabel metal3 18624 78960 18624 78960 0 Tile_X0Y1_FrameData_O[0]
rlabel metal2 18168 85512 18168 85512 0 Tile_X0Y1_FrameData_O[10]
rlabel metal2 20847 82572 20847 82572 0 Tile_X0Y1_FrameData_O[11]
rlabel metal2 21471 83076 21471 83076 0 Tile_X0Y1_FrameData_O[12]
rlabel metal2 21471 83580 21471 83580 0 Tile_X0Y1_FrameData_O[13]
rlabel metal2 21327 84084 21327 84084 0 Tile_X0Y1_FrameData_O[14]
rlabel metal4 20448 88620 20448 88620 0 Tile_X0Y1_FrameData_O[15]
rlabel metal2 21423 85092 21423 85092 0 Tile_X0Y1_FrameData_O[16]
rlabel metal2 21375 85596 21375 85596 0 Tile_X0Y1_FrameData_O[17]
rlabel metal2 21279 86100 21279 86100 0 Tile_X0Y1_FrameData_O[18]
rlabel metal2 21423 86604 21423 86604 0 Tile_X0Y1_FrameData_O[19]
rlabel metal2 21375 77532 21375 77532 0 Tile_X0Y1_FrameData_O[1]
rlabel metal2 21135 87108 21135 87108 0 Tile_X0Y1_FrameData_O[20]
rlabel metal2 21471 87612 21471 87612 0 Tile_X0Y1_FrameData_O[21]
rlabel metal2 21183 88116 21183 88116 0 Tile_X0Y1_FrameData_O[22]
rlabel metal2 21087 88620 21087 88620 0 Tile_X0Y1_FrameData_O[23]
rlabel metal2 21279 89124 21279 89124 0 Tile_X0Y1_FrameData_O[24]
rlabel metal2 21471 89628 21471 89628 0 Tile_X0Y1_FrameData_O[25]
rlabel metal2 21135 90132 21135 90132 0 Tile_X0Y1_FrameData_O[26]
rlabel metal2 21183 90636 21183 90636 0 Tile_X0Y1_FrameData_O[27]
rlabel metal2 21471 91140 21471 91140 0 Tile_X0Y1_FrameData_O[28]
rlabel metal2 21279 91644 21279 91644 0 Tile_X0Y1_FrameData_O[29]
rlabel metal2 21231 78036 21231 78036 0 Tile_X0Y1_FrameData_O[2]
rlabel metal2 21183 92148 21183 92148 0 Tile_X0Y1_FrameData_O[30]
rlabel metal2 21279 92652 21279 92652 0 Tile_X0Y1_FrameData_O[31]
rlabel metal3 20016 83328 20016 83328 0 Tile_X0Y1_FrameData_O[3]
rlabel metal2 21183 79044 21183 79044 0 Tile_X0Y1_FrameData_O[4]
rlabel metal2 20544 79506 20544 79506 0 Tile_X0Y1_FrameData_O[5]
rlabel metal2 20928 80220 20928 80220 0 Tile_X0Y1_FrameData_O[6]
rlabel via2 21519 80556 21519 80556 0 Tile_X0Y1_FrameData_O[7]
rlabel metal2 21279 81060 21279 81060 0 Tile_X0Y1_FrameData_O[8]
rlabel metal2 19887 81564 19887 81564 0 Tile_X0Y1_FrameData_O[9]
rlabel metal3 15840 618 15840 618 0 Tile_X0Y1_FrameStrobe[0]
rlabel metal2 2592 2562 2592 2562 0 Tile_X0Y1_FrameStrobe[10]
rlabel metal3 17952 534 17952 534 0 Tile_X0Y1_FrameStrobe[11]
rlabel metal3 17376 93912 17376 93912 0 Tile_X0Y1_FrameStrobe[12]
rlabel metal3 18336 282 18336 282 0 Tile_X0Y1_FrameStrobe[13]
rlabel metal3 18528 660 18528 660 0 Tile_X0Y1_FrameStrobe[14]
rlabel metal3 18720 618 18720 618 0 Tile_X0Y1_FrameStrobe[15]
rlabel metal3 18912 702 18912 702 0 Tile_X0Y1_FrameStrobe[16]
rlabel metal3 19104 114 19104 114 0 Tile_X0Y1_FrameStrobe[17]
rlabel metal3 19296 744 19296 744 0 Tile_X0Y1_FrameStrobe[18]
rlabel metal3 19488 744 19488 744 0 Tile_X0Y1_FrameStrobe[19]
rlabel metal3 16032 660 16032 660 0 Tile_X0Y1_FrameStrobe[1]
rlabel metal3 16224 156 16224 156 0 Tile_X0Y1_FrameStrobe[2]
rlabel metal3 16416 744 16416 744 0 Tile_X0Y1_FrameStrobe[3]
rlabel metal3 16608 240 16608 240 0 Tile_X0Y1_FrameStrobe[4]
rlabel metal3 16800 702 16800 702 0 Tile_X0Y1_FrameStrobe[5]
rlabel metal3 16992 114 16992 114 0 Tile_X0Y1_FrameStrobe[6]
rlabel metal3 17184 450 17184 450 0 Tile_X0Y1_FrameStrobe[7]
rlabel metal3 17376 996 17376 996 0 Tile_X0Y1_FrameStrobe[8]
rlabel metal3 17568 198 17568 198 0 Tile_X0Y1_FrameStrobe[9]
rlabel metal3 9024 22344 9024 22344 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame0_bit0.Q
rlabel metal2 10608 22512 10608 22512 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame0_bit1.Q
rlabel metal2 15888 49728 15888 49728 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame0_bit10.Q
rlabel metal2 17472 49980 17472 49980 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame0_bit11.Q
rlabel metal2 11952 43344 11952 43344 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame0_bit12.Q
rlabel metal2 10848 43512 10848 43512 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame0_bit13.Q
rlabel metal2 6816 41958 6816 41958 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame0_bit14.Q
rlabel metal2 5280 42042 5280 42042 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame0_bit15.Q
rlabel metal2 2496 46704 2496 46704 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame0_bit16.Q
rlabel metal2 3216 47460 3216 47460 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame0_bit17.Q
rlabel metal2 18624 48216 18624 48216 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame0_bit18.Q
rlabel metal2 19592 48720 19592 48720 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame0_bit19.Q
rlabel metal2 13632 16926 13632 16926 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame0_bit2.Q
rlabel metal3 15840 47712 15840 47712 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame0_bit20.Q
rlabel metal3 17280 47754 17280 47754 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame0_bit21.Q
rlabel metal2 10032 41412 10032 41412 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame0_bit22.Q
rlabel metal3 11232 49266 11232 49266 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame0_bit23.Q
rlabel via2 7504 35112 7504 35112 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame0_bit24.Q
rlabel metal2 7632 33852 7632 33852 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame0_bit25.Q
rlabel metal2 13920 22302 13920 22302 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame0_bit26.Q
rlabel metal2 14496 22470 14496 22470 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame0_bit27.Q
rlabel metal2 9888 35658 9888 35658 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame0_bit28.Q
rlabel metal2 9696 35406 9696 35406 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame0_bit29.Q
rlabel metal2 15264 16716 15264 16716 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame0_bit3.Q
rlabel metal2 9792 45444 9792 45444 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame0_bit30.Q
rlabel metal2 10560 45192 10560 45192 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame0_bit31.Q
rlabel metal2 11841 12432 11841 12432 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame0_bit4.Q
rlabel via2 13448 12432 13448 12432 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame0_bit5.Q
rlabel metal2 9072 33516 9072 33516 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame0_bit6.Q
rlabel metal3 10944 35070 10944 35070 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame0_bit7.Q
rlabel metal2 4800 35364 4800 35364 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame0_bit8.Q
rlabel metal3 5760 37380 5760 37380 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame0_bit9.Q
rlabel metal2 5449 45024 5449 45024 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit0.Q
rlabel metal2 4896 43596 4896 43596 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit1.Q
rlabel metal2 13344 16338 13344 16338 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit10.Q
rlabel metal2 14736 15708 14736 15708 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit11.Q
rlabel metal3 11904 9156 11904 9156 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit12.Q
rlabel metal3 14304 8232 14304 8232 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit13.Q
rlabel metal2 11040 27720 11040 27720 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit14.Q
rlabel metal2 11384 29064 11384 29064 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit15.Q
rlabel metal2 7392 20874 7392 20874 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit16.Q
rlabel metal2 8880 19908 8880 19908 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit17.Q
rlabel metal2 12816 13944 12816 13944 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit18.Q
rlabel metal2 14552 13944 14552 13944 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit19.Q
rlabel metal2 6136 45696 6136 45696 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit2.Q
rlabel metal3 12096 8652 12096 8652 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit20.Q
rlabel metal3 14016 9198 14016 9198 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit21.Q
rlabel metal3 9984 31794 9984 31794 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit22.Q
rlabel metal2 11568 31584 11568 31584 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit23.Q
rlabel metal3 8160 17514 8160 17514 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit24.Q
rlabel metal2 10320 17808 10320 17808 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit25.Q
rlabel metal3 12384 14490 12384 14490 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit26.Q
rlabel metal3 14304 15246 14304 15246 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit27.Q
rlabel metal3 11808 8442 11808 8442 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit28.Q
rlabel metal3 13824 8442 13824 8442 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit29.Q
rlabel metal2 5760 46704 5760 46704 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit3.Q
rlabel metal2 9264 33600 9264 33600 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit30.Q
rlabel via2 10952 33600 10952 33600 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit31.Q
rlabel metal2 6240 41160 6240 41160 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit4.Q
rlabel metal2 6432 29316 6432 29316 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit5.Q
rlabel metal2 6432 40488 6432 40488 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit6.Q
rlabel metal2 5184 38052 5184 38052 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit7.Q
rlabel metal2 6144 22974 6144 22974 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit8.Q
rlabel metal2 8168 23016 8168 23016 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit9.Q
rlabel metal2 18912 34524 18912 34524 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit0.Q
rlabel metal2 20208 35952 20208 35952 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit1.Q
rlabel metal2 14208 45738 14208 45738 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit10.Q
rlabel metal2 15560 45696 15560 45696 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit11.Q
rlabel metal3 6816 28770 6816 28770 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit12.Q
rlabel metal2 8664 29064 8664 29064 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit13.Q
rlabel metal2 16224 22512 16224 22512 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit14.Q
rlabel metal2 18096 22512 18096 22512 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit15.Q
rlabel via1 18528 38170 18528 38170 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit16.Q
rlabel metal2 20352 36876 20352 36876 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit17.Q
rlabel metal2 18048 43554 18048 43554 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit18.Q
rlabel metal2 19632 42168 19632 42168 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit19.Q
rlabel metal2 17664 45192 17664 45192 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit2.Q
rlabel metal2 9600 26082 9600 26082 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit20.Q
rlabel metal2 11640 26040 11640 26040 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit21.Q
rlabel metal2 18192 19992 18192 19992 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit22.Q
rlabel metal2 19944 19992 19944 19992 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit23.Q
rlabel metal2 13824 35154 13824 35154 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit24.Q
rlabel metal2 15176 35112 15176 35112 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit25.Q
rlabel metal3 13440 44730 13440 44730 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit26.Q
rlabel metal3 15072 44730 15072 44730 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit27.Q
rlabel metal2 6336 42714 6336 42714 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit28.Q
rlabel metal2 7944 42672 7944 42672 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit29.Q
rlabel metal2 19352 45696 19352 45696 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit3.Q
rlabel metal2 8688 44016 8688 44016 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit30.Q
rlabel metal2 10368 43806 10368 43806 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit31.Q
rlabel metal2 7584 26124 7584 26124 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit4.Q
rlabel metal2 9168 25998 9168 25998 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit5.Q
rlabel metal2 18432 19362 18432 19362 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit6.Q
rlabel metal3 19968 19026 19968 19026 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit7.Q
rlabel metal3 18528 31794 18528 31794 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit8.Q
rlabel metal2 20256 31626 20256 31626 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit9.Q
rlabel metal2 18240 40488 18240 40488 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame3_bit0.Q
rlabel metal3 20160 40194 20160 40194 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame3_bit1.Q
rlabel metal3 14688 38976 14688 38976 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame3_bit10.Q
rlabel metal2 15888 39144 15888 39144 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame3_bit11.Q
rlabel metal2 7008 30534 7008 30534 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame3_bit12.Q
rlabel metal2 8760 30576 8760 30576 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame3_bit13.Q
rlabel metal2 14913 26040 14913 26040 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame3_bit14.Q
rlabel via2 16808 26040 16808 26040 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame3_bit15.Q
rlabel metal2 18384 37464 18384 37464 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame3_bit16.Q
rlabel metal2 20016 37464 20016 37464 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame3_bit17.Q
rlabel metal2 17904 42672 17904 42672 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame3_bit18.Q
rlabel metal2 19496 42672 19496 42672 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame3_bit19.Q
rlabel metal3 17664 44730 17664 44730 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame3_bit2.Q
rlabel metal3 9312 24696 9312 24696 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame3_bit20.Q
rlabel metal2 11136 25368 11136 25368 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame3_bit21.Q
rlabel metal3 18528 14784 18528 14784 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame3_bit22.Q
rlabel metal2 20448 14196 20448 14196 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame3_bit23.Q
rlabel metal2 14112 34440 14112 34440 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame3_bit24.Q
rlabel metal2 15744 33852 15744 33852 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame3_bit25.Q
rlabel metal3 13440 46200 13440 46200 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame3_bit26.Q
rlabel metal3 14976 47166 14976 47166 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame3_bit27.Q
rlabel metal3 7488 27678 7488 27678 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame3_bit28.Q
rlabel metal2 7968 27804 7968 27804 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame3_bit29.Q
rlabel metal2 19872 45024 19872 45024 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame3_bit3.Q
rlabel metal2 16224 25410 16224 25410 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame3_bit30.Q
rlabel metal3 17760 25620 17760 25620 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame3_bit31.Q
rlabel metal3 7296 26376 7296 26376 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame3_bit4.Q
rlabel metal2 9456 25536 9456 25536 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame3_bit5.Q
rlabel metal3 18144 16002 18144 16002 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame3_bit6.Q
rlabel metal2 20256 16296 20256 16296 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame3_bit7.Q
rlabel metal2 18480 33012 18480 33012 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame3_bit8.Q
rlabel metal2 20064 33432 20064 33432 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame3_bit9.Q
rlabel metal2 9696 29946 9696 29946 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame4_bit0.Q
rlabel metal2 11136 27804 11136 27804 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame4_bit1.Q
rlabel via1 6931 12432 6931 12432 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame4_bit10.Q
rlabel metal2 5472 12516 5472 12516 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame4_bit11.Q
rlabel metal2 12144 19488 12144 19488 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame4_bit12.Q
rlabel metal2 10512 19992 10512 19992 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame4_bit13.Q
rlabel metal3 16704 17514 16704 17514 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame4_bit14.Q
rlabel metal2 15072 17808 15072 17808 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame4_bit15.Q
rlabel metal2 4472 24528 4472 24528 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame4_bit16.Q
rlabel metal3 2784 25200 2784 25200 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame4_bit17.Q
rlabel metal2 6048 22302 6048 22302 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame4_bit18.Q
rlabel metal2 7776 21756 7776 21756 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame4_bit19.Q
rlabel metal2 6024 9408 6024 9408 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame4_bit2.Q
rlabel metal3 16704 29400 16704 29400 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame4_bit20.Q
rlabel metal2 16320 27804 16320 27804 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame4_bit21.Q
rlabel metal2 19200 28560 19200 28560 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame4_bit22.Q
rlabel metal2 19872 28014 19872 28014 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame4_bit23.Q
rlabel metal2 6720 37212 6720 37212 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame4_bit24.Q
rlabel metal2 7989 36624 7989 36624 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame4_bit25.Q
rlabel via1 3270 33600 3270 33600 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame4_bit26.Q
rlabel metal2 3072 33558 3072 33558 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame4_bit27.Q
rlabel metal2 6576 29904 6576 29904 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame4_bit28.Q
rlabel metal3 8256 30534 8256 30534 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame4_bit29.Q
rlabel metal3 4512 8736 4512 8736 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame4_bit3.Q
rlabel metal2 16944 24528 16944 24528 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame4_bit30.Q
rlabel metal2 18624 24633 18624 24633 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame4_bit31.Q
rlabel metal2 12248 4872 12248 4872 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame4_bit4.Q
rlabel metal2 10656 4872 10656 4872 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame4_bit5.Q
rlabel metal2 17520 17808 17520 17808 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame4_bit6.Q
rlabel metal2 19200 17808 19200 17808 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame4_bit7.Q
rlabel metal2 5520 19320 5520 19320 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame4_bit8.Q
rlabel metal3 7200 18816 7200 18816 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame4_bit9.Q
rlabel metal2 3648 22386 3648 22386 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame5_bit0.Q
rlabel metal2 5280 22344 5280 22344 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame5_bit1.Q
rlabel metal2 4032 6636 4032 6636 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame5_bit10.Q
rlabel metal3 5856 8442 5856 8442 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame5_bit11.Q
rlabel metal3 13056 6006 13056 6006 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame5_bit12.Q
rlabel metal2 14448 5712 14448 5712 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame5_bit13.Q
rlabel via1 17864 14804 17864 14804 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame5_bit14.Q
rlabel metal3 17376 14028 17376 14028 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame5_bit15.Q
rlabel metal2 2688 19572 2688 19572 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame5_bit16.Q
rlabel metal2 4608 19362 4608 19362 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame5_bit17.Q
rlabel metal2 5040 13944 5040 13944 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame5_bit18.Q
rlabel via2 7112 13944 7112 13944 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame5_bit19.Q
rlabel metal3 2832 8148 2832 8148 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame5_bit2.Q
rlabel metal2 9168 9408 9168 9408 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame5_bit20.Q
rlabel metal2 10664 9408 10664 9408 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame5_bit21.Q
rlabel metal2 18240 13356 18240 13356 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame5_bit22.Q
rlabel metal2 19824 11592 19824 11592 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame5_bit23.Q
rlabel metal2 3072 23898 3072 23898 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame5_bit24.Q
rlabel metal3 3744 24318 3744 24318 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame5_bit25.Q
rlabel metal2 8976 16464 8976 16464 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame5_bit26.Q
rlabel metal3 10752 16338 10752 16338 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame5_bit27.Q
rlabel metal2 15216 13860 15216 13860 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame5_bit28.Q
rlabel metal2 16824 13944 16824 13944 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame5_bit29.Q
rlabel metal2 4032 7392 4032 7392 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame5_bit3.Q
rlabel metal2 13296 11760 13296 11760 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame5_bit30.Q
rlabel metal3 14976 11466 14976 11466 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame5_bit31.Q
rlabel metal2 10656 5124 10656 5124 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame5_bit4.Q
rlabel metal2 12432 3948 12432 3948 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame5_bit5.Q
rlabel metal2 15744 10416 15744 10416 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame5_bit6.Q
rlabel metal2 16952 10920 16952 10920 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame5_bit7.Q
rlabel metal2 3168 13440 3168 13440 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame5_bit8.Q
rlabel metal3 4704 16758 4704 16758 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame5_bit9.Q
rlabel metal2 2592 21000 2592 21000 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame6_bit0.Q
rlabel metal2 3848 21504 3848 21504 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame6_bit1.Q
rlabel metal3 6720 8022 6720 8022 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame6_bit10.Q
rlabel metal3 7872 8442 7872 8442 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame6_bit11.Q
rlabel metal2 9984 5334 9984 5334 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame6_bit12.Q
rlabel metal2 15624 4872 15624 4872 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame6_bit13.Q
rlabel metal2 8448 14826 8448 14826 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame6_bit14.Q
rlabel metal2 9936 14784 9936 14784 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame6_bit15.Q
rlabel metal2 2544 17136 2544 17136 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame6_bit16.Q
rlabel via2 4040 18480 4040 18480 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame6_bit17.Q
rlabel metal2 2640 13860 2640 13860 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame6_bit18.Q
rlabel via2 4136 13944 4136 13944 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame6_bit19.Q
rlabel metal2 2640 8904 2640 8904 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame6_bit2.Q
rlabel metal2 8736 7140 8736 7140 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame6_bit20.Q
rlabel metal2 10176 7224 10176 7224 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame6_bit21.Q
rlabel metal2 19248 8904 19248 8904 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame6_bit22.Q
rlabel metal2 19248 8148 19248 8148 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame6_bit23.Q
rlabel metal3 2784 16338 2784 16338 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame6_bit24.Q
rlabel via1 4616 16968 4616 16968 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame6_bit25.Q
rlabel metal2 7296 13146 7296 13146 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame6_bit26.Q
rlabel via2 9128 13944 9128 13944 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame6_bit27.Q
rlabel metal3 16128 7896 16128 7896 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame6_bit28.Q
rlabel metal3 17376 7938 17376 7938 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame6_bit29.Q
rlabel metal2 3848 12432 3848 12432 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame6_bit3.Q
rlabel metal2 17760 10416 17760 10416 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame6_bit30.Q
rlabel metal2 19448 12432 19448 12432 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame6_bit31.Q
rlabel metal3 8064 5754 8064 5754 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame6_bit4.Q
rlabel via2 9992 6384 9992 6384 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame6_bit5.Q
rlabel metal3 17760 8778 17760 8778 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame6_bit6.Q
rlabel metal3 19776 8022 19776 8022 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame6_bit7.Q
rlabel metal2 3120 14952 3120 14952 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame6_bit8.Q
rlabel metal2 4896 15624 4896 15624 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame6_bit9.Q
rlabel metal2 18336 26880 18336 26880 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit0.Q
rlabel metal2 20112 26880 20112 26880 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit1.Q
rlabel metal2 20256 20874 20256 20874 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit10.Q
rlabel metal2 19198 23814 19198 23814 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit11.Q
rlabel metal2 13920 31458 13920 31458 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit12.Q
rlabel metal2 13449 30618 13449 30618 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit13.Q
rlabel metal2 14880 29862 14880 29862 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit14.Q
rlabel metal2 12240 38136 12240 38136 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit15.Q
rlabel metal2 12096 38430 12096 38430 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit16.Q
rlabel metal2 13865 40488 13865 40488 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit17.Q
rlabel via2 9128 18480 9128 18480 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit18.Q
rlabel metal2 6912 17220 6912 17220 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit19.Q
rlabel metal3 17472 29190 17472 29190 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit2.Q
rlabel metal2 13976 18480 13976 18480 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit20.Q
rlabel metal2 12336 18480 12336 18480 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit21.Q
rlabel metal2 13016 10920 13016 10920 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit22.Q
rlabel metal2 11520 10878 11520 10878 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit23.Q
rlabel metal2 10992 20832 10992 20832 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit24.Q
rlabel metal2 9408 20874 9408 20874 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit25.Q
rlabel metal2 6000 10920 6000 10920 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit26.Q
rlabel metal2 8016 10416 8016 10416 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit27.Q
rlabel metal2 15393 6384 15393 6384 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit28.Q
rlabel via2 17000 6384 17000 6384 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit29.Q
rlabel metal2 18720 29820 18720 29820 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit3.Q
rlabel metal2 8304 11172 8304 11172 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit30.Q
rlabel metal2 10272 11802 10272 11802 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit31.Q
rlabel metal2 7928 24528 7928 24528 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit4.Q
rlabel metal2 6432 24570 6432 24570 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit5.Q
rlabel metal2 2688 27678 2688 27678 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit6.Q
rlabel metal3 2688 28434 2688 28434 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit7.Q
rlabel metal2 4320 27048 4320 27048 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit8.Q
rlabel metal2 19632 21504 19632 21504 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit9.Q
rlabel metal4 5664 38388 5664 38388 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit0.Q
rlabel metal2 8640 39018 8640 39018 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit1.Q
rlabel metal2 17938 36498 17938 36498 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit10.Q
rlabel metal2 15333 42672 15333 42672 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit11.Q
rlabel metal2 14880 41706 14880 41706 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit12.Q
rlabel metal2 15120 42000 15120 42000 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit13.Q
rlabel metal2 4992 32340 4992 32340 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit14.Q
rlabel metal2 6624 32340 6624 32340 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit15.Q
rlabel metal2 13728 23016 13728 23016 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit16.Q
rlabel via2 15368 23016 15368 23016 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit17.Q
rlabel metal2 15456 36624 15456 36624 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit18.Q
rlabel metal2 17424 35784 17424 35784 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit19.Q
rlabel metal2 3696 29064 3696 29064 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit2.Q
rlabel metal2 11040 45948 11040 45948 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit20.Q
rlabel metal2 12384 46536 12384 46536 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit21.Q
rlabel metal3 2688 38430 2688 38430 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit22.Q
rlabel metal2 4088 39648 4088 39648 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit23.Q
rlabel metal2 13728 32970 13728 32970 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit24.Q
rlabel metal2 14640 33432 14640 33432 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit25.Q
rlabel metal2 13056 42378 13056 42378 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit26.Q
rlabel metal2 11328 42000 11328 42000 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit27.Q
rlabel metal2 3704 36624 3704 36624 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit28.Q
rlabel metal2 2640 33852 2640 33852 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit29.Q
rlabel metal3 2784 29106 2784 29106 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit3.Q
rlabel metal2 4560 33096 4560 33096 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit30.Q
rlabel metal3 2784 32352 2784 32352 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit31.Q
rlabel metal2 3648 30072 3648 30072 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit4.Q
rlabel metal2 13584 20916 13584 20916 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit5.Q
rlabel metal2 13968 21336 13968 21336 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit6.Q
rlabel metal2 15456 21000 15456 21000 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit7.Q
rlabel metal2 17568 36582 17568 36582 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit8.Q
rlabel metal2 16416 35070 16416 35070 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit9.Q
rlabel metal2 8976 36624 8976 36624 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame9_bit10.Q
rlabel metal2 10431 36624 10431 36624 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame9_bit11.Q
rlabel metal2 15360 23856 15360 23856 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame9_bit12.Q
rlabel metal2 14016 23898 14016 23898 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame9_bit13.Q
rlabel metal2 11952 36120 11952 36120 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame9_bit14.Q
rlabel via1 14314 36643 14314 36643 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame9_bit15.Q
rlabel metal2 9512 47208 9512 47208 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame9_bit16.Q
rlabel metal2 7920 47208 7920 47208 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame9_bit17.Q
rlabel metal2 2640 38388 2640 38388 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame9_bit18.Q
rlabel metal2 4138 40488 4138 40488 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame9_bit19.Q
rlabel metal3 13536 30702 13536 30702 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame9_bit20.Q
rlabel via2 15272 32088 15272 32088 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame9_bit21.Q
rlabel via2 12392 41160 12392 41160 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame9_bit22.Q
rlabel metal2 10737 41160 10737 41160 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame9_bit23.Q
rlabel metal2 3648 35952 3648 35952 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame9_bit24.Q
rlabel metal2 2256 35952 2256 35952 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame9_bit25.Q
rlabel metal2 2544 44100 2544 44100 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame9_bit26.Q
rlabel metal2 3216 42084 3216 42084 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame9_bit27.Q
rlabel metal2 19496 41160 19496 41160 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame9_bit28.Q
rlabel metal3 17760 40530 17760 40530 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame9_bit29.Q
rlabel metal2 17912 30576 17912 30576 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame9_bit30.Q
rlabel metal2 16368 30576 16368 30576 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame9_bit31.Q
rlabel metal3 14928 15540 14928 15540 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.J_NS4_BEG10
rlabel metal2 13104 39564 13104 39564 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.J_NS4_BEG11
rlabel metal2 4320 22260 4320 22260 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.J_NS4_BEG12
rlabel metal2 18576 22260 18576 22260 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.J_NS4_BEG13
rlabel metal2 16320 13944 16320 13944 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.J_NS4_BEG14
rlabel metal2 15504 42756 15504 42756 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.J_NS4_BEG15
rlabel metal2 9024 21000 9024 21000 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.J_NS4_BEG4
rlabel metal3 19008 21042 19008 21042 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.J_NS4_BEG5
rlabel metal2 13632 19908 13632 19908 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.J_NS4_BEG6
rlabel metal4 14448 42252 14448 42252 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.J_NS4_BEG7
rlabel metal3 10176 17934 10176 17934 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.J_NS4_BEG8
rlabel metal2 14640 14952 14640 14952 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.J_NS4_BEG9
rlabel metal2 7080 32676 7080 32676 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.S1BEG0
rlabel metal2 15672 23268 15672 23268 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.S1BEG1
rlabel metal2 18096 35196 18096 35196 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.S1BEG2
rlabel metal2 12600 46452 12600 46452 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.S1BEG3
rlabel metal2 2112 43512 2112 43512 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.S2BEG0
rlabel metal2 17328 32844 17328 32844 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.S2BEG1
rlabel metal2 13344 42168 13344 42168 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.S2BEG2
rlabel metal2 5520 36372 5520 36372 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.S2BEG3
rlabel metal2 4728 34356 4728 34356 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.S2BEG4
rlabel metal2 19488 27048 19488 27048 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.S2BEG5
rlabel metal2 18816 30072 18816 30072 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.S2BEG6
rlabel metal2 8280 24612 8280 24612 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.S2BEG7
rlabel metal3 4464 18564 4464 18564 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.S4BEG0
rlabel metal3 19680 19908 19680 19908 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.S4BEG1
rlabel metal2 14592 29148 14592 29148 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.S4BEG2
rlabel metal2 13056 40488 13056 40488 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.S4BEG3
rlabel metal2 9528 18564 9528 18564 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.W1BEG0
rlabel metal2 14304 17724 14304 17724 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.W1BEG1
rlabel metal2 14496 9492 14496 9492 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.W1BEG2
rlabel metal2 11352 20748 11352 20748 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.W1BEG3
rlabel metal2 8112 10164 8112 10164 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.W2BEG0
rlabel metal2 17400 6468 17400 6468 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.W2BEG1
rlabel metal2 10680 11676 10680 11676 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.W2BEG2
rlabel metal4 4272 20748 4272 20748 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.W2BEG3
rlabel metal2 4896 11760 4896 11760 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.W2BEG4
rlabel metal2 10272 5628 10272 5628 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.W2BEG5
rlabel metal3 19680 8190 19680 8190 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.W2BEG6
rlabel metal2 5808 16464 5808 16464 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.W2BEG7
rlabel metal2 8280 8652 8280 8652 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.W2BEGb0
rlabel metal2 15960 4956 15960 4956 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.W2BEGb1
rlabel metal2 10200 14616 10200 14616 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.W2BEGb2
rlabel metal2 4296 18564 4296 18564 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.W2BEGb3
rlabel metal2 4416 13776 4416 13776 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.W2BEGb4
rlabel metal2 10632 7056 10632 7056 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.W2BEGb5
rlabel metal2 17664 9534 17664 9534 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.W2BEGb6
rlabel metal2 6144 16212 6144 16212 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.W2BEGb7
rlabel metal2 10968 17052 10968 17052 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.W6BEG0
rlabel metal2 17760 13272 17760 13272 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.W6BEG1
rlabel metal2 17112 17724 17112 17724 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.W6BEG10
rlabel metal3 4320 23730 4320 23730 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.W6BEG11
rlabel metal2 15384 11676 15384 11676 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.W6BEG2
rlabel metal2 11640 29820 11640 29820 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.W6BEG3
rlabel metal2 6168 9492 6168 9492 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.W6BEG4
rlabel metal2 12792 4956 12792 4956 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.W6BEG5
rlabel metal2 15072 17724 15072 17724 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.W6BEG6
rlabel metal2 8160 19320 8160 19320 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.W6BEG7
rlabel metal2 7320 12516 7320 12516 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.W6BEG8
rlabel metal2 12600 20076 12600 20076 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.W6BEG9
rlabel metal2 9528 14028 9528 14028 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.WW4BEG0
rlabel metal2 17856 8904 17856 8904 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.WW4BEG1
rlabel metal2 16032 14700 16032 14700 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.WW4BEG10
rlabel metal2 5040 19488 5040 19488 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.WW4BEG11
rlabel metal2 7920 13188 7920 13188 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.WW4BEG12
rlabel metal2 11256 9492 11256 9492 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.WW4BEG13
rlabel metal2 19248 12684 19248 12684 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.WW4BEG14
rlabel metal3 7200 24654 7200 24654 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.WW4BEG15
rlabel metal2 16704 11760 16704 11760 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.WW4BEG2
rlabel metal2 5424 22512 5424 22512 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.WW4BEG3
rlabel metal3 4608 9534 4608 9534 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.WW4BEG4
rlabel metal3 13344 5208 13344 5208 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.WW4BEG5
rlabel metal2 17400 11004 17400 11004 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.WW4BEG6
rlabel metal2 5520 17976 5520 17976 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.WW4BEG7
rlabel metal2 6912 9324 6912 9324 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.WW4BEG8
rlabel metal3 15072 6174 15072 6174 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.WW4BEG9
rlabel metal3 1824 912 1824 912 0 Tile_X0Y1_N1END[0]
rlabel metal2 2400 4032 2400 4032 0 Tile_X0Y1_N1END[1]
rlabel metal3 2208 1836 2208 1836 0 Tile_X0Y1_N1END[2]
rlabel metal3 2400 1038 2400 1038 0 Tile_X0Y1_N1END[3]
rlabel metal3 4128 534 4128 534 0 Tile_X0Y1_N2END[0]
rlabel metal3 4320 1332 4320 1332 0 Tile_X0Y1_N2END[1]
rlabel metal3 4512 954 4512 954 0 Tile_X0Y1_N2END[2]
rlabel metal3 4704 1332 4704 1332 0 Tile_X0Y1_N2END[3]
rlabel metal3 4896 450 4896 450 0 Tile_X0Y1_N2END[4]
rlabel metal3 5088 702 5088 702 0 Tile_X0Y1_N2END[5]
rlabel metal3 5280 534 5280 534 0 Tile_X0Y1_N2END[6]
rlabel metal3 5472 1290 5472 1290 0 Tile_X0Y1_N2END[7]
rlabel metal3 2592 912 2592 912 0 Tile_X0Y1_N2MID[0]
rlabel metal3 2784 954 2784 954 0 Tile_X0Y1_N2MID[1]
rlabel metal3 2976 954 2976 954 0 Tile_X0Y1_N2MID[2]
rlabel metal3 3168 1332 3168 1332 0 Tile_X0Y1_N2MID[3]
rlabel metal3 3360 954 3360 954 0 Tile_X0Y1_N2MID[4]
rlabel metal3 3552 1248 3552 1248 0 Tile_X0Y1_N2MID[5]
rlabel metal3 3744 1038 3744 1038 0 Tile_X0Y1_N2MID[6]
rlabel metal3 3936 702 3936 702 0 Tile_X0Y1_N2MID[7]
rlabel metal3 5664 1038 5664 1038 0 Tile_X0Y1_N4END[0]
rlabel metal3 7584 198 7584 198 0 Tile_X0Y1_N4END[10]
rlabel metal3 7776 744 7776 744 0 Tile_X0Y1_N4END[11]
rlabel metal2 6336 5544 6336 5544 0 Tile_X0Y1_N4END[12]
rlabel metal3 8160 744 8160 744 0 Tile_X0Y1_N4END[13]
rlabel metal3 8352 744 8352 744 0 Tile_X0Y1_N4END[14]
rlabel metal3 8544 744 8544 744 0 Tile_X0Y1_N4END[15]
rlabel metal3 5856 1332 5856 1332 0 Tile_X0Y1_N4END[1]
rlabel metal3 6048 954 6048 954 0 Tile_X0Y1_N4END[2]
rlabel metal3 6240 954 6240 954 0 Tile_X0Y1_N4END[3]
rlabel metal3 6432 996 6432 996 0 Tile_X0Y1_N4END[4]
rlabel metal3 6624 996 6624 996 0 Tile_X0Y1_N4END[5]
rlabel metal3 6816 954 6816 954 0 Tile_X0Y1_N4END[6]
rlabel metal3 7008 996 7008 996 0 Tile_X0Y1_N4END[7]
rlabel metal3 2784 93240 2784 93240 0 Tile_X0Y1_N4END[8]
rlabel metal2 3264 5502 3264 5502 0 Tile_X0Y1_N4END[9]
rlabel metal3 8736 870 8736 870 0 Tile_X0Y1_S1BEG[0]
rlabel metal3 8928 1248 8928 1248 0 Tile_X0Y1_S1BEG[1]
rlabel metal3 9120 870 9120 870 0 Tile_X0Y1_S1BEG[2]
rlabel metal3 9312 1248 9312 1248 0 Tile_X0Y1_S1BEG[3]
rlabel metal3 9504 870 9504 870 0 Tile_X0Y1_S2BEG[0]
rlabel metal3 9696 1248 9696 1248 0 Tile_X0Y1_S2BEG[1]
rlabel metal3 9888 870 9888 870 0 Tile_X0Y1_S2BEG[2]
rlabel metal3 10080 1248 10080 1248 0 Tile_X0Y1_S2BEG[3]
rlabel metal3 10272 870 10272 870 0 Tile_X0Y1_S2BEG[4]
rlabel metal3 10464 1248 10464 1248 0 Tile_X0Y1_S2BEG[5]
rlabel metal3 10656 870 10656 870 0 Tile_X0Y1_S2BEG[6]
rlabel metal3 10848 1248 10848 1248 0 Tile_X0Y1_S2BEG[7]
rlabel metal3 11040 870 11040 870 0 Tile_X0Y1_S2BEGb[0]
rlabel metal3 11232 912 11232 912 0 Tile_X0Y1_S2BEGb[1]
rlabel metal3 11424 870 11424 870 0 Tile_X0Y1_S2BEGb[2]
rlabel metal3 11616 870 11616 870 0 Tile_X0Y1_S2BEGb[3]
rlabel metal3 11808 912 11808 912 0 Tile_X0Y1_S2BEGb[4]
rlabel metal3 12000 870 12000 870 0 Tile_X0Y1_S2BEGb[5]
rlabel metal3 12192 870 12192 870 0 Tile_X0Y1_S2BEGb[6]
rlabel metal2 13080 1680 13080 1680 0 Tile_X0Y1_S2BEGb[7]
rlabel metal3 12576 1248 12576 1248 0 Tile_X0Y1_S4BEG[0]
rlabel metal3 14496 1248 14496 1248 0 Tile_X0Y1_S4BEG[10]
rlabel metal3 14688 912 14688 912 0 Tile_X0Y1_S4BEG[11]
rlabel metal3 14880 1248 14880 1248 0 Tile_X0Y1_S4BEG[12]
rlabel metal3 15072 828 15072 828 0 Tile_X0Y1_S4BEG[13]
rlabel metal3 15264 1248 15264 1248 0 Tile_X0Y1_S4BEG[14]
rlabel metal3 15456 828 15456 828 0 Tile_X0Y1_S4BEG[15]
rlabel metal3 12768 912 12768 912 0 Tile_X0Y1_S4BEG[1]
rlabel metal2 12984 2436 12984 2436 0 Tile_X0Y1_S4BEG[2]
rlabel metal3 13152 828 13152 828 0 Tile_X0Y1_S4BEG[3]
rlabel metal3 13344 1248 13344 1248 0 Tile_X0Y1_S4BEG[4]
rlabel metal3 13536 828 13536 828 0 Tile_X0Y1_S4BEG[5]
rlabel metal3 13728 1248 13728 1248 0 Tile_X0Y1_S4BEG[6]
rlabel metal3 13920 1038 13920 1038 0 Tile_X0Y1_S4BEG[7]
rlabel metal3 14112 1248 14112 1248 0 Tile_X0Y1_S4BEG[8]
rlabel metal3 14304 828 14304 828 0 Tile_X0Y1_S4BEG[9]
rlabel metal3 15648 324 15648 324 0 Tile_X0Y1_UserCLK
rlabel metal2 944 2772 944 2772 0 Tile_X0Y1_W1BEG[0]
rlabel metal2 840 2856 840 2856 0 Tile_X0Y1_W1BEG[1]
rlabel metal2 128 3444 128 3444 0 Tile_X0Y1_W1BEG[2]
rlabel metal2 1088 3780 1088 3780 0 Tile_X0Y1_W1BEG[3]
rlabel metal2 416 4116 416 4116 0 Tile_X0Y1_W2BEG[0]
rlabel metal2 224 4452 224 4452 0 Tile_X0Y1_W2BEG[1]
rlabel metal2 1400 4788 1400 4788 0 Tile_X0Y1_W2BEG[2]
rlabel metal2 512 5124 512 5124 0 Tile_X0Y1_W2BEG[3]
rlabel metal2 560 5460 560 5460 0 Tile_X0Y1_W2BEG[4]
rlabel metal2 176 5796 176 5796 0 Tile_X0Y1_W2BEG[5]
rlabel metal2 704 6132 704 6132 0 Tile_X0Y1_W2BEG[6]
rlabel metal2 320 6468 320 6468 0 Tile_X0Y1_W2BEG[7]
rlabel metal2 1472 6804 1472 6804 0 Tile_X0Y1_W2BEGb[0]
rlabel metal2 368 7140 368 7140 0 Tile_X0Y1_W2BEGb[1]
rlabel metal2 560 7476 560 7476 0 Tile_X0Y1_W2BEGb[2]
rlabel metal2 848 7812 848 7812 0 Tile_X0Y1_W2BEGb[3]
rlabel metal2 224 8148 224 8148 0 Tile_X0Y1_W2BEGb[4]
rlabel metal2 464 8484 464 8484 0 Tile_X0Y1_W2BEGb[5]
rlabel metal2 608 8820 608 8820 0 Tile_X0Y1_W2BEGb[6]
rlabel metal2 3768 6972 3768 6972 0 Tile_X0Y1_W2BEGb[7]
rlabel metal2 800 14868 800 14868 0 Tile_X0Y1_W6BEG[0]
rlabel metal2 320 18228 320 18228 0 Tile_X0Y1_W6BEG[10]
rlabel metal2 608 18564 608 18564 0 Tile_X0Y1_W6BEG[11]
rlabel metal2 224 15204 224 15204 0 Tile_X0Y1_W6BEG[1]
rlabel metal2 128 15540 128 15540 0 Tile_X0Y1_W6BEG[2]
rlabel metal2 704 15876 704 15876 0 Tile_X0Y1_W6BEG[3]
rlabel metal2 176 16212 176 16212 0 Tile_X0Y1_W6BEG[4]
rlabel metal2 800 16548 800 16548 0 Tile_X0Y1_W6BEG[5]
rlabel metal2 752 16884 752 16884 0 Tile_X0Y1_W6BEG[6]
rlabel metal2 4728 13860 4728 13860 0 Tile_X0Y1_W6BEG[7]
rlabel metal2 704 17556 704 17556 0 Tile_X0Y1_W6BEG[8]
rlabel metal2 944 17892 944 17892 0 Tile_X0Y1_W6BEG[9]
rlabel metal2 560 9492 560 9492 0 Tile_X0Y1_WW4BEG[0]
rlabel via2 80 12852 80 12852 0 Tile_X0Y1_WW4BEG[10]
rlabel metal2 608 13188 608 13188 0 Tile_X0Y1_WW4BEG[11]
rlabel metal2 944 13524 944 13524 0 Tile_X0Y1_WW4BEG[12]
rlabel via2 80 13860 80 13860 0 Tile_X0Y1_WW4BEG[13]
rlabel metal2 7200 14364 7200 14364 0 Tile_X0Y1_WW4BEG[14]
rlabel metal2 1328 14532 1328 14532 0 Tile_X0Y1_WW4BEG[15]
rlabel metal2 656 9828 656 9828 0 Tile_X0Y1_WW4BEG[1]
rlabel metal2 128 10164 128 10164 0 Tile_X0Y1_WW4BEG[2]
rlabel metal2 368 10500 368 10500 0 Tile_X0Y1_WW4BEG[3]
rlabel metal2 848 10836 848 10836 0 Tile_X0Y1_WW4BEG[4]
rlabel metal2 272 11172 272 11172 0 Tile_X0Y1_WW4BEG[5]
rlabel metal2 1040 11508 1040 11508 0 Tile_X0Y1_WW4BEG[6]
rlabel metal2 512 11844 512 11844 0 Tile_X0Y1_WW4BEG[7]
rlabel metal2 416 12180 416 12180 0 Tile_X0Y1_WW4BEG[8]
rlabel metal2 368 12516 368 12516 0 Tile_X0Y1_WW4BEG[9]
rlabel metal2 12480 60606 12480 60606 0 WEN_SRAM
rlabel metal2 4536 42504 4536 42504 0 _0000_
rlabel metal2 6672 40908 6672 40908 0 _0001_
rlabel metal3 7200 46200 7200 46200 0 _0002_
rlabel metal2 19944 73584 19944 73584 0 _0003_
rlabel metal2 12648 78456 12648 78456 0 _0004_
rlabel metal2 5496 79128 5496 79128 0 _0005_
rlabel via1 10760 58632 10760 58632 0 _0006_
rlabel via1 11230 45024 11230 45024 0 _0007_
rlabel via1 12670 35952 12670 35952 0 _0008_
rlabel metal2 14592 22302 14592 22302 0 _0009_
rlabel via1 7656 35112 7656 35112 0 _0010_
rlabel metal2 8640 63714 8640 63714 0 _0011_
rlabel metal2 19992 76944 19992 76944 0 _0012_
rlabel metal3 14400 85050 14400 85050 0 _0013_
rlabel metal3 7872 81606 7872 81606 0 _0014_
rlabel metal4 10560 53340 10560 53340 0 _0015_
rlabel metal3 17568 59304 17568 59304 0 _0016_
rlabel metal2 15672 82068 15672 82068 0 _0017_
rlabel metal2 6408 83748 6408 83748 0 _0018_
rlabel metal2 4728 32676 4728 32676 0 _0019_
rlabel metal2 4704 30366 4704 30366 0 _0020_
rlabel metal2 13917 19992 13917 19992 0 _0021_
rlabel metal2 15888 19404 15888 19404 0 _0022_
rlabel metal2 16032 35196 16032 35196 0 _0023_
rlabel metal2 18456 34944 18456 34944 0 _0024_
rlabel metal2 15888 42924 15888 42924 0 _0025_
rlabel metal2 16248 41412 16248 41412 0 _0026_
rlabel metal2 3384 25956 3384 25956 0 _0027_
rlabel metal2 4008 27384 4008 27384 0 _0028_
rlabel metal2 18528 18564 18528 18564 0 _0029_
rlabel metal2 20712 20160 20712 20160 0 _0030_
rlabel metal2 14196 29904 14196 29904 0 _0031_
rlabel metal2 15360 31500 15360 31500 0 _0032_
rlabel metal2 12960 38934 12960 38934 0 _0033_
rlabel metal3 13632 39018 13632 39018 0 _0034_
rlabel metal2 6432 44940 6432 44940 0 _0035_
rlabel via2 5658 45108 5658 45108 0 _0036_
rlabel metal2 7413 40488 7413 40488 0 _0037_
rlabel metal2 6984 74676 6984 74676 0 _0038_
rlabel metal2 17784 74676 17784 74676 0 _0039_
rlabel metal3 13248 86268 13248 86268 0 _0040_
rlabel via2 4243 54096 4243 54096 0 _0041_
rlabel metal2 6792 67536 6792 67536 0 _0042_
rlabel metal2 6000 39144 6000 39144 0 _0043_
rlabel metal2 7344 45654 7344 45654 0 _0044_
rlabel metal2 7248 44436 7248 44436 0 _0045_
rlabel metal2 7104 44856 7104 44856 0 _0046_
rlabel metal2 8208 45024 8208 45024 0 _0047_
rlabel metal2 6720 45696 6720 45696 0 _0048_
rlabel metal2 8855 45066 8855 45066 0 _0049_
rlabel metal2 8736 44898 8736 44898 0 _0050_
rlabel metal2 8520 44940 8520 44940 0 _0051_
rlabel metal3 9216 44688 9216 44688 0 _0052_
rlabel metal2 8496 42756 8496 42756 0 _0053_
rlabel metal2 8532 42672 8532 42672 0 _0054_
rlabel metal2 9408 42924 9408 42924 0 _0055_
rlabel metal2 9518 44058 9518 44058 0 _0056_
rlabel metal2 19392 72791 19392 72791 0 _0057_
rlabel metal2 19200 72912 19200 72912 0 _0058_
rlabel metal2 15456 74382 15456 74382 0 _0059_
rlabel metal2 13248 18480 13248 18480 0 _0060_
rlabel metal2 14304 22302 14304 22302 0 _0061_
rlabel metal2 14208 22386 14208 22386 0 _0062_
rlabel metal2 14784 23016 14784 23016 0 _0063_
rlabel metal2 12696 79884 12696 79884 0 _0064_
rlabel metal2 12768 79002 12768 79002 0 _0065_
rlabel metal3 13248 77364 13248 77364 0 _0066_
rlabel metal2 13365 35112 13365 35112 0 _0067_
rlabel via1 12287 35952 12287 35952 0 _0068_
rlabel metal2 12384 35994 12384 35994 0 _0069_
rlabel metal2 13440 36624 13440 36624 0 _0070_
rlabel metal2 3264 79758 3264 79758 0 _0071_
rlabel metal2 3216 79212 3216 79212 0 _0072_
rlabel metal2 8399 86520 8399 86520 0 _0073_
rlabel metal2 9984 20706 9984 20706 0 _0074_
rlabel metal3 10848 45654 10848 45654 0 _0075_
rlabel metal3 10368 45906 10368 45906 0 _0076_
rlabel metal2 11616 46536 11616 46536 0 _0077_
rlabel metal2 16080 19236 16080 19236 0 _0078_
rlabel metal2 15696 35112 15696 35112 0 _0079_
rlabel metal2 7104 42168 7104 42168 0 _0080_
rlabel metal2 4224 48216 4224 48216 0 _0081_
rlabel metal2 19056 41160 19056 41160 0 _0082_
rlabel metal4 17952 35112 17952 35112 0 _0083_
rlabel metal2 12768 39018 12768 39018 0 _0084_
rlabel metal2 12192 57624 12192 57624 0 _0085_
rlabel metal2 11520 58086 11520 58086 0 _0086_
rlabel metal2 10752 58842 10752 58842 0 _0087_
rlabel metal2 8784 17724 8784 17724 0 _0088_
rlabel via2 8067 35112 8067 35112 0 _0089_
rlabel metal2 7968 35070 7968 35070 0 _0090_
rlabel metal2 7584 34902 7584 34902 0 _0091_
rlabel metal2 7968 75306 7968 75306 0 _0092_
rlabel metal2 8736 75432 8736 75432 0 _0093_
rlabel metal3 17376 75306 17376 75306 0 _0094_
rlabel metal2 17660 75894 17660 75894 0 _0095_
rlabel metal2 12816 86520 12816 86520 0 _0096_
rlabel via1 13112 86520 13112 86520 0 _0097_
rlabel metal2 3683 54085 3683 54085 0 _0098_
rlabel metal2 4032 54264 4032 54264 0 _0099_
rlabel metal2 7488 69216 7488 69216 0 _0100_
rlabel metal2 7872 69384 7872 69384 0 _0101_
rlabel metal2 8640 63000 8640 63000 0 _0102_
rlabel metal2 8832 63210 8832 63210 0 _0103_
rlabel metal2 9168 63672 9168 63672 0 _0104_
rlabel metal3 9216 63546 9216 63546 0 _0105_
rlabel metal2 9408 63546 9408 63546 0 _0106_
rlabel metal2 9624 62580 9624 62580 0 _0107_
rlabel metal2 9600 63210 9600 63210 0 _0108_
rlabel metal2 20352 77490 20352 77490 0 _0109_
rlabel metal2 19632 78120 19632 78120 0 _0110_
rlabel metal2 20064 78456 20064 78456 0 _0111_
rlabel metal2 20009 77448 20009 77448 0 _0112_
rlabel metal2 19968 77700 19968 77700 0 _0113_
rlabel metal2 14976 78330 14976 78330 0 _0114_
rlabel metal4 18720 80724 18720 80724 0 _0115_
rlabel metal2 14551 84311 14551 84311 0 _0116_
rlabel metal2 13131 84336 13131 84336 0 _0117_
rlabel metal2 13032 84252 13032 84252 0 _0118_
rlabel metal2 13824 84462 13824 84462 0 _0119_
rlabel metal3 14304 85218 14304 85218 0 _0120_
rlabel metal2 14688 84378 14688 84378 0 _0121_
rlabel metal2 14832 84504 14832 84504 0 _0122_
rlabel metal2 7680 81312 7680 81312 0 _0123_
rlabel metal2 6549 80472 6549 80472 0 _0124_
rlabel metal2 6912 80556 6912 80556 0 _0125_
rlabel metal2 7392 80388 7392 80388 0 _0126_
rlabel metal2 8256 81354 8256 81354 0 _0127_
rlabel metal2 7968 82026 7968 82026 0 _0128_
rlabel metal3 8448 81606 8448 81606 0 _0129_
rlabel metal3 10080 52584 10080 52584 0 _0130_
rlabel metal2 10005 52584 10005 52584 0 _0131_
rlabel metal2 9888 51870 9888 51870 0 _0132_
rlabel via2 10373 51744 10373 51744 0 _0133_
rlabel metal2 10368 52038 10368 52038 0 _0134_
rlabel metal2 9984 52752 9984 52752 0 _0135_
rlabel metal2 10608 51996 10608 51996 0 _0136_
rlabel metal2 17664 58674 17664 58674 0 _0137_
rlabel metal2 15819 60144 15819 60144 0 _0138_
rlabel metal2 15840 57960 15840 57960 0 _0139_
rlabel metal2 17321 58716 17321 58716 0 _0140_
rlabel metal3 17376 59262 17376 59262 0 _0141_
rlabel metal2 17808 58632 17808 58632 0 _0142_
rlabel metal2 17904 58800 17904 58800 0 _0143_
rlabel metal2 14928 83496 14928 83496 0 _0144_
rlabel metal2 16728 81270 16728 81270 0 _0145_
rlabel metal2 17088 81228 17088 81228 0 _0146_
rlabel metal2 16464 81480 16464 81480 0 _0147_
rlabel metal2 16512 82908 16512 82908 0 _0148_
rlabel metal2 15792 81816 15792 81816 0 _0149_
rlabel metal2 16320 82866 16320 82866 0 _0150_
rlabel metal2 7632 83748 7632 83748 0 _0151_
rlabel metal2 7728 82236 7728 82236 0 _0152_
rlabel metal2 8736 83580 8736 83580 0 _0153_
rlabel metal2 7776 84252 7776 84252 0 _0154_
rlabel metal3 8544 84546 8544 84546 0 _0155_
rlabel metal3 7872 84756 7872 84756 0 _0156_
rlabel metal2 8400 84336 8400 84336 0 _0157_
rlabel metal3 13680 42168 13680 42168 0 _0158_
rlabel metal2 19632 40488 19632 40488 0 _0159_
rlabel metal2 19008 22260 19008 22260 0 _0160_
rlabel metal4 6000 23772 6000 23772 0 _0161_
rlabel metal2 8928 22260 8928 22260 0 _0162_
rlabel metal2 5280 21798 5280 21798 0 _0163_
rlabel metal2 8784 22260 8784 22260 0 _0164_
rlabel metal3 17088 27888 17088 27888 0 _0165_
rlabel metal2 17801 29064 17801 29064 0 _0166_
rlabel metal2 16992 26712 16992 26712 0 _0167_
rlabel metal2 20256 27594 20256 27594 0 _0168_
rlabel metal2 20016 28560 20016 28560 0 _0169_
rlabel metal2 20160 27510 20160 27510 0 _0170_
rlabel metal2 8352 36708 8352 36708 0 _0171_
rlabel metal2 7200 35784 7200 35784 0 _0172_
rlabel metal3 8256 36960 8256 36960 0 _0173_
rlabel metal2 2928 33348 2928 33348 0 _0174_
rlabel metal3 3360 33852 3360 33852 0 _0175_
rlabel metal2 3408 33348 3408 33348 0 _0176_
rlabel metal2 3648 28602 3648 28602 0 _0177_
rlabel metal3 4608 29022 4608 29022 0 _0178_
rlabel metal2 4512 28224 4512 28224 0 _0179_
rlabel metal2 4800 30618 4800 30618 0 _0180_
rlabel metal3 4512 30912 4512 30912 0 _0181_
rlabel metal2 3408 29169 3408 29169 0 _0182_
rlabel metal2 4872 29568 4872 29568 0 _0183_
rlabel metal2 4320 28434 4320 28434 0 _0184_
rlabel metal2 3977 28476 3977 28476 0 _0185_
rlabel metal2 3840 28140 3840 28140 0 _0186_
rlabel metal2 14400 19362 14400 19362 0 _0187_
rlabel metal2 14376 19488 14376 19488 0 _0188_
rlabel metal2 15312 19824 15312 19824 0 _0189_
rlabel metal4 15072 19740 15072 19740 0 _0190_
rlabel metal3 15264 19740 15264 19740 0 _0191_
rlabel metal2 15477 21504 15477 21504 0 _0192_
rlabel metal2 15504 21588 15504 21588 0 _0193_
rlabel metal3 16320 20832 16320 20832 0 _0194_
rlabel metal2 15929 21420 15929 21420 0 _0195_
rlabel metal2 15991 19992 15991 19992 0 _0196_
rlabel metal2 18528 36708 18528 36708 0 _0197_
rlabel metal2 15792 35952 15792 35952 0 _0198_
rlabel metal2 15600 35868 15600 35868 0 _0199_
rlabel metal3 18240 35994 18240 35994 0 _0200_
rlabel metal2 18048 36204 18048 36204 0 _0201_
rlabel metal2 16629 35112 16629 35112 0 _0202_
rlabel metal2 16656 35196 16656 35196 0 _0203_
rlabel metal2 17040 34440 17040 34440 0 _0204_
rlabel via2 17477 34524 17477 34524 0 _0205_
rlabel metal2 17520 34188 17520 34188 0 _0206_
rlabel metal3 15456 41538 15456 41538 0 _0207_
rlabel metal2 15576 41244 15576 41244 0 _0208_
rlabel metal2 13440 42462 13440 42462 0 _0209_
rlabel metal3 15936 42756 15936 42756 0 _0210_
rlabel metal2 15243 41412 15243 41412 0 _0211_
rlabel metal2 15483 42000 15483 42000 0 _0212_
rlabel metal2 15312 42042 15312 42042 0 _0213_
rlabel metal2 16224 42084 16224 42084 0 _0214_
rlabel via1 16026 42084 16026 42084 0 _0215_
rlabel metal2 15504 41748 15504 41748 0 _0216_
rlabel metal3 2592 27930 2592 27930 0 _0217_
rlabel metal2 3552 26334 3552 26334 0 _0218_
rlabel metal2 4416 25998 4416 25998 0 _0219_
rlabel metal2 4081 26040 4081 26040 0 _0220_
rlabel via1 4319 26040 4319 26040 0 _0221_
rlabel metal2 4080 23184 4080 23184 0 _0222_
rlabel metal2 5424 27636 5424 27636 0 _0223_
rlabel metal2 4416 27552 4416 27552 0 _0224_
rlabel metal2 5047 27468 5047 27468 0 _0225_
rlabel metal2 4663 25956 4663 25956 0 _0226_
rlabel metal2 20352 22890 20352 22890 0 _0227_
rlabel metal3 19200 22764 19200 22764 0 _0228_
rlabel metal2 19296 22596 19296 22596 0 _0229_
rlabel metal2 20448 21756 20448 21756 0 _0230_
rlabel metal2 20112 22428 20112 22428 0 _0231_
rlabel metal2 18816 18648 18816 18648 0 _0232_
rlabel metal2 18768 22512 18768 22512 0 _0233_
rlabel metal2 19584 23856 19584 23856 0 _0234_
rlabel metal2 19541 23940 19541 23940 0 _0235_
rlabel metal2 19913 22344 19913 22344 0 _0236_
rlabel metal2 13200 30576 13200 30576 0 _0237_
rlabel metal2 14438 30156 14438 30156 0 _0238_
rlabel metal2 14352 28980 14352 28980 0 _0239_
rlabel metal2 15456 29946 15456 29946 0 _0240_
rlabel metal2 14544 29064 14544 29064 0 _0241_
rlabel metal2 14640 29862 14640 29862 0 _0242_
rlabel metal2 14784 29946 14784 29946 0 _0243_
rlabel metal2 15360 31374 15360 31374 0 _0244_
rlabel metal3 14976 30744 14976 30744 0 _0245_
rlabel metal2 14791 28980 14791 28980 0 _0246_
rlabel metal2 12048 39648 12048 39648 0 _0247_
rlabel metal2 13824 39732 13824 39732 0 _0248_
rlabel metal2 13152 40488 13152 40488 0 _0249_
rlabel metal2 14088 39144 14088 39144 0 _0250_
rlabel metal2 13248 40530 13248 40530 0 _0251_
rlabel via2 12660 37464 12660 37464 0 _0252_
rlabel metal3 12768 37674 12768 37674 0 _0253_
rlabel metal2 13920 40152 13920 40152 0 _0254_
rlabel metal2 13056 37422 13056 37422 0 _0255_
rlabel metal2 12864 40614 12864 40614 0 _0256_
rlabel via1 5037 44226 5037 44226 0 _0257_
rlabel metal2 4368 45528 4368 45528 0 _0258_
rlabel metal2 5880 44184 5880 44184 0 _0259_
rlabel metal2 4704 44478 4704 44478 0 _0260_
rlabel via2 6348 44184 6348 44184 0 _0261_
rlabel via1 5514 44226 5514 44226 0 _0262_
rlabel metal2 4656 42924 4656 42924 0 _0263_
rlabel metal2 5419 43554 5419 43554 0 _0264_
rlabel metal2 5184 42924 5184 42924 0 _0265_
rlabel metal2 5520 43470 5520 43470 0 _0266_
rlabel metal4 5520 42840 5520 42840 0 _0267_
rlabel metal2 6048 43680 6048 43680 0 _0268_
rlabel metal2 5712 43512 5712 43512 0 _0269_
rlabel metal2 5305 45654 5305 45654 0 _0270_
rlabel metal3 5184 44436 5184 44436 0 _0271_
rlabel via1 5201 45024 5201 45024 0 _0272_
rlabel metal2 5088 45066 5088 45066 0 _0273_
rlabel via1 5020 45734 5020 45734 0 _0274_
rlabel via1 5724 45696 5724 45696 0 _0275_
rlabel metal2 5472 45780 5472 45780 0 _0276_
rlabel metal2 5952 45276 5952 45276 0 _0277_
rlabel metal3 5760 45612 5760 45612 0 _0278_
rlabel metal2 7584 40362 7584 40362 0 _0279_
rlabel metal2 5784 39648 5784 39648 0 _0280_
rlabel metal2 6994 40530 6994 40530 0 _0281_
rlabel metal2 6312 39648 6312 39648 0 _0282_
rlabel metal2 6624 39186 6624 39186 0 _0283_
rlabel metal2 5928 40992 5928 40992 0 _0284_
rlabel via1 6157 39732 6157 39732 0 _0285_
rlabel via2 7680 40476 7680 40476 0 _0286_
rlabel metal2 7200 38220 7200 38220 0 _0287_
rlabel metal2 5568 38178 5568 38178 0 _0288_
rlabel metal2 6768 38304 6768 38304 0 _0289_
rlabel metal2 5856 38220 5856 38220 0 _0290_
rlabel metal2 5451 38136 5451 38136 0 _0291_
rlabel metal3 6432 40530 6432 40530 0 _0292_
rlabel via1 6249 38976 6249 38976 0 _0293_
rlabel metal3 6144 38640 6144 38640 0 _0294_
rlabel metal2 5243 38220 5243 38220 0 _0295_
rlabel metal2 6672 38136 6672 38136 0 _0296_
rlabel metal2 19416 3192 19416 3192 0 net1
rlabel metal2 15480 13440 15480 13440 0 net10
rlabel metal2 13632 81312 13632 81312 0 net100
rlabel metal2 16176 81312 16176 81312 0 net101
rlabel metal2 2592 93030 2592 93030 0 net102
rlabel metal2 1920 93786 1920 93786 0 net103
rlabel metal3 10656 89250 10656 89250 0 net104
rlabel metal4 1872 89796 1872 89796 0 net105
rlabel metal3 2496 79296 2496 79296 0 net106
rlabel metal3 10752 87066 10752 87066 0 net107
rlabel via2 1632 86520 1632 86520 0 net108
rlabel metal2 1488 90804 1488 90804 0 net109
rlabel metal2 15264 54180 15264 54180 0 net11
rlabel metal2 1536 76776 1536 76776 0 net110
rlabel metal2 8880 74424 8880 74424 0 net111
rlabel metal4 11040 78498 11040 78498 0 net112
rlabel metal2 14400 67704 14400 67704 0 net113
rlabel metal2 9456 58632 9456 58632 0 net114
rlabel metal3 9696 81228 9696 81228 0 net115
rlabel via1 12304 79776 12304 79776 0 net116
rlabel metal2 8520 93912 8520 93912 0 net117
rlabel metal2 10536 94668 10536 94668 0 net118
rlabel metal2 11208 94668 11208 94668 0 net119
rlabel metal4 17616 37212 17616 37212 0 net12
rlabel metal4 12144 94164 12144 94164 0 net120
rlabel metal4 9552 60480 9552 60480 0 net121
rlabel metal3 7824 55524 7824 55524 0 net122
rlabel metal2 12360 94752 12360 94752 0 net123
rlabel metal4 13344 94752 13344 94752 0 net124
rlabel metal3 13056 94206 13056 94206 0 net125
rlabel metal2 5376 38976 5376 38976 0 net126
rlabel metal3 16224 51156 16224 51156 0 net127
rlabel metal2 9384 94668 9384 94668 0 net128
rlabel metal2 6336 41916 6336 41916 0 net129
rlabel metal3 20640 14028 20640 14028 0 net13
rlabel metal2 9768 94668 9768 94668 0 net130
rlabel metal3 19776 50190 19776 50190 0 net131
rlabel metal3 16416 48804 16416 48804 0 net132
rlabel metal2 10872 93912 10872 93912 0 net133
rlabel metal2 9120 58674 9120 58674 0 net134
rlabel metal2 15024 93660 15024 93660 0 net135
rlabel metal2 17184 80388 17184 80388 0 net136
rlabel metal2 13536 94500 13536 94500 0 net137
rlabel metal3 9504 17430 9504 17430 0 net138
rlabel metal2 14520 94752 14520 94752 0 net139
rlabel metal2 18984 4032 18984 4032 0 net14
rlabel metal2 13992 93912 13992 93912 0 net140
rlabel metal2 14760 94668 14760 94668 0 net141
rlabel metal2 10272 36456 10272 36456 0 net142
rlabel metal2 18576 15456 18576 15456 0 net143
rlabel metal4 2448 17976 2448 17976 0 net144
rlabel metal3 13536 38598 13536 38598 0 net145
rlabel metal2 7968 39060 7968 39060 0 net146
rlabel metal2 5592 18564 5592 18564 0 net147
rlabel metal2 18624 41160 18624 41160 0 net148
rlabel metal2 1608 16464 1608 16464 0 net149
rlabel metal2 19656 11172 19656 11172 0 net15
rlabel metal2 7344 38136 7344 38136 0 net150
rlabel metal2 1512 17976 1512 17976 0 net151
rlabel metal2 9576 24780 9576 24780 0 net152
rlabel metal2 1320 18312 1320 18312 0 net153
rlabel metal2 4992 21462 4992 21462 0 net154
rlabel metal2 16608 30534 16608 30534 0 net155
rlabel metal2 1560 13440 1560 13440 0 net156
rlabel metal2 8376 19488 8376 19488 0 net157
rlabel metal2 2280 14112 2280 14112 0 net158
rlabel metal2 1896 14112 1896 14112 0 net159
rlabel metal2 15240 14952 15240 14952 0 net16
rlabel metal2 1992 13860 1992 13860 0 net160
rlabel metal2 2784 39690 2784 39690 0 net161
rlabel metal3 7200 37002 7200 37002 0 net162
rlabel metal2 1800 29316 1800 29316 0 net163
rlabel metal2 5352 34356 5352 34356 0 net164
rlabel metal2 16896 25284 16896 25284 0 net165
rlabel metal2 19392 40404 19392 40404 0 net166
rlabel metal2 1800 25452 1800 25452 0 net167
rlabel metal3 2784 35406 2784 35406 0 net168
rlabel metal2 18864 19236 18864 19236 0 net169
rlabel metal4 18912 21672 18912 21672 0 net17
rlabel metal2 4800 37842 4800 37842 0 net170
rlabel metal2 1584 33180 1584 33180 0 net171
rlabel metal3 4080 33768 4080 33768 0 net172
rlabel metal2 2112 28854 2112 28854 0 net173
rlabel metal2 7248 28392 7248 28392 0 net174
rlabel metal2 19200 35952 19200 35952 0 net175
rlabel metal2 18096 42756 18096 42756 0 net176
rlabel metal2 4920 24780 4920 24780 0 net177
rlabel metal3 20064 21714 20064 21714 0 net178
rlabel metal2 14486 31500 14486 31500 0 net179
rlabel metal2 2400 60144 2400 60144 0 net18
rlabel metal2 1560 23184 1560 23184 0 net180
rlabel metal3 1824 18438 1824 18438 0 net181
rlabel metal2 18720 40446 18720 40446 0 net182
rlabel metal3 13632 37212 13632 37212 0 net183
rlabel metal2 7680 25998 7680 25998 0 net184
rlabel metal3 18528 19068 18528 19068 0 net185
rlabel metal2 14640 34440 14640 34440 0 net186
rlabel metal2 13968 45024 13968 45024 0 net187
rlabel metal2 7536 30660 7536 30660 0 net188
rlabel metal3 1632 20748 1632 20748 0 net189
rlabel metal4 14112 15372 14112 15372 0 net19
rlabel metal2 7104 33390 7104 33390 0 net190
rlabel metal2 13536 38136 13536 38136 0 net191
rlabel metal2 2376 36876 2376 36876 0 net192
rlabel metal2 13440 41916 13440 41916 0 net193
rlabel metal2 3648 38850 3648 38850 0 net194
rlabel metal2 13296 26880 13296 26880 0 net195
rlabel metal2 10704 37464 10704 37464 0 net196
rlabel metal2 1896 39900 1896 39900 0 net197
rlabel metal2 1488 39942 1488 39942 0 net198
rlabel metal2 16752 37464 16752 37464 0 net199
rlabel metal2 19032 4284 19032 4284 0 net2
rlabel metal2 18264 14952 18264 14952 0 net20
rlabel metal2 16656 42000 16656 42000 0 net200
rlabel metal2 9216 29148 9216 29148 0 net201
rlabel metal4 2064 33684 2064 33684 0 net202
rlabel metal2 1656 42840 1656 42840 0 net203
rlabel metal2 1872 39732 1872 39732 0 net204
rlabel metal3 1728 41412 1728 41412 0 net205
rlabel metal2 1992 43260 1992 43260 0 net206
rlabel metal2 2136 43680 2136 43680 0 net207
rlabel metal2 11280 42672 11280 42672 0 net208
rlabel metal2 1608 44352 1608 44352 0 net209
rlabel metal2 20712 13440 20712 13440 0 net21
rlabel metal3 2112 35616 2112 35616 0 net210
rlabel metal3 1248 40908 1248 40908 0 net211
rlabel metal2 2184 34356 2184 34356 0 net212
rlabel metal2 7632 34440 7632 34440 0 net213
rlabel metal2 9072 32928 9072 32928 0 net214
rlabel metal2 1752 34188 1752 34188 0 net215
rlabel metal2 1872 34818 1872 34818 0 net216
rlabel metal2 1944 35028 1944 35028 0 net217
rlabel metal4 1920 33180 1920 33180 0 net218
rlabel metal4 3024 33684 3024 33684 0 net219
rlabel metal2 17016 16464 17016 16464 0 net22
rlabel metal3 2400 35490 2400 35490 0 net220
rlabel metal2 1728 35574 1728 35574 0 net221
rlabel metal2 17400 2100 17400 2100 0 net222
rlabel metal2 8544 17850 8544 17850 0 net223
rlabel metal2 13440 22344 13440 22344 0 net224
rlabel metal2 12384 8694 12384 8694 0 net225
rlabel metal2 1824 1638 1824 1638 0 net226
rlabel metal2 3624 2100 3624 2100 0 net227
rlabel metal2 4680 2856 4680 2856 0 net228
rlabel metal2 4248 2100 4248 2100 0 net229
rlabel metal5 2400 19530 2400 19530 0 net23
rlabel metal2 4968 2772 4968 2772 0 net230
rlabel metal4 2592 48048 2592 48048 0 net231
rlabel metal3 18624 48594 18624 48594 0 net232
rlabel metal2 5304 2100 5304 2100 0 net233
rlabel metal2 5832 2856 5832 2856 0 net234
rlabel metal2 2136 2100 2136 2100 0 net235
rlabel metal2 2424 1680 2424 1680 0 net236
rlabel metal2 3000 1764 3000 1764 0 net237
rlabel metal2 3528 2772 3528 2772 0 net238
rlabel metal2 2712 2100 2712 2100 0 net239
rlabel metal2 17880 16464 17880 16464 0 net24
rlabel metal3 18240 48594 18240 48594 0 net240
rlabel metal2 15888 48048 15888 48048 0 net241
rlabel metal2 4392 2856 4392 2856 0 net242
rlabel metal2 7320 1764 7320 1764 0 net243
rlabel metal2 13632 14070 13632 14070 0 net244
rlabel metal3 13536 12180 13536 12180 0 net245
rlabel metal2 6264 2100 6264 2100 0 net246
rlabel metal2 6648 2100 6648 2100 0 net247
rlabel metal2 18048 69972 18048 69972 0 net248
rlabel metal3 16800 80556 16800 80556 0 net249
rlabel metal3 13344 17976 13344 17976 0 net25
rlabel metal2 6984 2100 6984 2100 0 net250
rlabel metal3 13056 20748 13056 20748 0 net251
rlabel metal2 17424 18648 17424 18648 0 net252
rlabel metal4 20880 22260 20880 22260 0 net253
rlabel metal4 16800 17052 16800 17052 0 net254
rlabel metal3 20160 17094 20160 17094 0 net255
rlabel metal4 8640 20160 8640 20160 0 net256
rlabel metal4 20352 18564 20352 18564 0 net257
rlabel metal4 13248 42840 13248 42840 0 net258
rlabel metal4 3504 53844 3504 53844 0 net259
rlabel metal2 14088 20160 14088 20160 0 net26
rlabel metal2 9312 21126 9312 21126 0 net260
rlabel metal2 8616 29736 8616 29736 0 net261
rlabel metal2 17280 23814 17280 23814 0 net262
rlabel metal3 18144 36960 18144 36960 0 net263
rlabel metal3 16272 39060 16272 39060 0 net264
rlabel metal2 16320 31458 16320 31458 0 net265
rlabel metal2 20496 15288 20496 15288 0 net266
rlabel metal2 16440 34188 16440 34188 0 net267
rlabel metal2 14976 46704 14976 46704 0 net268
rlabel metal3 16320 30870 16320 30870 0 net269
rlabel metal3 2784 59388 2784 59388 0 net27
rlabel metal4 18960 30660 18960 30660 0 net270
rlabel metal4 15504 31416 15504 31416 0 net271
rlabel metal4 8496 82992 8496 82992 0 net272
rlabel metal4 19872 35952 19872 35952 0 net273
rlabel metal3 19776 30618 19776 30618 0 net274
rlabel metal2 17088 56154 17088 56154 0 net275
rlabel metal4 14928 35784 14928 35784 0 net276
rlabel metal4 14880 34524 14880 34524 0 net277
rlabel metal4 12000 40824 12000 40824 0 net278
rlabel metal4 17856 34524 17856 34524 0 net279
rlabel metal2 18024 5040 18024 5040 0 net28
rlabel metal4 17280 33600 17280 33600 0 net280
rlabel metal4 13824 34356 13824 34356 0 net281
rlabel metal2 14400 40320 14400 40320 0 net282
rlabel metal2 14880 40488 14880 40488 0 net283
rlabel metal4 18192 38136 18192 38136 0 net284
rlabel metal4 17520 39732 17520 39732 0 net285
rlabel metal3 18528 39816 18528 39816 0 net286
rlabel metal3 19488 25872 19488 25872 0 net287
rlabel metal3 19440 18480 19440 18480 0 net288
rlabel metal2 20160 33054 20160 33054 0 net289
rlabel metal2 13440 5502 13440 5502 0 net29
rlabel metal4 21312 33180 21312 33180 0 net290
rlabel metal4 9216 29904 9216 29904 0 net291
rlabel metal2 20160 25326 20160 25326 0 net292
rlabel metal4 18432 93156 18432 93156 0 net293
rlabel metal4 19152 34944 19152 34944 0 net294
rlabel metal2 20784 41916 20784 41916 0 net295
rlabel metal2 20592 37968 20592 37968 0 net296
rlabel metal3 19776 45822 19776 45822 0 net297
rlabel metal2 11448 26124 11448 26124 0 net298
rlabel metal4 20352 19824 20352 19824 0 net299
rlabel metal2 10752 19950 10752 19950 0 net3
rlabel metal2 17664 17766 17664 17766 0 net30
rlabel metal2 15600 34944 15600 34944 0 net300
rlabel metal2 20064 49476 20064 49476 0 net301
rlabel metal3 14400 61950 14400 61950 0 net302
rlabel metal4 21024 61194 21024 61194 0 net303
rlabel metal4 17760 51828 17760 51828 0 net304
rlabel metal4 15312 52500 15312 52500 0 net305
rlabel metal2 20160 42714 20160 42714 0 net306
rlabel metal2 9288 53508 9288 53508 0 net307
rlabel metal2 20016 55524 20016 55524 0 net308
rlabel metal4 19056 55524 19056 55524 0 net309
rlabel metal2 16872 5544 16872 5544 0 net31
rlabel metal3 19872 56952 19872 56952 0 net310
rlabel metal3 16416 61740 16416 61740 0 net311
rlabel metal4 17712 56364 17712 56364 0 net312
rlabel metal4 17184 60480 17184 60480 0 net313
rlabel metal3 18336 59976 18336 59976 0 net314
rlabel metal4 13344 58296 13344 58296 0 net315
rlabel metal2 15360 57288 15360 57288 0 net316
rlabel metal2 20352 43428 20352 43428 0 net317
rlabel metal4 18624 64596 18624 64596 0 net318
rlabel metal3 14688 60102 14688 60102 0 net319
rlabel metal2 6960 8736 6960 8736 0 net32
rlabel metal3 19584 45234 19584 45234 0 net320
rlabel metal4 20784 19488 20784 19488 0 net321
rlabel metal4 21216 33306 21216 33306 0 net322
rlabel metal2 15936 45570 15936 45570 0 net323
rlabel metal4 16848 46452 16848 46452 0 net324
rlabel metal2 18768 34188 18768 34188 0 net325
rlabel metal2 15552 62874 15552 62874 0 net326
rlabel metal2 14688 61068 14688 61068 0 net327
rlabel metal2 17064 67620 17064 67620 0 net328
rlabel metal3 21408 79884 21408 79884 0 net329
rlabel metal2 15936 6510 15936 6510 0 net33
rlabel metal2 13896 83580 13896 83580 0 net330
rlabel metal2 2328 87948 2328 87948 0 net331
rlabel metal2 20160 74634 20160 74634 0 net332
rlabel metal3 13824 70140 13824 70140 0 net333
rlabel metal2 15024 73752 15024 73752 0 net334
rlabel metal2 14328 58044 14328 58044 0 net335
rlabel metal2 14688 70308 14688 70308 0 net336
rlabel metal2 18432 75180 18432 75180 0 net337
rlabel metal2 15600 73500 15600 73500 0 net338
rlabel metal2 14760 57960 14760 57960 0 net339
rlabel metal2 1560 75012 1560 75012 0 net34
rlabel metal2 2664 87864 2664 87864 0 net340
rlabel metal2 14880 73080 14880 73080 0 net341
rlabel metal2 17856 76524 17856 76524 0 net342
rlabel metal3 13056 79002 13056 79002 0 net343
rlabel metal2 14496 75222 14496 75222 0 net344
rlabel metal2 19776 79884 19776 79884 0 net345
rlabel metal2 14184 62580 14184 62580 0 net346
rlabel metal2 14184 61068 14184 61068 0 net347
rlabel metal3 15072 78330 15072 78330 0 net348
rlabel metal2 18960 82992 18960 82992 0 net349
rlabel metal2 2112 74970 2112 74970 0 net35
rlabel metal2 17208 55776 17208 55776 0 net350
rlabel metal2 10320 85260 10320 85260 0 net351
rlabel metal2 8088 60312 8088 60312 0 net352
rlabel metal2 14784 64008 14784 64008 0 net353
rlabel metal2 12960 63042 12960 63042 0 net354
rlabel metal3 20160 69846 20160 69846 0 net355
rlabel metal2 1848 54264 1848 54264 0 net356
rlabel metal2 2184 53508 2184 53508 0 net357
rlabel metal2 20064 71484 20064 71484 0 net358
rlabel metal2 16776 67116 16776 67116 0 net359
rlabel metal2 2568 75432 2568 75432 0 net36
rlabel metal2 16344 94836 16344 94836 0 net360
rlabel metal3 19776 94458 19776 94458 0 net361
rlabel metal2 19104 94206 19104 94206 0 net362
rlabel metal2 17688 94164 17688 94164 0 net363
rlabel metal2 19488 94248 19488 94248 0 net364
rlabel metal2 18816 93912 18816 93912 0 net365
rlabel metal2 19896 93912 19896 93912 0 net366
rlabel metal3 16032 88578 16032 88578 0 net367
rlabel metal2 19608 93912 19608 93912 0 net368
rlabel metal3 19584 92526 19584 92526 0 net369
rlabel metal2 7776 78918 7776 78918 0 net37
rlabel metal2 18600 92484 18600 92484 0 net370
rlabel metal2 15936 94584 15936 94584 0 net371
rlabel metal2 17064 90552 17064 90552 0 net372
rlabel metal3 17472 94668 17472 94668 0 net373
rlabel metal2 17760 94836 17760 94836 0 net374
rlabel metal2 20040 64092 20040 64092 0 net375
rlabel metal2 17472 93786 17472 93786 0 net376
rlabel metal2 17376 93702 17376 93702 0 net377
rlabel metal2 19200 93660 19200 93660 0 net378
rlabel metal2 19440 93744 19440 93744 0 net379
rlabel metal3 8832 77952 8832 77952 0 net38
rlabel metal2 10104 56532 10104 56532 0 net380
rlabel metal2 15264 73626 15264 73626 0 net381
rlabel metal2 2160 94416 2160 94416 0 net382
rlabel metal2 2016 93954 2016 93954 0 net383
rlabel metal5 1152 78888 1152 78888 0 net384
rlabel metal2 2400 94122 2400 94122 0 net385
rlabel metal4 1776 94836 1776 94836 0 net386
rlabel metal5 2112 80976 2112 80976 0 net387
rlabel metal5 2496 77616 2496 77616 0 net388
rlabel metal2 12096 73542 12096 73542 0 net389
rlabel metal2 5328 76482 5328 76482 0 net39
rlabel metal2 13752 75432 13752 75432 0 net390
rlabel metal2 10248 76944 10248 76944 0 net391
rlabel metal2 4584 41412 4584 41412 0 net392
rlabel metal2 14616 48888 14616 48888 0 net393
rlabel metal2 12456 42924 12456 42924 0 net394
rlabel metal4 4752 94164 4752 94164 0 net395
rlabel metal4 3696 94836 3696 94836 0 net396
rlabel metal2 19704 48804 19704 48804 0 net397
rlabel metal2 16632 31164 16632 31164 0 net398
rlabel metal2 8952 40236 8952 40236 0 net399
rlabel metal2 17280 14700 17280 14700 0 net4
rlabel metal3 13392 73584 13392 73584 0 net40
rlabel metal2 3240 94332 3240 94332 0 net400
rlabel metal3 17280 37170 17280 37170 0 net401
rlabel metal5 8064 66486 8064 66486 0 net402
rlabel metal2 9336 64092 9336 64092 0 net403
rlabel metal2 17376 93912 17376 93912 0 net404
rlabel metal2 13752 83412 13752 83412 0 net405
rlabel metal2 9192 81480 9192 81480 0 net406
rlabel metal2 3096 5544 3096 5544 0 net407
rlabel metal2 4200 94248 4200 94248 0 net408
rlabel metal2 6528 94206 6528 94206 0 net409
rlabel metal2 3189 54768 3189 54768 0 net41
rlabel metal4 5136 94836 5136 94836 0 net410
rlabel metal2 7320 91308 7320 91308 0 net411
rlabel metal2 6888 92064 6888 92064 0 net412
rlabel metal2 7704 91224 7704 91224 0 net413
rlabel metal2 5256 28560 5256 28560 0 net414
rlabel metal4 14160 35364 14160 35364 0 net415
rlabel metal2 15936 94794 15936 94794 0 net416
rlabel metal2 2160 51198 2160 51198 0 net417
rlabel metal5 1824 59514 1824 59514 0 net418
rlabel metal2 1440 53466 1440 53466 0 net419
rlabel metal2 8016 69888 8016 69888 0 net42
rlabel metal4 5088 63168 5088 63168 0 net420
rlabel metal3 2784 57036 2784 57036 0 net421
rlabel metal2 1440 53886 1440 53886 0 net422
rlabel metal2 1920 50988 1920 50988 0 net423
rlabel metal2 2160 56364 2160 56364 0 net424
rlabel metal3 2544 60480 2544 60480 0 net425
rlabel metal4 13248 63252 13248 63252 0 net426
rlabel metal2 18264 52668 18264 52668 0 net427
rlabel metal2 2592 57120 2592 57120 0 net428
rlabel metal3 2352 62328 2352 62328 0 net429
rlabel metal3 2064 77112 2064 77112 0 net43
rlabel metal2 1824 58716 1824 58716 0 net430
rlabel metal4 1776 59388 1776 59388 0 net431
rlabel metal3 4608 58842 4608 58842 0 net432
rlabel metal2 1440 60228 1440 60228 0 net433
rlabel metal2 14952 61404 14952 61404 0 net434
rlabel metal2 17472 54180 17472 54180 0 net435
rlabel metal2 3672 59556 3672 59556 0 net436
rlabel metal2 3216 68460 3216 68460 0 net437
rlabel metal3 6816 72828 6816 72828 0 net438
rlabel metal2 6600 61740 6600 61740 0 net439
rlabel metal2 15744 78120 15744 78120 0 net44
rlabel metal3 13056 69720 13056 69720 0 net440
rlabel metal4 1392 74172 1392 74172 0 net441
rlabel metal3 2688 69888 2688 69888 0 net442
rlabel metal2 6648 75768 6648 75768 0 net443
rlabel metal2 1440 71526 1440 71526 0 net444
rlabel metal3 1728 72366 1728 72366 0 net445
rlabel metal3 2496 64344 2496 64344 0 net446
rlabel metal2 2208 72114 2208 72114 0 net447
rlabel metal2 16056 70140 16056 70140 0 net448
rlabel metal2 6240 58632 6240 58632 0 net449
rlabel metal2 7824 73668 7824 73668 0 net45
rlabel metal2 14400 65982 14400 65982 0 net450
rlabel metal2 5064 61824 5064 61824 0 net451
rlabel metal2 3648 65436 3648 65436 0 net452
rlabel metal2 13536 68124 13536 68124 0 net453
rlabel metal2 15144 56448 15144 56448 0 net454
rlabel metal2 8184 59556 8184 59556 0 net455
rlabel metal4 15168 62832 15168 62832 0 net456
rlabel metal2 15000 58044 15000 58044 0 net457
rlabel metal2 2208 64470 2208 64470 0 net458
rlabel metal3 1728 66990 1728 66990 0 net459
rlabel metal2 6144 76734 6144 76734 0 net46
rlabel metal2 13824 65226 13824 65226 0 net460
rlabel metal3 9984 63084 9984 63084 0 net461
rlabel metal2 5832 58800 5832 58800 0 net462
rlabel metal2 1440 66066 1440 66066 0 net463
rlabel metal3 1824 65898 1824 65898 0 net464
rlabel metal2 3144 42168 3144 42168 0 net465
rlabel metal4 16944 77700 16944 77700 0 net466
rlabel metal4 14640 14784 14640 14784 0 net467
rlabel metal4 17856 87864 17856 87864 0 net468
rlabel metal4 16752 87948 16752 87948 0 net469
rlabel metal2 6336 75642 6336 75642 0 net47
rlabel metal4 20496 89628 20496 89628 0 net470
rlabel metal3 19392 88746 19392 88746 0 net471
rlabel metal2 17352 37380 17352 37380 0 net472
rlabel metal2 15720 38388 15720 38388 0 net473
rlabel metal3 19008 88830 19008 88830 0 net474
rlabel metal2 17064 34356 17064 34356 0 net475
rlabel metal4 20736 83580 20736 83580 0 net476
rlabel metal4 19344 62832 19344 62832 0 net477
rlabel metal4 14256 38724 14256 38724 0 net478
rlabel metal2 2088 39564 2088 39564 0 net479
rlabel metal3 13536 78120 13536 78120 0 net48
rlabel metal2 13344 40782 13344 40782 0 net480
rlabel metal4 20544 91140 20544 91140 0 net481
rlabel metal4 19104 34272 19104 34272 0 net482
rlabel metal4 19824 55356 19824 55356 0 net483
rlabel metal3 20544 46200 20544 46200 0 net484
rlabel metal2 15336 9660 15336 9660 0 net485
rlabel metal2 16728 40404 16728 40404 0 net486
rlabel metal4 20592 84252 20592 84252 0 net487
rlabel metal5 19728 18076 19728 18076 0 net488
rlabel metal4 21024 35784 21024 35784 0 net489
rlabel metal4 1824 63336 1824 63336 0 net49
rlabel metal4 19728 17976 19728 17976 0 net490
rlabel metal4 20448 86604 20448 86604 0 net491
rlabel metal2 7944 27048 7944 27048 0 net492
rlabel metal4 20160 33348 20160 33348 0 net493
rlabel metal2 2328 21336 2328 21336 0 net494
rlabel metal4 19392 38136 19392 38136 0 net495
rlabel metal5 17856 72744 17856 72744 0 net496
rlabel metal2 7824 31836 7824 31836 0 net497
rlabel metal2 15960 23604 15960 23604 0 net498
rlabel metal3 17664 6510 17664 6510 0 net499
rlabel metal2 14400 7014 14400 7014 0 net5
rlabel metal2 8688 72072 8688 72072 0 net50
rlabel metal2 9648 2604 9648 2604 0 net500
rlabel metal3 2208 43302 2208 43302 0 net501
rlabel metal3 17232 16968 17232 16968 0 net502
rlabel metal5 13056 38368 13056 38368 0 net503
rlabel metal4 9120 19908 9120 19908 0 net504
rlabel metal4 8928 2436 8928 2436 0 net505
rlabel metal4 18288 17892 18288 17892 0 net506
rlabel metal4 14064 17472 14064 17472 0 net507
rlabel metal3 8448 18648 8448 18648 0 net508
rlabel metal2 9696 1848 9696 1848 0 net509
rlabel metal3 12096 71610 12096 71610 0 net51
rlabel metal2 17448 53340 17448 53340 0 net510
rlabel metal4 11808 63672 11808 63672 0 net511
rlabel metal2 12192 2016 12192 2016 0 net512
rlabel metal2 6480 2436 6480 2436 0 net513
rlabel metal4 14112 21672 14112 21672 0 net514
rlabel metal4 15360 3444 15360 3444 0 net515
rlabel metal5 13440 11046 13440 11046 0 net516
rlabel metal2 14328 93912 14328 93912 0 net517
rlabel metal4 14928 83580 14928 83580 0 net518
rlabel metal3 15744 10248 15744 10248 0 net519
rlabel metal3 15648 76944 15648 76944 0 net52
rlabel metal2 14448 2688 14448 2688 0 net520
rlabel metal2 16128 1974 16128 1974 0 net521
rlabel metal2 15312 28812 15312 28812 0 net522
rlabel metal3 16608 17850 16608 17850 0 net523
rlabel metal2 4320 2310 4320 2310 0 net524
rlabel metal2 13344 2688 13344 2688 0 net525
rlabel metal3 14208 2142 14208 2142 0 net526
rlabel metal2 17736 93912 17736 93912 0 net527
rlabel metal2 16584 93912 16584 93912 0 net528
rlabel metal4 14592 2856 14592 2856 0 net529
rlabel metal2 8688 72912 8688 72912 0 net53
rlabel metal2 14976 2016 14976 2016 0 net530
rlabel metal3 14400 5964 14400 5964 0 net531
rlabel metal4 16800 1932 16800 1932 0 net532
rlabel metal4 3456 13188 3456 13188 0 net533
rlabel metal2 14136 17556 14136 17556 0 net534
rlabel metal2 2208 3402 2208 3402 0 net535
rlabel metal2 2592 4158 2592 4158 0 net536
rlabel metal3 2688 7098 2688 7098 0 net537
rlabel metal2 1440 3570 1440 3570 0 net538
rlabel metal2 5184 4956 5184 4956 0 net539
rlabel metal3 2208 80640 2208 80640 0 net54
rlabel metal3 2208 7098 2208 7098 0 net540
rlabel metal2 3360 5670 3360 5670 0 net541
rlabel metal2 2736 4956 2736 4956 0 net542
rlabel metal2 1824 4200 1824 4200 0 net543
rlabel metal2 1728 4242 1728 4242 0 net544
rlabel metal2 5184 7140 5184 7140 0 net545
rlabel metal2 15864 5124 15864 5124 0 net546
rlabel metal3 2400 4704 2400 4704 0 net547
rlabel metal2 5232 6552 5232 6552 0 net548
rlabel metal3 2400 8526 2400 8526 0 net549
rlabel metal3 13728 87402 13728 87402 0 net55
rlabel metal2 1824 5082 1824 5082 0 net550
rlabel metal3 1440 4788 1440 4788 0 net551
rlabel metal2 6024 16044 6024 16044 0 net552
rlabel metal2 10584 16800 10584 16800 0 net553
rlabel metal2 16440 17556 16440 17556 0 net554
rlabel metal2 10272 19320 10272 19320 0 net555
rlabel metal2 14520 13104 14520 13104 0 net556
rlabel metal2 4800 11676 4800 11676 0 net557
rlabel metal4 2976 15414 2976 15414 0 net558
rlabel metal2 5976 9660 5976 9660 0 net559
rlabel metal2 8208 69972 8208 69972 0 net56
rlabel metal2 8448 17052 8448 17052 0 net560
rlabel metal3 14400 16674 14400 16674 0 net561
rlabel metal2 5472 14028 5472 14028 0 net562
rlabel metal2 4560 13188 4560 13188 0 net563
rlabel metal2 1824 11886 1824 11886 0 net564
rlabel metal2 2208 5670 2208 5670 0 net565
rlabel metal2 15048 14532 15048 14532 0 net566
rlabel metal2 8352 13230 8352 13230 0 net567
rlabel metal2 7704 13020 7704 13020 0 net568
rlabel metal2 3744 9534 3744 9534 0 net569
rlabel metal2 18720 74424 18720 74424 0 net57
rlabel metal3 16608 13818 16608 13818 0 net570
rlabel metal3 6624 15372 6624 15372 0 net571
rlabel metal2 2592 6594 2592 6594 0 net572
rlabel metal3 2016 5376 2016 5376 0 net573
rlabel metal3 2112 5124 2112 5124 0 net574
rlabel metal2 1824 6426 1824 6426 0 net575
rlabel metal2 13128 5124 13128 5124 0 net576
rlabel metal3 16416 8778 16416 8778 0 net577
rlabel metal2 5640 16044 5640 16044 0 net578
rlabel metal3 1440 6510 1440 6510 0 net579
rlabel metal2 2400 88578 2400 88578 0 net58
rlabel metal2 14784 6132 14784 6132 0 net580
rlabel metal2 11904 60900 11904 60900 0 net581
rlabel metal2 21423 59892 21423 59892 0 net582
rlabel metal2 19968 59892 19968 59892 0 net583
rlabel metal3 2688 86268 2688 86268 0 net59
rlabel metal2 19272 8652 19272 8652 0 net6
rlabel metal2 8400 57036 8400 57036 0 net60
rlabel metal2 15984 58632 15984 58632 0 net61
rlabel metal2 14400 79044 14400 79044 0 net62
rlabel metal2 3312 60144 3312 60144 0 net623
rlabel metal2 16992 54684 16992 54684 0 net624
rlabel metal2 19200 63126 19200 63126 0 net625
rlabel metal2 4608 56238 4608 56238 0 net626
rlabel metal3 4176 53088 4176 53088 0 net627
rlabel metal2 4320 56280 4320 56280 0 net628
rlabel metal2 18768 63084 18768 63084 0 net629
rlabel metal2 7776 73752 7776 73752 0 net63
rlabel metal5 16032 62034 16032 62034 0 net630
rlabel metal2 8112 72912 8112 72912 0 net631
rlabel metal2 7800 37968 7800 37968 0 net632
rlabel metal2 16896 8820 16896 8820 0 net633
rlabel metal2 18000 18480 18000 18480 0 net634
rlabel metal2 4656 22344 4656 22344 0 net635
rlabel metal2 3552 21462 3552 21462 0 net636
rlabel metal4 5184 20244 5184 20244 0 net637
rlabel metal2 18624 17766 18624 17766 0 net638
rlabel metal2 18432 13104 18432 13104 0 net639
rlabel metal2 8544 62328 8544 62328 0 net64
rlabel metal2 4416 16212 4416 16212 0 net640
rlabel metal2 2496 38178 2496 38178 0 net641
rlabel metal2 2592 41160 2592 41160 0 net642
rlabel metal2 9312 37506 9312 37506 0 net643
rlabel metal2 15360 81228 15360 81228 0 net644
rlabel metal3 9168 63000 9168 63000 0 net645
rlabel metal2 9072 46536 9072 46536 0 net646
rlabel metal3 4512 32298 4512 32298 0 net647
rlabel metal2 13632 21504 13632 21504 0 net648
rlabel metal2 10944 42630 10944 42630 0 net649
rlabel metal3 18144 86310 18144 86310 0 net65
rlabel metal2 15192 36456 15192 36456 0 net650
rlabel metal2 14880 36750 14880 36750 0 net651
rlabel metal2 17616 75264 17616 75264 0 net652
rlabel metal2 18768 79800 18768 79800 0 net653
rlabel metal2 6720 73164 6720 73164 0 net654
rlabel metal2 11856 84336 11856 84336 0 net655
rlabel metal2 12672 77532 12672 77532 0 net656
rlabel metal2 13848 60312 13848 60312 0 net657
rlabel metal3 14688 8022 14688 8022 0 net658
rlabel metal2 16200 19824 16200 19824 0 net659
rlabel metal2 4104 80304 4104 80304 0 net66
rlabel metal2 17088 20076 17088 20076 0 net660
rlabel metal2 15168 8652 15168 8652 0 net661
rlabel metal3 13152 35700 13152 35700 0 net662
rlabel metal2 14640 58632 14640 58632 0 net663
rlabel metal2 11040 75264 11040 75264 0 net664
rlabel metal2 9600 72954 9600 72954 0 net665
rlabel metal2 10272 78288 10272 78288 0 net666
rlabel metal2 12336 53340 12336 53340 0 net667
rlabel metal3 11952 39144 11952 39144 0 net668
rlabel metal2 8208 11760 8208 11760 0 net669
rlabel metal3 13536 86982 13536 86982 0 net67
rlabel metal3 2496 9072 2496 9072 0 net670
rlabel metal3 17472 11088 17472 11088 0 net671
rlabel metal3 16128 11928 16128 11928 0 net672
rlabel metal2 2688 15456 2688 15456 0 net673
rlabel metal3 2784 17472 2784 17472 0 net674
rlabel metal2 2448 75936 2448 75936 0 net675
rlabel metal3 3024 60396 3024 60396 0 net676
rlabel metal2 3360 65394 3360 65394 0 net677
rlabel metal3 2304 54600 2304 54600 0 net678
rlabel metal2 19824 54768 19824 54768 0 net679
rlabel metal3 2832 81984 2832 81984 0 net68
rlabel metal3 1920 13116 1920 13116 0 net680
rlabel metal2 2552 19992 2552 19992 0 net681
rlabel metal2 16752 13272 16752 13272 0 net682
rlabel metal2 18144 11718 18144 11718 0 net683
rlabel metal2 10512 14700 10512 14700 0 net684
rlabel metal2 2544 73752 2544 73752 0 net685
rlabel metal2 2832 57792 2832 57792 0 net686
rlabel metal2 20256 63756 20256 63756 0 net687
rlabel metal2 13872 64680 13872 64680 0 net688
rlabel metal2 13344 63126 13344 63126 0 net689
rlabel metal5 1536 61320 1536 61320 0 net69
rlabel metal2 15264 61656 15264 61656 0 net690
rlabel metal2 10848 17724 10848 17724 0 net691
rlabel metal2 5376 13230 5376 13230 0 net692
rlabel metal4 15552 21336 15552 21336 0 net693
rlabel metal2 3168 25494 3168 25494 0 net694
rlabel metal2 16512 16968 16512 16968 0 net695
rlabel metal3 13056 41034 13056 41034 0 net696
rlabel metal2 5520 60144 5520 60144 0 net697
rlabel metal2 16320 60858 16320 60858 0 net698
rlabel via1 6648 66108 6648 66108 0 net699
rlabel metal3 16320 8904 16320 8904 0 net7
rlabel metal2 16080 56364 16080 56364 0 net70
rlabel metal2 16296 73500 16296 73500 0 net700
rlabel metal2 16224 80514 16224 80514 0 net701
rlabel metal3 13056 56448 13056 56448 0 net702
rlabel metal2 17712 15456 17712 15456 0 net703
rlabel metal2 16296 38052 16296 38052 0 net704
rlabel metal2 9312 30576 9312 30576 0 net705
rlabel metal2 15144 40572 15144 40572 0 net706
rlabel metal2 19248 38892 19248 38892 0 net707
rlabel metal3 15456 40572 15456 40572 0 net708
rlabel metal2 6384 53676 6384 53676 0 net709
rlabel metal2 4680 86016 4680 86016 0 net71
rlabel metal2 9384 88788 9384 88788 0 net710
rlabel metal2 15168 88074 15168 88074 0 net711
rlabel metal2 17952 82824 17952 82824 0 net712
rlabel metal2 13440 60018 13440 60018 0 net713
rlabel metal3 20256 32562 20256 32562 0 net714
rlabel metal4 18192 33180 18192 33180 0 net715
rlabel metal2 19680 20832 19680 20832 0 net716
rlabel metal2 17568 43428 17568 43428 0 net717
rlabel metal2 8832 42000 8832 42000 0 net718
rlabel metal3 14880 55062 14880 55062 0 net719
rlabel metal2 5376 87276 5376 87276 0 net72
rlabel metal2 2784 82866 2784 82866 0 net720
rlabel metal3 13152 89712 13152 89712 0 net721
rlabel metal2 7684 77448 7684 77448 0 net722
rlabel metal2 13824 57792 13824 57792 0 net723
rlabel metal3 12288 57288 12288 57288 0 net724
rlabel metal2 13632 7938 13632 7938 0 net725
rlabel metal2 14304 15456 14304 15456 0 net726
rlabel metal2 7728 16968 7728 16968 0 net727
rlabel metal3 8928 33936 8928 33936 0 net728
rlabel metal2 3984 42672 3984 42672 0 net729
rlabel metal2 3504 81018 3504 81018 0 net73
rlabel metal2 7056 20832 7056 20832 0 net730
rlabel metal2 10848 55734 10848 55734 0 net731
rlabel metal2 18240 70476 18240 70476 0 net732
rlabel metal2 12144 86520 12144 86520 0 net733
rlabel metal3 2784 80052 2784 80052 0 net734
rlabel metal2 10920 81480 10920 81480 0 net735
rlabel metal2 7848 59556 7848 59556 0 net736
rlabel metal2 7872 55566 7872 55566 0 net737
rlabel metal2 12480 13230 12480 13230 0 net738
rlabel metal2 14208 16590 14208 16590 0 net739
rlabel metal2 5208 80640 5208 80640 0 net74
rlabel metal2 10608 42000 10608 42000 0 net740
rlabel metal3 9792 35532 9792 35532 0 net741
rlabel metal2 8952 47796 8952 47796 0 net742
rlabel metal2 18336 51072 18336 51072 0 net743
rlabel metal4 16032 58380 16032 58380 0 net744
rlabel metal2 15408 58128 15408 58128 0 net745
rlabel metal2 10416 81984 10416 81984 0 net746
rlabel metal2 15648 57918 15648 57918 0 net747
rlabel metal2 11496 49644 11496 49644 0 net748
rlabel metal2 11136 47964 11136 47964 0 net749
rlabel metal2 4680 81144 4680 81144 0 net75
rlabel metal2 18768 23016 18768 23016 0 net750
rlabel metal2 1728 14784 1728 14784 0 net751
rlabel metal2 18480 14784 18480 14784 0 net752
rlabel metal2 16320 19320 16320 19320 0 net753
rlabel metal2 12432 20832 12432 20832 0 net754
rlabel metal3 6864 19068 6864 19068 0 net755
rlabel metal2 16848 16296 16848 16296 0 net756
rlabel metal3 17808 17976 17808 17976 0 net757
rlabel metal4 15504 17976 15504 17976 0 net758
rlabel metal4 16224 42672 16224 42672 0 net759
rlabel metal2 1560 84084 1560 84084 0 net76
rlabel metal3 14832 17976 14832 17976 0 net760
rlabel metal2 16224 40698 16224 40698 0 net761
rlabel metal2 1440 42126 1440 42126 0 net762
rlabel metal2 864 41160 864 41160 0 net763
rlabel metal2 13920 33474 13920 33474 0 net764
rlabel metal2 864 15456 864 15456 0 net765
rlabel metal2 18816 13860 18816 13860 0 net766
rlabel metal2 16656 19992 16656 19992 0 net767
rlabel metal3 15024 37296 15024 37296 0 net768
rlabel metal4 14688 38136 14688 38136 0 net769
rlabel metal2 1896 84084 1896 84084 0 net77
rlabel metal2 1920 22932 1920 22932 0 net770
rlabel metal3 13056 17976 13056 17976 0 net771
rlabel metal2 1248 11088 1248 11088 0 net772
rlabel metal3 1968 22512 1968 22512 0 net773
rlabel metal3 1248 18480 1248 18480 0 net774
rlabel metal2 14352 18480 14352 18480 0 net775
rlabel metal3 15072 22554 15072 22554 0 net776
rlabel metal2 13296 6384 13296 6384 0 net777
rlabel metal2 10848 19362 10848 19362 0 net778
rlabel metal2 13104 15456 13104 15456 0 net779
rlabel metal3 15648 84882 15648 84882 0 net78
rlabel metal3 16224 15162 16224 15162 0 net780
rlabel metal3 1920 21588 1920 21588 0 net781
rlabel metal2 15408 57120 15408 57120 0 net782
rlabel metal2 13680 55608 13680 55608 0 net783
rlabel metal3 2112 53718 2112 53718 0 net784
rlabel metal2 1344 73038 1344 73038 0 net785
rlabel metal4 2304 80724 2304 80724 0 net786
rlabel metal3 2016 56322 2016 56322 0 net787
rlabel metal2 18624 57162 18624 57162 0 net788
rlabel metal2 10608 63168 10608 63168 0 net789
rlabel metal2 10200 76860 10200 76860 0 net79
rlabel metal2 7968 61740 7968 61740 0 net790
rlabel metal2 17088 57120 17088 57120 0 net791
rlabel metal2 6480 82572 6480 82572 0 net792
rlabel metal2 1488 63840 1488 63840 0 net793
rlabel metal2 13368 82236 13368 82236 0 net794
rlabel metal2 16272 63840 16272 63840 0 net795
rlabel metal2 14112 75894 14112 75894 0 net796
rlabel metal2 14304 69888 14304 69888 0 net797
rlabel metal2 6242 56280 6242 56280 0 net798
rlabel metal2 13104 59304 13104 59304 0 net799
rlabel metal2 18528 13272 18528 13272 0 net8
rlabel metal2 2040 85596 2040 85596 0 net80
rlabel metal2 1728 61698 1728 61698 0 net800
rlabel metal2 1344 62328 1344 62328 0 net801
rlabel metal2 17088 63168 17088 63168 0 net802
rlabel metal2 19200 60144 19200 60144 0 net803
rlabel metal2 16560 59304 16560 59304 0 net804
rlabel metal4 16656 82068 16656 82068 0 net805
rlabel metal2 13824 57666 13824 57666 0 net806
rlabel metal2 10272 74256 10272 74256 0 net807
rlabel metal2 1536 69216 1536 69216 0 net808
rlabel metal2 3936 55650 3936 55650 0 net809
rlabel metal2 18528 82068 18528 82068 0 net81
rlabel metal2 1296 56280 1296 56280 0 net810
rlabel metal2 19056 58632 19056 58632 0 net811
rlabel metal2 16704 57792 16704 57792 0 net812
rlabel metal2 13776 61656 13776 61656 0 net813
rlabel metal2 14784 79842 14784 79842 0 net82
rlabel metal2 14424 83580 14424 83580 0 net83
rlabel metal2 1488 91602 1488 91602 0 net84
rlabel metal3 1632 90678 1632 90678 0 net85
rlabel metal2 2760 90888 2760 90888 0 net86
rlabel metal3 1632 77952 1632 77952 0 net87
rlabel metal5 2688 76902 2688 76902 0 net88
rlabel metal3 12192 63042 12192 63042 0 net89
rlabel metal2 19752 8904 19752 8904 0 net9
rlabel metal2 11760 64596 11760 64596 0 net90
rlabel metal2 18000 78960 18000 78960 0 net91
rlabel metal2 15096 73668 15096 73668 0 net92
rlabel metal3 2352 80724 2352 80724 0 net93
rlabel metal2 1488 92316 1488 92316 0 net94
rlabel metal2 1536 82740 1536 82740 0 net95
rlabel via2 2016 81984 2016 81984 0 net96
rlabel metal4 2736 83412 2736 83412 0 net97
rlabel metal4 9504 83748 9504 83748 0 net98
rlabel metal3 1680 83520 1680 83520 0 net99
<< properties >>
string FIXED_BBOX 0 0 21600 96768
<< end >>
