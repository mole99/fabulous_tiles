module IHP_SRAM (ADDR_SRAM0,
    ADDR_SRAM1,
    ADDR_SRAM2,
    ADDR_SRAM3,
    ADDR_SRAM4,
    ADDR_SRAM5,
    ADDR_SRAM6,
    ADDR_SRAM7,
    ADDR_SRAM8,
    ADDR_SRAM9,
    BM_SRAM0,
    BM_SRAM1,
    BM_SRAM10,
    BM_SRAM11,
    BM_SRAM12,
    BM_SRAM13,
    BM_SRAM14,
    BM_SRAM15,
    BM_SRAM16,
    BM_SRAM17,
    BM_SRAM18,
    BM_SRAM19,
    BM_SRAM2,
    BM_SRAM20,
    BM_SRAM21,
    BM_SRAM22,
    BM_SRAM23,
    BM_SRAM24,
    BM_SRAM25,
    BM_SRAM26,
    BM_SRAM27,
    BM_SRAM28,
    BM_SRAM29,
    BM_SRAM3,
    BM_SRAM30,
    BM_SRAM31,
    BM_SRAM4,
    BM_SRAM5,
    BM_SRAM6,
    BM_SRAM7,
    BM_SRAM8,
    BM_SRAM9,
    CLK_SRAM,
    CONFIGURED_top,
    DIN_SRAM0,
    DIN_SRAM1,
    DIN_SRAM10,
    DIN_SRAM11,
    DIN_SRAM12,
    DIN_SRAM13,
    DIN_SRAM14,
    DIN_SRAM15,
    DIN_SRAM16,
    DIN_SRAM17,
    DIN_SRAM18,
    DIN_SRAM19,
    DIN_SRAM2,
    DIN_SRAM20,
    DIN_SRAM21,
    DIN_SRAM22,
    DIN_SRAM23,
    DIN_SRAM24,
    DIN_SRAM25,
    DIN_SRAM26,
    DIN_SRAM27,
    DIN_SRAM28,
    DIN_SRAM29,
    DIN_SRAM3,
    DIN_SRAM30,
    DIN_SRAM31,
    DIN_SRAM4,
    DIN_SRAM5,
    DIN_SRAM6,
    DIN_SRAM7,
    DIN_SRAM8,
    DIN_SRAM9,
    DOUT_SRAM0,
    DOUT_SRAM1,
    DOUT_SRAM10,
    DOUT_SRAM11,
    DOUT_SRAM12,
    DOUT_SRAM13,
    DOUT_SRAM14,
    DOUT_SRAM15,
    DOUT_SRAM16,
    DOUT_SRAM17,
    DOUT_SRAM18,
    DOUT_SRAM19,
    DOUT_SRAM2,
    DOUT_SRAM20,
    DOUT_SRAM21,
    DOUT_SRAM22,
    DOUT_SRAM23,
    DOUT_SRAM24,
    DOUT_SRAM25,
    DOUT_SRAM26,
    DOUT_SRAM27,
    DOUT_SRAM28,
    DOUT_SRAM29,
    DOUT_SRAM3,
    DOUT_SRAM30,
    DOUT_SRAM31,
    DOUT_SRAM4,
    DOUT_SRAM5,
    DOUT_SRAM6,
    DOUT_SRAM7,
    DOUT_SRAM8,
    DOUT_SRAM9,
    MEN_SRAM,
    REN_SRAM,
    TIE_HIGH_SRAM,
    TIE_LOW_SRAM,
    Tile_X0Y0_UserCLKo,
    Tile_X0Y1_UserCLK,
    WEN_SRAM,
    Tile_X0Y0_E1END,
    Tile_X0Y0_E2END,
    Tile_X0Y0_E2MID,
    Tile_X0Y0_E6END,
    Tile_X0Y0_EE4END,
    Tile_X0Y0_FrameData,
    Tile_X0Y0_FrameData_O,
    Tile_X0Y0_FrameStrobe_O,
    Tile_X0Y0_N1BEG,
    Tile_X0Y0_N2BEG,
    Tile_X0Y0_N2BEGb,
    Tile_X0Y0_N4BEG,
    Tile_X0Y0_S1END,
    Tile_X0Y0_S2END,
    Tile_X0Y0_S2MID,
    Tile_X0Y0_S4END,
    Tile_X0Y0_W1BEG,
    Tile_X0Y0_W2BEG,
    Tile_X0Y0_W2BEGb,
    Tile_X0Y0_W6BEG,
    Tile_X0Y0_WW4BEG,
    Tile_X0Y1_E1END,
    Tile_X0Y1_E2END,
    Tile_X0Y1_E2MID,
    Tile_X0Y1_E6END,
    Tile_X0Y1_EE4END,
    Tile_X0Y1_FrameData,
    Tile_X0Y1_FrameData_O,
    Tile_X0Y1_FrameStrobe,
    Tile_X0Y1_N1END,
    Tile_X0Y1_N2END,
    Tile_X0Y1_N2MID,
    Tile_X0Y1_N4END,
    Tile_X0Y1_S1BEG,
    Tile_X0Y1_S2BEG,
    Tile_X0Y1_S2BEGb,
    Tile_X0Y1_S4BEG,
    Tile_X0Y1_W1BEG,
    Tile_X0Y1_W2BEG,
    Tile_X0Y1_W2BEGb,
    Tile_X0Y1_W6BEG,
    Tile_X0Y1_WW4BEG);
 output ADDR_SRAM0;
 output ADDR_SRAM1;
 output ADDR_SRAM2;
 output ADDR_SRAM3;
 output ADDR_SRAM4;
 output ADDR_SRAM5;
 output ADDR_SRAM6;
 output ADDR_SRAM7;
 output ADDR_SRAM8;
 output ADDR_SRAM9;
 output BM_SRAM0;
 output BM_SRAM1;
 output BM_SRAM10;
 output BM_SRAM11;
 output BM_SRAM12;
 output BM_SRAM13;
 output BM_SRAM14;
 output BM_SRAM15;
 output BM_SRAM16;
 output BM_SRAM17;
 output BM_SRAM18;
 output BM_SRAM19;
 output BM_SRAM2;
 output BM_SRAM20;
 output BM_SRAM21;
 output BM_SRAM22;
 output BM_SRAM23;
 output BM_SRAM24;
 output BM_SRAM25;
 output BM_SRAM26;
 output BM_SRAM27;
 output BM_SRAM28;
 output BM_SRAM29;
 output BM_SRAM3;
 output BM_SRAM30;
 output BM_SRAM31;
 output BM_SRAM4;
 output BM_SRAM5;
 output BM_SRAM6;
 output BM_SRAM7;
 output BM_SRAM8;
 output BM_SRAM9;
 output CLK_SRAM;
 input CONFIGURED_top;
 output DIN_SRAM0;
 output DIN_SRAM1;
 output DIN_SRAM10;
 output DIN_SRAM11;
 output DIN_SRAM12;
 output DIN_SRAM13;
 output DIN_SRAM14;
 output DIN_SRAM15;
 output DIN_SRAM16;
 output DIN_SRAM17;
 output DIN_SRAM18;
 output DIN_SRAM19;
 output DIN_SRAM2;
 output DIN_SRAM20;
 output DIN_SRAM21;
 output DIN_SRAM22;
 output DIN_SRAM23;
 output DIN_SRAM24;
 output DIN_SRAM25;
 output DIN_SRAM26;
 output DIN_SRAM27;
 output DIN_SRAM28;
 output DIN_SRAM29;
 output DIN_SRAM3;
 output DIN_SRAM30;
 output DIN_SRAM31;
 output DIN_SRAM4;
 output DIN_SRAM5;
 output DIN_SRAM6;
 output DIN_SRAM7;
 output DIN_SRAM8;
 output DIN_SRAM9;
 input DOUT_SRAM0;
 input DOUT_SRAM1;
 input DOUT_SRAM10;
 input DOUT_SRAM11;
 input DOUT_SRAM12;
 input DOUT_SRAM13;
 input DOUT_SRAM14;
 input DOUT_SRAM15;
 input DOUT_SRAM16;
 input DOUT_SRAM17;
 input DOUT_SRAM18;
 input DOUT_SRAM19;
 input DOUT_SRAM2;
 input DOUT_SRAM20;
 input DOUT_SRAM21;
 input DOUT_SRAM22;
 input DOUT_SRAM23;
 input DOUT_SRAM24;
 input DOUT_SRAM25;
 input DOUT_SRAM26;
 input DOUT_SRAM27;
 input DOUT_SRAM28;
 input DOUT_SRAM29;
 input DOUT_SRAM3;
 input DOUT_SRAM30;
 input DOUT_SRAM31;
 input DOUT_SRAM4;
 input DOUT_SRAM5;
 input DOUT_SRAM6;
 input DOUT_SRAM7;
 input DOUT_SRAM8;
 input DOUT_SRAM9;
 output MEN_SRAM;
 output REN_SRAM;
 output TIE_HIGH_SRAM;
 output TIE_LOW_SRAM;
 output Tile_X0Y0_UserCLKo;
 input Tile_X0Y1_UserCLK;
 output WEN_SRAM;
 input [3:0] Tile_X0Y0_E1END;
 input [7:0] Tile_X0Y0_E2END;
 input [7:0] Tile_X0Y0_E2MID;
 input [11:0] Tile_X0Y0_E6END;
 input [15:0] Tile_X0Y0_EE4END;
 input [31:0] Tile_X0Y0_FrameData;
 output [31:0] Tile_X0Y0_FrameData_O;
 output [19:0] Tile_X0Y0_FrameStrobe_O;
 output [3:0] Tile_X0Y0_N1BEG;
 output [7:0] Tile_X0Y0_N2BEG;
 output [7:0] Tile_X0Y0_N2BEGb;
 output [15:0] Tile_X0Y0_N4BEG;
 input [3:0] Tile_X0Y0_S1END;
 input [7:0] Tile_X0Y0_S2END;
 input [7:0] Tile_X0Y0_S2MID;
 input [15:0] Tile_X0Y0_S4END;
 output [3:0] Tile_X0Y0_W1BEG;
 output [7:0] Tile_X0Y0_W2BEG;
 output [7:0] Tile_X0Y0_W2BEGb;
 output [11:0] Tile_X0Y0_W6BEG;
 output [15:0] Tile_X0Y0_WW4BEG;
 input [3:0] Tile_X0Y1_E1END;
 input [7:0] Tile_X0Y1_E2END;
 input [7:0] Tile_X0Y1_E2MID;
 input [11:0] Tile_X0Y1_E6END;
 input [15:0] Tile_X0Y1_EE4END;
 input [31:0] Tile_X0Y1_FrameData;
 output [31:0] Tile_X0Y1_FrameData_O;
 input [19:0] Tile_X0Y1_FrameStrobe;
 input [3:0] Tile_X0Y1_N1END;
 input [7:0] Tile_X0Y1_N2END;
 input [7:0] Tile_X0Y1_N2MID;
 input [15:0] Tile_X0Y1_N4END;
 output [3:0] Tile_X0Y1_S1BEG;
 output [7:0] Tile_X0Y1_S2BEG;
 output [7:0] Tile_X0Y1_S2BEGb;
 output [15:0] Tile_X0Y1_S4BEG;
 output [3:0] Tile_X0Y1_W1BEG;
 output [7:0] Tile_X0Y1_W2BEG;
 output [7:0] Tile_X0Y1_W2BEGb;
 output [11:0] Tile_X0Y1_W6BEG;
 output [15:0] Tile_X0Y1_WW4BEG;

 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net583;
 wire net328;
 wire net329;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire net368;
 wire net369;
 wire net370;
 wire net371;
 wire net372;
 wire net373;
 wire net374;
 wire net375;
 wire net376;
 wire net377;
 wire net378;
 wire net379;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame0_bit0.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame0_bit1.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame0_bit10.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame0_bit11.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame0_bit12.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame0_bit13.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame0_bit14.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame0_bit15.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame0_bit16.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame0_bit17.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame0_bit18.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame0_bit19.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame0_bit2.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame0_bit20.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame0_bit21.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame0_bit22.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame0_bit23.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame0_bit24.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame0_bit25.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame0_bit26.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame0_bit27.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame0_bit28.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame0_bit29.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame0_bit3.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame0_bit30.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame0_bit31.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame0_bit4.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame0_bit5.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame0_bit6.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame0_bit7.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame0_bit8.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame0_bit9.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame1_bit0.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame1_bit1.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame1_bit10.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame1_bit11.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame1_bit12.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame1_bit13.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame1_bit14.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame1_bit15.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame1_bit16.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame1_bit17.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame1_bit18.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame1_bit19.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame1_bit2.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame1_bit20.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame1_bit21.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame1_bit22.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame1_bit23.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame1_bit24.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame1_bit25.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame1_bit26.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame1_bit27.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame1_bit28.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame1_bit29.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame1_bit3.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame1_bit30.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame1_bit31.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame1_bit4.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame1_bit5.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame1_bit6.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame1_bit7.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame1_bit8.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame1_bit9.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame2_bit0.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame2_bit1.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame2_bit10.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame2_bit11.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame2_bit12.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame2_bit13.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame2_bit14.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame2_bit15.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame2_bit16.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame2_bit17.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame2_bit18.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame2_bit19.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame2_bit2.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame2_bit20.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame2_bit21.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame2_bit22.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame2_bit23.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame2_bit24.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame2_bit25.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame2_bit26.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame2_bit27.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame2_bit28.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame2_bit29.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame2_bit3.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame2_bit30.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame2_bit31.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame2_bit4.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame2_bit5.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame2_bit6.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame2_bit7.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame2_bit8.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame2_bit9.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame3_bit0.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame3_bit1.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame3_bit10.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame3_bit11.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame3_bit12.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame3_bit13.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame3_bit14.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame3_bit15.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame3_bit16.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame3_bit17.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame3_bit18.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame3_bit19.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame3_bit2.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame3_bit20.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame3_bit21.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame3_bit22.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame3_bit23.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame3_bit24.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame3_bit25.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame3_bit26.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame3_bit27.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame3_bit28.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame3_bit29.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame3_bit3.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame3_bit30.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame3_bit31.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame3_bit4.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame3_bit5.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame3_bit6.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame3_bit7.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame3_bit8.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame3_bit9.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame4_bit0.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame4_bit1.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame4_bit10.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame4_bit11.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame4_bit12.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame4_bit13.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame4_bit14.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame4_bit15.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame4_bit16.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame4_bit17.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame4_bit18.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame4_bit19.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame4_bit2.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame4_bit20.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame4_bit21.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame4_bit22.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame4_bit23.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame4_bit24.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame4_bit25.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame4_bit26.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame4_bit27.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame4_bit28.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame4_bit29.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame4_bit3.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame4_bit30.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame4_bit31.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame4_bit4.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame4_bit5.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame4_bit6.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame4_bit7.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame4_bit8.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame4_bit9.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame5_bit0.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame5_bit1.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame5_bit10.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame5_bit11.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame5_bit12.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame5_bit13.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame5_bit14.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame5_bit15.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame5_bit16.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame5_bit17.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame5_bit18.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame5_bit19.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame5_bit2.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame5_bit20.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame5_bit21.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame5_bit22.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame5_bit23.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame5_bit24.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame5_bit25.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame5_bit26.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame5_bit27.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame5_bit28.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame5_bit29.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame5_bit3.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame5_bit30.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame5_bit31.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame5_bit4.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame5_bit5.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame5_bit6.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame5_bit7.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame5_bit8.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame5_bit9.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame6_bit0.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame6_bit1.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame6_bit10.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame6_bit11.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame6_bit12.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame6_bit13.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame6_bit14.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame6_bit15.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame6_bit16.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame6_bit17.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame6_bit18.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame6_bit19.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame6_bit2.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame6_bit20.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame6_bit21.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame6_bit22.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame6_bit23.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame6_bit24.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame6_bit25.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame6_bit26.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame6_bit27.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame6_bit28.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame6_bit29.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame6_bit3.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame6_bit30.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame6_bit31.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame6_bit4.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame6_bit5.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame6_bit6.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame6_bit7.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame6_bit8.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame6_bit9.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit0.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit1.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit10.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit11.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit12.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit13.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit14.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit15.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit16.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit17.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit18.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit19.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit2.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit20.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit21.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit22.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit23.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit24.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit25.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit26.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit27.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit28.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit29.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit3.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit30.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit31.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit4.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit5.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit6.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit7.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit8.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit9.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit0.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit1.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit10.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit11.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit12.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit13.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit14.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit15.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit16.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit17.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit18.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit19.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit2.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit20.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit21.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit22.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit23.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit24.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit25.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit26.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit27.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit28.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit29.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit3.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit30.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit31.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit4.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit5.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit6.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit7.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit8.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit9.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame9_bit22.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame9_bit23.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame9_bit24.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame9_bit25.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame9_bit26.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame9_bit27.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame9_bit28.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame9_bit29.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame9_bit30.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame9_bit31.Q ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS2_BEG0 ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS2_BEG1 ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS2_BEG2 ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS2_BEG3 ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS2_BEG4 ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS2_BEG5 ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS2_BEG6 ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS2_BEG7 ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG0 ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG1 ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG10 ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG11 ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG12 ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG13 ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG14 ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG15 ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG2 ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG3 ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG4 ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG5 ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG6 ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG7 ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG8 ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG9 ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.N1BEG0 ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.N1BEG1 ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.N1BEG2 ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.N1BEG3 ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.N1END0 ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.N1END1 ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.N1END2 ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.N1END3 ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.N2BEG0 ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.N2BEG1 ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.N2BEG2 ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.N2BEG3 ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.N2BEG4 ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.N2BEG5 ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.N2BEG6 ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.N2BEG7 ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.N2BEGb0 ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.N2BEGb1 ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.N2BEGb2 ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.N2BEGb3 ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.N2BEGb4 ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.N2BEGb5 ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.N2BEGb6 ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.N2BEGb7 ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.N4BEG0 ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.N4BEG1 ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.N4BEG2 ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.N4BEG3 ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.S2BEG0 ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.S2BEG1 ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.S2BEG2 ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.S2BEG3 ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.S2BEG4 ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.S2BEG5 ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.S2BEG6 ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.S2BEG7 ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.S4BEG0 ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.S4BEG1 ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.S4BEG2 ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.S4BEG3 ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.W1BEG0 ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.W1BEG1 ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.W1BEG2 ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.W1BEG3 ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.W2BEG0 ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.W2BEG1 ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.W2BEG2 ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.W2BEG3 ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.W2BEG4 ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.W2BEG5 ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.W2BEG6 ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.W2BEG7 ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.W2BEGb0 ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.W2BEGb1 ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.W2BEGb2 ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.W2BEGb3 ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.W2BEGb4 ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.W2BEGb5 ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.W2BEGb6 ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.W2BEGb7 ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.W6BEG0 ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.W6BEG1 ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.W6BEG10 ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.W6BEG11 ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.W6BEG2 ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.W6BEG3 ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.W6BEG4 ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.W6BEG5 ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.W6BEG6 ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.W6BEG7 ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.W6BEG8 ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.W6BEG9 ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.WW4BEG0 ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.WW4BEG1 ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.WW4BEG10 ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.WW4BEG11 ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.WW4BEG12 ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.WW4BEG13 ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.WW4BEG14 ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.WW4BEG15 ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.WW4BEG2 ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.WW4BEG3 ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.WW4BEG4 ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.WW4BEG5 ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.WW4BEG6 ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.WW4BEG7 ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.WW4BEG8 ;
 wire \Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.WW4BEG9 ;
 wire \Tile_X0Y0_IHP_SRAM_top.N4BEG_outbuf_10.A ;
 wire \Tile_X0Y0_IHP_SRAM_top.N4BEG_outbuf_11.A ;
 wire \Tile_X0Y0_IHP_SRAM_top.N4BEG_outbuf_8.A ;
 wire \Tile_X0Y0_IHP_SRAM_top.N4BEG_outbuf_9.A ;
 wire net380;
 wire net381;
 wire net382;
 wire net383;
 wire net384;
 wire net385;
 wire net386;
 wire net387;
 wire net388;
 wire net389;
 wire net390;
 wire net391;
 wire net392;
 wire net393;
 wire net394;
 wire net395;
 wire net396;
 wire net397;
 wire net398;
 wire net399;
 wire net400;
 wire net401;
 wire net402;
 wire net403;
 wire net404;
 wire net405;
 wire net406;
 wire net407;
 wire net408;
 wire net409;
 wire net410;
 wire net411;
 wire net412;
 wire net413;
 wire net414;
 wire net415;
 wire net416;
 wire net417;
 wire net418;
 wire net419;
 wire net420;
 wire net421;
 wire net422;
 wire net423;
 wire net424;
 wire net425;
 wire net426;
 wire net427;
 wire net428;
 wire net429;
 wire net430;
 wire net431;
 wire net432;
 wire net433;
 wire net434;
 wire net435;
 wire net436;
 wire net437;
 wire net438;
 wire net439;
 wire net440;
 wire net441;
 wire net442;
 wire net443;
 wire net444;
 wire net445;
 wire net446;
 wire net447;
 wire net448;
 wire net449;
 wire net450;
 wire net451;
 wire net452;
 wire net453;
 wire net454;
 wire net455;
 wire net456;
 wire net457;
 wire net458;
 wire net459;
 wire net460;
 wire net461;
 wire net462;
 wire net463;
 wire net464;
 wire net465;
 wire net466;
 wire net467;
 wire net468;
 wire net469;
 wire net470;
 wire net471;
 wire net472;
 wire net473;
 wire net474;
 wire net475;
 wire net476;
 wire net477;
 wire net478;
 wire net479;
 wire net480;
 wire net481;
 wire net482;
 wire net483;
 wire net484;
 wire net485;
 wire net486;
 wire net487;
 wire net488;
 wire net489;
 wire net490;
 wire net491;
 wire net492;
 wire net493;
 wire net494;
 wire net495;
 wire net496;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame0_bit0.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame0_bit1.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame0_bit10.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame0_bit11.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame0_bit12.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame0_bit13.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame0_bit14.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame0_bit15.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame0_bit16.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame0_bit17.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame0_bit18.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame0_bit19.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame0_bit2.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame0_bit20.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame0_bit21.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame0_bit22.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame0_bit23.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame0_bit24.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame0_bit25.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame0_bit26.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame0_bit27.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame0_bit28.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame0_bit29.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame0_bit3.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame0_bit30.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame0_bit31.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame0_bit4.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame0_bit5.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame0_bit6.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame0_bit7.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame0_bit8.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame0_bit9.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit0.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit1.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit10.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit11.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit12.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit13.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit14.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit15.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit16.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit17.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit18.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit19.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit2.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit20.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit21.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit22.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit23.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit24.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit25.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit26.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit27.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit28.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit29.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit3.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit30.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit31.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit4.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit5.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit6.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit7.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit8.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit9.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit0.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit1.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit10.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit11.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit12.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit13.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit14.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit15.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit16.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit17.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit18.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit19.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit2.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit20.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit21.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit22.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit23.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit24.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit25.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit26.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit27.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit28.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit29.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit3.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit30.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit31.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit4.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit5.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit6.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit7.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit8.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit9.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame3_bit0.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame3_bit1.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame3_bit10.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame3_bit11.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame3_bit12.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame3_bit13.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame3_bit14.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame3_bit15.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame3_bit16.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame3_bit17.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame3_bit18.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame3_bit19.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame3_bit2.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame3_bit20.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame3_bit21.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame3_bit22.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame3_bit23.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame3_bit24.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame3_bit25.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame3_bit26.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame3_bit27.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame3_bit28.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame3_bit29.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame3_bit3.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame3_bit30.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame3_bit31.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame3_bit4.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame3_bit5.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame3_bit6.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame3_bit7.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame3_bit8.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame3_bit9.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame4_bit0.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame4_bit1.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame4_bit10.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame4_bit11.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame4_bit12.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame4_bit13.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame4_bit14.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame4_bit15.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame4_bit16.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame4_bit17.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame4_bit18.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame4_bit19.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame4_bit2.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame4_bit20.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame4_bit21.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame4_bit22.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame4_bit23.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame4_bit24.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame4_bit25.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame4_bit26.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame4_bit27.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame4_bit28.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame4_bit29.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame4_bit3.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame4_bit30.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame4_bit31.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame4_bit4.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame4_bit5.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame4_bit6.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame4_bit7.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame4_bit8.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame4_bit9.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame5_bit0.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame5_bit1.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame5_bit10.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame5_bit11.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame5_bit12.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame5_bit13.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame5_bit14.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame5_bit15.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame5_bit16.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame5_bit17.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame5_bit18.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame5_bit19.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame5_bit2.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame5_bit20.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame5_bit21.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame5_bit22.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame5_bit23.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame5_bit24.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame5_bit25.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame5_bit26.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame5_bit27.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame5_bit28.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame5_bit29.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame5_bit3.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame5_bit30.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame5_bit31.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame5_bit4.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame5_bit5.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame5_bit6.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame5_bit7.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame5_bit8.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame5_bit9.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame6_bit0.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame6_bit1.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame6_bit10.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame6_bit11.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame6_bit12.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame6_bit13.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame6_bit14.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame6_bit15.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame6_bit16.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame6_bit17.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame6_bit18.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame6_bit19.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame6_bit2.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame6_bit20.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame6_bit21.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame6_bit22.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame6_bit23.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame6_bit24.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame6_bit25.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame6_bit26.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame6_bit27.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame6_bit28.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame6_bit29.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame6_bit3.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame6_bit30.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame6_bit31.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame6_bit4.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame6_bit5.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame6_bit6.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame6_bit7.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame6_bit8.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame6_bit9.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit0.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit1.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit10.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit11.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit12.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit13.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit14.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit15.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit16.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit17.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit18.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit19.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit2.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit20.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit21.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit22.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit23.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit24.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit25.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit26.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit27.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit28.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit29.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit3.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit30.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit31.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit4.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit5.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit6.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit7.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit8.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit9.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit0.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit1.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit10.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit11.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit12.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit13.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit14.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit15.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit16.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit17.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit18.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit19.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit2.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit20.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit21.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit22.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit23.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit24.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit25.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit26.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit27.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit28.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit29.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit3.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit30.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit31.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit4.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit5.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit6.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit7.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit8.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit9.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame9_bit10.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame9_bit11.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame9_bit12.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame9_bit13.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame9_bit14.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame9_bit15.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame9_bit16.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame9_bit17.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame9_bit18.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame9_bit19.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame9_bit20.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame9_bit21.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame9_bit22.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame9_bit23.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame9_bit24.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame9_bit25.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame9_bit26.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame9_bit27.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame9_bit28.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame9_bit29.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame9_bit30.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame9_bit31.Q ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.J_NS4_BEG10 ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.J_NS4_BEG11 ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.J_NS4_BEG12 ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.J_NS4_BEG13 ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.J_NS4_BEG14 ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.J_NS4_BEG15 ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.J_NS4_BEG4 ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.J_NS4_BEG5 ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.J_NS4_BEG6 ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.J_NS4_BEG7 ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.J_NS4_BEG8 ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.J_NS4_BEG9 ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.S1BEG0 ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.S1BEG1 ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.S1BEG2 ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.S1BEG3 ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.S2BEG0 ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.S2BEG1 ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.S2BEG2 ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.S2BEG3 ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.S2BEG4 ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.S2BEG5 ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.S2BEG6 ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.S2BEG7 ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.S4BEG0 ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.S4BEG1 ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.S4BEG2 ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.S4BEG3 ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.W1BEG0 ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.W1BEG1 ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.W1BEG2 ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.W1BEG3 ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.W2BEG0 ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.W2BEG1 ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.W2BEG2 ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.W2BEG3 ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.W2BEG4 ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.W2BEG5 ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.W2BEG6 ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.W2BEG7 ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.W2BEGb0 ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.W2BEGb1 ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.W2BEGb2 ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.W2BEGb3 ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.W2BEGb4 ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.W2BEGb5 ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.W2BEGb6 ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.W2BEGb7 ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.W6BEG0 ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.W6BEG1 ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.W6BEG10 ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.W6BEG11 ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.W6BEG2 ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.W6BEG3 ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.W6BEG4 ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.W6BEG5 ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.W6BEG6 ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.W6BEG7 ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.W6BEG8 ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.W6BEG9 ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.WW4BEG0 ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.WW4BEG1 ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.WW4BEG10 ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.WW4BEG11 ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.WW4BEG12 ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.WW4BEG13 ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.WW4BEG14 ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.WW4BEG15 ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.WW4BEG2 ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.WW4BEG3 ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.WW4BEG4 ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.WW4BEG5 ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.WW4BEG6 ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.WW4BEG7 ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.WW4BEG8 ;
 wire \Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.WW4BEG9 ;
 wire net497;
 wire net498;
 wire net499;
 wire net500;
 wire net501;
 wire net502;
 wire net503;
 wire net504;
 wire net505;
 wire net506;
 wire net507;
 wire net508;
 wire net509;
 wire net510;
 wire net511;
 wire net512;
 wire net513;
 wire net514;
 wire net515;
 wire net516;
 wire net517;
 wire net518;
 wire net519;
 wire net520;
 wire net521;
 wire net522;
 wire net523;
 wire net524;
 wire net525;
 wire net526;
 wire net527;
 wire net528;
 wire net529;
 wire net530;
 wire net531;
 wire net532;
 wire net533;
 wire net534;
 wire net535;
 wire net536;
 wire net537;
 wire net538;
 wire net539;
 wire net540;
 wire net541;
 wire net542;
 wire net543;
 wire net544;
 wire net545;
 wire net546;
 wire net547;
 wire net548;
 wire net549;
 wire net550;
 wire net551;
 wire net552;
 wire net553;
 wire net554;
 wire net555;
 wire net556;
 wire net557;
 wire net558;
 wire net559;
 wire net560;
 wire net561;
 wire net562;
 wire net563;
 wire net564;
 wire net565;
 wire net566;
 wire net567;
 wire net568;
 wire net569;
 wire net570;
 wire net571;
 wire net572;
 wire net573;
 wire net574;
 wire net575;
 wire net576;
 wire net577;
 wire net578;
 wire net579;
 wire net580;
 wire net581;
 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire net623;
 wire net624;
 wire net625;
 wire net626;
 wire net627;
 wire net628;
 wire net629;
 wire net630;
 wire net631;
 wire net632;
 wire net633;
 wire net634;
 wire net635;
 wire net636;
 wire net637;
 wire net638;
 wire net639;
 wire net640;
 wire net641;
 wire net642;
 wire net643;
 wire net644;
 wire net645;
 wire net646;
 wire net647;
 wire net648;
 wire net649;
 wire net650;
 wire net651;
 wire net652;
 wire net653;
 wire net654;
 wire net655;
 wire net656;
 wire net657;
 wire net658;
 wire net659;
 wire net660;
 wire net661;
 wire net662;
 wire net663;
 wire net664;
 wire net665;
 wire net666;
 wire net667;
 wire net668;
 wire net669;
 wire net670;
 wire net671;
 wire net672;
 wire net673;
 wire net674;
 wire net675;
 wire net676;
 wire net677;
 wire net678;
 wire net679;
 wire net680;
 wire net681;
 wire net682;
 wire net683;
 wire net684;
 wire net685;
 wire net686;
 wire net687;
 wire net688;
 wire net689;
 wire net690;
 wire net691;
 wire net692;
 wire net693;
 wire net694;
 wire net695;
 wire net696;
 wire net697;
 wire net698;
 wire net699;
 wire net700;
 wire net701;
 wire net702;
 wire net703;
 wire net704;
 wire net705;
 wire net706;
 wire net707;
 wire net708;
 wire net709;
 wire net710;
 wire net711;
 wire net712;
 wire net713;
 wire net714;
 wire net715;
 wire net716;
 wire net717;
 wire net718;
 wire net719;
 wire net720;
 wire net721;
 wire net722;
 wire net723;
 wire net724;
 wire net725;
 wire net726;
 wire net727;
 wire net728;
 wire net729;
 wire net730;
 wire net731;
 wire net732;
 wire net733;
 wire net734;
 wire net735;
 wire net736;
 wire net737;
 wire net738;
 wire net739;
 wire net740;
 wire net741;
 wire net742;
 wire net743;
 wire net744;
 wire net745;
 wire net746;
 wire net747;
 wire net748;
 wire net749;
 wire net750;
 wire net751;
 wire net752;
 wire net753;
 wire net754;
 wire net755;
 wire net756;
 wire net757;
 wire net758;
 wire net759;
 wire net760;
 wire net761;
 wire net762;
 wire net763;
 wire net764;
 wire net765;
 wire net766;
 wire net767;
 wire net768;
 wire net769;
 wire net770;
 wire net771;
 wire net772;
 wire net773;
 wire net774;
 wire net775;
 wire net776;
 wire net777;
 wire net778;
 wire net779;
 wire net780;
 wire net781;
 wire net782;
 wire net783;
 wire net784;
 wire net785;
 wire net786;
 wire net787;
 wire net788;
 wire net789;
 wire net790;
 wire net791;
 wire net792;
 wire net793;
 wire net794;
 wire net795;
 wire net796;
 wire net797;
 wire net798;
 wire net799;
 wire net800;
 wire net801;
 wire net802;
 wire net803;
 wire net804;
 wire net805;
 wire net806;
 wire net807;
 wire net808;
 wire net809;
 wire net810;
 wire net811;
 wire net812;
 wire net813;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net250;
 wire net582;

 sg13g2_inv_1 _0297_ (.Y(_0000_),
    .A(net157));
 sg13g2_inv_1 _0298_ (.Y(_0001_),
    .A(net151));
 sg13g2_inv_1 _0299_ (.Y(_0002_),
    .A(net128));
 sg13g2_inv_1 _0300_ (.Y(_0003_),
    .A(net57));
 sg13g2_inv_1 _0301_ (.Y(_0004_),
    .A(net58));
 sg13g2_inv_1 _0302_ (.Y(_0005_),
    .A(net59));
 sg13g2_inv_1 _0303_ (.Y(_0006_),
    .A(net54));
 sg13g2_inv_1 _0304_ (.Y(_0007_),
    .A(net167));
 sg13g2_inv_1 _0305_ (.Y(_0008_),
    .A(net166));
 sg13g2_inv_1 _0306_ (.Y(_0009_),
    .A(net165));
 sg13g2_inv_1 _0307_ (.Y(_0010_),
    .A(net162));
 sg13g2_inv_1 _0308_ (.Y(_0011_),
    .A(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit15.Q ));
 sg13g2_inv_1 _0309_ (.Y(_0012_),
    .A(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit18.Q ));
 sg13g2_inv_1 _0310_ (.Y(_0013_),
    .A(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit21.Q ));
 sg13g2_inv_1 _0311_ (.Y(_0014_),
    .A(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit24.Q ));
 sg13g2_inv_1 _0312_ (.Y(_0015_),
    .A(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit19.Q ));
 sg13g2_inv_1 _0313_ (.Y(_0016_),
    .A(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit22.Q ));
 sg13g2_inv_1 _0314_ (.Y(_0017_),
    .A(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit25.Q ));
 sg13g2_inv_1 _0315_ (.Y(_0018_),
    .A(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit28.Q ));
 sg13g2_inv_1 _0316_ (.Y(_0019_),
    .A(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit2.Q ));
 sg13g2_inv_1 _0317_ (.Y(_0020_),
    .A(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit3.Q ));
 sg13g2_inv_1 _0318_ (.Y(_0021_),
    .A(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit5.Q ));
 sg13g2_inv_1 _0319_ (.Y(_0022_),
    .A(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit6.Q ));
 sg13g2_inv_1 _0320_ (.Y(_0023_),
    .A(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit8.Q ));
 sg13g2_inv_1 _0321_ (.Y(_0024_),
    .A(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit9.Q ));
 sg13g2_inv_1 _0322_ (.Y(_0025_),
    .A(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit11.Q ));
 sg13g2_inv_1 _0323_ (.Y(_0026_),
    .A(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit12.Q ));
 sg13g2_inv_1 _0324_ (.Y(_0027_),
    .A(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit6.Q ));
 sg13g2_inv_1 _0325_ (.Y(_0028_),
    .A(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit7.Q ));
 sg13g2_inv_1 _0326_ (.Y(_0029_),
    .A(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit9.Q ));
 sg13g2_inv_1 _0327_ (.Y(_0030_),
    .A(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit10.Q ));
 sg13g2_inv_1 _0328_ (.Y(_0031_),
    .A(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit12.Q ));
 sg13g2_inv_1 _0329_ (.Y(_0032_),
    .A(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit13.Q ));
 sg13g2_inv_1 _0330_ (.Y(_0033_),
    .A(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit15.Q ));
 sg13g2_inv_1 _0331_ (.Y(_0034_),
    .A(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit16.Q ));
 sg13g2_inv_1 _0332_ (.Y(_0035_),
    .A(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit0.Q ));
 sg13g2_inv_1 _0333_ (.Y(_0036_),
    .A(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit3.Q ));
 sg13g2_inv_1 _0334_ (.Y(_0037_),
    .A(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit5.Q ));
 sg13g2_inv_1 _0335_ (.Y(_0038_),
    .A(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS2_BEG0 ));
 sg13g2_inv_1 _0336_ (.Y(_0039_),
    .A(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS2_BEG1 ));
 sg13g2_inv_1 _0337_ (.Y(_0040_),
    .A(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS2_BEG2 ));
 sg13g2_inv_1 _0338_ (.Y(_0041_),
    .A(net628));
 sg13g2_inv_1 _0339_ (.Y(_0042_),
    .A(net627));
 sg13g2_mux4_1 _0340_ (.S0(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit2.Q ),
    .A0(net53),
    .A1(net45),
    .A2(net64),
    .A3(net631),
    .S1(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit3.Q ),
    .X(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.S2BEG0 ));
 sg13g2_mux4_1 _0341_ (.S0(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame0_bit8.Q ),
    .A0(net235),
    .A1(net227),
    .A2(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.S2BEG0 ),
    .A3(net126),
    .S1(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame0_bit9.Q ),
    .X(_0043_));
 sg13g2_mux4_1 _0342_ (.S0(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame9_bit18.Q ),
    .A0(net161),
    .A1(net153),
    .A2(net171),
    .A3(net640),
    .S1(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame9_bit19.Q ),
    .X(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.N2BEGb0 ));
 sg13g2_mux4_1 _0343_ (.S0(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame0_bit9.Q ),
    .A0(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.N2BEGb0 ),
    .A1(net126),
    .A2(net235),
    .A3(net118),
    .S1(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame0_bit8.Q ),
    .X(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS2_BEG0 ));
 sg13g2_o21ai_1 _0344_ (.B1(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit29.Q ),
    .Y(_0044_),
    .A1(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit30.Q ),
    .A2(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.S2BEG0 ));
 sg13g2_nor2_1 _0345_ (.A(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit29.Q ),
    .B(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit30.Q ),
    .Y(_0045_));
 sg13g2_a22oi_1 _0346_ (.Y(_0046_),
    .B1(_0045_),
    .B2(net150),
    .A2(net129),
    .A1(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit30.Q ));
 sg13g2_nand3_1 _0347_ (.B(_0044_),
    .C(_0046_),
    .A(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit28.Q ),
    .Y(_0047_));
 sg13g2_nand2_1 _0348_ (.Y(_0048_),
    .A(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit30.Q ),
    .B(_0002_));
 sg13g2_o21ai_1 _0349_ (.B1(_0048_),
    .Y(_0049_),
    .A1(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit30.Q ),
    .A2(net149));
 sg13g2_nand3b_1 _0350_ (.B(net151),
    .C(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit29.Q ),
    .Y(_0050_),
    .A_N(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit30.Q ));
 sg13g2_o21ai_1 _0351_ (.B1(_0050_),
    .Y(_0051_),
    .A1(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit29.Q ),
    .A2(_0049_));
 sg13g2_o21ai_1 _0352_ (.B1(_0047_),
    .Y(_0052_),
    .A1(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit28.Q ),
    .A2(_0051_));
 sg13g2_mux4_1 _0353_ (.S0(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit28.Q ),
    .A0(net157),
    .A1(net160),
    .A2(net147),
    .A3(net148),
    .S1(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit29.Q ),
    .X(_0053_));
 sg13g2_mux4_1 _0354_ (.S0(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit28.Q ),
    .A0(net241),
    .A1(net229),
    .A2(net230),
    .A3(net154),
    .S1(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit29.Q ),
    .X(_0054_));
 sg13g2_mux2_1 _0355_ (.A0(_0054_),
    .A1(_0053_),
    .S(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit30.Q ),
    .X(_0055_));
 sg13g2_o21ai_1 _0356_ (.B1(net1),
    .Y(_0056_),
    .A1(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit31.Q ),
    .A2(_0055_));
 sg13g2_a21oi_1 _0357_ (.A1(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit31.Q ),
    .A2(_0052_),
    .Y(net326),
    .B1(_0056_));
 sg13g2_nand2b_1 _0358_ (.Y(_0057_),
    .B(net115),
    .A_N(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame0_bit26.Q ));
 sg13g2_nor3_1 _0359_ (.A(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame0_bit26.Q ),
    .B(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame0_bit27.Q ),
    .C(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.N1END1 ),
    .Y(_0058_));
 sg13g2_a221oi_1 _0360_ (.B2(_0057_),
    .C1(_0058_),
    .B1(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame0_bit27.Q ),
    .A1(_0003_),
    .Y(_0059_),
    .A2(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame0_bit26.Q ));
 sg13g2_mux4_1 _0361_ (.S0(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit28.Q ),
    .A0(net35),
    .A1(net65),
    .A2(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG13 ),
    .A3(_0059_),
    .S1(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit29.Q ),
    .X(_0060_));
 sg13g2_nand2b_1 _0362_ (.Y(_0061_),
    .B(_0060_),
    .A_N(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame0_bit26.Q ));
 sg13g2_nor3_1 _0363_ (.A(net224),
    .B(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame0_bit26.Q ),
    .C(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame0_bit27.Q ),
    .Y(_0062_));
 sg13g2_a221oi_1 _0364_ (.B2(_0061_),
    .C1(_0062_),
    .B1(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame0_bit27.Q ),
    .A1(_0009_),
    .Y(_0063_),
    .A2(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame0_bit26.Q ));
 sg13g2_mux4_1 _0365_ (.S0(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame9_bit13.Q ),
    .A0(net143),
    .A1(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.J_NS4_BEG13 ),
    .A2(net169),
    .A3(_0063_),
    .S1(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame9_bit12.Q ),
    .X(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.N1END1 ));
 sg13g2_mux4_1 _0366_ (.S0(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame0_bit2.Q ),
    .A0(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.N1END1 ),
    .A1(net248),
    .A2(net115),
    .A3(net135),
    .S1(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame0_bit3.Q ),
    .X(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG13 ));
 sg13g2_mux4_1 _0367_ (.S0(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame9_bit24.Q ),
    .A0(net35),
    .A1(net61),
    .A2(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG13 ),
    .A3(_0059_),
    .S1(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame9_bit25.Q ),
    .X(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.N1BEG1 ));
 sg13g2_nand2b_1 _0368_ (.Y(_0064_),
    .B(net116),
    .A_N(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame0_bit28.Q ));
 sg13g2_nor3_1 _0369_ (.A(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame0_bit28.Q ),
    .B(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame0_bit29.Q ),
    .C(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.N1END2 ),
    .Y(_0065_));
 sg13g2_a221oi_1 _0370_ (.B2(_0064_),
    .C1(_0065_),
    .B1(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame0_bit29.Q ),
    .A1(_0004_),
    .Y(_0066_),
    .A2(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame0_bit28.Q ));
 sg13g2_mux4_1 _0371_ (.S0(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit30.Q ),
    .A0(net36),
    .A1(net55),
    .A2(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG14 ),
    .A3(_0066_),
    .S1(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit31.Q ),
    .X(_0067_));
 sg13g2_nor3_1 _0372_ (.A(net225),
    .B(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame0_bit28.Q ),
    .C(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame0_bit29.Q ),
    .Y(_0068_));
 sg13g2_nand2b_1 _0373_ (.Y(_0069_),
    .B(_0067_),
    .A_N(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame0_bit28.Q ));
 sg13g2_a221oi_1 _0374_ (.B2(_0069_),
    .C1(_0068_),
    .B1(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame0_bit29.Q ),
    .A1(_0008_),
    .Y(_0070_),
    .A2(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame0_bit28.Q ));
 sg13g2_mux4_1 _0375_ (.S0(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame9_bit15.Q ),
    .A0(net144),
    .A1(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.J_NS4_BEG14 ),
    .A2(net170),
    .A3(_0070_),
    .S1(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame9_bit14.Q ),
    .X(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.N1END2 ));
 sg13g2_mux4_1 _0376_ (.S0(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame0_bit4.Q ),
    .A0(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.N1END2 ),
    .A1(net249),
    .A2(net116),
    .A3(net136),
    .S1(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame0_bit5.Q ),
    .X(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG14 ));
 sg13g2_mux4_1 _0377_ (.S0(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame9_bit26.Q ),
    .A0(net36),
    .A1(net62),
    .A2(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG14 ),
    .A3(_0066_),
    .S1(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame9_bit27.Q ),
    .X(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.N1BEG2 ));
 sg13g2_nand2b_1 _0378_ (.Y(_0071_),
    .B(net117),
    .A_N(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame0_bit30.Q ));
 sg13g2_nor3_1 _0379_ (.A(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame0_bit30.Q ),
    .B(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame0_bit31.Q ),
    .C(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.N1END3 ),
    .Y(_0072_));
 sg13g2_a221oi_1 _0380_ (.B2(_0071_),
    .C1(_0072_),
    .B1(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame0_bit31.Q ),
    .A1(_0005_),
    .Y(_0073_),
    .A2(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame0_bit30.Q ));
 sg13g2_mux4_1 _0381_ (.S0(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit0.Q ),
    .A0(net37),
    .A1(net56),
    .A2(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG15 ),
    .A3(_0073_),
    .S1(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit1.Q ),
    .X(_0074_));
 sg13g2_nor3_1 _0382_ (.A(net226),
    .B(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame0_bit30.Q ),
    .C(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame0_bit31.Q ),
    .Y(_0075_));
 sg13g2_nand2b_1 _0383_ (.Y(_0076_),
    .B(_0074_),
    .A_N(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame0_bit30.Q ));
 sg13g2_a221oi_1 _0384_ (.B2(_0076_),
    .C1(_0075_),
    .B1(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame0_bit31.Q ),
    .A1(_0007_),
    .Y(_0077_),
    .A2(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame0_bit30.Q ));
 sg13g2_mux4_1 _0385_ (.S0(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame9_bit17.Q ),
    .A0(net145),
    .A1(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.J_NS4_BEG15 ),
    .A2(net171),
    .A3(_0077_),
    .S1(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame9_bit16.Q ),
    .X(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.N1END3 ));
 sg13g2_mux4_1 _0386_ (.S0(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame0_bit6.Q ),
    .A0(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.N1END3 ),
    .A1(net250),
    .A2(net117),
    .A3(net137),
    .S1(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame0_bit7.Q ),
    .X(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG15 ));
 sg13g2_mux4_1 _0387_ (.S0(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame9_bit28.Q ),
    .A0(net37),
    .A1(net63),
    .A2(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG15 ),
    .A3(_0073_),
    .S1(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame9_bit29.Q ),
    .X(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.N1BEG3 ));
 sg13g2_mux4_1 _0388_ (.S0(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame9_bit30.Q ),
    .A0(net53),
    .A1(net45),
    .A2(net63),
    .A3(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS2_BEG0 ),
    .S1(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame9_bit31.Q ),
    .X(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.N2BEG0 ));
 sg13g2_mux4_1 _0389_ (.S0(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit4.Q ),
    .A0(net52),
    .A1(net44),
    .A2(net65),
    .A3(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS2_BEG1 ),
    .S1(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit5.Q ),
    .X(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.S2BEG1 ));
 sg13g2_mux4_1 _0390_ (.S0(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame0_bit10.Q ),
    .A0(net236),
    .A1(net228),
    .A2(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.S2BEG1 ),
    .A3(net127),
    .S1(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame0_bit11.Q ),
    .X(_0078_));
 sg13g2_mux4_1 _0391_ (.S0(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame9_bit20.Q ),
    .A0(net160),
    .A1(net152),
    .A2(net170),
    .A3(_0078_),
    .S1(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame9_bit21.Q ),
    .X(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.N2BEGb1 ));
 sg13g2_mux4_1 _0392_ (.S0(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame0_bit11.Q ),
    .A0(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.N2BEGb1 ),
    .A1(net127),
    .A2(net236),
    .A3(net119),
    .S1(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame0_bit10.Q ),
    .X(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS2_BEG1 ));
 sg13g2_mux4_1 _0393_ (.S0(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit0.Q ),
    .A0(net52),
    .A1(net44),
    .A2(net62),
    .A3(net630),
    .S1(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit1.Q ),
    .X(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.N2BEG1 ));
 sg13g2_mux4_1 _0394_ (.S0(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit6.Q ),
    .A0(net51),
    .A1(net43),
    .A2(net55),
    .A3(net629),
    .S1(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit7.Q ),
    .X(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.S2BEG2 ));
 sg13g2_mux4_1 _0395_ (.S0(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame0_bit13.Q ),
    .A0(net237),
    .A1(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.S2BEG2 ),
    .A2(net229),
    .A3(net128),
    .S1(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame0_bit12.Q ),
    .X(_0079_));
 sg13g2_mux4_1 _0396_ (.S0(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame9_bit23.Q ),
    .A0(net159),
    .A1(net169),
    .A2(net151),
    .A3(_0079_),
    .S1(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame9_bit22.Q ),
    .X(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.N2BEGb2 ));
 sg13g2_mux4_1 _0397_ (.S0(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame0_bit12.Q ),
    .A0(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.N2BEGb2 ),
    .A1(net237),
    .A2(net128),
    .A3(net120),
    .S1(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame0_bit13.Q ),
    .X(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS2_BEG2 ));
 sg13g2_mux4_1 _0398_ (.S0(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit2.Q ),
    .A0(net51),
    .A1(net43),
    .A2(net61),
    .A3(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS2_BEG2 ),
    .S1(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit3.Q ),
    .X(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.N2BEG2 ));
 sg13g2_mux4_1 _0399_ (.S0(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit8.Q ),
    .A0(net50),
    .A1(net42),
    .A2(net56),
    .A3(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS2_BEG3 ),
    .S1(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit9.Q ),
    .X(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.S2BEG3 ));
 sg13g2_mux4_1 _0400_ (.S0(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame0_bit15.Q ),
    .A0(net238),
    .A1(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.S2BEG3 ),
    .A2(net230),
    .A3(net129),
    .S1(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame0_bit14.Q ),
    .X(_0080_));
 sg13g2_mux4_1 _0401_ (.S0(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame9_bit25.Q ),
    .A0(net158),
    .A1(net168),
    .A2(net150),
    .A3(_0080_),
    .S1(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame9_bit24.Q ),
    .X(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.N2BEGb3 ));
 sg13g2_mux4_1 _0402_ (.S0(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame0_bit14.Q ),
    .A0(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.N2BEGb3 ),
    .A1(net238),
    .A2(net129),
    .A3(net121),
    .S1(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame0_bit15.Q ),
    .X(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS2_BEG3 ));
 sg13g2_mux4_1 _0403_ (.S0(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit4.Q ),
    .A0(net50),
    .A1(net42),
    .A2(net60),
    .A3(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS2_BEG3 ),
    .S1(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit5.Q ),
    .X(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.N2BEG3 ));
 sg13g2_mux4_1 _0404_ (.S0(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit11.Q ),
    .A0(net34),
    .A1(net41),
    .A2(net49),
    .A3(net626),
    .S1(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit10.Q ),
    .X(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.S2BEG4 ));
 sg13g2_mux4_1 _0405_ (.S0(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame0_bit16.Q ),
    .A0(net239),
    .A1(net231),
    .A2(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.S2BEG4 ),
    .A3(net130),
    .S1(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame0_bit17.Q ),
    .X(_0081_));
 sg13g2_mux4_1 _0406_ (.S0(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame9_bit26.Q ),
    .A0(net157),
    .A1(net149),
    .A2(net167),
    .A3(net636),
    .S1(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame9_bit27.Q ),
    .X(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.N2BEGb4 ));
 sg13g2_mux4_1 _0407_ (.S0(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame0_bit17.Q ),
    .A0(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.N2BEGb4 ),
    .A1(net130),
    .A2(net239),
    .A3(net122),
    .S1(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame0_bit16.Q ),
    .X(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS2_BEG4 ));
 sg13g2_mux4_1 _0408_ (.S0(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit6.Q ),
    .A0(net49),
    .A1(net41),
    .A2(net59),
    .A3(net627),
    .S1(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit7.Q ),
    .X(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.N2BEG4 ));
 sg13g2_mux4_1 _0409_ (.S0(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit12.Q ),
    .A0(net35),
    .A1(net48),
    .A2(net40),
    .A3(net625),
    .S1(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit13.Q ),
    .X(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.S2BEG5 ));
 sg13g2_mux4_1 _0410_ (.S0(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame0_bit18.Q ),
    .A0(net240),
    .A1(net232),
    .A2(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.S2BEG5 ),
    .A3(net131),
    .S1(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame0_bit19.Q ),
    .X(_0082_));
 sg13g2_mux4_1 _0411_ (.S0(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame9_bit29.Q ),
    .A0(net156),
    .A1(net166),
    .A2(net148),
    .A3(_0082_),
    .S1(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame9_bit28.Q ),
    .X(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.N2BEGb5 ));
 sg13g2_mux4_1 _0412_ (.S0(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame0_bit19.Q ),
    .A0(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.N2BEGb5 ),
    .A1(net131),
    .A2(net240),
    .A3(net123),
    .S1(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame0_bit18.Q ),
    .X(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS2_BEG5 ));
 sg13g2_mux4_1 _0413_ (.S0(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit8.Q ),
    .A0(net48),
    .A1(net40),
    .A2(net58),
    .A3(net625),
    .S1(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit9.Q ),
    .X(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.N2BEG5 ));
 sg13g2_mux4_1 _0414_ (.S0(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit14.Q ),
    .A0(net36),
    .A1(net47),
    .A2(net39),
    .A3(net624),
    .S1(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit15.Q ),
    .X(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.S2BEG6 ));
 sg13g2_mux4_1 _0415_ (.S0(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame0_bit20.Q ),
    .A0(net241),
    .A1(net233),
    .A2(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.S2BEG6 ),
    .A3(net132),
    .S1(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame0_bit21.Q ),
    .X(_0083_));
 sg13g2_mux4_1 _0416_ (.S0(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame9_bit31.Q ),
    .A0(net155),
    .A1(net165),
    .A2(net147),
    .A3(_0083_),
    .S1(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame9_bit30.Q ),
    .X(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.N2BEGb6 ));
 sg13g2_mux4_1 _0417_ (.S0(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame0_bit21.Q ),
    .A0(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.N2BEGb6 ),
    .A1(net132),
    .A2(net241),
    .A3(net124),
    .S1(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame0_bit20.Q ),
    .X(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS2_BEG6 ));
 sg13g2_mux4_1 _0418_ (.S0(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit10.Q ),
    .A0(net47),
    .A1(net39),
    .A2(net57),
    .A3(net624),
    .S1(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit11.Q ),
    .X(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.N2BEG6 ));
 sg13g2_mux4_1 _0419_ (.S0(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit16.Q ),
    .A0(net37),
    .A1(net46),
    .A2(net38),
    .A3(net623),
    .S1(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit17.Q ),
    .X(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.S2BEG7 ));
 sg13g2_mux4_1 _0420_ (.S0(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame0_bit22.Q ),
    .A0(net242),
    .A1(net234),
    .A2(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.S2BEG7 ),
    .A3(net133),
    .S1(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame0_bit23.Q ),
    .X(_0084_));
 sg13g2_mux4_1 _0421_ (.S0(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit0.Q ),
    .A0(net154),
    .A1(net146),
    .A2(net162),
    .A3(_0084_),
    .S1(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit1.Q ),
    .X(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.N2BEGb7 ));
 sg13g2_mux4_1 _0422_ (.S0(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame0_bit23.Q ),
    .A0(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.N2BEGb7 ),
    .A1(net133),
    .A2(net242),
    .A3(net125),
    .S1(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame0_bit22.Q ),
    .X(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS2_BEG7 ));
 sg13g2_mux4_1 _0423_ (.S0(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit12.Q ),
    .A0(net46),
    .A1(net38),
    .A2(net54),
    .A3(net623),
    .S1(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit13.Q ),
    .X(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.N2BEG7 ));
 sg13g2_nand2b_1 _0424_ (.Y(_0085_),
    .B(net114),
    .A_N(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame0_bit24.Q ));
 sg13g2_nor3_1 _0425_ (.A(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame0_bit24.Q ),
    .B(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame0_bit25.Q ),
    .C(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.N1END0 ),
    .Y(_0086_));
 sg13g2_a221oi_1 _0426_ (.B2(_0085_),
    .C1(_0086_),
    .B1(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame0_bit25.Q ),
    .A1(_0006_),
    .Y(_0087_),
    .A2(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame0_bit24.Q ));
 sg13g2_mux4_1 _0427_ (.S0(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit27.Q ),
    .A0(net34),
    .A1(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG12 ),
    .A2(net64),
    .A3(_0087_),
    .S1(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit26.Q ),
    .X(_0088_));
 sg13g2_nor3_1 _0428_ (.A(net223),
    .B(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame0_bit24.Q ),
    .C(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame0_bit25.Q ),
    .Y(_0089_));
 sg13g2_nand2b_1 _0429_ (.Y(_0090_),
    .B(_0088_),
    .A_N(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame0_bit24.Q ));
 sg13g2_a221oi_1 _0430_ (.B2(_0090_),
    .C1(_0089_),
    .B1(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame0_bit25.Q ),
    .A1(_0010_),
    .Y(_0091_),
    .A2(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame0_bit24.Q ));
 sg13g2_mux4_1 _0431_ (.S0(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame9_bit11.Q ),
    .A0(net142),
    .A1(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.J_NS4_BEG12 ),
    .A2(net168),
    .A3(_0091_),
    .S1(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame9_bit10.Q ),
    .X(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.N1END0 ));
 sg13g2_mux4_1 _0432_ (.S0(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit31.Q ),
    .A0(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.N1END0 ),
    .A1(net12),
    .A2(net114),
    .A3(net18),
    .S1(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit30.Q ),
    .X(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.W1BEG0 ));
 sg13g2_mux4_1 _0433_ (.S0(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame6_bit1.Q ),
    .A0(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.N1END1 ),
    .A1(net13),
    .A2(net115),
    .A3(net17),
    .S1(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame6_bit0.Q ),
    .X(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.W1BEG1 ));
 sg13g2_mux4_1 _0434_ (.S0(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame6_bit3.Q ),
    .A0(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.N1END2 ),
    .A1(net10),
    .A2(net116),
    .A3(net16),
    .S1(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame6_bit2.Q ),
    .X(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.W1BEG2 ));
 sg13g2_mux4_1 _0435_ (.S0(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame6_bit5.Q ),
    .A0(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.N1END3 ),
    .A1(net11),
    .A2(net117),
    .A3(net15),
    .S1(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame6_bit4.Q ),
    .X(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.W1BEG3 ));
 sg13g2_mux4_1 _0436_ (.S0(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame6_bit6.Q ),
    .A0(net10),
    .A1(net19),
    .A2(net631),
    .A3(net623),
    .S1(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame6_bit7.Q ),
    .X(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.W2BEG0 ));
 sg13g2_mux4_1 _0437_ (.S0(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame6_bit8.Q ),
    .A0(net11),
    .A1(net20),
    .A2(net630),
    .A3(net624),
    .S1(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame6_bit9.Q ),
    .X(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.W2BEG1 ));
 sg13g2_mux4_1 _0438_ (.S0(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame6_bit10.Q ),
    .A0(net12),
    .A1(net21),
    .A2(net629),
    .A3(net625),
    .S1(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame6_bit11.Q ),
    .X(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.W2BEG2 ));
 sg13g2_mux4_1 _0439_ (.S0(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame6_bit12.Q ),
    .A0(net13),
    .A1(net22),
    .A2(net628),
    .A3(net626),
    .S1(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame6_bit13.Q ),
    .X(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.W2BEG3 ));
 sg13g2_mux4_1 _0440_ (.S0(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame6_bit14.Q ),
    .A0(net15),
    .A1(net23),
    .A2(net628),
    .A3(net627),
    .S1(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame6_bit15.Q ),
    .X(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.W2BEG4 ));
 sg13g2_mux4_1 _0441_ (.S0(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame6_bit16.Q ),
    .A0(net16),
    .A1(net24),
    .A2(net629),
    .A3(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS2_BEG5 ),
    .S1(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame6_bit17.Q ),
    .X(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.W2BEG5 ));
 sg13g2_mux4_1 _0442_ (.S0(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame6_bit18.Q ),
    .A0(net17),
    .A1(net26),
    .A2(net630),
    .A3(net624),
    .S1(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame6_bit19.Q ),
    .X(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.W2BEG6 ));
 sg13g2_mux4_1 _0443_ (.S0(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame6_bit20.Q ),
    .A0(net18),
    .A1(net27),
    .A2(net631),
    .A3(net623),
    .S1(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame6_bit21.Q ),
    .X(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.W2BEG7 ));
 sg13g2_mux4_1 _0444_ (.S0(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame6_bit22.Q ),
    .A0(net10),
    .A1(net19),
    .A2(net631),
    .A3(net623),
    .S1(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame6_bit23.Q ),
    .X(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.W2BEGb0 ));
 sg13g2_mux4_1 _0445_ (.S0(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame6_bit24.Q ),
    .A0(net11),
    .A1(net20),
    .A2(net630),
    .A3(net624),
    .S1(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame6_bit25.Q ),
    .X(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.W2BEGb1 ));
 sg13g2_mux4_1 _0446_ (.S0(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame6_bit26.Q ),
    .A0(net12),
    .A1(net21),
    .A2(net629),
    .A3(net625),
    .S1(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame6_bit27.Q ),
    .X(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.W2BEGb2 ));
 sg13g2_mux4_1 _0447_ (.S0(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame6_bit28.Q ),
    .A0(net13),
    .A1(net22),
    .A2(net628),
    .A3(net626),
    .S1(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame6_bit29.Q ),
    .X(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.W2BEGb3 ));
 sg13g2_mux4_1 _0448_ (.S0(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame6_bit30.Q ),
    .A0(net15),
    .A1(net23),
    .A2(net628),
    .A3(net626),
    .S1(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame6_bit31.Q ),
    .X(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.W2BEGb4 ));
 sg13g2_mux4_1 _0449_ (.S0(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame5_bit0.Q ),
    .A0(net16),
    .A1(net24),
    .A2(net629),
    .A3(net625),
    .S1(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame5_bit1.Q ),
    .X(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.W2BEGb5 ));
 sg13g2_mux4_1 _0450_ (.S0(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame5_bit2.Q ),
    .A0(net17),
    .A1(net26),
    .A2(net630),
    .A3(net624),
    .S1(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame5_bit3.Q ),
    .X(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.W2BEGb6 ));
 sg13g2_mux4_1 _0451_ (.S0(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame5_bit4.Q ),
    .A0(net18),
    .A1(net27),
    .A2(net631),
    .A3(net623),
    .S1(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame5_bit5.Q ),
    .X(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.W2BEGb7 ));
 sg13g2_mux4_1 _0452_ (.S0(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame5_bit6.Q ),
    .A0(net10),
    .A1(net23),
    .A2(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG15 ),
    .A3(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS2_BEG7 ),
    .S1(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame5_bit7.Q ),
    .X(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.WW4BEG0 ));
 sg13g2_mux4_1 _0453_ (.S0(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame5_bit8.Q ),
    .A0(net11),
    .A1(net24),
    .A2(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG14 ),
    .A3(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS2_BEG6 ),
    .S1(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame5_bit9.Q ),
    .X(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.WW4BEG1 ));
 sg13g2_mux4_1 _0454_ (.S0(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame5_bit10.Q ),
    .A0(net12),
    .A1(net26),
    .A2(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG13 ),
    .A3(net625),
    .S1(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame5_bit11.Q ),
    .X(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.WW4BEG2 ));
 sg13g2_mux4_1 _0455_ (.S0(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame0_bit0.Q ),
    .A0(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.N1END0 ),
    .A1(net247),
    .A2(net114),
    .A3(net134),
    .S1(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame0_bit1.Q ),
    .X(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG12 ));
 sg13g2_mux4_1 _0456_ (.S0(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame5_bit12.Q ),
    .A0(net13),
    .A1(net27),
    .A2(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG12 ),
    .A3(net626),
    .S1(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame5_bit13.Q ),
    .X(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.WW4BEG3 ));
 sg13g2_mux4_1 _0457_ (.S0(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame1_bit30.Q ),
    .A0(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.N1END3 ),
    .A1(net250),
    .A2(net117),
    .A3(net137),
    .S1(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame1_bit31.Q ),
    .X(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG11 ));
 sg13g2_mux4_1 _0458_ (.S0(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame5_bit14.Q ),
    .A0(net15),
    .A1(net19),
    .A2(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG11 ),
    .A3(net628),
    .S1(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame5_bit15.Q ),
    .X(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.WW4BEG4 ));
 sg13g2_mux4_1 _0459_ (.S0(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame1_bit28.Q ),
    .A0(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.N1END2 ),
    .A1(net249),
    .A2(net116),
    .A3(net136),
    .S1(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame1_bit29.Q ),
    .X(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG10 ));
 sg13g2_mux4_1 _0460_ (.S0(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame5_bit16.Q ),
    .A0(net16),
    .A1(net19),
    .A2(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG10 ),
    .A3(net629),
    .S1(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame5_bit17.Q ),
    .X(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.WW4BEG5 ));
 sg13g2_mux4_1 _0461_ (.S0(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame1_bit26.Q ),
    .A0(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.N1END1 ),
    .A1(net248),
    .A2(net115),
    .A3(net135),
    .S1(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame1_bit27.Q ),
    .X(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG9 ));
 sg13g2_mux4_1 _0462_ (.S0(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame5_bit18.Q ),
    .A0(net17),
    .A1(net21),
    .A2(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG9 ),
    .A3(net630),
    .S1(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame5_bit19.Q ),
    .X(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.WW4BEG6 ));
 sg13g2_mux4_1 _0463_ (.S0(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame1_bit24.Q ),
    .A0(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.N1END0 ),
    .A1(net247),
    .A2(net114),
    .A3(net134),
    .S1(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame1_bit25.Q ),
    .X(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG8 ));
 sg13g2_mux4_1 _0464_ (.S0(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame5_bit20.Q ),
    .A0(net18),
    .A1(net22),
    .A2(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG8 ),
    .A3(net631),
    .S1(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame5_bit21.Q ),
    .X(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.WW4BEG7 ));
 sg13g2_mux4_1 _0465_ (.S0(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame1_bit22.Q ),
    .A0(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.N1END3 ),
    .A1(net250),
    .A2(net117),
    .A3(net137),
    .S1(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame1_bit23.Q ),
    .X(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG7 ));
 sg13g2_mux4_1 _0466_ (.S0(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame5_bit22.Q ),
    .A0(net15),
    .A1(net19),
    .A2(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG7 ),
    .A3(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS2_BEG7 ),
    .S1(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame5_bit23.Q ),
    .X(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.WW4BEG8 ));
 sg13g2_mux4_1 _0467_ (.S0(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame1_bit20.Q ),
    .A0(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.N1END2 ),
    .A1(net249),
    .A2(net116),
    .A3(net136),
    .S1(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame1_bit21.Q ),
    .X(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG6 ));
 sg13g2_mux4_1 _0468_ (.S0(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame5_bit24.Q ),
    .A0(net16),
    .A1(net20),
    .A2(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG6 ),
    .A3(net624),
    .S1(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame5_bit25.Q ),
    .X(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.WW4BEG9 ));
 sg13g2_mux4_1 _0469_ (.S0(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame1_bit18.Q ),
    .A0(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.N1END1 ),
    .A1(net248),
    .A2(net115),
    .A3(net135),
    .S1(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame1_bit19.Q ),
    .X(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG5 ));
 sg13g2_mux4_1 _0470_ (.S0(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame5_bit26.Q ),
    .A0(net17),
    .A1(net21),
    .A2(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG5 ),
    .A3(net625),
    .S1(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame5_bit27.Q ),
    .X(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.WW4BEG10 ));
 sg13g2_mux4_1 _0471_ (.S0(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame1_bit16.Q ),
    .A0(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.N1END0 ),
    .A1(net247),
    .A2(net114),
    .A3(net134),
    .S1(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame1_bit17.Q ),
    .X(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG4 ));
 sg13g2_mux4_1 _0472_ (.S0(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame5_bit28.Q ),
    .A0(net18),
    .A1(net22),
    .A2(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG4 ),
    .A3(net626),
    .S1(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame5_bit29.Q ),
    .X(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.WW4BEG11 ));
 sg13g2_mux4_1 _0473_ (.S0(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame1_bit14.Q ),
    .A0(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.N1END3 ),
    .A1(net250),
    .A2(net117),
    .A3(net137),
    .S1(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame1_bit15.Q ),
    .X(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG3 ));
 sg13g2_mux4_1 _0474_ (.S0(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame5_bit30.Q ),
    .A0(net10),
    .A1(net23),
    .A2(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG3 ),
    .A3(net628),
    .S1(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame5_bit31.Q ),
    .X(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.WW4BEG12 ));
 sg13g2_mux4_1 _0475_ (.S0(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame1_bit12.Q ),
    .A0(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.N1END2 ),
    .A1(net249),
    .A2(net116),
    .A3(net136),
    .S1(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame1_bit13.Q ),
    .X(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG2 ));
 sg13g2_mux4_1 _0476_ (.S0(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame4_bit0.Q ),
    .A0(net11),
    .A1(net24),
    .A2(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG2 ),
    .A3(net629),
    .S1(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame4_bit1.Q ),
    .X(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.WW4BEG13 ));
 sg13g2_mux4_1 _0477_ (.S0(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame1_bit10.Q ),
    .A0(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.N1END1 ),
    .A1(net248),
    .A2(net115),
    .A3(net135),
    .S1(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame1_bit11.Q ),
    .X(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG1 ));
 sg13g2_mux4_1 _0478_ (.S0(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame4_bit2.Q ),
    .A0(net12),
    .A1(net26),
    .A2(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG1 ),
    .A3(net630),
    .S1(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame4_bit3.Q ),
    .X(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.WW4BEG14 ));
 sg13g2_mux4_1 _0479_ (.S0(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame1_bit8.Q ),
    .A0(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.N1END0 ),
    .A1(net247),
    .A2(net114),
    .A3(net134),
    .S1(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame1_bit9.Q ),
    .X(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG0 ));
 sg13g2_mux4_1 _0480_ (.S0(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame4_bit4.Q ),
    .A0(net13),
    .A1(net27),
    .A2(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG0 ),
    .A3(net631),
    .S1(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame4_bit5.Q ),
    .X(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.WW4BEG15 ));
 sg13g2_mux4_1 _0481_ (.S0(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame4_bit6.Q ),
    .A0(net247),
    .A1(net134),
    .A2(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG11 ),
    .A3(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG15 ),
    .S1(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame4_bit7.Q ),
    .X(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.W6BEG0 ));
 sg13g2_mux4_1 _0482_ (.S0(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame4_bit8.Q ),
    .A0(net248),
    .A1(net135),
    .A2(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG10 ),
    .A3(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG14 ),
    .S1(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame4_bit9.Q ),
    .X(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.W6BEG1 ));
 sg13g2_mux4_1 _0483_ (.S0(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame4_bit10.Q ),
    .A0(net249),
    .A1(net136),
    .A2(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG9 ),
    .A3(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG13 ),
    .S1(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame4_bit11.Q ),
    .X(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.W6BEG2 ));
 sg13g2_mux4_1 _0484_ (.S0(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame4_bit12.Q ),
    .A0(net250),
    .A1(net137),
    .A2(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG8 ),
    .A3(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG12 ),
    .S1(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame4_bit13.Q ),
    .X(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.W6BEG3 ));
 sg13g2_mux4_1 _0485_ (.S0(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame4_bit15.Q ),
    .A0(net15),
    .A1(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG11 ),
    .A2(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG7 ),
    .A3(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS2_BEG0 ),
    .S1(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame4_bit14.Q ),
    .X(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.W6BEG4 ));
 sg13g2_mux4_1 _0486_ (.S0(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame4_bit17.Q ),
    .A0(net16),
    .A1(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG10 ),
    .A2(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG6 ),
    .A3(net630),
    .S1(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame4_bit16.Q ),
    .X(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.W6BEG5 ));
 sg13g2_mux4_1 _0487_ (.S0(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame4_bit18.Q ),
    .A0(net17),
    .A1(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG5 ),
    .A2(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG9 ),
    .A3(net629),
    .S1(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame4_bit19.Q ),
    .X(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.W6BEG6 ));
 sg13g2_mux4_1 _0488_ (.S0(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame4_bit20.Q ),
    .A0(net18),
    .A1(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG4 ),
    .A2(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG8 ),
    .A3(net628),
    .S1(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame4_bit21.Q ),
    .X(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.W6BEG7 ));
 sg13g2_mux4_1 _0489_ (.S0(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame4_bit23.Q ),
    .A0(net10),
    .A1(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG7 ),
    .A2(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG3 ),
    .A3(net626),
    .S1(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame4_bit22.Q ),
    .X(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.W6BEG8 ));
 sg13g2_mux4_1 _0490_ (.S0(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame4_bit25.Q ),
    .A0(net11),
    .A1(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG6 ),
    .A2(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG2 ),
    .A3(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS2_BEG5 ),
    .S1(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame4_bit24.Q ),
    .X(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.W6BEG9 ));
 sg13g2_mux4_1 _0491_ (.S0(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame4_bit27.Q ),
    .A0(net12),
    .A1(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG5 ),
    .A2(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG1 ),
    .A3(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS2_BEG6 ),
    .S1(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame4_bit26.Q ),
    .X(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.W6BEG10 ));
 sg13g2_mux4_1 _0492_ (.S0(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame4_bit29.Q ),
    .A0(net13),
    .A1(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG4 ),
    .A2(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG0 ),
    .A3(net623),
    .S1(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame4_bit28.Q ),
    .X(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.W6BEG11 ));
 sg13g2_mux4_1 _0493_ (.S0(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame4_bit30.Q ),
    .A0(net66),
    .A1(net80),
    .A2(net54),
    .A3(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG0 ),
    .S1(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame4_bit31.Q ),
    .X(net302));
 sg13g2_mux4_1 _0494_ (.S0(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame3_bit0.Q ),
    .A0(net73),
    .A1(net81),
    .A2(net57),
    .A3(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG1 ),
    .S1(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame3_bit1.Q ),
    .X(net303));
 sg13g2_mux4_1 _0495_ (.S0(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame3_bit2.Q ),
    .A0(net74),
    .A1(net67),
    .A2(net58),
    .A3(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG2 ),
    .S1(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame3_bit3.Q ),
    .X(net304));
 sg13g2_mux4_1 _0496_ (.S0(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame3_bit4.Q ),
    .A0(net75),
    .A1(net68),
    .A2(net59),
    .A3(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG3 ),
    .S1(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame3_bit5.Q ),
    .X(net305));
 sg13g2_mux4_1 _0497_ (.S0(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame3_bit6.Q ),
    .A0(net76),
    .A1(net69),
    .A2(net60),
    .A3(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG4 ),
    .S1(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame3_bit7.Q ),
    .X(net307));
 sg13g2_mux4_1 _0498_ (.S0(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame3_bit8.Q ),
    .A0(net77),
    .A1(net70),
    .A2(net61),
    .A3(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG5 ),
    .S1(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame3_bit9.Q ),
    .X(net308));
 sg13g2_mux4_1 _0499_ (.S0(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame3_bit10.Q ),
    .A0(net78),
    .A1(net71),
    .A2(net62),
    .A3(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG6 ),
    .S1(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame3_bit11.Q ),
    .X(net309));
 sg13g2_mux4_1 _0500_ (.S0(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame3_bit12.Q ),
    .A0(net79),
    .A1(net72),
    .A2(net63),
    .A3(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG7 ),
    .S1(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame3_bit13.Q ),
    .X(net310));
 sg13g2_mux4_1 _0501_ (.S0(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame3_bit14.Q ),
    .A0(net66),
    .A1(net80),
    .A2(net64),
    .A3(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG8 ),
    .S1(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame3_bit15.Q ),
    .X(net311));
 sg13g2_mux4_1 _0502_ (.S0(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame3_bit16.Q ),
    .A0(net73),
    .A1(net81),
    .A2(net65),
    .A3(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG9 ),
    .S1(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame3_bit17.Q ),
    .X(net312));
 sg13g2_mux4_1 _0503_ (.S0(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame3_bit18.Q ),
    .A0(net74),
    .A1(net67),
    .A2(net55),
    .A3(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG10 ),
    .S1(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame3_bit19.Q ),
    .X(net313));
 sg13g2_mux4_1 _0504_ (.S0(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame3_bit20.Q ),
    .A0(net75),
    .A1(net68),
    .A2(net56),
    .A3(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG11 ),
    .S1(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame3_bit21.Q ),
    .X(net314));
 sg13g2_mux4_1 _0505_ (.S0(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame3_bit22.Q ),
    .A0(net34),
    .A1(net76),
    .A2(net69),
    .A3(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG12 ),
    .S1(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame3_bit23.Q ),
    .X(net315));
 sg13g2_mux4_1 _0506_ (.S0(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame3_bit24.Q ),
    .A0(net35),
    .A1(net77),
    .A2(net70),
    .A3(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG13 ),
    .S1(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame3_bit25.Q ),
    .X(net316));
 sg13g2_mux4_1 _0507_ (.S0(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame3_bit26.Q ),
    .A0(net36),
    .A1(net78),
    .A2(net71),
    .A3(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG14 ),
    .S1(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame3_bit27.Q ),
    .X(net318));
 sg13g2_mux4_1 _0508_ (.S0(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame3_bit28.Q ),
    .A0(net37),
    .A1(net79),
    .A2(net72),
    .A3(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG15 ),
    .S1(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame3_bit29.Q ),
    .X(net319));
 sg13g2_mux4_1 _0509_ (.S0(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame3_bit30.Q ),
    .A0(net66),
    .A1(net80),
    .A2(net54),
    .A3(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG0 ),
    .S1(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame3_bit31.Q ),
    .X(net269));
 sg13g2_mux4_1 _0510_ (.S0(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame2_bit0.Q ),
    .A0(net73),
    .A1(net81),
    .A2(net57),
    .A3(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG1 ),
    .S1(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame2_bit1.Q ),
    .X(net270));
 sg13g2_mux4_1 _0511_ (.S0(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame2_bit2.Q ),
    .A0(net74),
    .A1(net67),
    .A2(net58),
    .A3(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG2 ),
    .S1(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame2_bit3.Q ),
    .X(net271));
 sg13g2_mux4_1 _0512_ (.S0(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame2_bit4.Q ),
    .A0(net75),
    .A1(net68),
    .A2(net59),
    .A3(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG3 ),
    .S1(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame2_bit5.Q ),
    .X(net272));
 sg13g2_mux4_1 _0513_ (.S0(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame2_bit6.Q ),
    .A0(net76),
    .A1(net69),
    .A2(net60),
    .A3(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG4 ),
    .S1(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame2_bit7.Q ),
    .X(net274));
 sg13g2_mux4_1 _0514_ (.S0(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame2_bit8.Q ),
    .A0(net77),
    .A1(net70),
    .A2(net61),
    .A3(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG5 ),
    .S1(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame2_bit9.Q ),
    .X(net275));
 sg13g2_mux4_1 _0515_ (.S0(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame2_bit10.Q ),
    .A0(net78),
    .A1(net71),
    .A2(net62),
    .A3(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG6 ),
    .S1(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame2_bit11.Q ),
    .X(net276));
 sg13g2_mux4_1 _0516_ (.S0(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame2_bit12.Q ),
    .A0(net79),
    .A1(net72),
    .A2(net63),
    .A3(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG7 ),
    .S1(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame2_bit13.Q ),
    .X(net277));
 sg13g2_mux4_1 _0517_ (.S0(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame2_bit14.Q ),
    .A0(net66),
    .A1(net80),
    .A2(net64),
    .A3(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG8 ),
    .S1(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame2_bit15.Q ),
    .X(net278));
 sg13g2_mux4_1 _0518_ (.S0(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame2_bit16.Q ),
    .A0(net73),
    .A1(net81),
    .A2(net65),
    .A3(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG9 ),
    .S1(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame2_bit17.Q ),
    .X(net279));
 sg13g2_mux4_1 _0519_ (.S0(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame2_bit18.Q ),
    .A0(net74),
    .A1(net67),
    .A2(net55),
    .A3(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG10 ),
    .S1(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame2_bit19.Q ),
    .X(net280));
 sg13g2_mux4_1 _0520_ (.S0(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame2_bit20.Q ),
    .A0(net75),
    .A1(net68),
    .A2(net56),
    .A3(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG11 ),
    .S1(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame2_bit21.Q ),
    .X(net281));
 sg13g2_mux4_1 _0521_ (.S0(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame2_bit22.Q ),
    .A0(net34),
    .A1(net76),
    .A2(net69),
    .A3(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG12 ),
    .S1(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame2_bit23.Q ),
    .X(net282));
 sg13g2_mux4_1 _0522_ (.S0(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame2_bit24.Q ),
    .A0(net35),
    .A1(net77),
    .A2(net70),
    .A3(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG13 ),
    .S1(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame2_bit25.Q ),
    .X(net283));
 sg13g2_mux4_1 _0523_ (.S0(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame2_bit26.Q ),
    .A0(net36),
    .A1(net78),
    .A2(net71),
    .A3(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG14 ),
    .S1(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame2_bit27.Q ),
    .X(net285));
 sg13g2_mux4_1 _0524_ (.S0(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame2_bit28.Q ),
    .A0(net37),
    .A1(net79),
    .A2(net72),
    .A3(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG15 ),
    .S1(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame2_bit29.Q ),
    .X(net286));
 sg13g2_nor3_1 _0525_ (.A(net46),
    .B(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame2_bit30.Q ),
    .C(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame2_bit31.Q ),
    .Y(_0092_));
 sg13g2_nand2b_1 _0526_ (.Y(_0093_),
    .B(net38),
    .A_N(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame2_bit31.Q ));
 sg13g2_a221oi_1 _0527_ (.B2(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame2_bit30.Q ),
    .C1(_0092_),
    .B1(_0093_),
    .A1(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame2_bit31.Q ),
    .Y(net256),
    .A2(_0038_));
 sg13g2_nor3_1 _0528_ (.A(net47),
    .B(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame1_bit0.Q ),
    .C(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame1_bit1.Q ),
    .Y(_0094_));
 sg13g2_nand2b_1 _0529_ (.Y(_0095_),
    .B(net39),
    .A_N(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame1_bit1.Q ));
 sg13g2_a221oi_1 _0530_ (.B2(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame1_bit0.Q ),
    .C1(_0094_),
    .B1(_0095_),
    .A1(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame1_bit1.Q ),
    .Y(net257),
    .A2(_0039_));
 sg13g2_nor3_1 _0531_ (.A(net48),
    .B(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame1_bit2.Q ),
    .C(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame1_bit3.Q ),
    .Y(_0096_));
 sg13g2_nand2b_1 _0532_ (.Y(_0097_),
    .B(net40),
    .A_N(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame1_bit3.Q ));
 sg13g2_a221oi_1 _0533_ (.B2(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame1_bit2.Q ),
    .C1(_0096_),
    .B1(_0097_),
    .A1(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame1_bit3.Q ),
    .Y(net258),
    .A2(_0040_));
 sg13g2_nor3_1 _0534_ (.A(net49),
    .B(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame1_bit4.Q ),
    .C(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame1_bit5.Q ),
    .Y(_0098_));
 sg13g2_nand2b_1 _0535_ (.Y(_0099_),
    .B(net41),
    .A_N(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame1_bit5.Q ));
 sg13g2_a221oi_1 _0536_ (.B2(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame1_bit4.Q ),
    .C1(_0098_),
    .B1(_0099_),
    .A1(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame1_bit5.Q ),
    .Y(net259),
    .A2(_0041_));
 sg13g2_nor3_1 _0537_ (.A(net50),
    .B(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame1_bit6.Q ),
    .C(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame1_bit7.Q ),
    .Y(_0100_));
 sg13g2_nand2b_1 _0538_ (.Y(_0101_),
    .B(net42),
    .A_N(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame1_bit7.Q ));
 sg13g2_a221oi_1 _0539_ (.B2(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame1_bit6.Q ),
    .C1(_0100_),
    .B1(_0101_),
    .A1(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame1_bit7.Q ),
    .Y(net260),
    .A2(_0042_));
 sg13g2_mux2_1 _0540_ (.A0(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG4 ),
    .A1(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG8 ),
    .S(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit14.Q ),
    .X(_0102_));
 sg13g2_nor2b_1 _0541_ (.A(net631),
    .B_N(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit14.Q ),
    .Y(_0103_));
 sg13g2_o21ai_1 _0542_ (.B1(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit15.Q ),
    .Y(_0104_),
    .A1(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit14.Q ),
    .A2(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG12 ));
 sg13g2_o21ai_1 _0543_ (.B1(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit16.Q ),
    .Y(_0105_),
    .A1(_0103_),
    .A2(_0104_));
 sg13g2_a21oi_1 _0544_ (.A1(_0011_),
    .A2(_0102_),
    .Y(_0106_),
    .B1(_0105_));
 sg13g2_mux4_1 _0545_ (.S0(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit14.Q ),
    .A0(net34),
    .A1(net66),
    .A2(net64),
    .A3(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG0 ),
    .S1(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit15.Q ),
    .X(_0107_));
 sg13g2_nor2_1 _0546_ (.A(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit16.Q ),
    .B(_0107_),
    .Y(_0108_));
 sg13g2_nor2_1 _0547_ (.A(_0106_),
    .B(_0108_),
    .Y(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.N4BEG0 ));
 sg13g2_mux2_1 _0548_ (.A0(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG5 ),
    .A1(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG9 ),
    .S(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit17.Q ),
    .X(_0109_));
 sg13g2_nor2b_1 _0549_ (.A(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS2_BEG1 ),
    .B_N(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit17.Q ),
    .Y(_0110_));
 sg13g2_o21ai_1 _0550_ (.B1(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit18.Q ),
    .Y(_0111_),
    .A1(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit17.Q ),
    .A2(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG13 ));
 sg13g2_o21ai_1 _0551_ (.B1(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit19.Q ),
    .Y(_0112_),
    .A1(_0110_),
    .A2(_0111_));
 sg13g2_a21oi_1 _0552_ (.A1(_0012_),
    .A2(_0109_),
    .Y(_0113_),
    .B1(_0112_));
 sg13g2_mux4_1 _0553_ (.S0(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit18.Q ),
    .A0(net35),
    .A1(net65),
    .A2(net73),
    .A3(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG1 ),
    .S1(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit17.Q ),
    .X(_0114_));
 sg13g2_nor2_1 _0554_ (.A(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit19.Q ),
    .B(_0114_),
    .Y(_0115_));
 sg13g2_nor2_1 _0555_ (.A(_0113_),
    .B(_0115_),
    .Y(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.N4BEG1 ));
 sg13g2_mux2_1 _0556_ (.A0(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG6 ),
    .A1(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG10 ),
    .S(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit20.Q ),
    .X(_0116_));
 sg13g2_nor2b_1 _0557_ (.A(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS2_BEG2 ),
    .B_N(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit20.Q ),
    .Y(_0117_));
 sg13g2_o21ai_1 _0558_ (.B1(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit21.Q ),
    .Y(_0118_),
    .A1(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit20.Q ),
    .A2(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG14 ));
 sg13g2_o21ai_1 _0559_ (.B1(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit22.Q ),
    .Y(_0119_),
    .A1(_0117_),
    .A2(_0118_));
 sg13g2_a21oi_1 _0560_ (.A1(_0013_),
    .A2(_0116_),
    .Y(_0120_),
    .B1(_0119_));
 sg13g2_mux4_1 _0561_ (.S0(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit21.Q ),
    .A0(net36),
    .A1(net55),
    .A2(net74),
    .A3(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG2 ),
    .S1(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit20.Q ),
    .X(_0121_));
 sg13g2_nor2_1 _0562_ (.A(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit22.Q ),
    .B(_0121_),
    .Y(_0122_));
 sg13g2_nor2_1 _0563_ (.A(_0120_),
    .B(_0122_),
    .Y(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.N4BEG2 ));
 sg13g2_mux2_1 _0564_ (.A0(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG7 ),
    .A1(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG11 ),
    .S(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit23.Q ),
    .X(_0123_));
 sg13g2_nor2b_1 _0565_ (.A(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS2_BEG3 ),
    .B_N(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit23.Q ),
    .Y(_0124_));
 sg13g2_o21ai_1 _0566_ (.B1(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit24.Q ),
    .Y(_0125_),
    .A1(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit23.Q ),
    .A2(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG15 ));
 sg13g2_o21ai_1 _0567_ (.B1(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit25.Q ),
    .Y(_0126_),
    .A1(_0124_),
    .A2(_0125_));
 sg13g2_a21oi_1 _0568_ (.A1(_0014_),
    .A2(_0123_),
    .Y(_0127_),
    .B1(_0126_));
 sg13g2_mux4_1 _0569_ (.S0(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit24.Q ),
    .A0(net37),
    .A1(net56),
    .A2(net75),
    .A3(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG3 ),
    .S1(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit23.Q ),
    .X(_0128_));
 sg13g2_nor2_1 _0570_ (.A(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit25.Q ),
    .B(_0128_),
    .Y(_0129_));
 sg13g2_nor2_1 _0571_ (.A(_0127_),
    .B(_0129_),
    .Y(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.N4BEG3 ));
 sg13g2_mux2_1 _0572_ (.A0(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG4 ),
    .A1(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG8 ),
    .S(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit18.Q ),
    .X(_0130_));
 sg13g2_nor2b_1 _0573_ (.A(net626),
    .B_N(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit18.Q ),
    .Y(_0131_));
 sg13g2_o21ai_1 _0574_ (.B1(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit19.Q ),
    .Y(_0132_),
    .A1(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit18.Q ),
    .A2(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG12 ));
 sg13g2_o21ai_1 _0575_ (.B1(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit20.Q ),
    .Y(_0133_),
    .A1(_0131_),
    .A2(_0132_));
 sg13g2_a21oi_1 _0576_ (.A1(_0015_),
    .A2(_0130_),
    .Y(_0134_),
    .B1(_0133_));
 sg13g2_mux4_1 _0577_ (.S0(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit18.Q ),
    .A0(net34),
    .A1(net69),
    .A2(net60),
    .A3(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG0 ),
    .S1(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit19.Q ),
    .X(_0135_));
 sg13g2_nor2_1 _0578_ (.A(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit20.Q ),
    .B(_0135_),
    .Y(_0136_));
 sg13g2_nor2_1 _0579_ (.A(_0134_),
    .B(_0136_),
    .Y(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.S4BEG0 ));
 sg13g2_mux2_1 _0580_ (.A0(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG5 ),
    .A1(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG9 ),
    .S(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit21.Q ),
    .X(_0137_));
 sg13g2_nor2b_1 _0581_ (.A(net625),
    .B_N(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit21.Q ),
    .Y(_0138_));
 sg13g2_o21ai_1 _0582_ (.B1(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit22.Q ),
    .Y(_0139_),
    .A1(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit21.Q ),
    .A2(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG13 ));
 sg13g2_o21ai_1 _0583_ (.B1(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit23.Q ),
    .Y(_0140_),
    .A1(_0138_),
    .A2(_0139_));
 sg13g2_a21oi_1 _0584_ (.A1(_0016_),
    .A2(_0137_),
    .Y(_0141_),
    .B1(_0140_));
 sg13g2_mux4_1 _0585_ (.S0(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit22.Q ),
    .A0(net35),
    .A1(net61),
    .A2(net70),
    .A3(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG1 ),
    .S1(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit21.Q ),
    .X(_0142_));
 sg13g2_nor2_1 _0586_ (.A(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit23.Q ),
    .B(_0142_),
    .Y(_0143_));
 sg13g2_nor2_1 _0587_ (.A(_0141_),
    .B(_0143_),
    .Y(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.S4BEG1 ));
 sg13g2_mux2_1 _0588_ (.A0(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG6 ),
    .A1(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG10 ),
    .S(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit24.Q ),
    .X(_0144_));
 sg13g2_nor2b_1 _0589_ (.A(net624),
    .B_N(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit24.Q ),
    .Y(_0145_));
 sg13g2_o21ai_1 _0590_ (.B1(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit25.Q ),
    .Y(_0146_),
    .A1(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit24.Q ),
    .A2(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG14 ));
 sg13g2_o21ai_1 _0591_ (.B1(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit26.Q ),
    .Y(_0147_),
    .A1(_0145_),
    .A2(_0146_));
 sg13g2_a21oi_1 _0592_ (.A1(_0017_),
    .A2(_0144_),
    .Y(_0148_),
    .B1(_0147_));
 sg13g2_mux4_1 _0593_ (.S0(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit25.Q ),
    .A0(net36),
    .A1(net62),
    .A2(net71),
    .A3(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG2 ),
    .S1(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit24.Q ),
    .X(_0149_));
 sg13g2_nor2_1 _0594_ (.A(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit26.Q ),
    .B(_0149_),
    .Y(_0150_));
 sg13g2_nor2_1 _0595_ (.A(_0148_),
    .B(_0150_),
    .Y(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.S4BEG2 ));
 sg13g2_mux2_1 _0596_ (.A0(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG7 ),
    .A1(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG11 ),
    .S(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit27.Q ),
    .X(_0151_));
 sg13g2_nor2b_1 _0597_ (.A(net623),
    .B_N(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit27.Q ),
    .Y(_0152_));
 sg13g2_o21ai_1 _0598_ (.B1(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit28.Q ),
    .Y(_0153_),
    .A1(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit27.Q ),
    .A2(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG15 ));
 sg13g2_o21ai_1 _0599_ (.B1(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit29.Q ),
    .Y(_0154_),
    .A1(_0152_),
    .A2(_0153_));
 sg13g2_a21oi_1 _0600_ (.A1(_0018_),
    .A2(_0151_),
    .Y(_0155_),
    .B1(_0154_));
 sg13g2_mux4_1 _0601_ (.S0(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit28.Q ),
    .A0(net37),
    .A1(net63),
    .A2(net72),
    .A3(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG3 ),
    .S1(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit27.Q ),
    .X(_0156_));
 sg13g2_nor2_1 _0602_ (.A(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit29.Q ),
    .B(_0156_),
    .Y(_0157_));
 sg13g2_nor2_1 _0603_ (.A(_0155_),
    .B(_0157_),
    .Y(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.S4BEG3 ));
 sg13g2_mux4_1 _0604_ (.S0(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame0_bit0.Q ),
    .A0(net223),
    .A1(net243),
    .A2(_0088_),
    .A3(net138),
    .S1(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame0_bit1.Q ),
    .X(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.J_NS4_BEG12 ));
 sg13g2_mux4_1 _0605_ (.S0(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame0_bit2.Q ),
    .A0(net224),
    .A1(net244),
    .A2(_0060_),
    .A3(net139),
    .S1(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame0_bit3.Q ),
    .X(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.J_NS4_BEG13 ));
 sg13g2_mux4_1 _0606_ (.S0(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame0_bit4.Q ),
    .A0(net225),
    .A1(net245),
    .A2(_0067_),
    .A3(net140),
    .S1(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame0_bit5.Q ),
    .X(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.J_NS4_BEG14 ));
 sg13g2_mux4_1 _0607_ (.S0(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame0_bit6.Q ),
    .A0(net226),
    .A1(net246),
    .A2(_0074_),
    .A3(net141),
    .S1(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame0_bit7.Q ),
    .X(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.J_NS4_BEG15 ));
 sg13g2_mux4_1 _0608_ (.S0(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame9_bit23.Q ),
    .A0(net34),
    .A1(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG12 ),
    .A2(net60),
    .A3(_0087_),
    .S1(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame9_bit22.Q ),
    .X(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.N1BEG0 ));
 sg13g2_mux4_1 _0609_ (.S0(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit14.Q ),
    .A0(net142),
    .A1(net172),
    .A2(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.J_NS4_BEG12 ),
    .A3(_0091_),
    .S1(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit15.Q ),
    .X(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.S1BEG0 ));
 sg13g2_mux4_1 _0610_ (.S0(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit16.Q ),
    .A0(net143),
    .A1(net173),
    .A2(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.J_NS4_BEG13 ),
    .A3(_0063_),
    .S1(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit17.Q ),
    .X(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.S1BEG1 ));
 sg13g2_mux4_1 _0611_ (.S0(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit18.Q ),
    .A0(net144),
    .A1(net163),
    .A2(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.J_NS4_BEG14 ),
    .A3(_0070_),
    .S1(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit19.Q ),
    .X(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.S1BEG2 ));
 sg13g2_mux4_1 _0612_ (.S0(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit20.Q ),
    .A0(net145),
    .A1(net164),
    .A2(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.J_NS4_BEG15 ),
    .A3(_0077_),
    .S1(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit21.Q ),
    .X(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.S1BEG3 ));
 sg13g2_mux4_1 _0613_ (.S0(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit22.Q ),
    .A0(net161),
    .A1(net153),
    .A2(net172),
    .A3(_0043_),
    .S1(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit23.Q ),
    .X(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.S2BEG0 ));
 sg13g2_mux4_1 _0614_ (.S0(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit24.Q ),
    .A0(net160),
    .A1(net152),
    .A2(net173),
    .A3(_0078_),
    .S1(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit25.Q ),
    .X(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.S2BEG1 ));
 sg13g2_mux4_1 _0615_ (.S0(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit27.Q ),
    .A0(net159),
    .A1(net163),
    .A2(net151),
    .A3(_0079_),
    .S1(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit26.Q ),
    .X(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.S2BEG2 ));
 sg13g2_mux4_1 _0616_ (.S0(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit29.Q ),
    .A0(net158),
    .A1(net164),
    .A2(net150),
    .A3(_0080_),
    .S1(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit28.Q ),
    .X(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.S2BEG3 ));
 sg13g2_mux4_1 _0617_ (.S0(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit31.Q ),
    .A0(net142),
    .A1(net149),
    .A2(net157),
    .A3(net635),
    .S1(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit30.Q ),
    .X(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.S2BEG4 ));
 sg13g2_mux4_1 _0618_ (.S0(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit0.Q ),
    .A0(net143),
    .A1(net156),
    .A2(net148),
    .A3(_0082_),
    .S1(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit1.Q ),
    .X(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.S2BEG5 ));
 sg13g2_mux4_1 _0619_ (.S0(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit2.Q ),
    .A0(net144),
    .A1(net155),
    .A2(net147),
    .A3(_0083_),
    .S1(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit3.Q ),
    .X(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.S2BEG6 ));
 sg13g2_mux4_1 _0620_ (.S0(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit5.Q ),
    .A0(net145),
    .A1(net146),
    .A2(net154),
    .A3(net632),
    .S1(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit4.Q ),
    .X(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.S2BEG7 ));
 sg13g2_mux4_1 _0621_ (.S0(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit19.Q ),
    .A0(net223),
    .A1(net14),
    .A2(_0088_),
    .A3(net31),
    .S1(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit18.Q ),
    .X(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.W1BEG0 ));
 sg13g2_mux4_1 _0622_ (.S0(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit21.Q ),
    .A0(net224),
    .A1(net25),
    .A2(_0060_),
    .A3(net30),
    .S1(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit20.Q ),
    .X(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.W1BEG1 ));
 sg13g2_mux4_1 _0623_ (.S0(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit23.Q ),
    .A0(net225),
    .A1(net2),
    .A2(_0067_),
    .A3(net29),
    .S1(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit22.Q ),
    .X(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.W1BEG2 ));
 sg13g2_mux4_1 _0624_ (.S0(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit25.Q ),
    .A0(net226),
    .A1(net3),
    .A2(_0074_),
    .A3(net28),
    .S1(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit24.Q ),
    .X(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.W1BEG3 ));
 sg13g2_mux4_1 _0625_ (.S0(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit26.Q ),
    .A0(net2),
    .A1(net32),
    .A2(net640),
    .A3(net632),
    .S1(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit27.Q ),
    .X(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.W2BEG0 ));
 sg13g2_mux4_1 _0626_ (.S0(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit28.Q ),
    .A0(net3),
    .A1(net33),
    .A2(net639),
    .A3(net633),
    .S1(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit29.Q ),
    .X(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.W2BEG1 ));
 sg13g2_mux4_1 _0627_ (.S0(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit30.Q ),
    .A0(net14),
    .A1(net4),
    .A2(net638),
    .A3(net634),
    .S1(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit31.Q ),
    .X(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.W2BEG2 ));
 sg13g2_mux4_1 _0628_ (.S0(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame6_bit0.Q ),
    .A0(net25),
    .A1(net5),
    .A2(net637),
    .A3(net636),
    .S1(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame6_bit1.Q ),
    .X(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.W2BEG3 ));
 sg13g2_mux4_1 _0629_ (.S0(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame6_bit2.Q ),
    .A0(net28),
    .A1(net6),
    .A2(net637),
    .A3(net635),
    .S1(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame6_bit3.Q ),
    .X(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.W2BEG4 ));
 sg13g2_mux4_1 _0630_ (.S0(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame6_bit4.Q ),
    .A0(net29),
    .A1(net7),
    .A2(net638),
    .A3(net634),
    .S1(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame6_bit5.Q ),
    .X(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.W2BEG5 ));
 sg13g2_mux4_1 _0631_ (.S0(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame6_bit6.Q ),
    .A0(net30),
    .A1(net8),
    .A2(net639),
    .A3(net633),
    .S1(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame6_bit7.Q ),
    .X(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.W2BEG6 ));
 sg13g2_mux4_1 _0632_ (.S0(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame6_bit8.Q ),
    .A0(net31),
    .A1(net9),
    .A2(net640),
    .A3(net632),
    .S1(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame6_bit9.Q ),
    .X(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.W2BEG7 ));
 sg13g2_mux4_1 _0633_ (.S0(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame6_bit10.Q ),
    .A0(net2),
    .A1(net32),
    .A2(net640),
    .A3(net632),
    .S1(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame6_bit11.Q ),
    .X(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.W2BEGb0 ));
 sg13g2_mux4_1 _0634_ (.S0(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame6_bit12.Q ),
    .A0(net3),
    .A1(net33),
    .A2(net639),
    .A3(net633),
    .S1(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame6_bit13.Q ),
    .X(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.W2BEGb1 ));
 sg13g2_mux4_1 _0635_ (.S0(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame6_bit14.Q ),
    .A0(net14),
    .A1(net4),
    .A2(net638),
    .A3(net634),
    .S1(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame6_bit15.Q ),
    .X(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.W2BEGb2 ));
 sg13g2_mux4_1 _0636_ (.S0(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame6_bit16.Q ),
    .A0(net25),
    .A1(net5),
    .A2(net637),
    .A3(net635),
    .S1(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame6_bit17.Q ),
    .X(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.W2BEGb3 ));
 sg13g2_mux4_1 _0637_ (.S0(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame6_bit18.Q ),
    .A0(net28),
    .A1(net6),
    .A2(net637),
    .A3(net635),
    .S1(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame6_bit19.Q ),
    .X(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.W2BEGb4 ));
 sg13g2_mux4_1 _0638_ (.S0(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame6_bit20.Q ),
    .A0(net29),
    .A1(net7),
    .A2(net638),
    .A3(net634),
    .S1(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame6_bit21.Q ),
    .X(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.W2BEGb5 ));
 sg13g2_mux4_1 _0639_ (.S0(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame6_bit22.Q ),
    .A0(net30),
    .A1(net8),
    .A2(net639),
    .A3(net633),
    .S1(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame6_bit23.Q ),
    .X(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.W2BEGb6 ));
 sg13g2_mux4_1 _0640_ (.S0(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame6_bit24.Q ),
    .A0(net31),
    .A1(net9),
    .A2(net640),
    .A3(net632),
    .S1(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame6_bit25.Q ),
    .X(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.W2BEGb7 ));
 sg13g2_mux4_1 _0641_ (.S0(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame6_bit26.Q ),
    .A0(net2),
    .A1(net6),
    .A2(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.J_NS4_BEG15 ),
    .A3(net632),
    .S1(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame6_bit27.Q ),
    .X(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.WW4BEG0 ));
 sg13g2_mux4_1 _0642_ (.S0(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame6_bit28.Q ),
    .A0(net3),
    .A1(net7),
    .A2(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.J_NS4_BEG14 ),
    .A3(net633),
    .S1(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame6_bit29.Q ),
    .X(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.WW4BEG1 ));
 sg13g2_mux4_1 _0643_ (.S0(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame6_bit30.Q ),
    .A0(net14),
    .A1(net8),
    .A2(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.J_NS4_BEG13 ),
    .A3(net634),
    .S1(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame6_bit31.Q ),
    .X(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.WW4BEG2 ));
 sg13g2_mux4_1 _0644_ (.S0(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame5_bit0.Q ),
    .A0(net25),
    .A1(net9),
    .A2(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.J_NS4_BEG12 ),
    .A3(net635),
    .S1(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame5_bit1.Q ),
    .X(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.WW4BEG3 ));
 sg13g2_mux4_1 _0645_ (.S0(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit30.Q ),
    .A0(net226),
    .A1(net246),
    .A2(_0074_),
    .A3(net141),
    .S1(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit31.Q ),
    .X(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.J_NS4_BEG11 ));
 sg13g2_mux4_1 _0646_ (.S0(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame5_bit2.Q ),
    .A0(net28),
    .A1(net32),
    .A2(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.J_NS4_BEG11 ),
    .A3(net637),
    .S1(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame5_bit3.Q ),
    .X(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.WW4BEG4 ));
 sg13g2_mux4_1 _0647_ (.S0(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit28.Q ),
    .A0(net225),
    .A1(net245),
    .A2(_0067_),
    .A3(net140),
    .S1(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit29.Q ),
    .X(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.J_NS4_BEG10 ));
 sg13g2_mux4_1 _0648_ (.S0(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame5_bit4.Q ),
    .A0(net29),
    .A1(net33),
    .A2(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.J_NS4_BEG10 ),
    .A3(net638),
    .S1(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame5_bit5.Q ),
    .X(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.WW4BEG5 ));
 sg13g2_mux4_1 _0649_ (.S0(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit26.Q ),
    .A0(net224),
    .A1(net244),
    .A2(_0060_),
    .A3(net139),
    .S1(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit27.Q ),
    .X(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.J_NS4_BEG9 ));
 sg13g2_mux4_1 _0650_ (.S0(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame5_bit6.Q ),
    .A0(net30),
    .A1(net4),
    .A2(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.J_NS4_BEG9 ),
    .A3(net639),
    .S1(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame5_bit7.Q ),
    .X(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.WW4BEG6 ));
 sg13g2_mux4_1 _0651_ (.S0(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit24.Q ),
    .A0(net223),
    .A1(net243),
    .A2(_0088_),
    .A3(net138),
    .S1(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit25.Q ),
    .X(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.J_NS4_BEG8 ));
 sg13g2_mux4_1 _0652_ (.S0(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame5_bit8.Q ),
    .A0(net31),
    .A1(net5),
    .A2(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.J_NS4_BEG8 ),
    .A3(net640),
    .S1(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame5_bit9.Q ),
    .X(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.WW4BEG7 ));
 sg13g2_mux4_1 _0653_ (.S0(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit22.Q ),
    .A0(net226),
    .A1(net246),
    .A2(_0074_),
    .A3(net141),
    .S1(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit23.Q ),
    .X(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.J_NS4_BEG7 ));
 sg13g2_mux4_1 _0654_ (.S0(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame5_bit10.Q ),
    .A0(net28),
    .A1(net32),
    .A2(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.J_NS4_BEG7 ),
    .A3(net632),
    .S1(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame5_bit11.Q ),
    .X(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.WW4BEG8 ));
 sg13g2_mux4_1 _0655_ (.S0(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit20.Q ),
    .A0(net225),
    .A1(net245),
    .A2(_0067_),
    .A3(net140),
    .S1(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit21.Q ),
    .X(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.J_NS4_BEG6 ));
 sg13g2_mux4_1 _0656_ (.S0(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame5_bit12.Q ),
    .A0(net29),
    .A1(net33),
    .A2(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.J_NS4_BEG6 ),
    .A3(net633),
    .S1(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame5_bit13.Q ),
    .X(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.WW4BEG9 ));
 sg13g2_mux4_1 _0657_ (.S0(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit18.Q ),
    .A0(net224),
    .A1(net244),
    .A2(_0060_),
    .A3(net139),
    .S1(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit19.Q ),
    .X(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.J_NS4_BEG5 ));
 sg13g2_mux4_1 _0658_ (.S0(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame5_bit14.Q ),
    .A0(net30),
    .A1(net4),
    .A2(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.J_NS4_BEG5 ),
    .A3(net634),
    .S1(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame5_bit15.Q ),
    .X(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.WW4BEG10 ));
 sg13g2_mux4_1 _0659_ (.S0(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit16.Q ),
    .A0(net223),
    .A1(net243),
    .A2(_0088_),
    .A3(net138),
    .S1(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit17.Q ),
    .X(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.J_NS4_BEG4 ));
 sg13g2_mux4_1 _0660_ (.S0(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame5_bit16.Q ),
    .A0(net31),
    .A1(net5),
    .A2(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.J_NS4_BEG4 ),
    .A3(net635),
    .S1(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame5_bit17.Q ),
    .X(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.WW4BEG11 ));
 sg13g2_mux4_1 _0661_ (.S0(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit14.Q ),
    .A0(net226),
    .A1(net246),
    .A2(_0074_),
    .A3(net141),
    .S1(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit15.Q ),
    .X(_0158_));
 sg13g2_mux4_1 _0662_ (.S0(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame5_bit18.Q ),
    .A0(net2),
    .A1(net6),
    .A2(_0158_),
    .A3(net637),
    .S1(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame5_bit19.Q ),
    .X(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.WW4BEG12 ));
 sg13g2_mux4_1 _0663_ (.S0(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit12.Q ),
    .A0(net225),
    .A1(net245),
    .A2(_0067_),
    .A3(net140),
    .S1(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit13.Q ),
    .X(_0159_));
 sg13g2_mux4_1 _0664_ (.S0(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame5_bit20.Q ),
    .A0(net3),
    .A1(net7),
    .A2(_0159_),
    .A3(net638),
    .S1(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame5_bit21.Q ),
    .X(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.WW4BEG13 ));
 sg13g2_mux4_1 _0665_ (.S0(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit10.Q ),
    .A0(net224),
    .A1(net244),
    .A2(_0060_),
    .A3(net139),
    .S1(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit11.Q ),
    .X(_0160_));
 sg13g2_mux4_1 _0666_ (.S0(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame5_bit22.Q ),
    .A0(net14),
    .A1(net8),
    .A2(_0160_),
    .A3(net639),
    .S1(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame5_bit23.Q ),
    .X(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.WW4BEG14 ));
 sg13g2_mux4_1 _0667_ (.S0(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit8.Q ),
    .A0(net223),
    .A1(net243),
    .A2(_0088_),
    .A3(net138),
    .S1(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit9.Q ),
    .X(_0161_));
 sg13g2_mux4_1 _0668_ (.S0(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame5_bit24.Q ),
    .A0(net25),
    .A1(net9),
    .A2(_0161_),
    .A3(_0043_),
    .S1(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame5_bit25.Q ),
    .X(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.WW4BEG15 ));
 sg13g2_mux4_1 _0669_ (.S0(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame5_bit26.Q ),
    .A0(net243),
    .A1(net138),
    .A2(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.J_NS4_BEG11 ),
    .A3(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.J_NS4_BEG15 ),
    .S1(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame5_bit27.Q ),
    .X(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.W6BEG0 ));
 sg13g2_mux4_1 _0670_ (.S0(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame5_bit28.Q ),
    .A0(net244),
    .A1(net139),
    .A2(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.J_NS4_BEG10 ),
    .A3(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.J_NS4_BEG14 ),
    .S1(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame5_bit29.Q ),
    .X(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.W6BEG1 ));
 sg13g2_mux4_1 _0671_ (.S0(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame5_bit30.Q ),
    .A0(net245),
    .A1(net140),
    .A2(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.J_NS4_BEG9 ),
    .A3(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.J_NS4_BEG13 ),
    .S1(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame5_bit31.Q ),
    .X(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.W6BEG2 ));
 sg13g2_mux4_1 _0672_ (.S0(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame4_bit0.Q ),
    .A0(net246),
    .A1(net141),
    .A2(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.J_NS4_BEG8 ),
    .A3(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.J_NS4_BEG12 ),
    .S1(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame4_bit1.Q ),
    .X(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.W6BEG3 ));
 sg13g2_mux4_1 _0673_ (.S0(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame4_bit3.Q ),
    .A0(net28),
    .A1(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.J_NS4_BEG11 ),
    .A2(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.J_NS4_BEG7 ),
    .A3(net640),
    .S1(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame4_bit2.Q ),
    .X(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.W6BEG4 ));
 sg13g2_mux4_1 _0674_ (.S0(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame4_bit5.Q ),
    .A0(net29),
    .A1(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.J_NS4_BEG10 ),
    .A2(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.J_NS4_BEG6 ),
    .A3(net639),
    .S1(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame4_bit4.Q ),
    .X(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.W6BEG5 ));
 sg13g2_mux4_1 _0675_ (.S0(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame4_bit6.Q ),
    .A0(net30),
    .A1(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.J_NS4_BEG5 ),
    .A2(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.J_NS4_BEG9 ),
    .A3(net638),
    .S1(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame4_bit7.Q ),
    .X(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.W6BEG6 ));
 sg13g2_mux4_1 _0676_ (.S0(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame4_bit8.Q ),
    .A0(net31),
    .A1(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.J_NS4_BEG4 ),
    .A2(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.J_NS4_BEG8 ),
    .A3(net637),
    .S1(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame4_bit9.Q ),
    .X(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.W6BEG7 ));
 sg13g2_mux4_1 _0677_ (.S0(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame4_bit11.Q ),
    .A0(net2),
    .A1(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.J_NS4_BEG7 ),
    .A2(_0158_),
    .A3(net635),
    .S1(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame4_bit10.Q ),
    .X(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.W6BEG8 ));
 sg13g2_mux4_1 _0678_ (.S0(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame4_bit13.Q ),
    .A0(net3),
    .A1(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.J_NS4_BEG6 ),
    .A2(_0159_),
    .A3(net634),
    .S1(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame4_bit12.Q ),
    .X(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.W6BEG9 ));
 sg13g2_mux4_1 _0679_ (.S0(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame4_bit15.Q ),
    .A0(net14),
    .A1(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.J_NS4_BEG5 ),
    .A2(_0160_),
    .A3(net633),
    .S1(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame4_bit14.Q ),
    .X(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.W6BEG10 ));
 sg13g2_mux4_1 _0680_ (.S0(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame4_bit17.Q ),
    .A0(net25),
    .A1(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.J_NS4_BEG4 ),
    .A2(_0161_),
    .A3(net632),
    .S1(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame4_bit16.Q ),
    .X(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.W6BEG11 ));
 sg13g2_nand3b_1 _0681_ (.B(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame4_bit19.Q ),
    .C(net640),
    .Y(_0162_),
    .A_N(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame4_bit18.Q ));
 sg13g2_nor2b_1 _0682_ (.A(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame4_bit18.Q ),
    .B_N(net154),
    .Y(_0163_));
 sg13g2_a21oi_1 _0683_ (.A1(net146),
    .A2(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame4_bit18.Q ),
    .Y(_0164_),
    .B1(_0163_));
 sg13g2_o21ai_1 _0684_ (.B1(_0162_),
    .Y(net251),
    .A1(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame4_bit19.Q ),
    .A2(_0164_));
 sg13g2_nand3b_1 _0685_ (.B(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame4_bit21.Q ),
    .C(_0078_),
    .Y(_0165_),
    .A_N(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame4_bit20.Q ));
 sg13g2_nor2b_1 _0686_ (.A(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame4_bit20.Q ),
    .B_N(net155),
    .Y(_0166_));
 sg13g2_a21oi_1 _0687_ (.A1(net147),
    .A2(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame4_bit20.Q ),
    .Y(_0167_),
    .B1(_0166_));
 sg13g2_o21ai_1 _0688_ (.B1(_0165_),
    .Y(net252),
    .A1(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame4_bit21.Q ),
    .A2(_0167_));
 sg13g2_nand3b_1 _0689_ (.B(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame4_bit23.Q ),
    .C(net638),
    .Y(_0168_),
    .A_N(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame4_bit22.Q ));
 sg13g2_nor2b_1 _0690_ (.A(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame4_bit22.Q ),
    .B_N(net156),
    .Y(_0169_));
 sg13g2_a21oi_1 _0691_ (.A1(net148),
    .A2(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame4_bit22.Q ),
    .Y(_0170_),
    .B1(_0169_));
 sg13g2_o21ai_1 _0692_ (.B1(_0168_),
    .Y(net253),
    .A1(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame4_bit23.Q ),
    .A2(_0170_));
 sg13g2_nand3b_1 _0693_ (.B(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame4_bit25.Q ),
    .C(net637),
    .Y(_0171_),
    .A_N(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame4_bit24.Q ));
 sg13g2_nor2_1 _0694_ (.A(_0000_),
    .B(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame4_bit24.Q ),
    .Y(_0172_));
 sg13g2_a21oi_1 _0695_ (.A1(net149),
    .A2(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame4_bit24.Q ),
    .Y(_0173_),
    .B1(_0172_));
 sg13g2_o21ai_1 _0696_ (.B1(_0171_),
    .Y(net254),
    .A1(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame4_bit25.Q ),
    .A2(_0173_));
 sg13g2_nand3b_1 _0697_ (.B(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame4_bit27.Q ),
    .C(net635),
    .Y(_0174_),
    .A_N(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame4_bit26.Q ));
 sg13g2_nor2b_1 _0698_ (.A(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame4_bit26.Q ),
    .B_N(net158),
    .Y(_0175_));
 sg13g2_a21oi_1 _0699_ (.A1(net150),
    .A2(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame4_bit26.Q ),
    .Y(_0176_),
    .B1(_0175_));
 sg13g2_o21ai_1 _0700_ (.B1(_0174_),
    .Y(net255),
    .A1(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame4_bit27.Q ),
    .A2(_0176_));
 sg13g2_mux4_1 _0701_ (.S0(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame4_bit28.Q ),
    .A0(net174),
    .A1(net188),
    .A2(net162),
    .A3(_0161_),
    .S1(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame4_bit29.Q ),
    .X(net261));
 sg13g2_mux4_1 _0702_ (.S0(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame4_bit30.Q ),
    .A0(net181),
    .A1(net189),
    .A2(net165),
    .A3(_0160_),
    .S1(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame4_bit31.Q ),
    .X(net262));
 sg13g2_mux4_1 _0703_ (.S0(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame3_bit0.Q ),
    .A0(net182),
    .A1(net175),
    .A2(net166),
    .A3(_0159_),
    .S1(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame3_bit1.Q ),
    .X(net273));
 sg13g2_mux4_1 _0704_ (.S0(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame3_bit2.Q ),
    .A0(net183),
    .A1(net176),
    .A2(net167),
    .A3(_0158_),
    .S1(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame3_bit3.Q ),
    .X(net284));
 sg13g2_mux4_1 _0705_ (.S0(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame3_bit4.Q ),
    .A0(net184),
    .A1(net177),
    .A2(net168),
    .A3(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.J_NS4_BEG4 ),
    .S1(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame3_bit5.Q ),
    .X(net287));
 sg13g2_mux4_1 _0706_ (.S0(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame3_bit6.Q ),
    .A0(net185),
    .A1(net178),
    .A2(net169),
    .A3(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.J_NS4_BEG5 ),
    .S1(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame3_bit7.Q ),
    .X(net288));
 sg13g2_mux4_1 _0707_ (.S0(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame3_bit8.Q ),
    .A0(net186),
    .A1(net179),
    .A2(net170),
    .A3(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.J_NS4_BEG6 ),
    .S1(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame3_bit9.Q ),
    .X(net289));
 sg13g2_mux4_1 _0708_ (.S0(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame3_bit10.Q ),
    .A0(net187),
    .A1(net180),
    .A2(net171),
    .A3(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.J_NS4_BEG7 ),
    .S1(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame3_bit11.Q ),
    .X(net290));
 sg13g2_mux4_1 _0709_ (.S0(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame3_bit12.Q ),
    .A0(net174),
    .A1(net188),
    .A2(net172),
    .A3(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.J_NS4_BEG8 ),
    .S1(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame3_bit13.Q ),
    .X(net291));
 sg13g2_mux4_1 _0710_ (.S0(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame3_bit14.Q ),
    .A0(net181),
    .A1(net189),
    .A2(net173),
    .A3(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.J_NS4_BEG9 ),
    .S1(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame3_bit15.Q ),
    .X(net292));
 sg13g2_mux4_1 _0711_ (.S0(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame3_bit16.Q ),
    .A0(net182),
    .A1(net175),
    .A2(net163),
    .A3(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.J_NS4_BEG10 ),
    .S1(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame3_bit17.Q ),
    .X(net263));
 sg13g2_mux4_1 _0712_ (.S0(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame3_bit18.Q ),
    .A0(net183),
    .A1(net176),
    .A2(net164),
    .A3(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.J_NS4_BEG11 ),
    .S1(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame3_bit19.Q ),
    .X(net264));
 sg13g2_mux4_1 _0713_ (.S0(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame3_bit20.Q ),
    .A0(net142),
    .A1(net184),
    .A2(net177),
    .A3(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.J_NS4_BEG12 ),
    .S1(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame3_bit21.Q ),
    .X(net265));
 sg13g2_mux4_1 _0714_ (.S0(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame3_bit22.Q ),
    .A0(net143),
    .A1(net185),
    .A2(net178),
    .A3(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.J_NS4_BEG13 ),
    .S1(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame3_bit23.Q ),
    .X(net266));
 sg13g2_mux4_1 _0715_ (.S0(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame3_bit24.Q ),
    .A0(net144),
    .A1(net186),
    .A2(net179),
    .A3(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.J_NS4_BEG14 ),
    .S1(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame3_bit25.Q ),
    .X(net267));
 sg13g2_mux4_1 _0716_ (.S0(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame3_bit26.Q ),
    .A0(net145),
    .A1(net187),
    .A2(net180),
    .A3(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.J_NS4_BEG15 ),
    .S1(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame3_bit27.Q ),
    .X(net268));
 sg13g2_mux4_1 _0717_ (.S0(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame3_bit28.Q ),
    .A0(net174),
    .A1(net188),
    .A2(net162),
    .A3(_0161_),
    .S1(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame3_bit29.Q ),
    .X(net294));
 sg13g2_mux4_1 _0718_ (.S0(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame3_bit30.Q ),
    .A0(net181),
    .A1(net189),
    .A2(net165),
    .A3(_0160_),
    .S1(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame3_bit31.Q ),
    .X(net295));
 sg13g2_mux4_1 _0719_ (.S0(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit0.Q ),
    .A0(net182),
    .A1(net175),
    .A2(net166),
    .A3(_0159_),
    .S1(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit1.Q ),
    .X(net306));
 sg13g2_mux4_1 _0720_ (.S0(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit2.Q ),
    .A0(net183),
    .A1(net176),
    .A2(net167),
    .A3(_0158_),
    .S1(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit3.Q ),
    .X(net317));
 sg13g2_mux4_1 _0721_ (.S0(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit4.Q ),
    .A0(net184),
    .A1(net177),
    .A2(net168),
    .A3(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.J_NS4_BEG4 ),
    .S1(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit5.Q ),
    .X(net320));
 sg13g2_mux4_1 _0722_ (.S0(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit6.Q ),
    .A0(net185),
    .A1(net178),
    .A2(net169),
    .A3(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.J_NS4_BEG5 ),
    .S1(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit7.Q ),
    .X(net321));
 sg13g2_mux4_1 _0723_ (.S0(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit8.Q ),
    .A0(net186),
    .A1(net179),
    .A2(net170),
    .A3(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.J_NS4_BEG6 ),
    .S1(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit9.Q ),
    .X(net322));
 sg13g2_mux4_1 _0724_ (.S0(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit10.Q ),
    .A0(net187),
    .A1(net180),
    .A2(net171),
    .A3(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.J_NS4_BEG7 ),
    .S1(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit11.Q ),
    .X(net323));
 sg13g2_mux4_1 _0725_ (.S0(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit12.Q ),
    .A0(net174),
    .A1(net188),
    .A2(net172),
    .A3(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.J_NS4_BEG8 ),
    .S1(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit13.Q ),
    .X(net324));
 sg13g2_mux4_1 _0726_ (.S0(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit14.Q ),
    .A0(net181),
    .A1(net189),
    .A2(net173),
    .A3(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.J_NS4_BEG9 ),
    .S1(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit15.Q ),
    .X(net325));
 sg13g2_mux4_1 _0727_ (.S0(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit16.Q ),
    .A0(net182),
    .A1(net175),
    .A2(net163),
    .A3(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.J_NS4_BEG10 ),
    .S1(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit17.Q ),
    .X(net296));
 sg13g2_mux4_1 _0728_ (.S0(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit18.Q ),
    .A0(net183),
    .A1(net176),
    .A2(net164),
    .A3(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.J_NS4_BEG11 ),
    .S1(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit19.Q ),
    .X(net297));
 sg13g2_mux4_1 _0729_ (.S0(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit20.Q ),
    .A0(net142),
    .A1(net184),
    .A2(net177),
    .A3(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.J_NS4_BEG12 ),
    .S1(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit21.Q ),
    .X(net298));
 sg13g2_mux4_1 _0730_ (.S0(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit22.Q ),
    .A0(net143),
    .A1(net185),
    .A2(net178),
    .A3(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.J_NS4_BEG13 ),
    .S1(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit23.Q ),
    .X(net299));
 sg13g2_mux4_1 _0731_ (.S0(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit24.Q ),
    .A0(net144),
    .A1(net186),
    .A2(net179),
    .A3(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.J_NS4_BEG14 ),
    .S1(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit25.Q ),
    .X(net300));
 sg13g2_mux4_1 _0732_ (.S0(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit26.Q ),
    .A0(net145),
    .A1(net187),
    .A2(net180),
    .A3(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.J_NS4_BEG15 ),
    .S1(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit27.Q ),
    .X(net301));
 sg13g2_o21ai_1 _0733_ (.B1(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit3.Q ),
    .Y(_0177_),
    .A1(net172),
    .A2(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit2.Q ));
 sg13g2_inv_1 _0734_ (.Y(_0178_),
    .A(_0177_));
 sg13g2_o21ai_1 _0735_ (.B1(_0178_),
    .Y(_0179_),
    .A1(_0019_),
    .A2(_0161_));
 sg13g2_mux2_1 _0736_ (.A0(net142),
    .A1(net174),
    .S(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit2.Q ),
    .X(_0180_));
 sg13g2_a21oi_1 _0737_ (.A1(_0020_),
    .A2(_0180_),
    .Y(_0181_),
    .B1(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit4.Q ));
 sg13g2_nor2_1 _0738_ (.A(_0019_),
    .B(_0043_),
    .Y(_0182_));
 sg13g2_o21ai_1 _0739_ (.B1(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit3.Q ),
    .Y(_0183_),
    .A1(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit2.Q ),
    .A2(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.J_NS4_BEG12 ));
 sg13g2_mux2_1 _0740_ (.A0(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.J_NS4_BEG4 ),
    .A1(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.J_NS4_BEG8 ),
    .S(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit2.Q ),
    .X(_0184_));
 sg13g2_o21ai_1 _0741_ (.B1(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit4.Q ),
    .Y(_0185_),
    .A1(_0182_),
    .A2(_0183_));
 sg13g2_a21oi_1 _0742_ (.A1(_0020_),
    .A2(_0184_),
    .Y(_0186_),
    .B1(_0185_));
 sg13g2_a21oi_1 _0743_ (.A1(_0179_),
    .A2(_0181_),
    .Y(\Tile_X0Y0_IHP_SRAM_top.N4BEG_outbuf_8.A ),
    .B1(_0186_));
 sg13g2_o21ai_1 _0744_ (.B1(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit6.Q ),
    .Y(_0187_),
    .A1(net173),
    .A2(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit5.Q ));
 sg13g2_inv_1 _0745_ (.Y(_0188_),
    .A(_0187_));
 sg13g2_o21ai_1 _0746_ (.B1(_0188_),
    .Y(_0189_),
    .A1(_0021_),
    .A2(_0160_));
 sg13g2_mux2_1 _0747_ (.A0(net143),
    .A1(net181),
    .S(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit5.Q ),
    .X(_0190_));
 sg13g2_a21oi_1 _0748_ (.A1(_0022_),
    .A2(_0190_),
    .Y(_0191_),
    .B1(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit7.Q ));
 sg13g2_nor2_1 _0749_ (.A(_0021_),
    .B(net639),
    .Y(_0192_));
 sg13g2_o21ai_1 _0750_ (.B1(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit6.Q ),
    .Y(_0193_),
    .A1(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit5.Q ),
    .A2(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.J_NS4_BEG13 ));
 sg13g2_mux2_1 _0751_ (.A0(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.J_NS4_BEG5 ),
    .A1(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.J_NS4_BEG9 ),
    .S(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit5.Q ),
    .X(_0194_));
 sg13g2_o21ai_1 _0752_ (.B1(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit7.Q ),
    .Y(_0195_),
    .A1(_0192_),
    .A2(_0193_));
 sg13g2_a21oi_1 _0753_ (.A1(_0022_),
    .A2(_0194_),
    .Y(_0196_),
    .B1(_0195_));
 sg13g2_a21oi_1 _0754_ (.A1(_0189_),
    .A2(_0191_),
    .Y(\Tile_X0Y0_IHP_SRAM_top.N4BEG_outbuf_9.A ),
    .B1(_0196_));
 sg13g2_o21ai_1 _0755_ (.B1(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit9.Q ),
    .Y(_0197_),
    .A1(net163),
    .A2(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit8.Q ));
 sg13g2_inv_1 _0756_ (.Y(_0198_),
    .A(_0197_));
 sg13g2_o21ai_1 _0757_ (.B1(_0198_),
    .Y(_0199_),
    .A1(_0023_),
    .A2(_0159_));
 sg13g2_mux2_1 _0758_ (.A0(net144),
    .A1(net182),
    .S(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit8.Q ),
    .X(_0200_));
 sg13g2_a21oi_1 _0759_ (.A1(_0024_),
    .A2(_0200_),
    .Y(_0201_),
    .B1(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit10.Q ));
 sg13g2_nor2_1 _0760_ (.A(_0023_),
    .B(_0079_),
    .Y(_0202_));
 sg13g2_o21ai_1 _0761_ (.B1(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit9.Q ),
    .Y(_0203_),
    .A1(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit8.Q ),
    .A2(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.J_NS4_BEG14 ));
 sg13g2_mux2_1 _0762_ (.A0(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.J_NS4_BEG6 ),
    .A1(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.J_NS4_BEG10 ),
    .S(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit8.Q ),
    .X(_0204_));
 sg13g2_o21ai_1 _0763_ (.B1(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit10.Q ),
    .Y(_0205_),
    .A1(_0202_),
    .A2(_0203_));
 sg13g2_a21oi_1 _0764_ (.A1(_0024_),
    .A2(_0204_),
    .Y(_0206_),
    .B1(_0205_));
 sg13g2_a21oi_1 _0765_ (.A1(_0199_),
    .A2(_0201_),
    .Y(\Tile_X0Y0_IHP_SRAM_top.N4BEG_outbuf_10.A ),
    .B1(_0206_));
 sg13g2_o21ai_1 _0766_ (.B1(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit12.Q ),
    .Y(_0207_),
    .A1(net164),
    .A2(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit11.Q ));
 sg13g2_inv_1 _0767_ (.Y(_0208_),
    .A(_0207_));
 sg13g2_o21ai_1 _0768_ (.B1(_0208_),
    .Y(_0209_),
    .A1(_0025_),
    .A2(_0158_));
 sg13g2_mux2_1 _0769_ (.A0(net145),
    .A1(net183),
    .S(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit11.Q ),
    .X(_0210_));
 sg13g2_a21oi_1 _0770_ (.A1(_0026_),
    .A2(_0210_),
    .Y(_0211_),
    .B1(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit13.Q ));
 sg13g2_nor2_1 _0771_ (.A(_0025_),
    .B(_0080_),
    .Y(_0212_));
 sg13g2_o21ai_1 _0772_ (.B1(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit12.Q ),
    .Y(_0213_),
    .A1(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit11.Q ),
    .A2(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.J_NS4_BEG15 ));
 sg13g2_mux2_1 _0773_ (.A0(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.J_NS4_BEG7 ),
    .A1(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.J_NS4_BEG11 ),
    .S(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit11.Q ),
    .X(_0214_));
 sg13g2_o21ai_1 _0774_ (.B1(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit13.Q ),
    .Y(_0215_),
    .A1(_0212_),
    .A2(_0213_));
 sg13g2_a21oi_1 _0775_ (.A1(_0026_),
    .A2(_0214_),
    .Y(_0216_),
    .B1(_0215_));
 sg13g2_a21oi_1 _0776_ (.A1(_0209_),
    .A2(_0211_),
    .Y(\Tile_X0Y0_IHP_SRAM_top.N4BEG_outbuf_11.A ),
    .B1(_0216_));
 sg13g2_o21ai_1 _0777_ (.B1(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit7.Q ),
    .Y(_0217_),
    .A1(net168),
    .A2(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit6.Q ));
 sg13g2_inv_1 _0778_ (.Y(_0218_),
    .A(_0217_));
 sg13g2_o21ai_1 _0779_ (.B1(_0218_),
    .Y(_0219_),
    .A1(_0027_),
    .A2(_0161_));
 sg13g2_mux2_1 _0780_ (.A0(net142),
    .A1(net177),
    .S(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit6.Q ),
    .X(_0220_));
 sg13g2_a21oi_1 _0781_ (.A1(_0028_),
    .A2(_0220_),
    .Y(_0221_),
    .B1(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit8.Q ));
 sg13g2_nor2_1 _0782_ (.A(_0027_),
    .B(net636),
    .Y(_0222_));
 sg13g2_o21ai_1 _0783_ (.B1(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit7.Q ),
    .Y(_0223_),
    .A1(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit6.Q ),
    .A2(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.J_NS4_BEG12 ));
 sg13g2_mux2_1 _0784_ (.A0(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.J_NS4_BEG4 ),
    .A1(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.J_NS4_BEG8 ),
    .S(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit6.Q ),
    .X(_0224_));
 sg13g2_o21ai_1 _0785_ (.B1(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit8.Q ),
    .Y(_0225_),
    .A1(_0222_),
    .A2(_0223_));
 sg13g2_a21oi_1 _0786_ (.A1(_0028_),
    .A2(_0224_),
    .Y(_0226_),
    .B1(_0225_));
 sg13g2_a21oi_1 _0787_ (.A1(_0219_),
    .A2(_0221_),
    .Y(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.S4BEG0 ),
    .B1(_0226_));
 sg13g2_o21ai_1 _0788_ (.B1(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit10.Q ),
    .Y(_0227_),
    .A1(net169),
    .A2(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit9.Q ));
 sg13g2_inv_1 _0789_ (.Y(_0228_),
    .A(_0227_));
 sg13g2_o21ai_1 _0790_ (.B1(_0228_),
    .Y(_0229_),
    .A1(_0029_),
    .A2(_0160_));
 sg13g2_mux2_1 _0791_ (.A0(net143),
    .A1(net178),
    .S(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit9.Q ),
    .X(_0230_));
 sg13g2_a21oi_1 _0792_ (.A1(_0030_),
    .A2(_0230_),
    .Y(_0231_),
    .B1(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit11.Q ));
 sg13g2_nor2_1 _0793_ (.A(_0029_),
    .B(net634),
    .Y(_0232_));
 sg13g2_o21ai_1 _0794_ (.B1(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit10.Q ),
    .Y(_0233_),
    .A1(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit9.Q ),
    .A2(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.J_NS4_BEG13 ));
 sg13g2_mux2_1 _0795_ (.A0(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.J_NS4_BEG5 ),
    .A1(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.J_NS4_BEG9 ),
    .S(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit9.Q ),
    .X(_0234_));
 sg13g2_o21ai_1 _0796_ (.B1(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit11.Q ),
    .Y(_0235_),
    .A1(_0232_),
    .A2(_0233_));
 sg13g2_a21oi_1 _0797_ (.A1(_0030_),
    .A2(_0234_),
    .Y(_0236_),
    .B1(_0235_));
 sg13g2_a21oi_1 _0798_ (.A1(_0229_),
    .A2(_0231_),
    .Y(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.S4BEG1 ),
    .B1(_0236_));
 sg13g2_o21ai_1 _0799_ (.B1(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit13.Q ),
    .Y(_0237_),
    .A1(net170),
    .A2(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit12.Q ));
 sg13g2_inv_1 _0800_ (.Y(_0238_),
    .A(_0237_));
 sg13g2_o21ai_1 _0801_ (.B1(_0238_),
    .Y(_0239_),
    .A1(_0031_),
    .A2(_0159_));
 sg13g2_mux2_1 _0802_ (.A0(net144),
    .A1(net179),
    .S(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit12.Q ),
    .X(_0240_));
 sg13g2_a21oi_1 _0803_ (.A1(_0032_),
    .A2(_0240_),
    .Y(_0241_),
    .B1(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit14.Q ));
 sg13g2_nor2_1 _0804_ (.A(_0031_),
    .B(net633),
    .Y(_0242_));
 sg13g2_o21ai_1 _0805_ (.B1(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit13.Q ),
    .Y(_0243_),
    .A1(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit12.Q ),
    .A2(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.J_NS4_BEG14 ));
 sg13g2_mux2_1 _0806_ (.A0(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.J_NS4_BEG6 ),
    .A1(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.J_NS4_BEG10 ),
    .S(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit12.Q ),
    .X(_0244_));
 sg13g2_o21ai_1 _0807_ (.B1(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit14.Q ),
    .Y(_0245_),
    .A1(_0242_),
    .A2(_0243_));
 sg13g2_a21oi_1 _0808_ (.A1(_0032_),
    .A2(_0244_),
    .Y(_0246_),
    .B1(_0245_));
 sg13g2_a21oi_1 _0809_ (.A1(_0239_),
    .A2(_0241_),
    .Y(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.S4BEG2 ),
    .B1(_0246_));
 sg13g2_o21ai_1 _0810_ (.B1(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit16.Q ),
    .Y(_0247_),
    .A1(net171),
    .A2(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit15.Q ));
 sg13g2_inv_1 _0811_ (.Y(_0248_),
    .A(_0247_));
 sg13g2_o21ai_1 _0812_ (.B1(_0248_),
    .Y(_0249_),
    .A1(_0033_),
    .A2(_0158_));
 sg13g2_mux2_1 _0813_ (.A0(net145),
    .A1(net180),
    .S(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit15.Q ),
    .X(_0250_));
 sg13g2_a21oi_1 _0814_ (.A1(_0034_),
    .A2(_0250_),
    .Y(_0251_),
    .B1(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit17.Q ));
 sg13g2_nor2_1 _0815_ (.A(_0033_),
    .B(_0084_),
    .Y(_0252_));
 sg13g2_o21ai_1 _0816_ (.B1(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit16.Q ),
    .Y(_0253_),
    .A1(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit15.Q ),
    .A2(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.J_NS4_BEG15 ));
 sg13g2_mux2_1 _0817_ (.A0(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.J_NS4_BEG7 ),
    .A1(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.J_NS4_BEG11 ),
    .S(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit15.Q ),
    .X(_0254_));
 sg13g2_o21ai_1 _0818_ (.B1(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit17.Q ),
    .Y(_0255_),
    .A1(_0252_),
    .A2(_0253_));
 sg13g2_a21oi_1 _0819_ (.A1(_0034_),
    .A2(_0254_),
    .Y(_0256_),
    .B1(_0255_));
 sg13g2_a21oi_1 _0820_ (.A1(_0249_),
    .A2(_0251_),
    .Y(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.S4BEG3 ),
    .B1(_0256_));
 sg13g2_nor2b_1 _0821_ (.A(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit2.Q ),
    .B_N(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit1.Q ),
    .Y(_0257_));
 sg13g2_nand2b_1 _0822_ (.Y(_0258_),
    .B(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit2.Q ),
    .A_N(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit1.Q ));
 sg13g2_nand2_1 _0823_ (.Y(_0259_),
    .A(net229),
    .B(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit0.Q ));
 sg13g2_or2_1 _0824_ (.X(_0260_),
    .B(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit2.Q ),
    .A(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit1.Q ));
 sg13g2_a21oi_1 _0825_ (.A1(net241),
    .A2(_0035_),
    .Y(_0261_),
    .B1(_0260_));
 sg13g2_nand2_1 _0826_ (.Y(_0262_),
    .A(net147),
    .B(_0035_));
 sg13g2_nand2_1 _0827_ (.Y(_0263_),
    .A(net148),
    .B(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit0.Q ));
 sg13g2_nand4_1 _0828_ (.B(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit2.Q ),
    .C(_0262_),
    .A(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit1.Q ),
    .Y(_0264_),
    .D(_0263_));
 sg13g2_a21oi_1 _0829_ (.A1(net160),
    .A2(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit0.Q ),
    .Y(_0265_),
    .B1(_0258_));
 sg13g2_o21ai_1 _0830_ (.B1(_0265_),
    .Y(_0266_),
    .A1(_0000_),
    .A2(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit0.Q ));
 sg13g2_and2_1 _0831_ (.A(net154),
    .B(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit0.Q ),
    .X(_0267_));
 sg13g2_a21oi_1 _0832_ (.A1(net230),
    .A2(_0035_),
    .Y(_0268_),
    .B1(_0267_));
 sg13g2_a22oi_1 _0833_ (.Y(_0269_),
    .B1(_0268_),
    .B2(_0257_),
    .A2(_0261_),
    .A1(_0259_));
 sg13g2_nand3_1 _0834_ (.B(_0266_),
    .C(_0269_),
    .A(_0264_),
    .Y(_0270_));
 sg13g2_nand2b_1 _0835_ (.Y(_0271_),
    .B(_0257_),
    .A_N(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.S2BEG0 ));
 sg13g2_or3_1 _0836_ (.A(net150),
    .B(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit1.Q ),
    .C(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit2.Q ),
    .X(_0272_));
 sg13g2_or2_1 _0837_ (.X(_0273_),
    .B(_0258_),
    .A(net129));
 sg13g2_nand4_1 _0838_ (.B(_0271_),
    .C(_0272_),
    .A(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit0.Q ),
    .Y(_0274_),
    .D(_0273_));
 sg13g2_nand2b_1 _0839_ (.Y(_0275_),
    .B(net151),
    .A_N(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit2.Q ));
 sg13g2_nor3_1 _0840_ (.A(net149),
    .B(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit1.Q ),
    .C(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit2.Q ),
    .Y(_0276_));
 sg13g2_a221oi_1 _0841_ (.B2(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit1.Q ),
    .C1(_0276_),
    .B1(_0275_),
    .A1(_0002_),
    .Y(_0277_),
    .A2(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit2.Q ));
 sg13g2_a21oi_1 _0842_ (.A1(_0035_),
    .A2(_0277_),
    .Y(_0278_),
    .B1(_0036_));
 sg13g2_a22oi_1 _0843_ (.Y(net327),
    .B1(_0274_),
    .B2(_0278_),
    .A2(_0270_),
    .A1(_0036_));
 sg13g2_mux4_1 _0844_ (.S0(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit4.Q ),
    .A0(net230),
    .A1(net154),
    .A2(net147),
    .A3(net148),
    .S1(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit6.Q ),
    .X(_0279_));
 sg13g2_nand2_1 _0845_ (.Y(_0280_),
    .A(net229),
    .B(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit4.Q ));
 sg13g2_nor2b_1 _0846_ (.A(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit4.Q ),
    .B_N(net241),
    .Y(_0281_));
 sg13g2_nor3_1 _0847_ (.A(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit5.Q ),
    .B(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit6.Q ),
    .C(_0281_),
    .Y(_0282_));
 sg13g2_nand2_1 _0848_ (.Y(_0283_),
    .A(_0037_),
    .B(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit6.Q ));
 sg13g2_nand2b_1 _0849_ (.Y(_0284_),
    .B(net157),
    .A_N(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit4.Q ));
 sg13g2_a21oi_1 _0850_ (.A1(net160),
    .A2(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit4.Q ),
    .Y(_0285_),
    .B1(_0283_));
 sg13g2_a22oi_1 _0851_ (.Y(_0286_),
    .B1(_0284_),
    .B2(_0285_),
    .A2(_0282_),
    .A1(_0280_));
 sg13g2_o21ai_1 _0852_ (.B1(_0286_),
    .Y(_0287_),
    .A1(_0037_),
    .A2(_0279_));
 sg13g2_nor3_1 _0853_ (.A(_0037_),
    .B(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit6.Q ),
    .C(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.S2BEG0 ),
    .Y(_0288_));
 sg13g2_nor3_1 _0854_ (.A(net150),
    .B(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit5.Q ),
    .C(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit6.Q ),
    .Y(_0289_));
 sg13g2_o21ai_1 _0855_ (.B1(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit4.Q ),
    .Y(_0290_),
    .A1(net129),
    .A2(_0283_));
 sg13g2_nor3_1 _0856_ (.A(_0288_),
    .B(_0289_),
    .C(_0290_),
    .Y(_0291_));
 sg13g2_a21oi_1 _0857_ (.A1(_0001_),
    .A2(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit5.Q ),
    .Y(_0292_),
    .B1(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit6.Q ));
 sg13g2_a21oi_1 _0858_ (.A1(net128),
    .A2(_0037_),
    .Y(_0293_),
    .B1(_0292_));
 sg13g2_nor3_1 _0859_ (.A(net149),
    .B(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit5.Q ),
    .C(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit6.Q ),
    .Y(_0294_));
 sg13g2_nor3_1 _0860_ (.A(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit4.Q ),
    .B(_0293_),
    .C(_0294_),
    .Y(_0295_));
 sg13g2_o21ai_1 _0861_ (.B1(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit7.Q ),
    .Y(_0296_),
    .A1(_0291_),
    .A2(_0295_));
 sg13g2_o21ai_1 _0862_ (.B1(_0296_),
    .Y(net581),
    .A1(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit7.Q ),
    .A2(_0287_));
 sg13g2_dlhq_1 _0863_ (.D(net106),
    .GATE(net745),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame0_bit31.Q ));
 sg13g2_dlhq_1 _0864_ (.D(net790),
    .GATE(net745),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame0_bit30.Q ));
 sg13g2_dlhq_1 _0865_ (.D(net792),
    .GATE(net745),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame0_bit29.Q ));
 sg13g2_dlhq_1 _0866_ (.D(net793),
    .GATE(net746),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame0_bit28.Q ));
 sg13g2_dlhq_1 _0867_ (.D(net794),
    .GATE(net747),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame0_bit27.Q ));
 sg13g2_dlhq_1 _0868_ (.D(net795),
    .GATE(net744),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame0_bit26.Q ));
 sg13g2_dlhq_1 _0869_ (.D(net796),
    .GATE(net748),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame0_bit25.Q ));
 sg13g2_dlhq_1 _0870_ (.D(net797),
    .GATE(net748),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame0_bit24.Q ));
 sg13g2_dlhq_1 _0871_ (.D(net798),
    .GATE(net743),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame0_bit23.Q ));
 sg13g2_dlhq_1 _0872_ (.D(net799),
    .GATE(net743),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame0_bit22.Q ));
 sg13g2_dlhq_1 _0873_ (.D(net800),
    .GATE(net744),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame0_bit21.Q ));
 sg13g2_dlhq_1 _0874_ (.D(net801),
    .GATE(net744),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame0_bit20.Q ));
 sg13g2_dlhq_1 _0875_ (.D(net803),
    .GATE(net743),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame0_bit19.Q ));
 sg13g2_dlhq_1 _0876_ (.D(net804),
    .GATE(net743),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame0_bit18.Q ));
 sg13g2_dlhq_1 _0877_ (.D(net805),
    .GATE(net744),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame0_bit17.Q ));
 sg13g2_dlhq_1 _0878_ (.D(net806),
    .GATE(net744),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame0_bit16.Q ));
 sg13g2_dlhq_1 _0879_ (.D(net88),
    .GATE(net744),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame0_bit15.Q ));
 sg13g2_dlhq_1 _0880_ (.D(net87),
    .GATE(net744),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame0_bit14.Q ));
 sg13g2_dlhq_1 _0881_ (.D(net809),
    .GATE(net745),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame0_bit13.Q ));
 sg13g2_dlhq_1 _0882_ (.D(net810),
    .GATE(net745),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame0_bit12.Q ));
 sg13g2_dlhq_1 _0883_ (.D(net811),
    .GATE(net745),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame0_bit11.Q ));
 sg13g2_dlhq_1 _0884_ (.D(net812),
    .GATE(net745),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame0_bit10.Q ));
 sg13g2_dlhq_1 _0885_ (.D(net782),
    .GATE(net743),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame0_bit9.Q ));
 sg13g2_dlhq_1 _0886_ (.D(net783),
    .GATE(net743),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame0_bit8.Q ));
 sg13g2_dlhq_1 _0887_ (.D(net111),
    .GATE(net746),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame0_bit7.Q ));
 sg13g2_dlhq_1 _0888_ (.D(net110),
    .GATE(net745),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame0_bit6.Q ));
 sg13g2_dlhq_1 _0889_ (.D(net109),
    .GATE(net746),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame0_bit5.Q ));
 sg13g2_dlhq_1 _0890_ (.D(net787),
    .GATE(net746),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame0_bit4.Q ));
 sg13g2_dlhq_1 _0891_ (.D(net788),
    .GATE(net747),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame0_bit3.Q ));
 sg13g2_dlhq_1 _0892_ (.D(net791),
    .GATE(net744),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame0_bit2.Q ));
 sg13g2_dlhq_1 _0893_ (.D(net802),
    .GATE(net743),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame0_bit1.Q ));
 sg13g2_dlhq_1 _0894_ (.D(net813),
    .GATE(net743),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame0_bit0.Q ));
 sg13g2_dlhq_1 _0895_ (.D(net106),
    .GATE(net734),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame1_bit31.Q ));
 sg13g2_dlhq_1 _0896_ (.D(net105),
    .GATE(net734),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame1_bit30.Q ));
 sg13g2_dlhq_1 _0897_ (.D(net103),
    .GATE(net735),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame1_bit29.Q ));
 sg13g2_dlhq_1 _0898_ (.D(net102),
    .GATE(net735),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame1_bit28.Q ));
 sg13g2_dlhq_1 _0899_ (.D(net794),
    .GATE(net733),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame1_bit27.Q ));
 sg13g2_dlhq_1 _0900_ (.D(net795),
    .GATE(net732),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame1_bit26.Q ));
 sg13g2_dlhq_1 _0901_ (.D(net796),
    .GATE(net731),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame1_bit25.Q ));
 sg13g2_dlhq_1 _0902_ (.D(net797),
    .GATE(net731),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame1_bit24.Q ));
 sg13g2_dlhq_1 _0903_ (.D(net97),
    .GATE(net734),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame1_bit23.Q ));
 sg13g2_dlhq_1 _0904_ (.D(net96),
    .GATE(net734),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame1_bit22.Q ));
 sg13g2_dlhq_1 _0905_ (.D(net95),
    .GATE(net734),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame1_bit21.Q ));
 sg13g2_dlhq_1 _0906_ (.D(net94),
    .GATE(net735),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame1_bit20.Q ));
 sg13g2_dlhq_1 _0907_ (.D(net92),
    .GATE(net733),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame1_bit19.Q ));
 sg13g2_dlhq_1 _0908_ (.D(net91),
    .GATE(net732),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame1_bit18.Q ));
 sg13g2_dlhq_1 _0909_ (.D(net805),
    .GATE(net731),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame1_bit17.Q ));
 sg13g2_dlhq_1 _0910_ (.D(net806),
    .GATE(net737),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame1_bit16.Q ));
 sg13g2_dlhq_1 _0911_ (.D(net88),
    .GATE(net734),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame1_bit15.Q ));
 sg13g2_dlhq_1 _0912_ (.D(net87),
    .GATE(net734),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame1_bit14.Q ));
 sg13g2_dlhq_1 _0913_ (.D(net809),
    .GATE(net735),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame1_bit13.Q ));
 sg13g2_dlhq_1 _0914_ (.D(net810),
    .GATE(net735),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame1_bit12.Q ));
 sg13g2_dlhq_1 _0915_ (.D(net811),
    .GATE(net732),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame1_bit11.Q ));
 sg13g2_dlhq_1 _0916_ (.D(net812),
    .GATE(net732),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame1_bit10.Q ));
 sg13g2_dlhq_1 _0917_ (.D(net782),
    .GATE(net731),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame1_bit9.Q ));
 sg13g2_dlhq_1 _0918_ (.D(net783),
    .GATE(net731),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame1_bit8.Q ));
 sg13g2_dlhq_1 _0919_ (.D(net784),
    .GATE(net732),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame1_bit7.Q ));
 sg13g2_dlhq_1 _0920_ (.D(net110),
    .GATE(net732),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame1_bit6.Q ));
 sg13g2_dlhq_1 _0921_ (.D(net786),
    .GATE(net731),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame1_bit5.Q ));
 sg13g2_dlhq_1 _0922_ (.D(net787),
    .GATE(net731),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame1_bit4.Q ));
 sg13g2_dlhq_1 _0923_ (.D(net107),
    .GATE(net733),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame1_bit3.Q ));
 sg13g2_dlhq_1 _0924_ (.D(net104),
    .GATE(net733),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame1_bit2.Q ));
 sg13g2_dlhq_1 _0925_ (.D(net93),
    .GATE(net732),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame1_bit1.Q ));
 sg13g2_dlhq_1 _0926_ (.D(net82),
    .GATE(net732),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame1_bit0.Q ));
 sg13g2_dlhq_1 _0927_ (.D(net789),
    .GATE(net722),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame2_bit31.Q ));
 sg13g2_dlhq_1 _0928_ (.D(net790),
    .GATE(net722),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame2_bit30.Q ));
 sg13g2_dlhq_1 _0929_ (.D(net792),
    .GATE(net720),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame2_bit29.Q ));
 sg13g2_dlhq_1 _0930_ (.D(net793),
    .GATE(net720),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame2_bit28.Q ));
 sg13g2_dlhq_1 _0931_ (.D(net101),
    .GATE(net722),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame2_bit27.Q ));
 sg13g2_dlhq_1 _0932_ (.D(net100),
    .GATE(net722),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame2_bit26.Q ));
 sg13g2_dlhq_1 _0933_ (.D(net796),
    .GATE(net723),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame2_bit25.Q ));
 sg13g2_dlhq_1 _0934_ (.D(net797),
    .GATE(net723),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame2_bit24.Q ));
 sg13g2_dlhq_1 _0935_ (.D(net798),
    .GATE(net723),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame2_bit23.Q ));
 sg13g2_dlhq_1 _0936_ (.D(net799),
    .GATE(net723),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame2_bit22.Q ));
 sg13g2_dlhq_1 _0937_ (.D(net95),
    .GATE(net720),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame2_bit21.Q ));
 sg13g2_dlhq_1 _0938_ (.D(net94),
    .GATE(net720),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame2_bit20.Q ));
 sg13g2_dlhq_1 _0939_ (.D(net803),
    .GATE(net721),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame2_bit19.Q ));
 sg13g2_dlhq_1 _0940_ (.D(net804),
    .GATE(net721),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame2_bit18.Q ));
 sg13g2_dlhq_1 _0941_ (.D(net805),
    .GATE(net721),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame2_bit17.Q ));
 sg13g2_dlhq_1 _0942_ (.D(net806),
    .GATE(net721),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame2_bit16.Q ));
 sg13g2_dlhq_1 _0943_ (.D(net807),
    .GATE(net723),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame2_bit15.Q ));
 sg13g2_dlhq_1 _0944_ (.D(net808),
    .GATE(net723),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame2_bit14.Q ));
 sg13g2_dlhq_1 _0945_ (.D(net86),
    .GATE(net720),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame2_bit13.Q ));
 sg13g2_dlhq_1 _0946_ (.D(net85),
    .GATE(net720),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame2_bit12.Q ));
 sg13g2_dlhq_1 _0947_ (.D(net84),
    .GATE(net722),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame2_bit11.Q ));
 sg13g2_dlhq_1 _0948_ (.D(net83),
    .GATE(net722),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame2_bit10.Q ));
 sg13g2_dlhq_1 _0949_ (.D(net782),
    .GATE(net719),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame2_bit9.Q ));
 sg13g2_dlhq_1 _0950_ (.D(net783),
    .GATE(net719),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame2_bit8.Q ));
 sg13g2_dlhq_1 _0951_ (.D(net784),
    .GATE(net723),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame2_bit7.Q ));
 sg13g2_dlhq_1 _0952_ (.D(net785),
    .GATE(net723),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame2_bit6.Q ));
 sg13g2_dlhq_1 _0953_ (.D(net109),
    .GATE(net720),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame2_bit5.Q ));
 sg13g2_dlhq_1 _0954_ (.D(net108),
    .GATE(net720),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame2_bit4.Q ));
 sg13g2_dlhq_1 _0955_ (.D(net107),
    .GATE(net721),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame2_bit3.Q ));
 sg13g2_dlhq_1 _0956_ (.D(net104),
    .GATE(net721),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame2_bit2.Q ));
 sg13g2_dlhq_1 _0957_ (.D(net802),
    .GATE(net722),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame2_bit1.Q ));
 sg13g2_dlhq_1 _0958_ (.D(net813),
    .GATE(net722),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame2_bit0.Q ));
 sg13g2_dlhq_1 _0959_ (.D(net789),
    .GATE(net709),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame3_bit31.Q ));
 sg13g2_dlhq_1 _0960_ (.D(net790),
    .GATE(net709),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame3_bit30.Q ));
 sg13g2_dlhq_1 _0961_ (.D(net103),
    .GATE(net712),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame3_bit29.Q ));
 sg13g2_dlhq_1 _0962_ (.D(net102),
    .GATE(net712),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame3_bit28.Q ));
 sg13g2_dlhq_1 _0963_ (.D(net101),
    .GATE(net712),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame3_bit27.Q ));
 sg13g2_dlhq_1 _0964_ (.D(net100),
    .GATE(net712),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame3_bit26.Q ));
 sg13g2_dlhq_1 _0965_ (.D(net796),
    .GATE(net709),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame3_bit25.Q ));
 sg13g2_dlhq_1 _0966_ (.D(net797),
    .GATE(net709),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame3_bit24.Q ));
 sg13g2_dlhq_1 _0967_ (.D(net798),
    .GATE(net709),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame3_bit23.Q ));
 sg13g2_dlhq_1 _0968_ (.D(net799),
    .GATE(net709),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame3_bit22.Q ));
 sg13g2_dlhq_1 _0969_ (.D(net800),
    .GATE(net710),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame3_bit21.Q ));
 sg13g2_dlhq_1 _0970_ (.D(net801),
    .GATE(net710),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame3_bit20.Q ));
 sg13g2_dlhq_1 _0971_ (.D(net803),
    .GATE(net711),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame3_bit19.Q ));
 sg13g2_dlhq_1 _0972_ (.D(net804),
    .GATE(net711),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame3_bit18.Q ));
 sg13g2_dlhq_1 _0973_ (.D(net805),
    .GATE(net711),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame3_bit17.Q ));
 sg13g2_dlhq_1 _0974_ (.D(net806),
    .GATE(net711),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame3_bit16.Q ));
 sg13g2_dlhq_1 _0975_ (.D(net807),
    .GATE(net713),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame3_bit15.Q ));
 sg13g2_dlhq_1 _0976_ (.D(net808),
    .GATE(net713),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame3_bit14.Q ));
 sg13g2_dlhq_1 _0977_ (.D(net86),
    .GATE(net710),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame3_bit13.Q ));
 sg13g2_dlhq_1 _0978_ (.D(net85),
    .GATE(net710),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame3_bit12.Q ));
 sg13g2_dlhq_1 _0979_ (.D(net84),
    .GATE(net712),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame3_bit11.Q ));
 sg13g2_dlhq_1 _0980_ (.D(net83),
    .GATE(net712),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame3_bit10.Q ));
 sg13g2_dlhq_1 _0981_ (.D(net782),
    .GATE(net708),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame3_bit9.Q ));
 sg13g2_dlhq_1 _0982_ (.D(net783),
    .GATE(net708),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame3_bit8.Q ));
 sg13g2_dlhq_1 _0983_ (.D(net784),
    .GATE(net709),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame3_bit7.Q ));
 sg13g2_dlhq_1 _0984_ (.D(net785),
    .GATE(net709),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame3_bit6.Q ));
 sg13g2_dlhq_1 _0985_ (.D(net786),
    .GATE(net710),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame3_bit5.Q ));
 sg13g2_dlhq_1 _0986_ (.D(net108),
    .GATE(net710),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame3_bit4.Q ));
 sg13g2_dlhq_1 _0987_ (.D(net788),
    .GATE(net711),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame3_bit3.Q ));
 sg13g2_dlhq_1 _0988_ (.D(net791),
    .GATE(net710),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame3_bit2.Q ));
 sg13g2_dlhq_1 _0989_ (.D(net802),
    .GATE(net712),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame3_bit1.Q ));
 sg13g2_dlhq_1 _0990_ (.D(net813),
    .GATE(net712),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame3_bit0.Q ));
 sg13g2_dlhq_1 _0991_ (.D(net789),
    .GATE(net698),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame4_bit31.Q ));
 sg13g2_dlhq_1 _0992_ (.D(net790),
    .GATE(net698),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame4_bit30.Q ));
 sg13g2_dlhq_1 _0993_ (.D(net792),
    .GATE(net699),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame4_bit29.Q ));
 sg13g2_dlhq_1 _0994_ (.D(net793),
    .GATE(net697),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame4_bit28.Q ));
 sg13g2_dlhq_1 _0995_ (.D(net794),
    .GATE(net698),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame4_bit27.Q ));
 sg13g2_dlhq_1 _0996_ (.D(net795),
    .GATE(net698),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame4_bit26.Q ));
 sg13g2_dlhq_1 _0997_ (.D(net796),
    .GATE(net700),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame4_bit25.Q ));
 sg13g2_dlhq_1 _0998_ (.D(net797),
    .GATE(net701),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame4_bit24.Q ));
 sg13g2_dlhq_1 _0999_ (.D(net798),
    .GATE(net700),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame4_bit23.Q ));
 sg13g2_dlhq_1 _1000_ (.D(net799),
    .GATE(net700),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame4_bit22.Q ));
 sg13g2_dlhq_1 _1001_ (.D(net800),
    .GATE(net697),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame4_bit21.Q ));
 sg13g2_dlhq_1 _1002_ (.D(net801),
    .GATE(net697),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame4_bit20.Q ));
 sg13g2_dlhq_1 _1003_ (.D(net803),
    .GATE(net698),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame4_bit19.Q ));
 sg13g2_dlhq_1 _1004_ (.D(net804),
    .GATE(net698),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame4_bit18.Q ));
 sg13g2_dlhq_1 _1005_ (.D(net805),
    .GATE(net698),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame4_bit17.Q ));
 sg13g2_dlhq_1 _1006_ (.D(net806),
    .GATE(net698),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame4_bit16.Q ));
 sg13g2_dlhq_1 _1007_ (.D(net807),
    .GATE(net700),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame4_bit15.Q ));
 sg13g2_dlhq_1 _1008_ (.D(net808),
    .GATE(net700),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame4_bit14.Q ));
 sg13g2_dlhq_1 _1009_ (.D(net809),
    .GATE(net697),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame4_bit13.Q ));
 sg13g2_dlhq_1 _1010_ (.D(net810),
    .GATE(net697),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame4_bit12.Q ));
 sg13g2_dlhq_1 _1011_ (.D(net811),
    .GATE(net701),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame4_bit11.Q ));
 sg13g2_dlhq_1 _1012_ (.D(net812),
    .GATE(net701),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame4_bit10.Q ));
 sg13g2_dlhq_1 _1013_ (.D(net782),
    .GATE(net700),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame4_bit9.Q ));
 sg13g2_dlhq_1 _1014_ (.D(net783),
    .GATE(net700),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame4_bit8.Q ));
 sg13g2_dlhq_1 _1015_ (.D(net784),
    .GATE(net700),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame4_bit7.Q ));
 sg13g2_dlhq_1 _1016_ (.D(net785),
    .GATE(net697),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame4_bit6.Q ));
 sg13g2_dlhq_1 _1017_ (.D(net786),
    .GATE(net697),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame4_bit5.Q ));
 sg13g2_dlhq_1 _1018_ (.D(net787),
    .GATE(net697),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame4_bit4.Q ));
 sg13g2_dlhq_1 _1019_ (.D(net788),
    .GATE(net702),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame4_bit3.Q ));
 sg13g2_dlhq_1 _1020_ (.D(net791),
    .GATE(net702),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame4_bit2.Q ));
 sg13g2_dlhq_1 _1021_ (.D(net802),
    .GATE(net699),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame4_bit1.Q ));
 sg13g2_dlhq_1 _1022_ (.D(net813),
    .GATE(net699),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame4_bit0.Q ));
 sg13g2_dlhq_1 _1023_ (.D(net789),
    .GATE(net685),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame5_bit31.Q ));
 sg13g2_dlhq_1 _1024_ (.D(net790),
    .GATE(net685),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame5_bit30.Q ));
 sg13g2_dlhq_1 _1025_ (.D(net792),
    .GATE(net685),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame5_bit29.Q ));
 sg13g2_dlhq_1 _1026_ (.D(net793),
    .GATE(net685),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame5_bit28.Q ));
 sg13g2_dlhq_1 _1027_ (.D(net794),
    .GATE(net687),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame5_bit27.Q ));
 sg13g2_dlhq_1 _1028_ (.D(net795),
    .GATE(net687),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame5_bit26.Q ));
 sg13g2_dlhq_1 _1029_ (.D(net796),
    .GATE(net688),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame5_bit25.Q ));
 sg13g2_dlhq_1 _1030_ (.D(net797),
    .GATE(net688),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame5_bit24.Q ));
 sg13g2_dlhq_1 _1031_ (.D(net798),
    .GATE(net685),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame5_bit23.Q ));
 sg13g2_dlhq_1 _1032_ (.D(net799),
    .GATE(net686),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame5_bit22.Q ));
 sg13g2_dlhq_1 _1033_ (.D(net800),
    .GATE(net686),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame5_bit21.Q ));
 sg13g2_dlhq_1 _1034_ (.D(net801),
    .GATE(net686),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame5_bit20.Q ));
 sg13g2_dlhq_1 _1035_ (.D(net803),
    .GATE(net687),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame5_bit19.Q ));
 sg13g2_dlhq_1 _1036_ (.D(net804),
    .GATE(net687),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame5_bit18.Q ));
 sg13g2_dlhq_1 _1037_ (.D(net90),
    .GATE(net688),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame5_bit17.Q ));
 sg13g2_dlhq_1 _1038_ (.D(net89),
    .GATE(net687),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame5_bit16.Q ));
 sg13g2_dlhq_1 _1039_ (.D(net807),
    .GATE(net685),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame5_bit15.Q ));
 sg13g2_dlhq_1 _1040_ (.D(net808),
    .GATE(net685),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame5_bit14.Q ));
 sg13g2_dlhq_1 _1041_ (.D(net809),
    .GATE(net686),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame5_bit13.Q ));
 sg13g2_dlhq_1 _1042_ (.D(net810),
    .GATE(net686),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame5_bit12.Q ));
 sg13g2_dlhq_1 _1043_ (.D(net811),
    .GATE(net687),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame5_bit11.Q ));
 sg13g2_dlhq_1 _1044_ (.D(net812),
    .GATE(net687),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame5_bit10.Q ));
 sg13g2_dlhq_1 _1045_ (.D(net113),
    .GATE(net688),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame5_bit9.Q ));
 sg13g2_dlhq_1 _1046_ (.D(net112),
    .GATE(net688),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame5_bit8.Q ));
 sg13g2_dlhq_1 _1047_ (.D(net784),
    .GATE(net686),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame5_bit7.Q ));
 sg13g2_dlhq_1 _1048_ (.D(net785),
    .GATE(net685),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame5_bit6.Q ));
 sg13g2_dlhq_1 _1049_ (.D(net786),
    .GATE(net686),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame5_bit5.Q ));
 sg13g2_dlhq_1 _1050_ (.D(net787),
    .GATE(net686),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame5_bit4.Q ));
 sg13g2_dlhq_1 _1051_ (.D(net788),
    .GATE(net690),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame5_bit3.Q ));
 sg13g2_dlhq_1 _1052_ (.D(net791),
    .GATE(net690),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame5_bit2.Q ));
 sg13g2_dlhq_1 _1053_ (.D(net802),
    .GATE(net690),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame5_bit1.Q ));
 sg13g2_dlhq_1 _1054_ (.D(net813),
    .GATE(net690),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame5_bit0.Q ));
 sg13g2_dlhq_1 _1055_ (.D(net789),
    .GATE(net675),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame6_bit31.Q ));
 sg13g2_dlhq_1 _1056_ (.D(net790),
    .GATE(net675),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame6_bit30.Q ));
 sg13g2_dlhq_1 _1057_ (.D(net792),
    .GATE(net678),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame6_bit29.Q ));
 sg13g2_dlhq_1 _1058_ (.D(net793),
    .GATE(net678),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame6_bit28.Q ));
 sg13g2_dlhq_1 _1059_ (.D(net794),
    .GATE(net677),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame6_bit27.Q ));
 sg13g2_dlhq_1 _1060_ (.D(net795),
    .GATE(net677),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame6_bit26.Q ));
 sg13g2_dlhq_1 _1061_ (.D(net796),
    .GATE(net675),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame6_bit25.Q ));
 sg13g2_dlhq_1 _1062_ (.D(net797),
    .GATE(net675),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame6_bit24.Q ));
 sg13g2_dlhq_1 _1063_ (.D(net798),
    .GATE(net675),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame6_bit23.Q ));
 sg13g2_dlhq_1 _1064_ (.D(net799),
    .GATE(net675),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame6_bit22.Q ));
 sg13g2_dlhq_1 _1065_ (.D(net800),
    .GATE(net676),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame6_bit21.Q ));
 sg13g2_dlhq_1 _1066_ (.D(net801),
    .GATE(net676),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame6_bit20.Q ));
 sg13g2_dlhq_1 _1067_ (.D(net803),
    .GATE(net679),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame6_bit19.Q ));
 sg13g2_dlhq_1 _1068_ (.D(net804),
    .GATE(net679),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame6_bit18.Q ));
 sg13g2_dlhq_1 _1069_ (.D(net90),
    .GATE(net678),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame6_bit17.Q ));
 sg13g2_dlhq_1 _1070_ (.D(net89),
    .GATE(net678),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame6_bit16.Q ));
 sg13g2_dlhq_1 _1071_ (.D(net807),
    .GATE(net678),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame6_bit15.Q ));
 sg13g2_dlhq_1 _1072_ (.D(net808),
    .GATE(net678),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame6_bit14.Q ));
 sg13g2_dlhq_1 _1073_ (.D(net809),
    .GATE(net675),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame6_bit13.Q ));
 sg13g2_dlhq_1 _1074_ (.D(net810),
    .GATE(net676),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame6_bit12.Q ));
 sg13g2_dlhq_1 _1075_ (.D(net811),
    .GATE(net677),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame6_bit11.Q ));
 sg13g2_dlhq_1 _1076_ (.D(net812),
    .GATE(net677),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame6_bit10.Q ));
 sg13g2_dlhq_1 _1077_ (.D(net782),
    .GATE(net679),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame6_bit9.Q ));
 sg13g2_dlhq_1 _1078_ (.D(net783),
    .GATE(net679),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame6_bit8.Q ));
 sg13g2_dlhq_1 _1079_ (.D(net784),
    .GATE(net676),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame6_bit7.Q ));
 sg13g2_dlhq_1 _1080_ (.D(net785),
    .GATE(net676),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame6_bit6.Q ));
 sg13g2_dlhq_1 _1081_ (.D(net786),
    .GATE(net675),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame6_bit5.Q ));
 sg13g2_dlhq_1 _1082_ (.D(net787),
    .GATE(net677),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame6_bit4.Q ));
 sg13g2_dlhq_1 _1083_ (.D(net788),
    .GATE(net679),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame6_bit3.Q ));
 sg13g2_dlhq_1 _1084_ (.D(net791),
    .GATE(net679),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame6_bit2.Q ));
 sg13g2_dlhq_1 _1085_ (.D(net802),
    .GATE(net679),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame6_bit1.Q ));
 sg13g2_dlhq_1 _1086_ (.D(net813),
    .GATE(net679),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame6_bit0.Q ));
 sg13g2_dlhq_1 _1087_ (.D(net789),
    .GATE(net667),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit31.Q ));
 sg13g2_dlhq_1 _1088_ (.D(net790),
    .GATE(net667),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit30.Q ));
 sg13g2_dlhq_1 _1089_ (.D(net792),
    .GATE(net664),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit29.Q ));
 sg13g2_dlhq_1 _1090_ (.D(net793),
    .GATE(net664),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit28.Q ));
 sg13g2_dlhq_1 _1091_ (.D(net794),
    .GATE(net664),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit27.Q ));
 sg13g2_dlhq_1 _1092_ (.D(net100),
    .GATE(net665),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit26.Q ));
 sg13g2_dlhq_1 _1093_ (.D(net99),
    .GATE(net665),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit25.Q ));
 sg13g2_dlhq_1 _1094_ (.D(net98),
    .GATE(net665),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit24.Q ));
 sg13g2_dlhq_1 _1095_ (.D(net798),
    .GATE(net663),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit23.Q ));
 sg13g2_dlhq_1 _1096_ (.D(net799),
    .GATE(net663),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit22.Q ));
 sg13g2_dlhq_1 _1097_ (.D(net800),
    .GATE(net663),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit21.Q ));
 sg13g2_dlhq_1 _1098_ (.D(net801),
    .GATE(net663),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit20.Q ));
 sg13g2_dlhq_1 _1099_ (.D(net803),
    .GATE(net663),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit19.Q ));
 sg13g2_dlhq_1 _1100_ (.D(net804),
    .GATE(net663),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit18.Q ));
 sg13g2_dlhq_1 _1101_ (.D(net805),
    .GATE(net664),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit17.Q ));
 sg13g2_dlhq_1 _1102_ (.D(net806),
    .GATE(net664),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit16.Q ));
 sg13g2_dlhq_1 _1103_ (.D(net807),
    .GATE(net664),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit15.Q ));
 sg13g2_dlhq_1 _1104_ (.D(net808),
    .GATE(net664),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit14.Q ));
 sg13g2_dlhq_1 _1105_ (.D(net809),
    .GATE(net665),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit13.Q ));
 sg13g2_dlhq_1 _1106_ (.D(net810),
    .GATE(net665),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit12.Q ));
 sg13g2_dlhq_1 _1107_ (.D(net811),
    .GATE(net663),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit11.Q ));
 sg13g2_dlhq_1 _1108_ (.D(net812),
    .GATE(net663),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit10.Q ));
 sg13g2_dlhq_1 _1109_ (.D(net782),
    .GATE(net666),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit9.Q ));
 sg13g2_dlhq_1 _1110_ (.D(net112),
    .GATE(net666),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit8.Q ));
 sg13g2_dlhq_1 _1111_ (.D(net111),
    .GATE(net666),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit7.Q ));
 sg13g2_dlhq_1 _1112_ (.D(net785),
    .GATE(net666),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit6.Q ));
 sg13g2_dlhq_1 _1113_ (.D(net786),
    .GATE(net666),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit5.Q ));
 sg13g2_dlhq_1 _1114_ (.D(net787),
    .GATE(net666),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit4.Q ));
 sg13g2_dlhq_1 _1115_ (.D(net788),
    .GATE(net665),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit3.Q ));
 sg13g2_dlhq_1 _1116_ (.D(net791),
    .GATE(net664),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit2.Q ));
 sg13g2_dlhq_1 _1117_ (.D(net802),
    .GATE(net666),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit1.Q ));
 sg13g2_dlhq_1 _1118_ (.D(net813),
    .GATE(net666),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit0.Q ));
 sg13g2_dlhq_1 _1119_ (.D(net789),
    .GATE(net655),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit31.Q ));
 sg13g2_dlhq_1 _1120_ (.D(net105),
    .GATE(net655),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit30.Q ));
 sg13g2_dlhq_1 _1121_ (.D(net792),
    .GATE(net653),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit29.Q ));
 sg13g2_dlhq_1 _1122_ (.D(net793),
    .GATE(net653),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit28.Q ));
 sg13g2_dlhq_1 _1123_ (.D(net794),
    .GATE(net657),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit27.Q ));
 sg13g2_dlhq_1 _1124_ (.D(net795),
    .GATE(net657),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit26.Q ));
 sg13g2_dlhq_1 _1125_ (.D(net99),
    .GATE(net654),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit25.Q ));
 sg13g2_dlhq_1 _1126_ (.D(net797),
    .GATE(net654),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit24.Q ));
 sg13g2_dlhq_1 _1127_ (.D(net97),
    .GATE(net654),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit23.Q ));
 sg13g2_dlhq_1 _1128_ (.D(net96),
    .GATE(net655),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit22.Q ));
 sg13g2_dlhq_1 _1129_ (.D(net800),
    .GATE(net655),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit21.Q ));
 sg13g2_dlhq_1 _1130_ (.D(net801),
    .GATE(net655),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit20.Q ));
 sg13g2_dlhq_1 _1131_ (.D(net803),
    .GATE(net653),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit19.Q ));
 sg13g2_dlhq_1 _1132_ (.D(net91),
    .GATE(net653),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit18.Q ));
 sg13g2_dlhq_1 _1133_ (.D(net805),
    .GATE(net653),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit17.Q ));
 sg13g2_dlhq_1 _1134_ (.D(net806),
    .GATE(net657),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit16.Q ));
 sg13g2_dlhq_1 _1135_ (.D(net807),
    .GATE(net657),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit15.Q ));
 sg13g2_dlhq_1 _1136_ (.D(net808),
    .GATE(net657),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit14.Q ));
 sg13g2_dlhq_1 _1137_ (.D(net809),
    .GATE(net657),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit13.Q ));
 sg13g2_dlhq_1 _1138_ (.D(net810),
    .GATE(net657),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit12.Q ));
 sg13g2_dlhq_1 _1139_ (.D(net811),
    .GATE(net652),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit11.Q ));
 sg13g2_dlhq_1 _1140_ (.D(net812),
    .GATE(net652),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit10.Q ));
 sg13g2_dlhq_1 _1141_ (.D(net782),
    .GATE(net652),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit9.Q ));
 sg13g2_dlhq_1 _1142_ (.D(net783),
    .GATE(net652),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit8.Q ));
 sg13g2_dlhq_1 _1143_ (.D(net784),
    .GATE(net652),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit7.Q ));
 sg13g2_dlhq_1 _1144_ (.D(net785),
    .GATE(net652),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit6.Q ));
 sg13g2_dlhq_1 _1145_ (.D(net786),
    .GATE(net652),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit5.Q ));
 sg13g2_dlhq_1 _1146_ (.D(net787),
    .GATE(net652),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit4.Q ));
 sg13g2_dlhq_1 _1147_ (.D(net788),
    .GATE(net654),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit3.Q ));
 sg13g2_dlhq_1 _1148_ (.D(net791),
    .GATE(net654),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit2.Q ));
 sg13g2_dlhq_1 _1149_ (.D(net93),
    .GATE(net654),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit1.Q ));
 sg13g2_dlhq_1 _1150_ (.D(net82),
    .GATE(net654),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit0.Q ));
 sg13g2_dlhq_1 _1151_ (.D(net106),
    .GATE(net644),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame9_bit31.Q ));
 sg13g2_dlhq_1 _1152_ (.D(net105),
    .GATE(net644),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame9_bit30.Q ));
 sg13g2_dlhq_1 _1153_ (.D(net103),
    .GATE(net645),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame9_bit29.Q ));
 sg13g2_dlhq_1 _1154_ (.D(net102),
    .GATE(net644),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame9_bit28.Q ));
 sg13g2_dlhq_1 _1155_ (.D(net101),
    .GATE(net644),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame9_bit27.Q ));
 sg13g2_dlhq_1 _1156_ (.D(net795),
    .GATE(net644),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame9_bit26.Q ));
 sg13g2_dlhq_1 _1157_ (.D(net796),
    .GATE(net644),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame9_bit25.Q ));
 sg13g2_dlhq_1 _1158_ (.D(net98),
    .GATE(net644),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame9_bit24.Q ));
 sg13g2_dlhq_1 _1159_ (.D(net798),
    .GATE(net645),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame9_bit23.Q ));
 sg13g2_dlhq_1 _1160_ (.D(net799),
    .GATE(net645),
    .Q(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame9_bit22.Q ));
 sg13g2_dlhq_1 _1161_ (.D(net214),
    .GATE(net740),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame0_bit31.Q ));
 sg13g2_dlhq_1 _1162_ (.D(net213),
    .GATE(net740),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame0_bit30.Q ));
 sg13g2_dlhq_1 _1163_ (.D(net211),
    .GATE(net741),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame0_bit29.Q ));
 sg13g2_dlhq_1 _1164_ (.D(net210),
    .GATE(net741),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame0_bit28.Q ));
 sg13g2_dlhq_1 _1165_ (.D(net762),
    .GATE(net739),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame0_bit27.Q ));
 sg13g2_dlhq_1 _1166_ (.D(net763),
    .GATE(net739),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame0_bit26.Q ));
 sg13g2_dlhq_1 _1167_ (.D(net207),
    .GATE(net742),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame0_bit25.Q ));
 sg13g2_dlhq_1 _1168_ (.D(net206),
    .GATE(net742),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame0_bit24.Q ));
 sg13g2_dlhq_1 _1169_ (.D(net766),
    .GATE(net738),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame0_bit23.Q ));
 sg13g2_dlhq_1 _1170_ (.D(net767),
    .GATE(net738),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame0_bit22.Q ));
 sg13g2_dlhq_1 _1171_ (.D(net768),
    .GATE(net738),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame0_bit21.Q ));
 sg13g2_dlhq_1 _1172_ (.D(net769),
    .GATE(net738),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame0_bit20.Q ));
 sg13g2_dlhq_1 _1173_ (.D(net771),
    .GATE(net739),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame0_bit19.Q ));
 sg13g2_dlhq_1 _1174_ (.D(net772),
    .GATE(net739),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame0_bit18.Q ));
 sg13g2_dlhq_1 _1175_ (.D(net773),
    .GATE(net740),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame0_bit17.Q ));
 sg13g2_dlhq_1 _1176_ (.D(net774),
    .GATE(net740),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame0_bit16.Q ));
 sg13g2_dlhq_1 _1177_ (.D(net775),
    .GATE(net740),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame0_bit15.Q ));
 sg13g2_dlhq_1 _1178_ (.D(net776),
    .GATE(net741),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame0_bit14.Q ));
 sg13g2_dlhq_1 _1179_ (.D(net777),
    .GATE(net740),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame0_bit13.Q ));
 sg13g2_dlhq_1 _1180_ (.D(net778),
    .GATE(net740),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame0_bit12.Q ));
 sg13g2_dlhq_1 _1181_ (.D(net779),
    .GATE(net738),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame0_bit11.Q ));
 sg13g2_dlhq_1 _1182_ (.D(net780),
    .GATE(net738),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame0_bit10.Q ));
 sg13g2_dlhq_1 _1183_ (.D(net221),
    .GATE(net742),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame0_bit9.Q ));
 sg13g2_dlhq_1 _1184_ (.D(net220),
    .GATE(net742),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame0_bit8.Q ));
 sg13g2_dlhq_1 _1185_ (.D(net752),
    .GATE(net741),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame0_bit7.Q ));
 sg13g2_dlhq_1 _1186_ (.D(net753),
    .GATE(net740),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame0_bit6.Q ));
 sg13g2_dlhq_1 _1187_ (.D(net754),
    .GATE(net738),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame0_bit5.Q ));
 sg13g2_dlhq_1 _1188_ (.D(net755),
    .GATE(net738),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame0_bit4.Q ));
 sg13g2_dlhq_1 _1189_ (.D(net756),
    .GATE(net739),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame0_bit3.Q ));
 sg13g2_dlhq_1 _1190_ (.D(net759),
    .GATE(net739),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame0_bit2.Q ));
 sg13g2_dlhq_1 _1191_ (.D(net770),
    .GATE(net739),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame0_bit1.Q ));
 sg13g2_dlhq_1 _1192_ (.D(net781),
    .GATE(net739),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame0_bit0.Q ));
 sg13g2_dlhq_1 _1193_ (.D(net214),
    .GATE(net728),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit31.Q ));
 sg13g2_dlhq_1 _1194_ (.D(net213),
    .GATE(net728),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit30.Q ));
 sg13g2_dlhq_1 _1195_ (.D(net760),
    .GATE(net725),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit29.Q ));
 sg13g2_dlhq_1 _1196_ (.D(net761),
    .GATE(net725),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit28.Q ));
 sg13g2_dlhq_1 _1197_ (.D(net762),
    .GATE(net726),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit27.Q ));
 sg13g2_dlhq_1 _1198_ (.D(net763),
    .GATE(net725),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit26.Q ));
 sg13g2_dlhq_1 _1199_ (.D(net764),
    .GATE(net727),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit25.Q ));
 sg13g2_dlhq_1 _1200_ (.D(net765),
    .GATE(net727),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit24.Q ));
 sg13g2_dlhq_1 _1201_ (.D(net766),
    .GATE(net728),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit23.Q ));
 sg13g2_dlhq_1 _1202_ (.D(net767),
    .GATE(net728),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit22.Q ));
 sg13g2_dlhq_1 _1203_ (.D(net768),
    .GATE(net725),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit21.Q ));
 sg13g2_dlhq_1 _1204_ (.D(net769),
    .GATE(net725),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit20.Q ));
 sg13g2_dlhq_1 _1205_ (.D(net771),
    .GATE(net726),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit19.Q ));
 sg13g2_dlhq_1 _1206_ (.D(net772),
    .GATE(net725),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit18.Q ));
 sg13g2_dlhq_1 _1207_ (.D(net773),
    .GATE(net730),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit17.Q ));
 sg13g2_dlhq_1 _1208_ (.D(net774),
    .GATE(net730),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit16.Q ));
 sg13g2_dlhq_1 _1209_ (.D(net196),
    .GATE(net728),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit15.Q ));
 sg13g2_dlhq_1 _1210_ (.D(net195),
    .GATE(net728),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit14.Q ));
 sg13g2_dlhq_1 _1211_ (.D(net777),
    .GATE(net725),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit13.Q ));
 sg13g2_dlhq_1 _1212_ (.D(net778),
    .GATE(net725),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit12.Q ));
 sg13g2_dlhq_1 _1213_ (.D(net779),
    .GATE(net726),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit11.Q ));
 sg13g2_dlhq_1 _1214_ (.D(net780),
    .GATE(net726),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit10.Q ));
 sg13g2_dlhq_1 _1215_ (.D(net221),
    .GATE(net727),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit9.Q ));
 sg13g2_dlhq_1 _1216_ (.D(net220),
    .GATE(net730),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit8.Q ));
 sg13g2_dlhq_1 _1217_ (.D(net752),
    .GATE(net729),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit7.Q ));
 sg13g2_dlhq_1 _1218_ (.D(net753),
    .GATE(net728),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit6.Q ));
 sg13g2_dlhq_1 _1219_ (.D(net217),
    .GATE(net728),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit5.Q ));
 sg13g2_dlhq_1 _1220_ (.D(net216),
    .GATE(net729),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit4.Q ));
 sg13g2_dlhq_1 _1221_ (.D(net215),
    .GATE(net731),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit3.Q ));
 sg13g2_dlhq_1 _1222_ (.D(net212),
    .GATE(net729),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit2.Q ));
 sg13g2_dlhq_1 _1223_ (.D(net770),
    .GATE(net729),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit1.Q ));
 sg13g2_dlhq_1 _1224_ (.D(net781),
    .GATE(net729),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit0.Q ));
 sg13g2_dlhq_1 _1225_ (.D(net214),
    .GATE(net718),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit31.Q ));
 sg13g2_dlhq_1 _1226_ (.D(net213),
    .GATE(net718),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit30.Q ));
 sg13g2_dlhq_1 _1227_ (.D(net760),
    .GATE(net718),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit29.Q ));
 sg13g2_dlhq_1 _1228_ (.D(net761),
    .GATE(net718),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit28.Q ));
 sg13g2_dlhq_1 _1229_ (.D(net762),
    .GATE(net717),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit27.Q ));
 sg13g2_dlhq_1 _1230_ (.D(net763),
    .GATE(net717),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit26.Q ));
 sg13g2_dlhq_1 _1231_ (.D(net207),
    .GATE(net714),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit25.Q ));
 sg13g2_dlhq_1 _1232_ (.D(net206),
    .GATE(net714),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit24.Q ));
 sg13g2_dlhq_1 _1233_ (.D(net766),
    .GATE(net716),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit23.Q ));
 sg13g2_dlhq_1 _1234_ (.D(net767),
    .GATE(net716),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit22.Q ));
 sg13g2_dlhq_1 _1235_ (.D(net203),
    .GATE(net714),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit21.Q ));
 sg13g2_dlhq_1 _1236_ (.D(net202),
    .GATE(net715),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit20.Q ));
 sg13g2_dlhq_1 _1237_ (.D(net200),
    .GATE(net717),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit19.Q ));
 sg13g2_dlhq_1 _1238_ (.D(net199),
    .GATE(net717),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit18.Q ));
 sg13g2_dlhq_1 _1239_ (.D(net198),
    .GATE(net714),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit17.Q ));
 sg13g2_dlhq_1 _1240_ (.D(net197),
    .GATE(net714),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit16.Q ));
 sg13g2_dlhq_1 _1241_ (.D(net775),
    .GATE(net716),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit15.Q ));
 sg13g2_dlhq_1 _1242_ (.D(net776),
    .GATE(net716),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit14.Q ));
 sg13g2_dlhq_1 _1243_ (.D(net777),
    .GATE(net715),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit13.Q ));
 sg13g2_dlhq_1 _1244_ (.D(net778),
    .GATE(net715),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit12.Q ));
 sg13g2_dlhq_1 _1245_ (.D(net779),
    .GATE(net717),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit11.Q ));
 sg13g2_dlhq_1 _1246_ (.D(net780),
    .GATE(net717),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit10.Q ));
 sg13g2_dlhq_1 _1247_ (.D(net750),
    .GATE(net714),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit9.Q ));
 sg13g2_dlhq_1 _1248_ (.D(net751),
    .GATE(net715),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit8.Q ));
 sg13g2_dlhq_1 _1249_ (.D(net752),
    .GATE(net716),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit7.Q ));
 sg13g2_dlhq_1 _1250_ (.D(net753),
    .GATE(net716),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit6.Q ));
 sg13g2_dlhq_1 _1251_ (.D(net754),
    .GATE(net714),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit5.Q ));
 sg13g2_dlhq_1 _1252_ (.D(net216),
    .GATE(net715),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit4.Q ));
 sg13g2_dlhq_1 _1253_ (.D(net215),
    .GATE(net717),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit3.Q ));
 sg13g2_dlhq_1 _1254_ (.D(net212),
    .GATE(net717),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit2.Q ));
 sg13g2_dlhq_1 _1255_ (.D(net770),
    .GATE(net715),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit1.Q ));
 sg13g2_dlhq_1 _1256_ (.D(net190),
    .GATE(net714),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit0.Q ));
 sg13g2_dlhq_1 _1257_ (.D(net757),
    .GATE(net704),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame3_bit31.Q ));
 sg13g2_dlhq_1 _1258_ (.D(net758),
    .GATE(net704),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame3_bit30.Q ));
 sg13g2_dlhq_1 _1259_ (.D(net760),
    .GATE(net706),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame3_bit29.Q ));
 sg13g2_dlhq_1 _1260_ (.D(net761),
    .GATE(net706),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame3_bit28.Q ));
 sg13g2_dlhq_1 _1261_ (.D(net209),
    .GATE(net708),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame3_bit27.Q ));
 sg13g2_dlhq_1 _1262_ (.D(net208),
    .GATE(net708),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame3_bit26.Q ));
 sg13g2_dlhq_1 _1263_ (.D(net764),
    .GATE(net707),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame3_bit25.Q ));
 sg13g2_dlhq_1 _1264_ (.D(net765),
    .GATE(net707),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame3_bit24.Q ));
 sg13g2_dlhq_1 _1265_ (.D(net766),
    .GATE(net703),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame3_bit23.Q ));
 sg13g2_dlhq_1 _1266_ (.D(net767),
    .GATE(net703),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame3_bit22.Q ));
 sg13g2_dlhq_1 _1267_ (.D(net768),
    .GATE(net706),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame3_bit21.Q ));
 sg13g2_dlhq_1 _1268_ (.D(net769),
    .GATE(net706),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame3_bit20.Q ));
 sg13g2_dlhq_1 _1269_ (.D(net200),
    .GATE(net706),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame3_bit19.Q ));
 sg13g2_dlhq_1 _1270_ (.D(net199),
    .GATE(net706),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame3_bit18.Q ));
 sg13g2_dlhq_1 _1271_ (.D(net198),
    .GATE(net707),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame3_bit17.Q ));
 sg13g2_dlhq_1 _1272_ (.D(net197),
    .GATE(net707),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame3_bit16.Q ));
 sg13g2_dlhq_1 _1273_ (.D(net196),
    .GATE(net704),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame3_bit15.Q ));
 sg13g2_dlhq_1 _1274_ (.D(net195),
    .GATE(net704),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame3_bit14.Q ));
 sg13g2_dlhq_1 _1275_ (.D(net194),
    .GATE(net705),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame3_bit13.Q ));
 sg13g2_dlhq_1 _1276_ (.D(net778),
    .GATE(net705),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame3_bit12.Q ));
 sg13g2_dlhq_1 _1277_ (.D(net192),
    .GATE(net704),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame3_bit11.Q ));
 sg13g2_dlhq_1 _1278_ (.D(net191),
    .GATE(net705),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame3_bit10.Q ));
 sg13g2_dlhq_1 _1279_ (.D(net750),
    .GATE(net707),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame3_bit9.Q ));
 sg13g2_dlhq_1 _1280_ (.D(net751),
    .GATE(net707),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame3_bit8.Q ));
 sg13g2_dlhq_1 _1281_ (.D(net752),
    .GATE(net703),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame3_bit7.Q ));
 sg13g2_dlhq_1 _1282_ (.D(net753),
    .GATE(net703),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame3_bit6.Q ));
 sg13g2_dlhq_1 _1283_ (.D(net754),
    .GATE(net706),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame3_bit5.Q ));
 sg13g2_dlhq_1 _1284_ (.D(net755),
    .GATE(net706),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame3_bit4.Q ));
 sg13g2_dlhq_1 _1285_ (.D(net756),
    .GATE(net703),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame3_bit3.Q ));
 sg13g2_dlhq_1 _1286_ (.D(net759),
    .GATE(net703),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame3_bit2.Q ));
 sg13g2_dlhq_1 _1287_ (.D(net770),
    .GATE(net703),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame3_bit1.Q ));
 sg13g2_dlhq_1 _1288_ (.D(net781),
    .GATE(net703),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame3_bit0.Q ));
 sg13g2_dlhq_1 _1289_ (.D(net757),
    .GATE(net695),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame4_bit31.Q ));
 sg13g2_dlhq_1 _1290_ (.D(net758),
    .GATE(net694),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame4_bit30.Q ));
 sg13g2_dlhq_1 _1291_ (.D(net211),
    .GATE(net694),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame4_bit29.Q ));
 sg13g2_dlhq_1 _1292_ (.D(net210),
    .GATE(net694),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame4_bit28.Q ));
 sg13g2_dlhq_1 _1293_ (.D(net762),
    .GATE(net694),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame4_bit27.Q ));
 sg13g2_dlhq_1 _1294_ (.D(net763),
    .GATE(net694),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame4_bit26.Q ));
 sg13g2_dlhq_1 _1295_ (.D(net207),
    .GATE(net696),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame4_bit25.Q ));
 sg13g2_dlhq_1 _1296_ (.D(net206),
    .GATE(net696),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame4_bit24.Q ));
 sg13g2_dlhq_1 _1297_ (.D(net766),
    .GATE(net695),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame4_bit23.Q ));
 sg13g2_dlhq_1 _1298_ (.D(net767),
    .GATE(net694),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame4_bit22.Q ));
 sg13g2_dlhq_1 _1299_ (.D(net768),
    .GATE(net693),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame4_bit21.Q ));
 sg13g2_dlhq_1 _1300_ (.D(net769),
    .GATE(net693),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame4_bit20.Q ));
 sg13g2_dlhq_1 _1301_ (.D(net771),
    .GATE(net693),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame4_bit19.Q ));
 sg13g2_dlhq_1 _1302_ (.D(net772),
    .GATE(net692),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame4_bit18.Q ));
 sg13g2_dlhq_1 _1303_ (.D(net773),
    .GATE(net694),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame4_bit17.Q ));
 sg13g2_dlhq_1 _1304_ (.D(net774),
    .GATE(net694),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame4_bit16.Q ));
 sg13g2_dlhq_1 _1305_ (.D(net775),
    .GATE(net693),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame4_bit15.Q ));
 sg13g2_dlhq_1 _1306_ (.D(net776),
    .GATE(net695),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame4_bit14.Q ));
 sg13g2_dlhq_1 _1307_ (.D(net777),
    .GATE(net693),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame4_bit13.Q ));
 sg13g2_dlhq_1 _1308_ (.D(net778),
    .GATE(net695),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame4_bit12.Q ));
 sg13g2_dlhq_1 _1309_ (.D(net779),
    .GATE(net692),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame4_bit11.Q ));
 sg13g2_dlhq_1 _1310_ (.D(net780),
    .GATE(net692),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame4_bit10.Q ));
 sg13g2_dlhq_1 _1311_ (.D(net750),
    .GATE(net693),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame4_bit9.Q ));
 sg13g2_dlhq_1 _1312_ (.D(net751),
    .GATE(net692),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame4_bit8.Q ));
 sg13g2_dlhq_1 _1313_ (.D(net752),
    .GATE(net695),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame4_bit7.Q ));
 sg13g2_dlhq_1 _1314_ (.D(net753),
    .GATE(net693),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame4_bit6.Q ));
 sg13g2_dlhq_1 _1315_ (.D(net754),
    .GATE(net692),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame4_bit5.Q ));
 sg13g2_dlhq_1 _1316_ (.D(net755),
    .GATE(net692),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame4_bit4.Q ));
 sg13g2_dlhq_1 _1317_ (.D(net756),
    .GATE(net692),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame4_bit3.Q ));
 sg13g2_dlhq_1 _1318_ (.D(net759),
    .GATE(net692),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame4_bit2.Q ));
 sg13g2_dlhq_1 _1319_ (.D(net201),
    .GATE(net696),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame4_bit1.Q ));
 sg13g2_dlhq_1 _1320_ (.D(net190),
    .GATE(net696),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame4_bit0.Q ));
 sg13g2_dlhq_1 _1321_ (.D(net757),
    .GATE(net682),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame5_bit31.Q ));
 sg13g2_dlhq_1 _1322_ (.D(net758),
    .GATE(net682),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame5_bit30.Q ));
 sg13g2_dlhq_1 _1323_ (.D(net760),
    .GATE(net682),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame5_bit29.Q ));
 sg13g2_dlhq_1 _1324_ (.D(net761),
    .GATE(net683),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame5_bit28.Q ));
 sg13g2_dlhq_1 _1325_ (.D(net762),
    .GATE(net683),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame5_bit27.Q ));
 sg13g2_dlhq_1 _1326_ (.D(net763),
    .GATE(net681),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame5_bit26.Q ));
 sg13g2_dlhq_1 _1327_ (.D(net764),
    .GATE(net681),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame5_bit25.Q ));
 sg13g2_dlhq_1 _1328_ (.D(net765),
    .GATE(net681),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame5_bit24.Q ));
 sg13g2_dlhq_1 _1329_ (.D(net766),
    .GATE(net683),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame5_bit23.Q ));
 sg13g2_dlhq_1 _1330_ (.D(net767),
    .GATE(net683),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame5_bit22.Q ));
 sg13g2_dlhq_1 _1331_ (.D(net768),
    .GATE(net681),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame5_bit21.Q ));
 sg13g2_dlhq_1 _1332_ (.D(net769),
    .GATE(net681),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame5_bit20.Q ));
 sg13g2_dlhq_1 _1333_ (.D(net771),
    .GATE(net684),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame5_bit19.Q ));
 sg13g2_dlhq_1 _1334_ (.D(net772),
    .GATE(net684),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame5_bit18.Q ));
 sg13g2_dlhq_1 _1335_ (.D(net773),
    .GATE(net681),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame5_bit17.Q ));
 sg13g2_dlhq_1 _1336_ (.D(net774),
    .GATE(net681),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame5_bit16.Q ));
 sg13g2_dlhq_1 _1337_ (.D(net775),
    .GATE(net682),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame5_bit15.Q ));
 sg13g2_dlhq_1 _1338_ (.D(net776),
    .GATE(net682),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame5_bit14.Q ));
 sg13g2_dlhq_1 _1339_ (.D(net777),
    .GATE(net682),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame5_bit13.Q ));
 sg13g2_dlhq_1 _1340_ (.D(net778),
    .GATE(net680),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame5_bit12.Q ));
 sg13g2_dlhq_1 _1341_ (.D(net779),
    .GATE(net680),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame5_bit11.Q ));
 sg13g2_dlhq_1 _1342_ (.D(net780),
    .GATE(net680),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame5_bit10.Q ));
 sg13g2_dlhq_1 _1343_ (.D(net750),
    .GATE(net684),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame5_bit9.Q ));
 sg13g2_dlhq_1 _1344_ (.D(net751),
    .GATE(net680),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame5_bit8.Q ));
 sg13g2_dlhq_1 _1345_ (.D(net752),
    .GATE(net682),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame5_bit7.Q ));
 sg13g2_dlhq_1 _1346_ (.D(net753),
    .GATE(net682),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame5_bit6.Q ));
 sg13g2_dlhq_1 _1347_ (.D(net754),
    .GATE(net680),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame5_bit5.Q ));
 sg13g2_dlhq_1 _1348_ (.D(net755),
    .GATE(net680),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame5_bit4.Q ));
 sg13g2_dlhq_1 _1349_ (.D(net756),
    .GATE(net680),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame5_bit3.Q ));
 sg13g2_dlhq_1 _1350_ (.D(net759),
    .GATE(net680),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame5_bit2.Q ));
 sg13g2_dlhq_1 _1351_ (.D(net770),
    .GATE(net691),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame5_bit1.Q ));
 sg13g2_dlhq_1 _1352_ (.D(net781),
    .GATE(net691),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame5_bit0.Q ));
 sg13g2_dlhq_1 _1353_ (.D(net757),
    .GATE(net672),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame6_bit31.Q ));
 sg13g2_dlhq_1 _1354_ (.D(net758),
    .GATE(net671),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame6_bit30.Q ));
 sg13g2_dlhq_1 _1355_ (.D(net760),
    .GATE(net671),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame6_bit29.Q ));
 sg13g2_dlhq_1 _1356_ (.D(net761),
    .GATE(net671),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame6_bit28.Q ));
 sg13g2_dlhq_1 _1357_ (.D(net762),
    .GATE(net669),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame6_bit27.Q ));
 sg13g2_dlhq_1 _1358_ (.D(net763),
    .GATE(net670),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame6_bit26.Q ));
 sg13g2_dlhq_1 _1359_ (.D(net764),
    .GATE(net673),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame6_bit25.Q ));
 sg13g2_dlhq_1 _1360_ (.D(net765),
    .GATE(net673),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame6_bit24.Q ));
 sg13g2_dlhq_1 _1361_ (.D(net766),
    .GATE(net671),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame6_bit23.Q ));
 sg13g2_dlhq_1 _1362_ (.D(net767),
    .GATE(net671),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame6_bit22.Q ));
 sg13g2_dlhq_1 _1363_ (.D(net768),
    .GATE(net669),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame6_bit21.Q ));
 sg13g2_dlhq_1 _1364_ (.D(net769),
    .GATE(net669),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame6_bit20.Q ));
 sg13g2_dlhq_1 _1365_ (.D(net771),
    .GATE(net673),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame6_bit19.Q ));
 sg13g2_dlhq_1 _1366_ (.D(net772),
    .GATE(net673),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame6_bit18.Q ));
 sg13g2_dlhq_1 _1367_ (.D(net773),
    .GATE(net674),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame6_bit17.Q ));
 sg13g2_dlhq_1 _1368_ (.D(net774),
    .GATE(net674),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame6_bit16.Q ));
 sg13g2_dlhq_1 _1369_ (.D(net775),
    .GATE(net672),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame6_bit15.Q ));
 sg13g2_dlhq_1 _1370_ (.D(net776),
    .GATE(net670),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame6_bit14.Q ));
 sg13g2_dlhq_1 _1371_ (.D(net777),
    .GATE(net671),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame6_bit13.Q ));
 sg13g2_dlhq_1 _1372_ (.D(net778),
    .GATE(net669),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame6_bit12.Q ));
 sg13g2_dlhq_1 _1373_ (.D(net779),
    .GATE(net669),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame6_bit11.Q ));
 sg13g2_dlhq_1 _1374_ (.D(net780),
    .GATE(net669),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame6_bit10.Q ));
 sg13g2_dlhq_1 _1375_ (.D(net750),
    .GATE(net670),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame6_bit9.Q ));
 sg13g2_dlhq_1 _1376_ (.D(net751),
    .GATE(net670),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame6_bit8.Q ));
 sg13g2_dlhq_1 _1377_ (.D(net752),
    .GATE(net671),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame6_bit7.Q ));
 sg13g2_dlhq_1 _1378_ (.D(net753),
    .GATE(net671),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame6_bit6.Q ));
 sg13g2_dlhq_1 _1379_ (.D(net754),
    .GATE(net669),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame6_bit5.Q ));
 sg13g2_dlhq_1 _1380_ (.D(net755),
    .GATE(net669),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame6_bit4.Q ));
 sg13g2_dlhq_1 _1381_ (.D(net756),
    .GATE(net670),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame6_bit3.Q ));
 sg13g2_dlhq_1 _1382_ (.D(net759),
    .GATE(net670),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame6_bit2.Q ));
 sg13g2_dlhq_1 _1383_ (.D(net770),
    .GATE(net674),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame6_bit1.Q ));
 sg13g2_dlhq_1 _1384_ (.D(net781),
    .GATE(net674),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame6_bit0.Q ));
 sg13g2_dlhq_1 _1385_ (.D(net757),
    .GATE(net658),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit31.Q ));
 sg13g2_dlhq_1 _1386_ (.D(net758),
    .GATE(net658),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit30.Q ));
 sg13g2_dlhq_1 _1387_ (.D(net760),
    .GATE(net661),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit29.Q ));
 sg13g2_dlhq_1 _1388_ (.D(net761),
    .GATE(net658),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit28.Q ));
 sg13g2_dlhq_1 _1389_ (.D(net762),
    .GATE(net658),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit27.Q ));
 sg13g2_dlhq_1 _1390_ (.D(net763),
    .GATE(net658),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit26.Q ));
 sg13g2_dlhq_1 _1391_ (.D(net764),
    .GATE(net659),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit25.Q ));
 sg13g2_dlhq_1 _1392_ (.D(net765),
    .GATE(net659),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit24.Q ));
 sg13g2_dlhq_1 _1393_ (.D(net766),
    .GATE(net661),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit23.Q ));
 sg13g2_dlhq_1 _1394_ (.D(net767),
    .GATE(net658),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit22.Q ));
 sg13g2_dlhq_1 _1395_ (.D(net768),
    .GATE(net658),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit21.Q ));
 sg13g2_dlhq_1 _1396_ (.D(net769),
    .GATE(net658),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit20.Q ));
 sg13g2_dlhq_1 _1397_ (.D(net771),
    .GATE(net659),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit19.Q ));
 sg13g2_dlhq_1 _1398_ (.D(net772),
    .GATE(net659),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit18.Q ));
 sg13g2_dlhq_1 _1399_ (.D(net773),
    .GATE(net662),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit17.Q ));
 sg13g2_dlhq_1 _1400_ (.D(net774),
    .GATE(net662),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit16.Q ));
 sg13g2_dlhq_1 _1401_ (.D(net196),
    .GATE(net662),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit15.Q ));
 sg13g2_dlhq_1 _1402_ (.D(net195),
    .GATE(net662),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit14.Q ));
 sg13g2_dlhq_1 _1403_ (.D(net194),
    .GATE(net668),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit13.Q ));
 sg13g2_dlhq_1 _1404_ (.D(net193),
    .GATE(net662),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit12.Q ));
 sg13g2_dlhq_1 _1405_ (.D(net779),
    .GATE(net660),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit11.Q ));
 sg13g2_dlhq_1 _1406_ (.D(net780),
    .GATE(net660),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit10.Q ));
 sg13g2_dlhq_1 _1407_ (.D(net750),
    .GATE(net660),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit9.Q ));
 sg13g2_dlhq_1 _1408_ (.D(net751),
    .GATE(net662),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit8.Q ));
 sg13g2_dlhq_1 _1409_ (.D(net219),
    .GATE(net662),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit7.Q ));
 sg13g2_dlhq_1 _1410_ (.D(net218),
    .GATE(net662),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit6.Q ));
 sg13g2_dlhq_1 _1411_ (.D(net754),
    .GATE(net659),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit5.Q ));
 sg13g2_dlhq_1 _1412_ (.D(net755),
    .GATE(net659),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit4.Q ));
 sg13g2_dlhq_1 _1413_ (.D(net756),
    .GATE(net660),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit3.Q ));
 sg13g2_dlhq_1 _1414_ (.D(net759),
    .GATE(net659),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit2.Q ));
 sg13g2_dlhq_1 _1415_ (.D(net770),
    .GATE(net660),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit1.Q ));
 sg13g2_dlhq_1 _1416_ (.D(net781),
    .GATE(net659),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit0.Q ));
 sg13g2_dlhq_1 _1417_ (.D(net757),
    .GATE(net647),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit31.Q ));
 sg13g2_dlhq_1 _1418_ (.D(net758),
    .GATE(net647),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit30.Q ));
 sg13g2_dlhq_1 _1419_ (.D(net211),
    .GATE(net649),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit29.Q ));
 sg13g2_dlhq_1 _1420_ (.D(net210),
    .GATE(net649),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit28.Q ));
 sg13g2_dlhq_1 _1421_ (.D(net209),
    .GATE(net649),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit27.Q ));
 sg13g2_dlhq_1 _1422_ (.D(net208),
    .GATE(net649),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit26.Q ));
 sg13g2_dlhq_1 _1423_ (.D(net764),
    .GATE(net647),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit25.Q ));
 sg13g2_dlhq_1 _1424_ (.D(net765),
    .GATE(net647),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit24.Q ));
 sg13g2_dlhq_1 _1425_ (.D(net205),
    .GATE(net647),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit23.Q ));
 sg13g2_dlhq_1 _1426_ (.D(net204),
    .GATE(net647),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit22.Q ));
 sg13g2_dlhq_1 _1427_ (.D(net768),
    .GATE(net651),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit21.Q ));
 sg13g2_dlhq_1 _1428_ (.D(net769),
    .GATE(net651),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit20.Q ));
 sg13g2_dlhq_1 _1429_ (.D(net200),
    .GATE(net650),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit19.Q ));
 sg13g2_dlhq_1 _1430_ (.D(net199),
    .GATE(net650),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit18.Q ));
 sg13g2_dlhq_1 _1431_ (.D(net773),
    .GATE(net648),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit17.Q ));
 sg13g2_dlhq_1 _1432_ (.D(net774),
    .GATE(net648),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit16.Q ));
 sg13g2_dlhq_1 _1433_ (.D(net775),
    .GATE(net649),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit15.Q ));
 sg13g2_dlhq_1 _1434_ (.D(net776),
    .GATE(net649),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit14.Q ));
 sg13g2_dlhq_1 _1435_ (.D(net777),
    .GATE(net651),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit13.Q ));
 sg13g2_dlhq_1 _1436_ (.D(net193),
    .GATE(net651),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit12.Q ));
 sg13g2_dlhq_1 _1437_ (.D(net192),
    .GATE(net651),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit11.Q ));
 sg13g2_dlhq_1 _1438_ (.D(net191),
    .GATE(net222),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit10.Q ));
 sg13g2_dlhq_1 _1439_ (.D(net750),
    .GATE(net650),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit9.Q ));
 sg13g2_dlhq_1 _1440_ (.D(net751),
    .GATE(net650),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit8.Q ));
 sg13g2_dlhq_1 _1441_ (.D(net752),
    .GATE(net648),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit7.Q ));
 sg13g2_dlhq_1 _1442_ (.D(net753),
    .GATE(net648),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit6.Q ));
 sg13g2_dlhq_1 _1443_ (.D(net754),
    .GATE(net648),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit5.Q ));
 sg13g2_dlhq_1 _1444_ (.D(net755),
    .GATE(net649),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit4.Q ));
 sg13g2_dlhq_1 _1445_ (.D(net756),
    .GATE(net649),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit3.Q ));
 sg13g2_dlhq_1 _1446_ (.D(net759),
    .GATE(net650),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit2.Q ));
 sg13g2_dlhq_1 _1447_ (.D(net770),
    .GATE(net647),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit1.Q ));
 sg13g2_dlhq_1 _1448_ (.D(net781),
    .GATE(net647),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit0.Q ));
 sg13g2_dlhq_1 _1449_ (.D(net757),
    .GATE(net641),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame9_bit31.Q ));
 sg13g2_dlhq_1 _1450_ (.D(net758),
    .GATE(net641),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame9_bit30.Q ));
 sg13g2_dlhq_1 _1451_ (.D(net760),
    .GATE(net641),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame9_bit29.Q ));
 sg13g2_dlhq_1 _1452_ (.D(net761),
    .GATE(net641),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame9_bit28.Q ));
 sg13g2_dlhq_1 _1453_ (.D(net762),
    .GATE(net642),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame9_bit27.Q ));
 sg13g2_dlhq_1 _1454_ (.D(net763),
    .GATE(net642),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame9_bit26.Q ));
 sg13g2_dlhq_1 _1455_ (.D(net764),
    .GATE(net642),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame9_bit25.Q ));
 sg13g2_dlhq_1 _1456_ (.D(net765),
    .GATE(net642),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame9_bit24.Q ));
 sg13g2_dlhq_1 _1457_ (.D(net205),
    .GATE(net642),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame9_bit23.Q ));
 sg13g2_dlhq_1 _1458_ (.D(net204),
    .GATE(net642),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame9_bit22.Q ));
 sg13g2_dlhq_1 _1459_ (.D(net203),
    .GATE(net641),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame9_bit21.Q ));
 sg13g2_dlhq_1 _1460_ (.D(net202),
    .GATE(net641),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame9_bit20.Q ));
 sg13g2_dlhq_1 _1461_ (.D(net771),
    .GATE(net641),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame9_bit19.Q ));
 sg13g2_dlhq_1 _1462_ (.D(net772),
    .GATE(net641),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame9_bit18.Q ));
 sg13g2_dlhq_1 _1463_ (.D(net773),
    .GATE(net646),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame9_bit17.Q ));
 sg13g2_dlhq_1 _1464_ (.D(net774),
    .GATE(net646),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame9_bit16.Q ));
 sg13g2_dlhq_1 _1465_ (.D(net775),
    .GATE(net643),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame9_bit15.Q ));
 sg13g2_dlhq_1 _1466_ (.D(net776),
    .GATE(net642),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame9_bit14.Q ));
 sg13g2_dlhq_1 _1467_ (.D(net777),
    .GATE(net643),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame9_bit13.Q ));
 sg13g2_dlhq_1 _1468_ (.D(net778),
    .GATE(net643),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame9_bit12.Q ));
 sg13g2_dlhq_1 _1469_ (.D(net192),
    .GATE(net642),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame9_bit11.Q ));
 sg13g2_dlhq_1 _1470_ (.D(net191),
    .GATE(net643),
    .Q(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame9_bit10.Q ));
 sg13g2_fill_1 FILLER_0_0 ();
 sg13g2_tiehi IHP_SRAM_583 (.L_HI(net583));
 sg13g2_buf_1 _1473_ (.A(Tile_X0Y1_UserCLK),
    .X(net293));
 sg13g2_buf_1 _1474_ (.A(net813),
    .X(net328));
 sg13g2_buf_1 _1475_ (.A(net802),
    .X(net339));
 sg13g2_buf_1 _1476_ (.A(net791),
    .X(net350));
 sg13g2_buf_1 _1477_ (.A(net788),
    .X(net353));
 sg13g2_buf_1 _1478_ (.A(net787),
    .X(net354));
 sg13g2_buf_1 _1479_ (.A(net786),
    .X(net355));
 sg13g2_buf_1 _1480_ (.A(net785),
    .X(net356));
 sg13g2_buf_1 _1481_ (.A(net784),
    .X(net357));
 sg13g2_buf_1 _1482_ (.A(net783),
    .X(net358));
 sg13g2_buf_1 _1483_ (.A(net113),
    .X(net359));
 sg13g2_buf_1 _1484_ (.A(net812),
    .X(net329));
 sg13g2_buf_1 _1485_ (.A(net811),
    .X(net330));
 sg13g2_buf_1 _1486_ (.A(net810),
    .X(net331));
 sg13g2_buf_1 _1487_ (.A(net809),
    .X(net332));
 sg13g2_buf_1 _1488_ (.A(net808),
    .X(net333));
 sg13g2_buf_1 _1489_ (.A(net807),
    .X(net334));
 sg13g2_buf_1 _1490_ (.A(net806),
    .X(net335));
 sg13g2_buf_1 _1491_ (.A(net805),
    .X(net336));
 sg13g2_buf_1 _1492_ (.A(net804),
    .X(net337));
 sg13g2_buf_1 _1493_ (.A(net92),
    .X(net338));
 sg13g2_buf_1 _1494_ (.A(net801),
    .X(net340));
 sg13g2_buf_1 _1495_ (.A(net800),
    .X(net341));
 sg13g2_buf_1 _1496_ (.A(net96),
    .X(net342));
 sg13g2_buf_1 _1497_ (.A(net97),
    .X(net343));
 sg13g2_buf_1 _1498_ (.A(net98),
    .X(net344));
 sg13g2_buf_1 _1499_ (.A(net99),
    .X(net345));
 sg13g2_buf_1 _1500_ (.A(net795),
    .X(net346));
 sg13g2_buf_1 _1501_ (.A(net794),
    .X(net347));
 sg13g2_buf_1 _1502_ (.A(net793),
    .X(net348));
 sg13g2_buf_1 _1503_ (.A(net792),
    .X(net349));
 sg13g2_buf_1 _1504_ (.A(net790),
    .X(net351));
 sg13g2_buf_1 _1505_ (.A(net789),
    .X(net352));
 sg13g2_buf_1 _1506_ (.A(net746),
    .X(net360));
 sg13g2_buf_1 _1507_ (.A(net734),
    .X(net371));
 sg13g2_buf_1 _1508_ (.A(net721),
    .X(net372));
 sg13g2_buf_1 _1509_ (.A(net710),
    .X(net373));
 sg13g2_buf_1 _1510_ (.A(net701),
    .X(net374));
 sg13g2_buf_1 _1511_ (.A(net687),
    .X(net375));
 sg13g2_buf_1 _1512_ (.A(net678),
    .X(net376));
 sg13g2_buf_1 _1513_ (.A(net667),
    .X(net377));
 sg13g2_buf_1 _1514_ (.A(net654),
    .X(net378));
 sg13g2_buf_1 _1515_ (.A(net644),
    .X(net379));
 sg13g2_buf_1 _1516_ (.A(Tile_X0Y1_FrameStrobe[10]),
    .X(net361));
 sg13g2_buf_1 _1517_ (.A(Tile_X0Y1_FrameStrobe[11]),
    .X(net362));
 sg13g2_buf_1 _1518_ (.A(Tile_X0Y1_FrameStrobe[12]),
    .X(net363));
 sg13g2_buf_1 _1519_ (.A(Tile_X0Y1_FrameStrobe[13]),
    .X(net364));
 sg13g2_buf_1 _1520_ (.A(Tile_X0Y1_FrameStrobe[14]),
    .X(net365));
 sg13g2_buf_1 _1521_ (.A(Tile_X0Y1_FrameStrobe[15]),
    .X(net366));
 sg13g2_buf_1 _1522_ (.A(Tile_X0Y1_FrameStrobe[16]),
    .X(net367));
 sg13g2_buf_1 _1523_ (.A(Tile_X0Y1_FrameStrobe[17]),
    .X(net368));
 sg13g2_buf_1 _1524_ (.A(Tile_X0Y1_FrameStrobe[18]),
    .X(net369));
 sg13g2_buf_1 _1525_ (.A(Tile_X0Y1_FrameStrobe[19]),
    .X(net370));
 sg13g2_buf_1 _1526_ (.A(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.N1BEG0 ),
    .X(net380));
 sg13g2_buf_1 _1527_ (.A(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.N1BEG1 ),
    .X(net381));
 sg13g2_buf_1 _1528_ (.A(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.N1BEG2 ),
    .X(net382));
 sg13g2_buf_1 _1529_ (.A(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.N1BEG3 ),
    .X(net383));
 sg13g2_buf_1 _1530_ (.A(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.N2BEG0 ),
    .X(net384));
 sg13g2_buf_1 _1531_ (.A(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.N2BEG1 ),
    .X(net385));
 sg13g2_buf_1 _1532_ (.A(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.N2BEG2 ),
    .X(net386));
 sg13g2_buf_1 _1533_ (.A(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.N2BEG3 ),
    .X(net387));
 sg13g2_buf_1 _1534_ (.A(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.N2BEG4 ),
    .X(net388));
 sg13g2_buf_1 _1535_ (.A(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.N2BEG5 ),
    .X(net389));
 sg13g2_buf_1 _1536_ (.A(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.N2BEG6 ),
    .X(net390));
 sg13g2_buf_1 _1537_ (.A(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.N2BEG7 ),
    .X(net391));
 sg13g2_buf_1 _1538_ (.A(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.N2BEGb0 ),
    .X(net392));
 sg13g2_buf_1 _1539_ (.A(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.N2BEGb1 ),
    .X(net393));
 sg13g2_buf_1 _1540_ (.A(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.N2BEGb2 ),
    .X(net394));
 sg13g2_buf_1 _1541_ (.A(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.N2BEGb3 ),
    .X(net395));
 sg13g2_buf_1 _1542_ (.A(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.N2BEGb4 ),
    .X(net396));
 sg13g2_buf_1 _1543_ (.A(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.N2BEGb5 ),
    .X(net397));
 sg13g2_buf_1 _1544_ (.A(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.N2BEGb6 ),
    .X(net398));
 sg13g2_buf_1 _1545_ (.A(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.N2BEGb7 ),
    .X(net399));
 sg13g2_buf_1 _1546_ (.A(Tile_X0Y1_N4END[8]),
    .X(net400));
 sg13g2_buf_1 _1547_ (.A(Tile_X0Y1_N4END[9]),
    .X(net407));
 sg13g2_buf_1 _1548_ (.A(Tile_X0Y1_N4END[10]),
    .X(net408));
 sg13g2_buf_1 _1549_ (.A(Tile_X0Y1_N4END[11]),
    .X(net409));
 sg13g2_buf_1 _1550_ (.A(Tile_X0Y1_N4END[12]),
    .X(net410));
 sg13g2_buf_1 _1551_ (.A(Tile_X0Y1_N4END[13]),
    .X(net411));
 sg13g2_buf_1 _1552_ (.A(Tile_X0Y1_N4END[14]),
    .X(net412));
 sg13g2_buf_1 _1553_ (.A(Tile_X0Y1_N4END[15]),
    .X(net413));
 sg13g2_buf_1 _1554_ (.A(\Tile_X0Y0_IHP_SRAM_top.N4BEG_outbuf_8.A ),
    .X(net414));
 sg13g2_buf_1 _1555_ (.A(\Tile_X0Y0_IHP_SRAM_top.N4BEG_outbuf_9.A ),
    .X(net415));
 sg13g2_buf_1 _1556_ (.A(\Tile_X0Y0_IHP_SRAM_top.N4BEG_outbuf_10.A ),
    .X(net401));
 sg13g2_buf_1 _1557_ (.A(\Tile_X0Y0_IHP_SRAM_top.N4BEG_outbuf_11.A ),
    .X(net402));
 sg13g2_buf_1 _1558_ (.A(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.N4BEG0 ),
    .X(net403));
 sg13g2_buf_1 _1559_ (.A(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.N4BEG1 ),
    .X(net404));
 sg13g2_buf_1 _1560_ (.A(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.N4BEG2 ),
    .X(net405));
 sg13g2_buf_1 _1561_ (.A(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.N4BEG3 ),
    .X(net406));
 sg13g2_buf_1 _1562_ (.A(Tile_X0Y1_UserCLK),
    .X(net416));
 sg13g2_buf_1 _1563_ (.A(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.W1BEG0 ),
    .X(net417));
 sg13g2_buf_1 _1564_ (.A(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.W1BEG1 ),
    .X(net418));
 sg13g2_buf_1 _1565_ (.A(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.W1BEG2 ),
    .X(net419));
 sg13g2_buf_1 _1566_ (.A(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.W1BEG3 ),
    .X(net420));
 sg13g2_buf_1 _1567_ (.A(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.W2BEG0 ),
    .X(net421));
 sg13g2_buf_1 _1568_ (.A(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.W2BEG1 ),
    .X(net422));
 sg13g2_buf_1 _1569_ (.A(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.W2BEG2 ),
    .X(net423));
 sg13g2_buf_1 _1570_ (.A(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.W2BEG3 ),
    .X(net424));
 sg13g2_buf_1 _1571_ (.A(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.W2BEG4 ),
    .X(net425));
 sg13g2_buf_1 _1572_ (.A(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.W2BEG5 ),
    .X(net426));
 sg13g2_buf_1 _1573_ (.A(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.W2BEG6 ),
    .X(net427));
 sg13g2_buf_1 _1574_ (.A(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.W2BEG7 ),
    .X(net428));
 sg13g2_buf_1 _1575_ (.A(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.W2BEGb0 ),
    .X(net429));
 sg13g2_buf_1 _1576_ (.A(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.W2BEGb1 ),
    .X(net430));
 sg13g2_buf_1 _1577_ (.A(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.W2BEGb2 ),
    .X(net431));
 sg13g2_buf_1 _1578_ (.A(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.W2BEGb3 ),
    .X(net432));
 sg13g2_buf_1 _1579_ (.A(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.W2BEGb4 ),
    .X(net433));
 sg13g2_buf_1 _1580_ (.A(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.W2BEGb5 ),
    .X(net434));
 sg13g2_buf_1 _1581_ (.A(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.W2BEGb6 ),
    .X(net435));
 sg13g2_buf_1 _1582_ (.A(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.W2BEGb7 ),
    .X(net436));
 sg13g2_buf_1 _1583_ (.A(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.W6BEG0 ),
    .X(net437));
 sg13g2_buf_1 _1584_ (.A(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.W6BEG1 ),
    .X(net440));
 sg13g2_buf_1 _1585_ (.A(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.W6BEG2 ),
    .X(net441));
 sg13g2_buf_1 _1586_ (.A(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.W6BEG3 ),
    .X(net442));
 sg13g2_buf_1 _1587_ (.A(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.W6BEG4 ),
    .X(net443));
 sg13g2_buf_1 _1588_ (.A(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.W6BEG5 ),
    .X(net444));
 sg13g2_buf_1 _1589_ (.A(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.W6BEG6 ),
    .X(net445));
 sg13g2_buf_1 _1590_ (.A(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.W6BEG7 ),
    .X(net446));
 sg13g2_buf_1 _1591_ (.A(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.W6BEG8 ),
    .X(net447));
 sg13g2_buf_1 _1592_ (.A(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.W6BEG9 ),
    .X(net448));
 sg13g2_buf_1 _1593_ (.A(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.W6BEG10 ),
    .X(net438));
 sg13g2_buf_1 _1594_ (.A(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.W6BEG11 ),
    .X(net439));
 sg13g2_buf_1 _1595_ (.A(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.WW4BEG0 ),
    .X(net449));
 sg13g2_buf_1 _1596_ (.A(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.WW4BEG1 ),
    .X(net456));
 sg13g2_buf_1 _1597_ (.A(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.WW4BEG2 ),
    .X(net457));
 sg13g2_buf_1 _1598_ (.A(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.WW4BEG3 ),
    .X(net458));
 sg13g2_buf_1 _1599_ (.A(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.WW4BEG4 ),
    .X(net459));
 sg13g2_buf_1 _1600_ (.A(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.WW4BEG5 ),
    .X(net460));
 sg13g2_buf_1 _1601_ (.A(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.WW4BEG6 ),
    .X(net461));
 sg13g2_buf_1 _1602_ (.A(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.WW4BEG7 ),
    .X(net462));
 sg13g2_buf_1 _1603_ (.A(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.WW4BEG8 ),
    .X(net463));
 sg13g2_buf_1 _1604_ (.A(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.WW4BEG9 ),
    .X(net464));
 sg13g2_buf_1 _1605_ (.A(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.WW4BEG10 ),
    .X(net450));
 sg13g2_buf_1 _1606_ (.A(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.WW4BEG11 ),
    .X(net451));
 sg13g2_buf_1 _1607_ (.A(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.WW4BEG12 ),
    .X(net452));
 sg13g2_buf_1 _1608_ (.A(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.WW4BEG13 ),
    .X(net453));
 sg13g2_buf_1 _1609_ (.A(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.WW4BEG14 ),
    .X(net454));
 sg13g2_buf_1 _1610_ (.A(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.WW4BEG15 ),
    .X(net455));
 sg13g2_buf_1 _1611_ (.A(net781),
    .X(net465));
 sg13g2_buf_1 _1612_ (.A(net201),
    .X(net476));
 sg13g2_buf_1 _1613_ (.A(net759),
    .X(net487));
 sg13g2_buf_1 _1614_ (.A(net756),
    .X(net490));
 sg13g2_buf_1 _1615_ (.A(net755),
    .X(net491));
 sg13g2_buf_1 _1616_ (.A(net217),
    .X(net492));
 sg13g2_buf_1 _1617_ (.A(net218),
    .X(net493));
 sg13g2_buf_1 _1618_ (.A(net219),
    .X(net494));
 sg13g2_buf_1 _1619_ (.A(net751),
    .X(net495));
 sg13g2_buf_1 _1620_ (.A(net750),
    .X(net496));
 sg13g2_buf_1 _1621_ (.A(net780),
    .X(net466));
 sg13g2_buf_1 _1622_ (.A(net779),
    .X(net467));
 sg13g2_buf_1 _1623_ (.A(net193),
    .X(net468));
 sg13g2_buf_1 _1624_ (.A(net194),
    .X(net469));
 sg13g2_buf_1 _1625_ (.A(net776),
    .X(net470));
 sg13g2_buf_1 _1626_ (.A(net775),
    .X(net471));
 sg13g2_buf_1 _1627_ (.A(net197),
    .X(net472));
 sg13g2_buf_1 _1628_ (.A(net198),
    .X(net473));
 sg13g2_buf_1 _1629_ (.A(net772),
    .X(net474));
 sg13g2_buf_1 _1630_ (.A(net771),
    .X(net475));
 sg13g2_buf_1 _1631_ (.A(net202),
    .X(net477));
 sg13g2_buf_1 _1632_ (.A(net203),
    .X(net478));
 sg13g2_buf_1 _1633_ (.A(net204),
    .X(net479));
 sg13g2_buf_1 _1634_ (.A(net205),
    .X(net480));
 sg13g2_buf_1 _1635_ (.A(net765),
    .X(net481));
 sg13g2_buf_1 _1636_ (.A(net764),
    .X(net482));
 sg13g2_buf_1 _1637_ (.A(net208),
    .X(net483));
 sg13g2_buf_1 _1638_ (.A(net209),
    .X(net484));
 sg13g2_buf_1 _1639_ (.A(net761),
    .X(net485));
 sg13g2_buf_1 _1640_ (.A(net760),
    .X(net486));
 sg13g2_buf_1 _1641_ (.A(net758),
    .X(net488));
 sg13g2_buf_1 _1642_ (.A(net757),
    .X(net489));
 sg13g2_buf_1 _1643_ (.A(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.S1BEG0 ),
    .X(net497));
 sg13g2_buf_1 _1644_ (.A(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.S1BEG1 ),
    .X(net498));
 sg13g2_buf_1 _1645_ (.A(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.S1BEG2 ),
    .X(net499));
 sg13g2_buf_1 _1646_ (.A(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.S1BEG3 ),
    .X(net500));
 sg13g2_buf_1 _1647_ (.A(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.S2BEG0 ),
    .X(net501));
 sg13g2_buf_1 _1648_ (.A(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.S2BEG1 ),
    .X(net502));
 sg13g2_buf_1 _1649_ (.A(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.S2BEG2 ),
    .X(net503));
 sg13g2_buf_1 _1650_ (.A(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.S2BEG3 ),
    .X(net504));
 sg13g2_buf_1 _1651_ (.A(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.S2BEG4 ),
    .X(net505));
 sg13g2_buf_1 _1652_ (.A(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.S2BEG5 ),
    .X(net506));
 sg13g2_buf_1 _1653_ (.A(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.S2BEG6 ),
    .X(net507));
 sg13g2_buf_1 _1654_ (.A(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.S2BEG7 ),
    .X(net508));
 sg13g2_buf_1 _1655_ (.A(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.S2BEG0 ),
    .X(net509));
 sg13g2_buf_1 _1656_ (.A(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.S2BEG1 ),
    .X(net510));
 sg13g2_buf_1 _1657_ (.A(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.S2BEG2 ),
    .X(net511));
 sg13g2_buf_1 _1658_ (.A(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.S2BEG3 ),
    .X(net512));
 sg13g2_buf_1 _1659_ (.A(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.S2BEG4 ),
    .X(net513));
 sg13g2_buf_1 _1660_ (.A(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.S2BEG5 ),
    .X(net514));
 sg13g2_buf_1 _1661_ (.A(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.S2BEG6 ),
    .X(net515));
 sg13g2_buf_1 _1662_ (.A(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.S2BEG7 ),
    .X(net516));
 sg13g2_buf_1 _1663_ (.A(Tile_X0Y0_S4END[8]),
    .X(net517));
 sg13g2_buf_1 _1664_ (.A(Tile_X0Y0_S4END[9]),
    .X(net524));
 sg13g2_buf_1 _1665_ (.A(Tile_X0Y0_S4END[10]),
    .X(net525));
 sg13g2_buf_1 _1666_ (.A(Tile_X0Y0_S4END[11]),
    .X(net526));
 sg13g2_buf_1 _1667_ (.A(Tile_X0Y0_S4END[12]),
    .X(net527));
 sg13g2_buf_1 _1668_ (.A(Tile_X0Y0_S4END[13]),
    .X(net528));
 sg13g2_buf_1 _1669_ (.A(Tile_X0Y0_S4END[14]),
    .X(net529));
 sg13g2_buf_1 _1670_ (.A(Tile_X0Y0_S4END[15]),
    .X(net530));
 sg13g2_buf_1 _1671_ (.A(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.S4BEG0 ),
    .X(net531));
 sg13g2_buf_1 _1672_ (.A(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.S4BEG1 ),
    .X(net532));
 sg13g2_buf_1 _1673_ (.A(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.S4BEG2 ),
    .X(net518));
 sg13g2_buf_1 _1674_ (.A(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.S4BEG3 ),
    .X(net519));
 sg13g2_buf_1 _1675_ (.A(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.S4BEG0 ),
    .X(net520));
 sg13g2_buf_1 _1676_ (.A(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.S4BEG1 ),
    .X(net521));
 sg13g2_buf_1 _1677_ (.A(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.S4BEG2 ),
    .X(net522));
 sg13g2_buf_1 _1678_ (.A(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.S4BEG3 ),
    .X(net523));
 sg13g2_buf_1 _1679_ (.A(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.W1BEG0 ),
    .X(net533));
 sg13g2_buf_1 _1680_ (.A(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.W1BEG1 ),
    .X(net534));
 sg13g2_buf_1 _1681_ (.A(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.W1BEG2 ),
    .X(net535));
 sg13g2_buf_1 _1682_ (.A(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.W1BEG3 ),
    .X(net536));
 sg13g2_buf_1 _1683_ (.A(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.W2BEG0 ),
    .X(net537));
 sg13g2_buf_1 _1684_ (.A(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.W2BEG1 ),
    .X(net538));
 sg13g2_buf_1 _1685_ (.A(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.W2BEG2 ),
    .X(net539));
 sg13g2_buf_1 _1686_ (.A(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.W2BEG3 ),
    .X(net540));
 sg13g2_buf_1 _1687_ (.A(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.W2BEG4 ),
    .X(net541));
 sg13g2_buf_1 _1688_ (.A(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.W2BEG5 ),
    .X(net542));
 sg13g2_buf_1 _1689_ (.A(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.W2BEG6 ),
    .X(net543));
 sg13g2_buf_1 _1690_ (.A(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.W2BEG7 ),
    .X(net544));
 sg13g2_buf_1 _1691_ (.A(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.W2BEGb0 ),
    .X(net545));
 sg13g2_buf_1 _1692_ (.A(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.W2BEGb1 ),
    .X(net546));
 sg13g2_buf_1 _1693_ (.A(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.W2BEGb2 ),
    .X(net547));
 sg13g2_buf_1 _1694_ (.A(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.W2BEGb3 ),
    .X(net548));
 sg13g2_buf_1 _1695_ (.A(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.W2BEGb4 ),
    .X(net549));
 sg13g2_buf_1 _1696_ (.A(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.W2BEGb5 ),
    .X(net550));
 sg13g2_buf_1 _1697_ (.A(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.W2BEGb6 ),
    .X(net551));
 sg13g2_buf_1 _1698_ (.A(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.W2BEGb7 ),
    .X(net552));
 sg13g2_buf_1 _1699_ (.A(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.W6BEG0 ),
    .X(net553));
 sg13g2_buf_1 _1700_ (.A(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.W6BEG1 ),
    .X(net556));
 sg13g2_buf_1 _1701_ (.A(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.W6BEG2 ),
    .X(net557));
 sg13g2_buf_1 _1702_ (.A(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.W6BEG3 ),
    .X(net558));
 sg13g2_buf_1 _1703_ (.A(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.W6BEG4 ),
    .X(net559));
 sg13g2_buf_1 _1704_ (.A(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.W6BEG5 ),
    .X(net560));
 sg13g2_buf_1 _1705_ (.A(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.W6BEG6 ),
    .X(net561));
 sg13g2_buf_1 _1706_ (.A(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.W6BEG7 ),
    .X(net562));
 sg13g2_buf_1 _1707_ (.A(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.W6BEG8 ),
    .X(net563));
 sg13g2_buf_1 _1708_ (.A(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.W6BEG9 ),
    .X(net564));
 sg13g2_buf_1 _1709_ (.A(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.W6BEG10 ),
    .X(net554));
 sg13g2_buf_1 _1710_ (.A(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.W6BEG11 ),
    .X(net555));
 sg13g2_buf_1 _1711_ (.A(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.WW4BEG0 ),
    .X(net565));
 sg13g2_buf_1 _1712_ (.A(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.WW4BEG1 ),
    .X(net572));
 sg13g2_buf_1 _1713_ (.A(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.WW4BEG2 ),
    .X(net573));
 sg13g2_buf_1 _1714_ (.A(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.WW4BEG3 ),
    .X(net574));
 sg13g2_buf_1 _1715_ (.A(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.WW4BEG4 ),
    .X(net575));
 sg13g2_buf_1 _1716_ (.A(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.WW4BEG5 ),
    .X(net576));
 sg13g2_buf_1 _1717_ (.A(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.WW4BEG6 ),
    .X(net577));
 sg13g2_buf_1 _1718_ (.A(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.WW4BEG7 ),
    .X(net578));
 sg13g2_buf_1 _1719_ (.A(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.WW4BEG8 ),
    .X(net579));
 sg13g2_buf_1 _1720_ (.A(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.WW4BEG9 ),
    .X(net580));
 sg13g2_buf_1 _1721_ (.A(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.WW4BEG10 ),
    .X(net566));
 sg13g2_buf_1 _1722_ (.A(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.WW4BEG11 ),
    .X(net567));
 sg13g2_buf_1 _1723_ (.A(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.WW4BEG12 ),
    .X(net568));
 sg13g2_buf_1 _1724_ (.A(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.WW4BEG13 ),
    .X(net569));
 sg13g2_buf_1 _1725_ (.A(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.WW4BEG14 ),
    .X(net570));
 sg13g2_buf_1 _1726_ (.A(\Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.WW4BEG15 ),
    .X(net571));
 sg13g2_buf_1 fanout623 (.A(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS2_BEG7 ),
    .X(net623));
 sg13g2_buf_1 fanout624 (.A(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS2_BEG6 ),
    .X(net624));
 sg13g2_buf_1 fanout625 (.A(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS2_BEG5 ),
    .X(net625));
 sg13g2_buf_1 fanout626 (.A(net627),
    .X(net626));
 sg13g2_buf_1 fanout627 (.A(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS2_BEG4 ),
    .X(net627));
 sg13g2_buf_1 fanout628 (.A(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS2_BEG3 ),
    .X(net628));
 sg13g2_buf_1 fanout629 (.A(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS2_BEG2 ),
    .X(net629));
 sg13g2_buf_1 fanout630 (.A(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS2_BEG1 ),
    .X(net630));
 sg13g2_buf_1 fanout631 (.A(\Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS2_BEG0 ),
    .X(net631));
 sg13g2_buf_1 fanout632 (.A(_0084_),
    .X(net632));
 sg13g2_buf_1 fanout633 (.A(_0083_),
    .X(net633));
 sg13g2_buf_1 fanout634 (.A(_0082_),
    .X(net634));
 sg13g2_buf_1 fanout635 (.A(net636),
    .X(net635));
 sg13g2_buf_1 fanout636 (.A(_0081_),
    .X(net636));
 sg13g2_buf_1 fanout637 (.A(_0080_),
    .X(net637));
 sg13g2_buf_1 fanout638 (.A(_0079_),
    .X(net638));
 sg13g2_buf_1 fanout639 (.A(_0078_),
    .X(net639));
 sg13g2_buf_1 fanout640 (.A(_0043_),
    .X(net640));
 sg13g2_buf_1 fanout641 (.A(net643),
    .X(net641));
 sg13g2_buf_1 fanout642 (.A(net643),
    .X(net642));
 sg13g2_buf_1 fanout643 (.A(net646),
    .X(net643));
 sg13g2_buf_1 fanout644 (.A(net645),
    .X(net644));
 sg13g2_buf_1 fanout645 (.A(net646),
    .X(net645));
 sg13g2_buf_1 fanout646 (.A(Tile_X0Y1_FrameStrobe[9]),
    .X(net646));
 sg13g2_buf_1 fanout647 (.A(net651),
    .X(net647));
 sg13g2_buf_1 fanout648 (.A(net651),
    .X(net648));
 sg13g2_buf_1 fanout649 (.A(net650),
    .X(net649));
 sg13g2_buf_1 fanout650 (.A(net651),
    .X(net650));
 sg13g2_buf_1 fanout651 (.A(net222),
    .X(net651));
 sg13g2_buf_1 fanout652 (.A(net656),
    .X(net652));
 sg13g2_buf_1 fanout653 (.A(net656),
    .X(net653));
 sg13g2_buf_1 fanout654 (.A(net656),
    .X(net654));
 sg13g2_buf_1 fanout655 (.A(net656),
    .X(net655));
 sg13g2_buf_1 fanout656 (.A(net657),
    .X(net656));
 sg13g2_buf_1 fanout657 (.A(net222),
    .X(net657));
 sg13g2_buf_1 fanout658 (.A(net661),
    .X(net658));
 sg13g2_buf_1 fanout659 (.A(net660),
    .X(net659));
 sg13g2_buf_1 fanout660 (.A(net661),
    .X(net660));
 sg13g2_buf_1 fanout661 (.A(net668),
    .X(net661));
 sg13g2_buf_1 fanout662 (.A(net668),
    .X(net662));
 sg13g2_buf_1 fanout663 (.A(net667),
    .X(net663));
 sg13g2_buf_1 fanout664 (.A(net665),
    .X(net664));
 sg13g2_buf_1 fanout665 (.A(net667),
    .X(net665));
 sg13g2_buf_1 fanout666 (.A(net667),
    .X(net666));
 sg13g2_buf_1 fanout667 (.A(net668),
    .X(net667));
 sg13g2_buf_1 fanout668 (.A(Tile_X0Y1_FrameStrobe[7]),
    .X(net668));
 sg13g2_buf_1 fanout669 (.A(net672),
    .X(net669));
 sg13g2_buf_1 fanout670 (.A(net672),
    .X(net670));
 sg13g2_buf_1 fanout671 (.A(net672),
    .X(net671));
 sg13g2_buf_1 fanout672 (.A(net673),
    .X(net672));
 sg13g2_buf_1 fanout673 (.A(net674),
    .X(net673));
 sg13g2_buf_1 fanout674 (.A(Tile_X0Y1_FrameStrobe[6]),
    .X(net674));
 sg13g2_buf_1 fanout675 (.A(net677),
    .X(net675));
 sg13g2_buf_1 fanout676 (.A(net677),
    .X(net676));
 sg13g2_buf_1 fanout677 (.A(net678),
    .X(net677));
 sg13g2_buf_1 fanout678 (.A(Tile_X0Y1_FrameStrobe[6]),
    .X(net678));
 sg13g2_buf_1 fanout679 (.A(Tile_X0Y1_FrameStrobe[6]),
    .X(net679));
 sg13g2_buf_1 fanout680 (.A(net681),
    .X(net680));
 sg13g2_buf_1 fanout681 (.A(net684),
    .X(net681));
 sg13g2_buf_1 fanout682 (.A(net684),
    .X(net682));
 sg13g2_buf_1 fanout683 (.A(net684),
    .X(net683));
 sg13g2_buf_1 fanout684 (.A(net691),
    .X(net684));
 sg13g2_buf_1 fanout685 (.A(net689),
    .X(net685));
 sg13g2_buf_1 fanout686 (.A(net689),
    .X(net686));
 sg13g2_buf_1 fanout687 (.A(net689),
    .X(net687));
 sg13g2_buf_1 fanout688 (.A(net689),
    .X(net688));
 sg13g2_buf_1 fanout689 (.A(net690),
    .X(net689));
 sg13g2_buf_1 fanout690 (.A(net691),
    .X(net690));
 sg13g2_buf_1 fanout691 (.A(Tile_X0Y1_FrameStrobe[5]),
    .X(net691));
 sg13g2_buf_1 fanout692 (.A(net693),
    .X(net692));
 sg13g2_buf_1 fanout693 (.A(net695),
    .X(net693));
 sg13g2_buf_1 fanout694 (.A(net695),
    .X(net694));
 sg13g2_buf_1 fanout695 (.A(net696),
    .X(net695));
 sg13g2_buf_1 fanout696 (.A(Tile_X0Y1_FrameStrobe[4]),
    .X(net696));
 sg13g2_buf_1 fanout697 (.A(net699),
    .X(net697));
 sg13g2_buf_1 fanout698 (.A(net699),
    .X(net698));
 sg13g2_buf_1 fanout699 (.A(net702),
    .X(net699));
 sg13g2_buf_1 fanout700 (.A(net701),
    .X(net700));
 sg13g2_buf_1 fanout701 (.A(net702),
    .X(net701));
 sg13g2_buf_1 fanout702 (.A(Tile_X0Y1_FrameStrobe[4]),
    .X(net702));
 sg13g2_buf_1 fanout703 (.A(net705),
    .X(net703));
 sg13g2_buf_1 fanout704 (.A(net705),
    .X(net704));
 sg13g2_buf_1 fanout705 (.A(net708),
    .X(net705));
 sg13g2_buf_1 fanout706 (.A(net708),
    .X(net706));
 sg13g2_buf_1 fanout707 (.A(net708),
    .X(net707));
 sg13g2_buf_1 fanout708 (.A(Tile_X0Y1_FrameStrobe[3]),
    .X(net708));
 sg13g2_buf_1 fanout709 (.A(net713),
    .X(net709));
 sg13g2_buf_1 fanout710 (.A(net713),
    .X(net710));
 sg13g2_buf_1 fanout711 (.A(net713),
    .X(net711));
 sg13g2_buf_1 fanout712 (.A(net713),
    .X(net712));
 sg13g2_buf_1 fanout713 (.A(Tile_X0Y1_FrameStrobe[3]),
    .X(net713));
 sg13g2_buf_1 fanout714 (.A(net715),
    .X(net714));
 sg13g2_buf_1 fanout715 (.A(net716),
    .X(net715));
 sg13g2_buf_1 fanout716 (.A(net719),
    .X(net716));
 sg13g2_buf_1 fanout717 (.A(net718),
    .X(net717));
 sg13g2_buf_1 fanout718 (.A(net719),
    .X(net718));
 sg13g2_buf_1 fanout719 (.A(net724),
    .X(net719));
 sg13g2_buf_1 fanout720 (.A(net724),
    .X(net720));
 sg13g2_buf_1 fanout721 (.A(net724),
    .X(net721));
 sg13g2_buf_1 fanout722 (.A(net724),
    .X(net722));
 sg13g2_buf_1 fanout723 (.A(net724),
    .X(net723));
 sg13g2_buf_1 fanout724 (.A(Tile_X0Y1_FrameStrobe[2]),
    .X(net724));
 sg13g2_buf_1 fanout725 (.A(net727),
    .X(net725));
 sg13g2_buf_1 fanout726 (.A(net727),
    .X(net726));
 sg13g2_buf_1 fanout727 (.A(net737),
    .X(net727));
 sg13g2_buf_1 fanout728 (.A(net730),
    .X(net728));
 sg13g2_buf_1 fanout729 (.A(net730),
    .X(net729));
 sg13g2_buf_1 fanout730 (.A(net737),
    .X(net730));
 sg13g2_buf_1 fanout731 (.A(net737),
    .X(net731));
 sg13g2_buf_1 fanout732 (.A(net736),
    .X(net732));
 sg13g2_buf_1 fanout733 (.A(net736),
    .X(net733));
 sg13g2_buf_1 fanout734 (.A(net736),
    .X(net734));
 sg13g2_buf_1 fanout735 (.A(net736),
    .X(net735));
 sg13g2_buf_1 fanout736 (.A(net737),
    .X(net736));
 sg13g2_buf_1 fanout737 (.A(Tile_X0Y1_FrameStrobe[1]),
    .X(net737));
 sg13g2_buf_1 fanout738 (.A(net749),
    .X(net738));
 sg13g2_buf_1 fanout739 (.A(net749),
    .X(net739));
 sg13g2_buf_1 fanout740 (.A(net741),
    .X(net740));
 sg13g2_buf_1 fanout741 (.A(net742),
    .X(net741));
 sg13g2_buf_1 fanout742 (.A(net749),
    .X(net742));
 sg13g2_buf_1 fanout743 (.A(net748),
    .X(net743));
 sg13g2_buf_1 fanout744 (.A(net747),
    .X(net744));
 sg13g2_buf_1 fanout745 (.A(net747),
    .X(net745));
 sg13g2_buf_1 fanout746 (.A(net747),
    .X(net746));
 sg13g2_buf_1 fanout747 (.A(net748),
    .X(net747));
 sg13g2_buf_1 fanout748 (.A(net749),
    .X(net748));
 sg13g2_buf_1 fanout749 (.A(Tile_X0Y1_FrameStrobe[0]),
    .X(net749));
 sg13g2_buf_1 fanout750 (.A(net221),
    .X(net750));
 sg13g2_buf_1 fanout751 (.A(net220),
    .X(net751));
 sg13g2_buf_1 fanout752 (.A(net219),
    .X(net752));
 sg13g2_buf_1 fanout753 (.A(net218),
    .X(net753));
 sg13g2_buf_1 fanout754 (.A(net217),
    .X(net754));
 sg13g2_buf_1 fanout755 (.A(net216),
    .X(net755));
 sg13g2_buf_1 fanout756 (.A(net215),
    .X(net756));
 sg13g2_buf_1 fanout757 (.A(net214),
    .X(net757));
 sg13g2_buf_1 fanout758 (.A(net213),
    .X(net758));
 sg13g2_buf_1 fanout759 (.A(net212),
    .X(net759));
 sg13g2_buf_1 fanout760 (.A(net211),
    .X(net760));
 sg13g2_buf_1 fanout761 (.A(net210),
    .X(net761));
 sg13g2_buf_1 fanout762 (.A(net209),
    .X(net762));
 sg13g2_buf_1 fanout763 (.A(net208),
    .X(net763));
 sg13g2_buf_1 fanout764 (.A(net207),
    .X(net764));
 sg13g2_buf_1 fanout765 (.A(net206),
    .X(net765));
 sg13g2_buf_1 fanout766 (.A(net205),
    .X(net766));
 sg13g2_buf_1 fanout767 (.A(net204),
    .X(net767));
 sg13g2_buf_1 fanout768 (.A(net203),
    .X(net768));
 sg13g2_buf_1 fanout769 (.A(net202),
    .X(net769));
 sg13g2_buf_1 fanout770 (.A(net201),
    .X(net770));
 sg13g2_buf_1 fanout771 (.A(net200),
    .X(net771));
 sg13g2_buf_1 fanout772 (.A(net199),
    .X(net772));
 sg13g2_buf_1 fanout773 (.A(net198),
    .X(net773));
 sg13g2_buf_1 fanout774 (.A(net197),
    .X(net774));
 sg13g2_buf_1 fanout775 (.A(net196),
    .X(net775));
 sg13g2_buf_1 fanout776 (.A(net195),
    .X(net776));
 sg13g2_buf_1 fanout777 (.A(net194),
    .X(net777));
 sg13g2_buf_1 fanout778 (.A(net193),
    .X(net778));
 sg13g2_buf_1 fanout779 (.A(net192),
    .X(net779));
 sg13g2_buf_1 fanout780 (.A(net191),
    .X(net780));
 sg13g2_buf_1 fanout781 (.A(net190),
    .X(net781));
 sg13g2_buf_1 fanout782 (.A(net113),
    .X(net782));
 sg13g2_buf_1 fanout783 (.A(net112),
    .X(net783));
 sg13g2_buf_1 fanout784 (.A(net111),
    .X(net784));
 sg13g2_buf_1 fanout785 (.A(net110),
    .X(net785));
 sg13g2_buf_1 fanout786 (.A(net109),
    .X(net786));
 sg13g2_buf_1 fanout787 (.A(net108),
    .X(net787));
 sg13g2_buf_1 fanout788 (.A(net107),
    .X(net788));
 sg13g2_buf_1 fanout789 (.A(net106),
    .X(net789));
 sg13g2_buf_1 fanout790 (.A(net105),
    .X(net790));
 sg13g2_buf_1 fanout791 (.A(net104),
    .X(net791));
 sg13g2_buf_1 fanout792 (.A(net103),
    .X(net792));
 sg13g2_buf_1 fanout793 (.A(net102),
    .X(net793));
 sg13g2_buf_1 fanout794 (.A(net101),
    .X(net794));
 sg13g2_buf_1 fanout795 (.A(net100),
    .X(net795));
 sg13g2_buf_1 fanout796 (.A(net99),
    .X(net796));
 sg13g2_buf_1 fanout797 (.A(net98),
    .X(net797));
 sg13g2_buf_1 fanout798 (.A(net97),
    .X(net798));
 sg13g2_buf_1 fanout799 (.A(net96),
    .X(net799));
 sg13g2_buf_1 fanout800 (.A(net95),
    .X(net800));
 sg13g2_buf_1 fanout801 (.A(net94),
    .X(net801));
 sg13g2_buf_1 fanout802 (.A(net93),
    .X(net802));
 sg13g2_buf_1 fanout803 (.A(net92),
    .X(net803));
 sg13g2_buf_1 fanout804 (.A(net91),
    .X(net804));
 sg13g2_buf_1 fanout805 (.A(net90),
    .X(net805));
 sg13g2_buf_1 fanout806 (.A(net89),
    .X(net806));
 sg13g2_buf_1 fanout807 (.A(net88),
    .X(net807));
 sg13g2_buf_1 fanout808 (.A(net87),
    .X(net808));
 sg13g2_buf_1 fanout809 (.A(net86),
    .X(net809));
 sg13g2_buf_1 fanout810 (.A(net85),
    .X(net810));
 sg13g2_buf_1 fanout811 (.A(net84),
    .X(net811));
 sg13g2_buf_1 fanout812 (.A(net83),
    .X(net812));
 sg13g2_buf_1 fanout813 (.A(net82),
    .X(net813));
 sg13g2_buf_1 input1 (.A(CONFIGURED_top),
    .X(net1));
 sg13g2_buf_1 input2 (.A(DOUT_SRAM0),
    .X(net2));
 sg13g2_buf_1 input3 (.A(DOUT_SRAM1),
    .X(net3));
 sg13g2_buf_1 input4 (.A(DOUT_SRAM10),
    .X(net4));
 sg13g2_buf_1 input5 (.A(DOUT_SRAM11),
    .X(net5));
 sg13g2_buf_1 input6 (.A(DOUT_SRAM12),
    .X(net6));
 sg13g2_buf_1 input7 (.A(DOUT_SRAM13),
    .X(net7));
 sg13g2_buf_1 input8 (.A(DOUT_SRAM14),
    .X(net8));
 sg13g2_buf_1 input9 (.A(DOUT_SRAM15),
    .X(net9));
 sg13g2_buf_1 input10 (.A(DOUT_SRAM16),
    .X(net10));
 sg13g2_buf_1 input11 (.A(DOUT_SRAM17),
    .X(net11));
 sg13g2_buf_1 input12 (.A(DOUT_SRAM18),
    .X(net12));
 sg13g2_buf_1 input13 (.A(DOUT_SRAM19),
    .X(net13));
 sg13g2_buf_1 input14 (.A(DOUT_SRAM2),
    .X(net14));
 sg13g2_buf_1 input15 (.A(DOUT_SRAM20),
    .X(net15));
 sg13g2_buf_1 input16 (.A(DOUT_SRAM21),
    .X(net16));
 sg13g2_buf_1 input17 (.A(DOUT_SRAM22),
    .X(net17));
 sg13g2_buf_1 input18 (.A(DOUT_SRAM23),
    .X(net18));
 sg13g2_buf_1 input19 (.A(DOUT_SRAM24),
    .X(net19));
 sg13g2_buf_1 input20 (.A(DOUT_SRAM25),
    .X(net20));
 sg13g2_buf_1 input21 (.A(DOUT_SRAM26),
    .X(net21));
 sg13g2_buf_1 input22 (.A(DOUT_SRAM27),
    .X(net22));
 sg13g2_buf_1 input23 (.A(DOUT_SRAM28),
    .X(net23));
 sg13g2_buf_1 input24 (.A(DOUT_SRAM29),
    .X(net24));
 sg13g2_buf_1 input25 (.A(DOUT_SRAM3),
    .X(net25));
 sg13g2_buf_1 input26 (.A(DOUT_SRAM30),
    .X(net26));
 sg13g2_buf_1 input27 (.A(DOUT_SRAM31),
    .X(net27));
 sg13g2_buf_1 input28 (.A(DOUT_SRAM4),
    .X(net28));
 sg13g2_buf_1 input29 (.A(DOUT_SRAM5),
    .X(net29));
 sg13g2_buf_1 input30 (.A(DOUT_SRAM6),
    .X(net30));
 sg13g2_buf_1 input31 (.A(DOUT_SRAM7),
    .X(net31));
 sg13g2_buf_1 input32 (.A(DOUT_SRAM8),
    .X(net32));
 sg13g2_buf_1 input33 (.A(DOUT_SRAM9),
    .X(net33));
 sg13g2_buf_1 input34 (.A(Tile_X0Y0_E1END[0]),
    .X(net34));
 sg13g2_buf_1 input35 (.A(Tile_X0Y0_E1END[1]),
    .X(net35));
 sg13g2_buf_1 input36 (.A(Tile_X0Y0_E1END[2]),
    .X(net36));
 sg13g2_buf_1 input37 (.A(Tile_X0Y0_E1END[3]),
    .X(net37));
 sg13g2_buf_1 input38 (.A(Tile_X0Y0_E2END[0]),
    .X(net38));
 sg13g2_buf_1 input39 (.A(Tile_X0Y0_E2END[1]),
    .X(net39));
 sg13g2_buf_1 input40 (.A(Tile_X0Y0_E2END[2]),
    .X(net40));
 sg13g2_buf_1 input41 (.A(Tile_X0Y0_E2END[3]),
    .X(net41));
 sg13g2_buf_1 input42 (.A(Tile_X0Y0_E2END[4]),
    .X(net42));
 sg13g2_buf_1 input43 (.A(Tile_X0Y0_E2END[5]),
    .X(net43));
 sg13g2_buf_1 input44 (.A(Tile_X0Y0_E2END[6]),
    .X(net44));
 sg13g2_buf_1 input45 (.A(Tile_X0Y0_E2END[7]),
    .X(net45));
 sg13g2_buf_1 input46 (.A(Tile_X0Y0_E2MID[0]),
    .X(net46));
 sg13g2_buf_1 input47 (.A(Tile_X0Y0_E2MID[1]),
    .X(net47));
 sg13g2_buf_1 input48 (.A(Tile_X0Y0_E2MID[2]),
    .X(net48));
 sg13g2_buf_1 input49 (.A(Tile_X0Y0_E2MID[3]),
    .X(net49));
 sg13g2_buf_1 input50 (.A(Tile_X0Y0_E2MID[4]),
    .X(net50));
 sg13g2_buf_1 input51 (.A(Tile_X0Y0_E2MID[5]),
    .X(net51));
 sg13g2_buf_1 input52 (.A(Tile_X0Y0_E2MID[6]),
    .X(net52));
 sg13g2_buf_1 input53 (.A(Tile_X0Y0_E2MID[7]),
    .X(net53));
 sg13g2_buf_1 input54 (.A(Tile_X0Y0_E6END[0]),
    .X(net54));
 sg13g2_buf_1 input55 (.A(Tile_X0Y0_E6END[10]),
    .X(net55));
 sg13g2_buf_1 input56 (.A(Tile_X0Y0_E6END[11]),
    .X(net56));
 sg13g2_buf_1 input57 (.A(Tile_X0Y0_E6END[1]),
    .X(net57));
 sg13g2_buf_1 input58 (.A(Tile_X0Y0_E6END[2]),
    .X(net58));
 sg13g2_buf_1 input59 (.A(Tile_X0Y0_E6END[3]),
    .X(net59));
 sg13g2_buf_1 input60 (.A(Tile_X0Y0_E6END[4]),
    .X(net60));
 sg13g2_buf_1 input61 (.A(Tile_X0Y0_E6END[5]),
    .X(net61));
 sg13g2_buf_1 input62 (.A(Tile_X0Y0_E6END[6]),
    .X(net62));
 sg13g2_buf_1 input63 (.A(Tile_X0Y0_E6END[7]),
    .X(net63));
 sg13g2_buf_1 input64 (.A(Tile_X0Y0_E6END[8]),
    .X(net64));
 sg13g2_buf_1 input65 (.A(Tile_X0Y0_E6END[9]),
    .X(net65));
 sg13g2_buf_1 input66 (.A(Tile_X0Y0_EE4END[0]),
    .X(net66));
 sg13g2_buf_1 input67 (.A(Tile_X0Y0_EE4END[10]),
    .X(net67));
 sg13g2_buf_1 input68 (.A(Tile_X0Y0_EE4END[11]),
    .X(net68));
 sg13g2_buf_1 input69 (.A(Tile_X0Y0_EE4END[12]),
    .X(net69));
 sg13g2_buf_1 input70 (.A(Tile_X0Y0_EE4END[13]),
    .X(net70));
 sg13g2_buf_1 input71 (.A(Tile_X0Y0_EE4END[14]),
    .X(net71));
 sg13g2_buf_1 input72 (.A(Tile_X0Y0_EE4END[15]),
    .X(net72));
 sg13g2_buf_1 input73 (.A(Tile_X0Y0_EE4END[1]),
    .X(net73));
 sg13g2_buf_1 input74 (.A(Tile_X0Y0_EE4END[2]),
    .X(net74));
 sg13g2_buf_1 input75 (.A(Tile_X0Y0_EE4END[3]),
    .X(net75));
 sg13g2_buf_1 input76 (.A(Tile_X0Y0_EE4END[4]),
    .X(net76));
 sg13g2_buf_1 input77 (.A(Tile_X0Y0_EE4END[5]),
    .X(net77));
 sg13g2_buf_1 input78 (.A(Tile_X0Y0_EE4END[6]),
    .X(net78));
 sg13g2_buf_1 input79 (.A(Tile_X0Y0_EE4END[7]),
    .X(net79));
 sg13g2_buf_1 input80 (.A(Tile_X0Y0_EE4END[8]),
    .X(net80));
 sg13g2_buf_1 input81 (.A(Tile_X0Y0_EE4END[9]),
    .X(net81));
 sg13g2_buf_1 input82 (.A(Tile_X0Y0_FrameData[0]),
    .X(net82));
 sg13g2_buf_1 input83 (.A(Tile_X0Y0_FrameData[10]),
    .X(net83));
 sg13g2_buf_1 input84 (.A(Tile_X0Y0_FrameData[11]),
    .X(net84));
 sg13g2_buf_1 input85 (.A(Tile_X0Y0_FrameData[12]),
    .X(net85));
 sg13g2_buf_1 input86 (.A(Tile_X0Y0_FrameData[13]),
    .X(net86));
 sg13g2_buf_1 input87 (.A(Tile_X0Y0_FrameData[14]),
    .X(net87));
 sg13g2_buf_1 input88 (.A(Tile_X0Y0_FrameData[15]),
    .X(net88));
 sg13g2_buf_1 input89 (.A(Tile_X0Y0_FrameData[16]),
    .X(net89));
 sg13g2_buf_1 input90 (.A(Tile_X0Y0_FrameData[17]),
    .X(net90));
 sg13g2_buf_1 input91 (.A(Tile_X0Y0_FrameData[18]),
    .X(net91));
 sg13g2_buf_1 input92 (.A(Tile_X0Y0_FrameData[19]),
    .X(net92));
 sg13g2_buf_1 input93 (.A(Tile_X0Y0_FrameData[1]),
    .X(net93));
 sg13g2_buf_1 input94 (.A(Tile_X0Y0_FrameData[20]),
    .X(net94));
 sg13g2_buf_1 input95 (.A(Tile_X0Y0_FrameData[21]),
    .X(net95));
 sg13g2_buf_1 input96 (.A(Tile_X0Y0_FrameData[22]),
    .X(net96));
 sg13g2_buf_1 input97 (.A(Tile_X0Y0_FrameData[23]),
    .X(net97));
 sg13g2_buf_1 input98 (.A(Tile_X0Y0_FrameData[24]),
    .X(net98));
 sg13g2_buf_1 input99 (.A(Tile_X0Y0_FrameData[25]),
    .X(net99));
 sg13g2_buf_1 input100 (.A(Tile_X0Y0_FrameData[26]),
    .X(net100));
 sg13g2_buf_1 input101 (.A(Tile_X0Y0_FrameData[27]),
    .X(net101));
 sg13g2_buf_1 input102 (.A(Tile_X0Y0_FrameData[28]),
    .X(net102));
 sg13g2_buf_1 input103 (.A(Tile_X0Y0_FrameData[29]),
    .X(net103));
 sg13g2_buf_1 input104 (.A(Tile_X0Y0_FrameData[2]),
    .X(net104));
 sg13g2_buf_1 input105 (.A(Tile_X0Y0_FrameData[30]),
    .X(net105));
 sg13g2_buf_1 input106 (.A(Tile_X0Y0_FrameData[31]),
    .X(net106));
 sg13g2_buf_1 input107 (.A(Tile_X0Y0_FrameData[3]),
    .X(net107));
 sg13g2_buf_1 input108 (.A(Tile_X0Y0_FrameData[4]),
    .X(net108));
 sg13g2_buf_1 input109 (.A(Tile_X0Y0_FrameData[5]),
    .X(net109));
 sg13g2_buf_1 input110 (.A(Tile_X0Y0_FrameData[6]),
    .X(net110));
 sg13g2_buf_1 input111 (.A(Tile_X0Y0_FrameData[7]),
    .X(net111));
 sg13g2_buf_1 input112 (.A(Tile_X0Y0_FrameData[8]),
    .X(net112));
 sg13g2_buf_1 input113 (.A(Tile_X0Y0_FrameData[9]),
    .X(net113));
 sg13g2_buf_1 input114 (.A(Tile_X0Y0_S1END[0]),
    .X(net114));
 sg13g2_buf_1 input115 (.A(Tile_X0Y0_S1END[1]),
    .X(net115));
 sg13g2_buf_1 input116 (.A(Tile_X0Y0_S1END[2]),
    .X(net116));
 sg13g2_buf_1 input117 (.A(Tile_X0Y0_S1END[3]),
    .X(net117));
 sg13g2_buf_1 input118 (.A(Tile_X0Y0_S2END[0]),
    .X(net118));
 sg13g2_buf_1 input119 (.A(Tile_X0Y0_S2END[1]),
    .X(net119));
 sg13g2_buf_1 input120 (.A(Tile_X0Y0_S2END[2]),
    .X(net120));
 sg13g2_buf_1 input121 (.A(Tile_X0Y0_S2END[3]),
    .X(net121));
 sg13g2_buf_1 input122 (.A(Tile_X0Y0_S2END[4]),
    .X(net122));
 sg13g2_buf_1 input123 (.A(Tile_X0Y0_S2END[5]),
    .X(net123));
 sg13g2_buf_1 input124 (.A(Tile_X0Y0_S2END[6]),
    .X(net124));
 sg13g2_buf_1 input125 (.A(Tile_X0Y0_S2END[7]),
    .X(net125));
 sg13g2_buf_1 input126 (.A(Tile_X0Y0_S2MID[0]),
    .X(net126));
 sg13g2_buf_1 input127 (.A(Tile_X0Y0_S2MID[1]),
    .X(net127));
 sg13g2_buf_1 input128 (.A(Tile_X0Y0_S2MID[2]),
    .X(net128));
 sg13g2_buf_1 input129 (.A(Tile_X0Y0_S2MID[3]),
    .X(net129));
 sg13g2_buf_1 input130 (.A(Tile_X0Y0_S2MID[4]),
    .X(net130));
 sg13g2_buf_1 input131 (.A(Tile_X0Y0_S2MID[5]),
    .X(net131));
 sg13g2_buf_1 input132 (.A(Tile_X0Y0_S2MID[6]),
    .X(net132));
 sg13g2_buf_1 input133 (.A(Tile_X0Y0_S2MID[7]),
    .X(net133));
 sg13g2_buf_1 input134 (.A(Tile_X0Y0_S4END[0]),
    .X(net134));
 sg13g2_buf_1 input135 (.A(Tile_X0Y0_S4END[1]),
    .X(net135));
 sg13g2_buf_1 input136 (.A(Tile_X0Y0_S4END[2]),
    .X(net136));
 sg13g2_buf_1 input137 (.A(Tile_X0Y0_S4END[3]),
    .X(net137));
 sg13g2_buf_1 input138 (.A(Tile_X0Y0_S4END[4]),
    .X(net138));
 sg13g2_buf_1 input139 (.A(Tile_X0Y0_S4END[5]),
    .X(net139));
 sg13g2_buf_1 input140 (.A(Tile_X0Y0_S4END[6]),
    .X(net140));
 sg13g2_buf_1 input141 (.A(Tile_X0Y0_S4END[7]),
    .X(net141));
 sg13g2_buf_1 input142 (.A(Tile_X0Y1_E1END[0]),
    .X(net142));
 sg13g2_buf_1 input143 (.A(Tile_X0Y1_E1END[1]),
    .X(net143));
 sg13g2_buf_1 input144 (.A(Tile_X0Y1_E1END[2]),
    .X(net144));
 sg13g2_buf_1 input145 (.A(Tile_X0Y1_E1END[3]),
    .X(net145));
 sg13g2_buf_1 input146 (.A(Tile_X0Y1_E2END[0]),
    .X(net146));
 sg13g2_buf_1 input147 (.A(Tile_X0Y1_E2END[1]),
    .X(net147));
 sg13g2_buf_1 input148 (.A(Tile_X0Y1_E2END[2]),
    .X(net148));
 sg13g2_buf_1 input149 (.A(Tile_X0Y1_E2END[3]),
    .X(net149));
 sg13g2_buf_1 input150 (.A(Tile_X0Y1_E2END[4]),
    .X(net150));
 sg13g2_buf_1 input151 (.A(Tile_X0Y1_E2END[5]),
    .X(net151));
 sg13g2_buf_1 input152 (.A(Tile_X0Y1_E2END[6]),
    .X(net152));
 sg13g2_buf_1 input153 (.A(Tile_X0Y1_E2END[7]),
    .X(net153));
 sg13g2_buf_1 input154 (.A(Tile_X0Y1_E2MID[0]),
    .X(net154));
 sg13g2_buf_1 input155 (.A(Tile_X0Y1_E2MID[1]),
    .X(net155));
 sg13g2_buf_1 input156 (.A(Tile_X0Y1_E2MID[2]),
    .X(net156));
 sg13g2_buf_1 input157 (.A(Tile_X0Y1_E2MID[3]),
    .X(net157));
 sg13g2_buf_1 input158 (.A(Tile_X0Y1_E2MID[4]),
    .X(net158));
 sg13g2_buf_1 input159 (.A(Tile_X0Y1_E2MID[5]),
    .X(net159));
 sg13g2_buf_1 input160 (.A(Tile_X0Y1_E2MID[6]),
    .X(net160));
 sg13g2_buf_1 input161 (.A(Tile_X0Y1_E2MID[7]),
    .X(net161));
 sg13g2_buf_1 input162 (.A(Tile_X0Y1_E6END[0]),
    .X(net162));
 sg13g2_buf_1 input163 (.A(Tile_X0Y1_E6END[10]),
    .X(net163));
 sg13g2_buf_1 input164 (.A(Tile_X0Y1_E6END[11]),
    .X(net164));
 sg13g2_buf_1 input165 (.A(Tile_X0Y1_E6END[1]),
    .X(net165));
 sg13g2_buf_1 input166 (.A(Tile_X0Y1_E6END[2]),
    .X(net166));
 sg13g2_buf_1 input167 (.A(Tile_X0Y1_E6END[3]),
    .X(net167));
 sg13g2_buf_1 input168 (.A(Tile_X0Y1_E6END[4]),
    .X(net168));
 sg13g2_buf_1 input169 (.A(Tile_X0Y1_E6END[5]),
    .X(net169));
 sg13g2_buf_1 input170 (.A(Tile_X0Y1_E6END[6]),
    .X(net170));
 sg13g2_buf_1 input171 (.A(Tile_X0Y1_E6END[7]),
    .X(net171));
 sg13g2_buf_1 input172 (.A(Tile_X0Y1_E6END[8]),
    .X(net172));
 sg13g2_buf_1 input173 (.A(Tile_X0Y1_E6END[9]),
    .X(net173));
 sg13g2_buf_1 input174 (.A(Tile_X0Y1_EE4END[0]),
    .X(net174));
 sg13g2_buf_1 input175 (.A(Tile_X0Y1_EE4END[10]),
    .X(net175));
 sg13g2_buf_1 input176 (.A(Tile_X0Y1_EE4END[11]),
    .X(net176));
 sg13g2_buf_1 input177 (.A(Tile_X0Y1_EE4END[12]),
    .X(net177));
 sg13g2_buf_1 input178 (.A(Tile_X0Y1_EE4END[13]),
    .X(net178));
 sg13g2_buf_1 input179 (.A(Tile_X0Y1_EE4END[14]),
    .X(net179));
 sg13g2_buf_1 input180 (.A(Tile_X0Y1_EE4END[15]),
    .X(net180));
 sg13g2_buf_1 input181 (.A(Tile_X0Y1_EE4END[1]),
    .X(net181));
 sg13g2_buf_1 input182 (.A(Tile_X0Y1_EE4END[2]),
    .X(net182));
 sg13g2_buf_1 input183 (.A(Tile_X0Y1_EE4END[3]),
    .X(net183));
 sg13g2_buf_1 input184 (.A(Tile_X0Y1_EE4END[4]),
    .X(net184));
 sg13g2_buf_1 input185 (.A(Tile_X0Y1_EE4END[5]),
    .X(net185));
 sg13g2_buf_1 input186 (.A(Tile_X0Y1_EE4END[6]),
    .X(net186));
 sg13g2_buf_1 input187 (.A(Tile_X0Y1_EE4END[7]),
    .X(net187));
 sg13g2_buf_1 input188 (.A(Tile_X0Y1_EE4END[8]),
    .X(net188));
 sg13g2_buf_1 input189 (.A(Tile_X0Y1_EE4END[9]),
    .X(net189));
 sg13g2_buf_1 input190 (.A(Tile_X0Y1_FrameData[0]),
    .X(net190));
 sg13g2_buf_1 input191 (.A(Tile_X0Y1_FrameData[10]),
    .X(net191));
 sg13g2_buf_1 input192 (.A(Tile_X0Y1_FrameData[11]),
    .X(net192));
 sg13g2_buf_1 input193 (.A(Tile_X0Y1_FrameData[12]),
    .X(net193));
 sg13g2_buf_1 input194 (.A(Tile_X0Y1_FrameData[13]),
    .X(net194));
 sg13g2_buf_1 input195 (.A(Tile_X0Y1_FrameData[14]),
    .X(net195));
 sg13g2_buf_1 input196 (.A(Tile_X0Y1_FrameData[15]),
    .X(net196));
 sg13g2_buf_1 input197 (.A(Tile_X0Y1_FrameData[16]),
    .X(net197));
 sg13g2_buf_1 input198 (.A(Tile_X0Y1_FrameData[17]),
    .X(net198));
 sg13g2_buf_1 input199 (.A(Tile_X0Y1_FrameData[18]),
    .X(net199));
 sg13g2_buf_1 input200 (.A(Tile_X0Y1_FrameData[19]),
    .X(net200));
 sg13g2_buf_1 input201 (.A(Tile_X0Y1_FrameData[1]),
    .X(net201));
 sg13g2_buf_1 input202 (.A(Tile_X0Y1_FrameData[20]),
    .X(net202));
 sg13g2_buf_1 input203 (.A(Tile_X0Y1_FrameData[21]),
    .X(net203));
 sg13g2_buf_1 input204 (.A(Tile_X0Y1_FrameData[22]),
    .X(net204));
 sg13g2_buf_1 input205 (.A(Tile_X0Y1_FrameData[23]),
    .X(net205));
 sg13g2_buf_1 input206 (.A(Tile_X0Y1_FrameData[24]),
    .X(net206));
 sg13g2_buf_1 input207 (.A(Tile_X0Y1_FrameData[25]),
    .X(net207));
 sg13g2_buf_1 input208 (.A(Tile_X0Y1_FrameData[26]),
    .X(net208));
 sg13g2_buf_1 input209 (.A(Tile_X0Y1_FrameData[27]),
    .X(net209));
 sg13g2_buf_1 input210 (.A(Tile_X0Y1_FrameData[28]),
    .X(net210));
 sg13g2_buf_1 input211 (.A(Tile_X0Y1_FrameData[29]),
    .X(net211));
 sg13g2_buf_1 input212 (.A(Tile_X0Y1_FrameData[2]),
    .X(net212));
 sg13g2_buf_1 input213 (.A(Tile_X0Y1_FrameData[30]),
    .X(net213));
 sg13g2_buf_1 input214 (.A(Tile_X0Y1_FrameData[31]),
    .X(net214));
 sg13g2_buf_1 input215 (.A(Tile_X0Y1_FrameData[3]),
    .X(net215));
 sg13g2_buf_1 input216 (.A(Tile_X0Y1_FrameData[4]),
    .X(net216));
 sg13g2_buf_1 input217 (.A(Tile_X0Y1_FrameData[5]),
    .X(net217));
 sg13g2_buf_1 input218 (.A(Tile_X0Y1_FrameData[6]),
    .X(net218));
 sg13g2_buf_1 input219 (.A(Tile_X0Y1_FrameData[7]),
    .X(net219));
 sg13g2_buf_1 input220 (.A(Tile_X0Y1_FrameData[8]),
    .X(net220));
 sg13g2_buf_1 input221 (.A(Tile_X0Y1_FrameData[9]),
    .X(net221));
 sg13g2_buf_1 input222 (.A(Tile_X0Y1_FrameStrobe[8]),
    .X(net222));
 sg13g2_buf_1 input223 (.A(Tile_X0Y1_N1END[0]),
    .X(net223));
 sg13g2_buf_1 input224 (.A(Tile_X0Y1_N1END[1]),
    .X(net224));
 sg13g2_buf_1 input225 (.A(Tile_X0Y1_N1END[2]),
    .X(net225));
 sg13g2_buf_1 input226 (.A(Tile_X0Y1_N1END[3]),
    .X(net226));
 sg13g2_buf_1 input227 (.A(Tile_X0Y1_N2END[0]),
    .X(net227));
 sg13g2_buf_1 input228 (.A(Tile_X0Y1_N2END[1]),
    .X(net228));
 sg13g2_buf_1 input229 (.A(Tile_X0Y1_N2END[2]),
    .X(net229));
 sg13g2_buf_1 input230 (.A(Tile_X0Y1_N2END[3]),
    .X(net230));
 sg13g2_buf_1 input231 (.A(Tile_X0Y1_N2END[4]),
    .X(net231));
 sg13g2_buf_1 input232 (.A(Tile_X0Y1_N2END[5]),
    .X(net232));
 sg13g2_buf_1 input233 (.A(Tile_X0Y1_N2END[6]),
    .X(net233));
 sg13g2_buf_1 input234 (.A(Tile_X0Y1_N2END[7]),
    .X(net234));
 sg13g2_buf_1 input235 (.A(Tile_X0Y1_N2MID[0]),
    .X(net235));
 sg13g2_buf_1 input236 (.A(Tile_X0Y1_N2MID[1]),
    .X(net236));
 sg13g2_buf_1 input237 (.A(Tile_X0Y1_N2MID[2]),
    .X(net237));
 sg13g2_buf_1 input238 (.A(Tile_X0Y1_N2MID[3]),
    .X(net238));
 sg13g2_buf_1 input239 (.A(Tile_X0Y1_N2MID[4]),
    .X(net239));
 sg13g2_buf_1 input240 (.A(Tile_X0Y1_N2MID[5]),
    .X(net240));
 sg13g2_buf_1 input241 (.A(Tile_X0Y1_N2MID[6]),
    .X(net241));
 sg13g2_buf_1 input242 (.A(Tile_X0Y1_N2MID[7]),
    .X(net242));
 sg13g2_buf_1 input243 (.A(Tile_X0Y1_N4END[0]),
    .X(net243));
 sg13g2_buf_1 input244 (.A(Tile_X0Y1_N4END[1]),
    .X(net244));
 sg13g2_buf_1 input245 (.A(Tile_X0Y1_N4END[2]),
    .X(net245));
 sg13g2_buf_1 input246 (.A(Tile_X0Y1_N4END[3]),
    .X(net246));
 sg13g2_buf_1 input247 (.A(Tile_X0Y1_N4END[4]),
    .X(net247));
 sg13g2_buf_1 input248 (.A(Tile_X0Y1_N4END[5]),
    .X(net248));
 sg13g2_buf_1 input249 (.A(Tile_X0Y1_N4END[6]),
    .X(net249));
 sg13g2_buf_1 input250 (.A(Tile_X0Y1_N4END[7]),
    .X(net250));
 sg13g2_buf_1 output251 (.A(net251),
    .X(ADDR_SRAM0));
 sg13g2_buf_1 output252 (.A(net252),
    .X(ADDR_SRAM1));
 sg13g2_buf_1 output253 (.A(net253),
    .X(ADDR_SRAM2));
 sg13g2_buf_1 output254 (.A(net254),
    .X(ADDR_SRAM3));
 sg13g2_buf_1 output255 (.A(net255),
    .X(ADDR_SRAM4));
 sg13g2_buf_1 output256 (.A(net256),
    .X(ADDR_SRAM5));
 sg13g2_buf_1 output257 (.A(net257),
    .X(ADDR_SRAM6));
 sg13g2_buf_1 output258 (.A(net258),
    .X(ADDR_SRAM7));
 sg13g2_buf_1 output259 (.A(net259),
    .X(ADDR_SRAM8));
 sg13g2_buf_1 output260 (.A(net260),
    .X(ADDR_SRAM9));
 sg13g2_buf_1 output261 (.A(net261),
    .X(BM_SRAM0));
 sg13g2_buf_1 output262 (.A(net262),
    .X(BM_SRAM1));
 sg13g2_buf_1 output263 (.A(net263),
    .X(BM_SRAM10));
 sg13g2_buf_1 output264 (.A(net264),
    .X(BM_SRAM11));
 sg13g2_buf_1 output265 (.A(net265),
    .X(BM_SRAM12));
 sg13g2_buf_1 output266 (.A(net266),
    .X(BM_SRAM13));
 sg13g2_buf_1 output267 (.A(net267),
    .X(BM_SRAM14));
 sg13g2_buf_1 output268 (.A(net268),
    .X(BM_SRAM15));
 sg13g2_buf_1 output269 (.A(net269),
    .X(BM_SRAM16));
 sg13g2_buf_1 output270 (.A(net270),
    .X(BM_SRAM17));
 sg13g2_buf_1 output271 (.A(net271),
    .X(BM_SRAM18));
 sg13g2_buf_1 output272 (.A(net272),
    .X(BM_SRAM19));
 sg13g2_buf_1 output273 (.A(net273),
    .X(BM_SRAM2));
 sg13g2_buf_1 output274 (.A(net274),
    .X(BM_SRAM20));
 sg13g2_buf_1 output275 (.A(net275),
    .X(BM_SRAM21));
 sg13g2_buf_1 output276 (.A(net276),
    .X(BM_SRAM22));
 sg13g2_buf_1 output277 (.A(net277),
    .X(BM_SRAM23));
 sg13g2_buf_1 output278 (.A(net278),
    .X(BM_SRAM24));
 sg13g2_buf_1 output279 (.A(net279),
    .X(BM_SRAM25));
 sg13g2_buf_1 output280 (.A(net280),
    .X(BM_SRAM26));
 sg13g2_buf_1 output281 (.A(net281),
    .X(BM_SRAM27));
 sg13g2_buf_1 output282 (.A(net282),
    .X(BM_SRAM28));
 sg13g2_buf_1 output283 (.A(net283),
    .X(BM_SRAM29));
 sg13g2_buf_1 output284 (.A(net284),
    .X(BM_SRAM3));
 sg13g2_buf_1 output285 (.A(net285),
    .X(BM_SRAM30));
 sg13g2_buf_1 output286 (.A(net286),
    .X(BM_SRAM31));
 sg13g2_buf_1 output287 (.A(net287),
    .X(BM_SRAM4));
 sg13g2_buf_1 output288 (.A(net288),
    .X(BM_SRAM5));
 sg13g2_buf_1 output289 (.A(net289),
    .X(BM_SRAM6));
 sg13g2_buf_1 output290 (.A(net290),
    .X(BM_SRAM7));
 sg13g2_buf_1 output291 (.A(net291),
    .X(BM_SRAM8));
 sg13g2_buf_1 output292 (.A(net292),
    .X(BM_SRAM9));
 sg13g2_buf_1 output293 (.A(net293),
    .X(CLK_SRAM));
 sg13g2_buf_1 output294 (.A(net294),
    .X(DIN_SRAM0));
 sg13g2_buf_1 output295 (.A(net295),
    .X(DIN_SRAM1));
 sg13g2_buf_1 output296 (.A(net296),
    .X(DIN_SRAM10));
 sg13g2_buf_1 output297 (.A(net297),
    .X(DIN_SRAM11));
 sg13g2_buf_1 output298 (.A(net298),
    .X(DIN_SRAM12));
 sg13g2_buf_1 output299 (.A(net299),
    .X(DIN_SRAM13));
 sg13g2_buf_1 output300 (.A(net300),
    .X(DIN_SRAM14));
 sg13g2_buf_1 output301 (.A(net301),
    .X(DIN_SRAM15));
 sg13g2_buf_1 output302 (.A(net302),
    .X(DIN_SRAM16));
 sg13g2_buf_1 output303 (.A(net303),
    .X(DIN_SRAM17));
 sg13g2_buf_1 output304 (.A(net304),
    .X(DIN_SRAM18));
 sg13g2_buf_1 output305 (.A(net305),
    .X(DIN_SRAM19));
 sg13g2_buf_1 output306 (.A(net306),
    .X(DIN_SRAM2));
 sg13g2_buf_1 output307 (.A(net307),
    .X(DIN_SRAM20));
 sg13g2_buf_1 output308 (.A(net308),
    .X(DIN_SRAM21));
 sg13g2_buf_1 output309 (.A(net309),
    .X(DIN_SRAM22));
 sg13g2_buf_1 output310 (.A(net310),
    .X(DIN_SRAM23));
 sg13g2_buf_1 output311 (.A(net311),
    .X(DIN_SRAM24));
 sg13g2_buf_1 output312 (.A(net312),
    .X(DIN_SRAM25));
 sg13g2_buf_1 output313 (.A(net313),
    .X(DIN_SRAM26));
 sg13g2_buf_1 output314 (.A(net314),
    .X(DIN_SRAM27));
 sg13g2_buf_1 output315 (.A(net315),
    .X(DIN_SRAM28));
 sg13g2_buf_1 output316 (.A(net316),
    .X(DIN_SRAM29));
 sg13g2_buf_1 output317 (.A(net317),
    .X(DIN_SRAM3));
 sg13g2_buf_1 output318 (.A(net318),
    .X(DIN_SRAM30));
 sg13g2_buf_1 output319 (.A(net319),
    .X(DIN_SRAM31));
 sg13g2_buf_1 output320 (.A(net320),
    .X(DIN_SRAM4));
 sg13g2_buf_1 output321 (.A(net321),
    .X(DIN_SRAM5));
 sg13g2_buf_1 output322 (.A(net322),
    .X(DIN_SRAM6));
 sg13g2_buf_1 output323 (.A(net323),
    .X(DIN_SRAM7));
 sg13g2_buf_1 output324 (.A(net324),
    .X(DIN_SRAM8));
 sg13g2_buf_1 output325 (.A(net325),
    .X(DIN_SRAM9));
 sg13g2_buf_1 output326 (.A(net326),
    .X(MEN_SRAM));
 sg13g2_buf_1 output327 (.A(net327),
    .X(REN_SRAM));
 sg13g2_buf_1 output328 (.A(net328),
    .X(Tile_X0Y0_FrameData_O[0]));
 sg13g2_buf_1 output329 (.A(net329),
    .X(Tile_X0Y0_FrameData_O[10]));
 sg13g2_buf_1 output330 (.A(net330),
    .X(Tile_X0Y0_FrameData_O[11]));
 sg13g2_buf_1 output331 (.A(net331),
    .X(Tile_X0Y0_FrameData_O[12]));
 sg13g2_buf_1 output332 (.A(net332),
    .X(Tile_X0Y0_FrameData_O[13]));
 sg13g2_buf_1 output333 (.A(net333),
    .X(Tile_X0Y0_FrameData_O[14]));
 sg13g2_buf_1 output334 (.A(net334),
    .X(Tile_X0Y0_FrameData_O[15]));
 sg13g2_buf_1 output335 (.A(net335),
    .X(Tile_X0Y0_FrameData_O[16]));
 sg13g2_buf_1 output336 (.A(net336),
    .X(Tile_X0Y0_FrameData_O[17]));
 sg13g2_buf_1 output337 (.A(net337),
    .X(Tile_X0Y0_FrameData_O[18]));
 sg13g2_buf_1 output338 (.A(net338),
    .X(Tile_X0Y0_FrameData_O[19]));
 sg13g2_buf_1 output339 (.A(net339),
    .X(Tile_X0Y0_FrameData_O[1]));
 sg13g2_buf_1 output340 (.A(net340),
    .X(Tile_X0Y0_FrameData_O[20]));
 sg13g2_buf_1 output341 (.A(net341),
    .X(Tile_X0Y0_FrameData_O[21]));
 sg13g2_buf_1 output342 (.A(net342),
    .X(Tile_X0Y0_FrameData_O[22]));
 sg13g2_buf_1 output343 (.A(net343),
    .X(Tile_X0Y0_FrameData_O[23]));
 sg13g2_buf_1 output344 (.A(net344),
    .X(Tile_X0Y0_FrameData_O[24]));
 sg13g2_buf_1 output345 (.A(net345),
    .X(Tile_X0Y0_FrameData_O[25]));
 sg13g2_buf_1 output346 (.A(net346),
    .X(Tile_X0Y0_FrameData_O[26]));
 sg13g2_buf_1 output347 (.A(net347),
    .X(Tile_X0Y0_FrameData_O[27]));
 sg13g2_buf_1 output348 (.A(net348),
    .X(Tile_X0Y0_FrameData_O[28]));
 sg13g2_buf_1 output349 (.A(net349),
    .X(Tile_X0Y0_FrameData_O[29]));
 sg13g2_buf_1 output350 (.A(net350),
    .X(Tile_X0Y0_FrameData_O[2]));
 sg13g2_buf_1 output351 (.A(net351),
    .X(Tile_X0Y0_FrameData_O[30]));
 sg13g2_buf_1 output352 (.A(net352),
    .X(Tile_X0Y0_FrameData_O[31]));
 sg13g2_buf_1 output353 (.A(net353),
    .X(Tile_X0Y0_FrameData_O[3]));
 sg13g2_buf_1 output354 (.A(net354),
    .X(Tile_X0Y0_FrameData_O[4]));
 sg13g2_buf_1 output355 (.A(net355),
    .X(Tile_X0Y0_FrameData_O[5]));
 sg13g2_buf_1 output356 (.A(net356),
    .X(Tile_X0Y0_FrameData_O[6]));
 sg13g2_buf_1 output357 (.A(net357),
    .X(Tile_X0Y0_FrameData_O[7]));
 sg13g2_buf_1 output358 (.A(net358),
    .X(Tile_X0Y0_FrameData_O[8]));
 sg13g2_buf_1 output359 (.A(net359),
    .X(Tile_X0Y0_FrameData_O[9]));
 sg13g2_buf_1 output360 (.A(net360),
    .X(Tile_X0Y0_FrameStrobe_O[0]));
 sg13g2_buf_1 output361 (.A(net361),
    .X(Tile_X0Y0_FrameStrobe_O[10]));
 sg13g2_buf_1 output362 (.A(net362),
    .X(Tile_X0Y0_FrameStrobe_O[11]));
 sg13g2_buf_1 output363 (.A(net363),
    .X(Tile_X0Y0_FrameStrobe_O[12]));
 sg13g2_buf_1 output364 (.A(net364),
    .X(Tile_X0Y0_FrameStrobe_O[13]));
 sg13g2_buf_1 output365 (.A(net365),
    .X(Tile_X0Y0_FrameStrobe_O[14]));
 sg13g2_buf_1 output366 (.A(net366),
    .X(Tile_X0Y0_FrameStrobe_O[15]));
 sg13g2_buf_1 output367 (.A(net367),
    .X(Tile_X0Y0_FrameStrobe_O[16]));
 sg13g2_buf_1 output368 (.A(net368),
    .X(Tile_X0Y0_FrameStrobe_O[17]));
 sg13g2_buf_1 output369 (.A(net369),
    .X(Tile_X0Y0_FrameStrobe_O[18]));
 sg13g2_buf_1 output370 (.A(net370),
    .X(Tile_X0Y0_FrameStrobe_O[19]));
 sg13g2_buf_1 output371 (.A(net371),
    .X(Tile_X0Y0_FrameStrobe_O[1]));
 sg13g2_buf_1 output372 (.A(net372),
    .X(Tile_X0Y0_FrameStrobe_O[2]));
 sg13g2_buf_1 output373 (.A(net373),
    .X(Tile_X0Y0_FrameStrobe_O[3]));
 sg13g2_buf_1 output374 (.A(net374),
    .X(Tile_X0Y0_FrameStrobe_O[4]));
 sg13g2_buf_1 output375 (.A(net375),
    .X(Tile_X0Y0_FrameStrobe_O[5]));
 sg13g2_buf_1 output376 (.A(net376),
    .X(Tile_X0Y0_FrameStrobe_O[6]));
 sg13g2_buf_1 output377 (.A(net377),
    .X(Tile_X0Y0_FrameStrobe_O[7]));
 sg13g2_buf_1 output378 (.A(net378),
    .X(Tile_X0Y0_FrameStrobe_O[8]));
 sg13g2_buf_1 output379 (.A(net379),
    .X(Tile_X0Y0_FrameStrobe_O[9]));
 sg13g2_buf_1 output380 (.A(net380),
    .X(Tile_X0Y0_N1BEG[0]));
 sg13g2_buf_1 output381 (.A(net381),
    .X(Tile_X0Y0_N1BEG[1]));
 sg13g2_buf_1 output382 (.A(net382),
    .X(Tile_X0Y0_N1BEG[2]));
 sg13g2_buf_1 output383 (.A(net383),
    .X(Tile_X0Y0_N1BEG[3]));
 sg13g2_buf_1 output384 (.A(net384),
    .X(Tile_X0Y0_N2BEG[0]));
 sg13g2_buf_1 output385 (.A(net385),
    .X(Tile_X0Y0_N2BEG[1]));
 sg13g2_buf_1 output386 (.A(net386),
    .X(Tile_X0Y0_N2BEG[2]));
 sg13g2_buf_1 output387 (.A(net387),
    .X(Tile_X0Y0_N2BEG[3]));
 sg13g2_buf_1 output388 (.A(net388),
    .X(Tile_X0Y0_N2BEG[4]));
 sg13g2_buf_1 output389 (.A(net389),
    .X(Tile_X0Y0_N2BEG[5]));
 sg13g2_buf_1 output390 (.A(net390),
    .X(Tile_X0Y0_N2BEG[6]));
 sg13g2_buf_1 output391 (.A(net391),
    .X(Tile_X0Y0_N2BEG[7]));
 sg13g2_buf_1 output392 (.A(net392),
    .X(Tile_X0Y0_N2BEGb[0]));
 sg13g2_buf_1 output393 (.A(net393),
    .X(Tile_X0Y0_N2BEGb[1]));
 sg13g2_buf_1 output394 (.A(net394),
    .X(Tile_X0Y0_N2BEGb[2]));
 sg13g2_buf_1 output395 (.A(net395),
    .X(Tile_X0Y0_N2BEGb[3]));
 sg13g2_buf_1 output396 (.A(net396),
    .X(Tile_X0Y0_N2BEGb[4]));
 sg13g2_buf_1 output397 (.A(net397),
    .X(Tile_X0Y0_N2BEGb[5]));
 sg13g2_buf_1 output398 (.A(net398),
    .X(Tile_X0Y0_N2BEGb[6]));
 sg13g2_buf_1 output399 (.A(net399),
    .X(Tile_X0Y0_N2BEGb[7]));
 sg13g2_buf_1 output400 (.A(net400),
    .X(Tile_X0Y0_N4BEG[0]));
 sg13g2_buf_1 output401 (.A(net401),
    .X(Tile_X0Y0_N4BEG[10]));
 sg13g2_buf_1 output402 (.A(net402),
    .X(Tile_X0Y0_N4BEG[11]));
 sg13g2_buf_1 output403 (.A(net403),
    .X(Tile_X0Y0_N4BEG[12]));
 sg13g2_buf_1 output404 (.A(net404),
    .X(Tile_X0Y0_N4BEG[13]));
 sg13g2_buf_1 output405 (.A(net405),
    .X(Tile_X0Y0_N4BEG[14]));
 sg13g2_buf_1 output406 (.A(net406),
    .X(Tile_X0Y0_N4BEG[15]));
 sg13g2_buf_1 output407 (.A(net407),
    .X(Tile_X0Y0_N4BEG[1]));
 sg13g2_buf_1 output408 (.A(net408),
    .X(Tile_X0Y0_N4BEG[2]));
 sg13g2_buf_1 output409 (.A(net409),
    .X(Tile_X0Y0_N4BEG[3]));
 sg13g2_buf_1 output410 (.A(net410),
    .X(Tile_X0Y0_N4BEG[4]));
 sg13g2_buf_1 output411 (.A(net411),
    .X(Tile_X0Y0_N4BEG[5]));
 sg13g2_buf_1 output412 (.A(net412),
    .X(Tile_X0Y0_N4BEG[6]));
 sg13g2_buf_1 output413 (.A(net413),
    .X(Tile_X0Y0_N4BEG[7]));
 sg13g2_buf_1 output414 (.A(net414),
    .X(Tile_X0Y0_N4BEG[8]));
 sg13g2_buf_1 output415 (.A(net415),
    .X(Tile_X0Y0_N4BEG[9]));
 sg13g2_buf_1 output416 (.A(net416),
    .X(Tile_X0Y0_UserCLKo));
 sg13g2_buf_1 output417 (.A(net417),
    .X(Tile_X0Y0_W1BEG[0]));
 sg13g2_buf_1 output418 (.A(net418),
    .X(Tile_X0Y0_W1BEG[1]));
 sg13g2_buf_1 output419 (.A(net419),
    .X(Tile_X0Y0_W1BEG[2]));
 sg13g2_buf_1 output420 (.A(net420),
    .X(Tile_X0Y0_W1BEG[3]));
 sg13g2_buf_1 output421 (.A(net421),
    .X(Tile_X0Y0_W2BEG[0]));
 sg13g2_buf_1 output422 (.A(net422),
    .X(Tile_X0Y0_W2BEG[1]));
 sg13g2_buf_1 output423 (.A(net423),
    .X(Tile_X0Y0_W2BEG[2]));
 sg13g2_buf_1 output424 (.A(net424),
    .X(Tile_X0Y0_W2BEG[3]));
 sg13g2_buf_1 output425 (.A(net425),
    .X(Tile_X0Y0_W2BEG[4]));
 sg13g2_buf_1 output426 (.A(net426),
    .X(Tile_X0Y0_W2BEG[5]));
 sg13g2_buf_1 output427 (.A(net427),
    .X(Tile_X0Y0_W2BEG[6]));
 sg13g2_buf_1 output428 (.A(net428),
    .X(Tile_X0Y0_W2BEG[7]));
 sg13g2_buf_1 output429 (.A(net429),
    .X(Tile_X0Y0_W2BEGb[0]));
 sg13g2_buf_1 output430 (.A(net430),
    .X(Tile_X0Y0_W2BEGb[1]));
 sg13g2_buf_1 output431 (.A(net431),
    .X(Tile_X0Y0_W2BEGb[2]));
 sg13g2_buf_1 output432 (.A(net432),
    .X(Tile_X0Y0_W2BEGb[3]));
 sg13g2_buf_1 output433 (.A(net433),
    .X(Tile_X0Y0_W2BEGb[4]));
 sg13g2_buf_1 output434 (.A(net434),
    .X(Tile_X0Y0_W2BEGb[5]));
 sg13g2_buf_1 output435 (.A(net435),
    .X(Tile_X0Y0_W2BEGb[6]));
 sg13g2_buf_1 output436 (.A(net436),
    .X(Tile_X0Y0_W2BEGb[7]));
 sg13g2_buf_1 output437 (.A(net437),
    .X(Tile_X0Y0_W6BEG[0]));
 sg13g2_buf_1 output438 (.A(net438),
    .X(Tile_X0Y0_W6BEG[10]));
 sg13g2_buf_1 output439 (.A(net439),
    .X(Tile_X0Y0_W6BEG[11]));
 sg13g2_buf_1 output440 (.A(net440),
    .X(Tile_X0Y0_W6BEG[1]));
 sg13g2_buf_1 output441 (.A(net441),
    .X(Tile_X0Y0_W6BEG[2]));
 sg13g2_buf_1 output442 (.A(net442),
    .X(Tile_X0Y0_W6BEG[3]));
 sg13g2_buf_1 output443 (.A(net443),
    .X(Tile_X0Y0_W6BEG[4]));
 sg13g2_buf_1 output444 (.A(net444),
    .X(Tile_X0Y0_W6BEG[5]));
 sg13g2_buf_1 output445 (.A(net445),
    .X(Tile_X0Y0_W6BEG[6]));
 sg13g2_buf_1 output446 (.A(net446),
    .X(Tile_X0Y0_W6BEG[7]));
 sg13g2_buf_1 output447 (.A(net447),
    .X(Tile_X0Y0_W6BEG[8]));
 sg13g2_buf_1 output448 (.A(net448),
    .X(Tile_X0Y0_W6BEG[9]));
 sg13g2_buf_1 output449 (.A(net449),
    .X(Tile_X0Y0_WW4BEG[0]));
 sg13g2_buf_1 output450 (.A(net450),
    .X(Tile_X0Y0_WW4BEG[10]));
 sg13g2_buf_1 output451 (.A(net451),
    .X(Tile_X0Y0_WW4BEG[11]));
 sg13g2_buf_1 output452 (.A(net452),
    .X(Tile_X0Y0_WW4BEG[12]));
 sg13g2_buf_1 output453 (.A(net453),
    .X(Tile_X0Y0_WW4BEG[13]));
 sg13g2_buf_1 output454 (.A(net454),
    .X(Tile_X0Y0_WW4BEG[14]));
 sg13g2_buf_1 output455 (.A(net455),
    .X(Tile_X0Y0_WW4BEG[15]));
 sg13g2_buf_1 output456 (.A(net456),
    .X(Tile_X0Y0_WW4BEG[1]));
 sg13g2_buf_1 output457 (.A(net457),
    .X(Tile_X0Y0_WW4BEG[2]));
 sg13g2_buf_1 output458 (.A(net458),
    .X(Tile_X0Y0_WW4BEG[3]));
 sg13g2_buf_1 output459 (.A(net459),
    .X(Tile_X0Y0_WW4BEG[4]));
 sg13g2_buf_1 output460 (.A(net460),
    .X(Tile_X0Y0_WW4BEG[5]));
 sg13g2_buf_1 output461 (.A(net461),
    .X(Tile_X0Y0_WW4BEG[6]));
 sg13g2_buf_1 output462 (.A(net462),
    .X(Tile_X0Y0_WW4BEG[7]));
 sg13g2_buf_1 output463 (.A(net463),
    .X(Tile_X0Y0_WW4BEG[8]));
 sg13g2_buf_1 output464 (.A(net464),
    .X(Tile_X0Y0_WW4BEG[9]));
 sg13g2_buf_1 output465 (.A(net465),
    .X(Tile_X0Y1_FrameData_O[0]));
 sg13g2_buf_1 output466 (.A(net466),
    .X(Tile_X0Y1_FrameData_O[10]));
 sg13g2_buf_1 output467 (.A(net467),
    .X(Tile_X0Y1_FrameData_O[11]));
 sg13g2_buf_1 output468 (.A(net468),
    .X(Tile_X0Y1_FrameData_O[12]));
 sg13g2_buf_1 output469 (.A(net469),
    .X(Tile_X0Y1_FrameData_O[13]));
 sg13g2_buf_1 output470 (.A(net470),
    .X(Tile_X0Y1_FrameData_O[14]));
 sg13g2_buf_1 output471 (.A(net471),
    .X(Tile_X0Y1_FrameData_O[15]));
 sg13g2_buf_1 output472 (.A(net472),
    .X(Tile_X0Y1_FrameData_O[16]));
 sg13g2_buf_1 output473 (.A(net473),
    .X(Tile_X0Y1_FrameData_O[17]));
 sg13g2_buf_1 output474 (.A(net474),
    .X(Tile_X0Y1_FrameData_O[18]));
 sg13g2_buf_1 output475 (.A(net475),
    .X(Tile_X0Y1_FrameData_O[19]));
 sg13g2_buf_1 output476 (.A(net476),
    .X(Tile_X0Y1_FrameData_O[1]));
 sg13g2_buf_1 output477 (.A(net477),
    .X(Tile_X0Y1_FrameData_O[20]));
 sg13g2_buf_1 output478 (.A(net478),
    .X(Tile_X0Y1_FrameData_O[21]));
 sg13g2_buf_1 output479 (.A(net479),
    .X(Tile_X0Y1_FrameData_O[22]));
 sg13g2_buf_1 output480 (.A(net480),
    .X(Tile_X0Y1_FrameData_O[23]));
 sg13g2_buf_1 output481 (.A(net481),
    .X(Tile_X0Y1_FrameData_O[24]));
 sg13g2_buf_1 output482 (.A(net482),
    .X(Tile_X0Y1_FrameData_O[25]));
 sg13g2_buf_1 output483 (.A(net483),
    .X(Tile_X0Y1_FrameData_O[26]));
 sg13g2_buf_1 output484 (.A(net484),
    .X(Tile_X0Y1_FrameData_O[27]));
 sg13g2_buf_1 output485 (.A(net485),
    .X(Tile_X0Y1_FrameData_O[28]));
 sg13g2_buf_1 output486 (.A(net486),
    .X(Tile_X0Y1_FrameData_O[29]));
 sg13g2_buf_1 output487 (.A(net487),
    .X(Tile_X0Y1_FrameData_O[2]));
 sg13g2_buf_1 output488 (.A(net488),
    .X(Tile_X0Y1_FrameData_O[30]));
 sg13g2_buf_1 output489 (.A(net489),
    .X(Tile_X0Y1_FrameData_O[31]));
 sg13g2_buf_1 output490 (.A(net490),
    .X(Tile_X0Y1_FrameData_O[3]));
 sg13g2_buf_1 output491 (.A(net491),
    .X(Tile_X0Y1_FrameData_O[4]));
 sg13g2_buf_1 output492 (.A(net492),
    .X(Tile_X0Y1_FrameData_O[5]));
 sg13g2_buf_1 output493 (.A(net493),
    .X(Tile_X0Y1_FrameData_O[6]));
 sg13g2_buf_1 output494 (.A(net494),
    .X(Tile_X0Y1_FrameData_O[7]));
 sg13g2_buf_1 output495 (.A(net495),
    .X(Tile_X0Y1_FrameData_O[8]));
 sg13g2_buf_1 output496 (.A(net496),
    .X(Tile_X0Y1_FrameData_O[9]));
 sg13g2_buf_1 output497 (.A(net497),
    .X(Tile_X0Y1_S1BEG[0]));
 sg13g2_buf_1 output498 (.A(net498),
    .X(Tile_X0Y1_S1BEG[1]));
 sg13g2_buf_1 output499 (.A(net499),
    .X(Tile_X0Y1_S1BEG[2]));
 sg13g2_buf_1 output500 (.A(net500),
    .X(Tile_X0Y1_S1BEG[3]));
 sg13g2_buf_1 output501 (.A(net501),
    .X(Tile_X0Y1_S2BEG[0]));
 sg13g2_buf_1 output502 (.A(net502),
    .X(Tile_X0Y1_S2BEG[1]));
 sg13g2_buf_1 output503 (.A(net503),
    .X(Tile_X0Y1_S2BEG[2]));
 sg13g2_buf_1 output504 (.A(net504),
    .X(Tile_X0Y1_S2BEG[3]));
 sg13g2_buf_1 output505 (.A(net505),
    .X(Tile_X0Y1_S2BEG[4]));
 sg13g2_buf_1 output506 (.A(net506),
    .X(Tile_X0Y1_S2BEG[5]));
 sg13g2_buf_1 output507 (.A(net507),
    .X(Tile_X0Y1_S2BEG[6]));
 sg13g2_buf_1 output508 (.A(net508),
    .X(Tile_X0Y1_S2BEG[7]));
 sg13g2_buf_1 output509 (.A(net509),
    .X(Tile_X0Y1_S2BEGb[0]));
 sg13g2_buf_1 output510 (.A(net510),
    .X(Tile_X0Y1_S2BEGb[1]));
 sg13g2_buf_1 output511 (.A(net511),
    .X(Tile_X0Y1_S2BEGb[2]));
 sg13g2_buf_1 output512 (.A(net512),
    .X(Tile_X0Y1_S2BEGb[3]));
 sg13g2_buf_1 output513 (.A(net513),
    .X(Tile_X0Y1_S2BEGb[4]));
 sg13g2_buf_1 output514 (.A(net514),
    .X(Tile_X0Y1_S2BEGb[5]));
 sg13g2_buf_1 output515 (.A(net515),
    .X(Tile_X0Y1_S2BEGb[6]));
 sg13g2_buf_1 output516 (.A(net516),
    .X(Tile_X0Y1_S2BEGb[7]));
 sg13g2_buf_1 output517 (.A(net517),
    .X(Tile_X0Y1_S4BEG[0]));
 sg13g2_buf_1 output518 (.A(net518),
    .X(Tile_X0Y1_S4BEG[10]));
 sg13g2_buf_1 output519 (.A(net519),
    .X(Tile_X0Y1_S4BEG[11]));
 sg13g2_buf_1 output520 (.A(net520),
    .X(Tile_X0Y1_S4BEG[12]));
 sg13g2_buf_1 output521 (.A(net521),
    .X(Tile_X0Y1_S4BEG[13]));
 sg13g2_buf_1 output522 (.A(net522),
    .X(Tile_X0Y1_S4BEG[14]));
 sg13g2_buf_1 output523 (.A(net523),
    .X(Tile_X0Y1_S4BEG[15]));
 sg13g2_buf_1 output524 (.A(net524),
    .X(Tile_X0Y1_S4BEG[1]));
 sg13g2_buf_1 output525 (.A(net525),
    .X(Tile_X0Y1_S4BEG[2]));
 sg13g2_buf_1 output526 (.A(net526),
    .X(Tile_X0Y1_S4BEG[3]));
 sg13g2_buf_1 output527 (.A(net527),
    .X(Tile_X0Y1_S4BEG[4]));
 sg13g2_buf_1 output528 (.A(net528),
    .X(Tile_X0Y1_S4BEG[5]));
 sg13g2_buf_1 output529 (.A(net529),
    .X(Tile_X0Y1_S4BEG[6]));
 sg13g2_buf_1 output530 (.A(net530),
    .X(Tile_X0Y1_S4BEG[7]));
 sg13g2_buf_1 output531 (.A(net531),
    .X(Tile_X0Y1_S4BEG[8]));
 sg13g2_buf_1 output532 (.A(net532),
    .X(Tile_X0Y1_S4BEG[9]));
 sg13g2_buf_1 output533 (.A(net533),
    .X(Tile_X0Y1_W1BEG[0]));
 sg13g2_buf_1 output534 (.A(net534),
    .X(Tile_X0Y1_W1BEG[1]));
 sg13g2_buf_1 output535 (.A(net535),
    .X(Tile_X0Y1_W1BEG[2]));
 sg13g2_buf_1 output536 (.A(net536),
    .X(Tile_X0Y1_W1BEG[3]));
 sg13g2_buf_1 output537 (.A(net537),
    .X(Tile_X0Y1_W2BEG[0]));
 sg13g2_buf_1 output538 (.A(net538),
    .X(Tile_X0Y1_W2BEG[1]));
 sg13g2_buf_1 output539 (.A(net539),
    .X(Tile_X0Y1_W2BEG[2]));
 sg13g2_buf_1 output540 (.A(net540),
    .X(Tile_X0Y1_W2BEG[3]));
 sg13g2_buf_1 output541 (.A(net541),
    .X(Tile_X0Y1_W2BEG[4]));
 sg13g2_buf_1 output542 (.A(net542),
    .X(Tile_X0Y1_W2BEG[5]));
 sg13g2_buf_1 output543 (.A(net543),
    .X(Tile_X0Y1_W2BEG[6]));
 sg13g2_buf_1 output544 (.A(net544),
    .X(Tile_X0Y1_W2BEG[7]));
 sg13g2_buf_1 output545 (.A(net545),
    .X(Tile_X0Y1_W2BEGb[0]));
 sg13g2_buf_1 output546 (.A(net546),
    .X(Tile_X0Y1_W2BEGb[1]));
 sg13g2_buf_1 output547 (.A(net547),
    .X(Tile_X0Y1_W2BEGb[2]));
 sg13g2_buf_1 output548 (.A(net548),
    .X(Tile_X0Y1_W2BEGb[3]));
 sg13g2_buf_1 output549 (.A(net549),
    .X(Tile_X0Y1_W2BEGb[4]));
 sg13g2_buf_1 output550 (.A(net550),
    .X(Tile_X0Y1_W2BEGb[5]));
 sg13g2_buf_1 output551 (.A(net551),
    .X(Tile_X0Y1_W2BEGb[6]));
 sg13g2_buf_1 output552 (.A(net552),
    .X(Tile_X0Y1_W2BEGb[7]));
 sg13g2_buf_1 output553 (.A(net553),
    .X(Tile_X0Y1_W6BEG[0]));
 sg13g2_buf_1 output554 (.A(net554),
    .X(Tile_X0Y1_W6BEG[10]));
 sg13g2_buf_1 output555 (.A(net555),
    .X(Tile_X0Y1_W6BEG[11]));
 sg13g2_buf_1 output556 (.A(net556),
    .X(Tile_X0Y1_W6BEG[1]));
 sg13g2_buf_1 output557 (.A(net557),
    .X(Tile_X0Y1_W6BEG[2]));
 sg13g2_buf_1 output558 (.A(net558),
    .X(Tile_X0Y1_W6BEG[3]));
 sg13g2_buf_1 output559 (.A(net559),
    .X(Tile_X0Y1_W6BEG[4]));
 sg13g2_buf_1 output560 (.A(net560),
    .X(Tile_X0Y1_W6BEG[5]));
 sg13g2_buf_1 output561 (.A(net561),
    .X(Tile_X0Y1_W6BEG[6]));
 sg13g2_buf_1 output562 (.A(net562),
    .X(Tile_X0Y1_W6BEG[7]));
 sg13g2_buf_1 output563 (.A(net563),
    .X(Tile_X0Y1_W6BEG[8]));
 sg13g2_buf_1 output564 (.A(net564),
    .X(Tile_X0Y1_W6BEG[9]));
 sg13g2_buf_1 output565 (.A(net565),
    .X(Tile_X0Y1_WW4BEG[0]));
 sg13g2_buf_1 output566 (.A(net566),
    .X(Tile_X0Y1_WW4BEG[10]));
 sg13g2_buf_1 output567 (.A(net567),
    .X(Tile_X0Y1_WW4BEG[11]));
 sg13g2_buf_1 output568 (.A(net568),
    .X(Tile_X0Y1_WW4BEG[12]));
 sg13g2_buf_1 output569 (.A(net569),
    .X(Tile_X0Y1_WW4BEG[13]));
 sg13g2_buf_1 output570 (.A(net570),
    .X(Tile_X0Y1_WW4BEG[14]));
 sg13g2_buf_1 output571 (.A(net571),
    .X(Tile_X0Y1_WW4BEG[15]));
 sg13g2_buf_1 output572 (.A(net572),
    .X(Tile_X0Y1_WW4BEG[1]));
 sg13g2_buf_1 output573 (.A(net573),
    .X(Tile_X0Y1_WW4BEG[2]));
 sg13g2_buf_1 output574 (.A(net574),
    .X(Tile_X0Y1_WW4BEG[3]));
 sg13g2_buf_1 output575 (.A(net575),
    .X(Tile_X0Y1_WW4BEG[4]));
 sg13g2_buf_1 output576 (.A(net576),
    .X(Tile_X0Y1_WW4BEG[5]));
 sg13g2_buf_1 output577 (.A(net577),
    .X(Tile_X0Y1_WW4BEG[6]));
 sg13g2_buf_1 output578 (.A(net578),
    .X(Tile_X0Y1_WW4BEG[7]));
 sg13g2_buf_1 output579 (.A(net579),
    .X(Tile_X0Y1_WW4BEG[8]));
 sg13g2_buf_1 output580 (.A(net580),
    .X(Tile_X0Y1_WW4BEG[9]));
 sg13g2_buf_1 output581 (.A(net581),
    .X(WEN_SRAM));
 sg13g2_tielo IHP_SRAM_582 (.L_LO(net582));
 sg13g2_decap_4 FILLER_0_69 ();
 sg13g2_decap_8 FILLER_0_161 ();
 sg13g2_fill_1 FILLER_0_168 ();
 sg13g2_decap_8 FILLER_0_173 ();
 sg13g2_decap_8 FILLER_0_180 ();
 sg13g2_decap_8 FILLER_0_187 ();
 sg13g2_decap_8 FILLER_0_194 ();
 sg13g2_fill_1 FILLER_1_4 ();
 sg13g2_fill_1 FILLER_1_13 ();
 sg13g2_fill_2 FILLER_1_18 ();
 sg13g2_fill_1 FILLER_1_20 ();
 sg13g2_decap_8 FILLER_1_53 ();
 sg13g2_decap_8 FILLER_1_60 ();
 sg13g2_decap_4 FILLER_1_67 ();
 sg13g2_fill_2 FILLER_1_71 ();
 sg13g2_decap_4 FILLER_1_77 ();
 sg13g2_decap_8 FILLER_1_105 ();
 sg13g2_decap_8 FILLER_1_112 ();
 sg13g2_decap_8 FILLER_1_151 ();
 sg13g2_decap_8 FILLER_1_158 ();
 sg13g2_decap_8 FILLER_1_165 ();
 sg13g2_decap_8 FILLER_1_172 ();
 sg13g2_decap_8 FILLER_1_179 ();
 sg13g2_decap_8 FILLER_1_186 ();
 sg13g2_decap_8 FILLER_1_193 ();
 sg13g2_fill_1 FILLER_1_200 ();
 sg13g2_decap_8 FILLER_2_28 ();
 sg13g2_decap_8 FILLER_2_35 ();
 sg13g2_decap_8 FILLER_2_42 ();
 sg13g2_decap_8 FILLER_2_49 ();
 sg13g2_decap_8 FILLER_2_56 ();
 sg13g2_decap_8 FILLER_2_63 ();
 sg13g2_decap_8 FILLER_2_70 ();
 sg13g2_decap_8 FILLER_2_77 ();
 sg13g2_decap_8 FILLER_2_84 ();
 sg13g2_decap_8 FILLER_2_91 ();
 sg13g2_decap_8 FILLER_2_98 ();
 sg13g2_decap_8 FILLER_2_105 ();
 sg13g2_decap_8 FILLER_2_112 ();
 sg13g2_decap_8 FILLER_2_119 ();
 sg13g2_decap_8 FILLER_2_126 ();
 sg13g2_decap_8 FILLER_2_133 ();
 sg13g2_decap_8 FILLER_2_140 ();
 sg13g2_decap_8 FILLER_2_147 ();
 sg13g2_decap_8 FILLER_2_154 ();
 sg13g2_decap_8 FILLER_2_161 ();
 sg13g2_decap_8 FILLER_2_168 ();
 sg13g2_decap_8 FILLER_2_175 ();
 sg13g2_decap_8 FILLER_2_182 ();
 sg13g2_decap_8 FILLER_2_189 ();
 sg13g2_fill_1 FILLER_2_196 ();
 sg13g2_decap_8 FILLER_3_20 ();
 sg13g2_decap_8 FILLER_3_27 ();
 sg13g2_decap_8 FILLER_3_34 ();
 sg13g2_decap_8 FILLER_3_41 ();
 sg13g2_decap_8 FILLER_3_48 ();
 sg13g2_decap_8 FILLER_3_55 ();
 sg13g2_decap_8 FILLER_3_62 ();
 sg13g2_decap_8 FILLER_3_69 ();
 sg13g2_decap_8 FILLER_3_76 ();
 sg13g2_decap_8 FILLER_3_83 ();
 sg13g2_decap_8 FILLER_3_90 ();
 sg13g2_decap_4 FILLER_3_97 ();
 sg13g2_decap_8 FILLER_3_118 ();
 sg13g2_decap_8 FILLER_3_125 ();
 sg13g2_decap_8 FILLER_3_132 ();
 sg13g2_decap_8 FILLER_3_139 ();
 sg13g2_decap_8 FILLER_3_146 ();
 sg13g2_decap_8 FILLER_3_153 ();
 sg13g2_decap_8 FILLER_3_160 ();
 sg13g2_decap_8 FILLER_3_167 ();
 sg13g2_decap_8 FILLER_3_174 ();
 sg13g2_decap_8 FILLER_3_181 ();
 sg13g2_decap_4 FILLER_3_188 ();
 sg13g2_fill_1 FILLER_3_192 ();
 sg13g2_decap_8 FILLER_4_20 ();
 sg13g2_decap_8 FILLER_4_27 ();
 sg13g2_decap_8 FILLER_4_34 ();
 sg13g2_decap_8 FILLER_4_41 ();
 sg13g2_decap_8 FILLER_4_48 ();
 sg13g2_fill_1 FILLER_4_55 ();
 sg13g2_decap_8 FILLER_4_73 ();
 sg13g2_fill_2 FILLER_4_80 ();
 sg13g2_decap_4 FILLER_4_128 ();
 sg13g2_decap_8 FILLER_4_157 ();
 sg13g2_decap_8 FILLER_4_164 ();
 sg13g2_decap_8 FILLER_4_171 ();
 sg13g2_decap_8 FILLER_4_178 ();
 sg13g2_decap_4 FILLER_4_185 ();
 sg13g2_decap_8 FILLER_5_24 ();
 sg13g2_fill_1 FILLER_5_31 ();
 sg13g2_fill_2 FILLER_5_40 ();
 sg13g2_fill_2 FILLER_5_97 ();
 sg13g2_fill_1 FILLER_5_99 ();
 sg13g2_decap_8 FILLER_5_176 ();
 sg13g2_fill_2 FILLER_5_183 ();
 sg13g2_fill_1 FILLER_6_16 ();
 sg13g2_fill_2 FILLER_6_25 ();
 sg13g2_fill_1 FILLER_6_27 ();
 sg13g2_decap_8 FILLER_6_45 ();
 sg13g2_fill_2 FILLER_6_52 ();
 sg13g2_fill_1 FILLER_6_54 ();
 sg13g2_fill_2 FILLER_6_72 ();
 sg13g2_decap_4 FILLER_6_99 ();
 sg13g2_decap_4 FILLER_6_120 ();
 sg13g2_fill_1 FILLER_6_124 ();
 sg13g2_fill_1 FILLER_6_146 ();
 sg13g2_decap_4 FILLER_6_172 ();
 sg13g2_fill_2 FILLER_6_176 ();
 sg13g2_fill_2 FILLER_6_195 ();
 sg13g2_fill_1 FILLER_7_41 ();
 sg13g2_fill_1 FILLER_7_59 ();
 sg13g2_decap_4 FILLER_7_115 ();
 sg13g2_fill_2 FILLER_7_119 ();
 sg13g2_fill_1 FILLER_7_189 ();
 sg13g2_fill_2 FILLER_7_194 ();
 sg13g2_fill_1 FILLER_7_196 ();
 sg13g2_fill_2 FILLER_8_0 ();
 sg13g2_fill_1 FILLER_8_36 ();
 sg13g2_fill_1 FILLER_8_54 ();
 sg13g2_decap_4 FILLER_8_72 ();
 sg13g2_fill_1 FILLER_8_76 ();
 sg13g2_fill_1 FILLER_8_94 ();
 sg13g2_decap_4 FILLER_8_112 ();
 sg13g2_fill_2 FILLER_8_150 ();
 sg13g2_fill_1 FILLER_8_152 ();
 sg13g2_fill_2 FILLER_8_178 ();
 sg13g2_fill_2 FILLER_9_25 ();
 sg13g2_fill_2 FILLER_9_94 ();
 sg13g2_fill_1 FILLER_9_113 ();
 sg13g2_decap_8 FILLER_9_135 ();
 sg13g2_fill_1 FILLER_9_146 ();
 sg13g2_fill_2 FILLER_10_4 ();
 sg13g2_fill_1 FILLER_10_6 ();
 sg13g2_fill_2 FILLER_10_28 ();
 sg13g2_fill_2 FILLER_10_55 ();
 sg13g2_decap_4 FILLER_10_61 ();
 sg13g2_fill_1 FILLER_10_65 ();
 sg13g2_decap_8 FILLER_10_108 ();
 sg13g2_fill_1 FILLER_10_115 ();
 sg13g2_fill_2 FILLER_10_141 ();
 sg13g2_fill_1 FILLER_10_143 ();
 sg13g2_fill_2 FILLER_10_194 ();
 sg13g2_fill_1 FILLER_10_196 ();
 sg13g2_fill_2 FILLER_11_4 ();
 sg13g2_fill_1 FILLER_11_6 ();
 sg13g2_fill_1 FILLER_11_15 ();
 sg13g2_fill_1 FILLER_11_54 ();
 sg13g2_decap_8 FILLER_11_76 ();
 sg13g2_decap_8 FILLER_11_83 ();
 sg13g2_decap_8 FILLER_11_90 ();
 sg13g2_fill_2 FILLER_11_97 ();
 sg13g2_fill_2 FILLER_11_154 ();
 sg13g2_fill_1 FILLER_11_173 ();
 sg13g2_fill_2 FILLER_11_195 ();
 sg13g2_fill_1 FILLER_12_88 ();
 sg13g2_fill_2 FILLER_12_127 ();
 sg13g2_fill_1 FILLER_12_146 ();
 sg13g2_fill_2 FILLER_12_172 ();
 sg13g2_fill_2 FILLER_12_191 ();
 sg13g2_fill_2 FILLER_13_8 ();
 sg13g2_fill_1 FILLER_13_31 ();
 sg13g2_fill_2 FILLER_13_57 ();
 sg13g2_fill_1 FILLER_13_59 ();
 sg13g2_decap_8 FILLER_13_102 ();
 sg13g2_decap_4 FILLER_13_151 ();
 sg13g2_fill_1 FILLER_14_37 ();
 sg13g2_fill_2 FILLER_14_71 ();
 sg13g2_decap_8 FILLER_14_94 ();
 sg13g2_decap_8 FILLER_14_101 ();
 sg13g2_fill_2 FILLER_14_108 ();
 sg13g2_fill_2 FILLER_14_194 ();
 sg13g2_fill_1 FILLER_14_196 ();
 sg13g2_fill_1 FILLER_15_29 ();
 sg13g2_fill_1 FILLER_15_47 ();
 sg13g2_fill_2 FILLER_15_65 ();
 sg13g2_fill_1 FILLER_15_67 ();
 sg13g2_decap_8 FILLER_15_80 ();
 sg13g2_fill_1 FILLER_15_121 ();
 sg13g2_decap_8 FILLER_15_139 ();
 sg13g2_fill_2 FILLER_15_146 ();
 sg13g2_fill_1 FILLER_15_148 ();
 sg13g2_fill_1 FILLER_15_174 ();
 sg13g2_fill_1 FILLER_15_196 ();
 sg13g2_fill_1 FILLER_16_12 ();
 sg13g2_fill_2 FILLER_16_42 ();
 sg13g2_fill_2 FILLER_16_90 ();
 sg13g2_fill_1 FILLER_16_96 ();
 sg13g2_decap_4 FILLER_16_118 ();
 sg13g2_fill_1 FILLER_16_122 ();
 sg13g2_fill_1 FILLER_16_182 ();
 sg13g2_fill_1 FILLER_16_200 ();
 sg13g2_fill_2 FILLER_17_0 ();
 sg13g2_fill_2 FILLER_17_95 ();
 sg13g2_fill_1 FILLER_17_97 ();
 sg13g2_fill_1 FILLER_17_119 ();
 sg13g2_decap_4 FILLER_17_141 ();
 sg13g2_fill_2 FILLER_17_145 ();
 sg13g2_fill_2 FILLER_17_176 ();
 sg13g2_fill_2 FILLER_17_199 ();
 sg13g2_fill_1 FILLER_18_0 ();
 sg13g2_fill_1 FILLER_18_18 ();
 sg13g2_fill_1 FILLER_18_61 ();
 sg13g2_fill_1 FILLER_18_66 ();
 sg13g2_fill_1 FILLER_18_101 ();
 sg13g2_fill_1 FILLER_18_123 ();
 sg13g2_fill_2 FILLER_18_141 ();
 sg13g2_fill_1 FILLER_18_143 ();
 sg13g2_fill_2 FILLER_18_199 ();
 sg13g2_fill_1 FILLER_19_4 ();
 sg13g2_fill_2 FILLER_19_22 ();
 sg13g2_fill_1 FILLER_19_24 ();
 sg13g2_fill_1 FILLER_19_58 ();
 sg13g2_fill_2 FILLER_19_63 ();
 sg13g2_fill_1 FILLER_19_82 ();
 sg13g2_decap_4 FILLER_19_121 ();
 sg13g2_fill_2 FILLER_19_163 ();
 sg13g2_fill_1 FILLER_19_165 ();
 sg13g2_fill_2 FILLER_19_199 ();
 sg13g2_fill_1 FILLER_20_17 ();
 sg13g2_fill_1 FILLER_20_39 ();
 sg13g2_fill_2 FILLER_20_78 ();
 sg13g2_fill_2 FILLER_20_105 ();
 sg13g2_decap_4 FILLER_20_124 ();
 sg13g2_fill_2 FILLER_20_166 ();
 sg13g2_fill_1 FILLER_21_21 ();
 sg13g2_fill_2 FILLER_21_55 ();
 sg13g2_fill_1 FILLER_21_95 ();
 sg13g2_decap_8 FILLER_21_100 ();
 sg13g2_decap_4 FILLER_21_107 ();
 sg13g2_decap_8 FILLER_21_128 ();
 sg13g2_fill_1 FILLER_21_139 ();
 sg13g2_fill_2 FILLER_21_194 ();
 sg13g2_fill_1 FILLER_21_196 ();
 sg13g2_fill_2 FILLER_22_45 ();
 sg13g2_fill_1 FILLER_22_64 ();
 sg13g2_decap_8 FILLER_22_90 ();
 sg13g2_fill_2 FILLER_22_97 ();
 sg13g2_fill_1 FILLER_22_171 ();
 sg13g2_fill_1 FILLER_23_0 ();
 sg13g2_fill_2 FILLER_23_43 ();
 sg13g2_fill_2 FILLER_23_98 ();
 sg13g2_decap_8 FILLER_23_117 ();
 sg13g2_decap_8 FILLER_23_124 ();
 sg13g2_fill_2 FILLER_23_131 ();
 sg13g2_fill_1 FILLER_23_143 ();
 sg13g2_fill_2 FILLER_23_149 ();
 sg13g2_fill_2 FILLER_23_176 ();
 sg13g2_fill_2 FILLER_23_199 ();
 sg13g2_fill_2 FILLER_24_21 ();
 sg13g2_fill_1 FILLER_24_23 ();
 sg13g2_fill_1 FILLER_24_62 ();
 sg13g2_fill_2 FILLER_24_126 ();
 sg13g2_fill_1 FILLER_24_155 ();
 sg13g2_fill_2 FILLER_25_25 ();
 sg13g2_fill_1 FILLER_25_27 ();
 sg13g2_fill_1 FILLER_25_45 ();
 sg13g2_decap_4 FILLER_25_109 ();
 sg13g2_fill_2 FILLER_25_178 ();
 sg13g2_fill_2 FILLER_26_37 ();
 sg13g2_fill_2 FILLER_26_61 ();
 sg13g2_fill_1 FILLER_26_63 ();
 sg13g2_fill_2 FILLER_26_115 ();
 sg13g2_fill_2 FILLER_26_159 ();
 sg13g2_fill_2 FILLER_27_4 ();
 sg13g2_fill_1 FILLER_27_6 ();
 sg13g2_fill_2 FILLER_27_83 ();
 sg13g2_fill_2 FILLER_27_106 ();
 sg13g2_fill_1 FILLER_27_108 ();
 sg13g2_decap_4 FILLER_27_126 ();
 sg13g2_fill_1 FILLER_27_143 ();
 sg13g2_fill_2 FILLER_27_178 ();
 sg13g2_fill_1 FILLER_27_200 ();
 sg13g2_fill_2 FILLER_28_4 ();
 sg13g2_fill_1 FILLER_28_6 ();
 sg13g2_fill_2 FILLER_28_53 ();
 sg13g2_fill_1 FILLER_28_55 ();
 sg13g2_fill_2 FILLER_28_106 ();
 sg13g2_fill_1 FILLER_28_108 ();
 sg13g2_fill_1 FILLER_28_151 ();
 sg13g2_fill_1 FILLER_29_0 ();
 sg13g2_fill_2 FILLER_29_47 ();
 sg13g2_fill_1 FILLER_29_49 ();
 sg13g2_fill_2 FILLER_29_67 ();
 sg13g2_fill_2 FILLER_29_94 ();
 sg13g2_fill_1 FILLER_29_96 ();
 sg13g2_fill_1 FILLER_29_131 ();
 sg13g2_fill_2 FILLER_29_157 ();
 sg13g2_fill_2 FILLER_29_179 ();
 sg13g2_fill_1 FILLER_29_200 ();
 sg13g2_fill_1 FILLER_30_0 ();
 sg13g2_fill_2 FILLER_30_51 ();
 sg13g2_fill_2 FILLER_30_124 ();
 sg13g2_fill_2 FILLER_31_4 ();
 sg13g2_fill_1 FILLER_31_6 ();
 sg13g2_fill_1 FILLER_31_32 ();
 sg13g2_fill_2 FILLER_31_37 ();
 sg13g2_fill_2 FILLER_31_64 ();
 sg13g2_fill_1 FILLER_31_66 ();
 sg13g2_fill_1 FILLER_31_105 ();
 sg13g2_decap_4 FILLER_31_123 ();
 sg13g2_fill_2 FILLER_31_127 ();
 sg13g2_fill_2 FILLER_31_133 ();
 sg13g2_fill_2 FILLER_32_0 ();
 sg13g2_fill_2 FILLER_32_41 ();
 sg13g2_fill_1 FILLER_32_47 ();
 sg13g2_fill_2 FILLER_32_107 ();
 sg13g2_fill_2 FILLER_32_138 ();
 sg13g2_fill_1 FILLER_32_140 ();
 sg13g2_fill_1 FILLER_32_200 ();
 sg13g2_fill_2 FILLER_33_0 ();
 sg13g2_fill_1 FILLER_33_2 ();
 sg13g2_fill_1 FILLER_33_71 ();
 sg13g2_fill_1 FILLER_33_97 ();
 sg13g2_fill_2 FILLER_33_127 ();
 sg13g2_fill_2 FILLER_33_168 ();
 sg13g2_fill_2 FILLER_33_199 ();
 sg13g2_fill_2 FILLER_34_49 ();
 sg13g2_fill_2 FILLER_34_85 ();
 sg13g2_fill_2 FILLER_34_121 ();
 sg13g2_fill_1 FILLER_34_123 ();
 sg13g2_fill_2 FILLER_34_141 ();
 sg13g2_fill_1 FILLER_34_143 ();
 sg13g2_fill_1 FILLER_34_161 ();
 sg13g2_fill_2 FILLER_35_0 ();
 sg13g2_fill_1 FILLER_35_2 ();
 sg13g2_fill_2 FILLER_35_20 ();
 sg13g2_fill_2 FILLER_35_27 ();
 sg13g2_fill_2 FILLER_35_135 ();
 sg13g2_fill_1 FILLER_35_200 ();
 sg13g2_fill_2 FILLER_36_12 ();
 sg13g2_fill_2 FILLER_36_55 ();
 sg13g2_fill_2 FILLER_36_78 ();
 sg13g2_fill_1 FILLER_36_80 ();
 sg13g2_fill_2 FILLER_36_110 ();
 sg13g2_fill_1 FILLER_36_112 ();
 sg13g2_decap_4 FILLER_36_130 ();
 sg13g2_fill_1 FILLER_36_134 ();
 sg13g2_fill_2 FILLER_36_144 ();
 sg13g2_fill_1 FILLER_36_196 ();
 sg13g2_fill_2 FILLER_37_0 ();
 sg13g2_fill_2 FILLER_37_85 ();
 sg13g2_fill_2 FILLER_37_112 ();
 sg13g2_fill_1 FILLER_37_114 ();
 sg13g2_decap_4 FILLER_37_119 ();
 sg13g2_fill_2 FILLER_37_163 ();
 sg13g2_fill_2 FILLER_37_191 ();
 sg13g2_fill_1 FILLER_38_122 ();
 sg13g2_fill_2 FILLER_38_179 ();
 sg13g2_fill_2 FILLER_39_0 ();
 sg13g2_fill_2 FILLER_39_56 ();
 sg13g2_fill_1 FILLER_39_75 ();
 sg13g2_fill_2 FILLER_39_110 ();
 sg13g2_fill_2 FILLER_39_129 ();
 sg13g2_fill_1 FILLER_39_182 ();
 sg13g2_fill_1 FILLER_39_200 ();
 sg13g2_fill_2 FILLER_40_68 ();
 sg13g2_fill_1 FILLER_40_82 ();
 sg13g2_fill_1 FILLER_40_87 ();
 sg13g2_fill_1 FILLER_40_109 ();
 sg13g2_decap_8 FILLER_40_118 ();
 sg13g2_decap_4 FILLER_40_125 ();
 sg13g2_fill_2 FILLER_40_171 ();
 sg13g2_fill_1 FILLER_40_173 ();
 sg13g2_fill_2 FILLER_40_199 ();
 sg13g2_fill_1 FILLER_41_62 ();
 sg13g2_fill_1 FILLER_41_77 ();
 sg13g2_fill_1 FILLER_41_150 ();
 sg13g2_fill_2 FILLER_41_176 ();
 sg13g2_fill_2 FILLER_41_199 ();
 sg13g2_decap_8 FILLER_42_105 ();
 sg13g2_decap_4 FILLER_42_112 ();
 sg13g2_fill_2 FILLER_42_116 ();
 sg13g2_fill_2 FILLER_42_152 ();
 sg13g2_fill_1 FILLER_42_154 ();
 sg13g2_fill_2 FILLER_42_199 ();
 sg13g2_fill_2 FILLER_43_8 ();
 sg13g2_fill_1 FILLER_43_10 ();
 sg13g2_fill_1 FILLER_43_45 ();
 sg13g2_decap_8 FILLER_43_105 ();
 sg13g2_fill_1 FILLER_43_112 ();
 sg13g2_fill_1 FILLER_43_134 ();
 sg13g2_fill_2 FILLER_43_156 ();
 sg13g2_fill_1 FILLER_43_188 ();
 sg13g2_fill_1 FILLER_44_8 ();
 sg13g2_fill_2 FILLER_44_26 ();
 sg13g2_fill_1 FILLER_44_90 ();
 sg13g2_fill_1 FILLER_44_151 ();
 sg13g2_fill_1 FILLER_44_200 ();
 sg13g2_fill_2 FILLER_45_8 ();
 sg13g2_fill_2 FILLER_45_31 ();
 sg13g2_fill_1 FILLER_45_33 ();
 sg13g2_fill_2 FILLER_45_140 ();
 sg13g2_fill_2 FILLER_46_8 ();
 sg13g2_fill_2 FILLER_46_35 ();
 sg13g2_fill_1 FILLER_46_37 ();
 sg13g2_fill_2 FILLER_46_98 ();
 sg13g2_fill_1 FILLER_46_100 ();
 sg13g2_fill_2 FILLER_46_146 ();
 sg13g2_fill_2 FILLER_46_199 ();
 sg13g2_fill_2 FILLER_47_75 ();
 sg13g2_fill_1 FILLER_47_77 ();
 sg13g2_fill_2 FILLER_47_116 ();
 sg13g2_fill_1 FILLER_47_118 ();
 sg13g2_fill_1 FILLER_47_173 ();
 sg13g2_fill_1 FILLER_47_178 ();
 sg13g2_fill_1 FILLER_47_200 ();
 sg13g2_fill_2 FILLER_48_38 ();
 sg13g2_decap_8 FILLER_48_65 ();
 sg13g2_fill_1 FILLER_48_72 ();
 sg13g2_decap_4 FILLER_48_81 ();
 sg13g2_fill_1 FILLER_48_85 ();
 sg13g2_decap_8 FILLER_48_90 ();
 sg13g2_fill_1 FILLER_48_97 ();
 sg13g2_fill_2 FILLER_48_123 ();
 sg13g2_fill_2 FILLER_48_146 ();
 sg13g2_fill_1 FILLER_48_156 ();
 sg13g2_fill_1 FILLER_48_161 ();
 sg13g2_fill_1 FILLER_48_200 ();
 sg13g2_fill_1 FILLER_49_12 ();
 sg13g2_decap_4 FILLER_49_98 ();
 sg13g2_fill_1 FILLER_49_102 ();
 sg13g2_fill_1 FILLER_49_163 ();
 sg13g2_fill_1 FILLER_49_181 ();
 sg13g2_fill_2 FILLER_49_199 ();
 sg13g2_fill_2 FILLER_50_12 ();
 sg13g2_fill_2 FILLER_50_64 ();
 sg13g2_decap_8 FILLER_50_104 ();
 sg13g2_fill_2 FILLER_50_155 ();
 sg13g2_fill_2 FILLER_50_174 ();
 sg13g2_fill_2 FILLER_51_12 ();
 sg13g2_decap_4 FILLER_51_35 ();
 sg13g2_fill_2 FILLER_51_70 ();
 sg13g2_fill_1 FILLER_51_72 ();
 sg13g2_decap_8 FILLER_51_106 ();
 sg13g2_decap_4 FILLER_51_113 ();
 sg13g2_fill_1 FILLER_51_117 ();
 sg13g2_fill_2 FILLER_51_137 ();
 sg13g2_fill_1 FILLER_51_139 ();
 sg13g2_fill_2 FILLER_51_173 ();
 sg13g2_fill_1 FILLER_51_175 ();
 sg13g2_fill_1 FILLER_52_34 ();
 sg13g2_fill_2 FILLER_52_39 ();
 sg13g2_fill_2 FILLER_52_63 ();
 sg13g2_decap_8 FILLER_52_120 ();
 sg13g2_fill_2 FILLER_52_127 ();
 sg13g2_fill_1 FILLER_52_129 ();
 sg13g2_fill_1 FILLER_52_196 ();
 sg13g2_fill_2 FILLER_53_0 ();
 sg13g2_fill_1 FILLER_53_23 ();
 sg13g2_decap_4 FILLER_53_62 ();
 sg13g2_fill_1 FILLER_53_66 ();
 sg13g2_decap_4 FILLER_53_101 ();
 sg13g2_fill_1 FILLER_53_105 ();
 sg13g2_fill_1 FILLER_53_159 ();
 sg13g2_fill_2 FILLER_53_194 ();
 sg13g2_fill_1 FILLER_53_196 ();
 sg13g2_fill_2 FILLER_54_12 ();
 sg13g2_decap_4 FILLER_54_83 ();
 sg13g2_fill_1 FILLER_54_87 ();
 sg13g2_fill_2 FILLER_54_195 ();
 sg13g2_fill_1 FILLER_55_8 ();
 sg13g2_fill_2 FILLER_55_30 ();
 sg13g2_fill_1 FILLER_55_32 ();
 sg13g2_fill_1 FILLER_55_53 ();
 sg13g2_decap_4 FILLER_55_75 ();
 sg13g2_fill_1 FILLER_55_79 ();
 sg13g2_fill_2 FILLER_55_97 ();
 sg13g2_fill_1 FILLER_55_99 ();
 sg13g2_decap_4 FILLER_55_129 ();
 sg13g2_fill_2 FILLER_55_133 ();
 sg13g2_fill_2 FILLER_55_195 ();
 sg13g2_fill_2 FILLER_56_8 ();
 sg13g2_fill_1 FILLER_56_10 ();
 sg13g2_fill_1 FILLER_56_32 ();
 sg13g2_fill_2 FILLER_56_93 ();
 sg13g2_decap_4 FILLER_56_99 ();
 sg13g2_fill_1 FILLER_56_103 ();
 sg13g2_fill_1 FILLER_56_181 ();
 sg13g2_fill_2 FILLER_56_199 ();
 sg13g2_decap_8 FILLER_57_8 ();
 sg13g2_fill_1 FILLER_57_15 ();
 sg13g2_fill_2 FILLER_57_56 ();
 sg13g2_fill_1 FILLER_57_64 ();
 sg13g2_fill_1 FILLER_57_82 ();
 sg13g2_fill_1 FILLER_57_108 ();
 sg13g2_decap_4 FILLER_57_113 ();
 sg13g2_decap_4 FILLER_57_121 ();
 sg13g2_fill_2 FILLER_57_125 ();
 sg13g2_fill_1 FILLER_57_148 ();
 sg13g2_fill_1 FILLER_57_153 ();
 sg13g2_fill_2 FILLER_57_171 ();
 sg13g2_fill_1 FILLER_57_173 ();
 sg13g2_fill_2 FILLER_57_195 ();
 sg13g2_decap_8 FILLER_58_8 ();
 sg13g2_decap_8 FILLER_58_15 ();
 sg13g2_decap_4 FILLER_58_22 ();
 sg13g2_fill_2 FILLER_58_26 ();
 sg13g2_fill_2 FILLER_58_72 ();
 sg13g2_decap_4 FILLER_58_129 ();
 sg13g2_fill_1 FILLER_58_133 ();
 sg13g2_decap_8 FILLER_58_155 ();
 sg13g2_decap_4 FILLER_58_162 ();
 sg13g2_fill_2 FILLER_58_166 ();
 sg13g2_fill_1 FILLER_59_0 ();
 sg13g2_decap_8 FILLER_59_18 ();
 sg13g2_fill_1 FILLER_59_29 ();
 sg13g2_fill_2 FILLER_59_67 ();
 sg13g2_fill_1 FILLER_59_69 ();
 sg13g2_decap_4 FILLER_59_122 ();
 sg13g2_decap_8 FILLER_59_164 ();
 sg13g2_fill_2 FILLER_59_171 ();
 sg13g2_fill_2 FILLER_59_190 ();
 sg13g2_fill_1 FILLER_59_192 ();
 sg13g2_decap_4 FILLER_60_0 ();
 sg13g2_decap_8 FILLER_60_42 ();
 sg13g2_fill_1 FILLER_60_49 ();
 sg13g2_decap_4 FILLER_60_91 ();
 sg13g2_fill_1 FILLER_60_95 ();
 sg13g2_fill_1 FILLER_60_99 ();
 sg13g2_fill_2 FILLER_60_117 ();
 sg13g2_fill_1 FILLER_60_119 ();
 sg13g2_decap_4 FILLER_60_171 ();
 sg13g2_fill_1 FILLER_60_192 ();
 sg13g2_decap_8 FILLER_61_0 ();
 sg13g2_fill_2 FILLER_61_7 ();
 sg13g2_decap_8 FILLER_61_51 ();
 sg13g2_decap_8 FILLER_61_58 ();
 sg13g2_decap_4 FILLER_61_65 ();
 sg13g2_fill_1 FILLER_61_69 ();
 sg13g2_decap_8 FILLER_61_74 ();
 sg13g2_fill_1 FILLER_61_81 ();
 sg13g2_fill_2 FILLER_61_86 ();
 sg13g2_fill_2 FILLER_61_92 ();
 sg13g2_fill_1 FILLER_61_94 ();
 sg13g2_decap_8 FILLER_61_103 ();
 sg13g2_decap_8 FILLER_61_110 ();
 sg13g2_decap_4 FILLER_61_117 ();
 sg13g2_fill_1 FILLER_61_121 ();
 sg13g2_decap_8 FILLER_61_139 ();
 sg13g2_decap_4 FILLER_61_146 ();
 sg13g2_decap_4 FILLER_61_188 ();
 sg13g2_fill_1 FILLER_61_192 ();
 sg13g2_decap_8 FILLER_62_0 ();
 sg13g2_decap_8 FILLER_62_7 ();
 sg13g2_decap_8 FILLER_62_14 ();
 sg13g2_decap_4 FILLER_62_21 ();
 sg13g2_fill_2 FILLER_62_25 ();
 sg13g2_decap_4 FILLER_62_31 ();
 sg13g2_fill_1 FILLER_62_85 ();
 sg13g2_fill_1 FILLER_62_90 ();
 sg13g2_decap_8 FILLER_62_129 ();
 sg13g2_decap_4 FILLER_62_136 ();
 sg13g2_fill_1 FILLER_62_140 ();
 sg13g2_decap_8 FILLER_62_166 ();
 sg13g2_fill_2 FILLER_62_173 ();
 sg13g2_fill_1 FILLER_62_200 ();
 sg13g2_decap_8 FILLER_63_0 ();
 sg13g2_fill_1 FILLER_63_7 ();
 sg13g2_decap_4 FILLER_63_25 ();
 sg13g2_decap_4 FILLER_63_46 ();
 sg13g2_fill_1 FILLER_63_50 ();
 sg13g2_fill_2 FILLER_63_85 ();
 sg13g2_decap_8 FILLER_63_129 ();
 sg13g2_fill_1 FILLER_63_136 ();
 sg13g2_decap_8 FILLER_63_175 ();
 sg13g2_decap_8 FILLER_63_182 ();
 sg13g2_decap_8 FILLER_64_0 ();
 sg13g2_fill_2 FILLER_64_7 ();
 sg13g2_fill_2 FILLER_64_26 ();
 sg13g2_fill_1 FILLER_64_28 ();
 sg13g2_decap_8 FILLER_64_46 ();
 sg13g2_decap_8 FILLER_64_53 ();
 sg13g2_decap_4 FILLER_64_60 ();
 sg13g2_fill_1 FILLER_64_64 ();
 sg13g2_fill_1 FILLER_64_103 ();
 sg13g2_fill_1 FILLER_64_108 ();
 sg13g2_fill_1 FILLER_64_117 ();
 sg13g2_decap_8 FILLER_64_173 ();
 sg13g2_decap_4 FILLER_65_8 ();
 sg13g2_fill_2 FILLER_65_12 ();
 sg13g2_decap_8 FILLER_65_18 ();
 sg13g2_decap_8 FILLER_65_25 ();
 sg13g2_fill_2 FILLER_65_32 ();
 sg13g2_decap_8 FILLER_65_68 ();
 sg13g2_decap_4 FILLER_65_75 ();
 sg13g2_fill_1 FILLER_65_79 ();
 sg13g2_decap_8 FILLER_65_118 ();
 sg13g2_fill_1 FILLER_65_125 ();
 sg13g2_decap_8 FILLER_65_143 ();
 sg13g2_fill_1 FILLER_65_188 ();
 sg13g2_fill_1 FILLER_66_8 ();
 sg13g2_decap_4 FILLER_66_42 ();
 sg13g2_fill_2 FILLER_66_46 ();
 sg13g2_fill_1 FILLER_66_86 ();
 sg13g2_fill_2 FILLER_66_122 ();
 sg13g2_fill_1 FILLER_66_124 ();
 sg13g2_fill_1 FILLER_66_176 ();
 sg13g2_fill_2 FILLER_66_194 ();
 sg13g2_fill_1 FILLER_66_196 ();
 sg13g2_decap_4 FILLER_67_21 ();
 sg13g2_decap_8 FILLER_67_63 ();
 sg13g2_fill_1 FILLER_67_70 ();
 sg13g2_fill_2 FILLER_67_194 ();
 sg13g2_fill_1 FILLER_67_196 ();
 sg13g2_fill_2 FILLER_68_4 ();
 sg13g2_fill_1 FILLER_68_6 ();
 sg13g2_fill_2 FILLER_68_11 ();
 sg13g2_fill_1 FILLER_68_13 ();
 sg13g2_fill_2 FILLER_68_35 ();
 sg13g2_fill_1 FILLER_68_37 ();
 sg13g2_fill_1 FILLER_68_55 ();
 sg13g2_fill_1 FILLER_68_77 ();
 sg13g2_fill_1 FILLER_68_83 ();
 sg13g2_decap_8 FILLER_68_101 ();
 sg13g2_decap_4 FILLER_68_108 ();
 sg13g2_fill_2 FILLER_68_112 ();
 sg13g2_decap_8 FILLER_68_122 ();
 sg13g2_fill_2 FILLER_68_129 ();
 sg13g2_fill_2 FILLER_68_177 ();
 sg13g2_fill_1 FILLER_68_200 ();
 sg13g2_fill_1 FILLER_69_4 ();
 sg13g2_decap_8 FILLER_69_72 ();
 sg13g2_decap_4 FILLER_69_79 ();
 sg13g2_fill_1 FILLER_69_83 ();
 sg13g2_fill_1 FILLER_69_126 ();
 sg13g2_fill_2 FILLER_69_198 ();
 sg13g2_fill_1 FILLER_69_200 ();
 sg13g2_fill_2 FILLER_70_0 ();
 sg13g2_fill_2 FILLER_70_49 ();
 sg13g2_fill_1 FILLER_70_51 ();
 sg13g2_decap_4 FILLER_70_107 ();
 sg13g2_fill_1 FILLER_70_111 ();
 sg13g2_fill_1 FILLER_70_146 ();
 sg13g2_fill_1 FILLER_70_164 ();
 sg13g2_fill_2 FILLER_70_182 ();
 sg13g2_fill_2 FILLER_71_0 ();
 sg13g2_fill_1 FILLER_71_27 ();
 sg13g2_fill_2 FILLER_71_53 ();
 sg13g2_fill_1 FILLER_71_55 ();
 sg13g2_fill_1 FILLER_71_73 ();
 sg13g2_fill_2 FILLER_71_95 ();
 sg13g2_fill_1 FILLER_71_97 ();
 sg13g2_decap_8 FILLER_71_119 ();
 sg13g2_fill_2 FILLER_71_126 ();
 sg13g2_fill_1 FILLER_71_128 ();
 sg13g2_fill_1 FILLER_71_192 ();
 sg13g2_fill_1 FILLER_72_4 ();
 sg13g2_fill_1 FILLER_72_22 ();
 sg13g2_decap_4 FILLER_72_48 ();
 sg13g2_fill_2 FILLER_72_73 ();
 sg13g2_fill_1 FILLER_72_75 ();
 sg13g2_decap_8 FILLER_72_97 ();
 sg13g2_decap_4 FILLER_72_104 ();
 sg13g2_fill_1 FILLER_72_167 ();
 sg13g2_decap_4 FILLER_73_62 ();
 sg13g2_fill_1 FILLER_73_66 ();
 sg13g2_fill_2 FILLER_73_88 ();
 sg13g2_fill_2 FILLER_73_145 ();
 sg13g2_fill_2 FILLER_73_198 ();
 sg13g2_fill_1 FILLER_73_200 ();
 sg13g2_fill_2 FILLER_74_0 ();
 sg13g2_fill_1 FILLER_74_2 ();
 sg13g2_fill_2 FILLER_74_20 ();
 sg13g2_fill_1 FILLER_74_22 ();
 sg13g2_decap_8 FILLER_74_82 ();
 sg13g2_fill_1 FILLER_74_89 ();
 sg13g2_fill_2 FILLER_74_138 ();
 sg13g2_fill_2 FILLER_74_157 ();
 sg13g2_fill_1 FILLER_74_159 ();
 sg13g2_fill_2 FILLER_74_198 ();
 sg13g2_fill_1 FILLER_74_200 ();
 sg13g2_fill_2 FILLER_75_8 ();
 sg13g2_fill_2 FILLER_75_56 ();
 sg13g2_fill_1 FILLER_75_96 ();
 sg13g2_fill_2 FILLER_75_108 ();
 sg13g2_decap_4 FILLER_75_114 ();
 sg13g2_fill_2 FILLER_75_118 ();
 sg13g2_fill_1 FILLER_75_128 ();
 sg13g2_fill_1 FILLER_75_146 ();
 sg13g2_fill_1 FILLER_75_181 ();
 sg13g2_fill_2 FILLER_75_199 ();
 sg13g2_fill_1 FILLER_76_21 ();
 sg13g2_fill_1 FILLER_76_68 ();
 sg13g2_fill_2 FILLER_76_77 ();
 sg13g2_fill_2 FILLER_76_96 ();
 sg13g2_fill_2 FILLER_76_123 ();
 sg13g2_fill_2 FILLER_76_159 ();
 sg13g2_fill_2 FILLER_76_199 ();
 sg13g2_fill_1 FILLER_77_8 ();
 sg13g2_fill_1 FILLER_77_47 ();
 sg13g2_fill_2 FILLER_77_65 ();
 sg13g2_decap_8 FILLER_77_71 ();
 sg13g2_decap_4 FILLER_77_78 ();
 sg13g2_fill_1 FILLER_77_120 ();
 sg13g2_fill_2 FILLER_77_129 ();
 sg13g2_fill_1 FILLER_77_139 ();
 sg13g2_fill_2 FILLER_77_175 ();
 sg13g2_fill_1 FILLER_77_177 ();
 sg13g2_fill_2 FILLER_77_199 ();
 sg13g2_fill_2 FILLER_78_21 ();
 sg13g2_fill_1 FILLER_78_23 ();
 sg13g2_fill_1 FILLER_78_91 ();
 sg13g2_decap_4 FILLER_78_109 ();
 sg13g2_fill_1 FILLER_78_113 ();
 sg13g2_fill_1 FILLER_78_139 ();
 sg13g2_fill_2 FILLER_78_178 ();
 sg13g2_fill_1 FILLER_78_180 ();
 sg13g2_fill_2 FILLER_78_198 ();
 sg13g2_fill_1 FILLER_78_200 ();
 sg13g2_fill_1 FILLER_79_4 ();
 sg13g2_fill_2 FILLER_79_47 ();
 sg13g2_fill_2 FILLER_79_108 ();
 sg13g2_fill_1 FILLER_79_148 ();
 sg13g2_fill_2 FILLER_79_199 ();
 sg13g2_fill_1 FILLER_80_21 ();
 sg13g2_fill_2 FILLER_80_43 ();
 sg13g2_fill_1 FILLER_80_45 ();
 sg13g2_fill_2 FILLER_80_88 ();
 sg13g2_fill_2 FILLER_80_111 ();
 sg13g2_fill_2 FILLER_80_138 ();
 sg13g2_fill_1 FILLER_80_178 ();
 sg13g2_fill_1 FILLER_80_196 ();
 sg13g2_fill_1 FILLER_81_4 ();
 sg13g2_fill_2 FILLER_81_26 ();
 sg13g2_fill_2 FILLER_81_93 ();
 sg13g2_fill_2 FILLER_81_112 ();
 sg13g2_decap_4 FILLER_81_118 ();
 sg13g2_fill_2 FILLER_81_168 ();
 sg13g2_fill_1 FILLER_81_170 ();
 sg13g2_fill_1 FILLER_81_196 ();
 sg13g2_fill_2 FILLER_82_0 ();
 sg13g2_fill_1 FILLER_82_2 ();
 sg13g2_fill_2 FILLER_82_45 ();
 sg13g2_fill_2 FILLER_82_90 ();
 sg13g2_fill_2 FILLER_82_113 ();
 sg13g2_fill_1 FILLER_82_115 ();
 sg13g2_fill_1 FILLER_82_153 ();
 sg13g2_fill_1 FILLER_82_200 ();
 sg13g2_fill_2 FILLER_83_8 ();
 sg13g2_fill_2 FILLER_83_56 ();
 sg13g2_fill_1 FILLER_83_58 ();
 sg13g2_fill_2 FILLER_83_84 ();
 sg13g2_decap_8 FILLER_83_107 ();
 sg13g2_fill_1 FILLER_83_114 ();
 sg13g2_fill_2 FILLER_83_157 ();
 sg13g2_fill_1 FILLER_83_159 ();
 sg13g2_fill_1 FILLER_83_177 ();
 sg13g2_fill_2 FILLER_83_195 ();
 sg13g2_fill_2 FILLER_84_0 ();
 sg13g2_fill_1 FILLER_84_2 ();
 sg13g2_fill_2 FILLER_84_28 ();
 sg13g2_decap_4 FILLER_84_106 ();
 sg13g2_fill_1 FILLER_84_143 ();
 sg13g2_fill_2 FILLER_84_199 ();
 sg13g2_fill_2 FILLER_85_12 ();
 sg13g2_fill_2 FILLER_85_35 ();
 sg13g2_fill_2 FILLER_85_54 ();
 sg13g2_fill_2 FILLER_85_68 ();
 sg13g2_fill_2 FILLER_85_87 ();
 sg13g2_fill_1 FILLER_85_89 ();
 sg13g2_decap_8 FILLER_85_107 ();
 sg13g2_decap_4 FILLER_85_114 ();
 sg13g2_fill_1 FILLER_85_118 ();
 sg13g2_fill_1 FILLER_85_140 ();
 sg13g2_fill_2 FILLER_85_170 ();
 sg13g2_fill_1 FILLER_86_4 ();
 sg13g2_fill_1 FILLER_86_85 ();
 sg13g2_fill_1 FILLER_86_128 ();
 sg13g2_fill_1 FILLER_86_200 ();
 sg13g2_fill_1 FILLER_87_0 ();
 sg13g2_fill_1 FILLER_87_63 ();
 sg13g2_fill_1 FILLER_87_85 ();
 sg13g2_fill_2 FILLER_87_158 ();
 sg13g2_fill_2 FILLER_87_198 ();
 sg13g2_fill_1 FILLER_87_200 ();
 sg13g2_fill_1 FILLER_88_25 ();
 sg13g2_fill_2 FILLER_88_93 ();
 sg13g2_fill_1 FILLER_88_95 ();
 sg13g2_fill_1 FILLER_88_113 ();
 sg13g2_fill_2 FILLER_88_139 ();
 sg13g2_fill_1 FILLER_88_162 ();
 sg13g2_fill_2 FILLER_88_167 ();
 sg13g2_fill_1 FILLER_88_169 ();
 sg13g2_fill_2 FILLER_88_187 ();
 sg13g2_fill_1 FILLER_88_189 ();
 sg13g2_fill_2 FILLER_88_194 ();
 sg13g2_fill_1 FILLER_88_196 ();
 sg13g2_fill_2 FILLER_89_0 ();
 sg13g2_fill_1 FILLER_89_74 ();
 sg13g2_decap_8 FILLER_89_100 ();
 sg13g2_fill_2 FILLER_89_124 ();
 sg13g2_fill_1 FILLER_89_130 ();
 sg13g2_fill_2 FILLER_89_198 ();
 sg13g2_fill_1 FILLER_89_200 ();
 sg13g2_fill_2 FILLER_90_0 ();
 sg13g2_fill_1 FILLER_90_2 ();
 sg13g2_fill_2 FILLER_90_20 ();
 sg13g2_fill_2 FILLER_90_85 ();
 sg13g2_decap_8 FILLER_90_108 ();
 sg13g2_fill_1 FILLER_90_115 ();
 sg13g2_fill_1 FILLER_90_137 ();
 sg13g2_fill_2 FILLER_90_159 ();
 sg13g2_fill_1 FILLER_90_161 ();
 sg13g2_fill_2 FILLER_90_191 ();
 sg13g2_fill_2 FILLER_91_29 ();
 sg13g2_fill_1 FILLER_91_31 ();
 sg13g2_fill_1 FILLER_91_61 ();
 sg13g2_fill_2 FILLER_91_84 ();
 sg13g2_fill_1 FILLER_91_107 ();
 sg13g2_fill_2 FILLER_91_129 ();
 sg13g2_fill_2 FILLER_91_148 ();
 sg13g2_fill_1 FILLER_91_150 ();
 sg13g2_fill_2 FILLER_91_172 ();
 sg13g2_fill_1 FILLER_91_174 ();
 sg13g2_fill_1 FILLER_91_200 ();
 sg13g2_fill_2 FILLER_92_4 ();
 sg13g2_fill_1 FILLER_92_6 ();
 sg13g2_fill_1 FILLER_92_15 ();
 sg13g2_fill_2 FILLER_92_54 ();
 sg13g2_fill_1 FILLER_92_56 ();
 sg13g2_fill_2 FILLER_92_74 ();
 sg13g2_fill_1 FILLER_92_76 ();
 sg13g2_fill_2 FILLER_92_136 ();
 sg13g2_fill_1 FILLER_92_138 ();
 sg13g2_fill_2 FILLER_92_164 ();
 sg13g2_fill_1 FILLER_92_166 ();
 sg13g2_fill_1 FILLER_92_196 ();
 sg13g2_fill_2 FILLER_93_49 ();
 sg13g2_fill_1 FILLER_93_51 ();
 sg13g2_decap_4 FILLER_93_101 ();
 sg13g2_fill_2 FILLER_93_109 ();
 sg13g2_fill_1 FILLER_93_111 ();
 sg13g2_fill_2 FILLER_93_163 ();
 sg13g2_fill_1 FILLER_93_165 ();
 sg13g2_fill_2 FILLER_93_176 ();
 sg13g2_fill_2 FILLER_93_199 ();
 sg13g2_fill_1 FILLER_94_0 ();
 sg13g2_fill_1 FILLER_94_56 ();
 sg13g2_fill_2 FILLER_94_82 ();
 sg13g2_fill_1 FILLER_94_84 ();
 sg13g2_fill_2 FILLER_94_119 ();
 sg13g2_fill_1 FILLER_94_196 ();
 sg13g2_fill_1 FILLER_95_0 ();
 sg13g2_fill_2 FILLER_95_39 ();
 sg13g2_fill_2 FILLER_95_96 ();
 sg13g2_fill_1 FILLER_95_144 ();
 sg13g2_fill_1 FILLER_95_157 ();
 sg13g2_fill_2 FILLER_95_175 ();
 sg13g2_fill_1 FILLER_96_21 ();
 sg13g2_fill_2 FILLER_96_67 ();
 sg13g2_fill_1 FILLER_96_111 ();
 sg13g2_fill_2 FILLER_96_133 ();
 sg13g2_fill_1 FILLER_96_135 ();
 sg13g2_fill_2 FILLER_96_157 ();
 sg13g2_fill_1 FILLER_96_159 ();
 sg13g2_fill_2 FILLER_96_194 ();
 sg13g2_fill_1 FILLER_96_196 ();
 sg13g2_fill_2 FILLER_97_12 ();
 sg13g2_fill_1 FILLER_97_14 ();
 sg13g2_fill_1 FILLER_97_83 ();
 sg13g2_decap_8 FILLER_97_105 ();
 sg13g2_decap_4 FILLER_97_112 ();
 sg13g2_fill_2 FILLER_97_116 ();
 sg13g2_fill_1 FILLER_98_21 ();
 sg13g2_fill_1 FILLER_98_93 ();
 sg13g2_fill_1 FILLER_98_111 ();
 sg13g2_fill_1 FILLER_98_133 ();
 sg13g2_fill_2 FILLER_99_0 ();
 sg13g2_fill_2 FILLER_99_48 ();
 sg13g2_fill_1 FILLER_99_50 ();
 sg13g2_fill_2 FILLER_99_106 ();
 sg13g2_fill_2 FILLER_99_125 ();
 sg13g2_fill_2 FILLER_100_8 ();
 sg13g2_fill_2 FILLER_100_44 ();
 sg13g2_fill_1 FILLER_100_46 ();
 sg13g2_fill_1 FILLER_100_81 ();
 sg13g2_fill_2 FILLER_100_141 ();
 sg13g2_fill_1 FILLER_100_143 ();
 sg13g2_fill_2 FILLER_101_17 ();
 sg13g2_fill_1 FILLER_101_62 ();
 sg13g2_fill_2 FILLER_101_138 ();
 sg13g2_fill_1 FILLER_101_140 ();
 sg13g2_fill_2 FILLER_102_26 ();
 sg13g2_fill_1 FILLER_102_65 ();
 sg13g2_fill_2 FILLER_102_95 ();
 sg13g2_fill_2 FILLER_102_101 ();
 sg13g2_fill_2 FILLER_102_128 ();
 sg13g2_fill_2 FILLER_102_198 ();
 sg13g2_fill_1 FILLER_102_200 ();
 sg13g2_fill_2 FILLER_103_0 ();
 sg13g2_fill_1 FILLER_103_2 ();
 sg13g2_fill_1 FILLER_103_32 ();
 sg13g2_fill_2 FILLER_103_100 ();
 sg13g2_fill_1 FILLER_103_102 ();
 sg13g2_fill_2 FILLER_103_107 ();
 sg13g2_fill_1 FILLER_103_109 ();
 sg13g2_fill_2 FILLER_103_158 ();
 sg13g2_fill_1 FILLER_103_160 ();
 sg13g2_fill_2 FILLER_103_186 ();
 sg13g2_fill_1 FILLER_103_188 ();
 sg13g2_fill_1 FILLER_104_4 ();
 sg13g2_fill_1 FILLER_104_116 ();
 sg13g2_fill_1 FILLER_104_142 ();
 sg13g2_fill_2 FILLER_104_198 ();
 sg13g2_fill_1 FILLER_104_200 ();
 sg13g2_fill_1 FILLER_105_81 ();
 sg13g2_fill_1 FILLER_105_103 ();
 sg13g2_fill_2 FILLER_105_125 ();
 sg13g2_fill_1 FILLER_105_127 ();
 sg13g2_fill_2 FILLER_105_167 ();
 sg13g2_fill_1 FILLER_105_169 ();
 sg13g2_fill_2 FILLER_105_199 ();
 sg13g2_fill_2 FILLER_106_0 ();
 sg13g2_fill_1 FILLER_106_2 ();
 sg13g2_fill_1 FILLER_106_72 ();
 sg13g2_fill_2 FILLER_106_101 ();
 sg13g2_fill_2 FILLER_106_124 ();
 sg13g2_fill_1 FILLER_106_126 ();
 sg13g2_fill_1 FILLER_106_177 ();
 sg13g2_fill_2 FILLER_106_199 ();
 sg13g2_fill_2 FILLER_107_0 ();
 sg13g2_fill_1 FILLER_107_2 ();
 sg13g2_fill_2 FILLER_107_58 ();
 sg13g2_decap_8 FILLER_107_94 ();
 sg13g2_decap_4 FILLER_107_101 ();
 sg13g2_fill_1 FILLER_107_126 ();
 sg13g2_fill_2 FILLER_107_131 ();
 sg13g2_fill_1 FILLER_107_133 ();
 sg13g2_fill_2 FILLER_107_161 ();
 sg13g2_fill_2 FILLER_108_0 ();
 sg13g2_fill_1 FILLER_108_2 ();
 sg13g2_fill_2 FILLER_108_20 ();
 sg13g2_fill_1 FILLER_108_86 ();
 sg13g2_decap_4 FILLER_108_125 ();
 sg13g2_fill_2 FILLER_108_137 ();
 sg13g2_fill_2 FILLER_108_148 ();
 sg13g2_fill_1 FILLER_108_150 ();
 sg13g2_fill_2 FILLER_109_12 ();
 sg13g2_fill_1 FILLER_109_14 ();
 sg13g2_fill_2 FILLER_109_78 ();
 sg13g2_fill_2 FILLER_109_118 ();
 sg13g2_fill_2 FILLER_109_169 ();
 sg13g2_fill_1 FILLER_109_171 ();
 sg13g2_fill_2 FILLER_110_0 ();
 sg13g2_fill_2 FILLER_110_40 ();
 sg13g2_fill_1 FILLER_110_64 ();
 sg13g2_fill_2 FILLER_110_141 ();
 sg13g2_fill_1 FILLER_110_143 ();
 sg13g2_fill_2 FILLER_110_199 ();
 sg13g2_fill_1 FILLER_111_4 ();
 sg13g2_fill_2 FILLER_111_30 ();
 sg13g2_fill_1 FILLER_111_32 ();
 sg13g2_fill_1 FILLER_111_50 ();
 sg13g2_fill_2 FILLER_111_59 ();
 sg13g2_fill_1 FILLER_111_61 ();
 sg13g2_fill_2 FILLER_111_113 ();
 sg13g2_fill_1 FILLER_111_115 ();
 sg13g2_fill_2 FILLER_111_198 ();
 sg13g2_fill_1 FILLER_111_200 ();
 sg13g2_fill_1 FILLER_112_0 ();
 sg13g2_fill_2 FILLER_112_89 ();
 sg13g2_fill_1 FILLER_112_91 ();
 sg13g2_fill_2 FILLER_112_129 ();
 sg13g2_fill_1 FILLER_112_131 ();
 sg13g2_fill_2 FILLER_112_166 ();
 sg13g2_fill_1 FILLER_112_168 ();
 sg13g2_fill_2 FILLER_112_190 ();
 sg13g2_fill_1 FILLER_112_192 ();
 sg13g2_fill_1 FILLER_113_58 ();
 sg13g2_fill_2 FILLER_113_97 ();
 sg13g2_decap_8 FILLER_113_130 ();
 sg13g2_decap_8 FILLER_113_137 ();
 sg13g2_decap_8 FILLER_113_144 ();
 sg13g2_fill_1 FILLER_113_168 ();
 sg13g2_fill_2 FILLER_113_190 ();
 sg13g2_fill_1 FILLER_113_192 ();
 sg13g2_fill_2 FILLER_114_4 ();
 sg13g2_fill_1 FILLER_114_6 ();
 sg13g2_fill_1 FILLER_114_15 ();
 sg13g2_fill_2 FILLER_114_75 ();
 sg13g2_fill_1 FILLER_114_77 ();
 sg13g2_fill_2 FILLER_114_116 ();
 sg13g2_fill_2 FILLER_114_198 ();
 sg13g2_fill_1 FILLER_114_200 ();
 sg13g2_fill_1 FILLER_115_33 ();
 sg13g2_decap_4 FILLER_115_55 ();
 sg13g2_fill_2 FILLER_115_59 ();
 sg13g2_decap_4 FILLER_115_78 ();
 sg13g2_fill_1 FILLER_115_82 ();
 sg13g2_fill_1 FILLER_115_95 ();
 sg13g2_decap_4 FILLER_115_159 ();
 sg13g2_fill_1 FILLER_115_180 ();
 sg13g2_decap_8 FILLER_116_53 ();
 sg13g2_decap_8 FILLER_116_60 ();
 sg13g2_decap_8 FILLER_116_67 ();
 sg13g2_decap_8 FILLER_116_74 ();
 sg13g2_decap_8 FILLER_116_81 ();
 sg13g2_decap_8 FILLER_116_88 ();
 sg13g2_decap_8 FILLER_116_95 ();
 sg13g2_decap_4 FILLER_116_102 ();
 sg13g2_fill_2 FILLER_116_161 ();
 sg13g2_decap_4 FILLER_116_180 ();
 sg13g2_fill_1 FILLER_116_184 ();
 sg13g2_decap_8 FILLER_117_32 ();
 sg13g2_decap_8 FILLER_117_39 ();
 sg13g2_decap_8 FILLER_117_46 ();
 sg13g2_decap_8 FILLER_117_53 ();
 sg13g2_decap_8 FILLER_117_60 ();
 sg13g2_decap_8 FILLER_117_67 ();
 sg13g2_decap_8 FILLER_117_74 ();
 sg13g2_decap_8 FILLER_117_81 ();
 sg13g2_decap_8 FILLER_117_88 ();
 sg13g2_decap_8 FILLER_117_95 ();
 sg13g2_decap_4 FILLER_117_102 ();
 sg13g2_decap_8 FILLER_117_123 ();
 sg13g2_decap_8 FILLER_117_130 ();
 sg13g2_decap_8 FILLER_117_154 ();
 sg13g2_decap_4 FILLER_117_161 ();
 sg13g2_decap_8 FILLER_117_169 ();
 sg13g2_decap_8 FILLER_117_176 ();
 sg13g2_decap_4 FILLER_117_183 ();
 sg13g2_fill_2 FILLER_117_187 ();
 sg13g2_decap_8 FILLER_118_20 ();
 sg13g2_decap_8 FILLER_118_27 ();
 sg13g2_decap_8 FILLER_118_34 ();
 sg13g2_decap_8 FILLER_118_41 ();
 sg13g2_decap_8 FILLER_118_48 ();
 sg13g2_decap_8 FILLER_118_55 ();
 sg13g2_decap_4 FILLER_118_62 ();
 sg13g2_fill_2 FILLER_118_66 ();
 sg13g2_decap_8 FILLER_118_76 ();
 sg13g2_decap_8 FILLER_118_83 ();
 sg13g2_decap_8 FILLER_118_90 ();
 sg13g2_decap_8 FILLER_118_97 ();
 sg13g2_decap_8 FILLER_118_104 ();
 sg13g2_decap_8 FILLER_118_111 ();
 sg13g2_decap_8 FILLER_118_118 ();
 sg13g2_decap_8 FILLER_118_125 ();
 sg13g2_decap_8 FILLER_118_132 ();
 sg13g2_decap_8 FILLER_118_139 ();
 sg13g2_decap_8 FILLER_118_146 ();
 sg13g2_decap_8 FILLER_118_153 ();
 sg13g2_decap_8 FILLER_118_160 ();
 sg13g2_decap_8 FILLER_118_167 ();
 sg13g2_decap_8 FILLER_118_174 ();
 sg13g2_decap_8 FILLER_118_181 ();
 sg13g2_decap_4 FILLER_118_188 ();
 sg13g2_fill_1 FILLER_118_192 ();
 sg13g2_decap_8 FILLER_119_20 ();
 sg13g2_decap_8 FILLER_119_27 ();
 sg13g2_decap_8 FILLER_119_34 ();
 sg13g2_decap_8 FILLER_119_41 ();
 sg13g2_decap_8 FILLER_119_48 ();
 sg13g2_decap_8 FILLER_119_55 ();
 sg13g2_decap_8 FILLER_119_62 ();
 sg13g2_decap_8 FILLER_119_73 ();
 sg13g2_decap_8 FILLER_119_80 ();
 sg13g2_decap_8 FILLER_119_87 ();
 sg13g2_decap_8 FILLER_119_94 ();
 sg13g2_decap_8 FILLER_119_101 ();
 sg13g2_decap_8 FILLER_119_108 ();
 sg13g2_decap_8 FILLER_119_115 ();
 sg13g2_decap_8 FILLER_119_122 ();
 sg13g2_decap_8 FILLER_119_129 ();
 sg13g2_decap_8 FILLER_119_136 ();
 sg13g2_decap_8 FILLER_119_143 ();
 sg13g2_decap_8 FILLER_119_150 ();
 sg13g2_decap_8 FILLER_119_157 ();
 sg13g2_decap_8 FILLER_119_164 ();
 sg13g2_decap_8 FILLER_119_171 ();
 sg13g2_decap_8 FILLER_119_178 ();
 sg13g2_decap_4 FILLER_119_185 ();
 sg13g2_decap_8 FILLER_120_20 ();
 sg13g2_decap_8 FILLER_120_27 ();
 sg13g2_decap_8 FILLER_120_34 ();
 sg13g2_decap_8 FILLER_120_41 ();
 sg13g2_decap_8 FILLER_120_48 ();
 sg13g2_decap_8 FILLER_120_55 ();
 sg13g2_decap_8 FILLER_120_62 ();
 sg13g2_decap_8 FILLER_120_69 ();
 sg13g2_decap_8 FILLER_120_76 ();
 sg13g2_decap_8 FILLER_120_83 ();
 sg13g2_decap_8 FILLER_120_90 ();
 sg13g2_decap_8 FILLER_120_97 ();
 sg13g2_decap_8 FILLER_120_104 ();
 sg13g2_decap_8 FILLER_120_111 ();
 sg13g2_decap_8 FILLER_120_118 ();
 sg13g2_decap_8 FILLER_120_125 ();
 sg13g2_decap_8 FILLER_120_132 ();
 sg13g2_decap_8 FILLER_120_139 ();
 sg13g2_decap_8 FILLER_120_146 ();
 sg13g2_decap_8 FILLER_120_153 ();
 sg13g2_decap_8 FILLER_120_160 ();
 sg13g2_decap_8 FILLER_120_167 ();
 sg13g2_decap_8 FILLER_120_174 ();
 sg13g2_decap_8 FILLER_121_24 ();
 sg13g2_decap_8 FILLER_121_31 ();
 sg13g2_decap_8 FILLER_121_38 ();
 sg13g2_decap_8 FILLER_121_45 ();
 sg13g2_decap_8 FILLER_121_52 ();
 sg13g2_decap_8 FILLER_121_59 ();
 sg13g2_decap_8 FILLER_121_66 ();
 sg13g2_decap_8 FILLER_121_73 ();
 sg13g2_decap_8 FILLER_121_80 ();
 sg13g2_decap_8 FILLER_121_87 ();
 sg13g2_decap_8 FILLER_121_94 ();
 sg13g2_decap_8 FILLER_121_101 ();
 sg13g2_decap_8 FILLER_121_108 ();
 sg13g2_decap_8 FILLER_121_115 ();
 sg13g2_decap_8 FILLER_121_122 ();
 sg13g2_decap_8 FILLER_121_129 ();
 sg13g2_decap_8 FILLER_121_136 ();
 sg13g2_decap_8 FILLER_121_143 ();
 sg13g2_decap_8 FILLER_121_150 ();
 sg13g2_decap_8 FILLER_121_157 ();
 sg13g2_decap_8 FILLER_121_164 ();
 sg13g2_fill_2 FILLER_121_171 ();
 sg13g2_fill_1 FILLER_122_24 ();
 sg13g2_decap_8 FILLER_122_105 ();
 sg13g2_decap_8 FILLER_122_112 ();
 sg13g2_fill_2 FILLER_122_135 ();
 sg13g2_decap_8 FILLER_122_149 ();
 sg13g2_fill_1 FILLER_122_200 ();
 sg13g2_fill_1 FILLER_123_0 ();
 sg13g2_decap_4 FILLER_123_145 ();
 sg13g2_fill_2 FILLER_123_149 ();
 sg13g2_fill_2 FILLER_123_199 ();
 assign TIE_HIGH_SRAM = net583;
 assign TIE_LOW_SRAM = net582;
endmodule
