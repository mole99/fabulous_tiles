VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO W_IO
  CLASS BLOCK ;
  FOREIGN W_IO ;
  ORIGIN 0.000 0.000 ;
  SIZE 68.640 BY 241.920 ;
  PIN A_I_top
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 11.980 0.450 12.380 ;
    END
  END A_I_top
  PIN A_O_top
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 6.940 0.450 7.340 ;
    END
  END A_O_top
  PIN A_T_top
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 17.020 0.450 17.420 ;
    END
  END A_T_top
  PIN A_config_C_bit0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 37.180 0.450 37.580 ;
    END
  END A_config_C_bit0
  PIN A_config_C_bit1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 42.220 0.450 42.620 ;
    END
  END A_config_C_bit1
  PIN A_config_C_bit2
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 47.260 0.450 47.660 ;
    END
  END A_config_C_bit2
  PIN A_config_C_bit3
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 52.300 0.450 52.700 ;
    END
  END A_config_C_bit3
  PIN B_I_top
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 27.100 0.450 27.500 ;
    END
  END B_I_top
  PIN B_O_top
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 22.060 0.450 22.460 ;
    END
  END B_O_top
  PIN B_T_top
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 32.140 0.450 32.540 ;
    END
  END B_T_top
  PIN B_config_C_bit0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 57.340 0.450 57.740 ;
    END
  END B_config_C_bit0
  PIN B_config_C_bit1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 62.380 0.450 62.780 ;
    END
  END B_config_C_bit1
  PIN B_config_C_bit2
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 67.420 0.450 67.820 ;
    END
  END B_config_C_bit2
  PIN B_config_C_bit3
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 72.460 0.450 72.860 ;
    END
  END B_config_C_bit3
  PIN E1BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 68.190 94.300 68.640 94.700 ;
    END
  END E1BEG[0]
  PIN E1BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 68.190 95.980 68.640 96.380 ;
    END
  END E1BEG[1]
  PIN E1BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 68.190 97.660 68.640 98.060 ;
    END
  END E1BEG[2]
  PIN E1BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 68.190 99.340 68.640 99.740 ;
    END
  END E1BEG[3]
  PIN E2BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 68.190 101.020 68.640 101.420 ;
    END
  END E2BEG[0]
  PIN E2BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 68.190 102.700 68.640 103.100 ;
    END
  END E2BEG[1]
  PIN E2BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 68.190 104.380 68.640 104.780 ;
    END
  END E2BEG[2]
  PIN E2BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 68.190 106.060 68.640 106.460 ;
    END
  END E2BEG[3]
  PIN E2BEG[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 68.190 107.740 68.640 108.140 ;
    END
  END E2BEG[4]
  PIN E2BEG[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 68.190 109.420 68.640 109.820 ;
    END
  END E2BEG[5]
  PIN E2BEG[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 68.190 111.100 68.640 111.500 ;
    END
  END E2BEG[6]
  PIN E2BEG[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 68.190 112.780 68.640 113.180 ;
    END
  END E2BEG[7]
  PIN E2BEGb[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 68.190 114.460 68.640 114.860 ;
    END
  END E2BEGb[0]
  PIN E2BEGb[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 68.190 116.140 68.640 116.540 ;
    END
  END E2BEGb[1]
  PIN E2BEGb[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 68.190 117.820 68.640 118.220 ;
    END
  END E2BEGb[2]
  PIN E2BEGb[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 68.190 119.500 68.640 119.900 ;
    END
  END E2BEGb[3]
  PIN E2BEGb[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 68.190 121.180 68.640 121.580 ;
    END
  END E2BEGb[4]
  PIN E2BEGb[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 68.190 122.860 68.640 123.260 ;
    END
  END E2BEGb[5]
  PIN E2BEGb[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 68.190 124.540 68.640 124.940 ;
    END
  END E2BEGb[6]
  PIN E2BEGb[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 68.190 126.220 68.640 126.620 ;
    END
  END E2BEGb[7]
  PIN E6BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 68.190 154.780 68.640 155.180 ;
    END
  END E6BEG[0]
  PIN E6BEG[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 68.190 171.580 68.640 171.980 ;
    END
  END E6BEG[10]
  PIN E6BEG[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 68.190 173.260 68.640 173.660 ;
    END
  END E6BEG[11]
  PIN E6BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 68.190 156.460 68.640 156.860 ;
    END
  END E6BEG[1]
  PIN E6BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 68.190 158.140 68.640 158.540 ;
    END
  END E6BEG[2]
  PIN E6BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 68.190 159.820 68.640 160.220 ;
    END
  END E6BEG[3]
  PIN E6BEG[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 68.190 161.500 68.640 161.900 ;
    END
  END E6BEG[4]
  PIN E6BEG[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 68.190 163.180 68.640 163.580 ;
    END
  END E6BEG[5]
  PIN E6BEG[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 68.190 164.860 68.640 165.260 ;
    END
  END E6BEG[6]
  PIN E6BEG[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 68.190 166.540 68.640 166.940 ;
    END
  END E6BEG[7]
  PIN E6BEG[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 68.190 168.220 68.640 168.620 ;
    END
  END E6BEG[8]
  PIN E6BEG[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 68.190 169.900 68.640 170.300 ;
    END
  END E6BEG[9]
  PIN EE4BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 68.190 127.900 68.640 128.300 ;
    END
  END EE4BEG[0]
  PIN EE4BEG[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 68.190 144.700 68.640 145.100 ;
    END
  END EE4BEG[10]
  PIN EE4BEG[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 68.190 146.380 68.640 146.780 ;
    END
  END EE4BEG[11]
  PIN EE4BEG[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 68.190 148.060 68.640 148.460 ;
    END
  END EE4BEG[12]
  PIN EE4BEG[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 68.190 149.740 68.640 150.140 ;
    END
  END EE4BEG[13]
  PIN EE4BEG[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 68.190 151.420 68.640 151.820 ;
    END
  END EE4BEG[14]
  PIN EE4BEG[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 68.190 153.100 68.640 153.500 ;
    END
  END EE4BEG[15]
  PIN EE4BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 68.190 129.580 68.640 129.980 ;
    END
  END EE4BEG[1]
  PIN EE4BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 68.190 131.260 68.640 131.660 ;
    END
  END EE4BEG[2]
  PIN EE4BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 68.190 132.940 68.640 133.340 ;
    END
  END EE4BEG[3]
  PIN EE4BEG[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 68.190 134.620 68.640 135.020 ;
    END
  END EE4BEG[4]
  PIN EE4BEG[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 68.190 136.300 68.640 136.700 ;
    END
  END EE4BEG[5]
  PIN EE4BEG[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 68.190 137.980 68.640 138.380 ;
    END
  END EE4BEG[6]
  PIN EE4BEG[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 68.190 139.660 68.640 140.060 ;
    END
  END EE4BEG[7]
  PIN EE4BEG[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 68.190 141.340 68.640 141.740 ;
    END
  END EE4BEG[8]
  PIN EE4BEG[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 68.190 143.020 68.640 143.420 ;
    END
  END EE4BEG[9]
  PIN FrameData[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 77.500 0.450 77.900 ;
    END
  END FrameData[0]
  PIN FrameData[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 127.900 0.450 128.300 ;
    END
  END FrameData[10]
  PIN FrameData[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 132.940 0.450 133.340 ;
    END
  END FrameData[11]
  PIN FrameData[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 137.980 0.450 138.380 ;
    END
  END FrameData[12]
  PIN FrameData[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 143.020 0.450 143.420 ;
    END
  END FrameData[13]
  PIN FrameData[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 148.060 0.450 148.460 ;
    END
  END FrameData[14]
  PIN FrameData[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 153.100 0.450 153.500 ;
    END
  END FrameData[15]
  PIN FrameData[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 158.140 0.450 158.540 ;
    END
  END FrameData[16]
  PIN FrameData[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 163.180 0.450 163.580 ;
    END
  END FrameData[17]
  PIN FrameData[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 168.220 0.450 168.620 ;
    END
  END FrameData[18]
  PIN FrameData[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 173.260 0.450 173.660 ;
    END
  END FrameData[19]
  PIN FrameData[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 82.540 0.450 82.940 ;
    END
  END FrameData[1]
  PIN FrameData[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 178.300 0.450 178.700 ;
    END
  END FrameData[20]
  PIN FrameData[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 183.340 0.450 183.740 ;
    END
  END FrameData[21]
  PIN FrameData[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 188.380 0.450 188.780 ;
    END
  END FrameData[22]
  PIN FrameData[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 193.420 0.450 193.820 ;
    END
  END FrameData[23]
  PIN FrameData[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 198.460 0.450 198.860 ;
    END
  END FrameData[24]
  PIN FrameData[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 203.500 0.450 203.900 ;
    END
  END FrameData[25]
  PIN FrameData[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 208.540 0.450 208.940 ;
    END
  END FrameData[26]
  PIN FrameData[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 213.580 0.450 213.980 ;
    END
  END FrameData[27]
  PIN FrameData[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 218.620 0.450 219.020 ;
    END
  END FrameData[28]
  PIN FrameData[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 223.660 0.450 224.060 ;
    END
  END FrameData[29]
  PIN FrameData[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 87.580 0.450 87.980 ;
    END
  END FrameData[2]
  PIN FrameData[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 228.700 0.450 229.100 ;
    END
  END FrameData[30]
  PIN FrameData[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 233.740 0.450 234.140 ;
    END
  END FrameData[31]
  PIN FrameData[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 92.620 0.450 93.020 ;
    END
  END FrameData[3]
  PIN FrameData[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 97.660 0.450 98.060 ;
    END
  END FrameData[4]
  PIN FrameData[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 102.700 0.450 103.100 ;
    END
  END FrameData[5]
  PIN FrameData[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 107.740 0.450 108.140 ;
    END
  END FrameData[6]
  PIN FrameData[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 112.780 0.450 113.180 ;
    END
  END FrameData[7]
  PIN FrameData[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 117.820 0.450 118.220 ;
    END
  END FrameData[8]
  PIN FrameData[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 122.860 0.450 123.260 ;
    END
  END FrameData[9]
  PIN FrameData_O[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 68.190 174.940 68.640 175.340 ;
    END
  END FrameData_O[0]
  PIN FrameData_O[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 68.190 191.740 68.640 192.140 ;
    END
  END FrameData_O[10]
  PIN FrameData_O[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 68.190 193.420 68.640 193.820 ;
    END
  END FrameData_O[11]
  PIN FrameData_O[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 68.190 195.100 68.640 195.500 ;
    END
  END FrameData_O[12]
  PIN FrameData_O[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 68.190 196.780 68.640 197.180 ;
    END
  END FrameData_O[13]
  PIN FrameData_O[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 68.190 198.460 68.640 198.860 ;
    END
  END FrameData_O[14]
  PIN FrameData_O[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 68.190 200.140 68.640 200.540 ;
    END
  END FrameData_O[15]
  PIN FrameData_O[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 68.190 201.820 68.640 202.220 ;
    END
  END FrameData_O[16]
  PIN FrameData_O[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 68.190 203.500 68.640 203.900 ;
    END
  END FrameData_O[17]
  PIN FrameData_O[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 68.190 205.180 68.640 205.580 ;
    END
  END FrameData_O[18]
  PIN FrameData_O[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 68.190 206.860 68.640 207.260 ;
    END
  END FrameData_O[19]
  PIN FrameData_O[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 68.190 176.620 68.640 177.020 ;
    END
  END FrameData_O[1]
  PIN FrameData_O[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 68.190 208.540 68.640 208.940 ;
    END
  END FrameData_O[20]
  PIN FrameData_O[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 68.190 210.220 68.640 210.620 ;
    END
  END FrameData_O[21]
  PIN FrameData_O[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 68.190 211.900 68.640 212.300 ;
    END
  END FrameData_O[22]
  PIN FrameData_O[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 68.190 213.580 68.640 213.980 ;
    END
  END FrameData_O[23]
  PIN FrameData_O[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 68.190 215.260 68.640 215.660 ;
    END
  END FrameData_O[24]
  PIN FrameData_O[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 68.190 216.940 68.640 217.340 ;
    END
  END FrameData_O[25]
  PIN FrameData_O[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 68.190 218.620 68.640 219.020 ;
    END
  END FrameData_O[26]
  PIN FrameData_O[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 68.190 220.300 68.640 220.700 ;
    END
  END FrameData_O[27]
  PIN FrameData_O[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 68.190 221.980 68.640 222.380 ;
    END
  END FrameData_O[28]
  PIN FrameData_O[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 68.190 223.660 68.640 224.060 ;
    END
  END FrameData_O[29]
  PIN FrameData_O[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 68.190 178.300 68.640 178.700 ;
    END
  END FrameData_O[2]
  PIN FrameData_O[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 68.190 225.340 68.640 225.740 ;
    END
  END FrameData_O[30]
  PIN FrameData_O[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 68.190 227.020 68.640 227.420 ;
    END
  END FrameData_O[31]
  PIN FrameData_O[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 68.190 179.980 68.640 180.380 ;
    END
  END FrameData_O[3]
  PIN FrameData_O[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 68.190 181.660 68.640 182.060 ;
    END
  END FrameData_O[4]
  PIN FrameData_O[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 68.190 183.340 68.640 183.740 ;
    END
  END FrameData_O[5]
  PIN FrameData_O[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 68.190 185.020 68.640 185.420 ;
    END
  END FrameData_O[6]
  PIN FrameData_O[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 68.190 186.700 68.640 187.100 ;
    END
  END FrameData_O[7]
  PIN FrameData_O[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 68.190 188.380 68.640 188.780 ;
    END
  END FrameData_O[8]
  PIN FrameData_O[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 68.190 190.060 68.640 190.460 ;
    END
  END FrameData_O[9]
  PIN FrameStrobe[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 7.960 0.000 8.360 0.400 ;
    END
  END FrameStrobe[0]
  PIN FrameStrobe[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 36.760 0.000 37.160 0.400 ;
    END
  END FrameStrobe[10]
  PIN FrameStrobe[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 39.640 0.000 40.040 0.400 ;
    END
  END FrameStrobe[11]
  PIN FrameStrobe[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 42.520 0.000 42.920 0.400 ;
    END
  END FrameStrobe[12]
  PIN FrameStrobe[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 45.400 0.000 45.800 0.400 ;
    END
  END FrameStrobe[13]
  PIN FrameStrobe[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 48.280 0.000 48.680 0.400 ;
    END
  END FrameStrobe[14]
  PIN FrameStrobe[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 51.160 0.000 51.560 0.400 ;
    END
  END FrameStrobe[15]
  PIN FrameStrobe[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 54.040 0.000 54.440 0.400 ;
    END
  END FrameStrobe[16]
  PIN FrameStrobe[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 56.920 0.000 57.320 0.400 ;
    END
  END FrameStrobe[17]
  PIN FrameStrobe[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 59.800 0.000 60.200 0.400 ;
    END
  END FrameStrobe[18]
  PIN FrameStrobe[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 62.680 0.000 63.080 0.400 ;
    END
  END FrameStrobe[19]
  PIN FrameStrobe[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 10.840 0.000 11.240 0.400 ;
    END
  END FrameStrobe[1]
  PIN FrameStrobe[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 13.720 0.000 14.120 0.400 ;
    END
  END FrameStrobe[2]
  PIN FrameStrobe[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 16.600 0.000 17.000 0.400 ;
    END
  END FrameStrobe[3]
  PIN FrameStrobe[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 19.480 0.000 19.880 0.400 ;
    END
  END FrameStrobe[4]
  PIN FrameStrobe[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 22.360 0.000 22.760 0.400 ;
    END
  END FrameStrobe[5]
  PIN FrameStrobe[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 25.240 0.000 25.640 0.400 ;
    END
  END FrameStrobe[6]
  PIN FrameStrobe[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 28.120 0.000 28.520 0.400 ;
    END
  END FrameStrobe[7]
  PIN FrameStrobe[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 31.000 0.000 31.400 0.400 ;
    END
  END FrameStrobe[8]
  PIN FrameStrobe[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 33.880 0.000 34.280 0.400 ;
    END
  END FrameStrobe[9]
  PIN FrameStrobe_O[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 7.960 241.520 8.360 241.920 ;
    END
  END FrameStrobe_O[0]
  PIN FrameStrobe_O[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 36.760 241.520 37.160 241.920 ;
    END
  END FrameStrobe_O[10]
  PIN FrameStrobe_O[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 39.640 241.520 40.040 241.920 ;
    END
  END FrameStrobe_O[11]
  PIN FrameStrobe_O[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 42.520 241.520 42.920 241.920 ;
    END
  END FrameStrobe_O[12]
  PIN FrameStrobe_O[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 45.400 241.520 45.800 241.920 ;
    END
  END FrameStrobe_O[13]
  PIN FrameStrobe_O[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 48.280 241.520 48.680 241.920 ;
    END
  END FrameStrobe_O[14]
  PIN FrameStrobe_O[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 51.160 241.520 51.560 241.920 ;
    END
  END FrameStrobe_O[15]
  PIN FrameStrobe_O[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 54.040 241.520 54.440 241.920 ;
    END
  END FrameStrobe_O[16]
  PIN FrameStrobe_O[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 56.920 241.520 57.320 241.920 ;
    END
  END FrameStrobe_O[17]
  PIN FrameStrobe_O[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 59.800 241.520 60.200 241.920 ;
    END
  END FrameStrobe_O[18]
  PIN FrameStrobe_O[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 62.680 241.520 63.080 241.920 ;
    END
  END FrameStrobe_O[19]
  PIN FrameStrobe_O[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 10.840 241.520 11.240 241.920 ;
    END
  END FrameStrobe_O[1]
  PIN FrameStrobe_O[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 13.720 241.520 14.120 241.920 ;
    END
  END FrameStrobe_O[2]
  PIN FrameStrobe_O[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 16.600 241.520 17.000 241.920 ;
    END
  END FrameStrobe_O[3]
  PIN FrameStrobe_O[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 19.480 241.520 19.880 241.920 ;
    END
  END FrameStrobe_O[4]
  PIN FrameStrobe_O[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 22.360 241.520 22.760 241.920 ;
    END
  END FrameStrobe_O[5]
  PIN FrameStrobe_O[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 25.240 241.520 25.640 241.920 ;
    END
  END FrameStrobe_O[6]
  PIN FrameStrobe_O[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 28.120 241.520 28.520 241.920 ;
    END
  END FrameStrobe_O[7]
  PIN FrameStrobe_O[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 31.000 241.520 31.400 241.920 ;
    END
  END FrameStrobe_O[8]
  PIN FrameStrobe_O[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 33.880 241.520 34.280 241.920 ;
    END
  END FrameStrobe_O[9]
  PIN UserCLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.633100 ;
    PORT
      LAYER Metal3 ;
        RECT 5.080 0.000 5.480 0.400 ;
    END
  END UserCLK
  PIN UserCLKo
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 5.080 241.520 5.480 241.920 ;
    END
  END UserCLKo
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal5 ;
        RECT 24.460 0.000 26.660 241.920 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal5 ;
        RECT 18.260 0.000 20.460 241.920 ;
    END
  END VPWR
  PIN W1END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 68.190 13.660 68.640 14.060 ;
    END
  END W1END[0]
  PIN W1END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 68.190 15.340 68.640 15.740 ;
    END
  END W1END[1]
  PIN W1END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 68.190 17.020 68.640 17.420 ;
    END
  END W1END[2]
  PIN W1END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 68.190 18.700 68.640 19.100 ;
    END
  END W1END[3]
  PIN W2END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 68.190 33.820 68.640 34.220 ;
    END
  END W2END[0]
  PIN W2END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 68.190 35.500 68.640 35.900 ;
    END
  END W2END[1]
  PIN W2END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 68.190 37.180 68.640 37.580 ;
    END
  END W2END[2]
  PIN W2END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 68.190 38.860 68.640 39.260 ;
    END
  END W2END[3]
  PIN W2END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 68.190 40.540 68.640 40.940 ;
    END
  END W2END[4]
  PIN W2END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 68.190 42.220 68.640 42.620 ;
    END
  END W2END[5]
  PIN W2END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 68.190 43.900 68.640 44.300 ;
    END
  END W2END[6]
  PIN W2END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 68.190 45.580 68.640 45.980 ;
    END
  END W2END[7]
  PIN W2MID[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 68.190 20.380 68.640 20.780 ;
    END
  END W2MID[0]
  PIN W2MID[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 68.190 22.060 68.640 22.460 ;
    END
  END W2MID[1]
  PIN W2MID[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 68.190 23.740 68.640 24.140 ;
    END
  END W2MID[2]
  PIN W2MID[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 68.190 25.420 68.640 25.820 ;
    END
  END W2MID[3]
  PIN W2MID[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 68.190 27.100 68.640 27.500 ;
    END
  END W2MID[4]
  PIN W2MID[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 68.190 28.780 68.640 29.180 ;
    END
  END W2MID[5]
  PIN W2MID[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 68.190 30.460 68.640 30.860 ;
    END
  END W2MID[6]
  PIN W2MID[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 68.190 32.140 68.640 32.540 ;
    END
  END W2MID[7]
  PIN W6END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 68.190 74.140 68.640 74.540 ;
    END
  END W6END[0]
  PIN W6END[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 68.190 90.940 68.640 91.340 ;
    END
  END W6END[10]
  PIN W6END[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 68.190 92.620 68.640 93.020 ;
    END
  END W6END[11]
  PIN W6END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 68.190 75.820 68.640 76.220 ;
    END
  END W6END[1]
  PIN W6END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 68.190 77.500 68.640 77.900 ;
    END
  END W6END[2]
  PIN W6END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 68.190 79.180 68.640 79.580 ;
    END
  END W6END[3]
  PIN W6END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 68.190 80.860 68.640 81.260 ;
    END
  END W6END[4]
  PIN W6END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 68.190 82.540 68.640 82.940 ;
    END
  END W6END[5]
  PIN W6END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 68.190 84.220 68.640 84.620 ;
    END
  END W6END[6]
  PIN W6END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 68.190 85.900 68.640 86.300 ;
    END
  END W6END[7]
  PIN W6END[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 68.190 87.580 68.640 87.980 ;
    END
  END W6END[8]
  PIN W6END[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 68.190 89.260 68.640 89.660 ;
    END
  END W6END[9]
  PIN WW4END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 68.190 47.260 68.640 47.660 ;
    END
  END WW4END[0]
  PIN WW4END[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 68.190 64.060 68.640 64.460 ;
    END
  END WW4END[10]
  PIN WW4END[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 68.190 65.740 68.640 66.140 ;
    END
  END WW4END[11]
  PIN WW4END[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 68.190 67.420 68.640 67.820 ;
    END
  END WW4END[12]
  PIN WW4END[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 68.190 69.100 68.640 69.500 ;
    END
  END WW4END[13]
  PIN WW4END[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 68.190 70.780 68.640 71.180 ;
    END
  END WW4END[14]
  PIN WW4END[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 68.190 72.460 68.640 72.860 ;
    END
  END WW4END[15]
  PIN WW4END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 68.190 48.940 68.640 49.340 ;
    END
  END WW4END[1]
  PIN WW4END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 68.190 50.620 68.640 51.020 ;
    END
  END WW4END[2]
  PIN WW4END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 68.190 52.300 68.640 52.700 ;
    END
  END WW4END[3]
  PIN WW4END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 68.190 53.980 68.640 54.380 ;
    END
  END WW4END[4]
  PIN WW4END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 68.190 55.660 68.640 56.060 ;
    END
  END WW4END[5]
  PIN WW4END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 68.190 57.340 68.640 57.740 ;
    END
  END WW4END[6]
  PIN WW4END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 68.190 59.020 68.640 59.420 ;
    END
  END WW4END[7]
  PIN WW4END[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 68.190 60.700 68.640 61.100 ;
    END
  END WW4END[8]
  PIN WW4END[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 68.190 62.380 68.640 62.780 ;
    END
  END WW4END[9]
  OBS
      LAYER GatPoly ;
        RECT 5.760 7.410 62.880 234.510 ;
      LAYER Metal1 ;
        RECT 5.760 7.340 62.880 234.580 ;
      LAYER Metal2 ;
        RECT 0.125 234.350 68.305 234.460 ;
        RECT 0.660 233.530 68.305 234.350 ;
        RECT 0.125 229.310 68.305 233.530 ;
        RECT 0.660 228.490 68.305 229.310 ;
        RECT 0.125 227.630 68.305 228.490 ;
        RECT 0.125 226.810 67.980 227.630 ;
        RECT 0.125 225.950 68.305 226.810 ;
        RECT 0.125 225.130 67.980 225.950 ;
        RECT 0.125 224.270 68.305 225.130 ;
        RECT 0.660 223.450 67.980 224.270 ;
        RECT 0.125 222.590 68.305 223.450 ;
        RECT 0.125 221.770 67.980 222.590 ;
        RECT 0.125 220.910 68.305 221.770 ;
        RECT 0.125 220.090 67.980 220.910 ;
        RECT 0.125 219.230 68.305 220.090 ;
        RECT 0.660 218.410 67.980 219.230 ;
        RECT 0.125 217.550 68.305 218.410 ;
        RECT 0.125 216.730 67.980 217.550 ;
        RECT 0.125 215.870 68.305 216.730 ;
        RECT 0.125 215.050 67.980 215.870 ;
        RECT 0.125 214.190 68.305 215.050 ;
        RECT 0.660 213.370 67.980 214.190 ;
        RECT 0.125 212.510 68.305 213.370 ;
        RECT 0.125 211.690 67.980 212.510 ;
        RECT 0.125 210.830 68.305 211.690 ;
        RECT 0.125 210.010 67.980 210.830 ;
        RECT 0.125 209.150 68.305 210.010 ;
        RECT 0.660 208.330 67.980 209.150 ;
        RECT 0.125 207.470 68.305 208.330 ;
        RECT 0.125 206.650 67.980 207.470 ;
        RECT 0.125 205.790 68.305 206.650 ;
        RECT 0.125 204.970 67.980 205.790 ;
        RECT 0.125 204.110 68.305 204.970 ;
        RECT 0.660 203.290 67.980 204.110 ;
        RECT 0.125 202.430 68.305 203.290 ;
        RECT 0.125 201.610 67.980 202.430 ;
        RECT 0.125 200.750 68.305 201.610 ;
        RECT 0.125 199.930 67.980 200.750 ;
        RECT 0.125 199.070 68.305 199.930 ;
        RECT 0.660 198.250 67.980 199.070 ;
        RECT 0.125 197.390 68.305 198.250 ;
        RECT 0.125 196.570 67.980 197.390 ;
        RECT 0.125 195.710 68.305 196.570 ;
        RECT 0.125 194.890 67.980 195.710 ;
        RECT 0.125 194.030 68.305 194.890 ;
        RECT 0.660 193.210 67.980 194.030 ;
        RECT 0.125 192.350 68.305 193.210 ;
        RECT 0.125 191.530 67.980 192.350 ;
        RECT 0.125 190.670 68.305 191.530 ;
        RECT 0.125 189.850 67.980 190.670 ;
        RECT 0.125 188.990 68.305 189.850 ;
        RECT 0.660 188.170 67.980 188.990 ;
        RECT 0.125 187.310 68.305 188.170 ;
        RECT 0.125 186.490 67.980 187.310 ;
        RECT 0.125 185.630 68.305 186.490 ;
        RECT 0.125 184.810 67.980 185.630 ;
        RECT 0.125 183.950 68.305 184.810 ;
        RECT 0.660 183.130 67.980 183.950 ;
        RECT 0.125 182.270 68.305 183.130 ;
        RECT 0.125 181.450 67.980 182.270 ;
        RECT 0.125 180.590 68.305 181.450 ;
        RECT 0.125 179.770 67.980 180.590 ;
        RECT 0.125 178.910 68.305 179.770 ;
        RECT 0.660 178.090 67.980 178.910 ;
        RECT 0.125 177.230 68.305 178.090 ;
        RECT 0.125 176.410 67.980 177.230 ;
        RECT 0.125 175.550 68.305 176.410 ;
        RECT 0.125 174.730 67.980 175.550 ;
        RECT 0.125 173.870 68.305 174.730 ;
        RECT 0.660 173.050 67.980 173.870 ;
        RECT 0.125 172.190 68.305 173.050 ;
        RECT 0.125 171.370 67.980 172.190 ;
        RECT 0.125 170.510 68.305 171.370 ;
        RECT 0.125 169.690 67.980 170.510 ;
        RECT 0.125 168.830 68.305 169.690 ;
        RECT 0.660 168.010 67.980 168.830 ;
        RECT 0.125 167.150 68.305 168.010 ;
        RECT 0.125 166.330 67.980 167.150 ;
        RECT 0.125 165.470 68.305 166.330 ;
        RECT 0.125 164.650 67.980 165.470 ;
        RECT 0.125 163.790 68.305 164.650 ;
        RECT 0.660 162.970 67.980 163.790 ;
        RECT 0.125 162.110 68.305 162.970 ;
        RECT 0.125 161.290 67.980 162.110 ;
        RECT 0.125 160.430 68.305 161.290 ;
        RECT 0.125 159.610 67.980 160.430 ;
        RECT 0.125 158.750 68.305 159.610 ;
        RECT 0.660 157.930 67.980 158.750 ;
        RECT 0.125 157.070 68.305 157.930 ;
        RECT 0.125 156.250 67.980 157.070 ;
        RECT 0.125 155.390 68.305 156.250 ;
        RECT 0.125 154.570 67.980 155.390 ;
        RECT 0.125 153.710 68.305 154.570 ;
        RECT 0.660 152.890 67.980 153.710 ;
        RECT 0.125 152.030 68.305 152.890 ;
        RECT 0.125 151.210 67.980 152.030 ;
        RECT 0.125 150.350 68.305 151.210 ;
        RECT 0.125 149.530 67.980 150.350 ;
        RECT 0.125 148.670 68.305 149.530 ;
        RECT 0.660 147.850 67.980 148.670 ;
        RECT 0.125 146.990 68.305 147.850 ;
        RECT 0.125 146.170 67.980 146.990 ;
        RECT 0.125 145.310 68.305 146.170 ;
        RECT 0.125 144.490 67.980 145.310 ;
        RECT 0.125 143.630 68.305 144.490 ;
        RECT 0.660 142.810 67.980 143.630 ;
        RECT 0.125 141.950 68.305 142.810 ;
        RECT 0.125 141.130 67.980 141.950 ;
        RECT 0.125 140.270 68.305 141.130 ;
        RECT 0.125 139.450 67.980 140.270 ;
        RECT 0.125 138.590 68.305 139.450 ;
        RECT 0.660 137.770 67.980 138.590 ;
        RECT 0.125 136.910 68.305 137.770 ;
        RECT 0.125 136.090 67.980 136.910 ;
        RECT 0.125 135.230 68.305 136.090 ;
        RECT 0.125 134.410 67.980 135.230 ;
        RECT 0.125 133.550 68.305 134.410 ;
        RECT 0.660 132.730 67.980 133.550 ;
        RECT 0.125 131.870 68.305 132.730 ;
        RECT 0.125 131.050 67.980 131.870 ;
        RECT 0.125 130.190 68.305 131.050 ;
        RECT 0.125 129.370 67.980 130.190 ;
        RECT 0.125 128.510 68.305 129.370 ;
        RECT 0.660 127.690 67.980 128.510 ;
        RECT 0.125 126.830 68.305 127.690 ;
        RECT 0.125 126.010 67.980 126.830 ;
        RECT 0.125 125.150 68.305 126.010 ;
        RECT 0.125 124.330 67.980 125.150 ;
        RECT 0.125 123.470 68.305 124.330 ;
        RECT 0.660 122.650 67.980 123.470 ;
        RECT 0.125 121.790 68.305 122.650 ;
        RECT 0.125 120.970 67.980 121.790 ;
        RECT 0.125 120.110 68.305 120.970 ;
        RECT 0.125 119.290 67.980 120.110 ;
        RECT 0.125 118.430 68.305 119.290 ;
        RECT 0.660 117.610 67.980 118.430 ;
        RECT 0.125 116.750 68.305 117.610 ;
        RECT 0.125 115.930 67.980 116.750 ;
        RECT 0.125 115.070 68.305 115.930 ;
        RECT 0.125 114.250 67.980 115.070 ;
        RECT 0.125 113.390 68.305 114.250 ;
        RECT 0.660 112.570 67.980 113.390 ;
        RECT 0.125 111.710 68.305 112.570 ;
        RECT 0.125 110.890 67.980 111.710 ;
        RECT 0.125 110.030 68.305 110.890 ;
        RECT 0.125 109.210 67.980 110.030 ;
        RECT 0.125 108.350 68.305 109.210 ;
        RECT 0.660 107.530 67.980 108.350 ;
        RECT 0.125 106.670 68.305 107.530 ;
        RECT 0.125 105.850 67.980 106.670 ;
        RECT 0.125 104.990 68.305 105.850 ;
        RECT 0.125 104.170 67.980 104.990 ;
        RECT 0.125 103.310 68.305 104.170 ;
        RECT 0.660 102.490 67.980 103.310 ;
        RECT 0.125 101.630 68.305 102.490 ;
        RECT 0.125 100.810 67.980 101.630 ;
        RECT 0.125 99.950 68.305 100.810 ;
        RECT 0.125 99.130 67.980 99.950 ;
        RECT 0.125 98.270 68.305 99.130 ;
        RECT 0.660 97.450 67.980 98.270 ;
        RECT 0.125 96.590 68.305 97.450 ;
        RECT 0.125 95.770 67.980 96.590 ;
        RECT 0.125 94.910 68.305 95.770 ;
        RECT 0.125 94.090 67.980 94.910 ;
        RECT 0.125 93.230 68.305 94.090 ;
        RECT 0.660 92.410 67.980 93.230 ;
        RECT 0.125 91.550 68.305 92.410 ;
        RECT 0.125 90.730 67.980 91.550 ;
        RECT 0.125 89.870 68.305 90.730 ;
        RECT 0.125 89.050 67.980 89.870 ;
        RECT 0.125 88.190 68.305 89.050 ;
        RECT 0.660 87.370 67.980 88.190 ;
        RECT 0.125 86.510 68.305 87.370 ;
        RECT 0.125 85.690 67.980 86.510 ;
        RECT 0.125 84.830 68.305 85.690 ;
        RECT 0.125 84.010 67.980 84.830 ;
        RECT 0.125 83.150 68.305 84.010 ;
        RECT 0.660 82.330 67.980 83.150 ;
        RECT 0.125 81.470 68.305 82.330 ;
        RECT 0.125 80.650 67.980 81.470 ;
        RECT 0.125 79.790 68.305 80.650 ;
        RECT 0.125 78.970 67.980 79.790 ;
        RECT 0.125 78.110 68.305 78.970 ;
        RECT 0.660 77.290 67.980 78.110 ;
        RECT 0.125 76.430 68.305 77.290 ;
        RECT 0.125 75.610 67.980 76.430 ;
        RECT 0.125 74.750 68.305 75.610 ;
        RECT 0.125 73.930 67.980 74.750 ;
        RECT 0.125 73.070 68.305 73.930 ;
        RECT 0.660 72.250 67.980 73.070 ;
        RECT 0.125 71.390 68.305 72.250 ;
        RECT 0.125 70.570 67.980 71.390 ;
        RECT 0.125 69.710 68.305 70.570 ;
        RECT 0.125 68.890 67.980 69.710 ;
        RECT 0.125 68.030 68.305 68.890 ;
        RECT 0.660 67.210 67.980 68.030 ;
        RECT 0.125 66.350 68.305 67.210 ;
        RECT 0.125 65.530 67.980 66.350 ;
        RECT 0.125 64.670 68.305 65.530 ;
        RECT 0.125 63.850 67.980 64.670 ;
        RECT 0.125 62.990 68.305 63.850 ;
        RECT 0.660 62.170 67.980 62.990 ;
        RECT 0.125 61.310 68.305 62.170 ;
        RECT 0.125 60.490 67.980 61.310 ;
        RECT 0.125 59.630 68.305 60.490 ;
        RECT 0.125 58.810 67.980 59.630 ;
        RECT 0.125 57.950 68.305 58.810 ;
        RECT 0.660 57.130 67.980 57.950 ;
        RECT 0.125 56.270 68.305 57.130 ;
        RECT 0.125 55.450 67.980 56.270 ;
        RECT 0.125 54.590 68.305 55.450 ;
        RECT 0.125 53.770 67.980 54.590 ;
        RECT 0.125 52.910 68.305 53.770 ;
        RECT 0.660 52.090 67.980 52.910 ;
        RECT 0.125 51.230 68.305 52.090 ;
        RECT 0.125 50.410 67.980 51.230 ;
        RECT 0.125 49.550 68.305 50.410 ;
        RECT 0.125 48.730 67.980 49.550 ;
        RECT 0.125 47.870 68.305 48.730 ;
        RECT 0.660 47.050 67.980 47.870 ;
        RECT 0.125 46.190 68.305 47.050 ;
        RECT 0.125 45.370 67.980 46.190 ;
        RECT 0.125 44.510 68.305 45.370 ;
        RECT 0.125 43.690 67.980 44.510 ;
        RECT 0.125 42.830 68.305 43.690 ;
        RECT 0.660 42.010 67.980 42.830 ;
        RECT 0.125 41.150 68.305 42.010 ;
        RECT 0.125 40.330 67.980 41.150 ;
        RECT 0.125 39.470 68.305 40.330 ;
        RECT 0.125 38.650 67.980 39.470 ;
        RECT 0.125 37.790 68.305 38.650 ;
        RECT 0.660 36.970 67.980 37.790 ;
        RECT 0.125 36.110 68.305 36.970 ;
        RECT 0.125 35.290 67.980 36.110 ;
        RECT 0.125 34.430 68.305 35.290 ;
        RECT 0.125 33.610 67.980 34.430 ;
        RECT 0.125 32.750 68.305 33.610 ;
        RECT 0.660 31.930 67.980 32.750 ;
        RECT 0.125 31.070 68.305 31.930 ;
        RECT 0.125 30.250 67.980 31.070 ;
        RECT 0.125 29.390 68.305 30.250 ;
        RECT 0.125 28.570 67.980 29.390 ;
        RECT 0.125 27.710 68.305 28.570 ;
        RECT 0.660 26.890 67.980 27.710 ;
        RECT 0.125 26.030 68.305 26.890 ;
        RECT 0.125 25.210 67.980 26.030 ;
        RECT 0.125 24.350 68.305 25.210 ;
        RECT 0.125 23.530 67.980 24.350 ;
        RECT 0.125 22.670 68.305 23.530 ;
        RECT 0.660 21.850 67.980 22.670 ;
        RECT 0.125 20.990 68.305 21.850 ;
        RECT 0.125 20.170 67.980 20.990 ;
        RECT 0.125 19.310 68.305 20.170 ;
        RECT 0.125 18.490 67.980 19.310 ;
        RECT 0.125 17.630 68.305 18.490 ;
        RECT 0.660 16.810 67.980 17.630 ;
        RECT 0.125 15.950 68.305 16.810 ;
        RECT 0.125 15.130 67.980 15.950 ;
        RECT 0.125 14.270 68.305 15.130 ;
        RECT 0.125 13.450 67.980 14.270 ;
        RECT 0.125 12.590 68.305 13.450 ;
        RECT 0.660 11.770 68.305 12.590 ;
        RECT 0.125 7.550 68.305 11.770 ;
        RECT 0.660 7.040 68.305 7.550 ;
      LAYER Metal3 ;
        RECT 0.380 241.310 4.870 241.820 ;
        RECT 5.690 241.310 7.750 241.820 ;
        RECT 8.570 241.310 10.630 241.820 ;
        RECT 11.450 241.310 13.510 241.820 ;
        RECT 14.330 241.310 16.390 241.820 ;
        RECT 17.210 241.310 19.270 241.820 ;
        RECT 20.090 241.310 22.150 241.820 ;
        RECT 22.970 241.310 25.030 241.820 ;
        RECT 25.850 241.310 27.910 241.820 ;
        RECT 28.730 241.310 30.790 241.820 ;
        RECT 31.610 241.310 33.670 241.820 ;
        RECT 34.490 241.310 36.550 241.820 ;
        RECT 37.370 241.310 39.430 241.820 ;
        RECT 40.250 241.310 42.310 241.820 ;
        RECT 43.130 241.310 45.190 241.820 ;
        RECT 46.010 241.310 48.070 241.820 ;
        RECT 48.890 241.310 50.950 241.820 ;
        RECT 51.770 241.310 53.830 241.820 ;
        RECT 54.650 241.310 56.710 241.820 ;
        RECT 57.530 241.310 59.590 241.820 ;
        RECT 60.410 241.310 62.470 241.820 ;
        RECT 63.290 241.310 68.260 241.820 ;
        RECT 0.380 0.610 68.260 241.310 ;
        RECT 0.380 0.400 4.870 0.610 ;
        RECT 5.690 0.400 7.750 0.610 ;
        RECT 8.570 0.400 10.630 0.610 ;
        RECT 11.450 0.400 13.510 0.610 ;
        RECT 14.330 0.400 16.390 0.610 ;
        RECT 17.210 0.400 19.270 0.610 ;
        RECT 20.090 0.400 22.150 0.610 ;
        RECT 22.970 0.400 25.030 0.610 ;
        RECT 25.850 0.400 27.910 0.610 ;
        RECT 28.730 0.400 30.790 0.610 ;
        RECT 31.610 0.400 33.670 0.610 ;
        RECT 34.490 0.400 36.550 0.610 ;
        RECT 37.370 0.400 39.430 0.610 ;
        RECT 40.250 0.400 42.310 0.610 ;
        RECT 43.130 0.400 45.190 0.610 ;
        RECT 46.010 0.400 48.070 0.610 ;
        RECT 48.890 0.400 50.950 0.610 ;
        RECT 51.770 0.400 53.830 0.610 ;
        RECT 54.650 0.400 56.710 0.610 ;
        RECT 57.530 0.400 59.590 0.610 ;
        RECT 60.410 0.400 62.470 0.610 ;
        RECT 63.290 0.400 68.260 0.610 ;
      LAYER Metal4 ;
        RECT 6.625 0.320 68.305 234.460 ;
      LAYER Metal5 ;
        RECT 7.100 0.695 18.050 232.405 ;
        RECT 20.670 0.695 24.250 232.405 ;
        RECT 26.870 0.695 68.260 232.405 ;
  END
END W_IO
END LIBRARY

