magic
tech sky130A
magscale 1 2
timestamp 1740383704
<< viali >>
rect 4169 8585 4203 8619
rect 4537 8585 4571 8619
rect 4905 8585 4939 8619
rect 5365 8585 5399 8619
rect 5641 8585 5675 8619
rect 6009 8585 6043 8619
rect 6745 8585 6779 8619
rect 7113 8585 7147 8619
rect 7573 8585 7607 8619
rect 7941 8585 7975 8619
rect 8217 8585 8251 8619
rect 8585 8585 8619 8619
rect 9321 8585 9355 8619
rect 9689 8585 9723 8619
rect 10057 8585 10091 8619
rect 10425 8585 10459 8619
rect 10793 8585 10827 8619
rect 11161 8585 11195 8619
rect 11989 8585 12023 8619
rect 12357 8585 12391 8619
rect 12725 8585 12759 8619
rect 13093 8585 13127 8619
rect 13461 8585 13495 8619
rect 13829 8585 13863 8619
rect 14289 8585 14323 8619
rect 24041 8585 24075 8619
rect 24593 8585 24627 8619
rect 24961 8585 24995 8619
rect 25697 8585 25731 8619
rect 27169 8585 27203 8619
rect 28273 8585 28307 8619
rect 28641 8585 28675 8619
rect 29009 8585 29043 8619
rect 30389 8585 30423 8619
rect 31125 8585 31159 8619
rect 4353 8449 4387 8483
rect 4721 8449 4755 8483
rect 5089 8449 5123 8483
rect 5181 8449 5215 8483
rect 5825 8449 5859 8483
rect 6193 8449 6227 8483
rect 6929 8449 6963 8483
rect 7297 8449 7331 8483
rect 7389 8449 7423 8483
rect 7757 8449 7791 8483
rect 8401 8449 8435 8483
rect 8769 8449 8803 8483
rect 9505 8449 9539 8483
rect 9873 8449 9907 8483
rect 10241 8449 10275 8483
rect 10609 8449 10643 8483
rect 10977 8449 11011 8483
rect 11345 8449 11379 8483
rect 11805 8449 11839 8483
rect 12173 8449 12207 8483
rect 12541 8449 12575 8483
rect 12909 8449 12943 8483
rect 13277 8449 13311 8483
rect 13645 8449 13679 8483
rect 14105 8449 14139 8483
rect 24225 8453 24259 8487
rect 24415 8449 24449 8483
rect 24777 8449 24811 8483
rect 25145 8449 25179 8483
rect 25513 8449 25547 8483
rect 25881 8449 25915 8483
rect 26249 8449 26283 8483
rect 26985 8449 27019 8483
rect 27353 8449 27387 8483
rect 27721 8449 27755 8483
rect 28089 8449 28123 8483
rect 28457 8449 28491 8483
rect 28825 8449 28859 8483
rect 29561 8449 29595 8483
rect 29929 8449 29963 8483
rect 30573 8449 30607 8483
rect 30941 8449 30975 8483
rect 31309 8449 31343 8483
rect 31677 8449 31711 8483
rect 25329 8313 25363 8347
rect 26065 8313 26099 8347
rect 26433 8313 26467 8347
rect 27537 8313 27571 8347
rect 27905 8313 27939 8347
rect 29745 8313 29779 8347
rect 30113 8313 30147 8347
rect 31493 8313 31527 8347
rect 31861 8245 31895 8279
rect 4353 8041 4387 8075
rect 5549 8041 5583 8075
rect 6285 8041 6319 8075
rect 6837 8041 6871 8075
rect 7757 8041 7791 8075
rect 8493 8041 8527 8075
rect 9321 8041 9355 8075
rect 9873 8041 9907 8075
rect 10977 8041 11011 8075
rect 11529 8041 11563 8075
rect 12081 8041 12115 8075
rect 26157 8041 26191 8075
rect 27353 8041 27387 8075
rect 28457 8041 28491 8075
rect 28825 8041 28859 8075
rect 29745 8041 29779 8075
rect 30665 8041 30699 8075
rect 31033 8041 31067 8075
rect 31401 8041 31435 8075
rect 4537 7837 4571 7871
rect 5365 7837 5399 7871
rect 6469 7837 6503 7871
rect 7021 7837 7055 7871
rect 7573 7837 7607 7871
rect 8677 7837 8711 7871
rect 9505 7837 9539 7871
rect 10057 7837 10091 7871
rect 11161 7837 11195 7871
rect 11713 7837 11747 7871
rect 12265 7837 12299 7871
rect 26341 7837 26375 7871
rect 27169 7837 27203 7871
rect 28273 7837 28307 7871
rect 28641 7837 28675 7871
rect 29561 7837 29595 7871
rect 30481 7837 30515 7871
rect 30849 7837 30883 7871
rect 31217 7837 31251 7871
rect 31585 7837 31619 7871
rect 31953 7837 31987 7871
rect 31769 7701 31803 7735
rect 32137 7701 32171 7735
rect 23121 7497 23155 7531
rect 24501 7497 24535 7531
rect 31493 7497 31527 7531
rect 26249 7429 26283 7463
rect 27445 7429 27479 7463
rect 22017 7361 22051 7395
rect 23213 7361 23247 7395
rect 23305 7361 23339 7395
rect 24593 7361 24627 7395
rect 24685 7361 24719 7395
rect 26341 7361 26375 7395
rect 27537 7361 27571 7395
rect 27629 7361 27663 7395
rect 31309 7361 31343 7395
rect 31677 7361 31711 7395
rect 23489 7225 23523 7259
rect 26525 7225 26559 7259
rect 22201 7157 22235 7191
rect 24869 7157 24903 7191
rect 27813 7157 27847 7191
rect 31861 7157 31895 7191
rect 4445 6953 4479 6987
rect 6285 6953 6319 6987
rect 12633 6953 12667 6987
rect 14381 6953 14415 6987
rect 16589 6953 16623 6987
rect 16865 6953 16899 6987
rect 19809 6953 19843 6987
rect 20729 6953 20763 6987
rect 26617 6953 26651 6987
rect 21373 6885 21407 6919
rect 24593 6885 24627 6919
rect 4261 6749 4295 6783
rect 6469 6749 6503 6783
rect 8033 6749 8067 6783
rect 10149 6749 10183 6783
rect 10241 6749 10275 6783
rect 10609 6749 10643 6783
rect 10701 6749 10735 6783
rect 11069 6749 11103 6783
rect 11345 6749 11379 6783
rect 11621 6749 11655 6783
rect 12817 6749 12851 6783
rect 13645 6749 13679 6783
rect 14565 6749 14599 6783
rect 15761 6749 15795 6783
rect 16221 6749 16255 6783
rect 16405 6749 16439 6783
rect 16681 6749 16715 6783
rect 16957 6749 16991 6783
rect 17325 6749 17359 6783
rect 17693 6749 17727 6783
rect 18429 6749 18463 6783
rect 19349 6749 19383 6783
rect 19625 6749 19659 6783
rect 19993 6749 20027 6783
rect 20913 6749 20947 6783
rect 21005 6749 21039 6783
rect 21189 6749 21223 6783
rect 21465 6749 21499 6783
rect 21741 6749 21775 6783
rect 23397 6749 23431 6783
rect 23673 6749 23707 6783
rect 24409 6749 24443 6783
rect 26065 6749 26099 6783
rect 26157 6749 26191 6783
rect 26433 6749 26467 6783
rect 31217 6749 31251 6783
rect 31585 6749 31619 6783
rect 31953 6749 31987 6783
rect 25973 6681 26007 6715
rect 7849 6613 7883 6647
rect 9965 6613 9999 6647
rect 10425 6613 10459 6647
rect 10885 6613 10919 6647
rect 11253 6613 11287 6647
rect 11529 6613 11563 6647
rect 11805 6613 11839 6647
rect 13461 6613 13495 6647
rect 15577 6613 15611 6647
rect 17141 6613 17175 6647
rect 17509 6613 17543 6647
rect 18245 6613 18279 6647
rect 19533 6613 19567 6647
rect 21649 6613 21683 6647
rect 23581 6613 23615 6647
rect 23857 6613 23891 6647
rect 26341 6613 26375 6647
rect 31401 6613 31435 6647
rect 31769 6613 31803 6647
rect 32137 6613 32171 6647
rect 5273 6409 5307 6443
rect 6653 6409 6687 6443
rect 7665 6409 7699 6443
rect 8401 6409 8435 6443
rect 8677 6409 8711 6443
rect 9229 6409 9263 6443
rect 10057 6409 10091 6443
rect 10333 6409 10367 6443
rect 28733 6409 28767 6443
rect 30849 6409 30883 6443
rect 31861 6409 31895 6443
rect 5457 6273 5491 6307
rect 6837 6273 6871 6307
rect 7849 6273 7883 6307
rect 8125 6273 8159 6307
rect 8217 6273 8251 6307
rect 8585 6273 8619 6307
rect 8861 6273 8895 6307
rect 9137 6273 9171 6307
rect 9413 6273 9447 6307
rect 9689 6273 9723 6307
rect 9781 6273 9815 6307
rect 10249 6277 10283 6311
rect 10517 6277 10551 6311
rect 10885 6273 10919 6307
rect 11253 6273 11287 6307
rect 22109 6273 22143 6307
rect 28549 6273 28583 6307
rect 31033 6273 31067 6307
rect 31309 6273 31343 6307
rect 31677 6273 31711 6307
rect 7941 6137 7975 6171
rect 9505 6137 9539 6171
rect 10701 6137 10735 6171
rect 31493 6137 31527 6171
rect 9965 6069 9999 6103
rect 11069 6069 11103 6103
rect 22293 6069 22327 6103
rect 6745 5865 6779 5899
rect 7389 5865 7423 5899
rect 7665 5865 7699 5899
rect 21649 5797 21683 5831
rect 31401 5797 31435 5831
rect 32137 5797 32171 5831
rect 6561 5661 6595 5695
rect 7205 5661 7239 5695
rect 7849 5661 7883 5695
rect 9137 5661 9171 5695
rect 16221 5661 16255 5695
rect 16405 5661 16439 5695
rect 21465 5661 21499 5695
rect 31217 5661 31251 5695
rect 31585 5661 31619 5695
rect 31953 5661 31987 5695
rect 8953 5525 8987 5559
rect 16589 5525 16623 5559
rect 31769 5525 31803 5559
rect 8493 5321 8527 5355
rect 21465 5321 21499 5355
rect 8677 5185 8711 5219
rect 15117 5185 15151 5219
rect 21281 5185 21315 5219
rect 31309 5185 31343 5219
rect 31677 5185 31711 5219
rect 15301 5049 15335 5083
rect 31493 4981 31527 5015
rect 31861 4981 31895 5015
rect 19533 4573 19567 4607
rect 22661 4573 22695 4607
rect 23765 4573 23799 4607
rect 31585 4573 31619 4607
rect 31953 4573 31987 4607
rect 19717 4437 19751 4471
rect 22845 4437 22879 4471
rect 23949 4437 23983 4471
rect 31769 4437 31803 4471
rect 32137 4437 32171 4471
rect 12449 4097 12483 4131
rect 12541 4097 12575 4131
rect 20913 4097 20947 4131
rect 31309 4097 31343 4131
rect 31677 4097 31711 4131
rect 12725 3893 12759 3927
rect 21097 3893 21131 3927
rect 31493 3893 31527 3927
rect 31861 3893 31895 3927
rect 6929 3689 6963 3723
rect 11805 3689 11839 3723
rect 15301 3689 15335 3723
rect 15669 3689 15703 3723
rect 15945 3689 15979 3723
rect 17601 3689 17635 3723
rect 17969 3689 18003 3723
rect 18153 3689 18187 3723
rect 19073 3689 19107 3723
rect 19441 3689 19475 3723
rect 19901 3689 19935 3723
rect 22017 3689 22051 3723
rect 25513 3689 25547 3723
rect 26157 3689 26191 3723
rect 10241 3621 10275 3655
rect 10885 3621 10919 3655
rect 15025 3621 15059 3655
rect 16773 3621 16807 3655
rect 19717 3621 19751 3655
rect 11161 3553 11195 3587
rect 17693 3553 17727 3587
rect 4721 3485 4755 3519
rect 6745 3485 6779 3519
rect 8217 3485 8251 3519
rect 9413 3485 9447 3519
rect 10333 3485 10367 3519
rect 10425 3485 10459 3519
rect 10701 3485 10735 3519
rect 11253 3485 11287 3519
rect 11345 3485 11379 3519
rect 11897 3485 11931 3519
rect 11989 3485 12023 3519
rect 12265 3485 12299 3519
rect 12541 3485 12575 3519
rect 14565 3485 14599 3519
rect 15393 3485 15427 3519
rect 15485 3485 15519 3519
rect 15761 3485 15795 3519
rect 16957 3485 16991 3519
rect 17049 3485 17083 3519
rect 17325 3485 17359 3519
rect 17785 3485 17819 3519
rect 18337 3485 18371 3519
rect 18613 3485 18647 3519
rect 18889 3485 18923 3519
rect 19257 3485 19291 3519
rect 19533 3485 19567 3519
rect 20177 3485 20211 3519
rect 21833 3485 21867 3519
rect 22201 3485 22235 3519
rect 22477 3485 22511 3519
rect 25329 3485 25363 3519
rect 25605 3485 25639 3519
rect 25973 3485 26007 3519
rect 31585 3485 31619 3519
rect 31953 3485 31987 3519
rect 4905 3349 4939 3383
rect 8401 3349 8435 3383
rect 9597 3349 9631 3383
rect 10609 3349 10643 3383
rect 11529 3349 11563 3383
rect 12173 3349 12207 3383
rect 12449 3349 12483 3383
rect 14749 3349 14783 3383
rect 16589 3349 16623 3383
rect 16681 3349 16715 3383
rect 16865 3349 16899 3383
rect 17233 3349 17267 3383
rect 17509 3349 17543 3383
rect 18521 3349 18555 3383
rect 18797 3349 18831 3383
rect 19993 3349 20027 3383
rect 22385 3349 22419 3383
rect 22661 3349 22695 3383
rect 25789 3349 25823 3383
rect 31769 3349 31803 3383
rect 32137 3349 32171 3383
rect 31309 3009 31343 3043
rect 31677 3009 31711 3043
rect 31493 2805 31527 2839
rect 31861 2805 31895 2839
rect 30573 2397 30607 2431
rect 30941 2397 30975 2431
rect 31309 2397 31343 2431
rect 31677 2397 31711 2431
rect 30757 2261 30791 2295
rect 31125 2261 31159 2295
rect 31493 2261 31527 2295
rect 31861 2261 31895 2295
<< metal1 >>
rect 15654 11092 15660 11144
rect 15712 11132 15718 11144
rect 22094 11132 22100 11144
rect 15712 11104 22100 11132
rect 15712 11092 15718 11104
rect 22094 11092 22100 11104
rect 22152 11092 22158 11144
rect 13630 10004 13636 10056
rect 13688 10044 13694 10056
rect 19334 10044 19340 10056
rect 13688 10016 19340 10044
rect 13688 10004 13694 10016
rect 19334 10004 19340 10016
rect 19392 10004 19398 10056
rect 25682 9596 25688 9648
rect 25740 9636 25746 9648
rect 26142 9636 26148 9648
rect 25740 9608 26148 9636
rect 25740 9596 25746 9608
rect 26142 9596 26148 9608
rect 26200 9596 26206 9648
rect 7650 9392 7656 9444
rect 7708 9432 7714 9444
rect 18782 9432 18788 9444
rect 7708 9404 18788 9432
rect 7708 9392 7714 9404
rect 18782 9392 18788 9404
rect 18840 9392 18846 9444
rect 8386 9256 8392 9308
rect 8444 9296 8450 9308
rect 12526 9296 12532 9308
rect 8444 9268 12532 9296
rect 8444 9256 8450 9268
rect 12526 9256 12532 9268
rect 12584 9256 12590 9308
rect 12802 9256 12808 9308
rect 12860 9296 12866 9308
rect 20990 9296 20996 9308
rect 12860 9268 20996 9296
rect 12860 9256 12866 9268
rect 20990 9256 20996 9268
rect 21048 9256 21054 9308
rect 10318 9188 10324 9240
rect 10376 9228 10382 9240
rect 17954 9228 17960 9240
rect 10376 9200 17960 9228
rect 10376 9188 10382 9200
rect 17954 9188 17960 9200
rect 18012 9188 18018 9240
rect 9858 9120 9864 9172
rect 9916 9160 9922 9172
rect 19242 9160 19248 9172
rect 9916 9132 19248 9160
rect 9916 9120 9922 9132
rect 19242 9120 19248 9132
rect 19300 9120 19306 9172
rect 10410 9052 10416 9104
rect 10468 9092 10474 9104
rect 18230 9092 18236 9104
rect 10468 9064 18236 9092
rect 10468 9052 10474 9064
rect 18230 9052 18236 9064
rect 18288 9052 18294 9104
rect 23474 9052 23480 9104
rect 23532 9092 23538 9104
rect 23750 9092 23756 9104
rect 23532 9064 23756 9092
rect 23532 9052 23538 9064
rect 23750 9052 23756 9064
rect 23808 9052 23814 9104
rect 27614 9052 27620 9104
rect 27672 9092 27678 9104
rect 28626 9092 28632 9104
rect 27672 9064 28632 9092
rect 27672 9052 27678 9064
rect 28626 9052 28632 9064
rect 28684 9052 28690 9104
rect 10594 8984 10600 9036
rect 10652 9024 10658 9036
rect 14090 9024 14096 9036
rect 10652 8996 14096 9024
rect 10652 8984 10658 8996
rect 14090 8984 14096 8996
rect 14148 8984 14154 9036
rect 21726 8984 21732 9036
rect 21784 9024 21790 9036
rect 28074 9024 28080 9036
rect 21784 8996 28080 9024
rect 21784 8984 21790 8996
rect 28074 8984 28080 8996
rect 28132 8984 28138 9036
rect 13722 8916 13728 8968
rect 13780 8956 13786 8968
rect 26878 8956 26884 8968
rect 13780 8928 26884 8956
rect 13780 8916 13786 8928
rect 26878 8916 26884 8928
rect 26936 8916 26942 8968
rect 27522 8916 27528 8968
rect 27580 8956 27586 8968
rect 31662 8956 31668 8968
rect 27580 8928 31668 8956
rect 27580 8916 27586 8928
rect 31662 8916 31668 8928
rect 31720 8916 31726 8968
rect 10962 8848 10968 8900
rect 11020 8888 11026 8900
rect 15562 8888 15568 8900
rect 11020 8860 15568 8888
rect 11020 8848 11026 8860
rect 15562 8848 15568 8860
rect 15620 8848 15626 8900
rect 17954 8848 17960 8900
rect 18012 8888 18018 8900
rect 25038 8888 25044 8900
rect 18012 8860 25044 8888
rect 18012 8848 18018 8860
rect 25038 8848 25044 8860
rect 25096 8848 25102 8900
rect 26694 8848 26700 8900
rect 26752 8888 26758 8900
rect 29914 8888 29920 8900
rect 26752 8860 29920 8888
rect 26752 8848 26758 8860
rect 29914 8848 29920 8860
rect 29972 8848 29978 8900
rect 11422 8780 11428 8832
rect 11480 8820 11486 8832
rect 13446 8820 13452 8832
rect 11480 8792 13452 8820
rect 11480 8780 11486 8792
rect 13446 8780 13452 8792
rect 13504 8780 13510 8832
rect 21266 8780 21272 8832
rect 21324 8820 21330 8832
rect 21542 8820 21548 8832
rect 21324 8792 21548 8820
rect 21324 8780 21330 8792
rect 21542 8780 21548 8792
rect 21600 8780 21606 8832
rect 23658 8780 23664 8832
rect 23716 8820 23722 8832
rect 28810 8820 28816 8832
rect 23716 8792 28816 8820
rect 23716 8780 23722 8792
rect 28810 8780 28816 8792
rect 28868 8780 28874 8832
rect 1104 8730 32568 8752
rect 1104 8678 3010 8730
rect 3062 8678 3074 8730
rect 3126 8678 3138 8730
rect 3190 8678 3202 8730
rect 3254 8678 3266 8730
rect 3318 8678 9010 8730
rect 9062 8678 9074 8730
rect 9126 8678 9138 8730
rect 9190 8678 9202 8730
rect 9254 8678 9266 8730
rect 9318 8678 15010 8730
rect 15062 8678 15074 8730
rect 15126 8678 15138 8730
rect 15190 8678 15202 8730
rect 15254 8678 15266 8730
rect 15318 8678 21010 8730
rect 21062 8678 21074 8730
rect 21126 8678 21138 8730
rect 21190 8678 21202 8730
rect 21254 8678 21266 8730
rect 21318 8678 27010 8730
rect 27062 8678 27074 8730
rect 27126 8678 27138 8730
rect 27190 8678 27202 8730
rect 27254 8678 27266 8730
rect 27318 8678 32568 8730
rect 1104 8656 32568 8678
rect 4157 8619 4215 8625
rect 4157 8585 4169 8619
rect 4203 8616 4215 8619
rect 4430 8616 4436 8628
rect 4203 8588 4436 8616
rect 4203 8585 4215 8588
rect 4157 8579 4215 8585
rect 4430 8576 4436 8588
rect 4488 8576 4494 8628
rect 4525 8619 4583 8625
rect 4525 8585 4537 8619
rect 4571 8616 4583 8619
rect 4706 8616 4712 8628
rect 4571 8588 4712 8616
rect 4571 8585 4583 8588
rect 4525 8579 4583 8585
rect 4706 8576 4712 8588
rect 4764 8576 4770 8628
rect 4893 8619 4951 8625
rect 4893 8585 4905 8619
rect 4939 8616 4951 8619
rect 4982 8616 4988 8628
rect 4939 8588 4988 8616
rect 4939 8585 4951 8588
rect 4893 8579 4951 8585
rect 4982 8576 4988 8588
rect 5040 8576 5046 8628
rect 5353 8619 5411 8625
rect 5353 8585 5365 8619
rect 5399 8616 5411 8619
rect 5534 8616 5540 8628
rect 5399 8588 5540 8616
rect 5399 8585 5411 8588
rect 5353 8579 5411 8585
rect 5534 8576 5540 8588
rect 5592 8576 5598 8628
rect 5629 8619 5687 8625
rect 5629 8585 5641 8619
rect 5675 8616 5687 8619
rect 5810 8616 5816 8628
rect 5675 8588 5816 8616
rect 5675 8585 5687 8588
rect 5629 8579 5687 8585
rect 5810 8576 5816 8588
rect 5868 8576 5874 8628
rect 5997 8619 6055 8625
rect 5997 8585 6009 8619
rect 6043 8616 6055 8619
rect 6362 8616 6368 8628
rect 6043 8588 6368 8616
rect 6043 8585 6055 8588
rect 5997 8579 6055 8585
rect 6362 8576 6368 8588
rect 6420 8576 6426 8628
rect 6733 8619 6791 8625
rect 6733 8585 6745 8619
rect 6779 8616 6791 8619
rect 6914 8616 6920 8628
rect 6779 8588 6920 8616
rect 6779 8585 6791 8588
rect 6733 8579 6791 8585
rect 6914 8576 6920 8588
rect 6972 8576 6978 8628
rect 7101 8619 7159 8625
rect 7101 8585 7113 8619
rect 7147 8616 7159 8619
rect 7190 8616 7196 8628
rect 7147 8588 7196 8616
rect 7147 8585 7159 8588
rect 7101 8579 7159 8585
rect 7190 8576 7196 8588
rect 7248 8576 7254 8628
rect 7561 8619 7619 8625
rect 7561 8585 7573 8619
rect 7607 8616 7619 8619
rect 7742 8616 7748 8628
rect 7607 8588 7748 8616
rect 7607 8585 7619 8588
rect 7561 8579 7619 8585
rect 7742 8576 7748 8588
rect 7800 8576 7806 8628
rect 7929 8619 7987 8625
rect 7929 8585 7941 8619
rect 7975 8616 7987 8619
rect 8018 8616 8024 8628
rect 7975 8588 8024 8616
rect 7975 8585 7987 8588
rect 7929 8579 7987 8585
rect 8018 8576 8024 8588
rect 8076 8576 8082 8628
rect 8205 8619 8263 8625
rect 8205 8585 8217 8619
rect 8251 8616 8263 8619
rect 8478 8616 8484 8628
rect 8251 8588 8484 8616
rect 8251 8585 8263 8588
rect 8205 8579 8263 8585
rect 8478 8576 8484 8588
rect 8536 8576 8542 8628
rect 8573 8619 8631 8625
rect 8573 8585 8585 8619
rect 8619 8616 8631 8619
rect 8754 8616 8760 8628
rect 8619 8588 8760 8616
rect 8619 8585 8631 8588
rect 8573 8579 8631 8585
rect 8754 8576 8760 8588
rect 8812 8576 8818 8628
rect 9309 8619 9367 8625
rect 9309 8585 9321 8619
rect 9355 8616 9367 8619
rect 9398 8616 9404 8628
rect 9355 8588 9404 8616
rect 9355 8585 9367 8588
rect 9309 8579 9367 8585
rect 9398 8576 9404 8588
rect 9456 8576 9462 8628
rect 9677 8619 9735 8625
rect 9677 8585 9689 8619
rect 9723 8616 9735 8619
rect 9950 8616 9956 8628
rect 9723 8588 9956 8616
rect 9723 8585 9735 8588
rect 9677 8579 9735 8585
rect 9950 8576 9956 8588
rect 10008 8576 10014 8628
rect 10045 8619 10103 8625
rect 10045 8585 10057 8619
rect 10091 8616 10103 8619
rect 10226 8616 10232 8628
rect 10091 8588 10232 8616
rect 10091 8585 10103 8588
rect 10045 8579 10103 8585
rect 10226 8576 10232 8588
rect 10284 8576 10290 8628
rect 10413 8619 10471 8625
rect 10413 8585 10425 8619
rect 10459 8616 10471 8619
rect 10502 8616 10508 8628
rect 10459 8588 10508 8616
rect 10459 8585 10471 8588
rect 10413 8579 10471 8585
rect 10502 8576 10508 8588
rect 10560 8576 10566 8628
rect 10781 8619 10839 8625
rect 10781 8585 10793 8619
rect 10827 8616 10839 8619
rect 11054 8616 11060 8628
rect 10827 8588 11060 8616
rect 10827 8585 10839 8588
rect 10781 8579 10839 8585
rect 11054 8576 11060 8588
rect 11112 8576 11118 8628
rect 11149 8619 11207 8625
rect 11149 8585 11161 8619
rect 11195 8616 11207 8619
rect 11606 8616 11612 8628
rect 11195 8588 11612 8616
rect 11195 8585 11207 8588
rect 11149 8579 11207 8585
rect 11606 8576 11612 8588
rect 11664 8576 11670 8628
rect 11977 8619 12035 8625
rect 11977 8585 11989 8619
rect 12023 8616 12035 8619
rect 12158 8616 12164 8628
rect 12023 8588 12164 8616
rect 12023 8585 12035 8588
rect 11977 8579 12035 8585
rect 12158 8576 12164 8588
rect 12216 8576 12222 8628
rect 12345 8619 12403 8625
rect 12345 8585 12357 8619
rect 12391 8616 12403 8619
rect 12434 8616 12440 8628
rect 12391 8588 12440 8616
rect 12391 8585 12403 8588
rect 12345 8579 12403 8585
rect 12434 8576 12440 8588
rect 12492 8576 12498 8628
rect 12710 8576 12716 8628
rect 12768 8576 12774 8628
rect 12986 8576 12992 8628
rect 13044 8616 13050 8628
rect 13081 8619 13139 8625
rect 13081 8616 13093 8619
rect 13044 8588 13093 8616
rect 13044 8576 13050 8588
rect 13081 8585 13093 8588
rect 13127 8585 13139 8619
rect 13081 8579 13139 8585
rect 13262 8576 13268 8628
rect 13320 8616 13326 8628
rect 13449 8619 13507 8625
rect 13449 8616 13461 8619
rect 13320 8588 13461 8616
rect 13320 8576 13326 8588
rect 13449 8585 13461 8588
rect 13495 8585 13507 8619
rect 13449 8579 13507 8585
rect 13538 8576 13544 8628
rect 13596 8616 13602 8628
rect 13817 8619 13875 8625
rect 13817 8616 13829 8619
rect 13596 8588 13829 8616
rect 13596 8576 13602 8588
rect 13817 8585 13829 8588
rect 13863 8585 13875 8619
rect 13817 8579 13875 8585
rect 13906 8576 13912 8628
rect 13964 8616 13970 8628
rect 14277 8619 14335 8625
rect 14277 8616 14289 8619
rect 13964 8588 14289 8616
rect 13964 8576 13970 8588
rect 14277 8585 14289 8588
rect 14323 8585 14335 8619
rect 14277 8579 14335 8585
rect 24026 8576 24032 8628
rect 24084 8576 24090 8628
rect 24136 8588 24348 8616
rect 10686 8548 10692 8560
rect 9508 8520 10692 8548
rect 4338 8440 4344 8492
rect 4396 8440 4402 8492
rect 4706 8440 4712 8492
rect 4764 8440 4770 8492
rect 5077 8483 5135 8489
rect 5077 8449 5089 8483
rect 5123 8449 5135 8483
rect 5077 8443 5135 8449
rect 5092 8412 5120 8443
rect 5166 8440 5172 8492
rect 5224 8440 5230 8492
rect 5810 8440 5816 8492
rect 5868 8440 5874 8492
rect 6178 8440 6184 8492
rect 6236 8440 6242 8492
rect 6917 8483 6975 8489
rect 6917 8449 6929 8483
rect 6963 8480 6975 8483
rect 7098 8480 7104 8492
rect 6963 8452 7104 8480
rect 6963 8449 6975 8452
rect 6917 8443 6975 8449
rect 7098 8440 7104 8452
rect 7156 8440 7162 8492
rect 7282 8440 7288 8492
rect 7340 8440 7346 8492
rect 7374 8440 7380 8492
rect 7432 8440 7438 8492
rect 7742 8440 7748 8492
rect 7800 8440 7806 8492
rect 8389 8483 8447 8489
rect 8389 8449 8401 8483
rect 8435 8480 8447 8483
rect 8662 8480 8668 8492
rect 8435 8452 8668 8480
rect 8435 8449 8447 8452
rect 8389 8443 8447 8449
rect 8662 8440 8668 8452
rect 8720 8440 8726 8492
rect 9508 8489 9536 8520
rect 10686 8508 10692 8520
rect 10744 8508 10750 8560
rect 11238 8508 11244 8560
rect 11296 8548 11302 8560
rect 11296 8520 13308 8548
rect 11296 8508 11302 8520
rect 8757 8483 8815 8489
rect 8757 8449 8769 8483
rect 8803 8449 8815 8483
rect 8757 8443 8815 8449
rect 9493 8483 9551 8489
rect 9493 8449 9505 8483
rect 9539 8449 9551 8483
rect 9493 8443 9551 8449
rect 8570 8412 8576 8424
rect 5092 8384 8576 8412
rect 8570 8372 8576 8384
rect 8628 8372 8634 8424
rect 8772 8344 8800 8443
rect 9858 8440 9864 8492
rect 9916 8440 9922 8492
rect 10229 8483 10287 8489
rect 10229 8449 10241 8483
rect 10275 8480 10287 8483
rect 10410 8480 10416 8492
rect 10275 8452 10416 8480
rect 10275 8449 10287 8452
rect 10229 8443 10287 8449
rect 10410 8440 10416 8452
rect 10468 8440 10474 8492
rect 10597 8483 10655 8489
rect 10597 8449 10609 8483
rect 10643 8449 10655 8483
rect 10597 8443 10655 8449
rect 10226 8344 10232 8356
rect 8772 8316 10232 8344
rect 10226 8304 10232 8316
rect 10284 8304 10290 8356
rect 10612 8344 10640 8443
rect 10962 8440 10968 8492
rect 11020 8440 11026 8492
rect 11333 8483 11391 8489
rect 11333 8449 11345 8483
rect 11379 8480 11391 8483
rect 11422 8480 11428 8492
rect 11379 8452 11428 8480
rect 11379 8449 11391 8452
rect 11333 8443 11391 8449
rect 11422 8440 11428 8452
rect 11480 8440 11486 8492
rect 11514 8440 11520 8492
rect 11572 8480 11578 8492
rect 11793 8483 11851 8489
rect 11793 8480 11805 8483
rect 11572 8452 11805 8480
rect 11572 8440 11578 8452
rect 11793 8449 11805 8452
rect 11839 8449 11851 8483
rect 11793 8443 11851 8449
rect 12158 8440 12164 8492
rect 12216 8440 12222 8492
rect 12526 8440 12532 8492
rect 12584 8440 12590 8492
rect 13280 8489 13308 8520
rect 16942 8508 16948 8560
rect 17000 8548 17006 8560
rect 24136 8548 24164 8588
rect 17000 8520 24164 8548
rect 24320 8548 24348 8588
rect 24394 8576 24400 8628
rect 24452 8616 24458 8628
rect 24581 8619 24639 8625
rect 24581 8616 24593 8619
rect 24452 8588 24593 8616
rect 24452 8576 24458 8588
rect 24581 8585 24593 8588
rect 24627 8585 24639 8619
rect 24581 8579 24639 8585
rect 24670 8576 24676 8628
rect 24728 8616 24734 8628
rect 24949 8619 25007 8625
rect 24949 8616 24961 8619
rect 24728 8588 24961 8616
rect 24728 8576 24734 8588
rect 24949 8585 24961 8588
rect 24995 8585 25007 8619
rect 24949 8579 25007 8585
rect 25038 8576 25044 8628
rect 25096 8576 25102 8628
rect 25130 8576 25136 8628
rect 25188 8616 25194 8628
rect 25685 8619 25743 8625
rect 25685 8616 25697 8619
rect 25188 8588 25697 8616
rect 25188 8576 25194 8588
rect 25685 8585 25697 8588
rect 25731 8585 25743 8619
rect 25685 8579 25743 8585
rect 26234 8576 26240 8628
rect 26292 8616 26298 8628
rect 27157 8619 27215 8625
rect 27157 8616 27169 8619
rect 26292 8588 27169 8616
rect 26292 8576 26298 8588
rect 27157 8585 27169 8588
rect 27203 8585 27215 8619
rect 27157 8579 27215 8585
rect 27430 8576 27436 8628
rect 27488 8616 27494 8628
rect 28261 8619 28319 8625
rect 28261 8616 28273 8619
rect 27488 8588 28273 8616
rect 27488 8576 27494 8588
rect 28261 8585 28273 8588
rect 28307 8585 28319 8619
rect 28261 8579 28319 8585
rect 28626 8576 28632 8628
rect 28684 8576 28690 8628
rect 28997 8619 29055 8625
rect 28997 8585 29009 8619
rect 29043 8585 29055 8619
rect 28997 8579 29055 8585
rect 24320 8520 24808 8548
rect 17000 8508 17006 8520
rect 12897 8483 12955 8489
rect 12897 8449 12909 8483
rect 12943 8449 12955 8483
rect 12897 8443 12955 8449
rect 13265 8483 13323 8489
rect 13265 8449 13277 8483
rect 13311 8449 13323 8483
rect 13265 8443 13323 8449
rect 11974 8372 11980 8424
rect 12032 8412 12038 8424
rect 12912 8412 12940 8443
rect 13354 8440 13360 8492
rect 13412 8480 13418 8492
rect 13633 8483 13691 8489
rect 13633 8480 13645 8483
rect 13412 8452 13645 8480
rect 13412 8440 13418 8452
rect 13633 8449 13645 8452
rect 13679 8449 13691 8483
rect 13633 8443 13691 8449
rect 14090 8440 14096 8492
rect 14148 8440 14154 8492
rect 24210 8444 24216 8496
rect 24268 8444 24274 8496
rect 24780 8489 24808 8520
rect 24403 8483 24461 8489
rect 24403 8449 24415 8483
rect 24449 8449 24461 8483
rect 24403 8443 24461 8449
rect 24765 8483 24823 8489
rect 24765 8449 24777 8483
rect 24811 8449 24823 8483
rect 25056 8480 25084 8576
rect 25222 8508 25228 8560
rect 25280 8548 25286 8560
rect 25280 8520 26188 8548
rect 25280 8508 25286 8520
rect 25133 8483 25191 8489
rect 25133 8480 25145 8483
rect 25056 8452 25145 8480
rect 24765 8443 24823 8449
rect 25133 8449 25145 8452
rect 25179 8449 25191 8483
rect 25133 8443 25191 8449
rect 12032 8384 12940 8412
rect 12032 8372 12038 8384
rect 13538 8372 13544 8424
rect 13596 8412 13602 8424
rect 16574 8412 16580 8424
rect 13596 8384 16580 8412
rect 13596 8372 13602 8384
rect 16574 8372 16580 8384
rect 16632 8372 16638 8424
rect 22370 8372 22376 8424
rect 22428 8412 22434 8424
rect 24412 8412 24440 8443
rect 25498 8440 25504 8492
rect 25556 8440 25562 8492
rect 25869 8483 25927 8489
rect 25869 8480 25881 8483
rect 25608 8452 25881 8480
rect 25608 8412 25636 8452
rect 25869 8449 25881 8452
rect 25915 8449 25927 8483
rect 25869 8443 25927 8449
rect 22428 8384 24440 8412
rect 24964 8384 25636 8412
rect 26160 8412 26188 8520
rect 26786 8508 26792 8560
rect 26844 8548 26850 8560
rect 26844 8520 27844 8548
rect 26844 8508 26850 8520
rect 26237 8483 26295 8489
rect 26237 8449 26249 8483
rect 26283 8480 26295 8483
rect 26326 8480 26332 8492
rect 26283 8452 26332 8480
rect 26283 8449 26295 8452
rect 26237 8443 26295 8449
rect 26326 8440 26332 8452
rect 26384 8440 26390 8492
rect 26510 8440 26516 8492
rect 26568 8480 26574 8492
rect 26973 8483 27031 8489
rect 26973 8480 26985 8483
rect 26568 8452 26985 8480
rect 26568 8440 26574 8452
rect 26973 8449 26985 8452
rect 27019 8449 27031 8483
rect 26973 8443 27031 8449
rect 27341 8483 27399 8489
rect 27341 8449 27353 8483
rect 27387 8449 27399 8483
rect 27341 8443 27399 8449
rect 27356 8412 27384 8443
rect 27706 8440 27712 8492
rect 27764 8440 27770 8492
rect 26160 8384 27384 8412
rect 22428 8372 22434 8384
rect 17494 8344 17500 8356
rect 10612 8316 17500 8344
rect 17494 8304 17500 8316
rect 17552 8304 17558 8356
rect 23382 8304 23388 8356
rect 23440 8344 23446 8356
rect 23440 8316 24716 8344
rect 23440 8304 23446 8316
rect 9950 8236 9956 8288
rect 10008 8276 10014 8288
rect 13998 8276 14004 8288
rect 10008 8248 14004 8276
rect 10008 8236 10014 8248
rect 13998 8236 14004 8248
rect 14056 8236 14062 8288
rect 24688 8276 24716 8316
rect 24964 8276 24992 8384
rect 25038 8304 25044 8356
rect 25096 8344 25102 8356
rect 25317 8347 25375 8353
rect 25317 8344 25329 8347
rect 25096 8316 25329 8344
rect 25096 8304 25102 8316
rect 25317 8313 25329 8316
rect 25363 8313 25375 8347
rect 25317 8307 25375 8313
rect 25406 8304 25412 8356
rect 25464 8344 25470 8356
rect 26053 8347 26111 8353
rect 26053 8344 26065 8347
rect 25464 8316 26065 8344
rect 25464 8304 25470 8316
rect 26053 8313 26065 8316
rect 26099 8313 26111 8347
rect 26053 8307 26111 8313
rect 26142 8304 26148 8356
rect 26200 8344 26206 8356
rect 26421 8347 26479 8353
rect 26421 8344 26433 8347
rect 26200 8316 26433 8344
rect 26200 8304 26206 8316
rect 26421 8313 26433 8316
rect 26467 8313 26479 8347
rect 26421 8307 26479 8313
rect 26602 8304 26608 8356
rect 26660 8344 26666 8356
rect 27525 8347 27583 8353
rect 27525 8344 27537 8347
rect 26660 8316 27537 8344
rect 26660 8304 26666 8316
rect 27525 8313 27537 8316
rect 27571 8313 27583 8347
rect 27816 8344 27844 8520
rect 27982 8508 27988 8560
rect 28040 8548 28046 8560
rect 29012 8548 29040 8579
rect 29546 8576 29552 8628
rect 29604 8616 29610 8628
rect 30377 8619 30435 8625
rect 30377 8616 30389 8619
rect 29604 8588 30389 8616
rect 29604 8576 29610 8588
rect 30377 8585 30389 8588
rect 30423 8585 30435 8619
rect 30377 8579 30435 8585
rect 31110 8576 31116 8628
rect 31168 8576 31174 8628
rect 28040 8520 29040 8548
rect 29104 8520 30972 8548
rect 28040 8508 28046 8520
rect 28074 8440 28080 8492
rect 28132 8440 28138 8492
rect 28445 8483 28503 8489
rect 28445 8449 28457 8483
rect 28491 8449 28503 8483
rect 28445 8443 28503 8449
rect 28460 8412 28488 8443
rect 28810 8440 28816 8492
rect 28868 8440 28874 8492
rect 28902 8440 28908 8492
rect 28960 8480 28966 8492
rect 29104 8480 29132 8520
rect 28960 8452 29132 8480
rect 28960 8440 28966 8452
rect 29546 8440 29552 8492
rect 29604 8440 29610 8492
rect 29914 8440 29920 8492
rect 29972 8440 29978 8492
rect 30558 8440 30564 8492
rect 30616 8440 30622 8492
rect 30944 8489 30972 8520
rect 30929 8483 30987 8489
rect 30929 8449 30941 8483
rect 30975 8449 30987 8483
rect 30929 8443 30987 8449
rect 31294 8440 31300 8492
rect 31352 8440 31358 8492
rect 31662 8440 31668 8492
rect 31720 8440 31726 8492
rect 28000 8384 28488 8412
rect 27893 8347 27951 8353
rect 27893 8344 27905 8347
rect 27816 8316 27905 8344
rect 27525 8307 27583 8313
rect 27893 8313 27905 8316
rect 27939 8313 27951 8347
rect 27893 8307 27951 8313
rect 24688 8248 24992 8276
rect 27614 8236 27620 8288
rect 27672 8276 27678 8288
rect 28000 8276 28028 8384
rect 28994 8372 29000 8424
rect 29052 8412 29058 8424
rect 29052 8384 30144 8412
rect 29052 8372 29058 8384
rect 28718 8304 28724 8356
rect 28776 8344 28782 8356
rect 30116 8353 30144 8384
rect 29733 8347 29791 8353
rect 29733 8344 29745 8347
rect 28776 8316 29745 8344
rect 28776 8304 28782 8316
rect 29733 8313 29745 8316
rect 29779 8313 29791 8347
rect 29733 8307 29791 8313
rect 30101 8347 30159 8353
rect 30101 8313 30113 8347
rect 30147 8313 30159 8347
rect 30101 8307 30159 8313
rect 31481 8347 31539 8353
rect 31481 8313 31493 8347
rect 31527 8344 31539 8347
rect 32582 8344 32588 8356
rect 31527 8316 32588 8344
rect 31527 8313 31539 8316
rect 31481 8307 31539 8313
rect 32582 8304 32588 8316
rect 32640 8304 32646 8356
rect 27672 8248 28028 8276
rect 27672 8236 27678 8248
rect 31846 8236 31852 8288
rect 31904 8236 31910 8288
rect 1104 8186 32568 8208
rect 1104 8134 1950 8186
rect 2002 8134 2014 8186
rect 2066 8134 2078 8186
rect 2130 8134 2142 8186
rect 2194 8134 2206 8186
rect 2258 8134 7950 8186
rect 8002 8134 8014 8186
rect 8066 8134 8078 8186
rect 8130 8134 8142 8186
rect 8194 8134 8206 8186
rect 8258 8134 13950 8186
rect 14002 8134 14014 8186
rect 14066 8134 14078 8186
rect 14130 8134 14142 8186
rect 14194 8134 14206 8186
rect 14258 8134 19950 8186
rect 20002 8134 20014 8186
rect 20066 8134 20078 8186
rect 20130 8134 20142 8186
rect 20194 8134 20206 8186
rect 20258 8134 25950 8186
rect 26002 8134 26014 8186
rect 26066 8134 26078 8186
rect 26130 8134 26142 8186
rect 26194 8134 26206 8186
rect 26258 8134 31950 8186
rect 32002 8134 32014 8186
rect 32066 8134 32078 8186
rect 32130 8134 32142 8186
rect 32194 8134 32206 8186
rect 32258 8134 32568 8186
rect 1104 8112 32568 8134
rect 4154 8032 4160 8084
rect 4212 8072 4218 8084
rect 4341 8075 4399 8081
rect 4341 8072 4353 8075
rect 4212 8044 4353 8072
rect 4212 8032 4218 8044
rect 4341 8041 4353 8044
rect 4387 8041 4399 8075
rect 4341 8035 4399 8041
rect 5258 8032 5264 8084
rect 5316 8072 5322 8084
rect 5537 8075 5595 8081
rect 5537 8072 5549 8075
rect 5316 8044 5549 8072
rect 5316 8032 5322 8044
rect 5537 8041 5549 8044
rect 5583 8041 5595 8075
rect 5537 8035 5595 8041
rect 6086 8032 6092 8084
rect 6144 8072 6150 8084
rect 6273 8075 6331 8081
rect 6273 8072 6285 8075
rect 6144 8044 6285 8072
rect 6144 8032 6150 8044
rect 6273 8041 6285 8044
rect 6319 8041 6331 8075
rect 6273 8035 6331 8041
rect 6638 8032 6644 8084
rect 6696 8072 6702 8084
rect 6825 8075 6883 8081
rect 6825 8072 6837 8075
rect 6696 8044 6837 8072
rect 6696 8032 6702 8044
rect 6825 8041 6837 8044
rect 6871 8041 6883 8075
rect 6825 8035 6883 8041
rect 7466 8032 7472 8084
rect 7524 8072 7530 8084
rect 7745 8075 7803 8081
rect 7745 8072 7757 8075
rect 7524 8044 7757 8072
rect 7524 8032 7530 8044
rect 7745 8041 7757 8044
rect 7791 8041 7803 8075
rect 7745 8035 7803 8041
rect 8294 8032 8300 8084
rect 8352 8072 8358 8084
rect 8481 8075 8539 8081
rect 8481 8072 8493 8075
rect 8352 8044 8493 8072
rect 8352 8032 8358 8044
rect 8481 8041 8493 8044
rect 8527 8041 8539 8075
rect 8481 8035 8539 8041
rect 8846 8032 8852 8084
rect 8904 8072 8910 8084
rect 9309 8075 9367 8081
rect 9309 8072 9321 8075
rect 8904 8044 9321 8072
rect 8904 8032 8910 8044
rect 9309 8041 9321 8044
rect 9355 8041 9367 8075
rect 9309 8035 9367 8041
rect 9674 8032 9680 8084
rect 9732 8072 9738 8084
rect 9861 8075 9919 8081
rect 9861 8072 9873 8075
rect 9732 8044 9873 8072
rect 9732 8032 9738 8044
rect 9861 8041 9873 8044
rect 9907 8041 9919 8075
rect 9861 8035 9919 8041
rect 10778 8032 10784 8084
rect 10836 8072 10842 8084
rect 10965 8075 11023 8081
rect 10965 8072 10977 8075
rect 10836 8044 10977 8072
rect 10836 8032 10842 8044
rect 10965 8041 10977 8044
rect 11011 8041 11023 8075
rect 10965 8035 11023 8041
rect 11330 8032 11336 8084
rect 11388 8072 11394 8084
rect 11517 8075 11575 8081
rect 11517 8072 11529 8075
rect 11388 8044 11529 8072
rect 11388 8032 11394 8044
rect 11517 8041 11529 8044
rect 11563 8041 11575 8075
rect 11517 8035 11575 8041
rect 11882 8032 11888 8084
rect 11940 8072 11946 8084
rect 12069 8075 12127 8081
rect 12069 8072 12081 8075
rect 11940 8044 12081 8072
rect 11940 8032 11946 8044
rect 12069 8041 12081 8044
rect 12115 8041 12127 8075
rect 12069 8035 12127 8041
rect 25866 8032 25872 8084
rect 25924 8072 25930 8084
rect 26145 8075 26203 8081
rect 26145 8072 26157 8075
rect 25924 8044 26157 8072
rect 25924 8032 25930 8044
rect 26145 8041 26157 8044
rect 26191 8041 26203 8075
rect 26145 8035 26203 8041
rect 27338 8032 27344 8084
rect 27396 8032 27402 8084
rect 28166 8032 28172 8084
rect 28224 8072 28230 8084
rect 28445 8075 28503 8081
rect 28445 8072 28457 8075
rect 28224 8044 28457 8072
rect 28224 8032 28230 8044
rect 28445 8041 28457 8044
rect 28491 8041 28503 8075
rect 28445 8035 28503 8041
rect 28534 8032 28540 8084
rect 28592 8072 28598 8084
rect 28813 8075 28871 8081
rect 28813 8072 28825 8075
rect 28592 8044 28825 8072
rect 28592 8032 28598 8044
rect 28813 8041 28825 8044
rect 28859 8041 28871 8075
rect 28813 8035 28871 8041
rect 29270 8032 29276 8084
rect 29328 8072 29334 8084
rect 29733 8075 29791 8081
rect 29733 8072 29745 8075
rect 29328 8044 29745 8072
rect 29328 8032 29334 8044
rect 29733 8041 29745 8044
rect 29779 8041 29791 8075
rect 29733 8035 29791 8041
rect 30650 8032 30656 8084
rect 30708 8032 30714 8084
rect 31018 8032 31024 8084
rect 31076 8032 31082 8084
rect 31386 8032 31392 8084
rect 31444 8032 31450 8084
rect 10042 7964 10048 8016
rect 10100 8004 10106 8016
rect 19334 8004 19340 8016
rect 10100 7976 19340 8004
rect 10100 7964 10106 7976
rect 19334 7964 19340 7976
rect 19392 7964 19398 8016
rect 8478 7896 8484 7948
rect 8536 7936 8542 7948
rect 20806 7936 20812 7948
rect 8536 7908 20812 7936
rect 8536 7896 8542 7908
rect 20806 7896 20812 7908
rect 20864 7896 20870 7948
rect 27614 7896 27620 7948
rect 27672 7936 27678 7948
rect 27672 7908 31616 7936
rect 27672 7896 27678 7908
rect 4525 7871 4583 7877
rect 4525 7837 4537 7871
rect 4571 7837 4583 7871
rect 4525 7831 4583 7837
rect 4540 7800 4568 7831
rect 5350 7828 5356 7880
rect 5408 7828 5414 7880
rect 6457 7871 6515 7877
rect 6457 7837 6469 7871
rect 6503 7868 6515 7871
rect 6914 7868 6920 7880
rect 6503 7840 6920 7868
rect 6503 7837 6515 7840
rect 6457 7831 6515 7837
rect 6914 7828 6920 7840
rect 6972 7828 6978 7880
rect 7009 7871 7067 7877
rect 7009 7837 7021 7871
rect 7055 7837 7067 7871
rect 7009 7831 7067 7837
rect 6270 7800 6276 7812
rect 4540 7772 6276 7800
rect 6270 7760 6276 7772
rect 6328 7760 6334 7812
rect 7024 7800 7052 7831
rect 7190 7828 7196 7880
rect 7248 7868 7254 7880
rect 7561 7871 7619 7877
rect 7561 7868 7573 7871
rect 7248 7840 7573 7868
rect 7248 7828 7254 7840
rect 7561 7837 7573 7840
rect 7607 7837 7619 7871
rect 7561 7831 7619 7837
rect 8662 7828 8668 7880
rect 8720 7828 8726 7880
rect 9490 7828 9496 7880
rect 9548 7828 9554 7880
rect 10042 7828 10048 7880
rect 10100 7828 10106 7880
rect 11149 7871 11207 7877
rect 11149 7837 11161 7871
rect 11195 7837 11207 7871
rect 11149 7831 11207 7837
rect 11701 7871 11759 7877
rect 11701 7837 11713 7871
rect 11747 7837 11759 7871
rect 11701 7831 11759 7837
rect 12253 7871 12311 7877
rect 12253 7837 12265 7871
rect 12299 7868 12311 7871
rect 12618 7868 12624 7880
rect 12299 7840 12624 7868
rect 12299 7837 12311 7840
rect 12253 7831 12311 7837
rect 9398 7800 9404 7812
rect 7024 7772 9404 7800
rect 9398 7760 9404 7772
rect 9456 7760 9462 7812
rect 11164 7732 11192 7831
rect 11716 7800 11744 7831
rect 12618 7828 12624 7840
rect 12676 7828 12682 7880
rect 25866 7828 25872 7880
rect 25924 7868 25930 7880
rect 26329 7871 26387 7877
rect 26329 7868 26341 7871
rect 25924 7840 26341 7868
rect 25924 7828 25930 7840
rect 26329 7837 26341 7840
rect 26375 7837 26387 7871
rect 26329 7831 26387 7837
rect 27157 7871 27215 7877
rect 27157 7837 27169 7871
rect 27203 7837 27215 7871
rect 27157 7831 27215 7837
rect 14366 7800 14372 7812
rect 11716 7772 14372 7800
rect 14366 7760 14372 7772
rect 14424 7760 14430 7812
rect 21450 7760 21456 7812
rect 21508 7800 21514 7812
rect 27172 7800 27200 7831
rect 28258 7828 28264 7880
rect 28316 7828 28322 7880
rect 28626 7828 28632 7880
rect 28684 7828 28690 7880
rect 29086 7828 29092 7880
rect 29144 7868 29150 7880
rect 29549 7871 29607 7877
rect 29549 7868 29561 7871
rect 29144 7840 29561 7868
rect 29144 7828 29150 7840
rect 29549 7837 29561 7840
rect 29595 7837 29607 7871
rect 29549 7831 29607 7837
rect 30466 7828 30472 7880
rect 30524 7828 30530 7880
rect 30650 7828 30656 7880
rect 30708 7868 30714 7880
rect 30837 7871 30895 7877
rect 30837 7868 30849 7871
rect 30708 7840 30849 7868
rect 30708 7828 30714 7840
rect 30837 7837 30849 7840
rect 30883 7837 30895 7871
rect 30837 7831 30895 7837
rect 30926 7828 30932 7880
rect 30984 7868 30990 7880
rect 31588 7877 31616 7908
rect 31205 7871 31263 7877
rect 31205 7868 31217 7871
rect 30984 7840 31217 7868
rect 30984 7828 30990 7840
rect 31205 7837 31217 7840
rect 31251 7837 31263 7871
rect 31205 7831 31263 7837
rect 31573 7871 31631 7877
rect 31573 7837 31585 7871
rect 31619 7837 31631 7871
rect 31573 7831 31631 7837
rect 31941 7871 31999 7877
rect 31941 7837 31953 7871
rect 31987 7837 31999 7871
rect 31941 7831 31999 7837
rect 21508 7772 27200 7800
rect 21508 7760 21514 7772
rect 28994 7760 29000 7812
rect 29052 7800 29058 7812
rect 31956 7800 31984 7831
rect 29052 7772 31984 7800
rect 29052 7760 29058 7772
rect 16482 7732 16488 7744
rect 11164 7704 16488 7732
rect 16482 7692 16488 7704
rect 16540 7692 16546 7744
rect 26234 7692 26240 7744
rect 26292 7732 26298 7744
rect 31294 7732 31300 7744
rect 26292 7704 31300 7732
rect 26292 7692 26298 7704
rect 31294 7692 31300 7704
rect 31352 7692 31358 7744
rect 31754 7692 31760 7744
rect 31812 7692 31818 7744
rect 32122 7692 32128 7744
rect 32180 7692 32186 7744
rect 1104 7642 32568 7664
rect 1104 7590 3010 7642
rect 3062 7590 3074 7642
rect 3126 7590 3138 7642
rect 3190 7590 3202 7642
rect 3254 7590 3266 7642
rect 3318 7590 9010 7642
rect 9062 7590 9074 7642
rect 9126 7590 9138 7642
rect 9190 7590 9202 7642
rect 9254 7590 9266 7642
rect 9318 7590 15010 7642
rect 15062 7590 15074 7642
rect 15126 7590 15138 7642
rect 15190 7590 15202 7642
rect 15254 7590 15266 7642
rect 15318 7590 21010 7642
rect 21062 7590 21074 7642
rect 21126 7590 21138 7642
rect 21190 7590 21202 7642
rect 21254 7590 21266 7642
rect 21318 7590 27010 7642
rect 27062 7590 27074 7642
rect 27126 7590 27138 7642
rect 27190 7590 27202 7642
rect 27254 7590 27266 7642
rect 27318 7590 32568 7642
rect 1104 7568 32568 7590
rect 23106 7488 23112 7540
rect 23164 7488 23170 7540
rect 24486 7488 24492 7540
rect 24544 7488 24550 7540
rect 28994 7528 29000 7540
rect 24596 7500 29000 7528
rect 10042 7420 10048 7472
rect 10100 7460 10106 7472
rect 10100 7432 16804 7460
rect 10100 7420 10106 7432
rect 10870 7352 10876 7404
rect 10928 7392 10934 7404
rect 16776 7392 16804 7432
rect 16850 7420 16856 7472
rect 16908 7460 16914 7472
rect 24596 7460 24624 7500
rect 28994 7488 29000 7500
rect 29052 7488 29058 7540
rect 31478 7488 31484 7540
rect 31536 7488 31542 7540
rect 16908 7432 24624 7460
rect 26237 7463 26295 7469
rect 16908 7420 16914 7432
rect 26237 7429 26249 7463
rect 26283 7460 26295 7463
rect 26418 7460 26424 7472
rect 26283 7432 26424 7460
rect 26283 7429 26295 7432
rect 26237 7423 26295 7429
rect 20806 7392 20812 7404
rect 10928 7364 16528 7392
rect 16776 7364 20812 7392
rect 10928 7352 10934 7364
rect 16500 7256 16528 7364
rect 20806 7352 20812 7364
rect 20864 7352 20870 7404
rect 22005 7395 22063 7401
rect 22005 7361 22017 7395
rect 22051 7392 22063 7395
rect 23106 7392 23112 7404
rect 22051 7364 23112 7392
rect 22051 7361 22063 7364
rect 22005 7355 22063 7361
rect 23106 7352 23112 7364
rect 23164 7352 23170 7404
rect 26344 7401 26372 7432
rect 26418 7420 26424 7432
rect 26476 7420 26482 7472
rect 26878 7420 26884 7472
rect 26936 7460 26942 7472
rect 27433 7463 27491 7469
rect 27433 7460 27445 7463
rect 26936 7432 27445 7460
rect 26936 7420 26942 7432
rect 27433 7429 27445 7432
rect 27479 7429 27491 7463
rect 27433 7423 27491 7429
rect 23201 7395 23259 7401
rect 23201 7361 23213 7395
rect 23247 7392 23259 7395
rect 23293 7395 23351 7401
rect 23293 7392 23305 7395
rect 23247 7364 23305 7392
rect 23247 7361 23259 7364
rect 23201 7355 23259 7361
rect 23293 7361 23305 7364
rect 23339 7361 23351 7395
rect 23293 7355 23351 7361
rect 24581 7395 24639 7401
rect 24581 7361 24593 7395
rect 24627 7392 24639 7395
rect 24673 7395 24731 7401
rect 24673 7392 24685 7395
rect 24627 7364 24685 7392
rect 24627 7361 24639 7364
rect 24581 7355 24639 7361
rect 24673 7361 24685 7364
rect 24719 7361 24731 7395
rect 24673 7355 24731 7361
rect 26329 7395 26387 7401
rect 26329 7361 26341 7395
rect 26375 7392 26387 7395
rect 27525 7395 27583 7401
rect 26375 7364 26409 7392
rect 26375 7361 26387 7364
rect 26329 7355 26387 7361
rect 27525 7361 27537 7395
rect 27571 7392 27583 7395
rect 27617 7395 27675 7401
rect 27617 7392 27629 7395
rect 27571 7364 27629 7392
rect 27571 7361 27583 7364
rect 27525 7355 27583 7361
rect 27617 7361 27629 7364
rect 27663 7361 27675 7395
rect 27617 7355 27675 7361
rect 31297 7395 31355 7401
rect 31297 7361 31309 7395
rect 31343 7361 31355 7395
rect 31297 7355 31355 7361
rect 31665 7395 31723 7401
rect 31665 7361 31677 7395
rect 31711 7361 31723 7395
rect 31665 7355 31723 7361
rect 16574 7284 16580 7336
rect 16632 7324 16638 7336
rect 31312 7324 31340 7355
rect 16632 7296 31340 7324
rect 16632 7284 16638 7296
rect 17402 7256 17408 7268
rect 16500 7228 17408 7256
rect 17402 7216 17408 7228
rect 17460 7216 17466 7268
rect 23477 7259 23535 7265
rect 23477 7225 23489 7259
rect 23523 7256 23535 7259
rect 26234 7256 26240 7268
rect 23523 7228 26240 7256
rect 23523 7225 23535 7228
rect 23477 7219 23535 7225
rect 26234 7216 26240 7228
rect 26292 7216 26298 7268
rect 26513 7259 26571 7265
rect 26513 7225 26525 7259
rect 26559 7256 26571 7259
rect 28902 7256 28908 7268
rect 26559 7228 28908 7256
rect 26559 7225 26571 7228
rect 26513 7219 26571 7225
rect 28902 7216 28908 7228
rect 28960 7216 28966 7268
rect 30374 7216 30380 7268
rect 30432 7256 30438 7268
rect 31680 7256 31708 7355
rect 30432 7228 31708 7256
rect 30432 7216 30438 7228
rect 10134 7148 10140 7200
rect 10192 7188 10198 7200
rect 17678 7188 17684 7200
rect 10192 7160 17684 7188
rect 10192 7148 10198 7160
rect 17678 7148 17684 7160
rect 17736 7148 17742 7200
rect 22189 7191 22247 7197
rect 22189 7157 22201 7191
rect 22235 7188 22247 7191
rect 23658 7188 23664 7200
rect 22235 7160 23664 7188
rect 22235 7157 22247 7160
rect 22189 7151 22247 7157
rect 23658 7148 23664 7160
rect 23716 7148 23722 7200
rect 24857 7191 24915 7197
rect 24857 7157 24869 7191
rect 24903 7188 24915 7191
rect 27430 7188 27436 7200
rect 24903 7160 27436 7188
rect 24903 7157 24915 7160
rect 24857 7151 24915 7157
rect 27430 7148 27436 7160
rect 27488 7148 27494 7200
rect 27801 7191 27859 7197
rect 27801 7157 27813 7191
rect 27847 7188 27859 7191
rect 30282 7188 30288 7200
rect 27847 7160 30288 7188
rect 27847 7157 27859 7160
rect 27801 7151 27859 7157
rect 30282 7148 30288 7160
rect 30340 7148 30346 7200
rect 31849 7191 31907 7197
rect 31849 7157 31861 7191
rect 31895 7188 31907 7191
rect 32766 7188 32772 7200
rect 31895 7160 32772 7188
rect 31895 7157 31907 7160
rect 31849 7151 31907 7157
rect 32766 7148 32772 7160
rect 32824 7148 32830 7200
rect 1104 7098 32568 7120
rect 1104 7046 1950 7098
rect 2002 7046 2014 7098
rect 2066 7046 2078 7098
rect 2130 7046 2142 7098
rect 2194 7046 2206 7098
rect 2258 7046 7950 7098
rect 8002 7046 8014 7098
rect 8066 7046 8078 7098
rect 8130 7046 8142 7098
rect 8194 7046 8206 7098
rect 8258 7046 13950 7098
rect 14002 7046 14014 7098
rect 14066 7046 14078 7098
rect 14130 7046 14142 7098
rect 14194 7046 14206 7098
rect 14258 7046 19950 7098
rect 20002 7046 20014 7098
rect 20066 7046 20078 7098
rect 20130 7046 20142 7098
rect 20194 7046 20206 7098
rect 20258 7046 25950 7098
rect 26002 7046 26014 7098
rect 26066 7046 26078 7098
rect 26130 7046 26142 7098
rect 26194 7046 26206 7098
rect 26258 7046 31950 7098
rect 32002 7046 32014 7098
rect 32066 7046 32078 7098
rect 32130 7046 32142 7098
rect 32194 7046 32206 7098
rect 32258 7046 32568 7098
rect 1104 7024 32568 7046
rect 4433 6987 4491 6993
rect 4433 6953 4445 6987
rect 4479 6984 4491 6987
rect 5350 6984 5356 6996
rect 4479 6956 5356 6984
rect 4479 6953 4491 6956
rect 4433 6947 4491 6953
rect 5350 6944 5356 6956
rect 5408 6944 5414 6996
rect 6270 6944 6276 6996
rect 6328 6944 6334 6996
rect 12618 6944 12624 6996
rect 12676 6944 12682 6996
rect 14366 6944 14372 6996
rect 14424 6944 14430 6996
rect 16574 6944 16580 6996
rect 16632 6944 16638 6996
rect 16850 6944 16856 6996
rect 16908 6944 16914 6996
rect 19242 6944 19248 6996
rect 19300 6984 19306 6996
rect 19797 6987 19855 6993
rect 19797 6984 19809 6987
rect 19300 6956 19809 6984
rect 19300 6944 19306 6956
rect 19797 6953 19809 6956
rect 19843 6953 19855 6987
rect 19797 6947 19855 6953
rect 20717 6987 20775 6993
rect 20717 6953 20729 6987
rect 20763 6984 20775 6987
rect 20806 6984 20812 6996
rect 20763 6956 20812 6984
rect 20763 6953 20775 6956
rect 20717 6947 20775 6953
rect 20806 6944 20812 6956
rect 20864 6944 20870 6996
rect 21818 6984 21824 6996
rect 21284 6956 21824 6984
rect 7098 6808 7104 6860
rect 7156 6848 7162 6860
rect 10962 6848 10968 6860
rect 7156 6820 10968 6848
rect 7156 6808 7162 6820
rect 10962 6808 10968 6820
rect 11020 6808 11026 6860
rect 20714 6848 20720 6860
rect 11072 6820 13584 6848
rect 4249 6783 4307 6789
rect 4249 6749 4261 6783
rect 4295 6749 4307 6783
rect 4249 6743 4307 6749
rect 4264 6712 4292 6743
rect 6454 6740 6460 6792
rect 6512 6740 6518 6792
rect 7834 6740 7840 6792
rect 7892 6780 7898 6792
rect 8021 6783 8079 6789
rect 8021 6780 8033 6783
rect 7892 6752 8033 6780
rect 7892 6740 7898 6752
rect 8021 6749 8033 6752
rect 8067 6749 8079 6783
rect 8021 6743 8079 6749
rect 10134 6740 10140 6792
rect 10192 6740 10198 6792
rect 10229 6783 10287 6789
rect 10229 6749 10241 6783
rect 10275 6780 10287 6783
rect 10410 6780 10416 6792
rect 10275 6752 10416 6780
rect 10275 6749 10287 6752
rect 10229 6743 10287 6749
rect 10410 6740 10416 6752
rect 10468 6740 10474 6792
rect 10597 6783 10655 6789
rect 10597 6749 10609 6783
rect 10643 6780 10655 6783
rect 10686 6780 10692 6792
rect 10643 6752 10692 6780
rect 10643 6749 10655 6752
rect 10597 6743 10655 6749
rect 10686 6740 10692 6752
rect 10744 6740 10750 6792
rect 11072 6789 11100 6820
rect 11057 6783 11115 6789
rect 11057 6749 11069 6783
rect 11103 6749 11115 6783
rect 11057 6743 11115 6749
rect 11333 6783 11391 6789
rect 11333 6749 11345 6783
rect 11379 6780 11391 6783
rect 11422 6780 11428 6792
rect 11379 6752 11428 6780
rect 11379 6749 11391 6752
rect 11333 6743 11391 6749
rect 11422 6740 11428 6752
rect 11480 6740 11486 6792
rect 11609 6783 11667 6789
rect 11609 6749 11621 6783
rect 11655 6780 11667 6783
rect 12066 6780 12072 6792
rect 11655 6752 12072 6780
rect 11655 6749 11667 6752
rect 11609 6743 11667 6749
rect 12066 6740 12072 6752
rect 12124 6740 12130 6792
rect 12802 6740 12808 6792
rect 12860 6740 12866 6792
rect 9674 6712 9680 6724
rect 4264 6684 9680 6712
rect 9674 6672 9680 6684
rect 9732 6672 9738 6724
rect 13354 6712 13360 6724
rect 10888 6684 13360 6712
rect 4338 6604 4344 6656
rect 4396 6644 4402 6656
rect 7837 6647 7895 6653
rect 7837 6644 7849 6647
rect 4396 6616 7849 6644
rect 4396 6604 4402 6616
rect 7837 6613 7849 6616
rect 7883 6613 7895 6647
rect 7837 6607 7895 6613
rect 9490 6604 9496 6656
rect 9548 6644 9554 6656
rect 9953 6647 10011 6653
rect 9953 6644 9965 6647
rect 9548 6616 9965 6644
rect 9548 6604 9554 6616
rect 9953 6613 9965 6616
rect 9999 6613 10011 6647
rect 9953 6607 10011 6613
rect 10413 6647 10471 6653
rect 10413 6613 10425 6647
rect 10459 6644 10471 6647
rect 10594 6644 10600 6656
rect 10459 6616 10600 6644
rect 10459 6613 10471 6616
rect 10413 6607 10471 6613
rect 10594 6604 10600 6616
rect 10652 6604 10658 6656
rect 10888 6653 10916 6684
rect 13354 6672 13360 6684
rect 13412 6672 13418 6724
rect 13556 6712 13584 6820
rect 13648 6820 17264 6848
rect 13648 6789 13676 6820
rect 13633 6783 13691 6789
rect 13633 6749 13645 6783
rect 13679 6749 13691 6783
rect 13633 6743 13691 6749
rect 14553 6783 14611 6789
rect 14553 6749 14565 6783
rect 14599 6780 14611 6783
rect 15654 6780 15660 6792
rect 14599 6752 15660 6780
rect 14599 6749 14611 6752
rect 14553 6743 14611 6749
rect 15654 6740 15660 6752
rect 15712 6740 15718 6792
rect 15746 6740 15752 6792
rect 15804 6740 15810 6792
rect 16114 6740 16120 6792
rect 16172 6780 16178 6792
rect 16209 6783 16267 6789
rect 16209 6780 16221 6783
rect 16172 6752 16221 6780
rect 16172 6740 16178 6752
rect 16209 6749 16221 6752
rect 16255 6780 16267 6783
rect 16393 6783 16451 6789
rect 16393 6780 16405 6783
rect 16255 6752 16405 6780
rect 16255 6749 16267 6752
rect 16209 6743 16267 6749
rect 16393 6749 16405 6752
rect 16439 6749 16451 6783
rect 16393 6743 16451 6749
rect 16666 6740 16672 6792
rect 16724 6780 16730 6792
rect 16945 6783 17003 6789
rect 16945 6780 16957 6783
rect 16724 6752 16957 6780
rect 16724 6740 16730 6752
rect 16945 6749 16957 6752
rect 16991 6749 17003 6783
rect 16945 6743 17003 6749
rect 16298 6712 16304 6724
rect 13556 6684 16304 6712
rect 16298 6672 16304 6684
rect 16356 6672 16362 6724
rect 16482 6672 16488 6724
rect 16540 6712 16546 6724
rect 17236 6712 17264 6820
rect 17328 6820 20720 6848
rect 17328 6789 17356 6820
rect 20714 6808 20720 6820
rect 20772 6808 20778 6860
rect 21284 6848 21312 6956
rect 21818 6944 21824 6956
rect 21876 6944 21882 6996
rect 26605 6987 26663 6993
rect 26605 6953 26617 6987
rect 26651 6984 26663 6987
rect 26694 6984 26700 6996
rect 26651 6956 26700 6984
rect 26651 6953 26663 6956
rect 26605 6947 26663 6953
rect 26694 6944 26700 6956
rect 26752 6944 26758 6996
rect 21361 6919 21419 6925
rect 21361 6885 21373 6919
rect 21407 6885 21419 6919
rect 21361 6879 21419 6885
rect 24581 6919 24639 6925
rect 24581 6885 24593 6919
rect 24627 6914 24639 6919
rect 24627 6886 24661 6914
rect 25884 6888 26096 6916
rect 24627 6885 24639 6886
rect 24581 6879 24639 6885
rect 20824 6820 21312 6848
rect 21376 6848 21404 6879
rect 22830 6848 22836 6860
rect 21376 6820 22836 6848
rect 17313 6783 17371 6789
rect 17313 6749 17325 6783
rect 17359 6749 17371 6783
rect 17313 6743 17371 6749
rect 17678 6740 17684 6792
rect 17736 6740 17742 6792
rect 18414 6740 18420 6792
rect 18472 6740 18478 6792
rect 19334 6740 19340 6792
rect 19392 6780 19398 6792
rect 19613 6783 19671 6789
rect 19613 6780 19625 6783
rect 19392 6752 19625 6780
rect 19392 6740 19398 6752
rect 19613 6749 19625 6752
rect 19659 6749 19671 6783
rect 19613 6743 19671 6749
rect 19978 6740 19984 6792
rect 20036 6740 20042 6792
rect 20824 6712 20852 6820
rect 22830 6808 22836 6820
rect 22888 6808 22894 6860
rect 23474 6808 23480 6860
rect 23532 6808 23538 6860
rect 24596 6848 24624 6879
rect 25884 6848 25912 6888
rect 24596 6820 25912 6848
rect 26068 6848 26096 6888
rect 29546 6848 29552 6860
rect 26068 6820 29552 6848
rect 29546 6808 29552 6820
rect 29604 6808 29610 6860
rect 30282 6808 30288 6860
rect 30340 6848 30346 6860
rect 30340 6820 31984 6848
rect 30340 6808 30346 6820
rect 20901 6783 20959 6789
rect 20901 6749 20913 6783
rect 20947 6749 20959 6783
rect 20901 6743 20959 6749
rect 16540 6684 17172 6712
rect 17236 6684 20852 6712
rect 20916 6712 20944 6743
rect 20990 6740 20996 6792
rect 21048 6780 21054 6792
rect 21177 6783 21235 6789
rect 21177 6780 21189 6783
rect 21048 6752 21189 6780
rect 21048 6740 21054 6752
rect 21177 6749 21189 6752
rect 21223 6749 21235 6783
rect 21177 6743 21235 6749
rect 21453 6783 21511 6789
rect 21453 6749 21465 6783
rect 21499 6780 21511 6783
rect 21634 6780 21640 6792
rect 21499 6752 21640 6780
rect 21499 6749 21511 6752
rect 21453 6743 21511 6749
rect 21634 6740 21640 6752
rect 21692 6780 21698 6792
rect 21729 6783 21787 6789
rect 21729 6780 21741 6783
rect 21692 6752 21741 6780
rect 21692 6740 21698 6752
rect 21729 6749 21741 6752
rect 21775 6749 21787 6783
rect 21729 6743 21787 6749
rect 23290 6740 23296 6792
rect 23348 6780 23354 6792
rect 23385 6783 23443 6789
rect 23385 6780 23397 6783
rect 23348 6752 23397 6780
rect 23348 6740 23354 6752
rect 23385 6749 23397 6752
rect 23431 6749 23443 6783
rect 23385 6743 23443 6749
rect 23492 6712 23520 6808
rect 23658 6740 23664 6792
rect 23716 6740 23722 6792
rect 24394 6740 24400 6792
rect 24452 6740 24458 6792
rect 26053 6783 26111 6789
rect 26053 6749 26065 6783
rect 26099 6776 26111 6783
rect 26145 6783 26203 6789
rect 26145 6776 26157 6783
rect 26099 6749 26157 6776
rect 26191 6749 26203 6783
rect 26053 6748 26203 6749
rect 26053 6743 26111 6748
rect 26145 6743 26203 6748
rect 26421 6783 26479 6789
rect 26421 6749 26433 6783
rect 26467 6780 26479 6783
rect 29362 6780 29368 6792
rect 26467 6752 29368 6780
rect 26467 6749 26479 6752
rect 26421 6743 26479 6749
rect 29362 6740 29368 6752
rect 29420 6740 29426 6792
rect 31205 6783 31263 6789
rect 31205 6749 31217 6783
rect 31251 6749 31263 6783
rect 31205 6743 31263 6749
rect 31573 6783 31631 6789
rect 31573 6749 31585 6783
rect 31619 6780 31631 6783
rect 31662 6780 31668 6792
rect 31619 6752 31668 6780
rect 31619 6749 31631 6752
rect 31573 6743 31631 6749
rect 20916 6684 23520 6712
rect 16540 6672 16546 6684
rect 10873 6647 10931 6653
rect 10873 6613 10885 6647
rect 10919 6613 10931 6647
rect 10873 6607 10931 6613
rect 11238 6604 11244 6656
rect 11296 6604 11302 6656
rect 11514 6604 11520 6656
rect 11572 6604 11578 6656
rect 11793 6647 11851 6653
rect 11793 6613 11805 6647
rect 11839 6644 11851 6647
rect 11974 6644 11980 6656
rect 11839 6616 11980 6644
rect 11839 6613 11851 6616
rect 11793 6607 11851 6613
rect 11974 6604 11980 6616
rect 12032 6604 12038 6656
rect 13446 6604 13452 6656
rect 13504 6604 13510 6656
rect 15562 6604 15568 6656
rect 15620 6604 15626 6656
rect 17144 6653 17172 6684
rect 25774 6672 25780 6724
rect 25832 6712 25838 6724
rect 25961 6715 26019 6721
rect 25961 6712 25973 6715
rect 25832 6684 25973 6712
rect 25832 6672 25838 6684
rect 25961 6681 25973 6684
rect 26007 6681 26019 6715
rect 30926 6712 30932 6724
rect 25961 6675 26019 6681
rect 26206 6684 30932 6712
rect 17129 6647 17187 6653
rect 17129 6613 17141 6647
rect 17175 6613 17187 6647
rect 17129 6607 17187 6613
rect 17494 6604 17500 6656
rect 17552 6604 17558 6656
rect 18230 6604 18236 6656
rect 18288 6604 18294 6656
rect 19518 6604 19524 6656
rect 19576 6604 19582 6656
rect 20806 6604 20812 6656
rect 20864 6644 20870 6656
rect 21542 6644 21548 6656
rect 20864 6616 21548 6644
rect 20864 6604 20870 6616
rect 21542 6604 21548 6616
rect 21600 6604 21606 6656
rect 21634 6604 21640 6656
rect 21692 6604 21698 6656
rect 22186 6604 22192 6656
rect 22244 6644 22250 6656
rect 22922 6644 22928 6656
rect 22244 6616 22928 6644
rect 22244 6604 22250 6616
rect 22922 6604 22928 6616
rect 22980 6604 22986 6656
rect 23566 6604 23572 6656
rect 23624 6604 23630 6656
rect 23842 6604 23848 6656
rect 23900 6604 23906 6656
rect 23934 6604 23940 6656
rect 23992 6644 23998 6656
rect 26206 6644 26234 6684
rect 30926 6672 30932 6684
rect 30984 6672 30990 6724
rect 23992 6616 26234 6644
rect 26329 6647 26387 6653
rect 23992 6604 23998 6616
rect 26329 6613 26341 6647
rect 26375 6644 26387 6647
rect 27614 6644 27620 6656
rect 26375 6616 27620 6644
rect 26375 6613 26387 6616
rect 26329 6607 26387 6613
rect 27614 6604 27620 6616
rect 27672 6604 27678 6656
rect 28718 6604 28724 6656
rect 28776 6644 28782 6656
rect 31220 6644 31248 6743
rect 31662 6740 31668 6752
rect 31720 6740 31726 6792
rect 31956 6789 31984 6820
rect 31941 6783 31999 6789
rect 31941 6749 31953 6783
rect 31987 6749 31999 6783
rect 31941 6743 31999 6749
rect 28776 6616 31248 6644
rect 28776 6604 28782 6616
rect 31386 6604 31392 6656
rect 31444 6604 31450 6656
rect 31754 6604 31760 6656
rect 31812 6604 31818 6656
rect 32125 6647 32183 6653
rect 32125 6613 32137 6647
rect 32171 6644 32183 6647
rect 32306 6644 32312 6656
rect 32171 6616 32312 6644
rect 32171 6613 32183 6616
rect 32125 6607 32183 6613
rect 32306 6604 32312 6616
rect 32364 6604 32370 6656
rect 1104 6554 32568 6576
rect 1104 6502 3010 6554
rect 3062 6502 3074 6554
rect 3126 6502 3138 6554
rect 3190 6502 3202 6554
rect 3254 6502 3266 6554
rect 3318 6502 9010 6554
rect 9062 6502 9074 6554
rect 9126 6502 9138 6554
rect 9190 6502 9202 6554
rect 9254 6502 9266 6554
rect 9318 6502 15010 6554
rect 15062 6502 15074 6554
rect 15126 6502 15138 6554
rect 15190 6502 15202 6554
rect 15254 6502 15266 6554
rect 15318 6502 21010 6554
rect 21062 6502 21074 6554
rect 21126 6502 21138 6554
rect 21190 6502 21202 6554
rect 21254 6502 21266 6554
rect 21318 6502 27010 6554
rect 27062 6502 27074 6554
rect 27126 6502 27138 6554
rect 27190 6502 27202 6554
rect 27254 6502 27266 6554
rect 27318 6502 32568 6554
rect 1104 6480 32568 6502
rect 5166 6400 5172 6452
rect 5224 6440 5230 6452
rect 5261 6443 5319 6449
rect 5261 6440 5273 6443
rect 5224 6412 5273 6440
rect 5224 6400 5230 6412
rect 5261 6409 5273 6412
rect 5307 6409 5319 6443
rect 5261 6403 5319 6409
rect 5810 6400 5816 6452
rect 5868 6440 5874 6452
rect 6641 6443 6699 6449
rect 6641 6440 6653 6443
rect 5868 6412 6653 6440
rect 5868 6400 5874 6412
rect 6641 6409 6653 6412
rect 6687 6409 6699 6443
rect 6641 6403 6699 6409
rect 6914 6400 6920 6452
rect 6972 6440 6978 6452
rect 7653 6443 7711 6449
rect 7653 6440 7665 6443
rect 6972 6412 7665 6440
rect 6972 6400 6978 6412
rect 7653 6409 7665 6412
rect 7699 6409 7711 6443
rect 7653 6403 7711 6409
rect 8386 6400 8392 6452
rect 8444 6400 8450 6452
rect 8662 6400 8668 6452
rect 8720 6400 8726 6452
rect 8754 6400 8760 6452
rect 8812 6440 8818 6452
rect 9217 6443 9275 6449
rect 9217 6440 9229 6443
rect 8812 6412 9229 6440
rect 8812 6400 8818 6412
rect 9217 6409 9229 6412
rect 9263 6409 9275 6443
rect 9217 6403 9275 6409
rect 9398 6400 9404 6452
rect 9456 6440 9462 6452
rect 10045 6443 10103 6449
rect 10045 6440 10057 6443
rect 9456 6412 10057 6440
rect 9456 6400 9462 6412
rect 10045 6409 10057 6412
rect 10091 6409 10103 6443
rect 10045 6403 10103 6409
rect 10318 6400 10324 6452
rect 10376 6400 10382 6452
rect 15838 6440 15844 6452
rect 10428 6412 15844 6440
rect 7558 6332 7564 6384
rect 7616 6372 7622 6384
rect 7616 6344 7972 6372
rect 7616 6332 7622 6344
rect 5445 6307 5503 6313
rect 5445 6273 5457 6307
rect 5491 6273 5503 6307
rect 5445 6267 5503 6273
rect 5460 6236 5488 6267
rect 6822 6264 6828 6316
rect 6880 6264 6886 6316
rect 7834 6264 7840 6316
rect 7892 6264 7898 6316
rect 7944 6304 7972 6344
rect 8113 6307 8171 6313
rect 8113 6304 8125 6307
rect 7944 6276 8125 6304
rect 8113 6273 8125 6276
rect 8159 6273 8171 6307
rect 8113 6267 8171 6273
rect 8205 6307 8263 6313
rect 8205 6273 8217 6307
rect 8251 6304 8263 6307
rect 8478 6304 8484 6316
rect 8251 6276 8484 6304
rect 8251 6273 8263 6276
rect 8205 6267 8263 6273
rect 8478 6264 8484 6276
rect 8536 6264 8542 6316
rect 8573 6307 8631 6313
rect 8573 6273 8585 6307
rect 8619 6304 8631 6307
rect 8846 6304 8852 6316
rect 8619 6276 8852 6304
rect 8619 6273 8631 6276
rect 8573 6267 8631 6273
rect 8846 6264 8852 6276
rect 8904 6264 8910 6316
rect 9125 6307 9183 6313
rect 9125 6273 9137 6307
rect 9171 6304 9183 6307
rect 9401 6307 9459 6313
rect 9401 6304 9413 6307
rect 9171 6276 9413 6304
rect 9171 6273 9183 6276
rect 9125 6267 9183 6273
rect 9401 6273 9413 6276
rect 9447 6304 9459 6307
rect 9582 6304 9588 6316
rect 9447 6276 9588 6304
rect 9447 6273 9459 6276
rect 9401 6267 9459 6273
rect 9582 6264 9588 6276
rect 9640 6264 9646 6316
rect 9677 6307 9735 6313
rect 9677 6273 9689 6307
rect 9723 6273 9735 6307
rect 9677 6267 9735 6273
rect 8938 6236 8944 6248
rect 5460 6208 8944 6236
rect 8938 6196 8944 6208
rect 8996 6196 9002 6248
rect 9692 6236 9720 6267
rect 9766 6264 9772 6316
rect 9824 6264 9830 6316
rect 10237 6311 10295 6317
rect 10237 6277 10249 6311
rect 10283 6308 10295 6311
rect 10283 6304 10364 6308
rect 10428 6304 10456 6412
rect 15838 6400 15844 6412
rect 15896 6400 15902 6452
rect 16298 6400 16304 6452
rect 16356 6440 16362 6452
rect 19794 6440 19800 6452
rect 16356 6412 19800 6440
rect 16356 6400 16362 6412
rect 19794 6400 19800 6412
rect 19852 6400 19858 6452
rect 19978 6400 19984 6452
rect 20036 6440 20042 6452
rect 23474 6440 23480 6452
rect 20036 6412 23480 6440
rect 20036 6400 20042 6412
rect 23474 6400 23480 6412
rect 23532 6400 23538 6452
rect 23658 6400 23664 6452
rect 23716 6440 23722 6452
rect 26418 6440 26424 6452
rect 23716 6412 26424 6440
rect 23716 6400 23722 6412
rect 26418 6400 26424 6412
rect 26476 6400 26482 6452
rect 28721 6443 28779 6449
rect 28721 6409 28733 6443
rect 28767 6440 28779 6443
rect 29086 6440 29092 6452
rect 28767 6412 29092 6440
rect 28767 6409 28779 6412
rect 28721 6403 28779 6409
rect 29086 6400 29092 6412
rect 29144 6400 29150 6452
rect 30558 6400 30564 6452
rect 30616 6440 30622 6452
rect 30837 6443 30895 6449
rect 30837 6440 30849 6443
rect 30616 6412 30849 6440
rect 30616 6400 30622 6412
rect 30837 6409 30849 6412
rect 30883 6409 30895 6443
rect 30837 6403 30895 6409
rect 31846 6400 31852 6452
rect 31904 6400 31910 6452
rect 10594 6332 10600 6384
rect 10652 6372 10658 6384
rect 12710 6372 12716 6384
rect 10652 6344 12716 6372
rect 10652 6332 10658 6344
rect 12710 6332 12716 6344
rect 12768 6332 12774 6384
rect 12802 6332 12808 6384
rect 12860 6372 12866 6384
rect 21358 6372 21364 6384
rect 12860 6344 21364 6372
rect 12860 6332 12866 6344
rect 21358 6332 21364 6344
rect 21416 6332 21422 6384
rect 21634 6332 21640 6384
rect 21692 6372 21698 6384
rect 30650 6372 30656 6384
rect 21692 6344 30656 6372
rect 21692 6332 21698 6344
rect 30650 6332 30656 6344
rect 30708 6332 30714 6384
rect 10505 6316 10563 6317
rect 10283 6280 10456 6304
rect 10283 6277 10295 6280
rect 10237 6271 10295 6277
rect 10336 6276 10456 6280
rect 10502 6264 10508 6316
rect 10560 6264 10566 6316
rect 10870 6264 10876 6316
rect 10928 6264 10934 6316
rect 11241 6307 11299 6313
rect 11241 6273 11253 6307
rect 11287 6304 11299 6307
rect 11790 6304 11796 6316
rect 11287 6276 11796 6304
rect 11287 6273 11299 6276
rect 11241 6267 11299 6273
rect 11790 6264 11796 6276
rect 11848 6264 11854 6316
rect 19610 6304 19616 6316
rect 12406 6276 19616 6304
rect 9950 6236 9956 6248
rect 9692 6208 9956 6236
rect 9950 6196 9956 6208
rect 10008 6196 10014 6248
rect 10410 6196 10416 6248
rect 10468 6236 10474 6248
rect 12406 6236 12434 6276
rect 19610 6264 19616 6276
rect 19668 6264 19674 6316
rect 21542 6264 21548 6316
rect 21600 6304 21606 6316
rect 22097 6307 22155 6313
rect 22097 6304 22109 6307
rect 21600 6276 22109 6304
rect 21600 6264 21606 6276
rect 22097 6273 22109 6276
rect 22143 6273 22155 6307
rect 22097 6267 22155 6273
rect 23290 6264 23296 6316
rect 23348 6304 23354 6316
rect 24302 6304 24308 6316
rect 23348 6276 24308 6304
rect 23348 6264 23354 6276
rect 24302 6264 24308 6276
rect 24360 6264 24366 6316
rect 24394 6264 24400 6316
rect 24452 6304 24458 6316
rect 27798 6304 27804 6316
rect 24452 6276 27804 6304
rect 24452 6264 24458 6276
rect 27798 6264 27804 6276
rect 27856 6264 27862 6316
rect 28537 6307 28595 6313
rect 28537 6273 28549 6307
rect 28583 6304 28595 6307
rect 30926 6304 30932 6316
rect 28583 6276 30932 6304
rect 28583 6273 28595 6276
rect 28537 6267 28595 6273
rect 30926 6264 30932 6276
rect 30984 6264 30990 6316
rect 31021 6307 31079 6313
rect 31021 6273 31033 6307
rect 31067 6273 31079 6307
rect 31021 6267 31079 6273
rect 10468 6208 12434 6236
rect 10468 6196 10474 6208
rect 19518 6196 19524 6248
rect 19576 6236 19582 6248
rect 30466 6236 30472 6248
rect 19576 6208 30472 6236
rect 19576 6196 19582 6208
rect 30466 6196 30472 6208
rect 30524 6196 30530 6248
rect 31036 6236 31064 6267
rect 31294 6264 31300 6316
rect 31352 6264 31358 6316
rect 31386 6264 31392 6316
rect 31444 6304 31450 6316
rect 31665 6307 31723 6313
rect 31665 6304 31677 6307
rect 31444 6276 31677 6304
rect 31444 6264 31450 6276
rect 31665 6273 31677 6276
rect 31711 6273 31723 6307
rect 31665 6267 31723 6273
rect 32490 6236 32496 6248
rect 31036 6208 32496 6236
rect 32490 6196 32496 6208
rect 32548 6196 32554 6248
rect 4706 6128 4712 6180
rect 4764 6168 4770 6180
rect 7929 6171 7987 6177
rect 7929 6168 7941 6171
rect 4764 6140 7941 6168
rect 4764 6128 4770 6140
rect 7929 6137 7941 6140
rect 7975 6137 7987 6171
rect 7929 6131 7987 6137
rect 8570 6128 8576 6180
rect 8628 6168 8634 6180
rect 9493 6171 9551 6177
rect 9493 6168 9505 6171
rect 8628 6140 9505 6168
rect 8628 6128 8634 6140
rect 9493 6137 9505 6140
rect 9539 6137 9551 6171
rect 9493 6131 9551 6137
rect 10689 6171 10747 6177
rect 10689 6137 10701 6171
rect 10735 6168 10747 6171
rect 10778 6168 10784 6180
rect 10735 6140 10784 6168
rect 10735 6137 10747 6140
rect 10689 6131 10747 6137
rect 10778 6128 10784 6140
rect 10836 6128 10842 6180
rect 12158 6168 12164 6180
rect 10888 6140 12164 6168
rect 6822 6060 6828 6112
rect 6880 6100 6886 6112
rect 9582 6100 9588 6112
rect 6880 6072 9588 6100
rect 6880 6060 6886 6072
rect 9582 6060 9588 6072
rect 9640 6060 9646 6112
rect 9953 6103 10011 6109
rect 9953 6069 9965 6103
rect 9999 6100 10011 6103
rect 10134 6100 10140 6112
rect 9999 6072 10140 6100
rect 9999 6069 10011 6072
rect 9953 6063 10011 6069
rect 10134 6060 10140 6072
rect 10192 6060 10198 6112
rect 10410 6060 10416 6112
rect 10468 6100 10474 6112
rect 10888 6100 10916 6140
rect 12158 6128 12164 6140
rect 12216 6128 12222 6180
rect 18414 6128 18420 6180
rect 18472 6168 18478 6180
rect 23198 6168 23204 6180
rect 18472 6140 23204 6168
rect 18472 6128 18478 6140
rect 23198 6128 23204 6140
rect 23256 6128 23262 6180
rect 23566 6128 23572 6180
rect 23624 6168 23630 6180
rect 28258 6168 28264 6180
rect 23624 6140 28264 6168
rect 23624 6128 23630 6140
rect 28258 6128 28264 6140
rect 28316 6128 28322 6180
rect 31478 6128 31484 6180
rect 31536 6128 31542 6180
rect 10468 6072 10916 6100
rect 10468 6060 10474 6072
rect 11054 6060 11060 6112
rect 11112 6060 11118 6112
rect 11146 6060 11152 6112
rect 11204 6100 11210 6112
rect 13630 6100 13636 6112
rect 11204 6072 13636 6100
rect 11204 6060 11210 6072
rect 13630 6060 13636 6072
rect 13688 6060 13694 6112
rect 15286 6060 15292 6112
rect 15344 6100 15350 6112
rect 17586 6100 17592 6112
rect 15344 6072 17592 6100
rect 15344 6060 15350 6072
rect 17586 6060 17592 6072
rect 17644 6060 17650 6112
rect 17678 6060 17684 6112
rect 17736 6100 17742 6112
rect 22186 6100 22192 6112
rect 17736 6072 22192 6100
rect 17736 6060 17742 6072
rect 22186 6060 22192 6072
rect 22244 6060 22250 6112
rect 22278 6060 22284 6112
rect 22336 6060 22342 6112
rect 23842 6060 23848 6112
rect 23900 6100 23906 6112
rect 28626 6100 28632 6112
rect 23900 6072 28632 6100
rect 23900 6060 23906 6072
rect 28626 6060 28632 6072
rect 28684 6060 28690 6112
rect 1104 6010 32568 6032
rect 1104 5958 1950 6010
rect 2002 5958 2014 6010
rect 2066 5958 2078 6010
rect 2130 5958 2142 6010
rect 2194 5958 2206 6010
rect 2258 5958 7950 6010
rect 8002 5958 8014 6010
rect 8066 5958 8078 6010
rect 8130 5958 8142 6010
rect 8194 5958 8206 6010
rect 8258 5958 13950 6010
rect 14002 5958 14014 6010
rect 14066 5958 14078 6010
rect 14130 5958 14142 6010
rect 14194 5958 14206 6010
rect 14258 5958 19950 6010
rect 20002 5958 20014 6010
rect 20066 5958 20078 6010
rect 20130 5958 20142 6010
rect 20194 5958 20206 6010
rect 20258 5958 25950 6010
rect 26002 5958 26014 6010
rect 26066 5958 26078 6010
rect 26130 5958 26142 6010
rect 26194 5958 26206 6010
rect 26258 5958 31950 6010
rect 32002 5958 32014 6010
rect 32066 5958 32078 6010
rect 32130 5958 32142 6010
rect 32194 5958 32206 6010
rect 32258 5958 32568 6010
rect 1104 5936 32568 5958
rect 6733 5899 6791 5905
rect 6733 5865 6745 5899
rect 6779 5896 6791 5899
rect 7190 5896 7196 5908
rect 6779 5868 7196 5896
rect 6779 5865 6791 5868
rect 6733 5859 6791 5865
rect 7190 5856 7196 5868
rect 7248 5856 7254 5908
rect 7374 5856 7380 5908
rect 7432 5856 7438 5908
rect 7653 5899 7711 5905
rect 7653 5865 7665 5899
rect 7699 5896 7711 5899
rect 7742 5896 7748 5908
rect 7699 5868 7748 5896
rect 7699 5865 7711 5868
rect 7653 5859 7711 5865
rect 7742 5856 7748 5868
rect 7800 5856 7806 5908
rect 7834 5856 7840 5908
rect 7892 5896 7898 5908
rect 7892 5868 8892 5896
rect 7892 5856 7898 5868
rect 8864 5828 8892 5868
rect 8938 5856 8944 5908
rect 8996 5896 9002 5908
rect 8996 5868 11376 5896
rect 8996 5856 9002 5868
rect 11348 5828 11376 5868
rect 11422 5856 11428 5908
rect 11480 5896 11486 5908
rect 15286 5896 15292 5908
rect 11480 5868 15292 5896
rect 11480 5856 11486 5868
rect 15286 5856 15292 5868
rect 15344 5856 15350 5908
rect 16758 5896 16764 5908
rect 15488 5868 16764 5896
rect 15488 5828 15516 5868
rect 16758 5856 16764 5868
rect 16816 5856 16822 5908
rect 17586 5856 17592 5908
rect 17644 5896 17650 5908
rect 20806 5896 20812 5908
rect 17644 5868 20812 5896
rect 17644 5856 17650 5868
rect 20806 5856 20812 5868
rect 20864 5856 20870 5908
rect 21358 5856 21364 5908
rect 21416 5896 21422 5908
rect 31294 5896 31300 5908
rect 21416 5868 31300 5896
rect 21416 5856 21422 5868
rect 31294 5856 31300 5868
rect 31352 5856 31358 5908
rect 16390 5828 16396 5840
rect 8864 5800 11284 5828
rect 11348 5800 15516 5828
rect 15672 5800 16396 5828
rect 11146 5760 11152 5772
rect 6564 5732 11152 5760
rect 6564 5701 6592 5732
rect 11146 5720 11152 5732
rect 11204 5720 11210 5772
rect 11256 5760 11284 5800
rect 15672 5760 15700 5800
rect 16390 5788 16396 5800
rect 16448 5788 16454 5840
rect 21637 5831 21695 5837
rect 21637 5797 21649 5831
rect 21683 5828 21695 5831
rect 21726 5828 21732 5840
rect 21683 5800 21732 5828
rect 21683 5797 21695 5800
rect 21637 5791 21695 5797
rect 21726 5788 21732 5800
rect 21784 5788 21790 5840
rect 22094 5828 22100 5840
rect 22066 5788 22100 5828
rect 22152 5788 22158 5840
rect 22278 5788 22284 5840
rect 22336 5828 22342 5840
rect 27522 5828 27528 5840
rect 22336 5800 27528 5828
rect 22336 5788 22342 5800
rect 27522 5788 27528 5800
rect 27580 5788 27586 5840
rect 31389 5831 31447 5837
rect 31389 5797 31401 5831
rect 31435 5828 31447 5831
rect 32030 5828 32036 5840
rect 31435 5800 32036 5828
rect 31435 5797 31447 5800
rect 31389 5791 31447 5797
rect 32030 5788 32036 5800
rect 32088 5788 32094 5840
rect 32122 5788 32128 5840
rect 32180 5788 32186 5840
rect 11256 5732 15700 5760
rect 15746 5720 15752 5772
rect 15804 5760 15810 5772
rect 22066 5760 22094 5788
rect 15804 5732 22094 5760
rect 15804 5720 15810 5732
rect 6549 5695 6607 5701
rect 6549 5661 6561 5695
rect 6595 5661 6607 5695
rect 6549 5655 6607 5661
rect 7006 5652 7012 5704
rect 7064 5692 7070 5704
rect 7193 5695 7251 5701
rect 7193 5692 7205 5695
rect 7064 5664 7205 5692
rect 7064 5652 7070 5664
rect 7193 5661 7205 5664
rect 7239 5661 7251 5695
rect 7193 5655 7251 5661
rect 7834 5652 7840 5704
rect 7892 5652 7898 5704
rect 9122 5652 9128 5704
rect 9180 5652 9186 5704
rect 13538 5692 13544 5704
rect 12406 5664 13544 5692
rect 9582 5584 9588 5636
rect 9640 5624 9646 5636
rect 12406 5624 12434 5664
rect 13538 5652 13544 5664
rect 13596 5652 13602 5704
rect 16206 5652 16212 5704
rect 16264 5692 16270 5704
rect 16393 5695 16451 5701
rect 16393 5692 16405 5695
rect 16264 5664 16405 5692
rect 16264 5652 16270 5664
rect 16393 5661 16405 5664
rect 16439 5661 16451 5695
rect 17126 5692 17132 5704
rect 16393 5655 16451 5661
rect 16500 5664 17132 5692
rect 9640 5596 12434 5624
rect 9640 5584 9646 5596
rect 6178 5516 6184 5568
rect 6236 5556 6242 5568
rect 8941 5559 8999 5565
rect 8941 5556 8953 5559
rect 6236 5528 8953 5556
rect 6236 5516 6242 5528
rect 8941 5525 8953 5528
rect 8987 5525 8999 5559
rect 8941 5519 8999 5525
rect 9674 5516 9680 5568
rect 9732 5556 9738 5568
rect 16500 5556 16528 5664
rect 17126 5652 17132 5664
rect 17184 5652 17190 5704
rect 20346 5652 20352 5704
rect 20404 5692 20410 5704
rect 21453 5695 21511 5701
rect 21453 5692 21465 5695
rect 20404 5664 21465 5692
rect 20404 5652 20410 5664
rect 21453 5661 21465 5664
rect 21499 5661 21511 5695
rect 21453 5655 21511 5661
rect 31202 5652 31208 5704
rect 31260 5652 31266 5704
rect 31294 5652 31300 5704
rect 31352 5692 31358 5704
rect 31573 5695 31631 5701
rect 31573 5692 31585 5695
rect 31352 5664 31585 5692
rect 31352 5652 31358 5664
rect 31573 5661 31585 5664
rect 31619 5661 31631 5695
rect 31573 5655 31631 5661
rect 31846 5652 31852 5704
rect 31904 5692 31910 5704
rect 31941 5695 31999 5701
rect 31941 5692 31953 5695
rect 31904 5664 31953 5692
rect 31904 5652 31910 5664
rect 31941 5661 31953 5664
rect 31987 5661 31999 5695
rect 31941 5655 31999 5661
rect 31662 5624 31668 5636
rect 16592 5596 31668 5624
rect 16592 5565 16620 5596
rect 31662 5584 31668 5596
rect 31720 5584 31726 5636
rect 9732 5528 16528 5556
rect 16577 5559 16635 5565
rect 9732 5516 9738 5528
rect 16577 5525 16589 5559
rect 16623 5525 16635 5559
rect 16577 5519 16635 5525
rect 31754 5516 31760 5568
rect 31812 5516 31818 5568
rect 1104 5466 32568 5488
rect 1104 5414 3010 5466
rect 3062 5414 3074 5466
rect 3126 5414 3138 5466
rect 3190 5414 3202 5466
rect 3254 5414 3266 5466
rect 3318 5414 9010 5466
rect 9062 5414 9074 5466
rect 9126 5414 9138 5466
rect 9190 5414 9202 5466
rect 9254 5414 9266 5466
rect 9318 5414 15010 5466
rect 15062 5414 15074 5466
rect 15126 5414 15138 5466
rect 15190 5414 15202 5466
rect 15254 5414 15266 5466
rect 15318 5414 21010 5466
rect 21062 5414 21074 5466
rect 21126 5414 21138 5466
rect 21190 5414 21202 5466
rect 21254 5414 21266 5466
rect 21318 5414 27010 5466
rect 27062 5414 27074 5466
rect 27126 5414 27138 5466
rect 27190 5414 27202 5466
rect 27254 5414 27266 5466
rect 27318 5414 32568 5466
rect 1104 5392 32568 5414
rect 7282 5312 7288 5364
rect 7340 5352 7346 5364
rect 8481 5355 8539 5361
rect 8481 5352 8493 5355
rect 7340 5324 8493 5352
rect 7340 5312 7346 5324
rect 8481 5321 8493 5324
rect 8527 5321 8539 5355
rect 8481 5315 8539 5321
rect 21450 5312 21456 5364
rect 21508 5312 21514 5364
rect 15378 5284 15384 5296
rect 8680 5256 15384 5284
rect 8680 5225 8708 5256
rect 15378 5244 15384 5256
rect 15436 5244 15442 5296
rect 19058 5244 19064 5296
rect 19116 5284 19122 5296
rect 19116 5256 26234 5284
rect 19116 5244 19122 5256
rect 8665 5219 8723 5225
rect 8665 5185 8677 5219
rect 8711 5185 8723 5219
rect 8665 5179 8723 5185
rect 9858 5176 9864 5228
rect 9916 5216 9922 5228
rect 15105 5219 15163 5225
rect 15105 5216 15117 5219
rect 9916 5188 15117 5216
rect 9916 5176 9922 5188
rect 15105 5185 15117 5188
rect 15151 5185 15163 5219
rect 15105 5179 15163 5185
rect 18414 5176 18420 5228
rect 18472 5216 18478 5228
rect 21269 5219 21327 5225
rect 21269 5216 21281 5219
rect 18472 5188 21281 5216
rect 18472 5176 18478 5188
rect 21269 5185 21281 5188
rect 21315 5185 21327 5219
rect 26206 5216 26234 5256
rect 31297 5219 31355 5225
rect 31297 5216 31309 5219
rect 26206 5188 31309 5216
rect 21269 5179 21327 5185
rect 31297 5185 31309 5188
rect 31343 5185 31355 5219
rect 31297 5179 31355 5185
rect 31662 5176 31668 5228
rect 31720 5176 31726 5228
rect 4614 5108 4620 5160
rect 4672 5148 4678 5160
rect 20898 5148 20904 5160
rect 4672 5120 20904 5148
rect 4672 5108 4678 5120
rect 20898 5108 20904 5120
rect 20956 5108 20962 5160
rect 15289 5083 15347 5089
rect 15289 5049 15301 5083
rect 15335 5080 15347 5083
rect 30374 5080 30380 5092
rect 15335 5052 30380 5080
rect 15335 5049 15347 5052
rect 15289 5043 15347 5049
rect 30374 5040 30380 5052
rect 30432 5040 30438 5092
rect 31478 4972 31484 5024
rect 31536 4972 31542 5024
rect 31849 5015 31907 5021
rect 31849 4981 31861 5015
rect 31895 5012 31907 5015
rect 32858 5012 32864 5024
rect 31895 4984 32864 5012
rect 31895 4981 31907 4984
rect 31849 4975 31907 4981
rect 32858 4972 32864 4984
rect 32916 4972 32922 5024
rect 1104 4922 32568 4944
rect 1104 4870 1950 4922
rect 2002 4870 2014 4922
rect 2066 4870 2078 4922
rect 2130 4870 2142 4922
rect 2194 4870 2206 4922
rect 2258 4870 7950 4922
rect 8002 4870 8014 4922
rect 8066 4870 8078 4922
rect 8130 4870 8142 4922
rect 8194 4870 8206 4922
rect 8258 4870 13950 4922
rect 14002 4870 14014 4922
rect 14066 4870 14078 4922
rect 14130 4870 14142 4922
rect 14194 4870 14206 4922
rect 14258 4870 19950 4922
rect 20002 4870 20014 4922
rect 20066 4870 20078 4922
rect 20130 4870 20142 4922
rect 20194 4870 20206 4922
rect 20258 4870 25950 4922
rect 26002 4870 26014 4922
rect 26066 4870 26078 4922
rect 26130 4870 26142 4922
rect 26194 4870 26206 4922
rect 26258 4870 31950 4922
rect 32002 4870 32014 4922
rect 32066 4870 32078 4922
rect 32130 4870 32142 4922
rect 32194 4870 32206 4922
rect 32258 4870 32568 4922
rect 1104 4848 32568 4870
rect 13814 4768 13820 4820
rect 13872 4808 13878 4820
rect 31386 4808 31392 4820
rect 13872 4780 31392 4808
rect 13872 4768 13878 4780
rect 31386 4768 31392 4780
rect 31444 4768 31450 4820
rect 15654 4700 15660 4752
rect 15712 4740 15718 4752
rect 31662 4740 31668 4752
rect 15712 4712 31668 4740
rect 15712 4700 15718 4712
rect 31662 4700 31668 4712
rect 31720 4700 31726 4752
rect 28718 4672 28724 4684
rect 22756 4644 28724 4672
rect 566 4564 572 4616
rect 624 4604 630 4616
rect 19521 4607 19579 4613
rect 19521 4604 19533 4607
rect 624 4576 19533 4604
rect 624 4564 630 4576
rect 19521 4573 19533 4576
rect 19567 4573 19579 4607
rect 22649 4607 22707 4613
rect 22649 4604 22661 4607
rect 19521 4567 19579 4573
rect 22066 4576 22661 4604
rect 16942 4496 16948 4548
rect 17000 4536 17006 4548
rect 22066 4536 22094 4576
rect 22649 4573 22661 4576
rect 22695 4573 22707 4607
rect 22649 4567 22707 4573
rect 17000 4508 22094 4536
rect 17000 4496 17006 4508
rect 19705 4471 19763 4477
rect 19705 4437 19717 4471
rect 19751 4468 19763 4471
rect 22756 4468 22784 4644
rect 28718 4632 28724 4644
rect 28776 4632 28782 4684
rect 23750 4564 23756 4616
rect 23808 4564 23814 4616
rect 28994 4564 29000 4616
rect 29052 4604 29058 4616
rect 31573 4607 31631 4613
rect 31573 4604 31585 4607
rect 29052 4576 31585 4604
rect 29052 4564 29058 4576
rect 31573 4573 31585 4576
rect 31619 4573 31631 4607
rect 31573 4567 31631 4573
rect 31938 4564 31944 4616
rect 31996 4564 32002 4616
rect 27706 4536 27712 4548
rect 22848 4508 27712 4536
rect 22848 4477 22876 4508
rect 27706 4496 27712 4508
rect 27764 4496 27770 4548
rect 19751 4440 22784 4468
rect 22833 4471 22891 4477
rect 19751 4437 19763 4440
rect 19705 4431 19763 4437
rect 22833 4437 22845 4471
rect 22879 4437 22891 4471
rect 22833 4431 22891 4437
rect 23937 4471 23995 4477
rect 23937 4437 23949 4471
rect 23983 4468 23995 4471
rect 24762 4468 24768 4480
rect 23983 4440 24768 4468
rect 23983 4437 23995 4440
rect 23937 4431 23995 4437
rect 24762 4428 24768 4440
rect 24820 4428 24826 4480
rect 31754 4428 31760 4480
rect 31812 4428 31818 4480
rect 32122 4428 32128 4480
rect 32180 4428 32186 4480
rect 1104 4378 32568 4400
rect 1104 4326 3010 4378
rect 3062 4326 3074 4378
rect 3126 4326 3138 4378
rect 3190 4326 3202 4378
rect 3254 4326 3266 4378
rect 3318 4326 9010 4378
rect 9062 4326 9074 4378
rect 9126 4326 9138 4378
rect 9190 4326 9202 4378
rect 9254 4326 9266 4378
rect 9318 4326 15010 4378
rect 15062 4326 15074 4378
rect 15126 4326 15138 4378
rect 15190 4326 15202 4378
rect 15254 4326 15266 4378
rect 15318 4326 21010 4378
rect 21062 4326 21074 4378
rect 21126 4326 21138 4378
rect 21190 4326 21202 4378
rect 21254 4326 21266 4378
rect 21318 4326 27010 4378
rect 27062 4326 27074 4378
rect 27126 4326 27138 4378
rect 27190 4326 27202 4378
rect 27254 4326 27266 4378
rect 27318 4326 32568 4378
rect 1104 4304 32568 4326
rect 19426 4224 19432 4276
rect 19484 4264 19490 4276
rect 31938 4264 31944 4276
rect 19484 4236 31944 4264
rect 19484 4224 19490 4236
rect 31938 4224 31944 4236
rect 31996 4224 32002 4276
rect 12434 4088 12440 4140
rect 12492 4128 12498 4140
rect 12529 4131 12587 4137
rect 12529 4128 12541 4131
rect 12492 4100 12541 4128
rect 12492 4088 12498 4100
rect 12529 4097 12541 4100
rect 12575 4097 12587 4131
rect 12529 4091 12587 4097
rect 17862 4088 17868 4140
rect 17920 4128 17926 4140
rect 19242 4128 19248 4140
rect 17920 4100 19248 4128
rect 17920 4088 17926 4100
rect 19242 4088 19248 4100
rect 19300 4088 19306 4140
rect 20898 4088 20904 4140
rect 20956 4088 20962 4140
rect 26878 4088 26884 4140
rect 26936 4128 26942 4140
rect 31297 4131 31355 4137
rect 31297 4128 31309 4131
rect 26936 4100 31309 4128
rect 26936 4088 26942 4100
rect 31297 4097 31309 4100
rect 31343 4097 31355 4131
rect 31297 4091 31355 4097
rect 31386 4088 31392 4140
rect 31444 4128 31450 4140
rect 31665 4131 31723 4137
rect 31665 4128 31677 4131
rect 31444 4100 31677 4128
rect 31444 4088 31450 4100
rect 31665 4097 31677 4100
rect 31711 4097 31723 4131
rect 31665 4091 31723 4097
rect 16390 4020 16396 4072
rect 16448 4060 16454 4072
rect 25498 4060 25504 4072
rect 16448 4032 25504 4060
rect 16448 4020 16454 4032
rect 25498 4020 25504 4032
rect 25556 4020 25562 4072
rect 7006 3952 7012 4004
rect 7064 3992 7070 4004
rect 31202 3992 31208 4004
rect 7064 3964 31208 3992
rect 7064 3952 7070 3964
rect 31202 3952 31208 3964
rect 31260 3952 31266 4004
rect 6914 3884 6920 3936
rect 6972 3924 6978 3936
rect 10686 3924 10692 3936
rect 6972 3896 10692 3924
rect 6972 3884 6978 3896
rect 10686 3884 10692 3896
rect 10744 3884 10750 3936
rect 12713 3927 12771 3933
rect 12713 3893 12725 3927
rect 12759 3924 12771 3927
rect 13814 3924 13820 3936
rect 12759 3896 13820 3924
rect 12759 3893 12771 3896
rect 12713 3887 12771 3893
rect 13814 3884 13820 3896
rect 13872 3884 13878 3936
rect 15930 3884 15936 3936
rect 15988 3924 15994 3936
rect 19794 3924 19800 3936
rect 15988 3896 19800 3924
rect 15988 3884 15994 3896
rect 19794 3884 19800 3896
rect 19852 3884 19858 3936
rect 21085 3927 21143 3933
rect 21085 3893 21097 3927
rect 21131 3924 21143 3927
rect 21358 3924 21364 3936
rect 21131 3896 21364 3924
rect 21131 3893 21143 3896
rect 21085 3887 21143 3893
rect 21358 3884 21364 3896
rect 21416 3884 21422 3936
rect 25498 3884 25504 3936
rect 25556 3924 25562 3936
rect 26510 3924 26516 3936
rect 25556 3896 26516 3924
rect 25556 3884 25562 3896
rect 26510 3884 26516 3896
rect 26568 3884 26574 3936
rect 31478 3884 31484 3936
rect 31536 3884 31542 3936
rect 31849 3927 31907 3933
rect 31849 3893 31861 3927
rect 31895 3924 31907 3927
rect 32858 3924 32864 3936
rect 31895 3896 32864 3924
rect 31895 3893 31907 3896
rect 31849 3887 31907 3893
rect 32858 3884 32864 3896
rect 32916 3884 32922 3936
rect 1104 3834 32568 3856
rect 1104 3782 1950 3834
rect 2002 3782 2014 3834
rect 2066 3782 2078 3834
rect 2130 3782 2142 3834
rect 2194 3782 2206 3834
rect 2258 3782 7950 3834
rect 8002 3782 8014 3834
rect 8066 3782 8078 3834
rect 8130 3782 8142 3834
rect 8194 3782 8206 3834
rect 8258 3782 13950 3834
rect 14002 3782 14014 3834
rect 14066 3782 14078 3834
rect 14130 3782 14142 3834
rect 14194 3782 14206 3834
rect 14258 3782 19950 3834
rect 20002 3782 20014 3834
rect 20066 3782 20078 3834
rect 20130 3782 20142 3834
rect 20194 3782 20206 3834
rect 20258 3782 25950 3834
rect 26002 3782 26014 3834
rect 26066 3782 26078 3834
rect 26130 3782 26142 3834
rect 26194 3782 26206 3834
rect 26258 3782 31950 3834
rect 32002 3782 32014 3834
rect 32066 3782 32078 3834
rect 32130 3782 32142 3834
rect 32194 3782 32206 3834
rect 32258 3782 32568 3834
rect 1104 3760 32568 3782
rect 6917 3723 6975 3729
rect 6917 3689 6929 3723
rect 6963 3720 6975 3723
rect 7006 3720 7012 3732
rect 6963 3692 7012 3720
rect 6963 3689 6975 3692
rect 6917 3683 6975 3689
rect 7006 3680 7012 3692
rect 7064 3680 7070 3732
rect 9582 3680 9588 3732
rect 9640 3720 9646 3732
rect 11793 3723 11851 3729
rect 11793 3720 11805 3723
rect 9640 3692 11805 3720
rect 9640 3680 9646 3692
rect 11793 3689 11805 3692
rect 11839 3689 11851 3723
rect 11793 3683 11851 3689
rect 14918 3680 14924 3732
rect 14976 3720 14982 3732
rect 15289 3723 15347 3729
rect 15289 3720 15301 3723
rect 14976 3692 15301 3720
rect 14976 3680 14982 3692
rect 15289 3689 15301 3692
rect 15335 3689 15347 3723
rect 15562 3720 15568 3732
rect 15289 3683 15347 3689
rect 15396 3692 15568 3720
rect 9398 3612 9404 3664
rect 9456 3652 9462 3664
rect 10229 3655 10287 3661
rect 10229 3652 10241 3655
rect 9456 3624 10241 3652
rect 9456 3612 9462 3624
rect 10229 3621 10241 3624
rect 10275 3621 10287 3655
rect 10229 3615 10287 3621
rect 10873 3655 10931 3661
rect 10873 3621 10885 3655
rect 10919 3652 10931 3655
rect 10919 3624 12434 3652
rect 10919 3621 10931 3624
rect 10873 3615 10931 3621
rect 1302 3544 1308 3596
rect 1360 3584 1366 3596
rect 1360 3556 6776 3584
rect 1360 3544 1366 3556
rect 1118 3476 1124 3528
rect 1176 3516 1182 3528
rect 6748 3525 6776 3556
rect 7466 3544 7472 3596
rect 7524 3584 7530 3596
rect 7524 3556 9444 3584
rect 7524 3544 7530 3556
rect 9416 3525 9444 3556
rect 9490 3544 9496 3596
rect 9548 3584 9554 3596
rect 11149 3587 11207 3593
rect 11149 3584 11161 3587
rect 9548 3556 11161 3584
rect 9548 3544 9554 3556
rect 11149 3553 11161 3556
rect 11195 3553 11207 3587
rect 12406 3584 12434 3624
rect 13722 3612 13728 3664
rect 13780 3652 13786 3664
rect 15013 3655 15071 3661
rect 15013 3652 15025 3655
rect 13780 3624 15025 3652
rect 13780 3612 13786 3624
rect 15013 3621 15025 3624
rect 15059 3652 15071 3655
rect 15396 3652 15424 3692
rect 15562 3680 15568 3692
rect 15620 3680 15626 3732
rect 15654 3680 15660 3732
rect 15712 3680 15718 3732
rect 15930 3680 15936 3732
rect 15988 3680 15994 3732
rect 16482 3680 16488 3732
rect 16540 3720 16546 3732
rect 17589 3723 17647 3729
rect 17589 3720 17601 3723
rect 16540 3692 17601 3720
rect 16540 3680 16546 3692
rect 17589 3689 17601 3692
rect 17635 3689 17647 3723
rect 17589 3683 17647 3689
rect 17954 3680 17960 3732
rect 18012 3680 18018 3732
rect 18138 3680 18144 3732
rect 18196 3720 18202 3732
rect 18874 3720 18880 3732
rect 18196 3692 18880 3720
rect 18196 3680 18202 3692
rect 18874 3680 18880 3692
rect 18932 3680 18938 3732
rect 19058 3680 19064 3732
rect 19116 3680 19122 3732
rect 19426 3680 19432 3732
rect 19484 3680 19490 3732
rect 19518 3680 19524 3732
rect 19576 3720 19582 3732
rect 19889 3723 19947 3729
rect 19889 3720 19901 3723
rect 19576 3692 19901 3720
rect 19576 3680 19582 3692
rect 19889 3689 19901 3692
rect 19935 3689 19947 3723
rect 19889 3683 19947 3689
rect 22005 3723 22063 3729
rect 22005 3689 22017 3723
rect 22051 3720 22063 3723
rect 24210 3720 24216 3732
rect 22051 3692 24216 3720
rect 22051 3689 22063 3692
rect 22005 3683 22063 3689
rect 24210 3680 24216 3692
rect 24268 3680 24274 3732
rect 25498 3680 25504 3732
rect 25556 3680 25562 3732
rect 25866 3680 25872 3732
rect 25924 3720 25930 3732
rect 26145 3723 26203 3729
rect 26145 3720 26157 3723
rect 25924 3692 26157 3720
rect 25924 3680 25930 3692
rect 26145 3689 26157 3692
rect 26191 3689 26203 3723
rect 26145 3683 26203 3689
rect 16761 3655 16819 3661
rect 15059 3624 15424 3652
rect 15488 3624 15884 3652
rect 15059 3621 15071 3624
rect 15013 3615 15071 3621
rect 15488 3584 15516 3624
rect 12406 3556 15516 3584
rect 15856 3584 15884 3624
rect 16761 3621 16773 3655
rect 16807 3652 16819 3655
rect 16807 3624 17356 3652
rect 16807 3621 16819 3624
rect 16761 3615 16819 3621
rect 15856 3556 17264 3584
rect 11149 3547 11207 3553
rect 4709 3519 4767 3525
rect 4709 3516 4721 3519
rect 1176 3488 4721 3516
rect 1176 3476 1182 3488
rect 4709 3485 4721 3488
rect 4755 3485 4767 3519
rect 4709 3479 4767 3485
rect 6733 3519 6791 3525
rect 6733 3485 6745 3519
rect 6779 3485 6791 3519
rect 6733 3479 6791 3485
rect 8205 3519 8263 3525
rect 8205 3485 8217 3519
rect 8251 3485 8263 3519
rect 8205 3479 8263 3485
rect 9401 3519 9459 3525
rect 9401 3485 9413 3519
rect 9447 3485 9459 3519
rect 9401 3479 9459 3485
rect 10321 3519 10379 3525
rect 10321 3485 10333 3519
rect 10367 3516 10379 3519
rect 10413 3519 10471 3525
rect 10413 3516 10425 3519
rect 10367 3488 10425 3516
rect 10367 3485 10379 3488
rect 10321 3479 10379 3485
rect 10413 3485 10425 3488
rect 10459 3485 10471 3519
rect 10413 3479 10471 3485
rect 1302 3408 1308 3460
rect 1360 3448 1366 3460
rect 8220 3448 8248 3479
rect 10686 3476 10692 3528
rect 10744 3476 10750 3528
rect 11241 3519 11299 3525
rect 11241 3485 11253 3519
rect 11287 3516 11299 3519
rect 11333 3519 11391 3525
rect 11333 3516 11345 3519
rect 11287 3488 11345 3516
rect 11287 3485 11299 3488
rect 11241 3479 11299 3485
rect 11333 3485 11345 3488
rect 11379 3485 11391 3519
rect 11333 3479 11391 3485
rect 11885 3519 11943 3525
rect 11885 3485 11897 3519
rect 11931 3516 11943 3519
rect 11977 3519 12035 3525
rect 11977 3516 11989 3519
rect 11931 3488 11989 3516
rect 11931 3485 11943 3488
rect 11885 3479 11943 3485
rect 11977 3485 11989 3488
rect 12023 3485 12035 3519
rect 11977 3479 12035 3485
rect 12066 3476 12072 3528
rect 12124 3516 12130 3528
rect 12253 3519 12311 3525
rect 12253 3516 12265 3519
rect 12124 3488 12265 3516
rect 12124 3476 12130 3488
rect 12253 3485 12265 3488
rect 12299 3516 12311 3519
rect 12529 3519 12587 3525
rect 12529 3516 12541 3519
rect 12299 3488 12541 3516
rect 12299 3485 12311 3488
rect 12253 3479 12311 3485
rect 12529 3485 12541 3488
rect 12575 3485 12587 3519
rect 12529 3479 12587 3485
rect 14550 3476 14556 3528
rect 14608 3476 14614 3528
rect 15381 3519 15439 3525
rect 15381 3485 15393 3519
rect 15427 3516 15439 3519
rect 15473 3519 15531 3525
rect 15473 3516 15485 3519
rect 15427 3488 15485 3516
rect 15427 3485 15439 3488
rect 15381 3479 15439 3485
rect 15473 3485 15485 3488
rect 15519 3485 15531 3519
rect 15473 3479 15531 3485
rect 15562 3476 15568 3528
rect 15620 3516 15626 3528
rect 15749 3519 15807 3525
rect 15749 3516 15761 3519
rect 15620 3488 15761 3516
rect 15620 3476 15626 3488
rect 15749 3485 15761 3488
rect 15795 3485 15807 3519
rect 16850 3516 16856 3528
rect 15749 3479 15807 3485
rect 16500 3488 16856 3516
rect 16390 3448 16396 3460
rect 1360 3420 8248 3448
rect 9600 3420 16396 3448
rect 1360 3408 1366 3420
rect 4890 3340 4896 3392
rect 4948 3340 4954 3392
rect 8386 3340 8392 3392
rect 8444 3340 8450 3392
rect 9600 3389 9628 3420
rect 16390 3408 16396 3420
rect 16448 3408 16454 3460
rect 9585 3383 9643 3389
rect 9585 3349 9597 3383
rect 9631 3349 9643 3383
rect 9585 3343 9643 3349
rect 10594 3340 10600 3392
rect 10652 3340 10658 3392
rect 11514 3340 11520 3392
rect 11572 3340 11578 3392
rect 12158 3340 12164 3392
rect 12216 3340 12222 3392
rect 12434 3340 12440 3392
rect 12492 3340 12498 3392
rect 14737 3383 14795 3389
rect 14737 3349 14749 3383
rect 14783 3380 14795 3383
rect 16500 3380 16528 3488
rect 16850 3476 16856 3488
rect 16908 3476 16914 3528
rect 16945 3519 17003 3525
rect 16945 3485 16957 3519
rect 16991 3516 17003 3519
rect 17037 3519 17095 3525
rect 17037 3516 17049 3519
rect 16991 3488 17049 3516
rect 16991 3485 17003 3488
rect 16945 3479 17003 3485
rect 17037 3485 17049 3488
rect 17083 3485 17095 3519
rect 17037 3479 17095 3485
rect 17236 3448 17264 3556
rect 17328 3525 17356 3624
rect 17402 3612 17408 3664
rect 17460 3652 17466 3664
rect 19705 3655 19763 3661
rect 17460 3624 18644 3652
rect 17460 3612 17466 3624
rect 17681 3587 17739 3593
rect 17681 3553 17693 3587
rect 17727 3584 17739 3587
rect 18616 3584 18644 3624
rect 19705 3621 19717 3655
rect 19751 3621 19763 3655
rect 19705 3615 19763 3621
rect 19720 3584 19748 3615
rect 19794 3612 19800 3664
rect 19852 3652 19858 3664
rect 31846 3652 31852 3664
rect 19852 3624 31852 3652
rect 19852 3612 19858 3624
rect 31846 3612 31852 3624
rect 31904 3612 31910 3664
rect 28994 3584 29000 3596
rect 17727 3556 18368 3584
rect 17727 3553 17739 3556
rect 17681 3547 17739 3553
rect 17313 3519 17371 3525
rect 17313 3485 17325 3519
rect 17359 3485 17371 3519
rect 17313 3479 17371 3485
rect 17770 3476 17776 3528
rect 17828 3476 17834 3528
rect 18340 3525 18368 3556
rect 18616 3556 19656 3584
rect 19720 3556 29000 3584
rect 18616 3525 18644 3556
rect 18325 3519 18383 3525
rect 18325 3485 18337 3519
rect 18371 3485 18383 3519
rect 18325 3479 18383 3485
rect 18601 3519 18659 3525
rect 18601 3485 18613 3519
rect 18647 3485 18659 3519
rect 18601 3479 18659 3485
rect 18874 3476 18880 3528
rect 18932 3476 18938 3528
rect 19242 3476 19248 3528
rect 19300 3476 19306 3528
rect 19518 3476 19524 3528
rect 19576 3476 19582 3528
rect 19628 3516 19656 3556
rect 28994 3544 29000 3556
rect 29052 3544 29058 3596
rect 20165 3519 20223 3525
rect 20165 3516 20177 3519
rect 19628 3488 20177 3516
rect 20165 3485 20177 3488
rect 20211 3485 20223 3519
rect 20165 3479 20223 3485
rect 21818 3476 21824 3528
rect 21876 3476 21882 3528
rect 22186 3476 22192 3528
rect 22244 3476 22250 3528
rect 22462 3476 22468 3528
rect 22520 3476 22526 3528
rect 23474 3476 23480 3528
rect 23532 3516 23538 3528
rect 25317 3519 25375 3525
rect 25317 3516 25329 3519
rect 23532 3488 25329 3516
rect 23532 3476 23538 3488
rect 25317 3485 25329 3488
rect 25363 3485 25375 3519
rect 25317 3479 25375 3485
rect 25590 3476 25596 3528
rect 25648 3476 25654 3528
rect 25682 3476 25688 3528
rect 25740 3516 25746 3528
rect 25961 3519 26019 3525
rect 25961 3516 25973 3519
rect 25740 3488 25973 3516
rect 25740 3476 25746 3488
rect 25961 3485 25973 3488
rect 26007 3485 26019 3519
rect 25961 3479 26019 3485
rect 31570 3476 31576 3528
rect 31628 3476 31634 3528
rect 31938 3476 31944 3528
rect 31996 3476 32002 3528
rect 31294 3448 31300 3460
rect 17236 3420 31300 3448
rect 31294 3408 31300 3420
rect 31352 3408 31358 3460
rect 14783 3352 16528 3380
rect 14783 3349 14795 3352
rect 14737 3343 14795 3349
rect 16574 3340 16580 3392
rect 16632 3340 16638 3392
rect 16666 3340 16672 3392
rect 16724 3340 16730 3392
rect 16850 3340 16856 3392
rect 16908 3340 16914 3392
rect 17218 3340 17224 3392
rect 17276 3340 17282 3392
rect 17494 3340 17500 3392
rect 17552 3340 17558 3392
rect 18506 3340 18512 3392
rect 18564 3340 18570 3392
rect 18782 3340 18788 3392
rect 18840 3340 18846 3392
rect 19242 3340 19248 3392
rect 19300 3380 19306 3392
rect 19981 3383 20039 3389
rect 19981 3380 19993 3383
rect 19300 3352 19993 3380
rect 19300 3340 19306 3352
rect 19981 3349 19993 3352
rect 20027 3349 20039 3383
rect 19981 3343 20039 3349
rect 22370 3340 22376 3392
rect 22428 3340 22434 3392
rect 22649 3383 22707 3389
rect 22649 3349 22661 3383
rect 22695 3380 22707 3383
rect 23382 3380 23388 3392
rect 22695 3352 23388 3380
rect 22695 3349 22707 3352
rect 22649 3343 22707 3349
rect 23382 3340 23388 3352
rect 23440 3340 23446 3392
rect 25777 3383 25835 3389
rect 25777 3349 25789 3383
rect 25823 3380 25835 3383
rect 26326 3380 26332 3392
rect 25823 3352 26332 3380
rect 25823 3349 25835 3352
rect 25777 3343 25835 3349
rect 26326 3340 26332 3352
rect 26384 3340 26390 3392
rect 31754 3340 31760 3392
rect 31812 3340 31818 3392
rect 32122 3340 32128 3392
rect 32180 3340 32186 3392
rect 1104 3290 32568 3312
rect 1104 3238 3010 3290
rect 3062 3238 3074 3290
rect 3126 3238 3138 3290
rect 3190 3238 3202 3290
rect 3254 3238 3266 3290
rect 3318 3238 9010 3290
rect 9062 3238 9074 3290
rect 9126 3238 9138 3290
rect 9190 3238 9202 3290
rect 9254 3238 9266 3290
rect 9318 3238 15010 3290
rect 15062 3238 15074 3290
rect 15126 3238 15138 3290
rect 15190 3238 15202 3290
rect 15254 3238 15266 3290
rect 15318 3238 21010 3290
rect 21062 3238 21074 3290
rect 21126 3238 21138 3290
rect 21190 3238 21202 3290
rect 21254 3238 21266 3290
rect 21318 3238 27010 3290
rect 27062 3238 27074 3290
rect 27126 3238 27138 3290
rect 27190 3238 27202 3290
rect 27254 3238 27266 3290
rect 27318 3238 32568 3290
rect 1104 3216 32568 3238
rect 4338 3136 4344 3188
rect 4396 3176 4402 3188
rect 14550 3176 14556 3188
rect 4396 3148 14556 3176
rect 4396 3136 4402 3148
rect 14550 3136 14556 3148
rect 14608 3136 14614 3188
rect 17494 3136 17500 3188
rect 17552 3176 17558 3188
rect 31938 3176 31944 3188
rect 17552 3148 31944 3176
rect 17552 3136 17558 3148
rect 31938 3136 31944 3148
rect 31996 3136 32002 3188
rect 9398 3068 9404 3120
rect 9456 3108 9462 3120
rect 12066 3108 12072 3120
rect 9456 3080 12072 3108
rect 9456 3068 9462 3080
rect 12066 3068 12072 3080
rect 12124 3068 12130 3120
rect 17218 3068 17224 3120
rect 17276 3108 17282 3120
rect 31570 3108 31576 3120
rect 17276 3080 31576 3108
rect 17276 3068 17282 3080
rect 31570 3068 31576 3080
rect 31628 3068 31634 3120
rect 5902 3000 5908 3052
rect 5960 3040 5966 3052
rect 16574 3040 16580 3052
rect 5960 3012 16580 3040
rect 5960 3000 5966 3012
rect 16574 3000 16580 3012
rect 16632 3040 16638 3052
rect 17770 3040 17776 3052
rect 16632 3012 17776 3040
rect 16632 3000 16638 3012
rect 17770 3000 17776 3012
rect 17828 3000 17834 3052
rect 18782 3000 18788 3052
rect 18840 3040 18846 3052
rect 26878 3040 26884 3052
rect 18840 3012 26884 3040
rect 18840 3000 18846 3012
rect 26878 3000 26884 3012
rect 26936 3000 26942 3052
rect 30374 3000 30380 3052
rect 30432 3040 30438 3052
rect 31297 3043 31355 3049
rect 31297 3040 31309 3043
rect 30432 3012 31309 3040
rect 30432 3000 30438 3012
rect 31297 3009 31309 3012
rect 31343 3009 31355 3043
rect 31297 3003 31355 3009
rect 31662 3000 31668 3052
rect 31720 3000 31726 3052
rect 10594 2864 10600 2916
rect 10652 2904 10658 2916
rect 31386 2904 31392 2916
rect 10652 2876 31392 2904
rect 10652 2864 10658 2876
rect 31386 2864 31392 2876
rect 31444 2864 31450 2916
rect 31481 2839 31539 2845
rect 31481 2805 31493 2839
rect 31527 2836 31539 2839
rect 31754 2836 31760 2848
rect 31527 2808 31760 2836
rect 31527 2805 31539 2808
rect 31481 2799 31539 2805
rect 31754 2796 31760 2808
rect 31812 2796 31818 2848
rect 31849 2839 31907 2845
rect 31849 2805 31861 2839
rect 31895 2836 31907 2839
rect 32858 2836 32864 2848
rect 31895 2808 32864 2836
rect 31895 2805 31907 2808
rect 31849 2799 31907 2805
rect 32858 2796 32864 2808
rect 32916 2796 32922 2848
rect 1104 2746 32568 2768
rect 1104 2694 1950 2746
rect 2002 2694 2014 2746
rect 2066 2694 2078 2746
rect 2130 2694 2142 2746
rect 2194 2694 2206 2746
rect 2258 2694 7950 2746
rect 8002 2694 8014 2746
rect 8066 2694 8078 2746
rect 8130 2694 8142 2746
rect 8194 2694 8206 2746
rect 8258 2694 13950 2746
rect 14002 2694 14014 2746
rect 14066 2694 14078 2746
rect 14130 2694 14142 2746
rect 14194 2694 14206 2746
rect 14258 2694 19950 2746
rect 20002 2694 20014 2746
rect 20066 2694 20078 2746
rect 20130 2694 20142 2746
rect 20194 2694 20206 2746
rect 20258 2694 25950 2746
rect 26002 2694 26014 2746
rect 26066 2694 26078 2746
rect 26130 2694 26142 2746
rect 26194 2694 26206 2746
rect 26258 2694 31950 2746
rect 32002 2694 32014 2746
rect 32066 2694 32078 2746
rect 32130 2694 32142 2746
rect 32194 2694 32206 2746
rect 32258 2694 32568 2746
rect 1104 2672 32568 2694
rect 12434 2592 12440 2644
rect 12492 2632 12498 2644
rect 12492 2604 31708 2632
rect 12492 2592 12498 2604
rect 12158 2524 12164 2576
rect 12216 2564 12222 2576
rect 12216 2536 30604 2564
rect 12216 2524 12222 2536
rect 11514 2456 11520 2508
rect 11572 2496 11578 2508
rect 30466 2496 30472 2508
rect 11572 2468 30472 2496
rect 11572 2456 11578 2468
rect 30466 2456 30472 2468
rect 30524 2456 30530 2508
rect 4890 2388 4896 2440
rect 4948 2428 4954 2440
rect 30576 2437 30604 2536
rect 30561 2431 30619 2437
rect 4948 2400 26740 2428
rect 4948 2388 4954 2400
rect 8386 2320 8392 2372
rect 8444 2360 8450 2372
rect 26712 2360 26740 2400
rect 30561 2397 30573 2431
rect 30607 2397 30619 2431
rect 30561 2391 30619 2397
rect 30834 2388 30840 2440
rect 30892 2428 30898 2440
rect 31680 2437 31708 2604
rect 30929 2431 30987 2437
rect 30929 2428 30941 2431
rect 30892 2400 30941 2428
rect 30892 2388 30898 2400
rect 30929 2397 30941 2400
rect 30975 2397 30987 2431
rect 30929 2391 30987 2397
rect 31297 2431 31355 2437
rect 31297 2397 31309 2431
rect 31343 2397 31355 2431
rect 31297 2391 31355 2397
rect 31665 2431 31723 2437
rect 31665 2397 31677 2431
rect 31711 2397 31723 2431
rect 31665 2391 31723 2397
rect 31312 2360 31340 2391
rect 8444 2332 22094 2360
rect 26712 2332 31340 2360
rect 8444 2320 8450 2332
rect 22066 2292 22094 2332
rect 30374 2292 30380 2304
rect 22066 2264 30380 2292
rect 30374 2252 30380 2264
rect 30432 2252 30438 2304
rect 30742 2252 30748 2304
rect 30800 2252 30806 2304
rect 31110 2252 31116 2304
rect 31168 2252 31174 2304
rect 31478 2252 31484 2304
rect 31536 2252 31542 2304
rect 31846 2252 31852 2304
rect 31904 2252 31910 2304
rect 1104 2202 32568 2224
rect 1104 2150 3010 2202
rect 3062 2150 3074 2202
rect 3126 2150 3138 2202
rect 3190 2150 3202 2202
rect 3254 2150 3266 2202
rect 3318 2150 9010 2202
rect 9062 2150 9074 2202
rect 9126 2150 9138 2202
rect 9190 2150 9202 2202
rect 9254 2150 9266 2202
rect 9318 2150 15010 2202
rect 15062 2150 15074 2202
rect 15126 2150 15138 2202
rect 15190 2150 15202 2202
rect 15254 2150 15266 2202
rect 15318 2150 21010 2202
rect 21062 2150 21074 2202
rect 21126 2150 21138 2202
rect 21190 2150 21202 2202
rect 21254 2150 21266 2202
rect 21318 2150 27010 2202
rect 27062 2150 27074 2202
rect 27126 2150 27138 2202
rect 27190 2150 27202 2202
rect 27254 2150 27266 2202
rect 27318 2150 32568 2202
rect 1104 2128 32568 2150
rect 12158 2048 12164 2100
rect 12216 2088 12222 2100
rect 25682 2088 25688 2100
rect 12216 2060 25688 2088
rect 12216 2048 12222 2060
rect 25682 2048 25688 2060
rect 25740 2048 25746 2100
rect 2774 144 2780 196
rect 2832 144 2838 196
rect 2792 116 2820 144
rect 22186 116 22192 128
rect 2792 88 22192 116
rect 22186 76 22192 88
rect 22244 76 22250 128
rect 1302 8 1308 60
rect 1360 48 1366 60
rect 21818 48 21824 60
rect 1360 20 21824 48
rect 1360 8 1366 20
rect 21818 8 21824 20
rect 21876 8 21882 60
<< via1 >>
rect 15660 11092 15712 11144
rect 22100 11092 22152 11144
rect 13636 10004 13688 10056
rect 19340 10004 19392 10056
rect 25688 9596 25740 9648
rect 26148 9596 26200 9648
rect 7656 9392 7708 9444
rect 18788 9392 18840 9444
rect 8392 9256 8444 9308
rect 12532 9256 12584 9308
rect 12808 9256 12860 9308
rect 20996 9256 21048 9308
rect 10324 9188 10376 9240
rect 17960 9188 18012 9240
rect 9864 9120 9916 9172
rect 19248 9120 19300 9172
rect 10416 9052 10468 9104
rect 18236 9052 18288 9104
rect 23480 9052 23532 9104
rect 23756 9052 23808 9104
rect 27620 9052 27672 9104
rect 28632 9052 28684 9104
rect 10600 8984 10652 9036
rect 14096 8984 14148 9036
rect 21732 8984 21784 9036
rect 28080 8984 28132 9036
rect 13728 8916 13780 8968
rect 26884 8916 26936 8968
rect 27528 8916 27580 8968
rect 31668 8916 31720 8968
rect 10968 8848 11020 8900
rect 15568 8848 15620 8900
rect 17960 8848 18012 8900
rect 25044 8848 25096 8900
rect 26700 8848 26752 8900
rect 29920 8848 29972 8900
rect 11428 8780 11480 8832
rect 13452 8780 13504 8832
rect 21272 8780 21324 8832
rect 21548 8780 21600 8832
rect 23664 8780 23716 8832
rect 28816 8780 28868 8832
rect 3010 8678 3062 8730
rect 3074 8678 3126 8730
rect 3138 8678 3190 8730
rect 3202 8678 3254 8730
rect 3266 8678 3318 8730
rect 9010 8678 9062 8730
rect 9074 8678 9126 8730
rect 9138 8678 9190 8730
rect 9202 8678 9254 8730
rect 9266 8678 9318 8730
rect 15010 8678 15062 8730
rect 15074 8678 15126 8730
rect 15138 8678 15190 8730
rect 15202 8678 15254 8730
rect 15266 8678 15318 8730
rect 21010 8678 21062 8730
rect 21074 8678 21126 8730
rect 21138 8678 21190 8730
rect 21202 8678 21254 8730
rect 21266 8678 21318 8730
rect 27010 8678 27062 8730
rect 27074 8678 27126 8730
rect 27138 8678 27190 8730
rect 27202 8678 27254 8730
rect 27266 8678 27318 8730
rect 4436 8576 4488 8628
rect 4712 8576 4764 8628
rect 4988 8576 5040 8628
rect 5540 8576 5592 8628
rect 5816 8576 5868 8628
rect 6368 8576 6420 8628
rect 6920 8576 6972 8628
rect 7196 8576 7248 8628
rect 7748 8576 7800 8628
rect 8024 8576 8076 8628
rect 8484 8576 8536 8628
rect 8760 8576 8812 8628
rect 9404 8576 9456 8628
rect 9956 8576 10008 8628
rect 10232 8576 10284 8628
rect 10508 8576 10560 8628
rect 11060 8576 11112 8628
rect 11612 8576 11664 8628
rect 12164 8576 12216 8628
rect 12440 8576 12492 8628
rect 12716 8619 12768 8628
rect 12716 8585 12725 8619
rect 12725 8585 12759 8619
rect 12759 8585 12768 8619
rect 12716 8576 12768 8585
rect 12992 8576 13044 8628
rect 13268 8576 13320 8628
rect 13544 8576 13596 8628
rect 13912 8576 13964 8628
rect 24032 8619 24084 8628
rect 24032 8585 24041 8619
rect 24041 8585 24075 8619
rect 24075 8585 24084 8619
rect 24032 8576 24084 8585
rect 4344 8483 4396 8492
rect 4344 8449 4353 8483
rect 4353 8449 4387 8483
rect 4387 8449 4396 8483
rect 4344 8440 4396 8449
rect 4712 8483 4764 8492
rect 4712 8449 4721 8483
rect 4721 8449 4755 8483
rect 4755 8449 4764 8483
rect 4712 8440 4764 8449
rect 5172 8483 5224 8492
rect 5172 8449 5181 8483
rect 5181 8449 5215 8483
rect 5215 8449 5224 8483
rect 5172 8440 5224 8449
rect 5816 8483 5868 8492
rect 5816 8449 5825 8483
rect 5825 8449 5859 8483
rect 5859 8449 5868 8483
rect 5816 8440 5868 8449
rect 6184 8483 6236 8492
rect 6184 8449 6193 8483
rect 6193 8449 6227 8483
rect 6227 8449 6236 8483
rect 6184 8440 6236 8449
rect 7104 8440 7156 8492
rect 7288 8483 7340 8492
rect 7288 8449 7297 8483
rect 7297 8449 7331 8483
rect 7331 8449 7340 8483
rect 7288 8440 7340 8449
rect 7380 8483 7432 8492
rect 7380 8449 7389 8483
rect 7389 8449 7423 8483
rect 7423 8449 7432 8483
rect 7380 8440 7432 8449
rect 7748 8483 7800 8492
rect 7748 8449 7757 8483
rect 7757 8449 7791 8483
rect 7791 8449 7800 8483
rect 7748 8440 7800 8449
rect 8668 8440 8720 8492
rect 10692 8508 10744 8560
rect 11244 8508 11296 8560
rect 8576 8372 8628 8424
rect 9864 8483 9916 8492
rect 9864 8449 9873 8483
rect 9873 8449 9907 8483
rect 9907 8449 9916 8483
rect 9864 8440 9916 8449
rect 10416 8440 10468 8492
rect 10232 8304 10284 8356
rect 10968 8483 11020 8492
rect 10968 8449 10977 8483
rect 10977 8449 11011 8483
rect 11011 8449 11020 8483
rect 10968 8440 11020 8449
rect 11428 8440 11480 8492
rect 11520 8440 11572 8492
rect 12164 8483 12216 8492
rect 12164 8449 12173 8483
rect 12173 8449 12207 8483
rect 12207 8449 12216 8483
rect 12164 8440 12216 8449
rect 12532 8483 12584 8492
rect 12532 8449 12541 8483
rect 12541 8449 12575 8483
rect 12575 8449 12584 8483
rect 12532 8440 12584 8449
rect 16948 8508 17000 8560
rect 24400 8576 24452 8628
rect 24676 8576 24728 8628
rect 25044 8576 25096 8628
rect 25136 8576 25188 8628
rect 26240 8576 26292 8628
rect 27436 8576 27488 8628
rect 28632 8619 28684 8628
rect 28632 8585 28641 8619
rect 28641 8585 28675 8619
rect 28675 8585 28684 8619
rect 28632 8576 28684 8585
rect 11980 8372 12032 8424
rect 13360 8440 13412 8492
rect 14096 8483 14148 8492
rect 14096 8449 14105 8483
rect 14105 8449 14139 8483
rect 14139 8449 14148 8483
rect 14096 8440 14148 8449
rect 24216 8487 24268 8496
rect 24216 8453 24225 8487
rect 24225 8453 24259 8487
rect 24259 8453 24268 8487
rect 24216 8444 24268 8453
rect 25228 8508 25280 8560
rect 13544 8372 13596 8424
rect 16580 8372 16632 8424
rect 22376 8372 22428 8424
rect 25504 8483 25556 8492
rect 25504 8449 25513 8483
rect 25513 8449 25547 8483
rect 25547 8449 25556 8483
rect 25504 8440 25556 8449
rect 26792 8508 26844 8560
rect 26332 8440 26384 8492
rect 26516 8440 26568 8492
rect 27712 8483 27764 8492
rect 27712 8449 27721 8483
rect 27721 8449 27755 8483
rect 27755 8449 27764 8483
rect 27712 8440 27764 8449
rect 17500 8304 17552 8356
rect 23388 8304 23440 8356
rect 9956 8236 10008 8288
rect 14004 8236 14056 8288
rect 25044 8304 25096 8356
rect 25412 8304 25464 8356
rect 26148 8304 26200 8356
rect 26608 8304 26660 8356
rect 27988 8508 28040 8560
rect 29552 8576 29604 8628
rect 31116 8619 31168 8628
rect 31116 8585 31125 8619
rect 31125 8585 31159 8619
rect 31159 8585 31168 8619
rect 31116 8576 31168 8585
rect 28080 8483 28132 8492
rect 28080 8449 28089 8483
rect 28089 8449 28123 8483
rect 28123 8449 28132 8483
rect 28080 8440 28132 8449
rect 28816 8483 28868 8492
rect 28816 8449 28825 8483
rect 28825 8449 28859 8483
rect 28859 8449 28868 8483
rect 28816 8440 28868 8449
rect 28908 8440 28960 8492
rect 29552 8483 29604 8492
rect 29552 8449 29561 8483
rect 29561 8449 29595 8483
rect 29595 8449 29604 8483
rect 29552 8440 29604 8449
rect 29920 8483 29972 8492
rect 29920 8449 29929 8483
rect 29929 8449 29963 8483
rect 29963 8449 29972 8483
rect 29920 8440 29972 8449
rect 30564 8483 30616 8492
rect 30564 8449 30573 8483
rect 30573 8449 30607 8483
rect 30607 8449 30616 8483
rect 30564 8440 30616 8449
rect 31300 8483 31352 8492
rect 31300 8449 31309 8483
rect 31309 8449 31343 8483
rect 31343 8449 31352 8483
rect 31300 8440 31352 8449
rect 31668 8483 31720 8492
rect 31668 8449 31677 8483
rect 31677 8449 31711 8483
rect 31711 8449 31720 8483
rect 31668 8440 31720 8449
rect 27620 8236 27672 8288
rect 29000 8372 29052 8424
rect 28724 8304 28776 8356
rect 32588 8304 32640 8356
rect 31852 8279 31904 8288
rect 31852 8245 31861 8279
rect 31861 8245 31895 8279
rect 31895 8245 31904 8279
rect 31852 8236 31904 8245
rect 1950 8134 2002 8186
rect 2014 8134 2066 8186
rect 2078 8134 2130 8186
rect 2142 8134 2194 8186
rect 2206 8134 2258 8186
rect 7950 8134 8002 8186
rect 8014 8134 8066 8186
rect 8078 8134 8130 8186
rect 8142 8134 8194 8186
rect 8206 8134 8258 8186
rect 13950 8134 14002 8186
rect 14014 8134 14066 8186
rect 14078 8134 14130 8186
rect 14142 8134 14194 8186
rect 14206 8134 14258 8186
rect 19950 8134 20002 8186
rect 20014 8134 20066 8186
rect 20078 8134 20130 8186
rect 20142 8134 20194 8186
rect 20206 8134 20258 8186
rect 25950 8134 26002 8186
rect 26014 8134 26066 8186
rect 26078 8134 26130 8186
rect 26142 8134 26194 8186
rect 26206 8134 26258 8186
rect 31950 8134 32002 8186
rect 32014 8134 32066 8186
rect 32078 8134 32130 8186
rect 32142 8134 32194 8186
rect 32206 8134 32258 8186
rect 4160 8032 4212 8084
rect 5264 8032 5316 8084
rect 6092 8032 6144 8084
rect 6644 8032 6696 8084
rect 7472 8032 7524 8084
rect 8300 8032 8352 8084
rect 8852 8032 8904 8084
rect 9680 8032 9732 8084
rect 10784 8032 10836 8084
rect 11336 8032 11388 8084
rect 11888 8032 11940 8084
rect 25872 8032 25924 8084
rect 27344 8075 27396 8084
rect 27344 8041 27353 8075
rect 27353 8041 27387 8075
rect 27387 8041 27396 8075
rect 27344 8032 27396 8041
rect 28172 8032 28224 8084
rect 28540 8032 28592 8084
rect 29276 8032 29328 8084
rect 30656 8075 30708 8084
rect 30656 8041 30665 8075
rect 30665 8041 30699 8075
rect 30699 8041 30708 8075
rect 30656 8032 30708 8041
rect 31024 8075 31076 8084
rect 31024 8041 31033 8075
rect 31033 8041 31067 8075
rect 31067 8041 31076 8075
rect 31024 8032 31076 8041
rect 31392 8075 31444 8084
rect 31392 8041 31401 8075
rect 31401 8041 31435 8075
rect 31435 8041 31444 8075
rect 31392 8032 31444 8041
rect 10048 7964 10100 8016
rect 19340 7964 19392 8016
rect 8484 7896 8536 7948
rect 20812 7896 20864 7948
rect 27620 7896 27672 7948
rect 5356 7871 5408 7880
rect 5356 7837 5365 7871
rect 5365 7837 5399 7871
rect 5399 7837 5408 7871
rect 5356 7828 5408 7837
rect 6920 7828 6972 7880
rect 6276 7760 6328 7812
rect 7196 7828 7248 7880
rect 8668 7871 8720 7880
rect 8668 7837 8677 7871
rect 8677 7837 8711 7871
rect 8711 7837 8720 7871
rect 8668 7828 8720 7837
rect 9496 7871 9548 7880
rect 9496 7837 9505 7871
rect 9505 7837 9539 7871
rect 9539 7837 9548 7871
rect 9496 7828 9548 7837
rect 10048 7871 10100 7880
rect 10048 7837 10057 7871
rect 10057 7837 10091 7871
rect 10091 7837 10100 7871
rect 10048 7828 10100 7837
rect 9404 7760 9456 7812
rect 12624 7828 12676 7880
rect 25872 7828 25924 7880
rect 14372 7760 14424 7812
rect 21456 7760 21508 7812
rect 28264 7871 28316 7880
rect 28264 7837 28273 7871
rect 28273 7837 28307 7871
rect 28307 7837 28316 7871
rect 28264 7828 28316 7837
rect 28632 7871 28684 7880
rect 28632 7837 28641 7871
rect 28641 7837 28675 7871
rect 28675 7837 28684 7871
rect 28632 7828 28684 7837
rect 29092 7828 29144 7880
rect 30472 7871 30524 7880
rect 30472 7837 30481 7871
rect 30481 7837 30515 7871
rect 30515 7837 30524 7871
rect 30472 7828 30524 7837
rect 30656 7828 30708 7880
rect 30932 7828 30984 7880
rect 29000 7760 29052 7812
rect 16488 7692 16540 7744
rect 26240 7692 26292 7744
rect 31300 7692 31352 7744
rect 31760 7735 31812 7744
rect 31760 7701 31769 7735
rect 31769 7701 31803 7735
rect 31803 7701 31812 7735
rect 31760 7692 31812 7701
rect 32128 7735 32180 7744
rect 32128 7701 32137 7735
rect 32137 7701 32171 7735
rect 32171 7701 32180 7735
rect 32128 7692 32180 7701
rect 3010 7590 3062 7642
rect 3074 7590 3126 7642
rect 3138 7590 3190 7642
rect 3202 7590 3254 7642
rect 3266 7590 3318 7642
rect 9010 7590 9062 7642
rect 9074 7590 9126 7642
rect 9138 7590 9190 7642
rect 9202 7590 9254 7642
rect 9266 7590 9318 7642
rect 15010 7590 15062 7642
rect 15074 7590 15126 7642
rect 15138 7590 15190 7642
rect 15202 7590 15254 7642
rect 15266 7590 15318 7642
rect 21010 7590 21062 7642
rect 21074 7590 21126 7642
rect 21138 7590 21190 7642
rect 21202 7590 21254 7642
rect 21266 7590 21318 7642
rect 27010 7590 27062 7642
rect 27074 7590 27126 7642
rect 27138 7590 27190 7642
rect 27202 7590 27254 7642
rect 27266 7590 27318 7642
rect 23112 7531 23164 7540
rect 23112 7497 23121 7531
rect 23121 7497 23155 7531
rect 23155 7497 23164 7531
rect 23112 7488 23164 7497
rect 24492 7531 24544 7540
rect 24492 7497 24501 7531
rect 24501 7497 24535 7531
rect 24535 7497 24544 7531
rect 24492 7488 24544 7497
rect 10048 7420 10100 7472
rect 10876 7352 10928 7404
rect 16856 7420 16908 7472
rect 29000 7488 29052 7540
rect 31484 7531 31536 7540
rect 31484 7497 31493 7531
rect 31493 7497 31527 7531
rect 31527 7497 31536 7531
rect 31484 7488 31536 7497
rect 20812 7352 20864 7404
rect 23112 7352 23164 7404
rect 26424 7420 26476 7472
rect 26884 7420 26936 7472
rect 16580 7284 16632 7336
rect 17408 7216 17460 7268
rect 26240 7216 26292 7268
rect 28908 7216 28960 7268
rect 30380 7216 30432 7268
rect 10140 7148 10192 7200
rect 17684 7148 17736 7200
rect 23664 7148 23716 7200
rect 27436 7148 27488 7200
rect 30288 7148 30340 7200
rect 32772 7148 32824 7200
rect 1950 7046 2002 7098
rect 2014 7046 2066 7098
rect 2078 7046 2130 7098
rect 2142 7046 2194 7098
rect 2206 7046 2258 7098
rect 7950 7046 8002 7098
rect 8014 7046 8066 7098
rect 8078 7046 8130 7098
rect 8142 7046 8194 7098
rect 8206 7046 8258 7098
rect 13950 7046 14002 7098
rect 14014 7046 14066 7098
rect 14078 7046 14130 7098
rect 14142 7046 14194 7098
rect 14206 7046 14258 7098
rect 19950 7046 20002 7098
rect 20014 7046 20066 7098
rect 20078 7046 20130 7098
rect 20142 7046 20194 7098
rect 20206 7046 20258 7098
rect 25950 7046 26002 7098
rect 26014 7046 26066 7098
rect 26078 7046 26130 7098
rect 26142 7046 26194 7098
rect 26206 7046 26258 7098
rect 31950 7046 32002 7098
rect 32014 7046 32066 7098
rect 32078 7046 32130 7098
rect 32142 7046 32194 7098
rect 32206 7046 32258 7098
rect 5356 6944 5408 6996
rect 6276 6987 6328 6996
rect 6276 6953 6285 6987
rect 6285 6953 6319 6987
rect 6319 6953 6328 6987
rect 6276 6944 6328 6953
rect 12624 6987 12676 6996
rect 12624 6953 12633 6987
rect 12633 6953 12667 6987
rect 12667 6953 12676 6987
rect 12624 6944 12676 6953
rect 14372 6987 14424 6996
rect 14372 6953 14381 6987
rect 14381 6953 14415 6987
rect 14415 6953 14424 6987
rect 14372 6944 14424 6953
rect 16580 6987 16632 6996
rect 16580 6953 16589 6987
rect 16589 6953 16623 6987
rect 16623 6953 16632 6987
rect 16580 6944 16632 6953
rect 16856 6987 16908 6996
rect 16856 6953 16865 6987
rect 16865 6953 16899 6987
rect 16899 6953 16908 6987
rect 16856 6944 16908 6953
rect 19248 6944 19300 6996
rect 20812 6944 20864 6996
rect 7104 6808 7156 6860
rect 10968 6808 11020 6860
rect 6460 6783 6512 6792
rect 6460 6749 6469 6783
rect 6469 6749 6503 6783
rect 6503 6749 6512 6783
rect 6460 6740 6512 6749
rect 7840 6740 7892 6792
rect 10140 6783 10192 6792
rect 10140 6749 10149 6783
rect 10149 6749 10183 6783
rect 10183 6749 10192 6783
rect 10140 6740 10192 6749
rect 10416 6740 10468 6792
rect 10692 6783 10744 6792
rect 10692 6749 10701 6783
rect 10701 6749 10735 6783
rect 10735 6749 10744 6783
rect 10692 6740 10744 6749
rect 11428 6740 11480 6792
rect 12072 6740 12124 6792
rect 12808 6783 12860 6792
rect 12808 6749 12817 6783
rect 12817 6749 12851 6783
rect 12851 6749 12860 6783
rect 12808 6740 12860 6749
rect 9680 6672 9732 6724
rect 4344 6604 4396 6656
rect 9496 6604 9548 6656
rect 10600 6604 10652 6656
rect 13360 6672 13412 6724
rect 15660 6740 15712 6792
rect 15752 6783 15804 6792
rect 15752 6749 15761 6783
rect 15761 6749 15795 6783
rect 15795 6749 15804 6783
rect 15752 6740 15804 6749
rect 16120 6740 16172 6792
rect 16672 6783 16724 6792
rect 16672 6749 16681 6783
rect 16681 6749 16715 6783
rect 16715 6749 16724 6783
rect 16672 6740 16724 6749
rect 16304 6672 16356 6724
rect 16488 6672 16540 6724
rect 20720 6808 20772 6860
rect 21824 6944 21876 6996
rect 26700 6944 26752 6996
rect 17684 6783 17736 6792
rect 17684 6749 17693 6783
rect 17693 6749 17727 6783
rect 17727 6749 17736 6783
rect 17684 6740 17736 6749
rect 18420 6783 18472 6792
rect 18420 6749 18429 6783
rect 18429 6749 18463 6783
rect 18463 6749 18472 6783
rect 18420 6740 18472 6749
rect 19340 6783 19392 6792
rect 19340 6749 19349 6783
rect 19349 6749 19383 6783
rect 19383 6749 19392 6783
rect 19340 6740 19392 6749
rect 19984 6783 20036 6792
rect 19984 6749 19993 6783
rect 19993 6749 20027 6783
rect 20027 6749 20036 6783
rect 19984 6740 20036 6749
rect 22836 6808 22888 6860
rect 23480 6808 23532 6860
rect 29552 6808 29604 6860
rect 30288 6808 30340 6860
rect 20996 6783 21048 6792
rect 20996 6749 21005 6783
rect 21005 6749 21039 6783
rect 21039 6749 21048 6783
rect 20996 6740 21048 6749
rect 21640 6740 21692 6792
rect 23296 6740 23348 6792
rect 23664 6783 23716 6792
rect 23664 6749 23673 6783
rect 23673 6749 23707 6783
rect 23707 6749 23716 6783
rect 23664 6740 23716 6749
rect 24400 6783 24452 6792
rect 24400 6749 24409 6783
rect 24409 6749 24443 6783
rect 24443 6749 24452 6783
rect 24400 6740 24452 6749
rect 29368 6740 29420 6792
rect 11244 6647 11296 6656
rect 11244 6613 11253 6647
rect 11253 6613 11287 6647
rect 11287 6613 11296 6647
rect 11244 6604 11296 6613
rect 11520 6647 11572 6656
rect 11520 6613 11529 6647
rect 11529 6613 11563 6647
rect 11563 6613 11572 6647
rect 11520 6604 11572 6613
rect 11980 6604 12032 6656
rect 13452 6647 13504 6656
rect 13452 6613 13461 6647
rect 13461 6613 13495 6647
rect 13495 6613 13504 6647
rect 13452 6604 13504 6613
rect 15568 6647 15620 6656
rect 15568 6613 15577 6647
rect 15577 6613 15611 6647
rect 15611 6613 15620 6647
rect 15568 6604 15620 6613
rect 25780 6672 25832 6724
rect 17500 6647 17552 6656
rect 17500 6613 17509 6647
rect 17509 6613 17543 6647
rect 17543 6613 17552 6647
rect 17500 6604 17552 6613
rect 18236 6647 18288 6656
rect 18236 6613 18245 6647
rect 18245 6613 18279 6647
rect 18279 6613 18288 6647
rect 18236 6604 18288 6613
rect 19524 6647 19576 6656
rect 19524 6613 19533 6647
rect 19533 6613 19567 6647
rect 19567 6613 19576 6647
rect 19524 6604 19576 6613
rect 20812 6604 20864 6656
rect 21548 6604 21600 6656
rect 21640 6647 21692 6656
rect 21640 6613 21649 6647
rect 21649 6613 21683 6647
rect 21683 6613 21692 6647
rect 21640 6604 21692 6613
rect 22192 6604 22244 6656
rect 22928 6604 22980 6656
rect 23572 6647 23624 6656
rect 23572 6613 23581 6647
rect 23581 6613 23615 6647
rect 23615 6613 23624 6647
rect 23572 6604 23624 6613
rect 23848 6647 23900 6656
rect 23848 6613 23857 6647
rect 23857 6613 23891 6647
rect 23891 6613 23900 6647
rect 23848 6604 23900 6613
rect 23940 6604 23992 6656
rect 30932 6672 30984 6724
rect 27620 6604 27672 6656
rect 28724 6604 28776 6656
rect 31668 6740 31720 6792
rect 31392 6647 31444 6656
rect 31392 6613 31401 6647
rect 31401 6613 31435 6647
rect 31435 6613 31444 6647
rect 31392 6604 31444 6613
rect 31760 6647 31812 6656
rect 31760 6613 31769 6647
rect 31769 6613 31803 6647
rect 31803 6613 31812 6647
rect 31760 6604 31812 6613
rect 32312 6604 32364 6656
rect 3010 6502 3062 6554
rect 3074 6502 3126 6554
rect 3138 6502 3190 6554
rect 3202 6502 3254 6554
rect 3266 6502 3318 6554
rect 9010 6502 9062 6554
rect 9074 6502 9126 6554
rect 9138 6502 9190 6554
rect 9202 6502 9254 6554
rect 9266 6502 9318 6554
rect 15010 6502 15062 6554
rect 15074 6502 15126 6554
rect 15138 6502 15190 6554
rect 15202 6502 15254 6554
rect 15266 6502 15318 6554
rect 21010 6502 21062 6554
rect 21074 6502 21126 6554
rect 21138 6502 21190 6554
rect 21202 6502 21254 6554
rect 21266 6502 21318 6554
rect 27010 6502 27062 6554
rect 27074 6502 27126 6554
rect 27138 6502 27190 6554
rect 27202 6502 27254 6554
rect 27266 6502 27318 6554
rect 5172 6400 5224 6452
rect 5816 6400 5868 6452
rect 6920 6400 6972 6452
rect 8392 6443 8444 6452
rect 8392 6409 8401 6443
rect 8401 6409 8435 6443
rect 8435 6409 8444 6443
rect 8392 6400 8444 6409
rect 8668 6443 8720 6452
rect 8668 6409 8677 6443
rect 8677 6409 8711 6443
rect 8711 6409 8720 6443
rect 8668 6400 8720 6409
rect 8760 6400 8812 6452
rect 9404 6400 9456 6452
rect 10324 6443 10376 6452
rect 10324 6409 10333 6443
rect 10333 6409 10367 6443
rect 10367 6409 10376 6443
rect 10324 6400 10376 6409
rect 7564 6332 7616 6384
rect 6828 6307 6880 6316
rect 6828 6273 6837 6307
rect 6837 6273 6871 6307
rect 6871 6273 6880 6307
rect 6828 6264 6880 6273
rect 7840 6307 7892 6316
rect 7840 6273 7849 6307
rect 7849 6273 7883 6307
rect 7883 6273 7892 6307
rect 7840 6264 7892 6273
rect 8484 6264 8536 6316
rect 8852 6307 8904 6316
rect 8852 6273 8861 6307
rect 8861 6273 8895 6307
rect 8895 6273 8904 6307
rect 8852 6264 8904 6273
rect 9588 6264 9640 6316
rect 8944 6196 8996 6248
rect 9772 6307 9824 6316
rect 9772 6273 9781 6307
rect 9781 6273 9815 6307
rect 9815 6273 9824 6307
rect 9772 6264 9824 6273
rect 15844 6400 15896 6452
rect 16304 6400 16356 6452
rect 19800 6400 19852 6452
rect 19984 6400 20036 6452
rect 23480 6400 23532 6452
rect 23664 6400 23716 6452
rect 26424 6400 26476 6452
rect 29092 6400 29144 6452
rect 30564 6400 30616 6452
rect 31852 6443 31904 6452
rect 31852 6409 31861 6443
rect 31861 6409 31895 6443
rect 31895 6409 31904 6443
rect 31852 6400 31904 6409
rect 10600 6332 10652 6384
rect 12716 6332 12768 6384
rect 12808 6332 12860 6384
rect 21364 6332 21416 6384
rect 21640 6332 21692 6384
rect 30656 6332 30708 6384
rect 10508 6311 10560 6316
rect 10508 6277 10517 6311
rect 10517 6277 10551 6311
rect 10551 6277 10560 6311
rect 10508 6264 10560 6277
rect 10876 6307 10928 6316
rect 10876 6273 10885 6307
rect 10885 6273 10919 6307
rect 10919 6273 10928 6307
rect 10876 6264 10928 6273
rect 11796 6264 11848 6316
rect 9956 6196 10008 6248
rect 10416 6196 10468 6248
rect 19616 6264 19668 6316
rect 21548 6264 21600 6316
rect 23296 6264 23348 6316
rect 24308 6264 24360 6316
rect 24400 6264 24452 6316
rect 27804 6264 27856 6316
rect 30932 6264 30984 6316
rect 19524 6196 19576 6248
rect 30472 6196 30524 6248
rect 31300 6307 31352 6316
rect 31300 6273 31309 6307
rect 31309 6273 31343 6307
rect 31343 6273 31352 6307
rect 31300 6264 31352 6273
rect 31392 6264 31444 6316
rect 32496 6196 32548 6248
rect 4712 6128 4764 6180
rect 8576 6128 8628 6180
rect 10784 6128 10836 6180
rect 6828 6060 6880 6112
rect 9588 6060 9640 6112
rect 10140 6060 10192 6112
rect 10416 6060 10468 6112
rect 12164 6128 12216 6180
rect 18420 6128 18472 6180
rect 23204 6128 23256 6180
rect 23572 6128 23624 6180
rect 28264 6128 28316 6180
rect 31484 6171 31536 6180
rect 31484 6137 31493 6171
rect 31493 6137 31527 6171
rect 31527 6137 31536 6171
rect 31484 6128 31536 6137
rect 11060 6103 11112 6112
rect 11060 6069 11069 6103
rect 11069 6069 11103 6103
rect 11103 6069 11112 6103
rect 11060 6060 11112 6069
rect 11152 6060 11204 6112
rect 13636 6060 13688 6112
rect 15292 6060 15344 6112
rect 17592 6060 17644 6112
rect 17684 6060 17736 6112
rect 22192 6060 22244 6112
rect 22284 6103 22336 6112
rect 22284 6069 22293 6103
rect 22293 6069 22327 6103
rect 22327 6069 22336 6103
rect 22284 6060 22336 6069
rect 23848 6060 23900 6112
rect 28632 6060 28684 6112
rect 1950 5958 2002 6010
rect 2014 5958 2066 6010
rect 2078 5958 2130 6010
rect 2142 5958 2194 6010
rect 2206 5958 2258 6010
rect 7950 5958 8002 6010
rect 8014 5958 8066 6010
rect 8078 5958 8130 6010
rect 8142 5958 8194 6010
rect 8206 5958 8258 6010
rect 13950 5958 14002 6010
rect 14014 5958 14066 6010
rect 14078 5958 14130 6010
rect 14142 5958 14194 6010
rect 14206 5958 14258 6010
rect 19950 5958 20002 6010
rect 20014 5958 20066 6010
rect 20078 5958 20130 6010
rect 20142 5958 20194 6010
rect 20206 5958 20258 6010
rect 25950 5958 26002 6010
rect 26014 5958 26066 6010
rect 26078 5958 26130 6010
rect 26142 5958 26194 6010
rect 26206 5958 26258 6010
rect 31950 5958 32002 6010
rect 32014 5958 32066 6010
rect 32078 5958 32130 6010
rect 32142 5958 32194 6010
rect 32206 5958 32258 6010
rect 7196 5856 7248 5908
rect 7380 5899 7432 5908
rect 7380 5865 7389 5899
rect 7389 5865 7423 5899
rect 7423 5865 7432 5899
rect 7380 5856 7432 5865
rect 7748 5856 7800 5908
rect 7840 5856 7892 5908
rect 8944 5856 8996 5908
rect 11428 5856 11480 5908
rect 15292 5856 15344 5908
rect 16764 5856 16816 5908
rect 17592 5856 17644 5908
rect 20812 5856 20864 5908
rect 21364 5856 21416 5908
rect 31300 5856 31352 5908
rect 11152 5720 11204 5772
rect 16396 5788 16448 5840
rect 21732 5788 21784 5840
rect 22100 5788 22152 5840
rect 22284 5788 22336 5840
rect 27528 5788 27580 5840
rect 32036 5788 32088 5840
rect 32128 5831 32180 5840
rect 32128 5797 32137 5831
rect 32137 5797 32171 5831
rect 32171 5797 32180 5831
rect 32128 5788 32180 5797
rect 15752 5720 15804 5772
rect 7012 5652 7064 5704
rect 7840 5695 7892 5704
rect 7840 5661 7849 5695
rect 7849 5661 7883 5695
rect 7883 5661 7892 5695
rect 7840 5652 7892 5661
rect 9128 5695 9180 5704
rect 9128 5661 9137 5695
rect 9137 5661 9171 5695
rect 9171 5661 9180 5695
rect 9128 5652 9180 5661
rect 9588 5584 9640 5636
rect 13544 5652 13596 5704
rect 16212 5695 16264 5704
rect 16212 5661 16221 5695
rect 16221 5661 16255 5695
rect 16255 5661 16264 5695
rect 16212 5652 16264 5661
rect 6184 5516 6236 5568
rect 9680 5516 9732 5568
rect 17132 5652 17184 5704
rect 20352 5652 20404 5704
rect 31208 5695 31260 5704
rect 31208 5661 31217 5695
rect 31217 5661 31251 5695
rect 31251 5661 31260 5695
rect 31208 5652 31260 5661
rect 31300 5652 31352 5704
rect 31852 5652 31904 5704
rect 31668 5584 31720 5636
rect 31760 5559 31812 5568
rect 31760 5525 31769 5559
rect 31769 5525 31803 5559
rect 31803 5525 31812 5559
rect 31760 5516 31812 5525
rect 3010 5414 3062 5466
rect 3074 5414 3126 5466
rect 3138 5414 3190 5466
rect 3202 5414 3254 5466
rect 3266 5414 3318 5466
rect 9010 5414 9062 5466
rect 9074 5414 9126 5466
rect 9138 5414 9190 5466
rect 9202 5414 9254 5466
rect 9266 5414 9318 5466
rect 15010 5414 15062 5466
rect 15074 5414 15126 5466
rect 15138 5414 15190 5466
rect 15202 5414 15254 5466
rect 15266 5414 15318 5466
rect 21010 5414 21062 5466
rect 21074 5414 21126 5466
rect 21138 5414 21190 5466
rect 21202 5414 21254 5466
rect 21266 5414 21318 5466
rect 27010 5414 27062 5466
rect 27074 5414 27126 5466
rect 27138 5414 27190 5466
rect 27202 5414 27254 5466
rect 27266 5414 27318 5466
rect 7288 5312 7340 5364
rect 21456 5355 21508 5364
rect 21456 5321 21465 5355
rect 21465 5321 21499 5355
rect 21499 5321 21508 5355
rect 21456 5312 21508 5321
rect 15384 5244 15436 5296
rect 19064 5244 19116 5296
rect 9864 5176 9916 5228
rect 18420 5176 18472 5228
rect 31668 5219 31720 5228
rect 31668 5185 31677 5219
rect 31677 5185 31711 5219
rect 31711 5185 31720 5219
rect 31668 5176 31720 5185
rect 4620 5108 4672 5160
rect 20904 5108 20956 5160
rect 30380 5040 30432 5092
rect 31484 5015 31536 5024
rect 31484 4981 31493 5015
rect 31493 4981 31527 5015
rect 31527 4981 31536 5015
rect 31484 4972 31536 4981
rect 32864 4972 32916 5024
rect 1950 4870 2002 4922
rect 2014 4870 2066 4922
rect 2078 4870 2130 4922
rect 2142 4870 2194 4922
rect 2206 4870 2258 4922
rect 7950 4870 8002 4922
rect 8014 4870 8066 4922
rect 8078 4870 8130 4922
rect 8142 4870 8194 4922
rect 8206 4870 8258 4922
rect 13950 4870 14002 4922
rect 14014 4870 14066 4922
rect 14078 4870 14130 4922
rect 14142 4870 14194 4922
rect 14206 4870 14258 4922
rect 19950 4870 20002 4922
rect 20014 4870 20066 4922
rect 20078 4870 20130 4922
rect 20142 4870 20194 4922
rect 20206 4870 20258 4922
rect 25950 4870 26002 4922
rect 26014 4870 26066 4922
rect 26078 4870 26130 4922
rect 26142 4870 26194 4922
rect 26206 4870 26258 4922
rect 31950 4870 32002 4922
rect 32014 4870 32066 4922
rect 32078 4870 32130 4922
rect 32142 4870 32194 4922
rect 32206 4870 32258 4922
rect 13820 4768 13872 4820
rect 31392 4768 31444 4820
rect 15660 4700 15712 4752
rect 31668 4700 31720 4752
rect 572 4564 624 4616
rect 16948 4496 17000 4548
rect 28724 4632 28776 4684
rect 23756 4607 23808 4616
rect 23756 4573 23765 4607
rect 23765 4573 23799 4607
rect 23799 4573 23808 4607
rect 23756 4564 23808 4573
rect 29000 4564 29052 4616
rect 31944 4607 31996 4616
rect 31944 4573 31953 4607
rect 31953 4573 31987 4607
rect 31987 4573 31996 4607
rect 31944 4564 31996 4573
rect 27712 4496 27764 4548
rect 24768 4428 24820 4480
rect 31760 4471 31812 4480
rect 31760 4437 31769 4471
rect 31769 4437 31803 4471
rect 31803 4437 31812 4471
rect 31760 4428 31812 4437
rect 32128 4471 32180 4480
rect 32128 4437 32137 4471
rect 32137 4437 32171 4471
rect 32171 4437 32180 4471
rect 32128 4428 32180 4437
rect 3010 4326 3062 4378
rect 3074 4326 3126 4378
rect 3138 4326 3190 4378
rect 3202 4326 3254 4378
rect 3266 4326 3318 4378
rect 9010 4326 9062 4378
rect 9074 4326 9126 4378
rect 9138 4326 9190 4378
rect 9202 4326 9254 4378
rect 9266 4326 9318 4378
rect 15010 4326 15062 4378
rect 15074 4326 15126 4378
rect 15138 4326 15190 4378
rect 15202 4326 15254 4378
rect 15266 4326 15318 4378
rect 21010 4326 21062 4378
rect 21074 4326 21126 4378
rect 21138 4326 21190 4378
rect 21202 4326 21254 4378
rect 21266 4326 21318 4378
rect 27010 4326 27062 4378
rect 27074 4326 27126 4378
rect 27138 4326 27190 4378
rect 27202 4326 27254 4378
rect 27266 4326 27318 4378
rect 19432 4224 19484 4276
rect 31944 4224 31996 4276
rect 12440 4131 12492 4140
rect 12440 4097 12449 4131
rect 12449 4097 12483 4131
rect 12483 4097 12492 4131
rect 12440 4088 12492 4097
rect 17868 4088 17920 4140
rect 19248 4088 19300 4140
rect 20904 4131 20956 4140
rect 20904 4097 20913 4131
rect 20913 4097 20947 4131
rect 20947 4097 20956 4131
rect 20904 4088 20956 4097
rect 26884 4088 26936 4140
rect 31392 4088 31444 4140
rect 16396 4020 16448 4072
rect 25504 4020 25556 4072
rect 7012 3952 7064 4004
rect 31208 3952 31260 4004
rect 6920 3884 6972 3936
rect 10692 3884 10744 3936
rect 13820 3884 13872 3936
rect 15936 3884 15988 3936
rect 19800 3884 19852 3936
rect 21364 3884 21416 3936
rect 25504 3884 25556 3936
rect 26516 3884 26568 3936
rect 31484 3927 31536 3936
rect 31484 3893 31493 3927
rect 31493 3893 31527 3927
rect 31527 3893 31536 3927
rect 31484 3884 31536 3893
rect 32864 3884 32916 3936
rect 1950 3782 2002 3834
rect 2014 3782 2066 3834
rect 2078 3782 2130 3834
rect 2142 3782 2194 3834
rect 2206 3782 2258 3834
rect 7950 3782 8002 3834
rect 8014 3782 8066 3834
rect 8078 3782 8130 3834
rect 8142 3782 8194 3834
rect 8206 3782 8258 3834
rect 13950 3782 14002 3834
rect 14014 3782 14066 3834
rect 14078 3782 14130 3834
rect 14142 3782 14194 3834
rect 14206 3782 14258 3834
rect 19950 3782 20002 3834
rect 20014 3782 20066 3834
rect 20078 3782 20130 3834
rect 20142 3782 20194 3834
rect 20206 3782 20258 3834
rect 25950 3782 26002 3834
rect 26014 3782 26066 3834
rect 26078 3782 26130 3834
rect 26142 3782 26194 3834
rect 26206 3782 26258 3834
rect 31950 3782 32002 3834
rect 32014 3782 32066 3834
rect 32078 3782 32130 3834
rect 32142 3782 32194 3834
rect 32206 3782 32258 3834
rect 7012 3680 7064 3732
rect 9588 3680 9640 3732
rect 14924 3680 14976 3732
rect 9404 3612 9456 3664
rect 1308 3544 1360 3596
rect 1124 3476 1176 3528
rect 7472 3544 7524 3596
rect 9496 3544 9548 3596
rect 13728 3612 13780 3664
rect 15568 3680 15620 3732
rect 15660 3723 15712 3732
rect 15660 3689 15669 3723
rect 15669 3689 15703 3723
rect 15703 3689 15712 3723
rect 15660 3680 15712 3689
rect 15936 3723 15988 3732
rect 15936 3689 15945 3723
rect 15945 3689 15979 3723
rect 15979 3689 15988 3723
rect 15936 3680 15988 3689
rect 16488 3680 16540 3732
rect 17960 3723 18012 3732
rect 17960 3689 17969 3723
rect 17969 3689 18003 3723
rect 18003 3689 18012 3723
rect 17960 3680 18012 3689
rect 18144 3723 18196 3732
rect 18144 3689 18153 3723
rect 18153 3689 18187 3723
rect 18187 3689 18196 3723
rect 18144 3680 18196 3689
rect 18880 3680 18932 3732
rect 19064 3723 19116 3732
rect 19064 3689 19073 3723
rect 19073 3689 19107 3723
rect 19107 3689 19116 3723
rect 19064 3680 19116 3689
rect 19432 3723 19484 3732
rect 19432 3689 19441 3723
rect 19441 3689 19475 3723
rect 19475 3689 19484 3723
rect 19432 3680 19484 3689
rect 19524 3680 19576 3732
rect 24216 3680 24268 3732
rect 25504 3723 25556 3732
rect 25504 3689 25513 3723
rect 25513 3689 25547 3723
rect 25547 3689 25556 3723
rect 25504 3680 25556 3689
rect 25872 3680 25924 3732
rect 1308 3408 1360 3460
rect 10692 3519 10744 3528
rect 10692 3485 10701 3519
rect 10701 3485 10735 3519
rect 10735 3485 10744 3519
rect 10692 3476 10744 3485
rect 12072 3476 12124 3528
rect 14556 3519 14608 3528
rect 14556 3485 14565 3519
rect 14565 3485 14599 3519
rect 14599 3485 14608 3519
rect 14556 3476 14608 3485
rect 15568 3476 15620 3528
rect 4896 3383 4948 3392
rect 4896 3349 4905 3383
rect 4905 3349 4939 3383
rect 4939 3349 4948 3383
rect 4896 3340 4948 3349
rect 8392 3383 8444 3392
rect 8392 3349 8401 3383
rect 8401 3349 8435 3383
rect 8435 3349 8444 3383
rect 8392 3340 8444 3349
rect 16396 3408 16448 3460
rect 10600 3383 10652 3392
rect 10600 3349 10609 3383
rect 10609 3349 10643 3383
rect 10643 3349 10652 3383
rect 10600 3340 10652 3349
rect 11520 3383 11572 3392
rect 11520 3349 11529 3383
rect 11529 3349 11563 3383
rect 11563 3349 11572 3383
rect 11520 3340 11572 3349
rect 12164 3383 12216 3392
rect 12164 3349 12173 3383
rect 12173 3349 12207 3383
rect 12207 3349 12216 3383
rect 12164 3340 12216 3349
rect 12440 3383 12492 3392
rect 12440 3349 12449 3383
rect 12449 3349 12483 3383
rect 12483 3349 12492 3383
rect 12440 3340 12492 3349
rect 16856 3476 16908 3528
rect 17408 3612 17460 3664
rect 19800 3612 19852 3664
rect 31852 3612 31904 3664
rect 17776 3519 17828 3528
rect 17776 3485 17785 3519
rect 17785 3485 17819 3519
rect 17819 3485 17828 3519
rect 17776 3476 17828 3485
rect 18880 3519 18932 3528
rect 18880 3485 18889 3519
rect 18889 3485 18923 3519
rect 18923 3485 18932 3519
rect 18880 3476 18932 3485
rect 19248 3519 19300 3528
rect 19248 3485 19257 3519
rect 19257 3485 19291 3519
rect 19291 3485 19300 3519
rect 19248 3476 19300 3485
rect 19524 3519 19576 3528
rect 19524 3485 19533 3519
rect 19533 3485 19567 3519
rect 19567 3485 19576 3519
rect 19524 3476 19576 3485
rect 29000 3544 29052 3596
rect 21824 3519 21876 3528
rect 21824 3485 21833 3519
rect 21833 3485 21867 3519
rect 21867 3485 21876 3519
rect 21824 3476 21876 3485
rect 22192 3519 22244 3528
rect 22192 3485 22201 3519
rect 22201 3485 22235 3519
rect 22235 3485 22244 3519
rect 22192 3476 22244 3485
rect 22468 3519 22520 3528
rect 22468 3485 22477 3519
rect 22477 3485 22511 3519
rect 22511 3485 22520 3519
rect 22468 3476 22520 3485
rect 23480 3476 23532 3528
rect 25596 3519 25648 3528
rect 25596 3485 25605 3519
rect 25605 3485 25639 3519
rect 25639 3485 25648 3519
rect 25596 3476 25648 3485
rect 25688 3476 25740 3528
rect 31576 3519 31628 3528
rect 31576 3485 31585 3519
rect 31585 3485 31619 3519
rect 31619 3485 31628 3519
rect 31576 3476 31628 3485
rect 31944 3519 31996 3528
rect 31944 3485 31953 3519
rect 31953 3485 31987 3519
rect 31987 3485 31996 3519
rect 31944 3476 31996 3485
rect 31300 3408 31352 3460
rect 16580 3383 16632 3392
rect 16580 3349 16589 3383
rect 16589 3349 16623 3383
rect 16623 3349 16632 3383
rect 16580 3340 16632 3349
rect 16672 3383 16724 3392
rect 16672 3349 16681 3383
rect 16681 3349 16715 3383
rect 16715 3349 16724 3383
rect 16672 3340 16724 3349
rect 16856 3383 16908 3392
rect 16856 3349 16865 3383
rect 16865 3349 16899 3383
rect 16899 3349 16908 3383
rect 16856 3340 16908 3349
rect 17224 3383 17276 3392
rect 17224 3349 17233 3383
rect 17233 3349 17267 3383
rect 17267 3349 17276 3383
rect 17224 3340 17276 3349
rect 17500 3383 17552 3392
rect 17500 3349 17509 3383
rect 17509 3349 17543 3383
rect 17543 3349 17552 3383
rect 17500 3340 17552 3349
rect 18512 3383 18564 3392
rect 18512 3349 18521 3383
rect 18521 3349 18555 3383
rect 18555 3349 18564 3383
rect 18512 3340 18564 3349
rect 18788 3383 18840 3392
rect 18788 3349 18797 3383
rect 18797 3349 18831 3383
rect 18831 3349 18840 3383
rect 18788 3340 18840 3349
rect 19248 3340 19300 3392
rect 22376 3383 22428 3392
rect 22376 3349 22385 3383
rect 22385 3349 22419 3383
rect 22419 3349 22428 3383
rect 22376 3340 22428 3349
rect 23388 3340 23440 3392
rect 26332 3340 26384 3392
rect 31760 3383 31812 3392
rect 31760 3349 31769 3383
rect 31769 3349 31803 3383
rect 31803 3349 31812 3383
rect 31760 3340 31812 3349
rect 32128 3383 32180 3392
rect 32128 3349 32137 3383
rect 32137 3349 32171 3383
rect 32171 3349 32180 3383
rect 32128 3340 32180 3349
rect 3010 3238 3062 3290
rect 3074 3238 3126 3290
rect 3138 3238 3190 3290
rect 3202 3238 3254 3290
rect 3266 3238 3318 3290
rect 9010 3238 9062 3290
rect 9074 3238 9126 3290
rect 9138 3238 9190 3290
rect 9202 3238 9254 3290
rect 9266 3238 9318 3290
rect 15010 3238 15062 3290
rect 15074 3238 15126 3290
rect 15138 3238 15190 3290
rect 15202 3238 15254 3290
rect 15266 3238 15318 3290
rect 21010 3238 21062 3290
rect 21074 3238 21126 3290
rect 21138 3238 21190 3290
rect 21202 3238 21254 3290
rect 21266 3238 21318 3290
rect 27010 3238 27062 3290
rect 27074 3238 27126 3290
rect 27138 3238 27190 3290
rect 27202 3238 27254 3290
rect 27266 3238 27318 3290
rect 4344 3136 4396 3188
rect 14556 3136 14608 3188
rect 17500 3136 17552 3188
rect 31944 3136 31996 3188
rect 9404 3068 9456 3120
rect 12072 3068 12124 3120
rect 17224 3068 17276 3120
rect 31576 3068 31628 3120
rect 5908 3000 5960 3052
rect 16580 3000 16632 3052
rect 17776 3000 17828 3052
rect 18788 3000 18840 3052
rect 26884 3000 26936 3052
rect 30380 3000 30432 3052
rect 31668 3043 31720 3052
rect 31668 3009 31677 3043
rect 31677 3009 31711 3043
rect 31711 3009 31720 3043
rect 31668 3000 31720 3009
rect 10600 2864 10652 2916
rect 31392 2864 31444 2916
rect 31760 2796 31812 2848
rect 32864 2796 32916 2848
rect 1950 2694 2002 2746
rect 2014 2694 2066 2746
rect 2078 2694 2130 2746
rect 2142 2694 2194 2746
rect 2206 2694 2258 2746
rect 7950 2694 8002 2746
rect 8014 2694 8066 2746
rect 8078 2694 8130 2746
rect 8142 2694 8194 2746
rect 8206 2694 8258 2746
rect 13950 2694 14002 2746
rect 14014 2694 14066 2746
rect 14078 2694 14130 2746
rect 14142 2694 14194 2746
rect 14206 2694 14258 2746
rect 19950 2694 20002 2746
rect 20014 2694 20066 2746
rect 20078 2694 20130 2746
rect 20142 2694 20194 2746
rect 20206 2694 20258 2746
rect 25950 2694 26002 2746
rect 26014 2694 26066 2746
rect 26078 2694 26130 2746
rect 26142 2694 26194 2746
rect 26206 2694 26258 2746
rect 31950 2694 32002 2746
rect 32014 2694 32066 2746
rect 32078 2694 32130 2746
rect 32142 2694 32194 2746
rect 32206 2694 32258 2746
rect 12440 2592 12492 2644
rect 12164 2524 12216 2576
rect 11520 2456 11572 2508
rect 30472 2456 30524 2508
rect 4896 2388 4948 2440
rect 8392 2320 8444 2372
rect 30840 2388 30892 2440
rect 30380 2252 30432 2304
rect 30748 2295 30800 2304
rect 30748 2261 30757 2295
rect 30757 2261 30791 2295
rect 30791 2261 30800 2295
rect 30748 2252 30800 2261
rect 31116 2295 31168 2304
rect 31116 2261 31125 2295
rect 31125 2261 31159 2295
rect 31159 2261 31168 2295
rect 31116 2252 31168 2261
rect 31484 2295 31536 2304
rect 31484 2261 31493 2295
rect 31493 2261 31527 2295
rect 31527 2261 31536 2295
rect 31484 2252 31536 2261
rect 31852 2295 31904 2304
rect 31852 2261 31861 2295
rect 31861 2261 31895 2295
rect 31895 2261 31904 2295
rect 31852 2252 31904 2261
rect 3010 2150 3062 2202
rect 3074 2150 3126 2202
rect 3138 2150 3190 2202
rect 3202 2150 3254 2202
rect 3266 2150 3318 2202
rect 9010 2150 9062 2202
rect 9074 2150 9126 2202
rect 9138 2150 9190 2202
rect 9202 2150 9254 2202
rect 9266 2150 9318 2202
rect 15010 2150 15062 2202
rect 15074 2150 15126 2202
rect 15138 2150 15190 2202
rect 15202 2150 15254 2202
rect 15266 2150 15318 2202
rect 21010 2150 21062 2202
rect 21074 2150 21126 2202
rect 21138 2150 21190 2202
rect 21202 2150 21254 2202
rect 21266 2150 21318 2202
rect 27010 2150 27062 2202
rect 27074 2150 27126 2202
rect 27138 2150 27190 2202
rect 27202 2150 27254 2202
rect 27266 2150 27318 2202
rect 12164 2048 12216 2100
rect 25688 2048 25740 2100
rect 2780 144 2832 196
rect 22192 76 22244 128
rect 1308 8 1360 60
rect 21824 8 21876 60
<< metal2 >>
rect 4158 11194 4214 11250
rect 4434 11194 4490 11250
rect 4710 11194 4766 11250
rect 4986 11194 5042 11250
rect 5262 11194 5318 11250
rect 5538 11194 5594 11250
rect 5814 11194 5870 11250
rect 6090 11194 6146 11250
rect 6366 11194 6422 11250
rect 6642 11194 6698 11250
rect 6918 11194 6974 11250
rect 7194 11194 7250 11250
rect 7470 11194 7526 11250
rect 7746 11194 7802 11250
rect 8022 11194 8078 11250
rect 8298 11194 8354 11250
rect 8574 11194 8630 11250
rect 8850 11194 8906 11250
rect 9126 11194 9182 11250
rect 9402 11194 9458 11250
rect 9678 11194 9734 11250
rect 9954 11194 10010 11250
rect 10230 11194 10286 11250
rect 10506 11194 10562 11250
rect 10782 11194 10838 11250
rect 11058 11194 11114 11250
rect 11334 11194 11390 11250
rect 11610 11194 11666 11250
rect 11886 11194 11942 11250
rect 12162 11194 12218 11250
rect 12438 11194 12494 11250
rect 12714 11194 12770 11250
rect 12990 11194 13046 11250
rect 13266 11194 13322 11250
rect 13542 11194 13598 11250
rect 13818 11194 13874 11250
rect 14094 11194 14150 11250
rect 14370 11194 14426 11250
rect 14646 11194 14702 11250
rect 14922 11194 14978 11250
rect 15198 11194 15254 11250
rect 15474 11194 15530 11250
rect 15750 11194 15806 11250
rect 16026 11194 16082 11250
rect 16302 11194 16358 11250
rect 16578 11194 16634 11250
rect 16854 11194 16910 11250
rect 17130 11194 17186 11250
rect 17406 11194 17462 11250
rect 17682 11194 17738 11250
rect 17958 11194 18014 11250
rect 18234 11194 18290 11250
rect 18510 11194 18566 11250
rect 18786 11194 18842 11250
rect 19062 11194 19118 11250
rect 19338 11194 19394 11250
rect 19614 11194 19670 11250
rect 19890 11194 19946 11250
rect 20166 11194 20222 11250
rect 20442 11194 20498 11250
rect 20718 11194 20774 11250
rect 20994 11194 21050 11250
rect 21270 11194 21326 11250
rect 21546 11194 21602 11250
rect 21822 11194 21878 11250
rect 22098 11194 22154 11250
rect 22374 11194 22430 11250
rect 22650 11194 22706 11250
rect 22926 11194 22982 11250
rect 23202 11194 23258 11250
rect 23478 11194 23534 11250
rect 23754 11194 23810 11250
rect 24030 11194 24086 11250
rect 24306 11194 24362 11250
rect 24582 11194 24638 11250
rect 24858 11194 24914 11250
rect 25134 11194 25190 11250
rect 25410 11194 25466 11250
rect 25686 11194 25742 11250
rect 25962 11194 26018 11250
rect 26238 11194 26294 11250
rect 26514 11194 26570 11250
rect 26790 11194 26846 11250
rect 27066 11194 27122 11250
rect 27342 11194 27398 11250
rect 27618 11194 27674 11250
rect 27894 11194 27950 11250
rect 28170 11194 28226 11250
rect 28446 11194 28502 11250
rect 28722 11194 28778 11250
rect 28998 11194 29054 11250
rect 29274 11194 29330 11250
rect 29550 11194 29606 11250
rect 3010 8732 3318 8741
rect 3010 8730 3016 8732
rect 3072 8730 3096 8732
rect 3152 8730 3176 8732
rect 3232 8730 3256 8732
rect 3312 8730 3318 8732
rect 3072 8678 3074 8730
rect 3254 8678 3256 8730
rect 3010 8676 3016 8678
rect 3072 8676 3096 8678
rect 3152 8676 3176 8678
rect 3232 8676 3256 8678
rect 3312 8676 3318 8678
rect 3010 8667 3318 8676
rect 1950 8188 2258 8197
rect 1950 8186 1956 8188
rect 2012 8186 2036 8188
rect 2092 8186 2116 8188
rect 2172 8186 2196 8188
rect 2252 8186 2258 8188
rect 2012 8134 2014 8186
rect 2194 8134 2196 8186
rect 1950 8132 1956 8134
rect 2012 8132 2036 8134
rect 2092 8132 2116 8134
rect 2172 8132 2196 8134
rect 2252 8132 2258 8134
rect 1950 8123 2258 8132
rect 4172 8090 4200 11194
rect 4448 8634 4476 11194
rect 4724 8634 4752 11194
rect 5000 8634 5028 11194
rect 4436 8628 4488 8634
rect 4436 8570 4488 8576
rect 4712 8628 4764 8634
rect 4712 8570 4764 8576
rect 4988 8628 5040 8634
rect 4988 8570 5040 8576
rect 4344 8492 4396 8498
rect 4344 8434 4396 8440
rect 4712 8492 4764 8498
rect 4712 8434 4764 8440
rect 5172 8492 5224 8498
rect 5172 8434 5224 8440
rect 4160 8084 4212 8090
rect 4160 8026 4212 8032
rect 3010 7644 3318 7653
rect 3010 7642 3016 7644
rect 3072 7642 3096 7644
rect 3152 7642 3176 7644
rect 3232 7642 3256 7644
rect 3312 7642 3318 7644
rect 3072 7590 3074 7642
rect 3254 7590 3256 7642
rect 3010 7588 3016 7590
rect 3072 7588 3096 7590
rect 3152 7588 3176 7590
rect 3232 7588 3256 7590
rect 3312 7588 3318 7590
rect 3010 7579 3318 7588
rect 1950 7100 2258 7109
rect 1950 7098 1956 7100
rect 2012 7098 2036 7100
rect 2092 7098 2116 7100
rect 2172 7098 2196 7100
rect 2252 7098 2258 7100
rect 2012 7046 2014 7098
rect 2194 7046 2196 7098
rect 1950 7044 1956 7046
rect 2012 7044 2036 7046
rect 2092 7044 2116 7046
rect 2172 7044 2196 7046
rect 2252 7044 2258 7046
rect 1950 7035 2258 7044
rect 4356 6662 4384 8434
rect 4344 6656 4396 6662
rect 570 6624 626 6633
rect 4344 6598 4396 6604
rect 570 6559 626 6568
rect 584 4622 612 6559
rect 3010 6556 3318 6565
rect 3010 6554 3016 6556
rect 3072 6554 3096 6556
rect 3152 6554 3176 6556
rect 3232 6554 3256 6556
rect 3312 6554 3318 6556
rect 3072 6502 3074 6554
rect 3254 6502 3256 6554
rect 3010 6500 3016 6502
rect 3072 6500 3096 6502
rect 3152 6500 3176 6502
rect 3232 6500 3256 6502
rect 3312 6500 3318 6502
rect 3010 6491 3318 6500
rect 4618 6216 4674 6225
rect 4724 6186 4752 8434
rect 5184 6458 5212 8434
rect 5276 8090 5304 11194
rect 5552 8634 5580 11194
rect 5828 8634 5856 11194
rect 5540 8628 5592 8634
rect 5540 8570 5592 8576
rect 5816 8628 5868 8634
rect 5816 8570 5868 8576
rect 5816 8492 5868 8498
rect 5816 8434 5868 8440
rect 5264 8084 5316 8090
rect 5264 8026 5316 8032
rect 5356 7880 5408 7886
rect 5356 7822 5408 7828
rect 5368 7002 5396 7822
rect 5356 6996 5408 7002
rect 5356 6938 5408 6944
rect 5828 6458 5856 8434
rect 6104 8090 6132 11194
rect 6380 8634 6408 11194
rect 6458 10840 6514 10849
rect 6458 10775 6514 10784
rect 6368 8628 6420 8634
rect 6368 8570 6420 8576
rect 6184 8492 6236 8498
rect 6184 8434 6236 8440
rect 6092 8084 6144 8090
rect 6092 8026 6144 8032
rect 5172 6452 5224 6458
rect 5172 6394 5224 6400
rect 5816 6452 5868 6458
rect 5816 6394 5868 6400
rect 4618 6151 4674 6160
rect 4712 6180 4764 6186
rect 1950 6012 2258 6021
rect 1950 6010 1956 6012
rect 2012 6010 2036 6012
rect 2092 6010 2116 6012
rect 2172 6010 2196 6012
rect 2252 6010 2258 6012
rect 2012 5958 2014 6010
rect 2194 5958 2196 6010
rect 1950 5956 1956 5958
rect 2012 5956 2036 5958
rect 2092 5956 2116 5958
rect 2172 5956 2196 5958
rect 2252 5956 2258 5958
rect 1950 5947 2258 5956
rect 3010 5468 3318 5477
rect 3010 5466 3016 5468
rect 3072 5466 3096 5468
rect 3152 5466 3176 5468
rect 3232 5466 3256 5468
rect 3312 5466 3318 5468
rect 3072 5414 3074 5466
rect 3254 5414 3256 5466
rect 3010 5412 3016 5414
rect 3072 5412 3096 5414
rect 3152 5412 3176 5414
rect 3232 5412 3256 5414
rect 3312 5412 3318 5414
rect 3010 5403 3318 5412
rect 1306 5264 1362 5273
rect 1306 5199 1362 5208
rect 572 4616 624 4622
rect 572 4558 624 4564
rect 1320 3602 1348 5199
rect 4632 5166 4660 6151
rect 4712 6122 4764 6128
rect 6196 5574 6224 8434
rect 6276 7812 6328 7818
rect 6276 7754 6328 7760
rect 6288 7002 6316 7754
rect 6276 6996 6328 7002
rect 6276 6938 6328 6944
rect 6472 6798 6500 10775
rect 6656 8090 6684 11194
rect 6932 8634 6960 11194
rect 7010 10432 7066 10441
rect 7010 10367 7066 10376
rect 6920 8628 6972 8634
rect 6920 8570 6972 8576
rect 6644 8084 6696 8090
rect 6644 8026 6696 8032
rect 6920 7880 6972 7886
rect 6920 7822 6972 7828
rect 6460 6792 6512 6798
rect 6460 6734 6512 6740
rect 6932 6458 6960 7822
rect 6920 6452 6972 6458
rect 6920 6394 6972 6400
rect 6828 6316 6880 6322
rect 6828 6258 6880 6264
rect 6840 6118 6868 6258
rect 6828 6112 6880 6118
rect 6828 6054 6880 6060
rect 7024 5710 7052 10367
rect 7208 8634 7236 11194
rect 7196 8628 7248 8634
rect 7196 8570 7248 8576
rect 7104 8492 7156 8498
rect 7104 8434 7156 8440
rect 7288 8492 7340 8498
rect 7288 8434 7340 8440
rect 7380 8492 7432 8498
rect 7380 8434 7432 8440
rect 7116 6866 7144 8434
rect 7196 7880 7248 7886
rect 7196 7822 7248 7828
rect 7104 6860 7156 6866
rect 7104 6802 7156 6808
rect 7208 5914 7236 7822
rect 7196 5908 7248 5914
rect 7196 5850 7248 5856
rect 7012 5704 7064 5710
rect 7012 5646 7064 5652
rect 6184 5568 6236 5574
rect 6184 5510 6236 5516
rect 7300 5370 7328 8434
rect 7392 5914 7420 8434
rect 7484 8090 7512 11194
rect 7562 9752 7618 9761
rect 7562 9687 7618 9696
rect 7472 8084 7524 8090
rect 7472 8026 7524 8032
rect 7576 6390 7604 9687
rect 7656 9444 7708 9450
rect 7656 9386 7708 9392
rect 7564 6384 7616 6390
rect 7564 6326 7616 6332
rect 7380 5908 7432 5914
rect 7380 5850 7432 5856
rect 7668 5692 7696 9386
rect 7760 8634 7788 11194
rect 7838 10024 7894 10033
rect 7838 9959 7894 9968
rect 7748 8628 7800 8634
rect 7748 8570 7800 8576
rect 7748 8492 7800 8498
rect 7748 8434 7800 8440
rect 7760 5914 7788 8434
rect 7852 6798 7880 9959
rect 8036 8634 8064 11194
rect 8024 8628 8076 8634
rect 8024 8570 8076 8576
rect 7950 8188 8258 8197
rect 7950 8186 7956 8188
rect 8012 8186 8036 8188
rect 8092 8186 8116 8188
rect 8172 8186 8196 8188
rect 8252 8186 8258 8188
rect 8012 8134 8014 8186
rect 8194 8134 8196 8186
rect 7950 8132 7956 8134
rect 8012 8132 8036 8134
rect 8092 8132 8116 8134
rect 8172 8132 8196 8134
rect 8252 8132 8258 8134
rect 7950 8123 8258 8132
rect 8312 8090 8340 11194
rect 8392 9308 8444 9314
rect 8392 9250 8444 9256
rect 8300 8084 8352 8090
rect 8300 8026 8352 8032
rect 7950 7100 8258 7109
rect 7950 7098 7956 7100
rect 8012 7098 8036 7100
rect 8092 7098 8116 7100
rect 8172 7098 8196 7100
rect 8252 7098 8258 7100
rect 8012 7046 8014 7098
rect 8194 7046 8196 7098
rect 7950 7044 7956 7046
rect 8012 7044 8036 7046
rect 8092 7044 8116 7046
rect 8172 7044 8196 7046
rect 8252 7044 8258 7046
rect 7950 7035 8258 7044
rect 7840 6792 7892 6798
rect 7840 6734 7892 6740
rect 8404 6458 8432 9250
rect 8484 8628 8536 8634
rect 8588 8616 8616 11194
rect 8864 9296 8892 11194
rect 8772 9268 8892 9296
rect 8772 8634 8800 9268
rect 9140 9194 9168 11194
rect 8864 9166 9168 9194
rect 8536 8588 8616 8616
rect 8760 8628 8812 8634
rect 8484 8570 8536 8576
rect 8760 8570 8812 8576
rect 8668 8492 8720 8498
rect 8720 8452 8800 8480
rect 8668 8434 8720 8440
rect 8576 8424 8628 8430
rect 8576 8366 8628 8372
rect 8484 7948 8536 7954
rect 8484 7890 8536 7896
rect 8392 6452 8444 6458
rect 8392 6394 8444 6400
rect 8496 6322 8524 7890
rect 7840 6316 7892 6322
rect 7840 6258 7892 6264
rect 8484 6316 8536 6322
rect 8484 6258 8536 6264
rect 7852 5914 7880 6258
rect 8588 6186 8616 8366
rect 8668 7880 8720 7886
rect 8668 7822 8720 7828
rect 8680 6458 8708 7822
rect 8772 6458 8800 8452
rect 8864 8090 8892 9166
rect 9010 8732 9318 8741
rect 9010 8730 9016 8732
rect 9072 8730 9096 8732
rect 9152 8730 9176 8732
rect 9232 8730 9256 8732
rect 9312 8730 9318 8732
rect 9072 8678 9074 8730
rect 9254 8678 9256 8730
rect 9010 8676 9016 8678
rect 9072 8676 9096 8678
rect 9152 8676 9176 8678
rect 9232 8676 9256 8678
rect 9312 8676 9318 8678
rect 9010 8667 9318 8676
rect 9416 8634 9444 11194
rect 9404 8628 9456 8634
rect 9404 8570 9456 8576
rect 9692 8090 9720 11194
rect 9864 9172 9916 9178
rect 9864 9114 9916 9120
rect 9876 8498 9904 9114
rect 9968 8634 9996 11194
rect 10046 9616 10102 9625
rect 10046 9551 10102 9560
rect 9956 8628 10008 8634
rect 9956 8570 10008 8576
rect 9864 8492 9916 8498
rect 9864 8434 9916 8440
rect 9956 8288 10008 8294
rect 9956 8230 10008 8236
rect 8852 8084 8904 8090
rect 8852 8026 8904 8032
rect 9680 8084 9732 8090
rect 9680 8026 9732 8032
rect 9496 7880 9548 7886
rect 9496 7822 9548 7828
rect 9404 7812 9456 7818
rect 9404 7754 9456 7760
rect 9010 7644 9318 7653
rect 9010 7642 9016 7644
rect 9072 7642 9096 7644
rect 9152 7642 9176 7644
rect 9232 7642 9256 7644
rect 9312 7642 9318 7644
rect 9072 7590 9074 7642
rect 9254 7590 9256 7642
rect 9010 7588 9016 7590
rect 9072 7588 9096 7590
rect 9152 7588 9176 7590
rect 9232 7588 9256 7590
rect 9312 7588 9318 7590
rect 9010 7579 9318 7588
rect 8850 7168 8906 7177
rect 8850 7103 8906 7112
rect 8668 6452 8720 6458
rect 8668 6394 8720 6400
rect 8760 6452 8812 6458
rect 8760 6394 8812 6400
rect 8864 6322 8892 7103
rect 9010 6556 9318 6565
rect 9010 6554 9016 6556
rect 9072 6554 9096 6556
rect 9152 6554 9176 6556
rect 9232 6554 9256 6556
rect 9312 6554 9318 6556
rect 9072 6502 9074 6554
rect 9254 6502 9256 6554
rect 9010 6500 9016 6502
rect 9072 6500 9096 6502
rect 9152 6500 9176 6502
rect 9232 6500 9256 6502
rect 9312 6500 9318 6502
rect 9010 6491 9318 6500
rect 9416 6458 9444 7754
rect 9508 6662 9536 7822
rect 9586 7712 9642 7721
rect 9586 7647 9642 7656
rect 9600 7426 9628 7647
rect 9600 7398 9720 7426
rect 9586 7304 9642 7313
rect 9586 7239 9642 7248
rect 9496 6656 9548 6662
rect 9496 6598 9548 6604
rect 9404 6452 9456 6458
rect 9404 6394 9456 6400
rect 9600 6322 9628 7239
rect 9692 7177 9720 7398
rect 9678 7168 9734 7177
rect 9678 7103 9734 7112
rect 9862 7032 9918 7041
rect 9862 6967 9918 6976
rect 9680 6724 9732 6730
rect 9680 6666 9732 6672
rect 8852 6316 8904 6322
rect 8852 6258 8904 6264
rect 9588 6316 9640 6322
rect 9588 6258 9640 6264
rect 8944 6248 8996 6254
rect 8944 6190 8996 6196
rect 9126 6216 9182 6225
rect 8576 6180 8628 6186
rect 8576 6122 8628 6128
rect 7950 6012 8258 6021
rect 7950 6010 7956 6012
rect 8012 6010 8036 6012
rect 8092 6010 8116 6012
rect 8172 6010 8196 6012
rect 8252 6010 8258 6012
rect 8012 5958 8014 6010
rect 8194 5958 8196 6010
rect 7950 5956 7956 5958
rect 8012 5956 8036 5958
rect 8092 5956 8116 5958
rect 8172 5956 8196 5958
rect 8252 5956 8258 5958
rect 7950 5947 8258 5956
rect 8956 5914 8984 6190
rect 9126 6151 9182 6160
rect 7748 5908 7800 5914
rect 7748 5850 7800 5856
rect 7840 5908 7892 5914
rect 7840 5850 7892 5856
rect 8944 5908 8996 5914
rect 8944 5850 8996 5856
rect 9140 5710 9168 6151
rect 9588 6112 9640 6118
rect 9588 6054 9640 6060
rect 7840 5704 7892 5710
rect 7668 5664 7840 5692
rect 7840 5646 7892 5652
rect 9128 5704 9180 5710
rect 9128 5646 9180 5652
rect 9600 5642 9628 6054
rect 9588 5636 9640 5642
rect 9588 5578 9640 5584
rect 9692 5574 9720 6666
rect 9770 6488 9826 6497
rect 9770 6423 9826 6432
rect 9784 6322 9812 6423
rect 9772 6316 9824 6322
rect 9772 6258 9824 6264
rect 9680 5568 9732 5574
rect 9680 5510 9732 5516
rect 9010 5468 9318 5477
rect 9010 5466 9016 5468
rect 9072 5466 9096 5468
rect 9152 5466 9176 5468
rect 9232 5466 9256 5468
rect 9312 5466 9318 5468
rect 9072 5414 9074 5466
rect 9254 5414 9256 5466
rect 9010 5412 9016 5414
rect 9072 5412 9096 5414
rect 9152 5412 9176 5414
rect 9232 5412 9256 5414
rect 9312 5412 9318 5414
rect 9010 5403 9318 5412
rect 7288 5364 7340 5370
rect 7288 5306 7340 5312
rect 6918 5264 6974 5273
rect 9876 5234 9904 6967
rect 9968 6254 9996 8230
rect 10060 8022 10088 9551
rect 10244 8634 10272 11194
rect 10324 9240 10376 9246
rect 10324 9182 10376 9188
rect 10232 8628 10284 8634
rect 10232 8570 10284 8576
rect 10336 8378 10364 9182
rect 10416 9104 10468 9110
rect 10416 9046 10468 9052
rect 10428 8498 10456 9046
rect 10520 8634 10548 11194
rect 10600 9036 10652 9042
rect 10600 8978 10652 8984
rect 10508 8628 10560 8634
rect 10508 8570 10560 8576
rect 10416 8492 10468 8498
rect 10416 8434 10468 8440
rect 10232 8356 10284 8362
rect 10336 8350 10548 8378
rect 10232 8298 10284 8304
rect 10048 8016 10100 8022
rect 10048 7958 10100 7964
rect 10048 7880 10100 7886
rect 10048 7822 10100 7828
rect 10060 7478 10088 7822
rect 10048 7472 10100 7478
rect 10048 7414 10100 7420
rect 10140 7200 10192 7206
rect 10140 7142 10192 7148
rect 10152 6798 10180 7142
rect 10140 6792 10192 6798
rect 10140 6734 10192 6740
rect 10244 6440 10272 8298
rect 10416 6792 10468 6798
rect 10416 6734 10468 6740
rect 10324 6452 10376 6458
rect 10244 6412 10324 6440
rect 10324 6394 10376 6400
rect 10428 6254 10456 6734
rect 10520 6322 10548 8350
rect 10612 6662 10640 8978
rect 10692 8560 10744 8566
rect 10692 8502 10744 8508
rect 10704 6882 10732 8502
rect 10796 8090 10824 11194
rect 10968 8900 11020 8906
rect 10968 8842 11020 8848
rect 10980 8498 11008 8842
rect 11072 8634 11100 11194
rect 11060 8628 11112 8634
rect 11060 8570 11112 8576
rect 11244 8560 11296 8566
rect 11244 8502 11296 8508
rect 10968 8492 11020 8498
rect 10968 8434 11020 8440
rect 10784 8084 10836 8090
rect 10784 8026 10836 8032
rect 10876 7404 10928 7410
rect 10876 7346 10928 7352
rect 10704 6854 10824 6882
rect 10692 6792 10744 6798
rect 10690 6760 10692 6769
rect 10744 6760 10746 6769
rect 10690 6695 10746 6704
rect 10600 6656 10652 6662
rect 10600 6598 10652 6604
rect 10598 6488 10654 6497
rect 10598 6423 10654 6432
rect 10612 6390 10640 6423
rect 10600 6384 10652 6390
rect 10600 6326 10652 6332
rect 10508 6316 10560 6322
rect 10508 6258 10560 6264
rect 9956 6248 10008 6254
rect 9956 6190 10008 6196
rect 10416 6248 10468 6254
rect 10416 6190 10468 6196
rect 10796 6186 10824 6854
rect 10888 6322 10916 7346
rect 10968 6860 11020 6866
rect 10968 6802 11020 6808
rect 10876 6316 10928 6322
rect 10876 6258 10928 6264
rect 10980 6202 11008 6802
rect 11256 6662 11284 8502
rect 11348 8090 11376 11194
rect 11428 8832 11480 8838
rect 11428 8774 11480 8780
rect 11440 8498 11468 8774
rect 11624 8634 11652 11194
rect 11794 9208 11850 9217
rect 11794 9143 11850 9152
rect 11612 8628 11664 8634
rect 11612 8570 11664 8576
rect 11428 8492 11480 8498
rect 11428 8434 11480 8440
rect 11520 8492 11572 8498
rect 11520 8434 11572 8440
rect 11336 8084 11388 8090
rect 11336 8026 11388 8032
rect 11428 6792 11480 6798
rect 11428 6734 11480 6740
rect 11244 6656 11296 6662
rect 11244 6598 11296 6604
rect 10784 6180 10836 6186
rect 10980 6174 11100 6202
rect 10784 6122 10836 6128
rect 11072 6118 11100 6174
rect 10140 6112 10192 6118
rect 10416 6112 10468 6118
rect 10192 6072 10416 6100
rect 10140 6054 10192 6060
rect 10416 6054 10468 6060
rect 11060 6112 11112 6118
rect 11060 6054 11112 6060
rect 11152 6112 11204 6118
rect 11152 6054 11204 6060
rect 11164 5778 11192 6054
rect 11440 5914 11468 6734
rect 11532 6662 11560 8434
rect 11520 6656 11572 6662
rect 11520 6598 11572 6604
rect 11808 6322 11836 9143
rect 11900 8090 11928 11194
rect 12070 8800 12126 8809
rect 12070 8735 12126 8744
rect 11980 8424 12032 8430
rect 11980 8366 12032 8372
rect 11888 8084 11940 8090
rect 11888 8026 11940 8032
rect 11992 6662 12020 8366
rect 12084 6798 12112 8735
rect 12176 8634 12204 11194
rect 12452 8634 12480 11194
rect 12532 9308 12584 9314
rect 12532 9250 12584 9256
rect 12164 8628 12216 8634
rect 12164 8570 12216 8576
rect 12440 8628 12492 8634
rect 12440 8570 12492 8576
rect 12544 8498 12572 9250
rect 12728 8634 12756 11194
rect 12808 9308 12860 9314
rect 12808 9250 12860 9256
rect 12716 8628 12768 8634
rect 12716 8570 12768 8576
rect 12820 8514 12848 9250
rect 13004 8634 13032 11194
rect 13280 8634 13308 11194
rect 13452 8832 13504 8838
rect 13452 8774 13504 8780
rect 12992 8628 13044 8634
rect 12992 8570 13044 8576
rect 13268 8628 13320 8634
rect 13268 8570 13320 8576
rect 12164 8492 12216 8498
rect 12164 8434 12216 8440
rect 12532 8492 12584 8498
rect 12532 8434 12584 8440
rect 12728 8486 12848 8514
rect 13360 8492 13412 8498
rect 12072 6792 12124 6798
rect 12072 6734 12124 6740
rect 11980 6656 12032 6662
rect 11980 6598 12032 6604
rect 11796 6316 11848 6322
rect 11796 6258 11848 6264
rect 12176 6186 12204 8434
rect 12624 7880 12676 7886
rect 12624 7822 12676 7828
rect 12636 7002 12664 7822
rect 12624 6996 12676 7002
rect 12624 6938 12676 6944
rect 12728 6390 12756 8486
rect 13360 8434 13412 8440
rect 12808 6792 12860 6798
rect 12808 6734 12860 6740
rect 12820 6390 12848 6734
rect 13372 6730 13400 8434
rect 13360 6724 13412 6730
rect 13360 6666 13412 6672
rect 13464 6662 13492 8774
rect 13556 8634 13584 11194
rect 13636 10056 13688 10062
rect 13636 9998 13688 10004
rect 13544 8628 13596 8634
rect 13544 8570 13596 8576
rect 13544 8424 13596 8430
rect 13544 8366 13596 8372
rect 13452 6656 13504 6662
rect 13452 6598 13504 6604
rect 12716 6384 12768 6390
rect 12438 6352 12494 6361
rect 12716 6326 12768 6332
rect 12808 6384 12860 6390
rect 12808 6326 12860 6332
rect 12438 6287 12494 6296
rect 12164 6180 12216 6186
rect 12164 6122 12216 6128
rect 11428 5908 11480 5914
rect 11428 5850 11480 5856
rect 11152 5772 11204 5778
rect 11152 5714 11204 5720
rect 6918 5199 6974 5208
rect 9864 5228 9916 5234
rect 4620 5160 4672 5166
rect 2870 5128 2926 5137
rect 4620 5102 4672 5108
rect 2870 5063 2926 5072
rect 1766 4992 1822 5001
rect 1766 4927 1822 4936
rect 1780 4593 1808 4927
rect 1950 4924 2258 4933
rect 1950 4922 1956 4924
rect 2012 4922 2036 4924
rect 2092 4922 2116 4924
rect 2172 4922 2196 4924
rect 2252 4922 2258 4924
rect 2012 4870 2014 4922
rect 2194 4870 2196 4922
rect 1950 4868 1956 4870
rect 2012 4868 2036 4870
rect 2092 4868 2116 4870
rect 2172 4868 2196 4870
rect 2252 4868 2258 4870
rect 1950 4859 2258 4868
rect 1766 4584 1822 4593
rect 1766 4519 1822 4528
rect 2884 4457 2912 5063
rect 2870 4448 2926 4457
rect 2870 4383 2926 4392
rect 3010 4380 3318 4389
rect 3010 4378 3016 4380
rect 3072 4378 3096 4380
rect 3152 4378 3176 4380
rect 3232 4378 3256 4380
rect 3312 4378 3318 4380
rect 3072 4326 3074 4378
rect 3254 4326 3256 4378
rect 3010 4324 3016 4326
rect 3072 4324 3096 4326
rect 3152 4324 3176 4326
rect 3232 4324 3256 4326
rect 3312 4324 3318 4326
rect 3010 4315 3318 4324
rect 6932 3942 6960 5199
rect 9864 5170 9916 5176
rect 7950 4924 8258 4933
rect 7950 4922 7956 4924
rect 8012 4922 8036 4924
rect 8092 4922 8116 4924
rect 8172 4922 8196 4924
rect 8252 4922 8258 4924
rect 8012 4870 8014 4922
rect 8194 4870 8196 4922
rect 7950 4868 7956 4870
rect 8012 4868 8036 4870
rect 8092 4868 8116 4870
rect 8172 4868 8196 4870
rect 8252 4868 8258 4870
rect 7950 4859 8258 4868
rect 9010 4380 9318 4389
rect 9010 4378 9016 4380
rect 9072 4378 9096 4380
rect 9152 4378 9176 4380
rect 9232 4378 9256 4380
rect 9312 4378 9318 4380
rect 9072 4326 9074 4378
rect 9254 4326 9256 4378
rect 9010 4324 9016 4326
rect 9072 4324 9096 4326
rect 9152 4324 9176 4326
rect 9232 4324 9256 4326
rect 9312 4324 9318 4326
rect 9010 4315 9318 4324
rect 12452 4146 12480 6287
rect 13556 5710 13584 8366
rect 13648 6118 13676 9998
rect 13726 9888 13782 9897
rect 13726 9823 13782 9832
rect 13740 8974 13768 9823
rect 13728 8968 13780 8974
rect 13728 8910 13780 8916
rect 13832 8616 13860 11194
rect 14108 9738 14136 11194
rect 14384 9761 14412 11194
rect 14660 10033 14688 11194
rect 14936 10849 14964 11194
rect 14922 10840 14978 10849
rect 14922 10775 14978 10784
rect 14646 10024 14702 10033
rect 14646 9959 14702 9968
rect 14016 9710 14136 9738
rect 14370 9752 14426 9761
rect 13912 8628 13964 8634
rect 13832 8588 13912 8616
rect 13912 8570 13964 8576
rect 14016 8294 14044 9710
rect 14370 9687 14426 9696
rect 14462 9480 14518 9489
rect 14462 9415 14518 9424
rect 14476 9081 14504 9415
rect 14462 9072 14518 9081
rect 14096 9036 14148 9042
rect 14462 9007 14518 9016
rect 14096 8978 14148 8984
rect 14108 8498 14136 8978
rect 15212 8922 15240 11194
rect 15488 9217 15516 11194
rect 15660 11144 15712 11150
rect 15660 11086 15712 11092
rect 15474 9208 15530 9217
rect 15474 9143 15530 9152
rect 15212 8894 15424 8922
rect 15010 8732 15318 8741
rect 15010 8730 15016 8732
rect 15072 8730 15096 8732
rect 15152 8730 15176 8732
rect 15232 8730 15256 8732
rect 15312 8730 15318 8732
rect 15072 8678 15074 8730
rect 15254 8678 15256 8730
rect 15010 8676 15016 8678
rect 15072 8676 15096 8678
rect 15152 8676 15176 8678
rect 15232 8676 15256 8678
rect 15312 8676 15318 8678
rect 15010 8667 15318 8676
rect 14096 8492 14148 8498
rect 14096 8434 14148 8440
rect 14004 8288 14056 8294
rect 14004 8230 14056 8236
rect 13950 8188 14258 8197
rect 13950 8186 13956 8188
rect 14012 8186 14036 8188
rect 14092 8186 14116 8188
rect 14172 8186 14196 8188
rect 14252 8186 14258 8188
rect 14012 8134 14014 8186
rect 14194 8134 14196 8186
rect 13950 8132 13956 8134
rect 14012 8132 14036 8134
rect 14092 8132 14116 8134
rect 14172 8132 14196 8134
rect 14252 8132 14258 8134
rect 13950 8123 14258 8132
rect 14830 8120 14886 8129
rect 14830 8055 14886 8064
rect 14372 7812 14424 7818
rect 14372 7754 14424 7760
rect 13950 7100 14258 7109
rect 13950 7098 13956 7100
rect 14012 7098 14036 7100
rect 14092 7098 14116 7100
rect 14172 7098 14196 7100
rect 14252 7098 14258 7100
rect 14012 7046 14014 7098
rect 14194 7046 14196 7098
rect 13950 7044 13956 7046
rect 14012 7044 14036 7046
rect 14092 7044 14116 7046
rect 14172 7044 14196 7046
rect 14252 7044 14258 7046
rect 13950 7035 14258 7044
rect 14384 7002 14412 7754
rect 14844 7721 14872 8055
rect 14830 7712 14886 7721
rect 14830 7647 14886 7656
rect 15010 7644 15318 7653
rect 15010 7642 15016 7644
rect 15072 7642 15096 7644
rect 15152 7642 15176 7644
rect 15232 7642 15256 7644
rect 15312 7642 15318 7644
rect 15072 7590 15074 7642
rect 15254 7590 15256 7642
rect 15010 7588 15016 7590
rect 15072 7588 15096 7590
rect 15152 7588 15176 7590
rect 15232 7588 15256 7590
rect 15312 7588 15318 7590
rect 15010 7579 15318 7588
rect 14372 6996 14424 7002
rect 14372 6938 14424 6944
rect 15010 6556 15318 6565
rect 15010 6554 15016 6556
rect 15072 6554 15096 6556
rect 15152 6554 15176 6556
rect 15232 6554 15256 6556
rect 15312 6554 15318 6556
rect 15072 6502 15074 6554
rect 15254 6502 15256 6554
rect 15010 6500 15016 6502
rect 15072 6500 15096 6502
rect 15152 6500 15176 6502
rect 15232 6500 15256 6502
rect 15312 6500 15318 6502
rect 15010 6491 15318 6500
rect 13636 6112 13688 6118
rect 13636 6054 13688 6060
rect 15292 6112 15344 6118
rect 15292 6054 15344 6060
rect 13950 6012 14258 6021
rect 13950 6010 13956 6012
rect 14012 6010 14036 6012
rect 14092 6010 14116 6012
rect 14172 6010 14196 6012
rect 14252 6010 14258 6012
rect 14012 5958 14014 6010
rect 14194 5958 14196 6010
rect 13950 5956 13956 5958
rect 14012 5956 14036 5958
rect 14092 5956 14116 5958
rect 14172 5956 14196 5958
rect 14252 5956 14258 5958
rect 13950 5947 14258 5956
rect 15304 5914 15332 6054
rect 15292 5908 15344 5914
rect 15292 5850 15344 5856
rect 13726 5808 13782 5817
rect 13726 5743 13782 5752
rect 13544 5704 13596 5710
rect 13544 5646 13596 5652
rect 12440 4140 12492 4146
rect 12440 4082 12492 4088
rect 9402 4040 9458 4049
rect 7012 4004 7064 4010
rect 9402 3975 9458 3984
rect 13634 4040 13690 4049
rect 13634 3975 13690 3984
rect 7012 3946 7064 3952
rect 6920 3936 6972 3942
rect 6920 3878 6972 3884
rect 1950 3836 2258 3845
rect 1950 3834 1956 3836
rect 2012 3834 2036 3836
rect 2092 3834 2116 3836
rect 2172 3834 2196 3836
rect 2252 3834 2258 3836
rect 2012 3782 2014 3834
rect 2194 3782 2196 3834
rect 1950 3780 1956 3782
rect 2012 3780 2036 3782
rect 2092 3780 2116 3782
rect 2172 3780 2196 3782
rect 2252 3780 2258 3782
rect 1950 3771 2258 3780
rect 7024 3738 7052 3946
rect 7950 3836 8258 3845
rect 7950 3834 7956 3836
rect 8012 3834 8036 3836
rect 8092 3834 8116 3836
rect 8172 3834 8196 3836
rect 8252 3834 8258 3836
rect 8012 3782 8014 3834
rect 8194 3782 8196 3834
rect 7950 3780 7956 3782
rect 8012 3780 8036 3782
rect 8092 3780 8116 3782
rect 8172 3780 8196 3782
rect 8252 3780 8258 3782
rect 7950 3771 8258 3780
rect 7012 3732 7064 3738
rect 7012 3674 7064 3680
rect 9416 3670 9444 3975
rect 10692 3936 10744 3942
rect 10692 3878 10744 3884
rect 9588 3732 9640 3738
rect 9588 3674 9640 3680
rect 9404 3664 9456 3670
rect 9404 3606 9456 3612
rect 1308 3596 1360 3602
rect 1308 3538 1360 3544
rect 7472 3596 7524 3602
rect 7472 3538 7524 3544
rect 9496 3596 9548 3602
rect 9496 3538 9548 3544
rect 1124 3528 1176 3534
rect 1124 3470 1176 3476
rect 1766 3496 1822 3505
rect 1136 1465 1164 3470
rect 1308 3460 1360 3466
rect 1766 3431 1822 3440
rect 1308 3402 1360 3408
rect 1320 2553 1348 3402
rect 1780 2825 1808 3431
rect 4896 3392 4948 3398
rect 1950 3360 2006 3369
rect 4896 3334 4948 3340
rect 1950 3295 2006 3304
rect 1964 2961 1992 3295
rect 3010 3292 3318 3301
rect 3010 3290 3016 3292
rect 3072 3290 3096 3292
rect 3152 3290 3176 3292
rect 3232 3290 3256 3292
rect 3312 3290 3318 3292
rect 3072 3238 3074 3290
rect 3254 3238 3256 3290
rect 3010 3236 3016 3238
rect 3072 3236 3096 3238
rect 3152 3236 3176 3238
rect 3232 3236 3256 3238
rect 3312 3236 3318 3238
rect 3010 3227 3318 3236
rect 4344 3188 4396 3194
rect 4344 3130 4396 3136
rect 1950 2952 2006 2961
rect 1950 2887 2006 2896
rect 1766 2816 1822 2825
rect 1766 2751 1822 2760
rect 1950 2748 2258 2757
rect 1950 2746 1956 2748
rect 2012 2746 2036 2748
rect 2092 2746 2116 2748
rect 2172 2746 2196 2748
rect 2252 2746 2258 2748
rect 2012 2694 2014 2746
rect 2194 2694 2196 2746
rect 1950 2692 1956 2694
rect 2012 2692 2036 2694
rect 2092 2692 2116 2694
rect 2172 2692 2196 2694
rect 2252 2692 2258 2694
rect 1950 2683 2258 2692
rect 1306 2544 1362 2553
rect 1306 2479 1362 2488
rect 3010 2204 3318 2213
rect 3010 2202 3016 2204
rect 3072 2202 3096 2204
rect 3152 2202 3176 2204
rect 3232 2202 3256 2204
rect 3312 2202 3318 2204
rect 3072 2150 3074 2202
rect 3254 2150 3256 2202
rect 3010 2148 3016 2150
rect 3072 2148 3096 2150
rect 3152 2148 3176 2150
rect 3232 2148 3256 2150
rect 3312 2148 3318 2150
rect 3010 2139 3318 2148
rect 1122 1456 1178 1465
rect 1122 1391 1178 1400
rect 2780 196 2832 202
rect 2780 138 2832 144
rect 1228 66 1348 82
rect 1228 60 1360 66
rect 1228 56 1308 60
rect 1214 54 1308 56
rect 1214 0 1270 54
rect 2792 56 2820 138
rect 4356 56 4384 3130
rect 4908 2446 4936 3334
rect 5908 3052 5960 3058
rect 5908 2994 5960 3000
rect 4896 2440 4948 2446
rect 4896 2382 4948 2388
rect 5920 56 5948 2994
rect 7484 56 7512 3538
rect 8392 3392 8444 3398
rect 8392 3334 8444 3340
rect 7950 2748 8258 2757
rect 7950 2746 7956 2748
rect 8012 2746 8036 2748
rect 8092 2746 8116 2748
rect 8172 2746 8196 2748
rect 8252 2746 8258 2748
rect 8012 2694 8014 2746
rect 8194 2694 8196 2746
rect 7950 2692 7956 2694
rect 8012 2692 8036 2694
rect 8092 2692 8116 2694
rect 8172 2692 8196 2694
rect 8252 2692 8258 2694
rect 7950 2683 8258 2692
rect 8404 2378 8432 3334
rect 9010 3292 9318 3301
rect 9010 3290 9016 3292
rect 9072 3290 9096 3292
rect 9152 3290 9176 3292
rect 9232 3290 9256 3292
rect 9312 3290 9318 3292
rect 9072 3238 9074 3290
rect 9254 3238 9256 3290
rect 9010 3236 9016 3238
rect 9072 3236 9096 3238
rect 9152 3236 9176 3238
rect 9232 3236 9256 3238
rect 9312 3236 9318 3238
rect 9010 3227 9318 3236
rect 9404 3120 9456 3126
rect 9404 3062 9456 3068
rect 9416 2417 9444 3062
rect 9402 2408 9458 2417
rect 8392 2372 8444 2378
rect 9402 2343 9458 2352
rect 8392 2314 8444 2320
rect 9010 2204 9318 2213
rect 9010 2202 9016 2204
rect 9072 2202 9096 2204
rect 9152 2202 9176 2204
rect 9232 2202 9256 2204
rect 9312 2202 9318 2204
rect 9072 2150 9074 2202
rect 9254 2150 9256 2202
rect 9010 2148 9016 2150
rect 9072 2148 9096 2150
rect 9152 2148 9176 2150
rect 9232 2148 9256 2150
rect 9312 2148 9318 2150
rect 9010 2139 9318 2148
rect 9508 1737 9536 3538
rect 9600 2009 9628 3674
rect 10704 3534 10732 3878
rect 10692 3528 10744 3534
rect 10692 3470 10744 3476
rect 12072 3528 12124 3534
rect 12072 3470 12124 3476
rect 10600 3392 10652 3398
rect 10600 3334 10652 3340
rect 11520 3392 11572 3398
rect 11520 3334 11572 3340
rect 10612 2922 10640 3334
rect 10600 2916 10652 2922
rect 10600 2858 10652 2864
rect 11532 2514 11560 3334
rect 12084 3126 12112 3470
rect 12164 3392 12216 3398
rect 12164 3334 12216 3340
rect 12440 3392 12492 3398
rect 12440 3334 12492 3340
rect 12072 3120 12124 3126
rect 12072 3062 12124 3068
rect 12176 2582 12204 3334
rect 12452 2650 12480 3334
rect 13648 2774 13676 3975
rect 13740 3670 13768 5743
rect 15010 5468 15318 5477
rect 15010 5466 15016 5468
rect 15072 5466 15096 5468
rect 15152 5466 15176 5468
rect 15232 5466 15256 5468
rect 15312 5466 15318 5468
rect 15072 5414 15074 5466
rect 15254 5414 15256 5466
rect 15010 5412 15016 5414
rect 15072 5412 15096 5414
rect 15152 5412 15176 5414
rect 15232 5412 15256 5414
rect 15312 5412 15318 5414
rect 15010 5403 15318 5412
rect 15396 5302 15424 8894
rect 15568 8900 15620 8906
rect 15568 8842 15620 8848
rect 15580 6662 15608 8842
rect 15672 6798 15700 11086
rect 15764 8786 15792 11194
rect 15764 8758 15884 8786
rect 15660 6792 15712 6798
rect 15660 6734 15712 6740
rect 15752 6792 15804 6798
rect 15752 6734 15804 6740
rect 15568 6656 15620 6662
rect 15568 6598 15620 6604
rect 15764 5778 15792 6734
rect 15856 6458 15884 8758
rect 15844 6452 15896 6458
rect 15844 6394 15896 6400
rect 16040 6225 16068 11194
rect 16118 9344 16174 9353
rect 16118 9279 16174 9288
rect 16132 6798 16160 9279
rect 16316 8514 16344 11194
rect 16316 8486 16436 8514
rect 16210 6896 16266 6905
rect 16210 6831 16266 6840
rect 16120 6792 16172 6798
rect 16120 6734 16172 6740
rect 16026 6216 16082 6225
rect 16026 6151 16082 6160
rect 15752 5772 15804 5778
rect 15752 5714 15804 5720
rect 16224 5710 16252 6831
rect 16304 6724 16356 6730
rect 16304 6666 16356 6672
rect 16316 6458 16344 6666
rect 16304 6452 16356 6458
rect 16304 6394 16356 6400
rect 16408 5846 16436 8486
rect 16592 8430 16620 11194
rect 16868 8514 16896 11194
rect 16776 8486 16896 8514
rect 16948 8560 17000 8566
rect 16948 8502 17000 8508
rect 16580 8424 16632 8430
rect 16580 8366 16632 8372
rect 16670 7848 16726 7857
rect 16670 7783 16726 7792
rect 16488 7744 16540 7750
rect 16488 7686 16540 7692
rect 16500 6730 16528 7686
rect 16580 7336 16632 7342
rect 16580 7278 16632 7284
rect 16592 7002 16620 7278
rect 16580 6996 16632 7002
rect 16580 6938 16632 6944
rect 16684 6798 16712 7783
rect 16672 6792 16724 6798
rect 16672 6734 16724 6740
rect 16488 6724 16540 6730
rect 16488 6666 16540 6672
rect 16776 5914 16804 8486
rect 16856 7472 16908 7478
rect 16856 7414 16908 7420
rect 16868 7002 16896 7414
rect 16856 6996 16908 7002
rect 16856 6938 16908 6944
rect 16764 5908 16816 5914
rect 16764 5850 16816 5856
rect 16396 5840 16448 5846
rect 16396 5782 16448 5788
rect 16212 5704 16264 5710
rect 16212 5646 16264 5652
rect 15384 5296 15436 5302
rect 16960 5250 16988 8502
rect 17144 5710 17172 11194
rect 17420 7274 17448 11194
rect 17500 8356 17552 8362
rect 17500 8298 17552 8304
rect 17408 7268 17460 7274
rect 17408 7210 17460 7216
rect 17512 6662 17540 8298
rect 17696 7206 17724 11194
rect 17972 9246 18000 11194
rect 18248 9330 18276 11194
rect 18156 9302 18276 9330
rect 17960 9240 18012 9246
rect 17960 9182 18012 9188
rect 17960 8900 18012 8906
rect 17960 8842 18012 8848
rect 17684 7200 17736 7206
rect 17684 7142 17736 7148
rect 17684 6792 17736 6798
rect 17684 6734 17736 6740
rect 17500 6656 17552 6662
rect 17500 6598 17552 6604
rect 17696 6118 17724 6734
rect 17592 6112 17644 6118
rect 17592 6054 17644 6060
rect 17684 6112 17736 6118
rect 17684 6054 17736 6060
rect 17604 5914 17632 6054
rect 17592 5908 17644 5914
rect 17592 5850 17644 5856
rect 17132 5704 17184 5710
rect 17132 5646 17184 5652
rect 15384 5238 15436 5244
rect 16868 5222 16988 5250
rect 13950 4924 14258 4933
rect 13950 4922 13956 4924
rect 14012 4922 14036 4924
rect 14092 4922 14116 4924
rect 14172 4922 14196 4924
rect 14252 4922 14258 4924
rect 14012 4870 14014 4922
rect 14194 4870 14196 4922
rect 13950 4868 13956 4870
rect 14012 4868 14036 4870
rect 14092 4868 14116 4870
rect 14172 4868 14196 4870
rect 14252 4868 14258 4870
rect 13950 4859 14258 4868
rect 13820 4820 13872 4826
rect 13820 4762 13872 4768
rect 13832 3942 13860 4762
rect 15660 4752 15712 4758
rect 15660 4694 15712 4700
rect 14922 4584 14978 4593
rect 14922 4519 14978 4528
rect 13820 3936 13872 3942
rect 13820 3878 13872 3884
rect 13950 3836 14258 3845
rect 13950 3834 13956 3836
rect 14012 3834 14036 3836
rect 14092 3834 14116 3836
rect 14172 3834 14196 3836
rect 14252 3834 14258 3836
rect 14012 3782 14014 3834
rect 14194 3782 14196 3834
rect 13950 3780 13956 3782
rect 14012 3780 14036 3782
rect 14092 3780 14116 3782
rect 14172 3780 14196 3782
rect 14252 3780 14258 3782
rect 13950 3771 14258 3780
rect 14936 3738 14964 4519
rect 15010 4380 15318 4389
rect 15010 4378 15016 4380
rect 15072 4378 15096 4380
rect 15152 4378 15176 4380
rect 15232 4378 15256 4380
rect 15312 4378 15318 4380
rect 15072 4326 15074 4378
rect 15254 4326 15256 4378
rect 15010 4324 15016 4326
rect 15072 4324 15096 4326
rect 15152 4324 15176 4326
rect 15232 4324 15256 4326
rect 15312 4324 15318 4326
rect 15010 4315 15318 4324
rect 15382 3904 15438 3913
rect 15382 3839 15438 3848
rect 14924 3732 14976 3738
rect 14924 3674 14976 3680
rect 13728 3664 13780 3670
rect 13728 3606 13780 3612
rect 14556 3528 14608 3534
rect 14556 3470 14608 3476
rect 14568 3194 14596 3470
rect 15010 3292 15318 3301
rect 15010 3290 15016 3292
rect 15072 3290 15096 3292
rect 15152 3290 15176 3292
rect 15232 3290 15256 3292
rect 15312 3290 15318 3292
rect 15072 3238 15074 3290
rect 15254 3238 15256 3290
rect 15010 3236 15016 3238
rect 15072 3236 15096 3238
rect 15152 3236 15176 3238
rect 15232 3236 15256 3238
rect 15312 3236 15318 3238
rect 15010 3227 15318 3236
rect 14556 3188 14608 3194
rect 14556 3130 14608 3136
rect 13648 2746 13768 2774
rect 12440 2644 12492 2650
rect 12440 2586 12492 2592
rect 12164 2576 12216 2582
rect 12164 2518 12216 2524
rect 11520 2508 11572 2514
rect 11520 2450 11572 2456
rect 12164 2100 12216 2106
rect 12164 2042 12216 2048
rect 9586 2000 9642 2009
rect 9586 1935 9642 1944
rect 9494 1728 9550 1737
rect 9494 1663 9550 1672
rect 9034 232 9090 241
rect 9034 167 9090 176
rect 9048 56 9076 167
rect 10598 96 10654 105
rect 1308 2 1360 8
rect 2778 0 2834 56
rect 4342 0 4398 56
rect 5906 0 5962 56
rect 7470 0 7526 56
rect 9034 0 9090 56
rect 12176 56 12204 2042
rect 13740 56 13768 2746
rect 13950 2748 14258 2757
rect 13950 2746 13956 2748
rect 14012 2746 14036 2748
rect 14092 2746 14116 2748
rect 14172 2746 14196 2748
rect 14252 2746 14258 2748
rect 14012 2694 14014 2746
rect 14194 2694 14196 2746
rect 13950 2692 13956 2694
rect 14012 2692 14036 2694
rect 14092 2692 14116 2694
rect 14172 2692 14196 2694
rect 14252 2692 14258 2694
rect 13950 2683 14258 2692
rect 15010 2204 15318 2213
rect 15010 2202 15016 2204
rect 15072 2202 15096 2204
rect 15152 2202 15176 2204
rect 15232 2202 15256 2204
rect 15312 2202 15318 2204
rect 15072 2150 15074 2202
rect 15254 2150 15256 2202
rect 15010 2148 15016 2150
rect 15072 2148 15096 2150
rect 15152 2148 15176 2150
rect 15232 2148 15256 2150
rect 15312 2148 15318 2150
rect 15010 2139 15318 2148
rect 15396 1986 15424 3839
rect 15672 3738 15700 4694
rect 16396 4072 16448 4078
rect 16396 4014 16448 4020
rect 15936 3936 15988 3942
rect 15936 3878 15988 3884
rect 15948 3738 15976 3878
rect 15568 3732 15620 3738
rect 15568 3674 15620 3680
rect 15660 3732 15712 3738
rect 15660 3674 15712 3680
rect 15936 3732 15988 3738
rect 15936 3674 15988 3680
rect 15580 3534 15608 3674
rect 15568 3528 15620 3534
rect 15568 3470 15620 3476
rect 16408 3466 16436 4014
rect 16488 3732 16540 3738
rect 16488 3674 16540 3680
rect 16500 3505 16528 3674
rect 16868 3534 16896 5222
rect 17866 5128 17922 5137
rect 17866 5063 17922 5072
rect 16948 4548 17000 4554
rect 16948 4490 17000 4496
rect 16856 3528 16908 3534
rect 16486 3496 16542 3505
rect 16396 3460 16448 3466
rect 16856 3470 16908 3476
rect 16486 3431 16542 3440
rect 16396 3402 16448 3408
rect 16580 3392 16632 3398
rect 16580 3334 16632 3340
rect 16672 3392 16724 3398
rect 16672 3334 16724 3340
rect 16856 3392 16908 3398
rect 16856 3334 16908 3340
rect 16592 3058 16620 3334
rect 16580 3052 16632 3058
rect 16580 2994 16632 3000
rect 16684 2961 16712 3334
rect 16868 3097 16896 3334
rect 16854 3088 16910 3097
rect 16854 3023 16910 3032
rect 16670 2952 16726 2961
rect 16670 2887 16726 2896
rect 16960 2258 16988 4490
rect 17880 4146 17908 5063
rect 17868 4140 17920 4146
rect 17868 4082 17920 4088
rect 17972 3738 18000 8842
rect 18156 7313 18184 9302
rect 18236 9104 18288 9110
rect 18236 9046 18288 9052
rect 18142 7304 18198 7313
rect 18142 7239 18198 7248
rect 18248 6662 18276 9046
rect 18524 8129 18552 11194
rect 18800 9450 18828 11194
rect 19076 10441 19104 11194
rect 19062 10432 19118 10441
rect 19062 10367 19118 10376
rect 19352 10062 19380 11194
rect 19340 10056 19392 10062
rect 19340 9998 19392 10004
rect 18788 9444 18840 9450
rect 18788 9386 18840 9392
rect 19248 9172 19300 9178
rect 19248 9114 19300 9120
rect 18510 8120 18566 8129
rect 18510 8055 18566 8064
rect 19260 7002 19288 9114
rect 19340 8016 19392 8022
rect 19340 7958 19392 7964
rect 19248 6996 19300 7002
rect 19248 6938 19300 6944
rect 19352 6798 19380 7958
rect 18420 6792 18472 6798
rect 18420 6734 18472 6740
rect 19340 6792 19392 6798
rect 19340 6734 19392 6740
rect 18236 6656 18288 6662
rect 18236 6598 18288 6604
rect 18432 6186 18460 6734
rect 19524 6656 19576 6662
rect 19524 6598 19576 6604
rect 19536 6254 19564 6598
rect 19628 6322 19656 11194
rect 19904 9194 19932 11194
rect 19720 9166 19932 9194
rect 19720 6769 19748 9166
rect 20180 9058 20208 11194
rect 19812 9030 20208 9058
rect 19706 6760 19762 6769
rect 19706 6695 19762 6704
rect 19812 6458 19840 9030
rect 20456 8945 20484 11194
rect 20732 9602 20760 11194
rect 20732 9574 20852 9602
rect 20718 9072 20774 9081
rect 20718 9007 20774 9016
rect 20442 8936 20498 8945
rect 20442 8871 20498 8880
rect 19950 8188 20258 8197
rect 19950 8186 19956 8188
rect 20012 8186 20036 8188
rect 20092 8186 20116 8188
rect 20172 8186 20196 8188
rect 20252 8186 20258 8188
rect 20012 8134 20014 8186
rect 20194 8134 20196 8186
rect 19950 8132 19956 8134
rect 20012 8132 20036 8134
rect 20092 8132 20116 8134
rect 20172 8132 20196 8134
rect 20252 8132 20258 8134
rect 19950 8123 20258 8132
rect 19950 7100 20258 7109
rect 19950 7098 19956 7100
rect 20012 7098 20036 7100
rect 20092 7098 20116 7100
rect 20172 7098 20196 7100
rect 20252 7098 20258 7100
rect 20012 7046 20014 7098
rect 20194 7046 20196 7098
rect 19950 7044 19956 7046
rect 20012 7044 20036 7046
rect 20092 7044 20116 7046
rect 20172 7044 20196 7046
rect 20252 7044 20258 7046
rect 19950 7035 20258 7044
rect 20732 6866 20760 9007
rect 20824 7954 20852 9574
rect 21008 9314 21036 11194
rect 20996 9308 21048 9314
rect 20996 9250 21048 9256
rect 20902 9208 20958 9217
rect 20902 9143 20958 9152
rect 20812 7948 20864 7954
rect 20812 7890 20864 7896
rect 20812 7404 20864 7410
rect 20812 7346 20864 7352
rect 20824 7002 20852 7346
rect 20812 6996 20864 7002
rect 20812 6938 20864 6944
rect 20720 6860 20772 6866
rect 20720 6802 20772 6808
rect 19984 6792 20036 6798
rect 20916 6780 20944 9143
rect 21284 8838 21312 11194
rect 21560 9058 21588 11194
rect 21638 9480 21694 9489
rect 21638 9415 21694 9424
rect 21376 9030 21588 9058
rect 21272 8832 21324 8838
rect 21272 8774 21324 8780
rect 21010 8732 21318 8741
rect 21010 8730 21016 8732
rect 21072 8730 21096 8732
rect 21152 8730 21176 8732
rect 21232 8730 21256 8732
rect 21312 8730 21318 8732
rect 21072 8678 21074 8730
rect 21254 8678 21256 8730
rect 21010 8676 21016 8678
rect 21072 8676 21096 8678
rect 21152 8676 21176 8678
rect 21232 8676 21256 8678
rect 21312 8676 21318 8678
rect 21010 8667 21318 8676
rect 21010 7644 21318 7653
rect 21010 7642 21016 7644
rect 21072 7642 21096 7644
rect 21152 7642 21176 7644
rect 21232 7642 21256 7644
rect 21312 7642 21318 7644
rect 21072 7590 21074 7642
rect 21254 7590 21256 7642
rect 21010 7588 21016 7590
rect 21072 7588 21096 7590
rect 21152 7588 21176 7590
rect 21232 7588 21256 7590
rect 21312 7588 21318 7590
rect 21010 7579 21318 7588
rect 20996 6792 21048 6798
rect 20916 6752 20996 6780
rect 19984 6734 20036 6740
rect 20996 6734 21048 6740
rect 19996 6458 20024 6734
rect 20812 6656 20864 6662
rect 20812 6598 20864 6604
rect 19800 6452 19852 6458
rect 19800 6394 19852 6400
rect 19984 6452 20036 6458
rect 19984 6394 20036 6400
rect 19616 6316 19668 6322
rect 19616 6258 19668 6264
rect 19524 6248 19576 6254
rect 19524 6190 19576 6196
rect 18420 6180 18472 6186
rect 18420 6122 18472 6128
rect 19950 6012 20258 6021
rect 19950 6010 19956 6012
rect 20012 6010 20036 6012
rect 20092 6010 20116 6012
rect 20172 6010 20196 6012
rect 20252 6010 20258 6012
rect 20012 5958 20014 6010
rect 20194 5958 20196 6010
rect 19950 5956 19956 5958
rect 20012 5956 20036 5958
rect 20092 5956 20116 5958
rect 20172 5956 20196 5958
rect 20252 5956 20258 5958
rect 19950 5947 20258 5956
rect 20824 5914 20852 6598
rect 21010 6556 21318 6565
rect 21010 6554 21016 6556
rect 21072 6554 21096 6556
rect 21152 6554 21176 6556
rect 21232 6554 21256 6556
rect 21312 6554 21318 6556
rect 21072 6502 21074 6554
rect 21254 6502 21256 6554
rect 21010 6500 21016 6502
rect 21072 6500 21096 6502
rect 21152 6500 21176 6502
rect 21232 6500 21256 6502
rect 21312 6500 21318 6502
rect 21010 6491 21318 6500
rect 21376 6390 21404 9030
rect 21548 8832 21600 8838
rect 21548 8774 21600 8780
rect 21456 7812 21508 7818
rect 21456 7754 21508 7760
rect 21364 6384 21416 6390
rect 21364 6326 21416 6332
rect 20812 5908 20864 5914
rect 20812 5850 20864 5856
rect 21364 5908 21416 5914
rect 21364 5850 21416 5856
rect 20352 5704 20404 5710
rect 20352 5646 20404 5652
rect 19064 5296 19116 5302
rect 19064 5238 19116 5244
rect 18420 5228 18472 5234
rect 18420 5170 18472 5176
rect 18142 4720 18198 4729
rect 18142 4655 18198 4664
rect 18156 3738 18184 4655
rect 17960 3732 18012 3738
rect 17960 3674 18012 3680
rect 18144 3732 18196 3738
rect 18144 3674 18196 3680
rect 17408 3664 17460 3670
rect 17406 3632 17408 3641
rect 17460 3632 17462 3641
rect 17406 3567 17462 3576
rect 17776 3528 17828 3534
rect 17776 3470 17828 3476
rect 17224 3392 17276 3398
rect 17224 3334 17276 3340
rect 17500 3392 17552 3398
rect 17500 3334 17552 3340
rect 17236 3126 17264 3334
rect 17512 3194 17540 3334
rect 17500 3188 17552 3194
rect 17500 3130 17552 3136
rect 17224 3120 17276 3126
rect 17224 3062 17276 3068
rect 17788 3058 17816 3470
rect 17776 3052 17828 3058
rect 17776 2994 17828 3000
rect 15304 1958 15424 1986
rect 16868 2230 16988 2258
rect 15304 56 15332 1958
rect 16868 56 16896 2230
rect 18432 56 18460 5170
rect 19076 3738 19104 5238
rect 19950 4924 20258 4933
rect 19950 4922 19956 4924
rect 20012 4922 20036 4924
rect 20092 4922 20116 4924
rect 20172 4922 20196 4924
rect 20252 4922 20258 4924
rect 20012 4870 20014 4922
rect 20194 4870 20196 4922
rect 19950 4868 19956 4870
rect 20012 4868 20036 4870
rect 20092 4868 20116 4870
rect 20172 4868 20196 4870
rect 20252 4868 20258 4870
rect 19950 4859 20258 4868
rect 19432 4276 19484 4282
rect 19432 4218 19484 4224
rect 19248 4140 19300 4146
rect 19248 4082 19300 4088
rect 18880 3732 18932 3738
rect 18880 3674 18932 3680
rect 19064 3732 19116 3738
rect 19064 3674 19116 3680
rect 18892 3534 18920 3674
rect 19260 3534 19288 4082
rect 19444 3738 19472 4218
rect 19522 4176 19578 4185
rect 19522 4111 19578 4120
rect 19536 3738 19564 4111
rect 19800 3936 19852 3942
rect 19800 3878 19852 3884
rect 19432 3732 19484 3738
rect 19432 3674 19484 3680
rect 19524 3732 19576 3738
rect 19524 3674 19576 3680
rect 19536 3534 19564 3674
rect 19812 3670 19840 3878
rect 19950 3836 20258 3845
rect 19950 3834 19956 3836
rect 20012 3834 20036 3836
rect 20092 3834 20116 3836
rect 20172 3834 20196 3836
rect 20252 3834 20258 3836
rect 20012 3782 20014 3834
rect 20194 3782 20196 3834
rect 19950 3780 19956 3782
rect 20012 3780 20036 3782
rect 20092 3780 20116 3782
rect 20172 3780 20196 3782
rect 20252 3780 20258 3782
rect 19950 3771 20258 3780
rect 19800 3664 19852 3670
rect 19800 3606 19852 3612
rect 18880 3528 18932 3534
rect 18510 3496 18566 3505
rect 18880 3470 18932 3476
rect 19248 3528 19300 3534
rect 19248 3470 19300 3476
rect 19524 3528 19576 3534
rect 19524 3470 19576 3476
rect 18510 3431 18566 3440
rect 18524 3398 18552 3431
rect 19260 3398 19288 3470
rect 18512 3392 18564 3398
rect 18512 3334 18564 3340
rect 18788 3392 18840 3398
rect 18788 3334 18840 3340
rect 19248 3392 19300 3398
rect 19248 3334 19300 3340
rect 18800 3058 18828 3334
rect 18788 3052 18840 3058
rect 18788 2994 18840 3000
rect 19950 2748 20258 2757
rect 19950 2746 19956 2748
rect 20012 2746 20036 2748
rect 20092 2746 20116 2748
rect 20172 2746 20196 2748
rect 20252 2746 20258 2748
rect 20012 2694 20014 2746
rect 20194 2694 20196 2746
rect 19950 2692 19956 2694
rect 20012 2692 20036 2694
rect 20092 2692 20116 2694
rect 20172 2692 20196 2694
rect 20252 2692 20258 2694
rect 19950 2683 20258 2692
rect 19996 56 20116 82
rect 10598 0 10654 40
rect 12162 0 12218 56
rect 13726 0 13782 56
rect 15290 0 15346 56
rect 16854 0 16910 56
rect 18418 0 18474 56
rect 19982 54 20116 56
rect 19982 0 20038 54
rect 20088 42 20116 54
rect 20364 42 20392 5646
rect 21010 5468 21318 5477
rect 21010 5466 21016 5468
rect 21072 5466 21096 5468
rect 21152 5466 21176 5468
rect 21232 5466 21256 5468
rect 21312 5466 21318 5468
rect 21072 5414 21074 5466
rect 21254 5414 21256 5466
rect 21010 5412 21016 5414
rect 21072 5412 21096 5414
rect 21152 5412 21176 5414
rect 21232 5412 21256 5414
rect 21312 5412 21318 5414
rect 21010 5403 21318 5412
rect 20904 5160 20956 5166
rect 20904 5102 20956 5108
rect 20916 4146 20944 5102
rect 21010 4380 21318 4389
rect 21010 4378 21016 4380
rect 21072 4378 21096 4380
rect 21152 4378 21176 4380
rect 21232 4378 21256 4380
rect 21312 4378 21318 4380
rect 21072 4326 21074 4378
rect 21254 4326 21256 4378
rect 21010 4324 21016 4326
rect 21072 4324 21096 4326
rect 21152 4324 21176 4326
rect 21232 4324 21256 4326
rect 21312 4324 21318 4326
rect 21010 4315 21318 4324
rect 20904 4140 20956 4146
rect 20904 4082 20956 4088
rect 21376 3942 21404 5850
rect 21468 5370 21496 7754
rect 21560 6662 21588 8774
rect 21652 6798 21680 9415
rect 21732 9036 21784 9042
rect 21732 8978 21784 8984
rect 21640 6792 21692 6798
rect 21640 6734 21692 6740
rect 21548 6656 21600 6662
rect 21548 6598 21600 6604
rect 21640 6656 21692 6662
rect 21640 6598 21692 6604
rect 21652 6390 21680 6598
rect 21640 6384 21692 6390
rect 21640 6326 21692 6332
rect 21548 6316 21600 6322
rect 21548 6258 21600 6264
rect 21456 5364 21508 5370
rect 21456 5306 21508 5312
rect 21364 3936 21416 3942
rect 21364 3878 21416 3884
rect 21010 3292 21318 3301
rect 21010 3290 21016 3292
rect 21072 3290 21096 3292
rect 21152 3290 21176 3292
rect 21232 3290 21256 3292
rect 21312 3290 21318 3292
rect 21072 3238 21074 3290
rect 21254 3238 21256 3290
rect 21010 3236 21016 3238
rect 21072 3236 21096 3238
rect 21152 3236 21176 3238
rect 21232 3236 21256 3238
rect 21312 3236 21318 3238
rect 21010 3227 21318 3236
rect 21010 2204 21318 2213
rect 21010 2202 21016 2204
rect 21072 2202 21096 2204
rect 21152 2202 21176 2204
rect 21232 2202 21256 2204
rect 21312 2202 21318 2204
rect 21072 2150 21074 2202
rect 21254 2150 21256 2202
rect 21010 2148 21016 2150
rect 21072 2148 21096 2150
rect 21152 2148 21176 2150
rect 21232 2148 21256 2150
rect 21312 2148 21318 2150
rect 21010 2139 21318 2148
rect 21560 56 21588 6258
rect 21744 5846 21772 8978
rect 21836 7002 21864 11194
rect 22112 11150 22140 11194
rect 22100 11144 22152 11150
rect 22100 11086 22152 11092
rect 22388 9058 22416 11194
rect 22664 9081 22692 11194
rect 22296 9030 22416 9058
rect 22650 9072 22706 9081
rect 21824 6996 21876 7002
rect 21824 6938 21876 6944
rect 22296 6914 22324 9030
rect 22650 9007 22706 9016
rect 22376 8424 22428 8430
rect 22376 8366 22428 8372
rect 22112 6886 22324 6914
rect 22112 5846 22140 6886
rect 22192 6656 22244 6662
rect 22192 6598 22244 6604
rect 22204 6118 22232 6598
rect 22192 6112 22244 6118
rect 22192 6054 22244 6060
rect 22284 6112 22336 6118
rect 22284 6054 22336 6060
rect 22296 5846 22324 6054
rect 21732 5840 21784 5846
rect 21732 5782 21784 5788
rect 22100 5840 22152 5846
rect 22100 5782 22152 5788
rect 22284 5840 22336 5846
rect 22284 5782 22336 5788
rect 21824 3528 21876 3534
rect 21824 3470 21876 3476
rect 22192 3528 22244 3534
rect 22192 3470 22244 3476
rect 21836 66 21864 3470
rect 22204 134 22232 3470
rect 22388 3398 22416 8366
rect 22836 6860 22888 6866
rect 22836 6802 22888 6808
rect 22848 6769 22876 6802
rect 22834 6760 22890 6769
rect 22834 6695 22890 6704
rect 22940 6662 22968 11194
rect 23110 8256 23166 8265
rect 23110 8191 23166 8200
rect 23124 7546 23152 8191
rect 23112 7540 23164 7546
rect 23112 7482 23164 7488
rect 23112 7404 23164 7410
rect 23112 7346 23164 7352
rect 22928 6656 22980 6662
rect 22928 6598 22980 6604
rect 22468 3528 22520 3534
rect 22468 3470 22520 3476
rect 22376 3392 22428 3398
rect 22376 3334 22428 3340
rect 22480 241 22508 3470
rect 22466 232 22522 241
rect 22466 167 22522 176
rect 22192 128 22244 134
rect 22192 70 22244 76
rect 21824 60 21876 66
rect 20088 14 20392 42
rect 21546 0 21602 56
rect 23124 56 23152 7346
rect 23216 6186 23244 11194
rect 23492 9738 23520 11194
rect 23492 9710 23612 9738
rect 23480 9104 23532 9110
rect 23480 9046 23532 9052
rect 23388 8356 23440 8362
rect 23388 8298 23440 8304
rect 23296 6792 23348 6798
rect 23296 6734 23348 6740
rect 23308 6322 23336 6734
rect 23296 6316 23348 6322
rect 23296 6258 23348 6264
rect 23204 6180 23256 6186
rect 23204 6122 23256 6128
rect 23400 3398 23428 8298
rect 23492 6866 23520 9046
rect 23480 6860 23532 6866
rect 23480 6802 23532 6808
rect 23584 6746 23612 9710
rect 23768 9110 23796 11194
rect 23756 9104 23808 9110
rect 23756 9046 23808 9052
rect 23664 8832 23716 8838
rect 23664 8774 23716 8780
rect 23676 7206 23704 8774
rect 24044 8634 24072 11194
rect 24032 8628 24084 8634
rect 24320 8616 24348 11194
rect 24400 8628 24452 8634
rect 24320 8588 24400 8616
rect 24032 8570 24084 8576
rect 24596 8616 24624 11194
rect 24676 8628 24728 8634
rect 24596 8588 24676 8616
rect 24400 8570 24452 8576
rect 24676 8570 24728 8576
rect 24872 8514 24900 11194
rect 25044 8900 25096 8906
rect 25044 8842 25096 8848
rect 25056 8634 25084 8842
rect 25148 8634 25176 11194
rect 25044 8628 25096 8634
rect 25044 8570 25096 8576
rect 25136 8628 25188 8634
rect 25136 8570 25188 8576
rect 25228 8560 25280 8566
rect 24216 8496 24268 8502
rect 24872 8486 25084 8514
rect 24216 8438 24268 8444
rect 23664 7200 23716 7206
rect 23664 7142 23716 7148
rect 23492 6718 23612 6746
rect 23664 6792 23716 6798
rect 23664 6734 23716 6740
rect 23938 6760 23994 6769
rect 23492 6458 23520 6718
rect 23572 6656 23624 6662
rect 23572 6598 23624 6604
rect 23480 6452 23532 6458
rect 23480 6394 23532 6400
rect 23584 6186 23612 6598
rect 23676 6458 23704 6734
rect 23938 6695 23994 6704
rect 23952 6662 23980 6695
rect 23848 6656 23900 6662
rect 23848 6598 23900 6604
rect 23940 6656 23992 6662
rect 23940 6598 23992 6604
rect 23664 6452 23716 6458
rect 23664 6394 23716 6400
rect 23572 6180 23624 6186
rect 23572 6122 23624 6128
rect 23860 6118 23888 6598
rect 23848 6112 23900 6118
rect 23848 6054 23900 6060
rect 23756 4616 23808 4622
rect 23756 4558 23808 4564
rect 23768 4049 23796 4558
rect 23754 4040 23810 4049
rect 23754 3975 23810 3984
rect 24228 3738 24256 8438
rect 25056 8362 25084 8486
rect 25148 8508 25228 8514
rect 25148 8502 25280 8508
rect 25148 8486 25268 8502
rect 25044 8356 25096 8362
rect 25044 8298 25096 8304
rect 25148 8242 25176 8486
rect 25424 8362 25452 11194
rect 25700 9654 25728 11194
rect 25688 9648 25740 9654
rect 25688 9590 25740 9596
rect 25504 8492 25556 8498
rect 25504 8434 25556 8440
rect 25412 8356 25464 8362
rect 25412 8298 25464 8304
rect 24780 8214 25176 8242
rect 24490 7984 24546 7993
rect 24490 7919 24546 7928
rect 24504 7546 24532 7919
rect 24492 7540 24544 7546
rect 24492 7482 24544 7488
rect 24400 6792 24452 6798
rect 24400 6734 24452 6740
rect 24412 6322 24440 6734
rect 24308 6316 24360 6322
rect 24308 6258 24360 6264
rect 24400 6316 24452 6322
rect 24400 6258 24452 6264
rect 24216 3732 24268 3738
rect 24216 3674 24268 3680
rect 23478 3632 23534 3641
rect 23478 3567 23534 3576
rect 23492 3534 23520 3567
rect 23480 3528 23532 3534
rect 23480 3470 23532 3476
rect 23388 3392 23440 3398
rect 23388 3334 23440 3340
rect 21824 2 21876 8
rect 23110 0 23166 56
rect 24320 42 24348 6258
rect 24780 4486 24808 8214
rect 24768 4480 24820 4486
rect 24768 4422 24820 4428
rect 25516 4078 25544 8434
rect 25976 8378 26004 11194
rect 26148 9648 26200 9654
rect 26148 9590 26200 9596
rect 25884 8350 26004 8378
rect 26160 8362 26188 9590
rect 26252 8634 26280 11194
rect 26528 8650 26556 11194
rect 26700 8900 26752 8906
rect 26700 8842 26752 8848
rect 26240 8628 26292 8634
rect 26528 8622 26648 8650
rect 26240 8570 26292 8576
rect 26422 8528 26478 8537
rect 26332 8492 26384 8498
rect 26422 8463 26478 8472
rect 26516 8492 26568 8498
rect 26332 8434 26384 8440
rect 26148 8356 26200 8362
rect 25884 8090 25912 8350
rect 26148 8298 26200 8304
rect 25950 8188 26258 8197
rect 25950 8186 25956 8188
rect 26012 8186 26036 8188
rect 26092 8186 26116 8188
rect 26172 8186 26196 8188
rect 26252 8186 26258 8188
rect 26012 8134 26014 8186
rect 26194 8134 26196 8186
rect 25950 8132 25956 8134
rect 26012 8132 26036 8134
rect 26092 8132 26116 8134
rect 26172 8132 26196 8134
rect 26252 8132 26258 8134
rect 25950 8123 26258 8132
rect 25872 8084 25924 8090
rect 25872 8026 25924 8032
rect 25872 7880 25924 7886
rect 25872 7822 25924 7828
rect 25778 7440 25834 7449
rect 25778 7375 25834 7384
rect 25792 6730 25820 7375
rect 25780 6724 25832 6730
rect 25780 6666 25832 6672
rect 25504 4072 25556 4078
rect 25504 4014 25556 4020
rect 25504 3936 25556 3942
rect 25504 3878 25556 3884
rect 25516 3738 25544 3878
rect 25884 3738 25912 7822
rect 26240 7744 26292 7750
rect 26240 7686 26292 7692
rect 26252 7274 26280 7686
rect 26240 7268 26292 7274
rect 26240 7210 26292 7216
rect 25950 7100 26258 7109
rect 25950 7098 25956 7100
rect 26012 7098 26036 7100
rect 26092 7098 26116 7100
rect 26172 7098 26196 7100
rect 26252 7098 26258 7100
rect 26012 7046 26014 7098
rect 26194 7046 26196 7098
rect 25950 7044 25956 7046
rect 26012 7044 26036 7046
rect 26092 7044 26116 7046
rect 26172 7044 26196 7046
rect 26252 7044 26258 7046
rect 25950 7035 26258 7044
rect 25950 6012 26258 6021
rect 25950 6010 25956 6012
rect 26012 6010 26036 6012
rect 26092 6010 26116 6012
rect 26172 6010 26196 6012
rect 26252 6010 26258 6012
rect 26012 5958 26014 6010
rect 26194 5958 26196 6010
rect 25950 5956 25956 5958
rect 26012 5956 26036 5958
rect 26092 5956 26116 5958
rect 26172 5956 26196 5958
rect 26252 5956 26258 5958
rect 25950 5947 26258 5956
rect 25950 4924 26258 4933
rect 25950 4922 25956 4924
rect 26012 4922 26036 4924
rect 26092 4922 26116 4924
rect 26172 4922 26196 4924
rect 26252 4922 26258 4924
rect 26012 4870 26014 4922
rect 26194 4870 26196 4922
rect 25950 4868 25956 4870
rect 26012 4868 26036 4870
rect 26092 4868 26116 4870
rect 26172 4868 26196 4870
rect 26252 4868 26258 4870
rect 25950 4859 26258 4868
rect 25950 3836 26258 3845
rect 25950 3834 25956 3836
rect 26012 3834 26036 3836
rect 26092 3834 26116 3836
rect 26172 3834 26196 3836
rect 26252 3834 26258 3836
rect 26012 3782 26014 3834
rect 26194 3782 26196 3834
rect 25950 3780 25956 3782
rect 26012 3780 26036 3782
rect 26092 3780 26116 3782
rect 26172 3780 26196 3782
rect 26252 3780 26258 3782
rect 25950 3771 26258 3780
rect 25504 3732 25556 3738
rect 25504 3674 25556 3680
rect 25872 3732 25924 3738
rect 25872 3674 25924 3680
rect 25596 3528 25648 3534
rect 25596 3470 25648 3476
rect 25688 3528 25740 3534
rect 25688 3470 25740 3476
rect 25608 105 25636 3470
rect 25700 2106 25728 3470
rect 26344 3398 26372 8434
rect 26436 7478 26464 8463
rect 26516 8434 26568 8440
rect 26424 7472 26476 7478
rect 26424 7414 26476 7420
rect 26424 6452 26476 6458
rect 26424 6394 26476 6400
rect 26332 3392 26384 3398
rect 26332 3334 26384 3340
rect 25950 2748 26258 2757
rect 25950 2746 25956 2748
rect 26012 2746 26036 2748
rect 26092 2746 26116 2748
rect 26172 2746 26196 2748
rect 26252 2746 26258 2748
rect 26012 2694 26014 2746
rect 26194 2694 26196 2746
rect 25950 2692 25956 2694
rect 26012 2692 26036 2694
rect 26092 2692 26116 2694
rect 26172 2692 26196 2694
rect 26252 2692 26258 2694
rect 25950 2683 26258 2692
rect 25688 2100 25740 2106
rect 25688 2042 25740 2048
rect 25594 96 25650 105
rect 24596 56 24716 82
rect 24596 54 24730 56
rect 24596 42 24624 54
rect 24320 14 24624 42
rect 24674 0 24730 54
rect 26252 56 26372 82
rect 25594 31 25650 40
rect 26238 54 26372 56
rect 26238 0 26294 54
rect 26344 42 26372 54
rect 26436 42 26464 6394
rect 26528 3942 26556 8434
rect 26620 8362 26648 8622
rect 26608 8356 26660 8362
rect 26608 8298 26660 8304
rect 26712 7002 26740 8842
rect 26804 8566 26832 11194
rect 27080 9466 27108 11194
rect 27356 9602 27384 11194
rect 27356 9574 27476 9602
rect 27080 9438 27384 9466
rect 26884 8968 26936 8974
rect 26884 8910 26936 8916
rect 26792 8560 26844 8566
rect 26792 8502 26844 8508
rect 26896 7478 26924 8910
rect 27010 8732 27318 8741
rect 27010 8730 27016 8732
rect 27072 8730 27096 8732
rect 27152 8730 27176 8732
rect 27232 8730 27256 8732
rect 27312 8730 27318 8732
rect 27072 8678 27074 8730
rect 27254 8678 27256 8730
rect 27010 8676 27016 8678
rect 27072 8676 27096 8678
rect 27152 8676 27176 8678
rect 27232 8676 27256 8678
rect 27312 8676 27318 8678
rect 27010 8667 27318 8676
rect 27356 8090 27384 9438
rect 27448 8634 27476 9574
rect 27632 9110 27660 11194
rect 27620 9104 27672 9110
rect 27620 9046 27672 9052
rect 27528 8968 27580 8974
rect 27528 8910 27580 8916
rect 27436 8628 27488 8634
rect 27436 8570 27488 8576
rect 27540 8344 27568 8910
rect 27908 8650 27936 11194
rect 28080 9036 28132 9042
rect 28080 8978 28132 8984
rect 27908 8622 28028 8650
rect 28000 8566 28028 8622
rect 27988 8560 28040 8566
rect 27988 8502 28040 8508
rect 28092 8498 28120 8978
rect 27712 8492 27764 8498
rect 27712 8434 27764 8440
rect 28080 8492 28132 8498
rect 28080 8434 28132 8440
rect 27448 8316 27568 8344
rect 27344 8084 27396 8090
rect 27344 8026 27396 8032
rect 27010 7644 27318 7653
rect 27010 7642 27016 7644
rect 27072 7642 27096 7644
rect 27152 7642 27176 7644
rect 27232 7642 27256 7644
rect 27312 7642 27318 7644
rect 27072 7590 27074 7642
rect 27254 7590 27256 7642
rect 27010 7588 27016 7590
rect 27072 7588 27096 7590
rect 27152 7588 27176 7590
rect 27232 7588 27256 7590
rect 27312 7588 27318 7590
rect 27010 7579 27318 7588
rect 26884 7472 26936 7478
rect 26884 7414 26936 7420
rect 27448 7206 27476 8316
rect 27620 8288 27672 8294
rect 27540 8236 27620 8242
rect 27540 8230 27672 8236
rect 27540 8214 27660 8230
rect 27436 7200 27488 7206
rect 27436 7142 27488 7148
rect 26700 6996 26752 7002
rect 26700 6938 26752 6944
rect 27010 6556 27318 6565
rect 27010 6554 27016 6556
rect 27072 6554 27096 6556
rect 27152 6554 27176 6556
rect 27232 6554 27256 6556
rect 27312 6554 27318 6556
rect 27072 6502 27074 6554
rect 27254 6502 27256 6554
rect 27010 6500 27016 6502
rect 27072 6500 27096 6502
rect 27152 6500 27176 6502
rect 27232 6500 27256 6502
rect 27312 6500 27318 6502
rect 27010 6491 27318 6500
rect 27540 5846 27568 8214
rect 27620 7948 27672 7954
rect 27620 7890 27672 7896
rect 27632 6662 27660 7890
rect 27620 6656 27672 6662
rect 27620 6598 27672 6604
rect 27528 5840 27580 5846
rect 27528 5782 27580 5788
rect 27010 5468 27318 5477
rect 27010 5466 27016 5468
rect 27072 5466 27096 5468
rect 27152 5466 27176 5468
rect 27232 5466 27256 5468
rect 27312 5466 27318 5468
rect 27072 5414 27074 5466
rect 27254 5414 27256 5466
rect 27010 5412 27016 5414
rect 27072 5412 27096 5414
rect 27152 5412 27176 5414
rect 27232 5412 27256 5414
rect 27312 5412 27318 5414
rect 27010 5403 27318 5412
rect 27724 4554 27752 8434
rect 28184 8090 28212 11194
rect 28172 8084 28224 8090
rect 28460 8072 28488 11194
rect 28632 9104 28684 9110
rect 28632 9046 28684 9052
rect 28644 8634 28672 9046
rect 28632 8628 28684 8634
rect 28632 8570 28684 8576
rect 28736 8362 28764 11194
rect 28816 8832 28868 8838
rect 28816 8774 28868 8780
rect 28828 8498 28856 8774
rect 28816 8492 28868 8498
rect 28816 8434 28868 8440
rect 28908 8492 28960 8498
rect 28908 8434 28960 8440
rect 28724 8356 28776 8362
rect 28724 8298 28776 8304
rect 28540 8084 28592 8090
rect 28460 8044 28540 8072
rect 28172 8026 28224 8032
rect 28540 8026 28592 8032
rect 28264 7880 28316 7886
rect 28264 7822 28316 7828
rect 28632 7880 28684 7886
rect 28632 7822 28684 7828
rect 27804 6316 27856 6322
rect 27804 6258 27856 6264
rect 27712 4548 27764 4554
rect 27712 4490 27764 4496
rect 27010 4380 27318 4389
rect 27010 4378 27016 4380
rect 27072 4378 27096 4380
rect 27152 4378 27176 4380
rect 27232 4378 27256 4380
rect 27312 4378 27318 4380
rect 27072 4326 27074 4378
rect 27254 4326 27256 4378
rect 27010 4324 27016 4326
rect 27072 4324 27096 4326
rect 27152 4324 27176 4326
rect 27232 4324 27256 4326
rect 27312 4324 27318 4326
rect 27010 4315 27318 4324
rect 26884 4140 26936 4146
rect 26884 4082 26936 4088
rect 26516 3936 26568 3942
rect 26516 3878 26568 3884
rect 26896 3058 26924 4082
rect 27010 3292 27318 3301
rect 27010 3290 27016 3292
rect 27072 3290 27096 3292
rect 27152 3290 27176 3292
rect 27232 3290 27256 3292
rect 27312 3290 27318 3292
rect 27072 3238 27074 3290
rect 27254 3238 27256 3290
rect 27010 3236 27016 3238
rect 27072 3236 27096 3238
rect 27152 3236 27176 3238
rect 27232 3236 27256 3238
rect 27312 3236 27318 3238
rect 27010 3227 27318 3236
rect 26884 3052 26936 3058
rect 26884 2994 26936 3000
rect 27010 2204 27318 2213
rect 27010 2202 27016 2204
rect 27072 2202 27096 2204
rect 27152 2202 27176 2204
rect 27232 2202 27256 2204
rect 27312 2202 27318 2204
rect 27072 2150 27074 2202
rect 27254 2150 27256 2202
rect 27010 2148 27016 2150
rect 27072 2148 27096 2150
rect 27152 2148 27176 2150
rect 27232 2148 27256 2150
rect 27312 2148 27318 2150
rect 27010 2139 27318 2148
rect 27816 56 27844 6258
rect 28276 6186 28304 7822
rect 28264 6180 28316 6186
rect 28264 6122 28316 6128
rect 28644 6118 28672 7822
rect 28920 7274 28948 8434
rect 29012 8430 29040 11194
rect 29000 8424 29052 8430
rect 29000 8366 29052 8372
rect 29288 8090 29316 11194
rect 29564 8634 29592 11194
rect 32310 9888 32366 9897
rect 32310 9823 32366 9832
rect 30654 9616 30710 9625
rect 30654 9551 30710 9560
rect 29920 8900 29972 8906
rect 29920 8842 29972 8848
rect 29552 8628 29604 8634
rect 29552 8570 29604 8576
rect 29932 8498 29960 8842
rect 29552 8492 29604 8498
rect 29552 8434 29604 8440
rect 29920 8492 29972 8498
rect 29920 8434 29972 8440
rect 30564 8492 30616 8498
rect 30564 8434 30616 8440
rect 29276 8084 29328 8090
rect 29276 8026 29328 8032
rect 29092 7880 29144 7886
rect 29092 7822 29144 7828
rect 29000 7812 29052 7818
rect 29000 7754 29052 7760
rect 29012 7546 29040 7754
rect 29000 7540 29052 7546
rect 29000 7482 29052 7488
rect 28908 7268 28960 7274
rect 28908 7210 28960 7216
rect 28724 6656 28776 6662
rect 28724 6598 28776 6604
rect 28632 6112 28684 6118
rect 28632 6054 28684 6060
rect 28736 4690 28764 6598
rect 29104 6458 29132 7822
rect 29564 6866 29592 8434
rect 30472 7880 30524 7886
rect 30472 7822 30524 7828
rect 30380 7268 30432 7274
rect 30380 7210 30432 7216
rect 30288 7200 30340 7206
rect 30288 7142 30340 7148
rect 30300 6866 30328 7142
rect 29552 6860 29604 6866
rect 29552 6802 29604 6808
rect 30288 6860 30340 6866
rect 30288 6802 30340 6808
rect 29368 6792 29420 6798
rect 29368 6734 29420 6740
rect 29092 6452 29144 6458
rect 29092 6394 29144 6400
rect 28724 4684 28776 4690
rect 28724 4626 28776 4632
rect 29000 4616 29052 4622
rect 29000 4558 29052 4564
rect 29012 3602 29040 4558
rect 29000 3596 29052 3602
rect 29000 3538 29052 3544
rect 29380 56 29408 6734
rect 30392 5098 30420 7210
rect 30484 6254 30512 7822
rect 30576 6458 30604 8434
rect 30668 8090 30696 9551
rect 31482 9344 31538 9353
rect 31482 9279 31538 9288
rect 31022 9072 31078 9081
rect 31022 9007 31078 9016
rect 31036 8090 31064 9007
rect 31390 8800 31446 8809
rect 31390 8735 31446 8744
rect 31116 8628 31168 8634
rect 31116 8570 31168 8576
rect 31128 8537 31156 8570
rect 31114 8528 31170 8537
rect 31114 8463 31170 8472
rect 31300 8492 31352 8498
rect 31300 8434 31352 8440
rect 30656 8084 30708 8090
rect 30656 8026 30708 8032
rect 31024 8084 31076 8090
rect 31024 8026 31076 8032
rect 30656 7880 30708 7886
rect 30656 7822 30708 7828
rect 30932 7880 30984 7886
rect 30932 7822 30984 7828
rect 30564 6452 30616 6458
rect 30564 6394 30616 6400
rect 30668 6390 30696 7822
rect 30944 6730 30972 7822
rect 31312 7750 31340 8434
rect 31404 8090 31432 8735
rect 31392 8084 31444 8090
rect 31392 8026 31444 8032
rect 31300 7744 31352 7750
rect 31300 7686 31352 7692
rect 31496 7546 31524 9279
rect 31668 8968 31720 8974
rect 31668 8910 31720 8916
rect 31680 8498 31708 8910
rect 31668 8492 31720 8498
rect 31668 8434 31720 8440
rect 31852 8288 31904 8294
rect 31852 8230 31904 8236
rect 31864 7993 31892 8230
rect 31950 8188 32258 8197
rect 31950 8186 31956 8188
rect 32012 8186 32036 8188
rect 32092 8186 32116 8188
rect 32172 8186 32196 8188
rect 32252 8186 32258 8188
rect 32012 8134 32014 8186
rect 32194 8134 32196 8186
rect 31950 8132 31956 8134
rect 32012 8132 32036 8134
rect 32092 8132 32116 8134
rect 32172 8132 32196 8134
rect 32252 8132 32258 8134
rect 31950 8123 32258 8132
rect 31850 7984 31906 7993
rect 31850 7919 31906 7928
rect 31760 7744 31812 7750
rect 32128 7744 32180 7750
rect 31760 7686 31812 7692
rect 32126 7712 32128 7721
rect 32180 7712 32182 7721
rect 31484 7540 31536 7546
rect 31484 7482 31536 7488
rect 31772 7449 31800 7686
rect 32126 7647 32182 7656
rect 31758 7440 31814 7449
rect 31758 7375 31814 7384
rect 31950 7100 32258 7109
rect 31950 7098 31956 7100
rect 32012 7098 32036 7100
rect 32092 7098 32116 7100
rect 32172 7098 32196 7100
rect 32252 7098 32258 7100
rect 32012 7046 32014 7098
rect 32194 7046 32196 7098
rect 31950 7044 31956 7046
rect 32012 7044 32036 7046
rect 32092 7044 32116 7046
rect 32172 7044 32196 7046
rect 32252 7044 32258 7046
rect 31950 7035 32258 7044
rect 31758 6896 31814 6905
rect 31758 6831 31814 6840
rect 31668 6792 31720 6798
rect 31668 6734 31720 6740
rect 30932 6724 30984 6730
rect 30932 6666 30984 6672
rect 31392 6656 31444 6662
rect 31390 6624 31392 6633
rect 31444 6624 31446 6633
rect 31390 6559 31446 6568
rect 30656 6384 30708 6390
rect 30656 6326 30708 6332
rect 30932 6316 30984 6322
rect 30932 6258 30984 6264
rect 31300 6316 31352 6322
rect 31300 6258 31352 6264
rect 31392 6316 31444 6322
rect 31392 6258 31444 6264
rect 30472 6248 30524 6254
rect 30472 6190 30524 6196
rect 30380 5092 30432 5098
rect 30380 5034 30432 5040
rect 30380 3052 30432 3058
rect 30380 2994 30432 3000
rect 30392 2310 30420 2994
rect 30484 2514 30880 2530
rect 30472 2508 30880 2514
rect 30524 2502 30880 2508
rect 30472 2450 30524 2456
rect 30852 2446 30880 2502
rect 30840 2440 30892 2446
rect 30840 2382 30892 2388
rect 30380 2304 30432 2310
rect 30380 2246 30432 2252
rect 30748 2304 30800 2310
rect 30748 2246 30800 2252
rect 30760 2009 30788 2246
rect 30746 2000 30802 2009
rect 30746 1935 30802 1944
rect 30944 56 30972 6258
rect 31312 5914 31340 6258
rect 31300 5908 31352 5914
rect 31300 5850 31352 5856
rect 31208 5704 31260 5710
rect 31208 5646 31260 5652
rect 31300 5704 31352 5710
rect 31300 5646 31352 5652
rect 31220 4010 31248 5646
rect 31208 4004 31260 4010
rect 31208 3946 31260 3952
rect 31312 3466 31340 5646
rect 31404 4826 31432 6258
rect 31482 6216 31538 6225
rect 31482 6151 31484 6160
rect 31536 6151 31538 6160
rect 31484 6122 31536 6128
rect 31680 5642 31708 6734
rect 31772 6662 31800 6831
rect 32324 6662 32352 9823
rect 32588 8356 32640 8362
rect 32588 8298 32640 8304
rect 32600 8265 32628 8298
rect 32586 8256 32642 8265
rect 32586 8191 32642 8200
rect 32772 7200 32824 7206
rect 32770 7168 32772 7177
rect 32824 7168 32826 7177
rect 32770 7103 32826 7112
rect 31760 6656 31812 6662
rect 31760 6598 31812 6604
rect 32312 6656 32364 6662
rect 32312 6598 32364 6604
rect 31852 6452 31904 6458
rect 31852 6394 31904 6400
rect 31864 6361 31892 6394
rect 31850 6352 31906 6361
rect 31850 6287 31906 6296
rect 32496 6248 32548 6254
rect 32496 6190 32548 6196
rect 31950 6012 32258 6021
rect 31950 6010 31956 6012
rect 32012 6010 32036 6012
rect 32092 6010 32116 6012
rect 32172 6010 32196 6012
rect 32252 6010 32258 6012
rect 32012 5958 32014 6010
rect 32194 5958 32196 6010
rect 31950 5956 31956 5958
rect 32012 5956 32036 5958
rect 32092 5956 32116 5958
rect 32172 5956 32196 5958
rect 32252 5956 32258 5958
rect 31950 5947 32258 5956
rect 32036 5840 32088 5846
rect 32128 5840 32180 5846
rect 32036 5782 32088 5788
rect 32126 5808 32128 5817
rect 32180 5808 32182 5817
rect 31852 5704 31904 5710
rect 31852 5646 31904 5652
rect 31668 5636 31720 5642
rect 31668 5578 31720 5584
rect 31760 5568 31812 5574
rect 31758 5536 31760 5545
rect 31812 5536 31814 5545
rect 31758 5471 31814 5480
rect 31668 5228 31720 5234
rect 31668 5170 31720 5176
rect 31484 5024 31536 5030
rect 31484 4966 31536 4972
rect 31392 4820 31444 4826
rect 31392 4762 31444 4768
rect 31496 4729 31524 4966
rect 31680 4758 31708 5170
rect 31668 4752 31720 4758
rect 31482 4720 31538 4729
rect 31668 4694 31720 4700
rect 31482 4655 31538 4664
rect 31760 4480 31812 4486
rect 31760 4422 31812 4428
rect 31772 4185 31800 4422
rect 31758 4176 31814 4185
rect 31392 4140 31444 4146
rect 31758 4111 31814 4120
rect 31392 4082 31444 4088
rect 31300 3460 31352 3466
rect 31300 3402 31352 3408
rect 31404 2922 31432 4082
rect 31484 3936 31536 3942
rect 31484 3878 31536 3884
rect 31496 3641 31524 3878
rect 31864 3670 31892 5646
rect 32048 5273 32076 5782
rect 32126 5743 32182 5752
rect 32034 5264 32090 5273
rect 32034 5199 32090 5208
rect 31950 4924 32258 4933
rect 31950 4922 31956 4924
rect 32012 4922 32036 4924
rect 32092 4922 32116 4924
rect 32172 4922 32196 4924
rect 32252 4922 32258 4924
rect 32012 4870 32014 4922
rect 32194 4870 32196 4922
rect 31950 4868 31956 4870
rect 32012 4868 32036 4870
rect 32092 4868 32116 4870
rect 32172 4868 32196 4870
rect 32252 4868 32258 4870
rect 31950 4859 32258 4868
rect 31944 4616 31996 4622
rect 31944 4558 31996 4564
rect 31956 4282 31984 4558
rect 32128 4480 32180 4486
rect 32126 4448 32128 4457
rect 32180 4448 32182 4457
rect 32126 4383 32182 4392
rect 31944 4276 31996 4282
rect 31944 4218 31996 4224
rect 31950 3836 32258 3845
rect 31950 3834 31956 3836
rect 32012 3834 32036 3836
rect 32092 3834 32116 3836
rect 32172 3834 32196 3836
rect 32252 3834 32258 3836
rect 32012 3782 32014 3834
rect 32194 3782 32196 3834
rect 31950 3780 31956 3782
rect 32012 3780 32036 3782
rect 32092 3780 32116 3782
rect 32172 3780 32196 3782
rect 32252 3780 32258 3782
rect 31950 3771 32258 3780
rect 31852 3664 31904 3670
rect 31482 3632 31538 3641
rect 31852 3606 31904 3612
rect 31482 3567 31538 3576
rect 31576 3528 31628 3534
rect 31944 3528 31996 3534
rect 31576 3470 31628 3476
rect 31666 3496 31722 3505
rect 31588 3126 31616 3470
rect 31944 3470 31996 3476
rect 31666 3431 31722 3440
rect 31576 3120 31628 3126
rect 31576 3062 31628 3068
rect 31680 3058 31708 3431
rect 31760 3392 31812 3398
rect 31760 3334 31812 3340
rect 31772 3097 31800 3334
rect 31956 3194 31984 3470
rect 32128 3392 32180 3398
rect 32126 3360 32128 3369
rect 32180 3360 32182 3369
rect 32126 3295 32182 3304
rect 31944 3188 31996 3194
rect 31944 3130 31996 3136
rect 31758 3088 31814 3097
rect 31668 3052 31720 3058
rect 31758 3023 31814 3032
rect 31668 2994 31720 3000
rect 31392 2916 31444 2922
rect 31392 2858 31444 2864
rect 31760 2848 31812 2854
rect 31760 2790 31812 2796
rect 31772 2553 31800 2790
rect 31950 2748 32258 2757
rect 31950 2746 31956 2748
rect 32012 2746 32036 2748
rect 32092 2746 32116 2748
rect 32172 2746 32196 2748
rect 32252 2746 32258 2748
rect 32012 2694 32014 2746
rect 32194 2694 32196 2746
rect 31950 2692 31956 2694
rect 32012 2692 32036 2694
rect 32092 2692 32116 2694
rect 32172 2692 32196 2694
rect 32252 2692 32258 2694
rect 31950 2683 32258 2692
rect 31758 2544 31814 2553
rect 31758 2479 31814 2488
rect 31116 2304 31168 2310
rect 31116 2246 31168 2252
rect 31484 2304 31536 2310
rect 31852 2304 31904 2310
rect 31484 2246 31536 2252
rect 31850 2272 31852 2281
rect 31904 2272 31906 2281
rect 31128 1737 31156 2246
rect 31114 1728 31170 1737
rect 31114 1663 31170 1672
rect 31496 1465 31524 2246
rect 31850 2207 31906 2216
rect 31482 1456 31538 1465
rect 31482 1391 31538 1400
rect 32508 56 32536 6190
rect 32864 5024 32916 5030
rect 32862 4992 32864 5001
rect 32916 4992 32918 5001
rect 32862 4927 32918 4936
rect 32864 3936 32916 3942
rect 32862 3904 32864 3913
rect 32916 3904 32918 3913
rect 32862 3839 32918 3848
rect 32864 2848 32916 2854
rect 32862 2816 32864 2825
rect 32916 2816 32918 2825
rect 32862 2751 32918 2760
rect 26344 14 26464 42
rect 27802 0 27858 56
rect 29366 0 29422 56
rect 30930 0 30986 56
rect 32494 0 32550 56
<< via2 >>
rect 3016 8730 3072 8732
rect 3096 8730 3152 8732
rect 3176 8730 3232 8732
rect 3256 8730 3312 8732
rect 3016 8678 3062 8730
rect 3062 8678 3072 8730
rect 3096 8678 3126 8730
rect 3126 8678 3138 8730
rect 3138 8678 3152 8730
rect 3176 8678 3190 8730
rect 3190 8678 3202 8730
rect 3202 8678 3232 8730
rect 3256 8678 3266 8730
rect 3266 8678 3312 8730
rect 3016 8676 3072 8678
rect 3096 8676 3152 8678
rect 3176 8676 3232 8678
rect 3256 8676 3312 8678
rect 1956 8186 2012 8188
rect 2036 8186 2092 8188
rect 2116 8186 2172 8188
rect 2196 8186 2252 8188
rect 1956 8134 2002 8186
rect 2002 8134 2012 8186
rect 2036 8134 2066 8186
rect 2066 8134 2078 8186
rect 2078 8134 2092 8186
rect 2116 8134 2130 8186
rect 2130 8134 2142 8186
rect 2142 8134 2172 8186
rect 2196 8134 2206 8186
rect 2206 8134 2252 8186
rect 1956 8132 2012 8134
rect 2036 8132 2092 8134
rect 2116 8132 2172 8134
rect 2196 8132 2252 8134
rect 3016 7642 3072 7644
rect 3096 7642 3152 7644
rect 3176 7642 3232 7644
rect 3256 7642 3312 7644
rect 3016 7590 3062 7642
rect 3062 7590 3072 7642
rect 3096 7590 3126 7642
rect 3126 7590 3138 7642
rect 3138 7590 3152 7642
rect 3176 7590 3190 7642
rect 3190 7590 3202 7642
rect 3202 7590 3232 7642
rect 3256 7590 3266 7642
rect 3266 7590 3312 7642
rect 3016 7588 3072 7590
rect 3096 7588 3152 7590
rect 3176 7588 3232 7590
rect 3256 7588 3312 7590
rect 1956 7098 2012 7100
rect 2036 7098 2092 7100
rect 2116 7098 2172 7100
rect 2196 7098 2252 7100
rect 1956 7046 2002 7098
rect 2002 7046 2012 7098
rect 2036 7046 2066 7098
rect 2066 7046 2078 7098
rect 2078 7046 2092 7098
rect 2116 7046 2130 7098
rect 2130 7046 2142 7098
rect 2142 7046 2172 7098
rect 2196 7046 2206 7098
rect 2206 7046 2252 7098
rect 1956 7044 2012 7046
rect 2036 7044 2092 7046
rect 2116 7044 2172 7046
rect 2196 7044 2252 7046
rect 570 6568 626 6624
rect 3016 6554 3072 6556
rect 3096 6554 3152 6556
rect 3176 6554 3232 6556
rect 3256 6554 3312 6556
rect 3016 6502 3062 6554
rect 3062 6502 3072 6554
rect 3096 6502 3126 6554
rect 3126 6502 3138 6554
rect 3138 6502 3152 6554
rect 3176 6502 3190 6554
rect 3190 6502 3202 6554
rect 3202 6502 3232 6554
rect 3256 6502 3266 6554
rect 3266 6502 3312 6554
rect 3016 6500 3072 6502
rect 3096 6500 3152 6502
rect 3176 6500 3232 6502
rect 3256 6500 3312 6502
rect 4618 6160 4674 6216
rect 6458 10784 6514 10840
rect 1956 6010 2012 6012
rect 2036 6010 2092 6012
rect 2116 6010 2172 6012
rect 2196 6010 2252 6012
rect 1956 5958 2002 6010
rect 2002 5958 2012 6010
rect 2036 5958 2066 6010
rect 2066 5958 2078 6010
rect 2078 5958 2092 6010
rect 2116 5958 2130 6010
rect 2130 5958 2142 6010
rect 2142 5958 2172 6010
rect 2196 5958 2206 6010
rect 2206 5958 2252 6010
rect 1956 5956 2012 5958
rect 2036 5956 2092 5958
rect 2116 5956 2172 5958
rect 2196 5956 2252 5958
rect 3016 5466 3072 5468
rect 3096 5466 3152 5468
rect 3176 5466 3232 5468
rect 3256 5466 3312 5468
rect 3016 5414 3062 5466
rect 3062 5414 3072 5466
rect 3096 5414 3126 5466
rect 3126 5414 3138 5466
rect 3138 5414 3152 5466
rect 3176 5414 3190 5466
rect 3190 5414 3202 5466
rect 3202 5414 3232 5466
rect 3256 5414 3266 5466
rect 3266 5414 3312 5466
rect 3016 5412 3072 5414
rect 3096 5412 3152 5414
rect 3176 5412 3232 5414
rect 3256 5412 3312 5414
rect 1306 5208 1362 5264
rect 7010 10376 7066 10432
rect 7562 9696 7618 9752
rect 7838 9968 7894 10024
rect 7956 8186 8012 8188
rect 8036 8186 8092 8188
rect 8116 8186 8172 8188
rect 8196 8186 8252 8188
rect 7956 8134 8002 8186
rect 8002 8134 8012 8186
rect 8036 8134 8066 8186
rect 8066 8134 8078 8186
rect 8078 8134 8092 8186
rect 8116 8134 8130 8186
rect 8130 8134 8142 8186
rect 8142 8134 8172 8186
rect 8196 8134 8206 8186
rect 8206 8134 8252 8186
rect 7956 8132 8012 8134
rect 8036 8132 8092 8134
rect 8116 8132 8172 8134
rect 8196 8132 8252 8134
rect 7956 7098 8012 7100
rect 8036 7098 8092 7100
rect 8116 7098 8172 7100
rect 8196 7098 8252 7100
rect 7956 7046 8002 7098
rect 8002 7046 8012 7098
rect 8036 7046 8066 7098
rect 8066 7046 8078 7098
rect 8078 7046 8092 7098
rect 8116 7046 8130 7098
rect 8130 7046 8142 7098
rect 8142 7046 8172 7098
rect 8196 7046 8206 7098
rect 8206 7046 8252 7098
rect 7956 7044 8012 7046
rect 8036 7044 8092 7046
rect 8116 7044 8172 7046
rect 8196 7044 8252 7046
rect 9016 8730 9072 8732
rect 9096 8730 9152 8732
rect 9176 8730 9232 8732
rect 9256 8730 9312 8732
rect 9016 8678 9062 8730
rect 9062 8678 9072 8730
rect 9096 8678 9126 8730
rect 9126 8678 9138 8730
rect 9138 8678 9152 8730
rect 9176 8678 9190 8730
rect 9190 8678 9202 8730
rect 9202 8678 9232 8730
rect 9256 8678 9266 8730
rect 9266 8678 9312 8730
rect 9016 8676 9072 8678
rect 9096 8676 9152 8678
rect 9176 8676 9232 8678
rect 9256 8676 9312 8678
rect 10046 9560 10102 9616
rect 9016 7642 9072 7644
rect 9096 7642 9152 7644
rect 9176 7642 9232 7644
rect 9256 7642 9312 7644
rect 9016 7590 9062 7642
rect 9062 7590 9072 7642
rect 9096 7590 9126 7642
rect 9126 7590 9138 7642
rect 9138 7590 9152 7642
rect 9176 7590 9190 7642
rect 9190 7590 9202 7642
rect 9202 7590 9232 7642
rect 9256 7590 9266 7642
rect 9266 7590 9312 7642
rect 9016 7588 9072 7590
rect 9096 7588 9152 7590
rect 9176 7588 9232 7590
rect 9256 7588 9312 7590
rect 8850 7112 8906 7168
rect 9016 6554 9072 6556
rect 9096 6554 9152 6556
rect 9176 6554 9232 6556
rect 9256 6554 9312 6556
rect 9016 6502 9062 6554
rect 9062 6502 9072 6554
rect 9096 6502 9126 6554
rect 9126 6502 9138 6554
rect 9138 6502 9152 6554
rect 9176 6502 9190 6554
rect 9190 6502 9202 6554
rect 9202 6502 9232 6554
rect 9256 6502 9266 6554
rect 9266 6502 9312 6554
rect 9016 6500 9072 6502
rect 9096 6500 9152 6502
rect 9176 6500 9232 6502
rect 9256 6500 9312 6502
rect 9586 7656 9642 7712
rect 9586 7248 9642 7304
rect 9678 7112 9734 7168
rect 9862 6976 9918 7032
rect 7956 6010 8012 6012
rect 8036 6010 8092 6012
rect 8116 6010 8172 6012
rect 8196 6010 8252 6012
rect 7956 5958 8002 6010
rect 8002 5958 8012 6010
rect 8036 5958 8066 6010
rect 8066 5958 8078 6010
rect 8078 5958 8092 6010
rect 8116 5958 8130 6010
rect 8130 5958 8142 6010
rect 8142 5958 8172 6010
rect 8196 5958 8206 6010
rect 8206 5958 8252 6010
rect 7956 5956 8012 5958
rect 8036 5956 8092 5958
rect 8116 5956 8172 5958
rect 8196 5956 8252 5958
rect 9126 6160 9182 6216
rect 9770 6432 9826 6488
rect 9016 5466 9072 5468
rect 9096 5466 9152 5468
rect 9176 5466 9232 5468
rect 9256 5466 9312 5468
rect 9016 5414 9062 5466
rect 9062 5414 9072 5466
rect 9096 5414 9126 5466
rect 9126 5414 9138 5466
rect 9138 5414 9152 5466
rect 9176 5414 9190 5466
rect 9190 5414 9202 5466
rect 9202 5414 9232 5466
rect 9256 5414 9266 5466
rect 9266 5414 9312 5466
rect 9016 5412 9072 5414
rect 9096 5412 9152 5414
rect 9176 5412 9232 5414
rect 9256 5412 9312 5414
rect 6918 5208 6974 5264
rect 10690 6740 10692 6760
rect 10692 6740 10744 6760
rect 10744 6740 10746 6760
rect 10690 6704 10746 6740
rect 10598 6432 10654 6488
rect 11794 9152 11850 9208
rect 12070 8744 12126 8800
rect 12438 6296 12494 6352
rect 2870 5072 2926 5128
rect 1766 4936 1822 4992
rect 1956 4922 2012 4924
rect 2036 4922 2092 4924
rect 2116 4922 2172 4924
rect 2196 4922 2252 4924
rect 1956 4870 2002 4922
rect 2002 4870 2012 4922
rect 2036 4870 2066 4922
rect 2066 4870 2078 4922
rect 2078 4870 2092 4922
rect 2116 4870 2130 4922
rect 2130 4870 2142 4922
rect 2142 4870 2172 4922
rect 2196 4870 2206 4922
rect 2206 4870 2252 4922
rect 1956 4868 2012 4870
rect 2036 4868 2092 4870
rect 2116 4868 2172 4870
rect 2196 4868 2252 4870
rect 1766 4528 1822 4584
rect 2870 4392 2926 4448
rect 3016 4378 3072 4380
rect 3096 4378 3152 4380
rect 3176 4378 3232 4380
rect 3256 4378 3312 4380
rect 3016 4326 3062 4378
rect 3062 4326 3072 4378
rect 3096 4326 3126 4378
rect 3126 4326 3138 4378
rect 3138 4326 3152 4378
rect 3176 4326 3190 4378
rect 3190 4326 3202 4378
rect 3202 4326 3232 4378
rect 3256 4326 3266 4378
rect 3266 4326 3312 4378
rect 3016 4324 3072 4326
rect 3096 4324 3152 4326
rect 3176 4324 3232 4326
rect 3256 4324 3312 4326
rect 7956 4922 8012 4924
rect 8036 4922 8092 4924
rect 8116 4922 8172 4924
rect 8196 4922 8252 4924
rect 7956 4870 8002 4922
rect 8002 4870 8012 4922
rect 8036 4870 8066 4922
rect 8066 4870 8078 4922
rect 8078 4870 8092 4922
rect 8116 4870 8130 4922
rect 8130 4870 8142 4922
rect 8142 4870 8172 4922
rect 8196 4870 8206 4922
rect 8206 4870 8252 4922
rect 7956 4868 8012 4870
rect 8036 4868 8092 4870
rect 8116 4868 8172 4870
rect 8196 4868 8252 4870
rect 9016 4378 9072 4380
rect 9096 4378 9152 4380
rect 9176 4378 9232 4380
rect 9256 4378 9312 4380
rect 9016 4326 9062 4378
rect 9062 4326 9072 4378
rect 9096 4326 9126 4378
rect 9126 4326 9138 4378
rect 9138 4326 9152 4378
rect 9176 4326 9190 4378
rect 9190 4326 9202 4378
rect 9202 4326 9232 4378
rect 9256 4326 9266 4378
rect 9266 4326 9312 4378
rect 9016 4324 9072 4326
rect 9096 4324 9152 4326
rect 9176 4324 9232 4326
rect 9256 4324 9312 4326
rect 13726 9832 13782 9888
rect 14922 10784 14978 10840
rect 14646 9968 14702 10024
rect 14370 9696 14426 9752
rect 14462 9424 14518 9480
rect 14462 9016 14518 9072
rect 15474 9152 15530 9208
rect 15016 8730 15072 8732
rect 15096 8730 15152 8732
rect 15176 8730 15232 8732
rect 15256 8730 15312 8732
rect 15016 8678 15062 8730
rect 15062 8678 15072 8730
rect 15096 8678 15126 8730
rect 15126 8678 15138 8730
rect 15138 8678 15152 8730
rect 15176 8678 15190 8730
rect 15190 8678 15202 8730
rect 15202 8678 15232 8730
rect 15256 8678 15266 8730
rect 15266 8678 15312 8730
rect 15016 8676 15072 8678
rect 15096 8676 15152 8678
rect 15176 8676 15232 8678
rect 15256 8676 15312 8678
rect 13956 8186 14012 8188
rect 14036 8186 14092 8188
rect 14116 8186 14172 8188
rect 14196 8186 14252 8188
rect 13956 8134 14002 8186
rect 14002 8134 14012 8186
rect 14036 8134 14066 8186
rect 14066 8134 14078 8186
rect 14078 8134 14092 8186
rect 14116 8134 14130 8186
rect 14130 8134 14142 8186
rect 14142 8134 14172 8186
rect 14196 8134 14206 8186
rect 14206 8134 14252 8186
rect 13956 8132 14012 8134
rect 14036 8132 14092 8134
rect 14116 8132 14172 8134
rect 14196 8132 14252 8134
rect 14830 8064 14886 8120
rect 13956 7098 14012 7100
rect 14036 7098 14092 7100
rect 14116 7098 14172 7100
rect 14196 7098 14252 7100
rect 13956 7046 14002 7098
rect 14002 7046 14012 7098
rect 14036 7046 14066 7098
rect 14066 7046 14078 7098
rect 14078 7046 14092 7098
rect 14116 7046 14130 7098
rect 14130 7046 14142 7098
rect 14142 7046 14172 7098
rect 14196 7046 14206 7098
rect 14206 7046 14252 7098
rect 13956 7044 14012 7046
rect 14036 7044 14092 7046
rect 14116 7044 14172 7046
rect 14196 7044 14252 7046
rect 14830 7656 14886 7712
rect 15016 7642 15072 7644
rect 15096 7642 15152 7644
rect 15176 7642 15232 7644
rect 15256 7642 15312 7644
rect 15016 7590 15062 7642
rect 15062 7590 15072 7642
rect 15096 7590 15126 7642
rect 15126 7590 15138 7642
rect 15138 7590 15152 7642
rect 15176 7590 15190 7642
rect 15190 7590 15202 7642
rect 15202 7590 15232 7642
rect 15256 7590 15266 7642
rect 15266 7590 15312 7642
rect 15016 7588 15072 7590
rect 15096 7588 15152 7590
rect 15176 7588 15232 7590
rect 15256 7588 15312 7590
rect 15016 6554 15072 6556
rect 15096 6554 15152 6556
rect 15176 6554 15232 6556
rect 15256 6554 15312 6556
rect 15016 6502 15062 6554
rect 15062 6502 15072 6554
rect 15096 6502 15126 6554
rect 15126 6502 15138 6554
rect 15138 6502 15152 6554
rect 15176 6502 15190 6554
rect 15190 6502 15202 6554
rect 15202 6502 15232 6554
rect 15256 6502 15266 6554
rect 15266 6502 15312 6554
rect 15016 6500 15072 6502
rect 15096 6500 15152 6502
rect 15176 6500 15232 6502
rect 15256 6500 15312 6502
rect 13956 6010 14012 6012
rect 14036 6010 14092 6012
rect 14116 6010 14172 6012
rect 14196 6010 14252 6012
rect 13956 5958 14002 6010
rect 14002 5958 14012 6010
rect 14036 5958 14066 6010
rect 14066 5958 14078 6010
rect 14078 5958 14092 6010
rect 14116 5958 14130 6010
rect 14130 5958 14142 6010
rect 14142 5958 14172 6010
rect 14196 5958 14206 6010
rect 14206 5958 14252 6010
rect 13956 5956 14012 5958
rect 14036 5956 14092 5958
rect 14116 5956 14172 5958
rect 14196 5956 14252 5958
rect 13726 5752 13782 5808
rect 9402 3984 9458 4040
rect 13634 3984 13690 4040
rect 1956 3834 2012 3836
rect 2036 3834 2092 3836
rect 2116 3834 2172 3836
rect 2196 3834 2252 3836
rect 1956 3782 2002 3834
rect 2002 3782 2012 3834
rect 2036 3782 2066 3834
rect 2066 3782 2078 3834
rect 2078 3782 2092 3834
rect 2116 3782 2130 3834
rect 2130 3782 2142 3834
rect 2142 3782 2172 3834
rect 2196 3782 2206 3834
rect 2206 3782 2252 3834
rect 1956 3780 2012 3782
rect 2036 3780 2092 3782
rect 2116 3780 2172 3782
rect 2196 3780 2252 3782
rect 7956 3834 8012 3836
rect 8036 3834 8092 3836
rect 8116 3834 8172 3836
rect 8196 3834 8252 3836
rect 7956 3782 8002 3834
rect 8002 3782 8012 3834
rect 8036 3782 8066 3834
rect 8066 3782 8078 3834
rect 8078 3782 8092 3834
rect 8116 3782 8130 3834
rect 8130 3782 8142 3834
rect 8142 3782 8172 3834
rect 8196 3782 8206 3834
rect 8206 3782 8252 3834
rect 7956 3780 8012 3782
rect 8036 3780 8092 3782
rect 8116 3780 8172 3782
rect 8196 3780 8252 3782
rect 1766 3440 1822 3496
rect 1950 3304 2006 3360
rect 3016 3290 3072 3292
rect 3096 3290 3152 3292
rect 3176 3290 3232 3292
rect 3256 3290 3312 3292
rect 3016 3238 3062 3290
rect 3062 3238 3072 3290
rect 3096 3238 3126 3290
rect 3126 3238 3138 3290
rect 3138 3238 3152 3290
rect 3176 3238 3190 3290
rect 3190 3238 3202 3290
rect 3202 3238 3232 3290
rect 3256 3238 3266 3290
rect 3266 3238 3312 3290
rect 3016 3236 3072 3238
rect 3096 3236 3152 3238
rect 3176 3236 3232 3238
rect 3256 3236 3312 3238
rect 1950 2896 2006 2952
rect 1766 2760 1822 2816
rect 1956 2746 2012 2748
rect 2036 2746 2092 2748
rect 2116 2746 2172 2748
rect 2196 2746 2252 2748
rect 1956 2694 2002 2746
rect 2002 2694 2012 2746
rect 2036 2694 2066 2746
rect 2066 2694 2078 2746
rect 2078 2694 2092 2746
rect 2116 2694 2130 2746
rect 2130 2694 2142 2746
rect 2142 2694 2172 2746
rect 2196 2694 2206 2746
rect 2206 2694 2252 2746
rect 1956 2692 2012 2694
rect 2036 2692 2092 2694
rect 2116 2692 2172 2694
rect 2196 2692 2252 2694
rect 1306 2488 1362 2544
rect 3016 2202 3072 2204
rect 3096 2202 3152 2204
rect 3176 2202 3232 2204
rect 3256 2202 3312 2204
rect 3016 2150 3062 2202
rect 3062 2150 3072 2202
rect 3096 2150 3126 2202
rect 3126 2150 3138 2202
rect 3138 2150 3152 2202
rect 3176 2150 3190 2202
rect 3190 2150 3202 2202
rect 3202 2150 3232 2202
rect 3256 2150 3266 2202
rect 3266 2150 3312 2202
rect 3016 2148 3072 2150
rect 3096 2148 3152 2150
rect 3176 2148 3232 2150
rect 3256 2148 3312 2150
rect 1122 1400 1178 1456
rect 7956 2746 8012 2748
rect 8036 2746 8092 2748
rect 8116 2746 8172 2748
rect 8196 2746 8252 2748
rect 7956 2694 8002 2746
rect 8002 2694 8012 2746
rect 8036 2694 8066 2746
rect 8066 2694 8078 2746
rect 8078 2694 8092 2746
rect 8116 2694 8130 2746
rect 8130 2694 8142 2746
rect 8142 2694 8172 2746
rect 8196 2694 8206 2746
rect 8206 2694 8252 2746
rect 7956 2692 8012 2694
rect 8036 2692 8092 2694
rect 8116 2692 8172 2694
rect 8196 2692 8252 2694
rect 9016 3290 9072 3292
rect 9096 3290 9152 3292
rect 9176 3290 9232 3292
rect 9256 3290 9312 3292
rect 9016 3238 9062 3290
rect 9062 3238 9072 3290
rect 9096 3238 9126 3290
rect 9126 3238 9138 3290
rect 9138 3238 9152 3290
rect 9176 3238 9190 3290
rect 9190 3238 9202 3290
rect 9202 3238 9232 3290
rect 9256 3238 9266 3290
rect 9266 3238 9312 3290
rect 9016 3236 9072 3238
rect 9096 3236 9152 3238
rect 9176 3236 9232 3238
rect 9256 3236 9312 3238
rect 9402 2352 9458 2408
rect 9016 2202 9072 2204
rect 9096 2202 9152 2204
rect 9176 2202 9232 2204
rect 9256 2202 9312 2204
rect 9016 2150 9062 2202
rect 9062 2150 9072 2202
rect 9096 2150 9126 2202
rect 9126 2150 9138 2202
rect 9138 2150 9152 2202
rect 9176 2150 9190 2202
rect 9190 2150 9202 2202
rect 9202 2150 9232 2202
rect 9256 2150 9266 2202
rect 9266 2150 9312 2202
rect 9016 2148 9072 2150
rect 9096 2148 9152 2150
rect 9176 2148 9232 2150
rect 9256 2148 9312 2150
rect 15016 5466 15072 5468
rect 15096 5466 15152 5468
rect 15176 5466 15232 5468
rect 15256 5466 15312 5468
rect 15016 5414 15062 5466
rect 15062 5414 15072 5466
rect 15096 5414 15126 5466
rect 15126 5414 15138 5466
rect 15138 5414 15152 5466
rect 15176 5414 15190 5466
rect 15190 5414 15202 5466
rect 15202 5414 15232 5466
rect 15256 5414 15266 5466
rect 15266 5414 15312 5466
rect 15016 5412 15072 5414
rect 15096 5412 15152 5414
rect 15176 5412 15232 5414
rect 15256 5412 15312 5414
rect 16118 9288 16174 9344
rect 16210 6840 16266 6896
rect 16026 6160 16082 6216
rect 16670 7792 16726 7848
rect 13956 4922 14012 4924
rect 14036 4922 14092 4924
rect 14116 4922 14172 4924
rect 14196 4922 14252 4924
rect 13956 4870 14002 4922
rect 14002 4870 14012 4922
rect 14036 4870 14066 4922
rect 14066 4870 14078 4922
rect 14078 4870 14092 4922
rect 14116 4870 14130 4922
rect 14130 4870 14142 4922
rect 14142 4870 14172 4922
rect 14196 4870 14206 4922
rect 14206 4870 14252 4922
rect 13956 4868 14012 4870
rect 14036 4868 14092 4870
rect 14116 4868 14172 4870
rect 14196 4868 14252 4870
rect 14922 4528 14978 4584
rect 13956 3834 14012 3836
rect 14036 3834 14092 3836
rect 14116 3834 14172 3836
rect 14196 3834 14252 3836
rect 13956 3782 14002 3834
rect 14002 3782 14012 3834
rect 14036 3782 14066 3834
rect 14066 3782 14078 3834
rect 14078 3782 14092 3834
rect 14116 3782 14130 3834
rect 14130 3782 14142 3834
rect 14142 3782 14172 3834
rect 14196 3782 14206 3834
rect 14206 3782 14252 3834
rect 13956 3780 14012 3782
rect 14036 3780 14092 3782
rect 14116 3780 14172 3782
rect 14196 3780 14252 3782
rect 15016 4378 15072 4380
rect 15096 4378 15152 4380
rect 15176 4378 15232 4380
rect 15256 4378 15312 4380
rect 15016 4326 15062 4378
rect 15062 4326 15072 4378
rect 15096 4326 15126 4378
rect 15126 4326 15138 4378
rect 15138 4326 15152 4378
rect 15176 4326 15190 4378
rect 15190 4326 15202 4378
rect 15202 4326 15232 4378
rect 15256 4326 15266 4378
rect 15266 4326 15312 4378
rect 15016 4324 15072 4326
rect 15096 4324 15152 4326
rect 15176 4324 15232 4326
rect 15256 4324 15312 4326
rect 15382 3848 15438 3904
rect 15016 3290 15072 3292
rect 15096 3290 15152 3292
rect 15176 3290 15232 3292
rect 15256 3290 15312 3292
rect 15016 3238 15062 3290
rect 15062 3238 15072 3290
rect 15096 3238 15126 3290
rect 15126 3238 15138 3290
rect 15138 3238 15152 3290
rect 15176 3238 15190 3290
rect 15190 3238 15202 3290
rect 15202 3238 15232 3290
rect 15256 3238 15266 3290
rect 15266 3238 15312 3290
rect 15016 3236 15072 3238
rect 15096 3236 15152 3238
rect 15176 3236 15232 3238
rect 15256 3236 15312 3238
rect 9586 1944 9642 2000
rect 9494 1672 9550 1728
rect 9034 176 9090 232
rect 10598 40 10654 96
rect 13956 2746 14012 2748
rect 14036 2746 14092 2748
rect 14116 2746 14172 2748
rect 14196 2746 14252 2748
rect 13956 2694 14002 2746
rect 14002 2694 14012 2746
rect 14036 2694 14066 2746
rect 14066 2694 14078 2746
rect 14078 2694 14092 2746
rect 14116 2694 14130 2746
rect 14130 2694 14142 2746
rect 14142 2694 14172 2746
rect 14196 2694 14206 2746
rect 14206 2694 14252 2746
rect 13956 2692 14012 2694
rect 14036 2692 14092 2694
rect 14116 2692 14172 2694
rect 14196 2692 14252 2694
rect 15016 2202 15072 2204
rect 15096 2202 15152 2204
rect 15176 2202 15232 2204
rect 15256 2202 15312 2204
rect 15016 2150 15062 2202
rect 15062 2150 15072 2202
rect 15096 2150 15126 2202
rect 15126 2150 15138 2202
rect 15138 2150 15152 2202
rect 15176 2150 15190 2202
rect 15190 2150 15202 2202
rect 15202 2150 15232 2202
rect 15256 2150 15266 2202
rect 15266 2150 15312 2202
rect 15016 2148 15072 2150
rect 15096 2148 15152 2150
rect 15176 2148 15232 2150
rect 15256 2148 15312 2150
rect 17866 5072 17922 5128
rect 16486 3440 16542 3496
rect 16854 3032 16910 3088
rect 16670 2896 16726 2952
rect 18142 7248 18198 7304
rect 19062 10376 19118 10432
rect 18510 8064 18566 8120
rect 19706 6704 19762 6760
rect 20718 9016 20774 9072
rect 20442 8880 20498 8936
rect 19956 8186 20012 8188
rect 20036 8186 20092 8188
rect 20116 8186 20172 8188
rect 20196 8186 20252 8188
rect 19956 8134 20002 8186
rect 20002 8134 20012 8186
rect 20036 8134 20066 8186
rect 20066 8134 20078 8186
rect 20078 8134 20092 8186
rect 20116 8134 20130 8186
rect 20130 8134 20142 8186
rect 20142 8134 20172 8186
rect 20196 8134 20206 8186
rect 20206 8134 20252 8186
rect 19956 8132 20012 8134
rect 20036 8132 20092 8134
rect 20116 8132 20172 8134
rect 20196 8132 20252 8134
rect 19956 7098 20012 7100
rect 20036 7098 20092 7100
rect 20116 7098 20172 7100
rect 20196 7098 20252 7100
rect 19956 7046 20002 7098
rect 20002 7046 20012 7098
rect 20036 7046 20066 7098
rect 20066 7046 20078 7098
rect 20078 7046 20092 7098
rect 20116 7046 20130 7098
rect 20130 7046 20142 7098
rect 20142 7046 20172 7098
rect 20196 7046 20206 7098
rect 20206 7046 20252 7098
rect 19956 7044 20012 7046
rect 20036 7044 20092 7046
rect 20116 7044 20172 7046
rect 20196 7044 20252 7046
rect 20902 9152 20958 9208
rect 21638 9424 21694 9480
rect 21016 8730 21072 8732
rect 21096 8730 21152 8732
rect 21176 8730 21232 8732
rect 21256 8730 21312 8732
rect 21016 8678 21062 8730
rect 21062 8678 21072 8730
rect 21096 8678 21126 8730
rect 21126 8678 21138 8730
rect 21138 8678 21152 8730
rect 21176 8678 21190 8730
rect 21190 8678 21202 8730
rect 21202 8678 21232 8730
rect 21256 8678 21266 8730
rect 21266 8678 21312 8730
rect 21016 8676 21072 8678
rect 21096 8676 21152 8678
rect 21176 8676 21232 8678
rect 21256 8676 21312 8678
rect 21016 7642 21072 7644
rect 21096 7642 21152 7644
rect 21176 7642 21232 7644
rect 21256 7642 21312 7644
rect 21016 7590 21062 7642
rect 21062 7590 21072 7642
rect 21096 7590 21126 7642
rect 21126 7590 21138 7642
rect 21138 7590 21152 7642
rect 21176 7590 21190 7642
rect 21190 7590 21202 7642
rect 21202 7590 21232 7642
rect 21256 7590 21266 7642
rect 21266 7590 21312 7642
rect 21016 7588 21072 7590
rect 21096 7588 21152 7590
rect 21176 7588 21232 7590
rect 21256 7588 21312 7590
rect 19956 6010 20012 6012
rect 20036 6010 20092 6012
rect 20116 6010 20172 6012
rect 20196 6010 20252 6012
rect 19956 5958 20002 6010
rect 20002 5958 20012 6010
rect 20036 5958 20066 6010
rect 20066 5958 20078 6010
rect 20078 5958 20092 6010
rect 20116 5958 20130 6010
rect 20130 5958 20142 6010
rect 20142 5958 20172 6010
rect 20196 5958 20206 6010
rect 20206 5958 20252 6010
rect 19956 5956 20012 5958
rect 20036 5956 20092 5958
rect 20116 5956 20172 5958
rect 20196 5956 20252 5958
rect 21016 6554 21072 6556
rect 21096 6554 21152 6556
rect 21176 6554 21232 6556
rect 21256 6554 21312 6556
rect 21016 6502 21062 6554
rect 21062 6502 21072 6554
rect 21096 6502 21126 6554
rect 21126 6502 21138 6554
rect 21138 6502 21152 6554
rect 21176 6502 21190 6554
rect 21190 6502 21202 6554
rect 21202 6502 21232 6554
rect 21256 6502 21266 6554
rect 21266 6502 21312 6554
rect 21016 6500 21072 6502
rect 21096 6500 21152 6502
rect 21176 6500 21232 6502
rect 21256 6500 21312 6502
rect 18142 4664 18198 4720
rect 17406 3612 17408 3632
rect 17408 3612 17460 3632
rect 17460 3612 17462 3632
rect 17406 3576 17462 3612
rect 19956 4922 20012 4924
rect 20036 4922 20092 4924
rect 20116 4922 20172 4924
rect 20196 4922 20252 4924
rect 19956 4870 20002 4922
rect 20002 4870 20012 4922
rect 20036 4870 20066 4922
rect 20066 4870 20078 4922
rect 20078 4870 20092 4922
rect 20116 4870 20130 4922
rect 20130 4870 20142 4922
rect 20142 4870 20172 4922
rect 20196 4870 20206 4922
rect 20206 4870 20252 4922
rect 19956 4868 20012 4870
rect 20036 4868 20092 4870
rect 20116 4868 20172 4870
rect 20196 4868 20252 4870
rect 19522 4120 19578 4176
rect 19956 3834 20012 3836
rect 20036 3834 20092 3836
rect 20116 3834 20172 3836
rect 20196 3834 20252 3836
rect 19956 3782 20002 3834
rect 20002 3782 20012 3834
rect 20036 3782 20066 3834
rect 20066 3782 20078 3834
rect 20078 3782 20092 3834
rect 20116 3782 20130 3834
rect 20130 3782 20142 3834
rect 20142 3782 20172 3834
rect 20196 3782 20206 3834
rect 20206 3782 20252 3834
rect 19956 3780 20012 3782
rect 20036 3780 20092 3782
rect 20116 3780 20172 3782
rect 20196 3780 20252 3782
rect 18510 3440 18566 3496
rect 19956 2746 20012 2748
rect 20036 2746 20092 2748
rect 20116 2746 20172 2748
rect 20196 2746 20252 2748
rect 19956 2694 20002 2746
rect 20002 2694 20012 2746
rect 20036 2694 20066 2746
rect 20066 2694 20078 2746
rect 20078 2694 20092 2746
rect 20116 2694 20130 2746
rect 20130 2694 20142 2746
rect 20142 2694 20172 2746
rect 20196 2694 20206 2746
rect 20206 2694 20252 2746
rect 19956 2692 20012 2694
rect 20036 2692 20092 2694
rect 20116 2692 20172 2694
rect 20196 2692 20252 2694
rect 21016 5466 21072 5468
rect 21096 5466 21152 5468
rect 21176 5466 21232 5468
rect 21256 5466 21312 5468
rect 21016 5414 21062 5466
rect 21062 5414 21072 5466
rect 21096 5414 21126 5466
rect 21126 5414 21138 5466
rect 21138 5414 21152 5466
rect 21176 5414 21190 5466
rect 21190 5414 21202 5466
rect 21202 5414 21232 5466
rect 21256 5414 21266 5466
rect 21266 5414 21312 5466
rect 21016 5412 21072 5414
rect 21096 5412 21152 5414
rect 21176 5412 21232 5414
rect 21256 5412 21312 5414
rect 21016 4378 21072 4380
rect 21096 4378 21152 4380
rect 21176 4378 21232 4380
rect 21256 4378 21312 4380
rect 21016 4326 21062 4378
rect 21062 4326 21072 4378
rect 21096 4326 21126 4378
rect 21126 4326 21138 4378
rect 21138 4326 21152 4378
rect 21176 4326 21190 4378
rect 21190 4326 21202 4378
rect 21202 4326 21232 4378
rect 21256 4326 21266 4378
rect 21266 4326 21312 4378
rect 21016 4324 21072 4326
rect 21096 4324 21152 4326
rect 21176 4324 21232 4326
rect 21256 4324 21312 4326
rect 21016 3290 21072 3292
rect 21096 3290 21152 3292
rect 21176 3290 21232 3292
rect 21256 3290 21312 3292
rect 21016 3238 21062 3290
rect 21062 3238 21072 3290
rect 21096 3238 21126 3290
rect 21126 3238 21138 3290
rect 21138 3238 21152 3290
rect 21176 3238 21190 3290
rect 21190 3238 21202 3290
rect 21202 3238 21232 3290
rect 21256 3238 21266 3290
rect 21266 3238 21312 3290
rect 21016 3236 21072 3238
rect 21096 3236 21152 3238
rect 21176 3236 21232 3238
rect 21256 3236 21312 3238
rect 21016 2202 21072 2204
rect 21096 2202 21152 2204
rect 21176 2202 21232 2204
rect 21256 2202 21312 2204
rect 21016 2150 21062 2202
rect 21062 2150 21072 2202
rect 21096 2150 21126 2202
rect 21126 2150 21138 2202
rect 21138 2150 21152 2202
rect 21176 2150 21190 2202
rect 21190 2150 21202 2202
rect 21202 2150 21232 2202
rect 21256 2150 21266 2202
rect 21266 2150 21312 2202
rect 21016 2148 21072 2150
rect 21096 2148 21152 2150
rect 21176 2148 21232 2150
rect 21256 2148 21312 2150
rect 22650 9016 22706 9072
rect 22834 6704 22890 6760
rect 23110 8200 23166 8256
rect 22466 176 22522 232
rect 23938 6704 23994 6760
rect 23754 3984 23810 4040
rect 24490 7928 24546 7984
rect 23478 3576 23534 3632
rect 26422 8472 26478 8528
rect 25956 8186 26012 8188
rect 26036 8186 26092 8188
rect 26116 8186 26172 8188
rect 26196 8186 26252 8188
rect 25956 8134 26002 8186
rect 26002 8134 26012 8186
rect 26036 8134 26066 8186
rect 26066 8134 26078 8186
rect 26078 8134 26092 8186
rect 26116 8134 26130 8186
rect 26130 8134 26142 8186
rect 26142 8134 26172 8186
rect 26196 8134 26206 8186
rect 26206 8134 26252 8186
rect 25956 8132 26012 8134
rect 26036 8132 26092 8134
rect 26116 8132 26172 8134
rect 26196 8132 26252 8134
rect 25778 7384 25834 7440
rect 25956 7098 26012 7100
rect 26036 7098 26092 7100
rect 26116 7098 26172 7100
rect 26196 7098 26252 7100
rect 25956 7046 26002 7098
rect 26002 7046 26012 7098
rect 26036 7046 26066 7098
rect 26066 7046 26078 7098
rect 26078 7046 26092 7098
rect 26116 7046 26130 7098
rect 26130 7046 26142 7098
rect 26142 7046 26172 7098
rect 26196 7046 26206 7098
rect 26206 7046 26252 7098
rect 25956 7044 26012 7046
rect 26036 7044 26092 7046
rect 26116 7044 26172 7046
rect 26196 7044 26252 7046
rect 25956 6010 26012 6012
rect 26036 6010 26092 6012
rect 26116 6010 26172 6012
rect 26196 6010 26252 6012
rect 25956 5958 26002 6010
rect 26002 5958 26012 6010
rect 26036 5958 26066 6010
rect 26066 5958 26078 6010
rect 26078 5958 26092 6010
rect 26116 5958 26130 6010
rect 26130 5958 26142 6010
rect 26142 5958 26172 6010
rect 26196 5958 26206 6010
rect 26206 5958 26252 6010
rect 25956 5956 26012 5958
rect 26036 5956 26092 5958
rect 26116 5956 26172 5958
rect 26196 5956 26252 5958
rect 25956 4922 26012 4924
rect 26036 4922 26092 4924
rect 26116 4922 26172 4924
rect 26196 4922 26252 4924
rect 25956 4870 26002 4922
rect 26002 4870 26012 4922
rect 26036 4870 26066 4922
rect 26066 4870 26078 4922
rect 26078 4870 26092 4922
rect 26116 4870 26130 4922
rect 26130 4870 26142 4922
rect 26142 4870 26172 4922
rect 26196 4870 26206 4922
rect 26206 4870 26252 4922
rect 25956 4868 26012 4870
rect 26036 4868 26092 4870
rect 26116 4868 26172 4870
rect 26196 4868 26252 4870
rect 25956 3834 26012 3836
rect 26036 3834 26092 3836
rect 26116 3834 26172 3836
rect 26196 3834 26252 3836
rect 25956 3782 26002 3834
rect 26002 3782 26012 3834
rect 26036 3782 26066 3834
rect 26066 3782 26078 3834
rect 26078 3782 26092 3834
rect 26116 3782 26130 3834
rect 26130 3782 26142 3834
rect 26142 3782 26172 3834
rect 26196 3782 26206 3834
rect 26206 3782 26252 3834
rect 25956 3780 26012 3782
rect 26036 3780 26092 3782
rect 26116 3780 26172 3782
rect 26196 3780 26252 3782
rect 25956 2746 26012 2748
rect 26036 2746 26092 2748
rect 26116 2746 26172 2748
rect 26196 2746 26252 2748
rect 25956 2694 26002 2746
rect 26002 2694 26012 2746
rect 26036 2694 26066 2746
rect 26066 2694 26078 2746
rect 26078 2694 26092 2746
rect 26116 2694 26130 2746
rect 26130 2694 26142 2746
rect 26142 2694 26172 2746
rect 26196 2694 26206 2746
rect 26206 2694 26252 2746
rect 25956 2692 26012 2694
rect 26036 2692 26092 2694
rect 26116 2692 26172 2694
rect 26196 2692 26252 2694
rect 25594 40 25650 96
rect 27016 8730 27072 8732
rect 27096 8730 27152 8732
rect 27176 8730 27232 8732
rect 27256 8730 27312 8732
rect 27016 8678 27062 8730
rect 27062 8678 27072 8730
rect 27096 8678 27126 8730
rect 27126 8678 27138 8730
rect 27138 8678 27152 8730
rect 27176 8678 27190 8730
rect 27190 8678 27202 8730
rect 27202 8678 27232 8730
rect 27256 8678 27266 8730
rect 27266 8678 27312 8730
rect 27016 8676 27072 8678
rect 27096 8676 27152 8678
rect 27176 8676 27232 8678
rect 27256 8676 27312 8678
rect 27016 7642 27072 7644
rect 27096 7642 27152 7644
rect 27176 7642 27232 7644
rect 27256 7642 27312 7644
rect 27016 7590 27062 7642
rect 27062 7590 27072 7642
rect 27096 7590 27126 7642
rect 27126 7590 27138 7642
rect 27138 7590 27152 7642
rect 27176 7590 27190 7642
rect 27190 7590 27202 7642
rect 27202 7590 27232 7642
rect 27256 7590 27266 7642
rect 27266 7590 27312 7642
rect 27016 7588 27072 7590
rect 27096 7588 27152 7590
rect 27176 7588 27232 7590
rect 27256 7588 27312 7590
rect 27016 6554 27072 6556
rect 27096 6554 27152 6556
rect 27176 6554 27232 6556
rect 27256 6554 27312 6556
rect 27016 6502 27062 6554
rect 27062 6502 27072 6554
rect 27096 6502 27126 6554
rect 27126 6502 27138 6554
rect 27138 6502 27152 6554
rect 27176 6502 27190 6554
rect 27190 6502 27202 6554
rect 27202 6502 27232 6554
rect 27256 6502 27266 6554
rect 27266 6502 27312 6554
rect 27016 6500 27072 6502
rect 27096 6500 27152 6502
rect 27176 6500 27232 6502
rect 27256 6500 27312 6502
rect 27016 5466 27072 5468
rect 27096 5466 27152 5468
rect 27176 5466 27232 5468
rect 27256 5466 27312 5468
rect 27016 5414 27062 5466
rect 27062 5414 27072 5466
rect 27096 5414 27126 5466
rect 27126 5414 27138 5466
rect 27138 5414 27152 5466
rect 27176 5414 27190 5466
rect 27190 5414 27202 5466
rect 27202 5414 27232 5466
rect 27256 5414 27266 5466
rect 27266 5414 27312 5466
rect 27016 5412 27072 5414
rect 27096 5412 27152 5414
rect 27176 5412 27232 5414
rect 27256 5412 27312 5414
rect 27016 4378 27072 4380
rect 27096 4378 27152 4380
rect 27176 4378 27232 4380
rect 27256 4378 27312 4380
rect 27016 4326 27062 4378
rect 27062 4326 27072 4378
rect 27096 4326 27126 4378
rect 27126 4326 27138 4378
rect 27138 4326 27152 4378
rect 27176 4326 27190 4378
rect 27190 4326 27202 4378
rect 27202 4326 27232 4378
rect 27256 4326 27266 4378
rect 27266 4326 27312 4378
rect 27016 4324 27072 4326
rect 27096 4324 27152 4326
rect 27176 4324 27232 4326
rect 27256 4324 27312 4326
rect 27016 3290 27072 3292
rect 27096 3290 27152 3292
rect 27176 3290 27232 3292
rect 27256 3290 27312 3292
rect 27016 3238 27062 3290
rect 27062 3238 27072 3290
rect 27096 3238 27126 3290
rect 27126 3238 27138 3290
rect 27138 3238 27152 3290
rect 27176 3238 27190 3290
rect 27190 3238 27202 3290
rect 27202 3238 27232 3290
rect 27256 3238 27266 3290
rect 27266 3238 27312 3290
rect 27016 3236 27072 3238
rect 27096 3236 27152 3238
rect 27176 3236 27232 3238
rect 27256 3236 27312 3238
rect 27016 2202 27072 2204
rect 27096 2202 27152 2204
rect 27176 2202 27232 2204
rect 27256 2202 27312 2204
rect 27016 2150 27062 2202
rect 27062 2150 27072 2202
rect 27096 2150 27126 2202
rect 27126 2150 27138 2202
rect 27138 2150 27152 2202
rect 27176 2150 27190 2202
rect 27190 2150 27202 2202
rect 27202 2150 27232 2202
rect 27256 2150 27266 2202
rect 27266 2150 27312 2202
rect 27016 2148 27072 2150
rect 27096 2148 27152 2150
rect 27176 2148 27232 2150
rect 27256 2148 27312 2150
rect 32310 9832 32366 9888
rect 30654 9560 30710 9616
rect 31482 9288 31538 9344
rect 31022 9016 31078 9072
rect 31390 8744 31446 8800
rect 31114 8472 31170 8528
rect 31956 8186 32012 8188
rect 32036 8186 32092 8188
rect 32116 8186 32172 8188
rect 32196 8186 32252 8188
rect 31956 8134 32002 8186
rect 32002 8134 32012 8186
rect 32036 8134 32066 8186
rect 32066 8134 32078 8186
rect 32078 8134 32092 8186
rect 32116 8134 32130 8186
rect 32130 8134 32142 8186
rect 32142 8134 32172 8186
rect 32196 8134 32206 8186
rect 32206 8134 32252 8186
rect 31956 8132 32012 8134
rect 32036 8132 32092 8134
rect 32116 8132 32172 8134
rect 32196 8132 32252 8134
rect 31850 7928 31906 7984
rect 32126 7692 32128 7712
rect 32128 7692 32180 7712
rect 32180 7692 32182 7712
rect 32126 7656 32182 7692
rect 31758 7384 31814 7440
rect 31956 7098 32012 7100
rect 32036 7098 32092 7100
rect 32116 7098 32172 7100
rect 32196 7098 32252 7100
rect 31956 7046 32002 7098
rect 32002 7046 32012 7098
rect 32036 7046 32066 7098
rect 32066 7046 32078 7098
rect 32078 7046 32092 7098
rect 32116 7046 32130 7098
rect 32130 7046 32142 7098
rect 32142 7046 32172 7098
rect 32196 7046 32206 7098
rect 32206 7046 32252 7098
rect 31956 7044 32012 7046
rect 32036 7044 32092 7046
rect 32116 7044 32172 7046
rect 32196 7044 32252 7046
rect 31758 6840 31814 6896
rect 31390 6604 31392 6624
rect 31392 6604 31444 6624
rect 31444 6604 31446 6624
rect 31390 6568 31446 6604
rect 30746 1944 30802 2000
rect 31482 6180 31538 6216
rect 31482 6160 31484 6180
rect 31484 6160 31536 6180
rect 31536 6160 31538 6180
rect 32586 8200 32642 8256
rect 32770 7148 32772 7168
rect 32772 7148 32824 7168
rect 32824 7148 32826 7168
rect 32770 7112 32826 7148
rect 31850 6296 31906 6352
rect 31956 6010 32012 6012
rect 32036 6010 32092 6012
rect 32116 6010 32172 6012
rect 32196 6010 32252 6012
rect 31956 5958 32002 6010
rect 32002 5958 32012 6010
rect 32036 5958 32066 6010
rect 32066 5958 32078 6010
rect 32078 5958 32092 6010
rect 32116 5958 32130 6010
rect 32130 5958 32142 6010
rect 32142 5958 32172 6010
rect 32196 5958 32206 6010
rect 32206 5958 32252 6010
rect 31956 5956 32012 5958
rect 32036 5956 32092 5958
rect 32116 5956 32172 5958
rect 32196 5956 32252 5958
rect 32126 5788 32128 5808
rect 32128 5788 32180 5808
rect 32180 5788 32182 5808
rect 31758 5516 31760 5536
rect 31760 5516 31812 5536
rect 31812 5516 31814 5536
rect 31758 5480 31814 5516
rect 31482 4664 31538 4720
rect 31758 4120 31814 4176
rect 32126 5752 32182 5788
rect 32034 5208 32090 5264
rect 31956 4922 32012 4924
rect 32036 4922 32092 4924
rect 32116 4922 32172 4924
rect 32196 4922 32252 4924
rect 31956 4870 32002 4922
rect 32002 4870 32012 4922
rect 32036 4870 32066 4922
rect 32066 4870 32078 4922
rect 32078 4870 32092 4922
rect 32116 4870 32130 4922
rect 32130 4870 32142 4922
rect 32142 4870 32172 4922
rect 32196 4870 32206 4922
rect 32206 4870 32252 4922
rect 31956 4868 32012 4870
rect 32036 4868 32092 4870
rect 32116 4868 32172 4870
rect 32196 4868 32252 4870
rect 32126 4428 32128 4448
rect 32128 4428 32180 4448
rect 32180 4428 32182 4448
rect 32126 4392 32182 4428
rect 31956 3834 32012 3836
rect 32036 3834 32092 3836
rect 32116 3834 32172 3836
rect 32196 3834 32252 3836
rect 31956 3782 32002 3834
rect 32002 3782 32012 3834
rect 32036 3782 32066 3834
rect 32066 3782 32078 3834
rect 32078 3782 32092 3834
rect 32116 3782 32130 3834
rect 32130 3782 32142 3834
rect 32142 3782 32172 3834
rect 32196 3782 32206 3834
rect 32206 3782 32252 3834
rect 31956 3780 32012 3782
rect 32036 3780 32092 3782
rect 32116 3780 32172 3782
rect 32196 3780 32252 3782
rect 31482 3576 31538 3632
rect 31666 3440 31722 3496
rect 32126 3340 32128 3360
rect 32128 3340 32180 3360
rect 32180 3340 32182 3360
rect 32126 3304 32182 3340
rect 31758 3032 31814 3088
rect 31956 2746 32012 2748
rect 32036 2746 32092 2748
rect 32116 2746 32172 2748
rect 32196 2746 32252 2748
rect 31956 2694 32002 2746
rect 32002 2694 32012 2746
rect 32036 2694 32066 2746
rect 32066 2694 32078 2746
rect 32078 2694 32092 2746
rect 32116 2694 32130 2746
rect 32130 2694 32142 2746
rect 32142 2694 32172 2746
rect 32196 2694 32206 2746
rect 32206 2694 32252 2746
rect 31956 2692 32012 2694
rect 32036 2692 32092 2694
rect 32116 2692 32172 2694
rect 32196 2692 32252 2694
rect 31758 2488 31814 2544
rect 31850 2252 31852 2272
rect 31852 2252 31904 2272
rect 31904 2252 31906 2272
rect 31114 1672 31170 1728
rect 31850 2216 31906 2252
rect 31482 1400 31538 1456
rect 32862 4972 32864 4992
rect 32864 4972 32916 4992
rect 32916 4972 32918 4992
rect 32862 4936 32918 4972
rect 32862 3884 32864 3904
rect 32864 3884 32916 3904
rect 32916 3884 32918 3904
rect 32862 3848 32918 3884
rect 32862 2796 32864 2816
rect 32864 2796 32916 2816
rect 32916 2796 32918 2816
rect 32862 2760 32918 2796
<< metal3 >>
rect 6453 10842 6519 10845
rect 14917 10842 14983 10845
rect 6453 10840 14983 10842
rect 6453 10784 6458 10840
rect 6514 10784 14922 10840
rect 14978 10784 14983 10840
rect 6453 10782 14983 10784
rect 6453 10779 6519 10782
rect 14917 10779 14983 10782
rect 7005 10434 7071 10437
rect 19057 10434 19123 10437
rect 7005 10432 19123 10434
rect 7005 10376 7010 10432
rect 7066 10376 19062 10432
rect 19118 10376 19123 10432
rect 7005 10374 19123 10376
rect 7005 10371 7071 10374
rect 19057 10371 19123 10374
rect 7833 10026 7899 10029
rect 14641 10026 14707 10029
rect 7833 10024 14707 10026
rect 7833 9968 7838 10024
rect 7894 9968 14646 10024
rect 14702 9968 14707 10024
rect 7833 9966 14707 9968
rect 7833 9963 7899 9966
rect 14641 9963 14707 9966
rect 0 9890 120 9920
rect 13721 9890 13787 9893
rect 0 9888 13787 9890
rect 0 9832 13726 9888
rect 13782 9832 13787 9888
rect 0 9830 13787 9832
rect 0 9800 120 9830
rect 13721 9827 13787 9830
rect 32305 9890 32371 9893
rect 33630 9890 33750 9920
rect 32305 9888 33750 9890
rect 32305 9832 32310 9888
rect 32366 9832 33750 9888
rect 32305 9830 33750 9832
rect 32305 9827 32371 9830
rect 33630 9800 33750 9830
rect 7557 9754 7623 9757
rect 14365 9754 14431 9757
rect 7557 9752 14431 9754
rect 7557 9696 7562 9752
rect 7618 9696 14370 9752
rect 14426 9696 14431 9752
rect 7557 9694 14431 9696
rect 7557 9691 7623 9694
rect 14365 9691 14431 9694
rect 0 9618 120 9648
rect 10041 9618 10107 9621
rect 0 9616 10107 9618
rect 0 9560 10046 9616
rect 10102 9560 10107 9616
rect 0 9558 10107 9560
rect 0 9528 120 9558
rect 10041 9555 10107 9558
rect 30649 9618 30715 9621
rect 33630 9618 33750 9648
rect 30649 9616 33750 9618
rect 30649 9560 30654 9616
rect 30710 9560 33750 9616
rect 30649 9558 33750 9560
rect 30649 9555 30715 9558
rect 33630 9528 33750 9558
rect 14457 9482 14523 9485
rect 21633 9482 21699 9485
rect 14457 9480 21699 9482
rect 14457 9424 14462 9480
rect 14518 9424 21638 9480
rect 21694 9424 21699 9480
rect 14457 9422 21699 9424
rect 14457 9419 14523 9422
rect 21633 9419 21699 9422
rect 0 9346 120 9376
rect 16113 9346 16179 9349
rect 0 9344 16179 9346
rect 0 9288 16118 9344
rect 16174 9288 16179 9344
rect 0 9286 16179 9288
rect 0 9256 120 9286
rect 16113 9283 16179 9286
rect 31477 9346 31543 9349
rect 33630 9346 33750 9376
rect 31477 9344 33750 9346
rect 31477 9288 31482 9344
rect 31538 9288 33750 9344
rect 31477 9286 33750 9288
rect 31477 9283 31543 9286
rect 33630 9256 33750 9286
rect 11789 9210 11855 9213
rect 15469 9210 15535 9213
rect 20897 9210 20963 9213
rect 11789 9208 15535 9210
rect 11789 9152 11794 9208
rect 11850 9152 15474 9208
rect 15530 9152 15535 9208
rect 11789 9150 15535 9152
rect 11789 9147 11855 9150
rect 15469 9147 15535 9150
rect 20486 9208 20963 9210
rect 20486 9152 20902 9208
rect 20958 9152 20963 9208
rect 20486 9150 20963 9152
rect 0 9074 120 9104
rect 14457 9074 14523 9077
rect 20486 9074 20546 9150
rect 20897 9147 20963 9150
rect 0 9072 14523 9074
rect 0 9016 14462 9072
rect 14518 9016 14523 9072
rect 0 9014 14523 9016
rect 0 8984 120 9014
rect 14457 9011 14523 9014
rect 14598 9014 20546 9074
rect 20713 9074 20779 9077
rect 22645 9074 22711 9077
rect 20713 9072 22711 9074
rect 20713 9016 20718 9072
rect 20774 9016 22650 9072
rect 22706 9016 22711 9072
rect 20713 9014 22711 9016
rect 14598 8938 14658 9014
rect 20713 9011 20779 9014
rect 22645 9011 22711 9014
rect 31017 9074 31083 9077
rect 33630 9074 33750 9104
rect 31017 9072 33750 9074
rect 31017 9016 31022 9072
rect 31078 9016 33750 9072
rect 31017 9014 33750 9016
rect 31017 9011 31083 9014
rect 33630 8984 33750 9014
rect 20437 8938 20503 8941
rect 2730 8878 14658 8938
rect 14782 8936 20503 8938
rect 14782 8880 20442 8936
rect 20498 8880 20503 8936
rect 14782 8878 20503 8880
rect 0 8802 120 8832
rect 2730 8802 2790 8878
rect 0 8742 2790 8802
rect 12065 8802 12131 8805
rect 14782 8802 14842 8878
rect 20437 8875 20503 8878
rect 12065 8800 14842 8802
rect 12065 8744 12070 8800
rect 12126 8744 14842 8800
rect 12065 8742 14842 8744
rect 31385 8802 31451 8805
rect 33630 8802 33750 8832
rect 31385 8800 33750 8802
rect 31385 8744 31390 8800
rect 31446 8744 33750 8800
rect 31385 8742 33750 8744
rect 0 8712 120 8742
rect 12065 8739 12131 8742
rect 31385 8739 31451 8742
rect 3006 8736 3322 8737
rect 3006 8672 3012 8736
rect 3076 8672 3092 8736
rect 3156 8672 3172 8736
rect 3236 8672 3252 8736
rect 3316 8672 3322 8736
rect 3006 8671 3322 8672
rect 9006 8736 9322 8737
rect 9006 8672 9012 8736
rect 9076 8672 9092 8736
rect 9156 8672 9172 8736
rect 9236 8672 9252 8736
rect 9316 8672 9322 8736
rect 9006 8671 9322 8672
rect 15006 8736 15322 8737
rect 15006 8672 15012 8736
rect 15076 8672 15092 8736
rect 15156 8672 15172 8736
rect 15236 8672 15252 8736
rect 15316 8672 15322 8736
rect 15006 8671 15322 8672
rect 21006 8736 21322 8737
rect 21006 8672 21012 8736
rect 21076 8672 21092 8736
rect 21156 8672 21172 8736
rect 21236 8672 21252 8736
rect 21316 8672 21322 8736
rect 21006 8671 21322 8672
rect 27006 8736 27322 8737
rect 27006 8672 27012 8736
rect 27076 8672 27092 8736
rect 27156 8672 27172 8736
rect 27236 8672 27252 8736
rect 27316 8672 27322 8736
rect 33630 8712 33750 8742
rect 27006 8671 27322 8672
rect 0 8530 120 8560
rect 26417 8530 26483 8533
rect 0 8528 26483 8530
rect 0 8472 26422 8528
rect 26478 8472 26483 8528
rect 0 8470 26483 8472
rect 0 8440 120 8470
rect 26417 8467 26483 8470
rect 31109 8530 31175 8533
rect 33630 8530 33750 8560
rect 31109 8528 33750 8530
rect 31109 8472 31114 8528
rect 31170 8472 33750 8528
rect 31109 8470 33750 8472
rect 31109 8467 31175 8470
rect 33630 8440 33750 8470
rect 1718 8334 2514 8394
rect 0 8258 120 8288
rect 1718 8258 1778 8334
rect 0 8198 1778 8258
rect 2454 8258 2514 8334
rect 7790 8334 8402 8394
rect 7790 8258 7850 8334
rect 2454 8198 7850 8258
rect 8342 8258 8402 8334
rect 13678 8334 14474 8394
rect 13678 8258 13738 8334
rect 8342 8198 13738 8258
rect 14414 8258 14474 8334
rect 19750 8334 20546 8394
rect 19750 8258 19810 8334
rect 14414 8198 19810 8258
rect 20486 8258 20546 8334
rect 23105 8258 23171 8261
rect 20486 8256 23171 8258
rect 20486 8200 23110 8256
rect 23166 8200 23171 8256
rect 20486 8198 23171 8200
rect 0 8168 120 8198
rect 23105 8195 23171 8198
rect 32581 8258 32647 8261
rect 33630 8258 33750 8288
rect 32581 8256 33750 8258
rect 32581 8200 32586 8256
rect 32642 8200 33750 8256
rect 32581 8198 33750 8200
rect 32581 8195 32647 8198
rect 1946 8192 2262 8193
rect 1946 8128 1952 8192
rect 2016 8128 2032 8192
rect 2096 8128 2112 8192
rect 2176 8128 2192 8192
rect 2256 8128 2262 8192
rect 1946 8127 2262 8128
rect 7946 8192 8262 8193
rect 7946 8128 7952 8192
rect 8016 8128 8032 8192
rect 8096 8128 8112 8192
rect 8176 8128 8192 8192
rect 8256 8128 8262 8192
rect 7946 8127 8262 8128
rect 13946 8192 14262 8193
rect 13946 8128 13952 8192
rect 14016 8128 14032 8192
rect 14096 8128 14112 8192
rect 14176 8128 14192 8192
rect 14256 8128 14262 8192
rect 13946 8127 14262 8128
rect 19946 8192 20262 8193
rect 19946 8128 19952 8192
rect 20016 8128 20032 8192
rect 20096 8128 20112 8192
rect 20176 8128 20192 8192
rect 20256 8128 20262 8192
rect 19946 8127 20262 8128
rect 25946 8192 26262 8193
rect 25946 8128 25952 8192
rect 26016 8128 26032 8192
rect 26096 8128 26112 8192
rect 26176 8128 26192 8192
rect 26256 8128 26262 8192
rect 25946 8127 26262 8128
rect 31946 8192 32262 8193
rect 31946 8128 31952 8192
rect 32016 8128 32032 8192
rect 32096 8128 32112 8192
rect 32176 8128 32192 8192
rect 32256 8128 32262 8192
rect 33630 8168 33750 8198
rect 31946 8127 32262 8128
rect 14825 8122 14891 8125
rect 18505 8122 18571 8125
rect 14825 8120 18571 8122
rect 14825 8064 14830 8120
rect 14886 8064 18510 8120
rect 18566 8064 18571 8120
rect 14825 8062 18571 8064
rect 14825 8059 14891 8062
rect 18505 8059 18571 8062
rect 0 7986 120 8016
rect 24485 7986 24551 7989
rect 0 7984 24551 7986
rect 0 7928 24490 7984
rect 24546 7928 24551 7984
rect 0 7926 24551 7928
rect 0 7896 120 7926
rect 24485 7923 24551 7926
rect 31845 7986 31911 7989
rect 33630 7986 33750 8016
rect 31845 7984 33750 7986
rect 31845 7928 31850 7984
rect 31906 7928 33750 7984
rect 31845 7926 33750 7928
rect 31845 7923 31911 7926
rect 33630 7896 33750 7926
rect 16665 7850 16731 7853
rect 2730 7848 16731 7850
rect 2730 7792 16670 7848
rect 16726 7792 16731 7848
rect 2730 7790 16731 7792
rect 0 7714 120 7744
rect 2730 7714 2790 7790
rect 16665 7787 16731 7790
rect 0 7654 2790 7714
rect 9581 7714 9647 7717
rect 14825 7714 14891 7717
rect 9581 7712 14891 7714
rect 9581 7656 9586 7712
rect 9642 7656 14830 7712
rect 14886 7656 14891 7712
rect 9581 7654 14891 7656
rect 0 7624 120 7654
rect 9581 7651 9647 7654
rect 14825 7651 14891 7654
rect 32121 7714 32187 7717
rect 33630 7714 33750 7744
rect 32121 7712 33750 7714
rect 32121 7656 32126 7712
rect 32182 7656 33750 7712
rect 32121 7654 33750 7656
rect 32121 7651 32187 7654
rect 3006 7648 3322 7649
rect 3006 7584 3012 7648
rect 3076 7584 3092 7648
rect 3156 7584 3172 7648
rect 3236 7584 3252 7648
rect 3316 7584 3322 7648
rect 3006 7583 3322 7584
rect 9006 7648 9322 7649
rect 9006 7584 9012 7648
rect 9076 7584 9092 7648
rect 9156 7584 9172 7648
rect 9236 7584 9252 7648
rect 9316 7584 9322 7648
rect 9006 7583 9322 7584
rect 15006 7648 15322 7649
rect 15006 7584 15012 7648
rect 15076 7584 15092 7648
rect 15156 7584 15172 7648
rect 15236 7584 15252 7648
rect 15316 7584 15322 7648
rect 15006 7583 15322 7584
rect 21006 7648 21322 7649
rect 21006 7584 21012 7648
rect 21076 7584 21092 7648
rect 21156 7584 21172 7648
rect 21236 7584 21252 7648
rect 21316 7584 21322 7648
rect 21006 7583 21322 7584
rect 27006 7648 27322 7649
rect 27006 7584 27012 7648
rect 27076 7584 27092 7648
rect 27156 7584 27172 7648
rect 27236 7584 27252 7648
rect 27316 7584 27322 7648
rect 33630 7624 33750 7654
rect 27006 7583 27322 7584
rect 0 7442 120 7472
rect 25773 7442 25839 7445
rect 0 7440 25839 7442
rect 0 7384 25778 7440
rect 25834 7384 25839 7440
rect 0 7382 25839 7384
rect 0 7352 120 7382
rect 25773 7379 25839 7382
rect 31753 7442 31819 7445
rect 33630 7442 33750 7472
rect 31753 7440 33750 7442
rect 31753 7384 31758 7440
rect 31814 7384 33750 7440
rect 31753 7382 33750 7384
rect 31753 7379 31819 7382
rect 33630 7352 33750 7382
rect 9581 7306 9647 7309
rect 18137 7306 18203 7309
rect 1718 7246 8402 7306
rect 0 7170 120 7200
rect 1718 7170 1778 7246
rect 0 7110 1778 7170
rect 0 7080 120 7110
rect 1946 7104 2262 7105
rect 1946 7040 1952 7104
rect 2016 7040 2032 7104
rect 2096 7040 2112 7104
rect 2176 7040 2192 7104
rect 2256 7040 2262 7104
rect 1946 7039 2262 7040
rect 7946 7104 8262 7105
rect 7946 7040 7952 7104
rect 8016 7040 8032 7104
rect 8096 7040 8112 7104
rect 8176 7040 8192 7104
rect 8256 7040 8262 7104
rect 7946 7039 8262 7040
rect 8342 7034 8402 7246
rect 9581 7304 18203 7306
rect 9581 7248 9586 7304
rect 9642 7248 18142 7304
rect 18198 7248 18203 7304
rect 9581 7246 18203 7248
rect 9581 7243 9647 7246
rect 18137 7243 18203 7246
rect 8845 7170 8911 7173
rect 9673 7170 9739 7173
rect 8845 7168 9739 7170
rect 8845 7112 8850 7168
rect 8906 7112 9678 7168
rect 9734 7112 9739 7168
rect 8845 7110 9739 7112
rect 8845 7107 8911 7110
rect 9673 7107 9739 7110
rect 32765 7170 32831 7173
rect 33630 7170 33750 7200
rect 32765 7168 33750 7170
rect 32765 7112 32770 7168
rect 32826 7112 33750 7168
rect 32765 7110 33750 7112
rect 32765 7107 32831 7110
rect 13946 7104 14262 7105
rect 13946 7040 13952 7104
rect 14016 7040 14032 7104
rect 14096 7040 14112 7104
rect 14176 7040 14192 7104
rect 14256 7040 14262 7104
rect 13946 7039 14262 7040
rect 19946 7104 20262 7105
rect 19946 7040 19952 7104
rect 20016 7040 20032 7104
rect 20096 7040 20112 7104
rect 20176 7040 20192 7104
rect 20256 7040 20262 7104
rect 19946 7039 20262 7040
rect 25946 7104 26262 7105
rect 25946 7040 25952 7104
rect 26016 7040 26032 7104
rect 26096 7040 26112 7104
rect 26176 7040 26192 7104
rect 26256 7040 26262 7104
rect 25946 7039 26262 7040
rect 31946 7104 32262 7105
rect 31946 7040 31952 7104
rect 32016 7040 32032 7104
rect 32096 7040 32112 7104
rect 32176 7040 32192 7104
rect 32256 7040 32262 7104
rect 33630 7080 33750 7110
rect 31946 7039 32262 7040
rect 9857 7034 9923 7037
rect 8342 7032 9923 7034
rect 8342 6976 9862 7032
rect 9918 6976 9923 7032
rect 8342 6974 9923 6976
rect 9857 6971 9923 6974
rect 0 6898 120 6928
rect 16205 6898 16271 6901
rect 0 6896 16271 6898
rect 0 6840 16210 6896
rect 16266 6840 16271 6896
rect 0 6838 16271 6840
rect 0 6808 120 6838
rect 16205 6835 16271 6838
rect 31753 6898 31819 6901
rect 33630 6898 33750 6928
rect 31753 6896 33750 6898
rect 31753 6840 31758 6896
rect 31814 6840 33750 6896
rect 31753 6838 33750 6840
rect 31753 6835 31819 6838
rect 33630 6808 33750 6838
rect 10685 6762 10751 6765
rect 19701 6762 19767 6765
rect 10685 6760 19767 6762
rect 10685 6704 10690 6760
rect 10746 6704 19706 6760
rect 19762 6704 19767 6760
rect 10685 6702 19767 6704
rect 10685 6699 10751 6702
rect 19701 6699 19767 6702
rect 22829 6762 22895 6765
rect 23933 6762 23999 6765
rect 22829 6760 23999 6762
rect 22829 6704 22834 6760
rect 22890 6704 23938 6760
rect 23994 6704 23999 6760
rect 22829 6702 23999 6704
rect 22829 6699 22895 6702
rect 23933 6699 23999 6702
rect 0 6626 120 6656
rect 565 6626 631 6629
rect 0 6624 631 6626
rect 0 6568 570 6624
rect 626 6568 631 6624
rect 0 6566 631 6568
rect 0 6536 120 6566
rect 565 6563 631 6566
rect 31385 6626 31451 6629
rect 33630 6626 33750 6656
rect 31385 6624 33750 6626
rect 31385 6568 31390 6624
rect 31446 6568 33750 6624
rect 31385 6566 33750 6568
rect 31385 6563 31451 6566
rect 3006 6560 3322 6561
rect 3006 6496 3012 6560
rect 3076 6496 3092 6560
rect 3156 6496 3172 6560
rect 3236 6496 3252 6560
rect 3316 6496 3322 6560
rect 3006 6495 3322 6496
rect 9006 6560 9322 6561
rect 9006 6496 9012 6560
rect 9076 6496 9092 6560
rect 9156 6496 9172 6560
rect 9236 6496 9252 6560
rect 9316 6496 9322 6560
rect 9006 6495 9322 6496
rect 15006 6560 15322 6561
rect 15006 6496 15012 6560
rect 15076 6496 15092 6560
rect 15156 6496 15172 6560
rect 15236 6496 15252 6560
rect 15316 6496 15322 6560
rect 15006 6495 15322 6496
rect 21006 6560 21322 6561
rect 21006 6496 21012 6560
rect 21076 6496 21092 6560
rect 21156 6496 21172 6560
rect 21236 6496 21252 6560
rect 21316 6496 21322 6560
rect 21006 6495 21322 6496
rect 27006 6560 27322 6561
rect 27006 6496 27012 6560
rect 27076 6496 27092 6560
rect 27156 6496 27172 6560
rect 27236 6496 27252 6560
rect 27316 6496 27322 6560
rect 33630 6536 33750 6566
rect 27006 6495 27322 6496
rect 9765 6490 9831 6493
rect 10593 6490 10659 6493
rect 9765 6488 10659 6490
rect 9765 6432 9770 6488
rect 9826 6432 10598 6488
rect 10654 6432 10659 6488
rect 9765 6430 10659 6432
rect 9765 6427 9831 6430
rect 10593 6427 10659 6430
rect 0 6354 120 6384
rect 12433 6354 12499 6357
rect 0 6352 12499 6354
rect 0 6296 12438 6352
rect 12494 6296 12499 6352
rect 0 6294 12499 6296
rect 0 6264 120 6294
rect 12433 6291 12499 6294
rect 31845 6354 31911 6357
rect 33630 6354 33750 6384
rect 31845 6352 33750 6354
rect 31845 6296 31850 6352
rect 31906 6296 33750 6352
rect 31845 6294 33750 6296
rect 31845 6291 31911 6294
rect 33630 6264 33750 6294
rect 4613 6218 4679 6221
rect 1718 6216 4679 6218
rect 1718 6160 4618 6216
rect 4674 6160 4679 6216
rect 1718 6158 4679 6160
rect 0 6082 120 6112
rect 1718 6082 1778 6158
rect 4613 6155 4679 6158
rect 9121 6218 9187 6221
rect 16021 6218 16087 6221
rect 9121 6216 16087 6218
rect 9121 6160 9126 6216
rect 9182 6160 16026 6216
rect 16082 6160 16087 6216
rect 9121 6158 16087 6160
rect 9121 6155 9187 6158
rect 16021 6155 16087 6158
rect 31477 6218 31543 6221
rect 31477 6216 32690 6218
rect 31477 6160 31482 6216
rect 31538 6160 32690 6216
rect 31477 6158 32690 6160
rect 31477 6155 31543 6158
rect 0 6022 1778 6082
rect 32630 6082 32690 6158
rect 33630 6082 33750 6112
rect 32630 6022 33750 6082
rect 0 5992 120 6022
rect 1946 6016 2262 6017
rect 1946 5952 1952 6016
rect 2016 5952 2032 6016
rect 2096 5952 2112 6016
rect 2176 5952 2192 6016
rect 2256 5952 2262 6016
rect 1946 5951 2262 5952
rect 7946 6016 8262 6017
rect 7946 5952 7952 6016
rect 8016 5952 8032 6016
rect 8096 5952 8112 6016
rect 8176 5952 8192 6016
rect 8256 5952 8262 6016
rect 7946 5951 8262 5952
rect 13946 6016 14262 6017
rect 13946 5952 13952 6016
rect 14016 5952 14032 6016
rect 14096 5952 14112 6016
rect 14176 5952 14192 6016
rect 14256 5952 14262 6016
rect 13946 5951 14262 5952
rect 19946 6016 20262 6017
rect 19946 5952 19952 6016
rect 20016 5952 20032 6016
rect 20096 5952 20112 6016
rect 20176 5952 20192 6016
rect 20256 5952 20262 6016
rect 19946 5951 20262 5952
rect 25946 6016 26262 6017
rect 25946 5952 25952 6016
rect 26016 5952 26032 6016
rect 26096 5952 26112 6016
rect 26176 5952 26192 6016
rect 26256 5952 26262 6016
rect 25946 5951 26262 5952
rect 31946 6016 32262 6017
rect 31946 5952 31952 6016
rect 32016 5952 32032 6016
rect 32096 5952 32112 6016
rect 32176 5952 32192 6016
rect 32256 5952 32262 6016
rect 33630 5992 33750 6022
rect 31946 5951 32262 5952
rect 0 5810 120 5840
rect 13721 5810 13787 5813
rect 0 5808 13787 5810
rect 0 5752 13726 5808
rect 13782 5752 13787 5808
rect 0 5750 13787 5752
rect 0 5720 120 5750
rect 13721 5747 13787 5750
rect 32121 5810 32187 5813
rect 33630 5810 33750 5840
rect 32121 5808 33750 5810
rect 32121 5752 32126 5808
rect 32182 5752 33750 5808
rect 32121 5750 33750 5752
rect 32121 5747 32187 5750
rect 33630 5720 33750 5750
rect 0 5538 120 5568
rect 31753 5538 31819 5541
rect 33630 5538 33750 5568
rect 0 5478 2790 5538
rect 0 5448 120 5478
rect 0 5266 120 5296
rect 1301 5266 1367 5269
rect 0 5264 1367 5266
rect 0 5208 1306 5264
rect 1362 5208 1367 5264
rect 0 5206 1367 5208
rect 2730 5266 2790 5478
rect 31753 5536 33750 5538
rect 31753 5480 31758 5536
rect 31814 5480 33750 5536
rect 31753 5478 33750 5480
rect 31753 5475 31819 5478
rect 3006 5472 3322 5473
rect 3006 5408 3012 5472
rect 3076 5408 3092 5472
rect 3156 5408 3172 5472
rect 3236 5408 3252 5472
rect 3316 5408 3322 5472
rect 3006 5407 3322 5408
rect 9006 5472 9322 5473
rect 9006 5408 9012 5472
rect 9076 5408 9092 5472
rect 9156 5408 9172 5472
rect 9236 5408 9252 5472
rect 9316 5408 9322 5472
rect 9006 5407 9322 5408
rect 15006 5472 15322 5473
rect 15006 5408 15012 5472
rect 15076 5408 15092 5472
rect 15156 5408 15172 5472
rect 15236 5408 15252 5472
rect 15316 5408 15322 5472
rect 15006 5407 15322 5408
rect 21006 5472 21322 5473
rect 21006 5408 21012 5472
rect 21076 5408 21092 5472
rect 21156 5408 21172 5472
rect 21236 5408 21252 5472
rect 21316 5408 21322 5472
rect 21006 5407 21322 5408
rect 27006 5472 27322 5473
rect 27006 5408 27012 5472
rect 27076 5408 27092 5472
rect 27156 5408 27172 5472
rect 27236 5408 27252 5472
rect 27316 5408 27322 5472
rect 33630 5448 33750 5478
rect 27006 5407 27322 5408
rect 6913 5266 6979 5269
rect 2730 5264 6979 5266
rect 2730 5208 6918 5264
rect 6974 5208 6979 5264
rect 2730 5206 6979 5208
rect 0 5176 120 5206
rect 1301 5203 1367 5206
rect 6913 5203 6979 5206
rect 32029 5266 32095 5269
rect 33630 5266 33750 5296
rect 32029 5264 33750 5266
rect 32029 5208 32034 5264
rect 32090 5208 33750 5264
rect 32029 5206 33750 5208
rect 32029 5203 32095 5206
rect 33630 5176 33750 5206
rect 2865 5130 2931 5133
rect 17861 5130 17927 5133
rect 2865 5128 17927 5130
rect 2865 5072 2870 5128
rect 2926 5072 17866 5128
rect 17922 5072 17927 5128
rect 2865 5070 17927 5072
rect 2865 5067 2931 5070
rect 17861 5067 17927 5070
rect 0 4994 120 5024
rect 1761 4994 1827 4997
rect 0 4992 1827 4994
rect 0 4936 1766 4992
rect 1822 4936 1827 4992
rect 0 4934 1827 4936
rect 0 4904 120 4934
rect 1761 4931 1827 4934
rect 32857 4994 32923 4997
rect 33630 4994 33750 5024
rect 32857 4992 33750 4994
rect 32857 4936 32862 4992
rect 32918 4936 33750 4992
rect 32857 4934 33750 4936
rect 32857 4931 32923 4934
rect 1946 4928 2262 4929
rect 1946 4864 1952 4928
rect 2016 4864 2032 4928
rect 2096 4864 2112 4928
rect 2176 4864 2192 4928
rect 2256 4864 2262 4928
rect 1946 4863 2262 4864
rect 7946 4928 8262 4929
rect 7946 4864 7952 4928
rect 8016 4864 8032 4928
rect 8096 4864 8112 4928
rect 8176 4864 8192 4928
rect 8256 4864 8262 4928
rect 7946 4863 8262 4864
rect 13946 4928 14262 4929
rect 13946 4864 13952 4928
rect 14016 4864 14032 4928
rect 14096 4864 14112 4928
rect 14176 4864 14192 4928
rect 14256 4864 14262 4928
rect 13946 4863 14262 4864
rect 19946 4928 20262 4929
rect 19946 4864 19952 4928
rect 20016 4864 20032 4928
rect 20096 4864 20112 4928
rect 20176 4864 20192 4928
rect 20256 4864 20262 4928
rect 19946 4863 20262 4864
rect 25946 4928 26262 4929
rect 25946 4864 25952 4928
rect 26016 4864 26032 4928
rect 26096 4864 26112 4928
rect 26176 4864 26192 4928
rect 26256 4864 26262 4928
rect 25946 4863 26262 4864
rect 31946 4928 32262 4929
rect 31946 4864 31952 4928
rect 32016 4864 32032 4928
rect 32096 4864 32112 4928
rect 32176 4864 32192 4928
rect 32256 4864 32262 4928
rect 33630 4904 33750 4934
rect 31946 4863 32262 4864
rect 0 4722 120 4752
rect 18137 4722 18203 4725
rect 0 4720 18203 4722
rect 0 4664 18142 4720
rect 18198 4664 18203 4720
rect 0 4662 18203 4664
rect 0 4632 120 4662
rect 18137 4659 18203 4662
rect 31477 4722 31543 4725
rect 33630 4722 33750 4752
rect 31477 4720 33750 4722
rect 31477 4664 31482 4720
rect 31538 4664 33750 4720
rect 31477 4662 33750 4664
rect 31477 4659 31543 4662
rect 33630 4632 33750 4662
rect 1761 4586 1827 4589
rect 14917 4586 14983 4589
rect 1761 4584 14983 4586
rect 1761 4528 1766 4584
rect 1822 4528 14922 4584
rect 14978 4528 14983 4584
rect 1761 4526 14983 4528
rect 1761 4523 1827 4526
rect 14917 4523 14983 4526
rect 0 4450 120 4480
rect 2865 4450 2931 4453
rect 0 4448 2931 4450
rect 0 4392 2870 4448
rect 2926 4392 2931 4448
rect 0 4390 2931 4392
rect 0 4360 120 4390
rect 2865 4387 2931 4390
rect 32121 4450 32187 4453
rect 33630 4450 33750 4480
rect 32121 4448 33750 4450
rect 32121 4392 32126 4448
rect 32182 4392 33750 4448
rect 32121 4390 33750 4392
rect 32121 4387 32187 4390
rect 3006 4384 3322 4385
rect 3006 4320 3012 4384
rect 3076 4320 3092 4384
rect 3156 4320 3172 4384
rect 3236 4320 3252 4384
rect 3316 4320 3322 4384
rect 3006 4319 3322 4320
rect 9006 4384 9322 4385
rect 9006 4320 9012 4384
rect 9076 4320 9092 4384
rect 9156 4320 9172 4384
rect 9236 4320 9252 4384
rect 9316 4320 9322 4384
rect 9006 4319 9322 4320
rect 15006 4384 15322 4385
rect 15006 4320 15012 4384
rect 15076 4320 15092 4384
rect 15156 4320 15172 4384
rect 15236 4320 15252 4384
rect 15316 4320 15322 4384
rect 15006 4319 15322 4320
rect 21006 4384 21322 4385
rect 21006 4320 21012 4384
rect 21076 4320 21092 4384
rect 21156 4320 21172 4384
rect 21236 4320 21252 4384
rect 21316 4320 21322 4384
rect 21006 4319 21322 4320
rect 27006 4384 27322 4385
rect 27006 4320 27012 4384
rect 27076 4320 27092 4384
rect 27156 4320 27172 4384
rect 27236 4320 27252 4384
rect 27316 4320 27322 4384
rect 33630 4360 33750 4390
rect 27006 4319 27322 4320
rect 0 4178 120 4208
rect 19517 4178 19583 4181
rect 0 4176 19583 4178
rect 0 4120 19522 4176
rect 19578 4120 19583 4176
rect 0 4118 19583 4120
rect 0 4088 120 4118
rect 19517 4115 19583 4118
rect 31753 4178 31819 4181
rect 33630 4178 33750 4208
rect 31753 4176 33750 4178
rect 31753 4120 31758 4176
rect 31814 4120 33750 4176
rect 31753 4118 33750 4120
rect 31753 4115 31819 4118
rect 33630 4088 33750 4118
rect 9397 4042 9463 4045
rect 1718 4040 9463 4042
rect 1718 3984 9402 4040
rect 9458 3984 9463 4040
rect 1718 3982 9463 3984
rect 0 3906 120 3936
rect 1718 3906 1778 3982
rect 9397 3979 9463 3982
rect 13629 4042 13695 4045
rect 23749 4042 23815 4045
rect 13629 4040 14474 4042
rect 13629 3984 13634 4040
rect 13690 3984 14474 4040
rect 13629 3982 14474 3984
rect 13629 3979 13695 3982
rect 0 3846 1778 3906
rect 0 3816 120 3846
rect 1946 3840 2262 3841
rect 1946 3776 1952 3840
rect 2016 3776 2032 3840
rect 2096 3776 2112 3840
rect 2176 3776 2192 3840
rect 2256 3776 2262 3840
rect 1946 3775 2262 3776
rect 7946 3840 8262 3841
rect 7946 3776 7952 3840
rect 8016 3776 8032 3840
rect 8096 3776 8112 3840
rect 8176 3776 8192 3840
rect 8256 3776 8262 3840
rect 7946 3775 8262 3776
rect 13946 3840 14262 3841
rect 13946 3776 13952 3840
rect 14016 3776 14032 3840
rect 14096 3776 14112 3840
rect 14176 3776 14192 3840
rect 14256 3776 14262 3840
rect 13946 3775 14262 3776
rect 14414 3770 14474 3982
rect 18462 4040 23815 4042
rect 18462 3984 23754 4040
rect 23810 3984 23815 4040
rect 18462 3982 23815 3984
rect 15377 3906 15443 3909
rect 18462 3906 18522 3982
rect 23749 3979 23815 3982
rect 15377 3904 18522 3906
rect 15377 3848 15382 3904
rect 15438 3848 18522 3904
rect 15377 3846 18522 3848
rect 32857 3906 32923 3909
rect 33630 3906 33750 3936
rect 32857 3904 33750 3906
rect 32857 3848 32862 3904
rect 32918 3848 33750 3904
rect 32857 3846 33750 3848
rect 15377 3843 15443 3846
rect 32857 3843 32923 3846
rect 19946 3840 20262 3841
rect 19946 3776 19952 3840
rect 20016 3776 20032 3840
rect 20096 3776 20112 3840
rect 20176 3776 20192 3840
rect 20256 3776 20262 3840
rect 19946 3775 20262 3776
rect 25946 3840 26262 3841
rect 25946 3776 25952 3840
rect 26016 3776 26032 3840
rect 26096 3776 26112 3840
rect 26176 3776 26192 3840
rect 26256 3776 26262 3840
rect 25946 3775 26262 3776
rect 31946 3840 32262 3841
rect 31946 3776 31952 3840
rect 32016 3776 32032 3840
rect 32096 3776 32112 3840
rect 32176 3776 32192 3840
rect 32256 3776 32262 3840
rect 33630 3816 33750 3846
rect 31946 3775 32262 3776
rect 14414 3710 17970 3770
rect 0 3634 120 3664
rect 17401 3634 17467 3637
rect 0 3632 17467 3634
rect 0 3576 17406 3632
rect 17462 3576 17467 3632
rect 0 3574 17467 3576
rect 17910 3634 17970 3710
rect 23473 3634 23539 3637
rect 17910 3632 23539 3634
rect 17910 3576 23478 3632
rect 23534 3576 23539 3632
rect 17910 3574 23539 3576
rect 0 3544 120 3574
rect 17401 3571 17467 3574
rect 23473 3571 23539 3574
rect 31477 3634 31543 3637
rect 33630 3634 33750 3664
rect 31477 3632 33750 3634
rect 31477 3576 31482 3632
rect 31538 3576 33750 3632
rect 31477 3574 33750 3576
rect 31477 3571 31543 3574
rect 33630 3544 33750 3574
rect 1761 3498 1827 3501
rect 16481 3498 16547 3501
rect 1761 3496 16547 3498
rect 1761 3440 1766 3496
rect 1822 3440 16486 3496
rect 16542 3440 16547 3496
rect 1761 3438 16547 3440
rect 1761 3435 1827 3438
rect 16481 3435 16547 3438
rect 18505 3498 18571 3501
rect 31661 3498 31727 3501
rect 18505 3496 31727 3498
rect 18505 3440 18510 3496
rect 18566 3440 31666 3496
rect 31722 3440 31727 3496
rect 18505 3438 31727 3440
rect 18505 3435 18571 3438
rect 31661 3435 31727 3438
rect 0 3362 120 3392
rect 1945 3362 2011 3365
rect 0 3360 2011 3362
rect 0 3304 1950 3360
rect 2006 3304 2011 3360
rect 0 3302 2011 3304
rect 0 3272 120 3302
rect 1945 3299 2011 3302
rect 32121 3362 32187 3365
rect 33630 3362 33750 3392
rect 32121 3360 33750 3362
rect 32121 3304 32126 3360
rect 32182 3304 33750 3360
rect 32121 3302 33750 3304
rect 32121 3299 32187 3302
rect 3006 3296 3322 3297
rect 3006 3232 3012 3296
rect 3076 3232 3092 3296
rect 3156 3232 3172 3296
rect 3236 3232 3252 3296
rect 3316 3232 3322 3296
rect 3006 3231 3322 3232
rect 9006 3296 9322 3297
rect 9006 3232 9012 3296
rect 9076 3232 9092 3296
rect 9156 3232 9172 3296
rect 9236 3232 9252 3296
rect 9316 3232 9322 3296
rect 9006 3231 9322 3232
rect 15006 3296 15322 3297
rect 15006 3232 15012 3296
rect 15076 3232 15092 3296
rect 15156 3232 15172 3296
rect 15236 3232 15252 3296
rect 15316 3232 15322 3296
rect 15006 3231 15322 3232
rect 21006 3296 21322 3297
rect 21006 3232 21012 3296
rect 21076 3232 21092 3296
rect 21156 3232 21172 3296
rect 21236 3232 21252 3296
rect 21316 3232 21322 3296
rect 21006 3231 21322 3232
rect 27006 3296 27322 3297
rect 27006 3232 27012 3296
rect 27076 3232 27092 3296
rect 27156 3232 27172 3296
rect 27236 3232 27252 3296
rect 27316 3232 27322 3296
rect 33630 3272 33750 3302
rect 27006 3231 27322 3232
rect 0 3090 120 3120
rect 16849 3090 16915 3093
rect 0 3088 16915 3090
rect 0 3032 16854 3088
rect 16910 3032 16915 3088
rect 0 3030 16915 3032
rect 0 3000 120 3030
rect 16849 3027 16915 3030
rect 31753 3090 31819 3093
rect 33630 3090 33750 3120
rect 31753 3088 33750 3090
rect 31753 3032 31758 3088
rect 31814 3032 33750 3088
rect 31753 3030 33750 3032
rect 31753 3027 31819 3030
rect 33630 3000 33750 3030
rect 1945 2954 2011 2957
rect 16665 2954 16731 2957
rect 1945 2952 16731 2954
rect 1945 2896 1950 2952
rect 2006 2896 16670 2952
rect 16726 2896 16731 2952
rect 1945 2894 16731 2896
rect 1945 2891 2011 2894
rect 16665 2891 16731 2894
rect 0 2818 120 2848
rect 1761 2818 1827 2821
rect 0 2816 1827 2818
rect 0 2760 1766 2816
rect 1822 2760 1827 2816
rect 0 2758 1827 2760
rect 0 2728 120 2758
rect 1761 2755 1827 2758
rect 32857 2818 32923 2821
rect 33630 2818 33750 2848
rect 32857 2816 33750 2818
rect 32857 2760 32862 2816
rect 32918 2760 33750 2816
rect 32857 2758 33750 2760
rect 32857 2755 32923 2758
rect 1946 2752 2262 2753
rect 1946 2688 1952 2752
rect 2016 2688 2032 2752
rect 2096 2688 2112 2752
rect 2176 2688 2192 2752
rect 2256 2688 2262 2752
rect 1946 2687 2262 2688
rect 7946 2752 8262 2753
rect 7946 2688 7952 2752
rect 8016 2688 8032 2752
rect 8096 2688 8112 2752
rect 8176 2688 8192 2752
rect 8256 2688 8262 2752
rect 7946 2687 8262 2688
rect 13946 2752 14262 2753
rect 13946 2688 13952 2752
rect 14016 2688 14032 2752
rect 14096 2688 14112 2752
rect 14176 2688 14192 2752
rect 14256 2688 14262 2752
rect 13946 2687 14262 2688
rect 19946 2752 20262 2753
rect 19946 2688 19952 2752
rect 20016 2688 20032 2752
rect 20096 2688 20112 2752
rect 20176 2688 20192 2752
rect 20256 2688 20262 2752
rect 19946 2687 20262 2688
rect 25946 2752 26262 2753
rect 25946 2688 25952 2752
rect 26016 2688 26032 2752
rect 26096 2688 26112 2752
rect 26176 2688 26192 2752
rect 26256 2688 26262 2752
rect 25946 2687 26262 2688
rect 31946 2752 32262 2753
rect 31946 2688 31952 2752
rect 32016 2688 32032 2752
rect 32096 2688 32112 2752
rect 32176 2688 32192 2752
rect 32256 2688 32262 2752
rect 33630 2728 33750 2758
rect 31946 2687 32262 2688
rect 0 2546 120 2576
rect 1301 2546 1367 2549
rect 0 2544 1367 2546
rect 0 2488 1306 2544
rect 1362 2488 1367 2544
rect 0 2486 1367 2488
rect 0 2456 120 2486
rect 1301 2483 1367 2486
rect 31753 2546 31819 2549
rect 33630 2546 33750 2576
rect 31753 2544 33750 2546
rect 31753 2488 31758 2544
rect 31814 2488 33750 2544
rect 31753 2486 33750 2488
rect 31753 2483 31819 2486
rect 33630 2456 33750 2486
rect 9397 2410 9463 2413
rect 2822 2408 9463 2410
rect 2822 2352 9402 2408
rect 9458 2352 9463 2408
rect 2822 2350 9463 2352
rect 0 2274 120 2304
rect 2822 2274 2882 2350
rect 9397 2347 9463 2350
rect 0 2214 2882 2274
rect 31845 2274 31911 2277
rect 33630 2274 33750 2304
rect 31845 2272 33750 2274
rect 31845 2216 31850 2272
rect 31906 2216 33750 2272
rect 31845 2214 33750 2216
rect 0 2184 120 2214
rect 31845 2211 31911 2214
rect 3006 2208 3322 2209
rect 3006 2144 3012 2208
rect 3076 2144 3092 2208
rect 3156 2144 3172 2208
rect 3236 2144 3252 2208
rect 3316 2144 3322 2208
rect 3006 2143 3322 2144
rect 9006 2208 9322 2209
rect 9006 2144 9012 2208
rect 9076 2144 9092 2208
rect 9156 2144 9172 2208
rect 9236 2144 9252 2208
rect 9316 2144 9322 2208
rect 9006 2143 9322 2144
rect 15006 2208 15322 2209
rect 15006 2144 15012 2208
rect 15076 2144 15092 2208
rect 15156 2144 15172 2208
rect 15236 2144 15252 2208
rect 15316 2144 15322 2208
rect 15006 2143 15322 2144
rect 21006 2208 21322 2209
rect 21006 2144 21012 2208
rect 21076 2144 21092 2208
rect 21156 2144 21172 2208
rect 21236 2144 21252 2208
rect 21316 2144 21322 2208
rect 21006 2143 21322 2144
rect 27006 2208 27322 2209
rect 27006 2144 27012 2208
rect 27076 2144 27092 2208
rect 27156 2144 27172 2208
rect 27236 2144 27252 2208
rect 27316 2144 27322 2208
rect 33630 2184 33750 2214
rect 27006 2143 27322 2144
rect 0 2002 120 2032
rect 9581 2002 9647 2005
rect 0 2000 9647 2002
rect 0 1944 9586 2000
rect 9642 1944 9647 2000
rect 0 1942 9647 1944
rect 0 1912 120 1942
rect 9581 1939 9647 1942
rect 30741 2002 30807 2005
rect 33630 2002 33750 2032
rect 30741 2000 33750 2002
rect 30741 1944 30746 2000
rect 30802 1944 33750 2000
rect 30741 1942 33750 1944
rect 30741 1939 30807 1942
rect 33630 1912 33750 1942
rect 0 1730 120 1760
rect 9489 1730 9555 1733
rect 0 1728 9555 1730
rect 0 1672 9494 1728
rect 9550 1672 9555 1728
rect 0 1670 9555 1672
rect 0 1640 120 1670
rect 9489 1667 9555 1670
rect 31109 1730 31175 1733
rect 33630 1730 33750 1760
rect 31109 1728 33750 1730
rect 31109 1672 31114 1728
rect 31170 1672 33750 1728
rect 31109 1670 33750 1672
rect 31109 1667 31175 1670
rect 33630 1640 33750 1670
rect 0 1458 120 1488
rect 1117 1458 1183 1461
rect 0 1456 1183 1458
rect 0 1400 1122 1456
rect 1178 1400 1183 1456
rect 0 1398 1183 1400
rect 0 1368 120 1398
rect 1117 1395 1183 1398
rect 31477 1458 31543 1461
rect 33630 1458 33750 1488
rect 31477 1456 33750 1458
rect 31477 1400 31482 1456
rect 31538 1400 33750 1456
rect 31477 1398 33750 1400
rect 31477 1395 31543 1398
rect 33630 1368 33750 1398
rect 9029 234 9095 237
rect 22461 234 22527 237
rect 9029 232 22527 234
rect 9029 176 9034 232
rect 9090 176 22466 232
rect 22522 176 22527 232
rect 9029 174 22527 176
rect 9029 171 9095 174
rect 22461 171 22527 174
rect 10593 98 10659 101
rect 25589 98 25655 101
rect 10593 96 25655 98
rect 10593 40 10598 96
rect 10654 40 25594 96
rect 25650 40 25655 96
rect 10593 38 25655 40
rect 10593 35 10659 38
rect 25589 35 25655 38
<< via3 >>
rect 3012 8732 3076 8736
rect 3012 8676 3016 8732
rect 3016 8676 3072 8732
rect 3072 8676 3076 8732
rect 3012 8672 3076 8676
rect 3092 8732 3156 8736
rect 3092 8676 3096 8732
rect 3096 8676 3152 8732
rect 3152 8676 3156 8732
rect 3092 8672 3156 8676
rect 3172 8732 3236 8736
rect 3172 8676 3176 8732
rect 3176 8676 3232 8732
rect 3232 8676 3236 8732
rect 3172 8672 3236 8676
rect 3252 8732 3316 8736
rect 3252 8676 3256 8732
rect 3256 8676 3312 8732
rect 3312 8676 3316 8732
rect 3252 8672 3316 8676
rect 9012 8732 9076 8736
rect 9012 8676 9016 8732
rect 9016 8676 9072 8732
rect 9072 8676 9076 8732
rect 9012 8672 9076 8676
rect 9092 8732 9156 8736
rect 9092 8676 9096 8732
rect 9096 8676 9152 8732
rect 9152 8676 9156 8732
rect 9092 8672 9156 8676
rect 9172 8732 9236 8736
rect 9172 8676 9176 8732
rect 9176 8676 9232 8732
rect 9232 8676 9236 8732
rect 9172 8672 9236 8676
rect 9252 8732 9316 8736
rect 9252 8676 9256 8732
rect 9256 8676 9312 8732
rect 9312 8676 9316 8732
rect 9252 8672 9316 8676
rect 15012 8732 15076 8736
rect 15012 8676 15016 8732
rect 15016 8676 15072 8732
rect 15072 8676 15076 8732
rect 15012 8672 15076 8676
rect 15092 8732 15156 8736
rect 15092 8676 15096 8732
rect 15096 8676 15152 8732
rect 15152 8676 15156 8732
rect 15092 8672 15156 8676
rect 15172 8732 15236 8736
rect 15172 8676 15176 8732
rect 15176 8676 15232 8732
rect 15232 8676 15236 8732
rect 15172 8672 15236 8676
rect 15252 8732 15316 8736
rect 15252 8676 15256 8732
rect 15256 8676 15312 8732
rect 15312 8676 15316 8732
rect 15252 8672 15316 8676
rect 21012 8732 21076 8736
rect 21012 8676 21016 8732
rect 21016 8676 21072 8732
rect 21072 8676 21076 8732
rect 21012 8672 21076 8676
rect 21092 8732 21156 8736
rect 21092 8676 21096 8732
rect 21096 8676 21152 8732
rect 21152 8676 21156 8732
rect 21092 8672 21156 8676
rect 21172 8732 21236 8736
rect 21172 8676 21176 8732
rect 21176 8676 21232 8732
rect 21232 8676 21236 8732
rect 21172 8672 21236 8676
rect 21252 8732 21316 8736
rect 21252 8676 21256 8732
rect 21256 8676 21312 8732
rect 21312 8676 21316 8732
rect 21252 8672 21316 8676
rect 27012 8732 27076 8736
rect 27012 8676 27016 8732
rect 27016 8676 27072 8732
rect 27072 8676 27076 8732
rect 27012 8672 27076 8676
rect 27092 8732 27156 8736
rect 27092 8676 27096 8732
rect 27096 8676 27152 8732
rect 27152 8676 27156 8732
rect 27092 8672 27156 8676
rect 27172 8732 27236 8736
rect 27172 8676 27176 8732
rect 27176 8676 27232 8732
rect 27232 8676 27236 8732
rect 27172 8672 27236 8676
rect 27252 8732 27316 8736
rect 27252 8676 27256 8732
rect 27256 8676 27312 8732
rect 27312 8676 27316 8732
rect 27252 8672 27316 8676
rect 1952 8188 2016 8192
rect 1952 8132 1956 8188
rect 1956 8132 2012 8188
rect 2012 8132 2016 8188
rect 1952 8128 2016 8132
rect 2032 8188 2096 8192
rect 2032 8132 2036 8188
rect 2036 8132 2092 8188
rect 2092 8132 2096 8188
rect 2032 8128 2096 8132
rect 2112 8188 2176 8192
rect 2112 8132 2116 8188
rect 2116 8132 2172 8188
rect 2172 8132 2176 8188
rect 2112 8128 2176 8132
rect 2192 8188 2256 8192
rect 2192 8132 2196 8188
rect 2196 8132 2252 8188
rect 2252 8132 2256 8188
rect 2192 8128 2256 8132
rect 7952 8188 8016 8192
rect 7952 8132 7956 8188
rect 7956 8132 8012 8188
rect 8012 8132 8016 8188
rect 7952 8128 8016 8132
rect 8032 8188 8096 8192
rect 8032 8132 8036 8188
rect 8036 8132 8092 8188
rect 8092 8132 8096 8188
rect 8032 8128 8096 8132
rect 8112 8188 8176 8192
rect 8112 8132 8116 8188
rect 8116 8132 8172 8188
rect 8172 8132 8176 8188
rect 8112 8128 8176 8132
rect 8192 8188 8256 8192
rect 8192 8132 8196 8188
rect 8196 8132 8252 8188
rect 8252 8132 8256 8188
rect 8192 8128 8256 8132
rect 13952 8188 14016 8192
rect 13952 8132 13956 8188
rect 13956 8132 14012 8188
rect 14012 8132 14016 8188
rect 13952 8128 14016 8132
rect 14032 8188 14096 8192
rect 14032 8132 14036 8188
rect 14036 8132 14092 8188
rect 14092 8132 14096 8188
rect 14032 8128 14096 8132
rect 14112 8188 14176 8192
rect 14112 8132 14116 8188
rect 14116 8132 14172 8188
rect 14172 8132 14176 8188
rect 14112 8128 14176 8132
rect 14192 8188 14256 8192
rect 14192 8132 14196 8188
rect 14196 8132 14252 8188
rect 14252 8132 14256 8188
rect 14192 8128 14256 8132
rect 19952 8188 20016 8192
rect 19952 8132 19956 8188
rect 19956 8132 20012 8188
rect 20012 8132 20016 8188
rect 19952 8128 20016 8132
rect 20032 8188 20096 8192
rect 20032 8132 20036 8188
rect 20036 8132 20092 8188
rect 20092 8132 20096 8188
rect 20032 8128 20096 8132
rect 20112 8188 20176 8192
rect 20112 8132 20116 8188
rect 20116 8132 20172 8188
rect 20172 8132 20176 8188
rect 20112 8128 20176 8132
rect 20192 8188 20256 8192
rect 20192 8132 20196 8188
rect 20196 8132 20252 8188
rect 20252 8132 20256 8188
rect 20192 8128 20256 8132
rect 25952 8188 26016 8192
rect 25952 8132 25956 8188
rect 25956 8132 26012 8188
rect 26012 8132 26016 8188
rect 25952 8128 26016 8132
rect 26032 8188 26096 8192
rect 26032 8132 26036 8188
rect 26036 8132 26092 8188
rect 26092 8132 26096 8188
rect 26032 8128 26096 8132
rect 26112 8188 26176 8192
rect 26112 8132 26116 8188
rect 26116 8132 26172 8188
rect 26172 8132 26176 8188
rect 26112 8128 26176 8132
rect 26192 8188 26256 8192
rect 26192 8132 26196 8188
rect 26196 8132 26252 8188
rect 26252 8132 26256 8188
rect 26192 8128 26256 8132
rect 31952 8188 32016 8192
rect 31952 8132 31956 8188
rect 31956 8132 32012 8188
rect 32012 8132 32016 8188
rect 31952 8128 32016 8132
rect 32032 8188 32096 8192
rect 32032 8132 32036 8188
rect 32036 8132 32092 8188
rect 32092 8132 32096 8188
rect 32032 8128 32096 8132
rect 32112 8188 32176 8192
rect 32112 8132 32116 8188
rect 32116 8132 32172 8188
rect 32172 8132 32176 8188
rect 32112 8128 32176 8132
rect 32192 8188 32256 8192
rect 32192 8132 32196 8188
rect 32196 8132 32252 8188
rect 32252 8132 32256 8188
rect 32192 8128 32256 8132
rect 3012 7644 3076 7648
rect 3012 7588 3016 7644
rect 3016 7588 3072 7644
rect 3072 7588 3076 7644
rect 3012 7584 3076 7588
rect 3092 7644 3156 7648
rect 3092 7588 3096 7644
rect 3096 7588 3152 7644
rect 3152 7588 3156 7644
rect 3092 7584 3156 7588
rect 3172 7644 3236 7648
rect 3172 7588 3176 7644
rect 3176 7588 3232 7644
rect 3232 7588 3236 7644
rect 3172 7584 3236 7588
rect 3252 7644 3316 7648
rect 3252 7588 3256 7644
rect 3256 7588 3312 7644
rect 3312 7588 3316 7644
rect 3252 7584 3316 7588
rect 9012 7644 9076 7648
rect 9012 7588 9016 7644
rect 9016 7588 9072 7644
rect 9072 7588 9076 7644
rect 9012 7584 9076 7588
rect 9092 7644 9156 7648
rect 9092 7588 9096 7644
rect 9096 7588 9152 7644
rect 9152 7588 9156 7644
rect 9092 7584 9156 7588
rect 9172 7644 9236 7648
rect 9172 7588 9176 7644
rect 9176 7588 9232 7644
rect 9232 7588 9236 7644
rect 9172 7584 9236 7588
rect 9252 7644 9316 7648
rect 9252 7588 9256 7644
rect 9256 7588 9312 7644
rect 9312 7588 9316 7644
rect 9252 7584 9316 7588
rect 15012 7644 15076 7648
rect 15012 7588 15016 7644
rect 15016 7588 15072 7644
rect 15072 7588 15076 7644
rect 15012 7584 15076 7588
rect 15092 7644 15156 7648
rect 15092 7588 15096 7644
rect 15096 7588 15152 7644
rect 15152 7588 15156 7644
rect 15092 7584 15156 7588
rect 15172 7644 15236 7648
rect 15172 7588 15176 7644
rect 15176 7588 15232 7644
rect 15232 7588 15236 7644
rect 15172 7584 15236 7588
rect 15252 7644 15316 7648
rect 15252 7588 15256 7644
rect 15256 7588 15312 7644
rect 15312 7588 15316 7644
rect 15252 7584 15316 7588
rect 21012 7644 21076 7648
rect 21012 7588 21016 7644
rect 21016 7588 21072 7644
rect 21072 7588 21076 7644
rect 21012 7584 21076 7588
rect 21092 7644 21156 7648
rect 21092 7588 21096 7644
rect 21096 7588 21152 7644
rect 21152 7588 21156 7644
rect 21092 7584 21156 7588
rect 21172 7644 21236 7648
rect 21172 7588 21176 7644
rect 21176 7588 21232 7644
rect 21232 7588 21236 7644
rect 21172 7584 21236 7588
rect 21252 7644 21316 7648
rect 21252 7588 21256 7644
rect 21256 7588 21312 7644
rect 21312 7588 21316 7644
rect 21252 7584 21316 7588
rect 27012 7644 27076 7648
rect 27012 7588 27016 7644
rect 27016 7588 27072 7644
rect 27072 7588 27076 7644
rect 27012 7584 27076 7588
rect 27092 7644 27156 7648
rect 27092 7588 27096 7644
rect 27096 7588 27152 7644
rect 27152 7588 27156 7644
rect 27092 7584 27156 7588
rect 27172 7644 27236 7648
rect 27172 7588 27176 7644
rect 27176 7588 27232 7644
rect 27232 7588 27236 7644
rect 27172 7584 27236 7588
rect 27252 7644 27316 7648
rect 27252 7588 27256 7644
rect 27256 7588 27312 7644
rect 27312 7588 27316 7644
rect 27252 7584 27316 7588
rect 1952 7100 2016 7104
rect 1952 7044 1956 7100
rect 1956 7044 2012 7100
rect 2012 7044 2016 7100
rect 1952 7040 2016 7044
rect 2032 7100 2096 7104
rect 2032 7044 2036 7100
rect 2036 7044 2092 7100
rect 2092 7044 2096 7100
rect 2032 7040 2096 7044
rect 2112 7100 2176 7104
rect 2112 7044 2116 7100
rect 2116 7044 2172 7100
rect 2172 7044 2176 7100
rect 2112 7040 2176 7044
rect 2192 7100 2256 7104
rect 2192 7044 2196 7100
rect 2196 7044 2252 7100
rect 2252 7044 2256 7100
rect 2192 7040 2256 7044
rect 7952 7100 8016 7104
rect 7952 7044 7956 7100
rect 7956 7044 8012 7100
rect 8012 7044 8016 7100
rect 7952 7040 8016 7044
rect 8032 7100 8096 7104
rect 8032 7044 8036 7100
rect 8036 7044 8092 7100
rect 8092 7044 8096 7100
rect 8032 7040 8096 7044
rect 8112 7100 8176 7104
rect 8112 7044 8116 7100
rect 8116 7044 8172 7100
rect 8172 7044 8176 7100
rect 8112 7040 8176 7044
rect 8192 7100 8256 7104
rect 8192 7044 8196 7100
rect 8196 7044 8252 7100
rect 8252 7044 8256 7100
rect 8192 7040 8256 7044
rect 13952 7100 14016 7104
rect 13952 7044 13956 7100
rect 13956 7044 14012 7100
rect 14012 7044 14016 7100
rect 13952 7040 14016 7044
rect 14032 7100 14096 7104
rect 14032 7044 14036 7100
rect 14036 7044 14092 7100
rect 14092 7044 14096 7100
rect 14032 7040 14096 7044
rect 14112 7100 14176 7104
rect 14112 7044 14116 7100
rect 14116 7044 14172 7100
rect 14172 7044 14176 7100
rect 14112 7040 14176 7044
rect 14192 7100 14256 7104
rect 14192 7044 14196 7100
rect 14196 7044 14252 7100
rect 14252 7044 14256 7100
rect 14192 7040 14256 7044
rect 19952 7100 20016 7104
rect 19952 7044 19956 7100
rect 19956 7044 20012 7100
rect 20012 7044 20016 7100
rect 19952 7040 20016 7044
rect 20032 7100 20096 7104
rect 20032 7044 20036 7100
rect 20036 7044 20092 7100
rect 20092 7044 20096 7100
rect 20032 7040 20096 7044
rect 20112 7100 20176 7104
rect 20112 7044 20116 7100
rect 20116 7044 20172 7100
rect 20172 7044 20176 7100
rect 20112 7040 20176 7044
rect 20192 7100 20256 7104
rect 20192 7044 20196 7100
rect 20196 7044 20252 7100
rect 20252 7044 20256 7100
rect 20192 7040 20256 7044
rect 25952 7100 26016 7104
rect 25952 7044 25956 7100
rect 25956 7044 26012 7100
rect 26012 7044 26016 7100
rect 25952 7040 26016 7044
rect 26032 7100 26096 7104
rect 26032 7044 26036 7100
rect 26036 7044 26092 7100
rect 26092 7044 26096 7100
rect 26032 7040 26096 7044
rect 26112 7100 26176 7104
rect 26112 7044 26116 7100
rect 26116 7044 26172 7100
rect 26172 7044 26176 7100
rect 26112 7040 26176 7044
rect 26192 7100 26256 7104
rect 26192 7044 26196 7100
rect 26196 7044 26252 7100
rect 26252 7044 26256 7100
rect 26192 7040 26256 7044
rect 31952 7100 32016 7104
rect 31952 7044 31956 7100
rect 31956 7044 32012 7100
rect 32012 7044 32016 7100
rect 31952 7040 32016 7044
rect 32032 7100 32096 7104
rect 32032 7044 32036 7100
rect 32036 7044 32092 7100
rect 32092 7044 32096 7100
rect 32032 7040 32096 7044
rect 32112 7100 32176 7104
rect 32112 7044 32116 7100
rect 32116 7044 32172 7100
rect 32172 7044 32176 7100
rect 32112 7040 32176 7044
rect 32192 7100 32256 7104
rect 32192 7044 32196 7100
rect 32196 7044 32252 7100
rect 32252 7044 32256 7100
rect 32192 7040 32256 7044
rect 3012 6556 3076 6560
rect 3012 6500 3016 6556
rect 3016 6500 3072 6556
rect 3072 6500 3076 6556
rect 3012 6496 3076 6500
rect 3092 6556 3156 6560
rect 3092 6500 3096 6556
rect 3096 6500 3152 6556
rect 3152 6500 3156 6556
rect 3092 6496 3156 6500
rect 3172 6556 3236 6560
rect 3172 6500 3176 6556
rect 3176 6500 3232 6556
rect 3232 6500 3236 6556
rect 3172 6496 3236 6500
rect 3252 6556 3316 6560
rect 3252 6500 3256 6556
rect 3256 6500 3312 6556
rect 3312 6500 3316 6556
rect 3252 6496 3316 6500
rect 9012 6556 9076 6560
rect 9012 6500 9016 6556
rect 9016 6500 9072 6556
rect 9072 6500 9076 6556
rect 9012 6496 9076 6500
rect 9092 6556 9156 6560
rect 9092 6500 9096 6556
rect 9096 6500 9152 6556
rect 9152 6500 9156 6556
rect 9092 6496 9156 6500
rect 9172 6556 9236 6560
rect 9172 6500 9176 6556
rect 9176 6500 9232 6556
rect 9232 6500 9236 6556
rect 9172 6496 9236 6500
rect 9252 6556 9316 6560
rect 9252 6500 9256 6556
rect 9256 6500 9312 6556
rect 9312 6500 9316 6556
rect 9252 6496 9316 6500
rect 15012 6556 15076 6560
rect 15012 6500 15016 6556
rect 15016 6500 15072 6556
rect 15072 6500 15076 6556
rect 15012 6496 15076 6500
rect 15092 6556 15156 6560
rect 15092 6500 15096 6556
rect 15096 6500 15152 6556
rect 15152 6500 15156 6556
rect 15092 6496 15156 6500
rect 15172 6556 15236 6560
rect 15172 6500 15176 6556
rect 15176 6500 15232 6556
rect 15232 6500 15236 6556
rect 15172 6496 15236 6500
rect 15252 6556 15316 6560
rect 15252 6500 15256 6556
rect 15256 6500 15312 6556
rect 15312 6500 15316 6556
rect 15252 6496 15316 6500
rect 21012 6556 21076 6560
rect 21012 6500 21016 6556
rect 21016 6500 21072 6556
rect 21072 6500 21076 6556
rect 21012 6496 21076 6500
rect 21092 6556 21156 6560
rect 21092 6500 21096 6556
rect 21096 6500 21152 6556
rect 21152 6500 21156 6556
rect 21092 6496 21156 6500
rect 21172 6556 21236 6560
rect 21172 6500 21176 6556
rect 21176 6500 21232 6556
rect 21232 6500 21236 6556
rect 21172 6496 21236 6500
rect 21252 6556 21316 6560
rect 21252 6500 21256 6556
rect 21256 6500 21312 6556
rect 21312 6500 21316 6556
rect 21252 6496 21316 6500
rect 27012 6556 27076 6560
rect 27012 6500 27016 6556
rect 27016 6500 27072 6556
rect 27072 6500 27076 6556
rect 27012 6496 27076 6500
rect 27092 6556 27156 6560
rect 27092 6500 27096 6556
rect 27096 6500 27152 6556
rect 27152 6500 27156 6556
rect 27092 6496 27156 6500
rect 27172 6556 27236 6560
rect 27172 6500 27176 6556
rect 27176 6500 27232 6556
rect 27232 6500 27236 6556
rect 27172 6496 27236 6500
rect 27252 6556 27316 6560
rect 27252 6500 27256 6556
rect 27256 6500 27312 6556
rect 27312 6500 27316 6556
rect 27252 6496 27316 6500
rect 1952 6012 2016 6016
rect 1952 5956 1956 6012
rect 1956 5956 2012 6012
rect 2012 5956 2016 6012
rect 1952 5952 2016 5956
rect 2032 6012 2096 6016
rect 2032 5956 2036 6012
rect 2036 5956 2092 6012
rect 2092 5956 2096 6012
rect 2032 5952 2096 5956
rect 2112 6012 2176 6016
rect 2112 5956 2116 6012
rect 2116 5956 2172 6012
rect 2172 5956 2176 6012
rect 2112 5952 2176 5956
rect 2192 6012 2256 6016
rect 2192 5956 2196 6012
rect 2196 5956 2252 6012
rect 2252 5956 2256 6012
rect 2192 5952 2256 5956
rect 7952 6012 8016 6016
rect 7952 5956 7956 6012
rect 7956 5956 8012 6012
rect 8012 5956 8016 6012
rect 7952 5952 8016 5956
rect 8032 6012 8096 6016
rect 8032 5956 8036 6012
rect 8036 5956 8092 6012
rect 8092 5956 8096 6012
rect 8032 5952 8096 5956
rect 8112 6012 8176 6016
rect 8112 5956 8116 6012
rect 8116 5956 8172 6012
rect 8172 5956 8176 6012
rect 8112 5952 8176 5956
rect 8192 6012 8256 6016
rect 8192 5956 8196 6012
rect 8196 5956 8252 6012
rect 8252 5956 8256 6012
rect 8192 5952 8256 5956
rect 13952 6012 14016 6016
rect 13952 5956 13956 6012
rect 13956 5956 14012 6012
rect 14012 5956 14016 6012
rect 13952 5952 14016 5956
rect 14032 6012 14096 6016
rect 14032 5956 14036 6012
rect 14036 5956 14092 6012
rect 14092 5956 14096 6012
rect 14032 5952 14096 5956
rect 14112 6012 14176 6016
rect 14112 5956 14116 6012
rect 14116 5956 14172 6012
rect 14172 5956 14176 6012
rect 14112 5952 14176 5956
rect 14192 6012 14256 6016
rect 14192 5956 14196 6012
rect 14196 5956 14252 6012
rect 14252 5956 14256 6012
rect 14192 5952 14256 5956
rect 19952 6012 20016 6016
rect 19952 5956 19956 6012
rect 19956 5956 20012 6012
rect 20012 5956 20016 6012
rect 19952 5952 20016 5956
rect 20032 6012 20096 6016
rect 20032 5956 20036 6012
rect 20036 5956 20092 6012
rect 20092 5956 20096 6012
rect 20032 5952 20096 5956
rect 20112 6012 20176 6016
rect 20112 5956 20116 6012
rect 20116 5956 20172 6012
rect 20172 5956 20176 6012
rect 20112 5952 20176 5956
rect 20192 6012 20256 6016
rect 20192 5956 20196 6012
rect 20196 5956 20252 6012
rect 20252 5956 20256 6012
rect 20192 5952 20256 5956
rect 25952 6012 26016 6016
rect 25952 5956 25956 6012
rect 25956 5956 26012 6012
rect 26012 5956 26016 6012
rect 25952 5952 26016 5956
rect 26032 6012 26096 6016
rect 26032 5956 26036 6012
rect 26036 5956 26092 6012
rect 26092 5956 26096 6012
rect 26032 5952 26096 5956
rect 26112 6012 26176 6016
rect 26112 5956 26116 6012
rect 26116 5956 26172 6012
rect 26172 5956 26176 6012
rect 26112 5952 26176 5956
rect 26192 6012 26256 6016
rect 26192 5956 26196 6012
rect 26196 5956 26252 6012
rect 26252 5956 26256 6012
rect 26192 5952 26256 5956
rect 31952 6012 32016 6016
rect 31952 5956 31956 6012
rect 31956 5956 32012 6012
rect 32012 5956 32016 6012
rect 31952 5952 32016 5956
rect 32032 6012 32096 6016
rect 32032 5956 32036 6012
rect 32036 5956 32092 6012
rect 32092 5956 32096 6012
rect 32032 5952 32096 5956
rect 32112 6012 32176 6016
rect 32112 5956 32116 6012
rect 32116 5956 32172 6012
rect 32172 5956 32176 6012
rect 32112 5952 32176 5956
rect 32192 6012 32256 6016
rect 32192 5956 32196 6012
rect 32196 5956 32252 6012
rect 32252 5956 32256 6012
rect 32192 5952 32256 5956
rect 3012 5468 3076 5472
rect 3012 5412 3016 5468
rect 3016 5412 3072 5468
rect 3072 5412 3076 5468
rect 3012 5408 3076 5412
rect 3092 5468 3156 5472
rect 3092 5412 3096 5468
rect 3096 5412 3152 5468
rect 3152 5412 3156 5468
rect 3092 5408 3156 5412
rect 3172 5468 3236 5472
rect 3172 5412 3176 5468
rect 3176 5412 3232 5468
rect 3232 5412 3236 5468
rect 3172 5408 3236 5412
rect 3252 5468 3316 5472
rect 3252 5412 3256 5468
rect 3256 5412 3312 5468
rect 3312 5412 3316 5468
rect 3252 5408 3316 5412
rect 9012 5468 9076 5472
rect 9012 5412 9016 5468
rect 9016 5412 9072 5468
rect 9072 5412 9076 5468
rect 9012 5408 9076 5412
rect 9092 5468 9156 5472
rect 9092 5412 9096 5468
rect 9096 5412 9152 5468
rect 9152 5412 9156 5468
rect 9092 5408 9156 5412
rect 9172 5468 9236 5472
rect 9172 5412 9176 5468
rect 9176 5412 9232 5468
rect 9232 5412 9236 5468
rect 9172 5408 9236 5412
rect 9252 5468 9316 5472
rect 9252 5412 9256 5468
rect 9256 5412 9312 5468
rect 9312 5412 9316 5468
rect 9252 5408 9316 5412
rect 15012 5468 15076 5472
rect 15012 5412 15016 5468
rect 15016 5412 15072 5468
rect 15072 5412 15076 5468
rect 15012 5408 15076 5412
rect 15092 5468 15156 5472
rect 15092 5412 15096 5468
rect 15096 5412 15152 5468
rect 15152 5412 15156 5468
rect 15092 5408 15156 5412
rect 15172 5468 15236 5472
rect 15172 5412 15176 5468
rect 15176 5412 15232 5468
rect 15232 5412 15236 5468
rect 15172 5408 15236 5412
rect 15252 5468 15316 5472
rect 15252 5412 15256 5468
rect 15256 5412 15312 5468
rect 15312 5412 15316 5468
rect 15252 5408 15316 5412
rect 21012 5468 21076 5472
rect 21012 5412 21016 5468
rect 21016 5412 21072 5468
rect 21072 5412 21076 5468
rect 21012 5408 21076 5412
rect 21092 5468 21156 5472
rect 21092 5412 21096 5468
rect 21096 5412 21152 5468
rect 21152 5412 21156 5468
rect 21092 5408 21156 5412
rect 21172 5468 21236 5472
rect 21172 5412 21176 5468
rect 21176 5412 21232 5468
rect 21232 5412 21236 5468
rect 21172 5408 21236 5412
rect 21252 5468 21316 5472
rect 21252 5412 21256 5468
rect 21256 5412 21312 5468
rect 21312 5412 21316 5468
rect 21252 5408 21316 5412
rect 27012 5468 27076 5472
rect 27012 5412 27016 5468
rect 27016 5412 27072 5468
rect 27072 5412 27076 5468
rect 27012 5408 27076 5412
rect 27092 5468 27156 5472
rect 27092 5412 27096 5468
rect 27096 5412 27152 5468
rect 27152 5412 27156 5468
rect 27092 5408 27156 5412
rect 27172 5468 27236 5472
rect 27172 5412 27176 5468
rect 27176 5412 27232 5468
rect 27232 5412 27236 5468
rect 27172 5408 27236 5412
rect 27252 5468 27316 5472
rect 27252 5412 27256 5468
rect 27256 5412 27312 5468
rect 27312 5412 27316 5468
rect 27252 5408 27316 5412
rect 1952 4924 2016 4928
rect 1952 4868 1956 4924
rect 1956 4868 2012 4924
rect 2012 4868 2016 4924
rect 1952 4864 2016 4868
rect 2032 4924 2096 4928
rect 2032 4868 2036 4924
rect 2036 4868 2092 4924
rect 2092 4868 2096 4924
rect 2032 4864 2096 4868
rect 2112 4924 2176 4928
rect 2112 4868 2116 4924
rect 2116 4868 2172 4924
rect 2172 4868 2176 4924
rect 2112 4864 2176 4868
rect 2192 4924 2256 4928
rect 2192 4868 2196 4924
rect 2196 4868 2252 4924
rect 2252 4868 2256 4924
rect 2192 4864 2256 4868
rect 7952 4924 8016 4928
rect 7952 4868 7956 4924
rect 7956 4868 8012 4924
rect 8012 4868 8016 4924
rect 7952 4864 8016 4868
rect 8032 4924 8096 4928
rect 8032 4868 8036 4924
rect 8036 4868 8092 4924
rect 8092 4868 8096 4924
rect 8032 4864 8096 4868
rect 8112 4924 8176 4928
rect 8112 4868 8116 4924
rect 8116 4868 8172 4924
rect 8172 4868 8176 4924
rect 8112 4864 8176 4868
rect 8192 4924 8256 4928
rect 8192 4868 8196 4924
rect 8196 4868 8252 4924
rect 8252 4868 8256 4924
rect 8192 4864 8256 4868
rect 13952 4924 14016 4928
rect 13952 4868 13956 4924
rect 13956 4868 14012 4924
rect 14012 4868 14016 4924
rect 13952 4864 14016 4868
rect 14032 4924 14096 4928
rect 14032 4868 14036 4924
rect 14036 4868 14092 4924
rect 14092 4868 14096 4924
rect 14032 4864 14096 4868
rect 14112 4924 14176 4928
rect 14112 4868 14116 4924
rect 14116 4868 14172 4924
rect 14172 4868 14176 4924
rect 14112 4864 14176 4868
rect 14192 4924 14256 4928
rect 14192 4868 14196 4924
rect 14196 4868 14252 4924
rect 14252 4868 14256 4924
rect 14192 4864 14256 4868
rect 19952 4924 20016 4928
rect 19952 4868 19956 4924
rect 19956 4868 20012 4924
rect 20012 4868 20016 4924
rect 19952 4864 20016 4868
rect 20032 4924 20096 4928
rect 20032 4868 20036 4924
rect 20036 4868 20092 4924
rect 20092 4868 20096 4924
rect 20032 4864 20096 4868
rect 20112 4924 20176 4928
rect 20112 4868 20116 4924
rect 20116 4868 20172 4924
rect 20172 4868 20176 4924
rect 20112 4864 20176 4868
rect 20192 4924 20256 4928
rect 20192 4868 20196 4924
rect 20196 4868 20252 4924
rect 20252 4868 20256 4924
rect 20192 4864 20256 4868
rect 25952 4924 26016 4928
rect 25952 4868 25956 4924
rect 25956 4868 26012 4924
rect 26012 4868 26016 4924
rect 25952 4864 26016 4868
rect 26032 4924 26096 4928
rect 26032 4868 26036 4924
rect 26036 4868 26092 4924
rect 26092 4868 26096 4924
rect 26032 4864 26096 4868
rect 26112 4924 26176 4928
rect 26112 4868 26116 4924
rect 26116 4868 26172 4924
rect 26172 4868 26176 4924
rect 26112 4864 26176 4868
rect 26192 4924 26256 4928
rect 26192 4868 26196 4924
rect 26196 4868 26252 4924
rect 26252 4868 26256 4924
rect 26192 4864 26256 4868
rect 31952 4924 32016 4928
rect 31952 4868 31956 4924
rect 31956 4868 32012 4924
rect 32012 4868 32016 4924
rect 31952 4864 32016 4868
rect 32032 4924 32096 4928
rect 32032 4868 32036 4924
rect 32036 4868 32092 4924
rect 32092 4868 32096 4924
rect 32032 4864 32096 4868
rect 32112 4924 32176 4928
rect 32112 4868 32116 4924
rect 32116 4868 32172 4924
rect 32172 4868 32176 4924
rect 32112 4864 32176 4868
rect 32192 4924 32256 4928
rect 32192 4868 32196 4924
rect 32196 4868 32252 4924
rect 32252 4868 32256 4924
rect 32192 4864 32256 4868
rect 3012 4380 3076 4384
rect 3012 4324 3016 4380
rect 3016 4324 3072 4380
rect 3072 4324 3076 4380
rect 3012 4320 3076 4324
rect 3092 4380 3156 4384
rect 3092 4324 3096 4380
rect 3096 4324 3152 4380
rect 3152 4324 3156 4380
rect 3092 4320 3156 4324
rect 3172 4380 3236 4384
rect 3172 4324 3176 4380
rect 3176 4324 3232 4380
rect 3232 4324 3236 4380
rect 3172 4320 3236 4324
rect 3252 4380 3316 4384
rect 3252 4324 3256 4380
rect 3256 4324 3312 4380
rect 3312 4324 3316 4380
rect 3252 4320 3316 4324
rect 9012 4380 9076 4384
rect 9012 4324 9016 4380
rect 9016 4324 9072 4380
rect 9072 4324 9076 4380
rect 9012 4320 9076 4324
rect 9092 4380 9156 4384
rect 9092 4324 9096 4380
rect 9096 4324 9152 4380
rect 9152 4324 9156 4380
rect 9092 4320 9156 4324
rect 9172 4380 9236 4384
rect 9172 4324 9176 4380
rect 9176 4324 9232 4380
rect 9232 4324 9236 4380
rect 9172 4320 9236 4324
rect 9252 4380 9316 4384
rect 9252 4324 9256 4380
rect 9256 4324 9312 4380
rect 9312 4324 9316 4380
rect 9252 4320 9316 4324
rect 15012 4380 15076 4384
rect 15012 4324 15016 4380
rect 15016 4324 15072 4380
rect 15072 4324 15076 4380
rect 15012 4320 15076 4324
rect 15092 4380 15156 4384
rect 15092 4324 15096 4380
rect 15096 4324 15152 4380
rect 15152 4324 15156 4380
rect 15092 4320 15156 4324
rect 15172 4380 15236 4384
rect 15172 4324 15176 4380
rect 15176 4324 15232 4380
rect 15232 4324 15236 4380
rect 15172 4320 15236 4324
rect 15252 4380 15316 4384
rect 15252 4324 15256 4380
rect 15256 4324 15312 4380
rect 15312 4324 15316 4380
rect 15252 4320 15316 4324
rect 21012 4380 21076 4384
rect 21012 4324 21016 4380
rect 21016 4324 21072 4380
rect 21072 4324 21076 4380
rect 21012 4320 21076 4324
rect 21092 4380 21156 4384
rect 21092 4324 21096 4380
rect 21096 4324 21152 4380
rect 21152 4324 21156 4380
rect 21092 4320 21156 4324
rect 21172 4380 21236 4384
rect 21172 4324 21176 4380
rect 21176 4324 21232 4380
rect 21232 4324 21236 4380
rect 21172 4320 21236 4324
rect 21252 4380 21316 4384
rect 21252 4324 21256 4380
rect 21256 4324 21312 4380
rect 21312 4324 21316 4380
rect 21252 4320 21316 4324
rect 27012 4380 27076 4384
rect 27012 4324 27016 4380
rect 27016 4324 27072 4380
rect 27072 4324 27076 4380
rect 27012 4320 27076 4324
rect 27092 4380 27156 4384
rect 27092 4324 27096 4380
rect 27096 4324 27152 4380
rect 27152 4324 27156 4380
rect 27092 4320 27156 4324
rect 27172 4380 27236 4384
rect 27172 4324 27176 4380
rect 27176 4324 27232 4380
rect 27232 4324 27236 4380
rect 27172 4320 27236 4324
rect 27252 4380 27316 4384
rect 27252 4324 27256 4380
rect 27256 4324 27312 4380
rect 27312 4324 27316 4380
rect 27252 4320 27316 4324
rect 1952 3836 2016 3840
rect 1952 3780 1956 3836
rect 1956 3780 2012 3836
rect 2012 3780 2016 3836
rect 1952 3776 2016 3780
rect 2032 3836 2096 3840
rect 2032 3780 2036 3836
rect 2036 3780 2092 3836
rect 2092 3780 2096 3836
rect 2032 3776 2096 3780
rect 2112 3836 2176 3840
rect 2112 3780 2116 3836
rect 2116 3780 2172 3836
rect 2172 3780 2176 3836
rect 2112 3776 2176 3780
rect 2192 3836 2256 3840
rect 2192 3780 2196 3836
rect 2196 3780 2252 3836
rect 2252 3780 2256 3836
rect 2192 3776 2256 3780
rect 7952 3836 8016 3840
rect 7952 3780 7956 3836
rect 7956 3780 8012 3836
rect 8012 3780 8016 3836
rect 7952 3776 8016 3780
rect 8032 3836 8096 3840
rect 8032 3780 8036 3836
rect 8036 3780 8092 3836
rect 8092 3780 8096 3836
rect 8032 3776 8096 3780
rect 8112 3836 8176 3840
rect 8112 3780 8116 3836
rect 8116 3780 8172 3836
rect 8172 3780 8176 3836
rect 8112 3776 8176 3780
rect 8192 3836 8256 3840
rect 8192 3780 8196 3836
rect 8196 3780 8252 3836
rect 8252 3780 8256 3836
rect 8192 3776 8256 3780
rect 13952 3836 14016 3840
rect 13952 3780 13956 3836
rect 13956 3780 14012 3836
rect 14012 3780 14016 3836
rect 13952 3776 14016 3780
rect 14032 3836 14096 3840
rect 14032 3780 14036 3836
rect 14036 3780 14092 3836
rect 14092 3780 14096 3836
rect 14032 3776 14096 3780
rect 14112 3836 14176 3840
rect 14112 3780 14116 3836
rect 14116 3780 14172 3836
rect 14172 3780 14176 3836
rect 14112 3776 14176 3780
rect 14192 3836 14256 3840
rect 14192 3780 14196 3836
rect 14196 3780 14252 3836
rect 14252 3780 14256 3836
rect 14192 3776 14256 3780
rect 19952 3836 20016 3840
rect 19952 3780 19956 3836
rect 19956 3780 20012 3836
rect 20012 3780 20016 3836
rect 19952 3776 20016 3780
rect 20032 3836 20096 3840
rect 20032 3780 20036 3836
rect 20036 3780 20092 3836
rect 20092 3780 20096 3836
rect 20032 3776 20096 3780
rect 20112 3836 20176 3840
rect 20112 3780 20116 3836
rect 20116 3780 20172 3836
rect 20172 3780 20176 3836
rect 20112 3776 20176 3780
rect 20192 3836 20256 3840
rect 20192 3780 20196 3836
rect 20196 3780 20252 3836
rect 20252 3780 20256 3836
rect 20192 3776 20256 3780
rect 25952 3836 26016 3840
rect 25952 3780 25956 3836
rect 25956 3780 26012 3836
rect 26012 3780 26016 3836
rect 25952 3776 26016 3780
rect 26032 3836 26096 3840
rect 26032 3780 26036 3836
rect 26036 3780 26092 3836
rect 26092 3780 26096 3836
rect 26032 3776 26096 3780
rect 26112 3836 26176 3840
rect 26112 3780 26116 3836
rect 26116 3780 26172 3836
rect 26172 3780 26176 3836
rect 26112 3776 26176 3780
rect 26192 3836 26256 3840
rect 26192 3780 26196 3836
rect 26196 3780 26252 3836
rect 26252 3780 26256 3836
rect 26192 3776 26256 3780
rect 31952 3836 32016 3840
rect 31952 3780 31956 3836
rect 31956 3780 32012 3836
rect 32012 3780 32016 3836
rect 31952 3776 32016 3780
rect 32032 3836 32096 3840
rect 32032 3780 32036 3836
rect 32036 3780 32092 3836
rect 32092 3780 32096 3836
rect 32032 3776 32096 3780
rect 32112 3836 32176 3840
rect 32112 3780 32116 3836
rect 32116 3780 32172 3836
rect 32172 3780 32176 3836
rect 32112 3776 32176 3780
rect 32192 3836 32256 3840
rect 32192 3780 32196 3836
rect 32196 3780 32252 3836
rect 32252 3780 32256 3836
rect 32192 3776 32256 3780
rect 3012 3292 3076 3296
rect 3012 3236 3016 3292
rect 3016 3236 3072 3292
rect 3072 3236 3076 3292
rect 3012 3232 3076 3236
rect 3092 3292 3156 3296
rect 3092 3236 3096 3292
rect 3096 3236 3152 3292
rect 3152 3236 3156 3292
rect 3092 3232 3156 3236
rect 3172 3292 3236 3296
rect 3172 3236 3176 3292
rect 3176 3236 3232 3292
rect 3232 3236 3236 3292
rect 3172 3232 3236 3236
rect 3252 3292 3316 3296
rect 3252 3236 3256 3292
rect 3256 3236 3312 3292
rect 3312 3236 3316 3292
rect 3252 3232 3316 3236
rect 9012 3292 9076 3296
rect 9012 3236 9016 3292
rect 9016 3236 9072 3292
rect 9072 3236 9076 3292
rect 9012 3232 9076 3236
rect 9092 3292 9156 3296
rect 9092 3236 9096 3292
rect 9096 3236 9152 3292
rect 9152 3236 9156 3292
rect 9092 3232 9156 3236
rect 9172 3292 9236 3296
rect 9172 3236 9176 3292
rect 9176 3236 9232 3292
rect 9232 3236 9236 3292
rect 9172 3232 9236 3236
rect 9252 3292 9316 3296
rect 9252 3236 9256 3292
rect 9256 3236 9312 3292
rect 9312 3236 9316 3292
rect 9252 3232 9316 3236
rect 15012 3292 15076 3296
rect 15012 3236 15016 3292
rect 15016 3236 15072 3292
rect 15072 3236 15076 3292
rect 15012 3232 15076 3236
rect 15092 3292 15156 3296
rect 15092 3236 15096 3292
rect 15096 3236 15152 3292
rect 15152 3236 15156 3292
rect 15092 3232 15156 3236
rect 15172 3292 15236 3296
rect 15172 3236 15176 3292
rect 15176 3236 15232 3292
rect 15232 3236 15236 3292
rect 15172 3232 15236 3236
rect 15252 3292 15316 3296
rect 15252 3236 15256 3292
rect 15256 3236 15312 3292
rect 15312 3236 15316 3292
rect 15252 3232 15316 3236
rect 21012 3292 21076 3296
rect 21012 3236 21016 3292
rect 21016 3236 21072 3292
rect 21072 3236 21076 3292
rect 21012 3232 21076 3236
rect 21092 3292 21156 3296
rect 21092 3236 21096 3292
rect 21096 3236 21152 3292
rect 21152 3236 21156 3292
rect 21092 3232 21156 3236
rect 21172 3292 21236 3296
rect 21172 3236 21176 3292
rect 21176 3236 21232 3292
rect 21232 3236 21236 3292
rect 21172 3232 21236 3236
rect 21252 3292 21316 3296
rect 21252 3236 21256 3292
rect 21256 3236 21312 3292
rect 21312 3236 21316 3292
rect 21252 3232 21316 3236
rect 27012 3292 27076 3296
rect 27012 3236 27016 3292
rect 27016 3236 27072 3292
rect 27072 3236 27076 3292
rect 27012 3232 27076 3236
rect 27092 3292 27156 3296
rect 27092 3236 27096 3292
rect 27096 3236 27152 3292
rect 27152 3236 27156 3292
rect 27092 3232 27156 3236
rect 27172 3292 27236 3296
rect 27172 3236 27176 3292
rect 27176 3236 27232 3292
rect 27232 3236 27236 3292
rect 27172 3232 27236 3236
rect 27252 3292 27316 3296
rect 27252 3236 27256 3292
rect 27256 3236 27312 3292
rect 27312 3236 27316 3292
rect 27252 3232 27316 3236
rect 1952 2748 2016 2752
rect 1952 2692 1956 2748
rect 1956 2692 2012 2748
rect 2012 2692 2016 2748
rect 1952 2688 2016 2692
rect 2032 2748 2096 2752
rect 2032 2692 2036 2748
rect 2036 2692 2092 2748
rect 2092 2692 2096 2748
rect 2032 2688 2096 2692
rect 2112 2748 2176 2752
rect 2112 2692 2116 2748
rect 2116 2692 2172 2748
rect 2172 2692 2176 2748
rect 2112 2688 2176 2692
rect 2192 2748 2256 2752
rect 2192 2692 2196 2748
rect 2196 2692 2252 2748
rect 2252 2692 2256 2748
rect 2192 2688 2256 2692
rect 7952 2748 8016 2752
rect 7952 2692 7956 2748
rect 7956 2692 8012 2748
rect 8012 2692 8016 2748
rect 7952 2688 8016 2692
rect 8032 2748 8096 2752
rect 8032 2692 8036 2748
rect 8036 2692 8092 2748
rect 8092 2692 8096 2748
rect 8032 2688 8096 2692
rect 8112 2748 8176 2752
rect 8112 2692 8116 2748
rect 8116 2692 8172 2748
rect 8172 2692 8176 2748
rect 8112 2688 8176 2692
rect 8192 2748 8256 2752
rect 8192 2692 8196 2748
rect 8196 2692 8252 2748
rect 8252 2692 8256 2748
rect 8192 2688 8256 2692
rect 13952 2748 14016 2752
rect 13952 2692 13956 2748
rect 13956 2692 14012 2748
rect 14012 2692 14016 2748
rect 13952 2688 14016 2692
rect 14032 2748 14096 2752
rect 14032 2692 14036 2748
rect 14036 2692 14092 2748
rect 14092 2692 14096 2748
rect 14032 2688 14096 2692
rect 14112 2748 14176 2752
rect 14112 2692 14116 2748
rect 14116 2692 14172 2748
rect 14172 2692 14176 2748
rect 14112 2688 14176 2692
rect 14192 2748 14256 2752
rect 14192 2692 14196 2748
rect 14196 2692 14252 2748
rect 14252 2692 14256 2748
rect 14192 2688 14256 2692
rect 19952 2748 20016 2752
rect 19952 2692 19956 2748
rect 19956 2692 20012 2748
rect 20012 2692 20016 2748
rect 19952 2688 20016 2692
rect 20032 2748 20096 2752
rect 20032 2692 20036 2748
rect 20036 2692 20092 2748
rect 20092 2692 20096 2748
rect 20032 2688 20096 2692
rect 20112 2748 20176 2752
rect 20112 2692 20116 2748
rect 20116 2692 20172 2748
rect 20172 2692 20176 2748
rect 20112 2688 20176 2692
rect 20192 2748 20256 2752
rect 20192 2692 20196 2748
rect 20196 2692 20252 2748
rect 20252 2692 20256 2748
rect 20192 2688 20256 2692
rect 25952 2748 26016 2752
rect 25952 2692 25956 2748
rect 25956 2692 26012 2748
rect 26012 2692 26016 2748
rect 25952 2688 26016 2692
rect 26032 2748 26096 2752
rect 26032 2692 26036 2748
rect 26036 2692 26092 2748
rect 26092 2692 26096 2748
rect 26032 2688 26096 2692
rect 26112 2748 26176 2752
rect 26112 2692 26116 2748
rect 26116 2692 26172 2748
rect 26172 2692 26176 2748
rect 26112 2688 26176 2692
rect 26192 2748 26256 2752
rect 26192 2692 26196 2748
rect 26196 2692 26252 2748
rect 26252 2692 26256 2748
rect 26192 2688 26256 2692
rect 31952 2748 32016 2752
rect 31952 2692 31956 2748
rect 31956 2692 32012 2748
rect 32012 2692 32016 2748
rect 31952 2688 32016 2692
rect 32032 2748 32096 2752
rect 32032 2692 32036 2748
rect 32036 2692 32092 2748
rect 32092 2692 32096 2748
rect 32032 2688 32096 2692
rect 32112 2748 32176 2752
rect 32112 2692 32116 2748
rect 32116 2692 32172 2748
rect 32172 2692 32176 2748
rect 32112 2688 32176 2692
rect 32192 2748 32256 2752
rect 32192 2692 32196 2748
rect 32196 2692 32252 2748
rect 32252 2692 32256 2748
rect 32192 2688 32256 2692
rect 3012 2204 3076 2208
rect 3012 2148 3016 2204
rect 3016 2148 3072 2204
rect 3072 2148 3076 2204
rect 3012 2144 3076 2148
rect 3092 2204 3156 2208
rect 3092 2148 3096 2204
rect 3096 2148 3152 2204
rect 3152 2148 3156 2204
rect 3092 2144 3156 2148
rect 3172 2204 3236 2208
rect 3172 2148 3176 2204
rect 3176 2148 3232 2204
rect 3232 2148 3236 2204
rect 3172 2144 3236 2148
rect 3252 2204 3316 2208
rect 3252 2148 3256 2204
rect 3256 2148 3312 2204
rect 3312 2148 3316 2204
rect 3252 2144 3316 2148
rect 9012 2204 9076 2208
rect 9012 2148 9016 2204
rect 9016 2148 9072 2204
rect 9072 2148 9076 2204
rect 9012 2144 9076 2148
rect 9092 2204 9156 2208
rect 9092 2148 9096 2204
rect 9096 2148 9152 2204
rect 9152 2148 9156 2204
rect 9092 2144 9156 2148
rect 9172 2204 9236 2208
rect 9172 2148 9176 2204
rect 9176 2148 9232 2204
rect 9232 2148 9236 2204
rect 9172 2144 9236 2148
rect 9252 2204 9316 2208
rect 9252 2148 9256 2204
rect 9256 2148 9312 2204
rect 9312 2148 9316 2204
rect 9252 2144 9316 2148
rect 15012 2204 15076 2208
rect 15012 2148 15016 2204
rect 15016 2148 15072 2204
rect 15072 2148 15076 2204
rect 15012 2144 15076 2148
rect 15092 2204 15156 2208
rect 15092 2148 15096 2204
rect 15096 2148 15152 2204
rect 15152 2148 15156 2204
rect 15092 2144 15156 2148
rect 15172 2204 15236 2208
rect 15172 2148 15176 2204
rect 15176 2148 15232 2204
rect 15232 2148 15236 2204
rect 15172 2144 15236 2148
rect 15252 2204 15316 2208
rect 15252 2148 15256 2204
rect 15256 2148 15312 2204
rect 15312 2148 15316 2204
rect 15252 2144 15316 2148
rect 21012 2204 21076 2208
rect 21012 2148 21016 2204
rect 21016 2148 21072 2204
rect 21072 2148 21076 2204
rect 21012 2144 21076 2148
rect 21092 2204 21156 2208
rect 21092 2148 21096 2204
rect 21096 2148 21152 2204
rect 21152 2148 21156 2204
rect 21092 2144 21156 2148
rect 21172 2204 21236 2208
rect 21172 2148 21176 2204
rect 21176 2148 21232 2204
rect 21232 2148 21236 2204
rect 21172 2144 21236 2148
rect 21252 2204 21316 2208
rect 21252 2148 21256 2204
rect 21256 2148 21312 2204
rect 21312 2148 21316 2204
rect 21252 2144 21316 2148
rect 27012 2204 27076 2208
rect 27012 2148 27016 2204
rect 27016 2148 27072 2204
rect 27072 2148 27076 2204
rect 27012 2144 27076 2148
rect 27092 2204 27156 2208
rect 27092 2148 27096 2204
rect 27096 2148 27152 2204
rect 27152 2148 27156 2204
rect 27092 2144 27156 2148
rect 27172 2204 27236 2208
rect 27172 2148 27176 2204
rect 27176 2148 27232 2204
rect 27232 2148 27236 2204
rect 27172 2144 27236 2148
rect 27252 2204 27316 2208
rect 27252 2148 27256 2204
rect 27256 2148 27312 2204
rect 27312 2148 27316 2204
rect 27252 2144 27316 2148
<< metal4 >>
rect 1944 8192 2264 11250
rect 1944 8128 1952 8192
rect 2016 8128 2032 8192
rect 2096 8128 2112 8192
rect 2176 8128 2192 8192
rect 2256 8128 2264 8192
rect 1944 7104 2264 8128
rect 1944 7040 1952 7104
rect 2016 7040 2032 7104
rect 2096 7040 2112 7104
rect 2176 7040 2192 7104
rect 2256 7040 2264 7104
rect 1944 6016 2264 7040
rect 1944 5952 1952 6016
rect 2016 5952 2032 6016
rect 2096 5952 2112 6016
rect 2176 5952 2192 6016
rect 2256 5952 2264 6016
rect 1944 4928 2264 5952
rect 1944 4864 1952 4928
rect 2016 4864 2032 4928
rect 2096 4864 2112 4928
rect 2176 4864 2192 4928
rect 2256 4864 2264 4928
rect 1944 3840 2264 4864
rect 1944 3776 1952 3840
rect 2016 3776 2032 3840
rect 2096 3776 2112 3840
rect 2176 3776 2192 3840
rect 2256 3776 2264 3840
rect 1944 2752 2264 3776
rect 1944 2688 1952 2752
rect 2016 2688 2032 2752
rect 2096 2688 2112 2752
rect 2176 2688 2192 2752
rect 2256 2688 2264 2752
rect 1944 0 2264 2688
rect 3004 8736 3324 11250
rect 3004 8672 3012 8736
rect 3076 8672 3092 8736
rect 3156 8672 3172 8736
rect 3236 8672 3252 8736
rect 3316 8672 3324 8736
rect 3004 7648 3324 8672
rect 3004 7584 3012 7648
rect 3076 7584 3092 7648
rect 3156 7584 3172 7648
rect 3236 7584 3252 7648
rect 3316 7584 3324 7648
rect 3004 6560 3324 7584
rect 3004 6496 3012 6560
rect 3076 6496 3092 6560
rect 3156 6496 3172 6560
rect 3236 6496 3252 6560
rect 3316 6496 3324 6560
rect 3004 5472 3324 6496
rect 3004 5408 3012 5472
rect 3076 5408 3092 5472
rect 3156 5408 3172 5472
rect 3236 5408 3252 5472
rect 3316 5408 3324 5472
rect 3004 4384 3324 5408
rect 3004 4320 3012 4384
rect 3076 4320 3092 4384
rect 3156 4320 3172 4384
rect 3236 4320 3252 4384
rect 3316 4320 3324 4384
rect 3004 3296 3324 4320
rect 3004 3232 3012 3296
rect 3076 3232 3092 3296
rect 3156 3232 3172 3296
rect 3236 3232 3252 3296
rect 3316 3232 3324 3296
rect 3004 2208 3324 3232
rect 3004 2144 3012 2208
rect 3076 2144 3092 2208
rect 3156 2144 3172 2208
rect 3236 2144 3252 2208
rect 3316 2144 3324 2208
rect 3004 0 3324 2144
rect 7944 8192 8264 11250
rect 7944 8128 7952 8192
rect 8016 8128 8032 8192
rect 8096 8128 8112 8192
rect 8176 8128 8192 8192
rect 8256 8128 8264 8192
rect 7944 7104 8264 8128
rect 7944 7040 7952 7104
rect 8016 7040 8032 7104
rect 8096 7040 8112 7104
rect 8176 7040 8192 7104
rect 8256 7040 8264 7104
rect 7944 6016 8264 7040
rect 7944 5952 7952 6016
rect 8016 5952 8032 6016
rect 8096 5952 8112 6016
rect 8176 5952 8192 6016
rect 8256 5952 8264 6016
rect 7944 4928 8264 5952
rect 7944 4864 7952 4928
rect 8016 4864 8032 4928
rect 8096 4864 8112 4928
rect 8176 4864 8192 4928
rect 8256 4864 8264 4928
rect 7944 3840 8264 4864
rect 7944 3776 7952 3840
rect 8016 3776 8032 3840
rect 8096 3776 8112 3840
rect 8176 3776 8192 3840
rect 8256 3776 8264 3840
rect 7944 2752 8264 3776
rect 7944 2688 7952 2752
rect 8016 2688 8032 2752
rect 8096 2688 8112 2752
rect 8176 2688 8192 2752
rect 8256 2688 8264 2752
rect 7944 0 8264 2688
rect 9004 8736 9324 11250
rect 9004 8672 9012 8736
rect 9076 8672 9092 8736
rect 9156 8672 9172 8736
rect 9236 8672 9252 8736
rect 9316 8672 9324 8736
rect 9004 7648 9324 8672
rect 9004 7584 9012 7648
rect 9076 7584 9092 7648
rect 9156 7584 9172 7648
rect 9236 7584 9252 7648
rect 9316 7584 9324 7648
rect 9004 6560 9324 7584
rect 9004 6496 9012 6560
rect 9076 6496 9092 6560
rect 9156 6496 9172 6560
rect 9236 6496 9252 6560
rect 9316 6496 9324 6560
rect 9004 5472 9324 6496
rect 9004 5408 9012 5472
rect 9076 5408 9092 5472
rect 9156 5408 9172 5472
rect 9236 5408 9252 5472
rect 9316 5408 9324 5472
rect 9004 4384 9324 5408
rect 9004 4320 9012 4384
rect 9076 4320 9092 4384
rect 9156 4320 9172 4384
rect 9236 4320 9252 4384
rect 9316 4320 9324 4384
rect 9004 3296 9324 4320
rect 9004 3232 9012 3296
rect 9076 3232 9092 3296
rect 9156 3232 9172 3296
rect 9236 3232 9252 3296
rect 9316 3232 9324 3296
rect 9004 2208 9324 3232
rect 9004 2144 9012 2208
rect 9076 2144 9092 2208
rect 9156 2144 9172 2208
rect 9236 2144 9252 2208
rect 9316 2144 9324 2208
rect 9004 0 9324 2144
rect 13944 8192 14264 11250
rect 13944 8128 13952 8192
rect 14016 8128 14032 8192
rect 14096 8128 14112 8192
rect 14176 8128 14192 8192
rect 14256 8128 14264 8192
rect 13944 7104 14264 8128
rect 13944 7040 13952 7104
rect 14016 7040 14032 7104
rect 14096 7040 14112 7104
rect 14176 7040 14192 7104
rect 14256 7040 14264 7104
rect 13944 6016 14264 7040
rect 13944 5952 13952 6016
rect 14016 5952 14032 6016
rect 14096 5952 14112 6016
rect 14176 5952 14192 6016
rect 14256 5952 14264 6016
rect 13944 4928 14264 5952
rect 13944 4864 13952 4928
rect 14016 4864 14032 4928
rect 14096 4864 14112 4928
rect 14176 4864 14192 4928
rect 14256 4864 14264 4928
rect 13944 3840 14264 4864
rect 13944 3776 13952 3840
rect 14016 3776 14032 3840
rect 14096 3776 14112 3840
rect 14176 3776 14192 3840
rect 14256 3776 14264 3840
rect 13944 2752 14264 3776
rect 13944 2688 13952 2752
rect 14016 2688 14032 2752
rect 14096 2688 14112 2752
rect 14176 2688 14192 2752
rect 14256 2688 14264 2752
rect 13944 0 14264 2688
rect 15004 8736 15324 11250
rect 15004 8672 15012 8736
rect 15076 8672 15092 8736
rect 15156 8672 15172 8736
rect 15236 8672 15252 8736
rect 15316 8672 15324 8736
rect 15004 7648 15324 8672
rect 15004 7584 15012 7648
rect 15076 7584 15092 7648
rect 15156 7584 15172 7648
rect 15236 7584 15252 7648
rect 15316 7584 15324 7648
rect 15004 6560 15324 7584
rect 15004 6496 15012 6560
rect 15076 6496 15092 6560
rect 15156 6496 15172 6560
rect 15236 6496 15252 6560
rect 15316 6496 15324 6560
rect 15004 5472 15324 6496
rect 15004 5408 15012 5472
rect 15076 5408 15092 5472
rect 15156 5408 15172 5472
rect 15236 5408 15252 5472
rect 15316 5408 15324 5472
rect 15004 4384 15324 5408
rect 15004 4320 15012 4384
rect 15076 4320 15092 4384
rect 15156 4320 15172 4384
rect 15236 4320 15252 4384
rect 15316 4320 15324 4384
rect 15004 3296 15324 4320
rect 15004 3232 15012 3296
rect 15076 3232 15092 3296
rect 15156 3232 15172 3296
rect 15236 3232 15252 3296
rect 15316 3232 15324 3296
rect 15004 2208 15324 3232
rect 15004 2144 15012 2208
rect 15076 2144 15092 2208
rect 15156 2144 15172 2208
rect 15236 2144 15252 2208
rect 15316 2144 15324 2208
rect 15004 0 15324 2144
rect 19944 8192 20264 11250
rect 19944 8128 19952 8192
rect 20016 8128 20032 8192
rect 20096 8128 20112 8192
rect 20176 8128 20192 8192
rect 20256 8128 20264 8192
rect 19944 7104 20264 8128
rect 19944 7040 19952 7104
rect 20016 7040 20032 7104
rect 20096 7040 20112 7104
rect 20176 7040 20192 7104
rect 20256 7040 20264 7104
rect 19944 6016 20264 7040
rect 19944 5952 19952 6016
rect 20016 5952 20032 6016
rect 20096 5952 20112 6016
rect 20176 5952 20192 6016
rect 20256 5952 20264 6016
rect 19944 4928 20264 5952
rect 19944 4864 19952 4928
rect 20016 4864 20032 4928
rect 20096 4864 20112 4928
rect 20176 4864 20192 4928
rect 20256 4864 20264 4928
rect 19944 3840 20264 4864
rect 19944 3776 19952 3840
rect 20016 3776 20032 3840
rect 20096 3776 20112 3840
rect 20176 3776 20192 3840
rect 20256 3776 20264 3840
rect 19944 2752 20264 3776
rect 19944 2688 19952 2752
rect 20016 2688 20032 2752
rect 20096 2688 20112 2752
rect 20176 2688 20192 2752
rect 20256 2688 20264 2752
rect 19944 0 20264 2688
rect 21004 8736 21324 11250
rect 21004 8672 21012 8736
rect 21076 8672 21092 8736
rect 21156 8672 21172 8736
rect 21236 8672 21252 8736
rect 21316 8672 21324 8736
rect 21004 7648 21324 8672
rect 21004 7584 21012 7648
rect 21076 7584 21092 7648
rect 21156 7584 21172 7648
rect 21236 7584 21252 7648
rect 21316 7584 21324 7648
rect 21004 6560 21324 7584
rect 21004 6496 21012 6560
rect 21076 6496 21092 6560
rect 21156 6496 21172 6560
rect 21236 6496 21252 6560
rect 21316 6496 21324 6560
rect 21004 5472 21324 6496
rect 21004 5408 21012 5472
rect 21076 5408 21092 5472
rect 21156 5408 21172 5472
rect 21236 5408 21252 5472
rect 21316 5408 21324 5472
rect 21004 4384 21324 5408
rect 21004 4320 21012 4384
rect 21076 4320 21092 4384
rect 21156 4320 21172 4384
rect 21236 4320 21252 4384
rect 21316 4320 21324 4384
rect 21004 3296 21324 4320
rect 21004 3232 21012 3296
rect 21076 3232 21092 3296
rect 21156 3232 21172 3296
rect 21236 3232 21252 3296
rect 21316 3232 21324 3296
rect 21004 2208 21324 3232
rect 21004 2144 21012 2208
rect 21076 2144 21092 2208
rect 21156 2144 21172 2208
rect 21236 2144 21252 2208
rect 21316 2144 21324 2208
rect 21004 0 21324 2144
rect 25944 8192 26264 11250
rect 25944 8128 25952 8192
rect 26016 8128 26032 8192
rect 26096 8128 26112 8192
rect 26176 8128 26192 8192
rect 26256 8128 26264 8192
rect 25944 7104 26264 8128
rect 25944 7040 25952 7104
rect 26016 7040 26032 7104
rect 26096 7040 26112 7104
rect 26176 7040 26192 7104
rect 26256 7040 26264 7104
rect 25944 6016 26264 7040
rect 25944 5952 25952 6016
rect 26016 5952 26032 6016
rect 26096 5952 26112 6016
rect 26176 5952 26192 6016
rect 26256 5952 26264 6016
rect 25944 4928 26264 5952
rect 25944 4864 25952 4928
rect 26016 4864 26032 4928
rect 26096 4864 26112 4928
rect 26176 4864 26192 4928
rect 26256 4864 26264 4928
rect 25944 3840 26264 4864
rect 25944 3776 25952 3840
rect 26016 3776 26032 3840
rect 26096 3776 26112 3840
rect 26176 3776 26192 3840
rect 26256 3776 26264 3840
rect 25944 2752 26264 3776
rect 25944 2688 25952 2752
rect 26016 2688 26032 2752
rect 26096 2688 26112 2752
rect 26176 2688 26192 2752
rect 26256 2688 26264 2752
rect 25944 0 26264 2688
rect 27004 8736 27324 11250
rect 27004 8672 27012 8736
rect 27076 8672 27092 8736
rect 27156 8672 27172 8736
rect 27236 8672 27252 8736
rect 27316 8672 27324 8736
rect 27004 7648 27324 8672
rect 27004 7584 27012 7648
rect 27076 7584 27092 7648
rect 27156 7584 27172 7648
rect 27236 7584 27252 7648
rect 27316 7584 27324 7648
rect 27004 6560 27324 7584
rect 27004 6496 27012 6560
rect 27076 6496 27092 6560
rect 27156 6496 27172 6560
rect 27236 6496 27252 6560
rect 27316 6496 27324 6560
rect 27004 5472 27324 6496
rect 27004 5408 27012 5472
rect 27076 5408 27092 5472
rect 27156 5408 27172 5472
rect 27236 5408 27252 5472
rect 27316 5408 27324 5472
rect 27004 4384 27324 5408
rect 27004 4320 27012 4384
rect 27076 4320 27092 4384
rect 27156 4320 27172 4384
rect 27236 4320 27252 4384
rect 27316 4320 27324 4384
rect 27004 3296 27324 4320
rect 27004 3232 27012 3296
rect 27076 3232 27092 3296
rect 27156 3232 27172 3296
rect 27236 3232 27252 3296
rect 27316 3232 27324 3296
rect 27004 2208 27324 3232
rect 27004 2144 27012 2208
rect 27076 2144 27092 2208
rect 27156 2144 27172 2208
rect 27236 2144 27252 2208
rect 27316 2144 27324 2208
rect 27004 0 27324 2144
rect 31944 8192 32264 11250
rect 31944 8128 31952 8192
rect 32016 8128 32032 8192
rect 32096 8128 32112 8192
rect 32176 8128 32192 8192
rect 32256 8128 32264 8192
rect 31944 7104 32264 8128
rect 31944 7040 31952 7104
rect 32016 7040 32032 7104
rect 32096 7040 32112 7104
rect 32176 7040 32192 7104
rect 32256 7040 32264 7104
rect 31944 6016 32264 7040
rect 31944 5952 31952 6016
rect 32016 5952 32032 6016
rect 32096 5952 32112 6016
rect 32176 5952 32192 6016
rect 32256 5952 32264 6016
rect 31944 4928 32264 5952
rect 31944 4864 31952 4928
rect 32016 4864 32032 4928
rect 32096 4864 32112 4928
rect 32176 4864 32192 4928
rect 32256 4864 32264 4928
rect 31944 3840 32264 4864
rect 31944 3776 31952 3840
rect 32016 3776 32032 3840
rect 32096 3776 32112 3840
rect 32176 3776 32192 3840
rect 32256 3776 32264 3840
rect 31944 2752 32264 3776
rect 31944 2688 31952 2752
rect 32016 2688 32032 2752
rect 32096 2688 32112 2752
rect 32176 2688 32192 2752
rect 32256 2688 32264 2752
rect 31944 0 32264 2688
use sky130_fd_sc_hd__buf_1  _00_
timestamp -3599
transform 1 0 4692 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _01_
timestamp -3599
transform 1 0 11316 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _02_
timestamp -3599
transform 1 0 11960 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _03_
timestamp -3599
transform 1 0 12236 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _04_
timestamp -3599
transform 1 0 8188 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _05_
timestamp -3599
transform 1 0 18308 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _06_
timestamp -3599
transform 1 0 17020 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _07_
timestamp -3599
transform 1 0 17296 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _08_
timestamp -3599
transform 1 0 18584 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _09_
timestamp -3599
transform 1 0 10396 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _10_
timestamp -3599
transform 1 0 19504 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _11_
timestamp -3599
transform 1 0 19228 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _12_
timestamp -3599
transform 1 0 18860 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _13_
timestamp -3599
transform 1 0 15456 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _14_
timestamp -3599
transform 1 0 6716 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _15_
timestamp -3599
transform -1 0 10948 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _16_
timestamp -3599
transform 1 0 15732 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _17_
timestamp -3599
transform 1 0 20884 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _18_
timestamp -3599
transform 1 0 12512 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _19_
timestamp -3599
transform 1 0 19504 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _20_
timestamp -3599
transform 1 0 16376 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _21_
timestamp -3599
transform 1 0 15088 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _22_
timestamp -3599
transform -1 0 26404 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _23_
timestamp -3599
transform 1 0 16652 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _24_
timestamp -3599
transform -1 0 24932 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _25_
timestamp -3599
transform -1 0 23552 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _26_
timestamp -3599
transform -1 0 26588 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _27_
timestamp -3599
transform 1 0 21160 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _28_
timestamp -3599
transform 1 0 21436 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _29_
timestamp -3599
transform 1 0 16376 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _30_
timestamp -3599
transform 1 0 19320 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _31_
timestamp -3599
transform -1 0 27876 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _32_
timestamp -3599
transform -1 0 22448 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _33_
timestamp -3599
transform 1 0 14536 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _34_
timestamp -3599
transform -1 0 18032 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _35_
timestamp -3599
transform 1 0 9384 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _36_
timestamp -3599
transform -1 0 22724 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _37_
timestamp -3599
transform -1 0 25852 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _38_
timestamp -3599
transform -1 0 26220 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _39_
timestamp -3599
transform -1 0 25576 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _40_
timestamp -3599
transform -1 0 24012 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _41_
timestamp -3599
transform -1 0 22908 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _42_
timestamp -3599
transform -1 0 21528 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _43_
timestamp -3599
transform -1 0 21712 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _44_
timestamp -3599
transform -1 0 22356 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _45_
timestamp -3599
transform -1 0 22264 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _46_
timestamp -3599
transform -1 0 23644 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _47_
timestamp -3599
transform -1 0 23920 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _48_
timestamp -3599
transform -1 0 24656 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _49_
timestamp -3599
transform -1 0 26680 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _50_
timestamp -3599
transform -1 0 28796 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _51_
timestamp -3599
transform 1 0 30820 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _52_
timestamp -3599
transform 1 0 6256 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _53_
timestamp -3599
transform 1 0 7820 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _54_
timestamp -3599
transform 1 0 7912 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _55_
timestamp -3599
transform 1 0 9476 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _56_
timestamp -3599
transform -1 0 4508 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _57_
timestamp -3599
transform 1 0 5244 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _58_
timestamp -3599
transform 1 0 6624 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _59_
timestamp -3599
transform 1 0 7636 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _60_
timestamp -3599
transform 1 0 8924 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _61_
timestamp -3599
transform 1 0 10028 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _62_
timestamp -3599
transform 1 0 11040 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _63_
timestamp -3599
transform 1 0 8464 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _64_
timestamp -3599
transform -1 0 6808 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _65_
timestamp -3599
transform -1 0 7452 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _66_
timestamp -3599
transform 1 0 7636 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _67_
timestamp -3599
transform 1 0 8648 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _68_
timestamp -3599
transform 1 0 9200 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _69_
timestamp -3599
transform 1 0 10304 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _70_
timestamp -3599
transform 1 0 9936 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _71_
timestamp -3599
transform 1 0 10672 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _72_
timestamp -3599
transform -1 0 20976 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _73_
timestamp -3599
transform 1 0 19780 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _74_
timestamp -3599
transform 1 0 18216 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _75_
timestamp -3599
transform 1 0 17480 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _76_
timestamp -3599
transform 1 0 17112 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _77_
timestamp -3599
transform 1 0 15548 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _78_
timestamp -3599
transform 1 0 14352 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _79_
timestamp -3599
transform 1 0 13432 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _80_
timestamp -3599
transform 1 0 12604 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _81_
timestamp -3599
transform -1 0 11592 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _82_
timestamp -3599
transform -1 0 10028 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _83_
timestamp -3599
transform -1 0 8464 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _84_
timestamp -3599
transform -1 0 11868 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _85_
timestamp -3599
transform -1 0 11316 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _86_
timestamp -3599
transform -1 0 10948 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _87_
timestamp -3599
transform -1 0 10488 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _88_
timestamp -3599
transform 1 0 21804 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1
timestamp -3599
transform -1 0 19964 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_2
timestamp -3599
transform -1 0 20148 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_3
timestamp -3599
transform 1 0 18124 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_4
timestamp -3599
transform 1 0 14996 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_5
timestamp -3599
transform -1 0 12512 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_6
timestamp -3599
transform -1 0 11316 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_7
timestamp -3599
transform 1 0 16192 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_8
timestamp -3599
transform 1 0 25944 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_9
timestamp -3599
transform -1 0 17112 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_10
timestamp -3599
transform -1 0 24656 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_11
timestamp -3599
transform -1 0 23276 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_12
timestamp -3599
transform -1 0 26312 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_13
timestamp -3599
transform 1 0 20976 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_14
timestamp -3599
transform -1 0 21896 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_15
timestamp -3599
transform 1 0 16192 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_16
timestamp -3599
transform -1 0 11960 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_17
timestamp -3599
transform -1 0 19780 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_18
timestamp -3599
transform -1 0 27600 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_19
timestamp -3599
transform -1 0 12696 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_20
timestamp -3599
transform -1 0 17756 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_21
timestamp -3599
transform -1 0 17020 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_22
timestamp -3599
transform -1 0 16836 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_23
timestamp -3599
transform -1 0 20332 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_24
timestamp -3599
transform 1 0 10212 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_25
timestamp -3599
transform -1 0 16652 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_26
timestamp -3599
transform -1 0 9200 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_27
timestamp -3599
transform -1 0 8648 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_28
timestamp -3599
transform -1 0 10672 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_29
timestamp -3599
transform 1 0 15272 0 1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3
timestamp 1636964856
transform 1 0 1380 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15
timestamp 1636964856
transform 1 0 2484 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27
timestamp -3599
transform 1 0 3588 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29
timestamp 1636964856
transform 1 0 3772 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41
timestamp 1636964856
transform 1 0 4876 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_53
timestamp -3599
transform 1 0 5980 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57
timestamp 1636964856
transform 1 0 6348 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69
timestamp 1636964856
transform 1 0 7452 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_81
timestamp -3599
transform 1 0 8556 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85
timestamp 1636964856
transform 1 0 8924 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_97
timestamp 1636964856
transform 1 0 10028 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_109
timestamp -3599
transform 1 0 11132 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_113
timestamp 1636964856
transform 1 0 11500 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_125
timestamp 1636964856
transform 1 0 12604 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_137
timestamp -3599
transform 1 0 13708 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_141
timestamp 1636964856
transform 1 0 14076 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_153
timestamp 1636964856
transform 1 0 15180 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_165
timestamp -3599
transform 1 0 16284 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_169
timestamp 1636964856
transform 1 0 16652 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_181
timestamp 1636964856
transform 1 0 17756 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_193
timestamp -3599
transform 1 0 18860 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_197
timestamp 1636964856
transform 1 0 19228 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_209
timestamp 1636964856
transform 1 0 20332 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_221
timestamp -3599
transform 1 0 21436 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_225
timestamp 1636964856
transform 1 0 21804 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_237
timestamp 1636964856
transform 1 0 22908 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_249
timestamp -3599
transform 1 0 24012 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_253
timestamp 1636964856
transform 1 0 24380 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_265
timestamp 1636964856
transform 1 0 25484 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_277
timestamp -3599
transform 1 0 26588 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_281
timestamp 1636964856
transform 1 0 26956 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_293
timestamp 1636964856
transform 1 0 28060 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_305
timestamp -3599
transform 1 0 29164 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_309
timestamp -3599
transform 1 0 29532 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_317
timestamp -3599
transform 1 0 30268 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_337
timestamp -3599
transform 1 0 32108 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_1_3
timestamp 1636964856
transform 1 0 1380 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_15
timestamp 1636964856
transform 1 0 2484 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_27
timestamp 1636964856
transform 1 0 3588 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_39
timestamp 1636964856
transform 1 0 4692 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_51
timestamp -3599
transform 1 0 5796 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_55
timestamp -3599
transform 1 0 6164 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_57
timestamp 1636964856
transform 1 0 6348 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_69
timestamp 1636964856
transform 1 0 7452 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_81
timestamp 1636964856
transform 1 0 8556 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_93
timestamp 1636964856
transform 1 0 9660 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_105
timestamp -3599
transform 1 0 10764 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_111
timestamp -3599
transform 1 0 11316 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_113
timestamp 1636964856
transform 1 0 11500 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_125
timestamp 1636964856
transform 1 0 12604 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_137
timestamp 1636964856
transform 1 0 13708 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_149
timestamp 1636964856
transform 1 0 14812 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_161
timestamp -3599
transform 1 0 15916 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_167
timestamp -3599
transform 1 0 16468 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_169
timestamp 1636964856
transform 1 0 16652 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_181
timestamp 1636964856
transform 1 0 17756 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_193
timestamp 1636964856
transform 1 0 18860 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_205
timestamp 1636964856
transform 1 0 19964 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_217
timestamp -3599
transform 1 0 21068 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_223
timestamp -3599
transform 1 0 21620 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_225
timestamp 1636964856
transform 1 0 21804 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_237
timestamp 1636964856
transform 1 0 22908 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_249
timestamp 1636964856
transform 1 0 24012 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_261
timestamp 1636964856
transform 1 0 25116 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_273
timestamp -3599
transform 1 0 26220 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_279
timestamp -3599
transform 1 0 26772 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_281
timestamp 1636964856
transform 1 0 26956 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_293
timestamp 1636964856
transform 1 0 28060 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_305
timestamp 1636964856
transform 1 0 29164 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_317
timestamp -3599
transform 1 0 30268 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_1_325
timestamp -3599
transform 1 0 31004 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_1_337
timestamp -3599
transform 1 0 32108 0 -1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3
timestamp 1636964856
transform 1 0 1380 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_15
timestamp 1636964856
transform 1 0 2484 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_2_27
timestamp -3599
transform 1 0 3588 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_2_29
timestamp -3599
transform 1 0 3772 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_2_37
timestamp -3599
transform 1 0 4508 0 1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_2_42
timestamp 1636964856
transform 1 0 4968 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_54
timestamp -3599
transform 1 0 6072 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_60
timestamp -3599
transform 1 0 6624 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_64
timestamp 1636964856
transform 1 0 6992 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_2_76
timestamp -3599
transform 1 0 8096 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_80
timestamp -3599
transform 1 0 8464 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_85
timestamp -3599
transform 1 0 8924 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_89
timestamp -3599
transform 1 0 9292 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_2_93
timestamp -3599
transform 1 0 9660 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_2_107
timestamp -3599
transform 1 0 10948 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_114
timestamp -3599
transform 1 0 11592 0 1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_2_126
timestamp 1636964856
transform 1 0 12696 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_2_138
timestamp -3599
transform 1 0 13800 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_141
timestamp -3599
transform 1 0 14076 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_145
timestamp -3599
transform 1 0 14444 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_149
timestamp -3599
transform 1 0 14812 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_2_153
timestamp -3599
transform 1 0 15180 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_162
timestamp -3599
transform 1 0 16008 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_166
timestamp -3599
transform 1 0 16376 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_2_184
timestamp -3599
transform 1 0 18032 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_209
timestamp 1636964856
transform 1 0 20332 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_2_221
timestamp -3599
transform 1 0 21436 0 1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_2_235
timestamp 1636964856
transform 1 0 22724 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_2_247
timestamp -3599
transform 1 0 23828 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_251
timestamp -3599
transform 1 0 24196 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_2_253
timestamp -3599
transform 1 0 24380 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_2_261
timestamp -3599
transform 1 0 25116 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_2_269
timestamp -3599
transform 1 0 25852 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_273
timestamp 1636964856
transform 1 0 26220 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_285
timestamp 1636964856
transform 1 0 27324 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_2_297
timestamp -3599
transform 1 0 28428 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_2_305
timestamp -3599
transform 1 0 29164 0 1 3264
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_2_309
timestamp 1636964856
transform 1 0 29532 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_2_321
timestamp -3599
transform 1 0 30636 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_2_329
timestamp -3599
transform 1 0 31372 0 1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3
timestamp 1636964856
transform 1 0 1380 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_15
timestamp 1636964856
transform 1 0 2484 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_27
timestamp 1636964856
transform 1 0 3588 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_39
timestamp 1636964856
transform 1 0 4692 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_3_51
timestamp -3599
transform 1 0 5796 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_55
timestamp -3599
transform 1 0 6164 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_57
timestamp 1636964856
transform 1 0 6348 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_69
timestamp 1636964856
transform 1 0 7452 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_81
timestamp 1636964856
transform 1 0 8556 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_93
timestamp 1636964856
transform 1 0 9660 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_105
timestamp -3599
transform 1 0 10764 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_111
timestamp -3599
transform 1 0 11316 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_3_113
timestamp -3599
transform 1 0 11500 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_3_121
timestamp -3599
transform 1 0 12236 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_127
timestamp 1636964856
transform 1 0 12788 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_139
timestamp 1636964856
transform 1 0 13892 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_151
timestamp 1636964856
transform 1 0 14996 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_3_163
timestamp -3599
transform 1 0 16100 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_167
timestamp -3599
transform 1 0 16468 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_169
timestamp 1636964856
transform 1 0 16652 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_181
timestamp 1636964856
transform 1 0 17756 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_193
timestamp 1636964856
transform 1 0 18860 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_3_205
timestamp -3599
transform 1 0 19964 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_3_213
timestamp -3599
transform 1 0 20700 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_3_218
timestamp -3599
transform 1 0 21160 0 -1 4352
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_3_225
timestamp 1636964856
transform 1 0 21804 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_237
timestamp 1636964856
transform 1 0 22908 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_249
timestamp 1636964856
transform 1 0 24012 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_261
timestamp 1636964856
transform 1 0 25116 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_273
timestamp -3599
transform 1 0 26220 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_279
timestamp -3599
transform 1 0 26772 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_281
timestamp 1636964856
transform 1 0 26956 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_293
timestamp 1636964856
transform 1 0 28060 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_305
timestamp 1636964856
transform 1 0 29164 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_3_317
timestamp -3599
transform 1 0 30268 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_3_325
timestamp -3599
transform 1 0 31004 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_3_337
timestamp -3599
transform 1 0 32108 0 -1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3
timestamp 1636964856
transform 1 0 1380 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_15
timestamp 1636964856
transform 1 0 2484 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_4_27
timestamp -3599
transform 1 0 3588 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_29
timestamp 1636964856
transform 1 0 3772 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_41
timestamp 1636964856
transform 1 0 4876 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_53
timestamp 1636964856
transform 1 0 5980 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_65
timestamp 1636964856
transform 1 0 7084 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_77
timestamp -3599
transform 1 0 8188 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_83
timestamp -3599
transform 1 0 8740 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_85
timestamp 1636964856
transform 1 0 8924 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_97
timestamp 1636964856
transform 1 0 10028 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_109
timestamp 1636964856
transform 1 0 11132 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_121
timestamp 1636964856
transform 1 0 12236 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_133
timestamp -3599
transform 1 0 13340 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_139
timestamp -3599
transform 1 0 13892 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_141
timestamp 1636964856
transform 1 0 14076 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_153
timestamp 1636964856
transform 1 0 15180 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_165
timestamp 1636964856
transform 1 0 16284 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_177
timestamp 1636964856
transform 1 0 17388 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_189
timestamp -3599
transform 1 0 18492 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_195
timestamp -3599
transform 1 0 19044 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_4_197
timestamp -3599
transform 1 0 19228 0 1 4352
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_4_203
timestamp 1636964856
transform 1 0 19780 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_215
timestamp 1636964856
transform 1 0 20884 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_227
timestamp -3599
transform 1 0 21988 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_233
timestamp -3599
transform 1 0 22540 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_4_237
timestamp -3599
transform 1 0 22908 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_4_245
timestamp -3599
transform 1 0 23644 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_4_249
timestamp -3599
transform 1 0 24012 0 1 4352
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_4_253
timestamp 1636964856
transform 1 0 24380 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_265
timestamp 1636964856
transform 1 0 25484 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_277
timestamp 1636964856
transform 1 0 26588 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_289
timestamp 1636964856
transform 1 0 27692 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_301
timestamp -3599
transform 1 0 28796 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_307
timestamp -3599
transform 1 0 29348 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_309
timestamp 1636964856
transform 1 0 29532 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_4_321
timestamp -3599
transform 1 0 30636 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_4_329
timestamp -3599
transform 1 0 31372 0 1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3
timestamp 1636964856
transform 1 0 1380 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_15
timestamp 1636964856
transform 1 0 2484 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_27
timestamp 1636964856
transform 1 0 3588 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_39
timestamp 1636964856
transform 1 0 4692 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_5_51
timestamp -3599
transform 1 0 5796 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_55
timestamp -3599
transform 1 0 6164 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_57
timestamp 1636964856
transform 1 0 6348 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_5_69
timestamp -3599
transform 1 0 7452 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_5_77
timestamp -3599
transform 1 0 8188 0 -1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_5_83
timestamp 1636964856
transform 1 0 8740 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_95
timestamp 1636964856
transform 1 0 9844 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_5_107
timestamp -3599
transform 1 0 10948 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_111
timestamp -3599
transform 1 0 11316 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_113
timestamp 1636964856
transform 1 0 11500 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_125
timestamp 1636964856
transform 1 0 12604 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_137
timestamp 1636964856
transform 1 0 13708 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_5_149
timestamp -3599
transform 1 0 14812 0 -1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_5_155
timestamp 1636964856
transform 1 0 15364 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_5_167
timestamp -3599
transform 1 0 16468 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_169
timestamp 1636964856
transform 1 0 16652 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_181
timestamp 1636964856
transform 1 0 17756 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_193
timestamp 1636964856
transform 1 0 18860 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_205
timestamp 1636964856
transform 1 0 19964 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_5_217
timestamp -3599
transform 1 0 21068 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_222
timestamp -3599
transform 1 0 21528 0 -1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_5_225
timestamp 1636964856
transform 1 0 21804 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_237
timestamp 1636964856
transform 1 0 22908 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_249
timestamp 1636964856
transform 1 0 24012 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_261
timestamp 1636964856
transform 1 0 25116 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_273
timestamp -3599
transform 1 0 26220 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_279
timestamp -3599
transform 1 0 26772 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_281
timestamp 1636964856
transform 1 0 26956 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_293
timestamp 1636964856
transform 1 0 28060 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_305
timestamp 1636964856
transform 1 0 29164 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_5_317
timestamp -3599
transform 1 0 30268 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_5_325
timestamp -3599
transform 1 0 31004 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_5_337
timestamp -3599
transform 1 0 32108 0 -1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3
timestamp 1636964856
transform 1 0 1380 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_15
timestamp 1636964856
transform 1 0 2484 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_6_27
timestamp -3599
transform 1 0 3588 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_29
timestamp 1636964856
transform 1 0 3772 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_41
timestamp 1636964856
transform 1 0 4876 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_53
timestamp -3599
transform 1 0 5980 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_6_62
timestamp -3599
transform 1 0 6808 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_6_69
timestamp -3599
transform 1 0 7452 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_6_74
timestamp -3599
transform 1 0 7912 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_6_82
timestamp -3599
transform 1 0 8648 0 1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_6_88
timestamp 1636964856
transform 1 0 9200 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_100
timestamp 1636964856
transform 1 0 10304 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_112
timestamp 1636964856
transform 1 0 11408 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_124
timestamp 1636964856
transform 1 0 12512 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_6_136
timestamp -3599
transform 1 0 13616 0 1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_6_141
timestamp 1636964856
transform 1 0 14076 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_6_153
timestamp -3599
transform 1 0 15180 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_6_161
timestamp -3599
transform 1 0 15916 0 1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_6_169
timestamp 1636964856
transform 1 0 16652 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_181
timestamp 1636964856
transform 1 0 17756 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_6_193
timestamp -3599
transform 1 0 18860 0 1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_6_197
timestamp 1636964856
transform 1 0 19228 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_209
timestamp 1636964856
transform 1 0 20332 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_224
timestamp 1636964856
transform 1 0 21712 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_236
timestamp 1636964856
transform 1 0 22816 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_6_248
timestamp -3599
transform 1 0 23920 0 1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_6_253
timestamp 1636964856
transform 1 0 24380 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_265
timestamp 1636964856
transform 1 0 25484 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_277
timestamp 1636964856
transform 1 0 26588 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_289
timestamp 1636964856
transform 1 0 27692 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_301
timestamp -3599
transform 1 0 28796 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_307
timestamp -3599
transform 1 0 29348 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_309
timestamp 1636964856
transform 1 0 29532 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_321
timestamp -3599
transform 1 0 30636 0 1 5440
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3
timestamp 1636964856
transform 1 0 1380 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_15
timestamp 1636964856
transform 1 0 2484 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_27
timestamp 1636964856
transform 1 0 3588 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_39
timestamp -3599
transform 1 0 4692 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_7_48
timestamp -3599
transform 1 0 5520 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_7_57
timestamp -3599
transform 1 0 6348 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_7_63
timestamp -3599
transform 1 0 6900 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_7_85
timestamp -3599
transform 1 0 8924 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_7_103
timestamp -3599
transform 1 0 10580 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_7_107
timestamp -3599
transform 1 0 10948 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_7_111
timestamp -3599
transform 1 0 11316 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_113
timestamp 1636964856
transform 1 0 11500 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_125
timestamp 1636964856
transform 1 0 12604 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_137
timestamp 1636964856
transform 1 0 13708 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_149
timestamp 1636964856
transform 1 0 14812 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_161
timestamp -3599
transform 1 0 15916 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_167
timestamp -3599
transform 1 0 16468 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_169
timestamp 1636964856
transform 1 0 16652 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_181
timestamp 1636964856
transform 1 0 17756 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_193
timestamp 1636964856
transform 1 0 18860 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_205
timestamp 1636964856
transform 1 0 19964 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_217
timestamp -3599
transform 1 0 21068 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_223
timestamp -3599
transform 1 0 21620 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_7_225
timestamp -3599
transform 1 0 21804 0 -1 6528
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_7_231
timestamp 1636964856
transform 1 0 22356 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_243
timestamp 1636964856
transform 1 0 23460 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_255
timestamp 1636964856
transform 1 0 24564 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_267
timestamp 1636964856
transform 1 0 25668 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_7_279
timestamp -3599
transform 1 0 26772 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_281
timestamp 1636964856
transform 1 0 26956 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_293
timestamp -3599
transform 1 0 28060 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_297
timestamp -3599
transform 1 0 28428 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_301
timestamp 1636964856
transform 1 0 28796 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_7_313
timestamp -3599
transform 1 0 29900 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_7_321
timestamp -3599
transform 1 0 30636 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_326
timestamp -3599
transform 1 0 31096 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_337
timestamp -3599
transform 1 0 32108 0 -1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3
timestamp 1636964856
transform 1 0 1380 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_15
timestamp 1636964856
transform 1 0 2484 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_8_27
timestamp -3599
transform 1 0 3588 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_29
timestamp -3599
transform 1 0 3772 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_33
timestamp -3599
transform 1 0 4140 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_37
timestamp 1636964856
transform 1 0 4508 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_49
timestamp -3599
transform 1 0 5612 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_55
timestamp -3599
transform 1 0 6164 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_59
timestamp 1636964856
transform 1 0 6532 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_8_71
timestamp -3599
transform 1 0 7636 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_8_76
timestamp -3599
transform 1 0 8096 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_8_85
timestamp -3599
transform 1 0 8924 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_8_93
timestamp -3599
transform 1 0 9660 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_8_107
timestamp -3599
transform 1 0 10948 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_8_117
timestamp -3599
transform 1 0 11868 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_8_128
timestamp -3599
transform 1 0 12880 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_8_137
timestamp -3599
transform 1 0 13708 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_141
timestamp -3599
transform 1 0 14076 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_8_147
timestamp -3599
transform 1 0 14628 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_8_155
timestamp -3599
transform 1 0 15364 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_160
timestamp -3599
transform 1 0 15824 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_177
timestamp -3599
transform 1 0 17388 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_181
timestamp -3599
transform 1 0 17756 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_185
timestamp -3599
transform 1 0 18124 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_8_189
timestamp -3599
transform 1 0 18492 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_195
timestamp -3599
transform 1 0 19044 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_8_197
timestamp -3599
transform 1 0 19228 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_8_206
timestamp -3599
transform 1 0 20056 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_212
timestamp -3599
transform 1 0 20608 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_226
timestamp 1636964856
transform 1 0 21896 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_8_238
timestamp -3599
transform 1 0 23000 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_248
timestamp -3599
transform 1 0 23920 0 1 6528
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_8_256
timestamp 1636964856
transform 1 0 24656 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_8_268
timestamp -3599
transform 1 0 25760 0 1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_8_278
timestamp 1636964856
transform 1 0 26680 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_290
timestamp 1636964856
transform 1 0 27784 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_302
timestamp -3599
transform 1 0 28888 0 1 6528
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_8_309
timestamp 1636964856
transform 1 0 29532 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_321
timestamp -3599
transform 1 0 30636 0 1 6528
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3
timestamp 1636964856
transform 1 0 1380 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_15
timestamp 1636964856
transform 1 0 2484 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_27
timestamp 1636964856
transform 1 0 3588 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_39
timestamp 1636964856
transform 1 0 4692 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_9_51
timestamp -3599
transform 1 0 5796 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_55
timestamp -3599
transform 1 0 6164 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_57
timestamp 1636964856
transform 1 0 6348 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_69
timestamp 1636964856
transform 1 0 7452 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_81
timestamp 1636964856
transform 1 0 8556 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_93
timestamp 1636964856
transform 1 0 9660 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_105
timestamp -3599
transform 1 0 10764 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_111
timestamp -3599
transform 1 0 11316 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_113
timestamp 1636964856
transform 1 0 11500 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_125
timestamp 1636964856
transform 1 0 12604 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_137
timestamp 1636964856
transform 1 0 13708 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_149
timestamp 1636964856
transform 1 0 14812 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_161
timestamp -3599
transform 1 0 15916 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_167
timestamp -3599
transform 1 0 16468 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_169
timestamp 1636964856
transform 1 0 16652 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_181
timestamp 1636964856
transform 1 0 17756 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_193
timestamp 1636964856
transform 1 0 18860 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_205
timestamp 1636964856
transform 1 0 19964 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_217
timestamp -3599
transform 1 0 21068 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_223
timestamp -3599
transform 1 0 21620 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_225
timestamp -3599
transform 1 0 21804 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_9_230
timestamp -3599
transform 1 0 22264 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_9_238
timestamp -3599
transform 1 0 23000 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_9_244
timestamp -3599
transform 1 0 23552 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_9_252
timestamp -3599
transform 1 0 24288 0 -1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_9_259
timestamp 1636964856
transform 1 0 24932 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_9_271
timestamp -3599
transform 1 0 26036 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_9_277
timestamp -3599
transform 1 0 26588 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_9_281
timestamp -3599
transform 1 0 26956 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_285
timestamp -3599
transform 1 0 27324 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_291
timestamp 1636964856
transform 1 0 27876 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_303
timestamp 1636964856
transform 1 0 28980 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_315
timestamp 1636964856
transform 1 0 30084 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_9_327
timestamp -3599
transform 1 0 31188 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_337
timestamp -3599
transform 1 0 32108 0 -1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_10_3
timestamp 1636964856
transform 1 0 1380 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_15
timestamp 1636964856
transform 1 0 2484 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_10_27
timestamp -3599
transform 1 0 3588 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_29
timestamp -3599
transform 1 0 3772 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_33
timestamp -3599
transform 1 0 4140 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_10_38
timestamp -3599
transform 1 0 4600 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_10_50
timestamp -3599
transform 1 0 5704 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_54
timestamp -3599
transform 1 0 6072 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_59
timestamp -3599
transform 1 0 6532 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_65
timestamp -3599
transform 1 0 7084 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_69
timestamp -3599
transform 1 0 7452 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_74
timestamp -3599
transform 1 0 7912 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_78
timestamp -3599
transform 1 0 8280 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_10_83
timestamp -3599
transform 1 0 8740 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_10_85
timestamp -3599
transform 1 0 8924 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_10_92
timestamp -3599
transform 1 0 9568 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_10_98
timestamp -3599
transform 1 0 10120 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_10_110
timestamp -3599
transform 1 0 11224 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_116
timestamp -3599
transform 1 0 11776 0 1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_10_122
timestamp 1636964856
transform 1 0 12328 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_134
timestamp -3599
transform 1 0 13432 0 1 7616
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_10_141
timestamp 1636964856
transform 1 0 14076 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_153
timestamp 1636964856
transform 1 0 15180 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_165
timestamp 1636964856
transform 1 0 16284 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_177
timestamp 1636964856
transform 1 0 17388 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_189
timestamp -3599
transform 1 0 18492 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_195
timestamp -3599
transform 1 0 19044 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_197
timestamp 1636964856
transform 1 0 19228 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_209
timestamp 1636964856
transform 1 0 20332 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_221
timestamp 1636964856
transform 1 0 21436 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_233
timestamp 1636964856
transform 1 0 22540 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_245
timestamp -3599
transform 1 0 23644 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_251
timestamp -3599
transform 1 0 24196 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_253
timestamp 1636964856
transform 1 0 24380 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_265
timestamp -3599
transform 1 0 25484 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_10_275
timestamp -3599
transform 1 0 26404 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_10_287
timestamp -3599
transform 1 0 27508 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_10_303
timestamp -3599
transform 1 0 28980 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_307
timestamp -3599
transform 1 0 29348 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_10_313
timestamp -3599
transform 1 0 29900 0 1 7616
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_11_3
timestamp 1636964856
transform 1 0 1380 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_15
timestamp 1636964856
transform 1 0 2484 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_11_27
timestamp -3599
transform 1 0 3588 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_11_29
timestamp -3599
transform 1 0 3772 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_57
timestamp -3599
transform 1 0 6348 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_85
timestamp -3599
transform 1 0 8924 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_113
timestamp -3599
transform 1 0 11500 0 -1 8704
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_11_145
timestamp 1636964856
transform 1 0 14444 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_11_157
timestamp -3599
transform 1 0 15548 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_11_165
timestamp -3599
transform 1 0 16284 0 -1 8704
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_11_169
timestamp 1636964856
transform 1 0 16652 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_181
timestamp 1636964856
transform 1 0 17756 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_11_193
timestamp -3599
transform 1 0 18860 0 -1 8704
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_11_197
timestamp 1636964856
transform 1 0 19228 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_209
timestamp 1636964856
transform 1 0 20332 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_11_221
timestamp -3599
transform 1 0 21436 0 -1 8704
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_11_225
timestamp 1636964856
transform 1 0 21804 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_237
timestamp 1636964856
transform 1 0 22908 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_11_277
timestamp -3599
transform 1 0 26588 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_305
timestamp -3599
transform 1 0 29164 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_321
timestamp -3599
transform 1 0 30636 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_11_337
timestamp -3599
transform 1 0 32108 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  output1
timestamp -3599
transform 1 0 31280 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output2
timestamp -3599
transform 1 0 31556 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output3
timestamp -3599
transform 1 0 31924 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output4
timestamp -3599
transform 1 0 31280 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output5
timestamp -3599
transform 1 0 31648 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output6
timestamp -3599
transform 1 0 31188 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output7
timestamp -3599
transform 1 0 31556 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output8
timestamp -3599
transform 1 0 31924 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output9
timestamp -3599
transform 1 0 31280 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output10
timestamp -3599
transform 1 0 31648 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output11
timestamp -3599
transform 1 0 31188 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output12
timestamp -3599
transform 1 0 30912 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output13
timestamp -3599
transform 1 0 31556 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output14
timestamp -3599
transform 1 0 31648 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output15
timestamp -3599
transform 1 0 31556 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output16
timestamp -3599
transform 1 0 31924 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output17
timestamp -3599
transform 1 0 31648 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output18
timestamp -3599
transform 1 0 31280 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output19
timestamp -3599
transform 1 0 30912 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output20
timestamp -3599
transform 1 0 31188 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output21
timestamp -3599
transform 1 0 30820 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output22
timestamp -3599
transform 1 0 31280 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output23
timestamp -3599
transform 1 0 30544 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output24
timestamp -3599
transform 1 0 30452 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output25
timestamp -3599
transform 1 0 31924 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output26
timestamp -3599
transform 1 0 31648 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output27
timestamp -3599
transform 1 0 31280 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output28
timestamp -3599
transform 1 0 31648 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output29
timestamp -3599
transform 1 0 31556 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output30
timestamp -3599
transform 1 0 31924 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output31
timestamp -3599
transform 1 0 31280 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output32
timestamp -3599
transform 1 0 31648 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output33
timestamp -3599
transform 1 0 24380 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output34
timestamp -3599
transform 1 0 27140 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output35
timestamp -3599
transform 1 0 28060 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output36
timestamp -3599
transform 1 0 28428 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output37
timestamp -3599
transform 1 0 28796 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output38
timestamp -3599
transform 1 0 28244 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output39
timestamp -3599
transform 1 0 28612 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output40
timestamp -3599
transform 1 0 29532 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output41
timestamp -3599
transform 1 0 29900 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output42
timestamp -3599
transform 1 0 29532 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output43
timestamp -3599
transform -1 0 30636 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output44
timestamp -3599
transform 1 0 24748 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output45
timestamp -3599
transform 1 0 25116 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output46
timestamp -3599
transform 1 0 25484 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output47
timestamp -3599
transform 1 0 25852 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output48
timestamp -3599
transform 1 0 26220 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output49
timestamp -3599
transform -1 0 26404 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output50
timestamp -3599
transform 1 0 26956 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output51
timestamp -3599
transform 1 0 27324 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output52
timestamp -3599
transform 1 0 27692 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output53
timestamp -3599
transform -1 0 4600 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output54
timestamp -3599
transform -1 0 4416 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output55
timestamp -3599
transform -1 0 4784 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output56
timestamp -3599
transform -1 0 5152 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output57
timestamp -3599
transform 1 0 5336 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output58
timestamp -3599
transform 1 0 5152 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output59
timestamp -3599
transform -1 0 5888 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output60
timestamp -3599
transform -1 0 6532 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output61
timestamp -3599
transform -1 0 6256 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output62
timestamp -3599
transform -1 0 7084 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output63
timestamp -3599
transform -1 0 6992 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output64
timestamp -3599
transform -1 0 7360 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output65
timestamp -3599
transform 1 0 7544 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output66
timestamp -3599
transform 1 0 7360 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output67
timestamp -3599
transform 1 0 7728 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output68
timestamp -3599
transform -1 0 8740 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output69
timestamp -3599
transform -1 0 8464 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output70
timestamp -3599
transform -1 0 8832 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output71
timestamp -3599
transform -1 0 9568 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output72
timestamp -3599
transform -1 0 9568 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output73
timestamp -3599
transform -1 0 10120 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output74
timestamp -3599
transform 1 0 12144 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output75
timestamp -3599
transform 1 0 12512 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output76
timestamp -3599
transform 1 0 12880 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output77
timestamp -3599
transform 1 0 13248 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output78
timestamp -3599
transform 1 0 13616 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output79
timestamp -3599
transform 1 0 14076 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output80
timestamp -3599
transform -1 0 9936 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output81
timestamp -3599
transform -1 0 10304 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output82
timestamp -3599
transform -1 0 10672 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output83
timestamp -3599
transform -1 0 11224 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output84
timestamp -3599
transform -1 0 11040 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output85
timestamp -3599
transform -1 0 11776 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output86
timestamp -3599
transform -1 0 11408 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output87
timestamp -3599
transform -1 0 12328 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output88
timestamp -3599
transform 1 0 11776 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  output89
timestamp -3599
transform -1 0 24288 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Left_12
timestamp -3599
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Right_0
timestamp -3599
transform -1 0 32568 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Left_13
timestamp -3599
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Right_1
timestamp -3599
transform -1 0 32568 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Left_14
timestamp -3599
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Right_2
timestamp -3599
transform -1 0 32568 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Left_15
timestamp -3599
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Right_3
timestamp -3599
transform -1 0 32568 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Left_16
timestamp -3599
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Right_4
timestamp -3599
transform -1 0 32568 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Left_17
timestamp -3599
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Right_5
timestamp -3599
transform -1 0 32568 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Left_18
timestamp -3599
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Right_6
timestamp -3599
transform -1 0 32568 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Left_19
timestamp -3599
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Right_7
timestamp -3599
transform -1 0 32568 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Left_20
timestamp -3599
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Right_8
timestamp -3599
transform -1 0 32568 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Left_21
timestamp -3599
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Right_9
timestamp -3599
transform -1 0 32568 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_Left_22
timestamp -3599
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_Right_10
timestamp -3599
transform -1 0 32568 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_Left_23
timestamp -3599
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_Right_11
timestamp -3599
transform -1 0 32568 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_24
timestamp -3599
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_25
timestamp -3599
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_26
timestamp -3599
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_27
timestamp -3599
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_28
timestamp -3599
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_29
timestamp -3599
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_30
timestamp -3599
transform 1 0 19136 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_31
timestamp -3599
transform 1 0 21712 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_32
timestamp -3599
transform 1 0 24288 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_33
timestamp -3599
transform 1 0 26864 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_34
timestamp -3599
transform 1 0 29440 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_35
timestamp -3599
transform 1 0 32016 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_36
timestamp -3599
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_37
timestamp -3599
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_38
timestamp -3599
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_39
timestamp -3599
transform 1 0 21712 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_40
timestamp -3599
transform 1 0 26864 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_41
timestamp -3599
transform 1 0 32016 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_42
timestamp -3599
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_43
timestamp -3599
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_44
timestamp -3599
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_45
timestamp -3599
transform 1 0 19136 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_46
timestamp -3599
transform 1 0 24288 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_47
timestamp -3599
transform 1 0 29440 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_48
timestamp -3599
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_49
timestamp -3599
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_50
timestamp -3599
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_51
timestamp -3599
transform 1 0 21712 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_52
timestamp -3599
transform 1 0 26864 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_53
timestamp -3599
transform 1 0 32016 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_54
timestamp -3599
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_55
timestamp -3599
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_56
timestamp -3599
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_57
timestamp -3599
transform 1 0 19136 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_58
timestamp -3599
transform 1 0 24288 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_59
timestamp -3599
transform 1 0 29440 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_60
timestamp -3599
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_61
timestamp -3599
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_62
timestamp -3599
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_63
timestamp -3599
transform 1 0 21712 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_64
timestamp -3599
transform 1 0 26864 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_65
timestamp -3599
transform 1 0 32016 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_66
timestamp -3599
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_67
timestamp -3599
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_68
timestamp -3599
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_69
timestamp -3599
transform 1 0 19136 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_70
timestamp -3599
transform 1 0 24288 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_71
timestamp -3599
transform 1 0 29440 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_72
timestamp -3599
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_73
timestamp -3599
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_74
timestamp -3599
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_75
timestamp -3599
transform 1 0 21712 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_76
timestamp -3599
transform 1 0 26864 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_77
timestamp -3599
transform 1 0 32016 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_78
timestamp -3599
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_79
timestamp -3599
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_80
timestamp -3599
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_81
timestamp -3599
transform 1 0 19136 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_82
timestamp -3599
transform 1 0 24288 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_83
timestamp -3599
transform 1 0 29440 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_84
timestamp -3599
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_85
timestamp -3599
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_86
timestamp -3599
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_87
timestamp -3599
transform 1 0 21712 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_88
timestamp -3599
transform 1 0 26864 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_89
timestamp -3599
transform 1 0 32016 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_90
timestamp -3599
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_91
timestamp -3599
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_92
timestamp -3599
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_93
timestamp -3599
transform 1 0 19136 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_94
timestamp -3599
transform 1 0 24288 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_95
timestamp -3599
transform 1 0 29440 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_96
timestamp -3599
transform 1 0 3680 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_97
timestamp -3599
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_98
timestamp -3599
transform 1 0 8832 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_99
timestamp -3599
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_100
timestamp -3599
transform 1 0 13984 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_101
timestamp -3599
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_102
timestamp -3599
transform 1 0 19136 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_103
timestamp -3599
transform 1 0 21712 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_104
timestamp -3599
transform 1 0 24288 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_105
timestamp -3599
transform 1 0 26864 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_106
timestamp -3599
transform 1 0 29440 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_107
timestamp -3599
transform 1 0 32016 0 -1 8704
box -38 -48 130 592
<< labels >>
flabel metal3 s 0 1368 120 1488 0 FreeSans 480 0 0 0 FrameData[0]
port 0 nsew signal input
flabel metal3 s 0 4088 120 4208 0 FreeSans 480 0 0 0 FrameData[10]
port 1 nsew signal input
flabel metal3 s 0 4360 120 4480 0 FreeSans 480 0 0 0 FrameData[11]
port 2 nsew signal input
flabel metal3 s 0 4632 120 4752 0 FreeSans 480 0 0 0 FrameData[12]
port 3 nsew signal input
flabel metal3 s 0 4904 120 5024 0 FreeSans 480 0 0 0 FrameData[13]
port 4 nsew signal input
flabel metal3 s 0 5176 120 5296 0 FreeSans 480 0 0 0 FrameData[14]
port 5 nsew signal input
flabel metal3 s 0 5448 120 5568 0 FreeSans 480 0 0 0 FrameData[15]
port 6 nsew signal input
flabel metal3 s 0 5720 120 5840 0 FreeSans 480 0 0 0 FrameData[16]
port 7 nsew signal input
flabel metal3 s 0 5992 120 6112 0 FreeSans 480 0 0 0 FrameData[17]
port 8 nsew signal input
flabel metal3 s 0 6264 120 6384 0 FreeSans 480 0 0 0 FrameData[18]
port 9 nsew signal input
flabel metal3 s 0 6536 120 6656 0 FreeSans 480 0 0 0 FrameData[19]
port 10 nsew signal input
flabel metal3 s 0 1640 120 1760 0 FreeSans 480 0 0 0 FrameData[1]
port 11 nsew signal input
flabel metal3 s 0 6808 120 6928 0 FreeSans 480 0 0 0 FrameData[20]
port 12 nsew signal input
flabel metal3 s 0 7080 120 7200 0 FreeSans 480 0 0 0 FrameData[21]
port 13 nsew signal input
flabel metal3 s 0 7352 120 7472 0 FreeSans 480 0 0 0 FrameData[22]
port 14 nsew signal input
flabel metal3 s 0 7624 120 7744 0 FreeSans 480 0 0 0 FrameData[23]
port 15 nsew signal input
flabel metal3 s 0 7896 120 8016 0 FreeSans 480 0 0 0 FrameData[24]
port 16 nsew signal input
flabel metal3 s 0 8168 120 8288 0 FreeSans 480 0 0 0 FrameData[25]
port 17 nsew signal input
flabel metal3 s 0 8440 120 8560 0 FreeSans 480 0 0 0 FrameData[26]
port 18 nsew signal input
flabel metal3 s 0 8712 120 8832 0 FreeSans 480 0 0 0 FrameData[27]
port 19 nsew signal input
flabel metal3 s 0 8984 120 9104 0 FreeSans 480 0 0 0 FrameData[28]
port 20 nsew signal input
flabel metal3 s 0 9256 120 9376 0 FreeSans 480 0 0 0 FrameData[29]
port 21 nsew signal input
flabel metal3 s 0 1912 120 2032 0 FreeSans 480 0 0 0 FrameData[2]
port 22 nsew signal input
flabel metal3 s 0 9528 120 9648 0 FreeSans 480 0 0 0 FrameData[30]
port 23 nsew signal input
flabel metal3 s 0 9800 120 9920 0 FreeSans 480 0 0 0 FrameData[31]
port 24 nsew signal input
flabel metal3 s 0 2184 120 2304 0 FreeSans 480 0 0 0 FrameData[3]
port 25 nsew signal input
flabel metal3 s 0 2456 120 2576 0 FreeSans 480 0 0 0 FrameData[4]
port 26 nsew signal input
flabel metal3 s 0 2728 120 2848 0 FreeSans 480 0 0 0 FrameData[5]
port 27 nsew signal input
flabel metal3 s 0 3000 120 3120 0 FreeSans 480 0 0 0 FrameData[6]
port 28 nsew signal input
flabel metal3 s 0 3272 120 3392 0 FreeSans 480 0 0 0 FrameData[7]
port 29 nsew signal input
flabel metal3 s 0 3544 120 3664 0 FreeSans 480 0 0 0 FrameData[8]
port 30 nsew signal input
flabel metal3 s 0 3816 120 3936 0 FreeSans 480 0 0 0 FrameData[9]
port 31 nsew signal input
flabel metal3 s 33630 1368 33750 1488 0 FreeSans 480 0 0 0 FrameData_O[0]
port 32 nsew signal output
flabel metal3 s 33630 4088 33750 4208 0 FreeSans 480 0 0 0 FrameData_O[10]
port 33 nsew signal output
flabel metal3 s 33630 4360 33750 4480 0 FreeSans 480 0 0 0 FrameData_O[11]
port 34 nsew signal output
flabel metal3 s 33630 4632 33750 4752 0 FreeSans 480 0 0 0 FrameData_O[12]
port 35 nsew signal output
flabel metal3 s 33630 4904 33750 5024 0 FreeSans 480 0 0 0 FrameData_O[13]
port 36 nsew signal output
flabel metal3 s 33630 5176 33750 5296 0 FreeSans 480 0 0 0 FrameData_O[14]
port 37 nsew signal output
flabel metal3 s 33630 5448 33750 5568 0 FreeSans 480 0 0 0 FrameData_O[15]
port 38 nsew signal output
flabel metal3 s 33630 5720 33750 5840 0 FreeSans 480 0 0 0 FrameData_O[16]
port 39 nsew signal output
flabel metal3 s 33630 5992 33750 6112 0 FreeSans 480 0 0 0 FrameData_O[17]
port 40 nsew signal output
flabel metal3 s 33630 6264 33750 6384 0 FreeSans 480 0 0 0 FrameData_O[18]
port 41 nsew signal output
flabel metal3 s 33630 6536 33750 6656 0 FreeSans 480 0 0 0 FrameData_O[19]
port 42 nsew signal output
flabel metal3 s 33630 1640 33750 1760 0 FreeSans 480 0 0 0 FrameData_O[1]
port 43 nsew signal output
flabel metal3 s 33630 6808 33750 6928 0 FreeSans 480 0 0 0 FrameData_O[20]
port 44 nsew signal output
flabel metal3 s 33630 7080 33750 7200 0 FreeSans 480 0 0 0 FrameData_O[21]
port 45 nsew signal output
flabel metal3 s 33630 7352 33750 7472 0 FreeSans 480 0 0 0 FrameData_O[22]
port 46 nsew signal output
flabel metal3 s 33630 7624 33750 7744 0 FreeSans 480 0 0 0 FrameData_O[23]
port 47 nsew signal output
flabel metal3 s 33630 7896 33750 8016 0 FreeSans 480 0 0 0 FrameData_O[24]
port 48 nsew signal output
flabel metal3 s 33630 8168 33750 8288 0 FreeSans 480 0 0 0 FrameData_O[25]
port 49 nsew signal output
flabel metal3 s 33630 8440 33750 8560 0 FreeSans 480 0 0 0 FrameData_O[26]
port 50 nsew signal output
flabel metal3 s 33630 8712 33750 8832 0 FreeSans 480 0 0 0 FrameData_O[27]
port 51 nsew signal output
flabel metal3 s 33630 8984 33750 9104 0 FreeSans 480 0 0 0 FrameData_O[28]
port 52 nsew signal output
flabel metal3 s 33630 9256 33750 9376 0 FreeSans 480 0 0 0 FrameData_O[29]
port 53 nsew signal output
flabel metal3 s 33630 1912 33750 2032 0 FreeSans 480 0 0 0 FrameData_O[2]
port 54 nsew signal output
flabel metal3 s 33630 9528 33750 9648 0 FreeSans 480 0 0 0 FrameData_O[30]
port 55 nsew signal output
flabel metal3 s 33630 9800 33750 9920 0 FreeSans 480 0 0 0 FrameData_O[31]
port 56 nsew signal output
flabel metal3 s 33630 2184 33750 2304 0 FreeSans 480 0 0 0 FrameData_O[3]
port 57 nsew signal output
flabel metal3 s 33630 2456 33750 2576 0 FreeSans 480 0 0 0 FrameData_O[4]
port 58 nsew signal output
flabel metal3 s 33630 2728 33750 2848 0 FreeSans 480 0 0 0 FrameData_O[5]
port 59 nsew signal output
flabel metal3 s 33630 3000 33750 3120 0 FreeSans 480 0 0 0 FrameData_O[6]
port 60 nsew signal output
flabel metal3 s 33630 3272 33750 3392 0 FreeSans 480 0 0 0 FrameData_O[7]
port 61 nsew signal output
flabel metal3 s 33630 3544 33750 3664 0 FreeSans 480 0 0 0 FrameData_O[8]
port 62 nsew signal output
flabel metal3 s 33630 3816 33750 3936 0 FreeSans 480 0 0 0 FrameData_O[9]
port 63 nsew signal output
flabel metal2 s 2778 0 2834 56 0 FreeSans 224 0 0 0 FrameStrobe[0]
port 64 nsew signal input
flabel metal2 s 18418 0 18474 56 0 FreeSans 224 0 0 0 FrameStrobe[10]
port 65 nsew signal input
flabel metal2 s 19982 0 20038 56 0 FreeSans 224 0 0 0 FrameStrobe[11]
port 66 nsew signal input
flabel metal2 s 21546 0 21602 56 0 FreeSans 224 0 0 0 FrameStrobe[12]
port 67 nsew signal input
flabel metal2 s 23110 0 23166 56 0 FreeSans 224 0 0 0 FrameStrobe[13]
port 68 nsew signal input
flabel metal2 s 24674 0 24730 56 0 FreeSans 224 0 0 0 FrameStrobe[14]
port 69 nsew signal input
flabel metal2 s 26238 0 26294 56 0 FreeSans 224 0 0 0 FrameStrobe[15]
port 70 nsew signal input
flabel metal2 s 27802 0 27858 56 0 FreeSans 224 0 0 0 FrameStrobe[16]
port 71 nsew signal input
flabel metal2 s 29366 0 29422 56 0 FreeSans 224 0 0 0 FrameStrobe[17]
port 72 nsew signal input
flabel metal2 s 30930 0 30986 56 0 FreeSans 224 0 0 0 FrameStrobe[18]
port 73 nsew signal input
flabel metal2 s 32494 0 32550 56 0 FreeSans 224 0 0 0 FrameStrobe[19]
port 74 nsew signal input
flabel metal2 s 4342 0 4398 56 0 FreeSans 224 0 0 0 FrameStrobe[1]
port 75 nsew signal input
flabel metal2 s 5906 0 5962 56 0 FreeSans 224 0 0 0 FrameStrobe[2]
port 76 nsew signal input
flabel metal2 s 7470 0 7526 56 0 FreeSans 224 0 0 0 FrameStrobe[3]
port 77 nsew signal input
flabel metal2 s 9034 0 9090 56 0 FreeSans 224 0 0 0 FrameStrobe[4]
port 78 nsew signal input
flabel metal2 s 10598 0 10654 56 0 FreeSans 224 0 0 0 FrameStrobe[5]
port 79 nsew signal input
flabel metal2 s 12162 0 12218 56 0 FreeSans 224 0 0 0 FrameStrobe[6]
port 80 nsew signal input
flabel metal2 s 13726 0 13782 56 0 FreeSans 224 0 0 0 FrameStrobe[7]
port 81 nsew signal input
flabel metal2 s 15290 0 15346 56 0 FreeSans 224 0 0 0 FrameStrobe[8]
port 82 nsew signal input
flabel metal2 s 16854 0 16910 56 0 FreeSans 224 0 0 0 FrameStrobe[9]
port 83 nsew signal input
flabel metal2 s 24306 11194 24362 11250 0 FreeSans 224 0 0 0 FrameStrobe_O[0]
port 84 nsew signal output
flabel metal2 s 27066 11194 27122 11250 0 FreeSans 224 0 0 0 FrameStrobe_O[10]
port 85 nsew signal output
flabel metal2 s 27342 11194 27398 11250 0 FreeSans 224 0 0 0 FrameStrobe_O[11]
port 86 nsew signal output
flabel metal2 s 27618 11194 27674 11250 0 FreeSans 224 0 0 0 FrameStrobe_O[12]
port 87 nsew signal output
flabel metal2 s 27894 11194 27950 11250 0 FreeSans 224 0 0 0 FrameStrobe_O[13]
port 88 nsew signal output
flabel metal2 s 28170 11194 28226 11250 0 FreeSans 224 0 0 0 FrameStrobe_O[14]
port 89 nsew signal output
flabel metal2 s 28446 11194 28502 11250 0 FreeSans 224 0 0 0 FrameStrobe_O[15]
port 90 nsew signal output
flabel metal2 s 28722 11194 28778 11250 0 FreeSans 224 0 0 0 FrameStrobe_O[16]
port 91 nsew signal output
flabel metal2 s 28998 11194 29054 11250 0 FreeSans 224 0 0 0 FrameStrobe_O[17]
port 92 nsew signal output
flabel metal2 s 29274 11194 29330 11250 0 FreeSans 224 0 0 0 FrameStrobe_O[18]
port 93 nsew signal output
flabel metal2 s 29550 11194 29606 11250 0 FreeSans 224 0 0 0 FrameStrobe_O[19]
port 94 nsew signal output
flabel metal2 s 24582 11194 24638 11250 0 FreeSans 224 0 0 0 FrameStrobe_O[1]
port 95 nsew signal output
flabel metal2 s 24858 11194 24914 11250 0 FreeSans 224 0 0 0 FrameStrobe_O[2]
port 96 nsew signal output
flabel metal2 s 25134 11194 25190 11250 0 FreeSans 224 0 0 0 FrameStrobe_O[3]
port 97 nsew signal output
flabel metal2 s 25410 11194 25466 11250 0 FreeSans 224 0 0 0 FrameStrobe_O[4]
port 98 nsew signal output
flabel metal2 s 25686 11194 25742 11250 0 FreeSans 224 0 0 0 FrameStrobe_O[5]
port 99 nsew signal output
flabel metal2 s 25962 11194 26018 11250 0 FreeSans 224 0 0 0 FrameStrobe_O[6]
port 100 nsew signal output
flabel metal2 s 26238 11194 26294 11250 0 FreeSans 224 0 0 0 FrameStrobe_O[7]
port 101 nsew signal output
flabel metal2 s 26514 11194 26570 11250 0 FreeSans 224 0 0 0 FrameStrobe_O[8]
port 102 nsew signal output
flabel metal2 s 26790 11194 26846 11250 0 FreeSans 224 0 0 0 FrameStrobe_O[9]
port 103 nsew signal output
flabel metal2 s 4158 11194 4214 11250 0 FreeSans 224 0 0 0 N1BEG[0]
port 104 nsew signal output
flabel metal2 s 4434 11194 4490 11250 0 FreeSans 224 0 0 0 N1BEG[1]
port 105 nsew signal output
flabel metal2 s 4710 11194 4766 11250 0 FreeSans 224 0 0 0 N1BEG[2]
port 106 nsew signal output
flabel metal2 s 4986 11194 5042 11250 0 FreeSans 224 0 0 0 N1BEG[3]
port 107 nsew signal output
flabel metal2 s 5262 11194 5318 11250 0 FreeSans 224 0 0 0 N2BEG[0]
port 108 nsew signal output
flabel metal2 s 5538 11194 5594 11250 0 FreeSans 224 0 0 0 N2BEG[1]
port 109 nsew signal output
flabel metal2 s 5814 11194 5870 11250 0 FreeSans 224 0 0 0 N2BEG[2]
port 110 nsew signal output
flabel metal2 s 6090 11194 6146 11250 0 FreeSans 224 0 0 0 N2BEG[3]
port 111 nsew signal output
flabel metal2 s 6366 11194 6422 11250 0 FreeSans 224 0 0 0 N2BEG[4]
port 112 nsew signal output
flabel metal2 s 6642 11194 6698 11250 0 FreeSans 224 0 0 0 N2BEG[5]
port 113 nsew signal output
flabel metal2 s 6918 11194 6974 11250 0 FreeSans 224 0 0 0 N2BEG[6]
port 114 nsew signal output
flabel metal2 s 7194 11194 7250 11250 0 FreeSans 224 0 0 0 N2BEG[7]
port 115 nsew signal output
flabel metal2 s 7470 11194 7526 11250 0 FreeSans 224 0 0 0 N2BEGb[0]
port 116 nsew signal output
flabel metal2 s 7746 11194 7802 11250 0 FreeSans 224 0 0 0 N2BEGb[1]
port 117 nsew signal output
flabel metal2 s 8022 11194 8078 11250 0 FreeSans 224 0 0 0 N2BEGb[2]
port 118 nsew signal output
flabel metal2 s 8298 11194 8354 11250 0 FreeSans 224 0 0 0 N2BEGb[3]
port 119 nsew signal output
flabel metal2 s 8574 11194 8630 11250 0 FreeSans 224 0 0 0 N2BEGb[4]
port 120 nsew signal output
flabel metal2 s 8850 11194 8906 11250 0 FreeSans 224 0 0 0 N2BEGb[5]
port 121 nsew signal output
flabel metal2 s 9126 11194 9182 11250 0 FreeSans 224 0 0 0 N2BEGb[6]
port 122 nsew signal output
flabel metal2 s 9402 11194 9458 11250 0 FreeSans 224 0 0 0 N2BEGb[7]
port 123 nsew signal output
flabel metal2 s 9678 11194 9734 11250 0 FreeSans 224 0 0 0 N4BEG[0]
port 124 nsew signal output
flabel metal2 s 12438 11194 12494 11250 0 FreeSans 224 0 0 0 N4BEG[10]
port 125 nsew signal output
flabel metal2 s 12714 11194 12770 11250 0 FreeSans 224 0 0 0 N4BEG[11]
port 126 nsew signal output
flabel metal2 s 12990 11194 13046 11250 0 FreeSans 224 0 0 0 N4BEG[12]
port 127 nsew signal output
flabel metal2 s 13266 11194 13322 11250 0 FreeSans 224 0 0 0 N4BEG[13]
port 128 nsew signal output
flabel metal2 s 13542 11194 13598 11250 0 FreeSans 224 0 0 0 N4BEG[14]
port 129 nsew signal output
flabel metal2 s 13818 11194 13874 11250 0 FreeSans 224 0 0 0 N4BEG[15]
port 130 nsew signal output
flabel metal2 s 9954 11194 10010 11250 0 FreeSans 224 0 0 0 N4BEG[1]
port 131 nsew signal output
flabel metal2 s 10230 11194 10286 11250 0 FreeSans 224 0 0 0 N4BEG[2]
port 132 nsew signal output
flabel metal2 s 10506 11194 10562 11250 0 FreeSans 224 0 0 0 N4BEG[3]
port 133 nsew signal output
flabel metal2 s 10782 11194 10838 11250 0 FreeSans 224 0 0 0 N4BEG[4]
port 134 nsew signal output
flabel metal2 s 11058 11194 11114 11250 0 FreeSans 224 0 0 0 N4BEG[5]
port 135 nsew signal output
flabel metal2 s 11334 11194 11390 11250 0 FreeSans 224 0 0 0 N4BEG[6]
port 136 nsew signal output
flabel metal2 s 11610 11194 11666 11250 0 FreeSans 224 0 0 0 N4BEG[7]
port 137 nsew signal output
flabel metal2 s 11886 11194 11942 11250 0 FreeSans 224 0 0 0 N4BEG[8]
port 138 nsew signal output
flabel metal2 s 12162 11194 12218 11250 0 FreeSans 224 0 0 0 N4BEG[9]
port 139 nsew signal output
flabel metal2 s 14094 11194 14150 11250 0 FreeSans 224 0 0 0 S1END[0]
port 140 nsew signal input
flabel metal2 s 14370 11194 14426 11250 0 FreeSans 224 0 0 0 S1END[1]
port 141 nsew signal input
flabel metal2 s 14646 11194 14702 11250 0 FreeSans 224 0 0 0 S1END[2]
port 142 nsew signal input
flabel metal2 s 14922 11194 14978 11250 0 FreeSans 224 0 0 0 S1END[3]
port 143 nsew signal input
flabel metal2 s 17406 11194 17462 11250 0 FreeSans 224 0 0 0 S2END[0]
port 144 nsew signal input
flabel metal2 s 17682 11194 17738 11250 0 FreeSans 224 0 0 0 S2END[1]
port 145 nsew signal input
flabel metal2 s 17958 11194 18014 11250 0 FreeSans 224 0 0 0 S2END[2]
port 146 nsew signal input
flabel metal2 s 18234 11194 18290 11250 0 FreeSans 224 0 0 0 S2END[3]
port 147 nsew signal input
flabel metal2 s 18510 11194 18566 11250 0 FreeSans 224 0 0 0 S2END[4]
port 148 nsew signal input
flabel metal2 s 18786 11194 18842 11250 0 FreeSans 224 0 0 0 S2END[5]
port 149 nsew signal input
flabel metal2 s 19062 11194 19118 11250 0 FreeSans 224 0 0 0 S2END[6]
port 150 nsew signal input
flabel metal2 s 19338 11194 19394 11250 0 FreeSans 224 0 0 0 S2END[7]
port 151 nsew signal input
flabel metal2 s 15198 11194 15254 11250 0 FreeSans 224 0 0 0 S2MID[0]
port 152 nsew signal input
flabel metal2 s 15474 11194 15530 11250 0 FreeSans 224 0 0 0 S2MID[1]
port 153 nsew signal input
flabel metal2 s 15750 11194 15806 11250 0 FreeSans 224 0 0 0 S2MID[2]
port 154 nsew signal input
flabel metal2 s 16026 11194 16082 11250 0 FreeSans 224 0 0 0 S2MID[3]
port 155 nsew signal input
flabel metal2 s 16302 11194 16358 11250 0 FreeSans 224 0 0 0 S2MID[4]
port 156 nsew signal input
flabel metal2 s 16578 11194 16634 11250 0 FreeSans 224 0 0 0 S2MID[5]
port 157 nsew signal input
flabel metal2 s 16854 11194 16910 11250 0 FreeSans 224 0 0 0 S2MID[6]
port 158 nsew signal input
flabel metal2 s 17130 11194 17186 11250 0 FreeSans 224 0 0 0 S2MID[7]
port 159 nsew signal input
flabel metal2 s 19614 11194 19670 11250 0 FreeSans 224 0 0 0 S4END[0]
port 160 nsew signal input
flabel metal2 s 22374 11194 22430 11250 0 FreeSans 224 0 0 0 S4END[10]
port 161 nsew signal input
flabel metal2 s 22650 11194 22706 11250 0 FreeSans 224 0 0 0 S4END[11]
port 162 nsew signal input
flabel metal2 s 22926 11194 22982 11250 0 FreeSans 224 0 0 0 S4END[12]
port 163 nsew signal input
flabel metal2 s 23202 11194 23258 11250 0 FreeSans 224 0 0 0 S4END[13]
port 164 nsew signal input
flabel metal2 s 23478 11194 23534 11250 0 FreeSans 224 0 0 0 S4END[14]
port 165 nsew signal input
flabel metal2 s 23754 11194 23810 11250 0 FreeSans 224 0 0 0 S4END[15]
port 166 nsew signal input
flabel metal2 s 19890 11194 19946 11250 0 FreeSans 224 0 0 0 S4END[1]
port 167 nsew signal input
flabel metal2 s 20166 11194 20222 11250 0 FreeSans 224 0 0 0 S4END[2]
port 168 nsew signal input
flabel metal2 s 20442 11194 20498 11250 0 FreeSans 224 0 0 0 S4END[3]
port 169 nsew signal input
flabel metal2 s 20718 11194 20774 11250 0 FreeSans 224 0 0 0 S4END[4]
port 170 nsew signal input
flabel metal2 s 20994 11194 21050 11250 0 FreeSans 224 0 0 0 S4END[5]
port 171 nsew signal input
flabel metal2 s 21270 11194 21326 11250 0 FreeSans 224 0 0 0 S4END[6]
port 172 nsew signal input
flabel metal2 s 21546 11194 21602 11250 0 FreeSans 224 0 0 0 S4END[7]
port 173 nsew signal input
flabel metal2 s 21822 11194 21878 11250 0 FreeSans 224 0 0 0 S4END[8]
port 174 nsew signal input
flabel metal2 s 22098 11194 22154 11250 0 FreeSans 224 0 0 0 S4END[9]
port 175 nsew signal input
flabel metal2 s 1214 0 1270 56 0 FreeSans 224 0 0 0 UserCLK
port 176 nsew signal input
flabel metal2 s 24030 11194 24086 11250 0 FreeSans 224 0 0 0 UserCLKo
port 177 nsew signal output
flabel metal4 s 3004 0 3324 11250 0 FreeSans 1920 90 0 0 VGND
port 178 nsew ground bidirectional
flabel metal4 s 3004 0 3324 60 0 FreeSans 480 0 0 0 VGND
port 178 nsew ground bidirectional
flabel metal4 s 3004 11190 3324 11250 0 FreeSans 480 0 0 0 VGND
port 178 nsew ground bidirectional
flabel metal4 s 9004 0 9324 11250 0 FreeSans 1920 90 0 0 VGND
port 178 nsew ground bidirectional
flabel metal4 s 9004 0 9324 60 0 FreeSans 480 0 0 0 VGND
port 178 nsew ground bidirectional
flabel metal4 s 9004 11190 9324 11250 0 FreeSans 480 0 0 0 VGND
port 178 nsew ground bidirectional
flabel metal4 s 15004 0 15324 11250 0 FreeSans 1920 90 0 0 VGND
port 178 nsew ground bidirectional
flabel metal4 s 15004 0 15324 60 0 FreeSans 480 0 0 0 VGND
port 178 nsew ground bidirectional
flabel metal4 s 15004 11190 15324 11250 0 FreeSans 480 0 0 0 VGND
port 178 nsew ground bidirectional
flabel metal4 s 21004 0 21324 11250 0 FreeSans 1920 90 0 0 VGND
port 178 nsew ground bidirectional
flabel metal4 s 21004 0 21324 60 0 FreeSans 480 0 0 0 VGND
port 178 nsew ground bidirectional
flabel metal4 s 21004 11190 21324 11250 0 FreeSans 480 0 0 0 VGND
port 178 nsew ground bidirectional
flabel metal4 s 27004 0 27324 11250 0 FreeSans 1920 90 0 0 VGND
port 178 nsew ground bidirectional
flabel metal4 s 27004 0 27324 60 0 FreeSans 480 0 0 0 VGND
port 178 nsew ground bidirectional
flabel metal4 s 27004 11190 27324 11250 0 FreeSans 480 0 0 0 VGND
port 178 nsew ground bidirectional
flabel metal4 s 1944 0 2264 11250 0 FreeSans 1920 90 0 0 VPWR
port 179 nsew power bidirectional
flabel metal4 s 1944 0 2264 60 0 FreeSans 480 0 0 0 VPWR
port 179 nsew power bidirectional
flabel metal4 s 1944 11190 2264 11250 0 FreeSans 480 0 0 0 VPWR
port 179 nsew power bidirectional
flabel metal4 s 7944 0 8264 11250 0 FreeSans 1920 90 0 0 VPWR
port 179 nsew power bidirectional
flabel metal4 s 7944 0 8264 60 0 FreeSans 480 0 0 0 VPWR
port 179 nsew power bidirectional
flabel metal4 s 7944 11190 8264 11250 0 FreeSans 480 0 0 0 VPWR
port 179 nsew power bidirectional
flabel metal4 s 13944 0 14264 11250 0 FreeSans 1920 90 0 0 VPWR
port 179 nsew power bidirectional
flabel metal4 s 13944 0 14264 60 0 FreeSans 480 0 0 0 VPWR
port 179 nsew power bidirectional
flabel metal4 s 13944 11190 14264 11250 0 FreeSans 480 0 0 0 VPWR
port 179 nsew power bidirectional
flabel metal4 s 19944 0 20264 11250 0 FreeSans 1920 90 0 0 VPWR
port 179 nsew power bidirectional
flabel metal4 s 19944 0 20264 60 0 FreeSans 480 0 0 0 VPWR
port 179 nsew power bidirectional
flabel metal4 s 19944 11190 20264 11250 0 FreeSans 480 0 0 0 VPWR
port 179 nsew power bidirectional
flabel metal4 s 25944 0 26264 11250 0 FreeSans 1920 90 0 0 VPWR
port 179 nsew power bidirectional
flabel metal4 s 25944 0 26264 60 0 FreeSans 480 0 0 0 VPWR
port 179 nsew power bidirectional
flabel metal4 s 25944 11190 26264 11250 0 FreeSans 480 0 0 0 VPWR
port 179 nsew power bidirectional
flabel metal4 s 31944 0 32264 11250 0 FreeSans 1920 90 0 0 VPWR
port 179 nsew power bidirectional
flabel metal4 s 31944 0 32264 60 0 FreeSans 480 0 0 0 VPWR
port 179 nsew power bidirectional
flabel metal4 s 31944 11190 32264 11250 0 FreeSans 480 0 0 0 VPWR
port 179 nsew power bidirectional
rlabel metal1 16836 8704 16836 8704 0 VGND
rlabel metal1 16836 8160 16836 8160 0 VPWR
rlabel metal3 620 1428 620 1428 0 FrameData[0]
rlabel metal2 19550 3825 19550 3825 0 FrameData[10]
rlabel metal2 19274 3808 19274 3808 0 FrameData[11]
rlabel metal2 18170 4199 18170 4199 0 FrameData[12]
rlabel metal3 942 4964 942 4964 0 FrameData[13]
rlabel metal3 712 5236 712 5236 0 FrameData[14]
rlabel metal3 1425 5508 1425 5508 0 FrameData[15]
rlabel metal1 14398 3638 14398 3638 0 FrameData[16]
rlabel metal3 919 6052 919 6052 0 FrameData[17]
rlabel metal2 12466 5219 12466 5219 0 FrameData[18]
rlabel metal3 344 6596 344 6596 0 FrameData[19]
rlabel metal3 4806 1700 4806 1700 0 FrameData[1]
rlabel metal2 16238 6273 16238 6273 0 FrameData[20]
rlabel metal3 919 7140 919 7140 0 FrameData[21]
rlabel metal1 25898 6698 25898 6698 0 FrameData[22]
rlabel metal2 16698 7293 16698 7293 0 FrameData[23]
rlabel metal2 24518 7735 24518 7735 0 FrameData[24]
rlabel metal3 919 8228 919 8228 0 FrameData[25]
rlabel metal1 26358 7446 26358 7446 0 FrameData[26]
rlabel metal2 20976 6766 20976 6766 0 FrameData[27]
rlabel metal1 21574 6766 21574 6766 0 FrameData[28]
rlabel metal1 16192 6766 16192 6766 0 FrameData[29]
rlabel metal3 4852 1972 4852 1972 0 FrameData[2]
rlabel metal2 19366 7378 19366 7378 0 FrameData[30]
rlabel metal1 27186 7446 27186 7446 0 FrameData[31]
rlabel metal3 1471 2244 1471 2244 0 FrameData[3]
rlabel metal3 712 2516 712 2516 0 FrameData[4]
rlabel metal3 942 2788 942 2788 0 FrameData[5]
rlabel metal2 16882 3213 16882 3213 0 FrameData[6]
rlabel metal3 1034 3332 1034 3332 0 FrameData[7]
rlabel metal1 18630 3570 18630 3570 0 FrameData[8]
rlabel metal3 919 3876 919 3876 0 FrameData[9]
rlabel metal2 31510 1853 31510 1853 0 FrameData_O[0]
rlabel metal3 32723 4148 32723 4148 0 FrameData_O[10]
rlabel metal3 32907 4420 32907 4420 0 FrameData_O[11]
rlabel metal3 32585 4692 32585 4692 0 FrameData_O[12]
rlabel metal3 33275 4964 33275 4964 0 FrameData_O[13]
rlabel metal3 32861 5236 32861 5236 0 FrameData_O[14]
rlabel metal3 32723 5508 32723 5508 0 FrameData_O[15]
rlabel metal3 32907 5780 32907 5780 0 FrameData_O[16]
rlabel metal3 33160 6052 33160 6052 0 FrameData_O[17]
rlabel metal3 32769 6324 32769 6324 0 FrameData_O[18]
rlabel via2 31418 6613 31418 6613 0 FrameData_O[19]
rlabel metal2 31142 1989 31142 1989 0 FrameData_O[1]
rlabel metal2 31786 6749 31786 6749 0 FrameData_O[20]
rlabel metal3 33229 7140 33229 7140 0 FrameData_O[21]
rlabel metal3 32723 7412 32723 7412 0 FrameData_O[22]
rlabel metal3 32907 7684 32907 7684 0 FrameData_O[23]
rlabel metal3 32769 7956 32769 7956 0 FrameData_O[24]
rlabel metal3 33137 8228 33137 8228 0 FrameData_O[25]
rlabel metal3 32401 8500 32401 8500 0 FrameData_O[26]
rlabel metal2 31418 8415 31418 8415 0 FrameData_O[27]
rlabel metal2 31050 8551 31050 8551 0 FrameData_O[28]
rlabel metal2 31510 8415 31510 8415 0 FrameData_O[29]
rlabel metal2 30774 2125 30774 2125 0 FrameData_O[2]
rlabel metal2 30682 8823 30682 8823 0 FrameData_O[30]
rlabel metal1 32246 6630 32246 6630 0 FrameData_O[31]
rlabel metal3 32769 2244 32769 2244 0 FrameData_O[3]
rlabel metal3 32723 2516 32723 2516 0 FrameData_O[4]
rlabel metal3 33275 2788 33275 2788 0 FrameData_O[5]
rlabel metal3 32723 3060 32723 3060 0 FrameData_O[6]
rlabel metal3 32907 3332 32907 3332 0 FrameData_O[7]
rlabel metal3 32585 3604 32585 3604 0 FrameData_O[8]
rlabel metal3 33275 3876 33275 3876 0 FrameData_O[9]
rlabel metal2 2806 106 2806 106 0 FrameStrobe[0]
rlabel metal1 19872 5202 19872 5202 0 FrameStrobe[10]
rlabel metal2 20010 55 20010 55 0 FrameStrobe[11]
rlabel metal2 21574 3166 21574 3166 0 FrameStrobe[12]
rlabel metal1 22586 7378 22586 7378 0 FrameStrobe[13]
rlabel metal1 23828 6290 23828 6290 0 FrameStrobe[14]
rlabel metal2 23690 6596 23690 6596 0 FrameStrobe[15]
rlabel metal2 24426 6528 24426 6528 0 FrameStrobe[16]
rlabel metal1 27922 6766 27922 6766 0 FrameStrobe[17]
rlabel metal1 29762 6290 29762 6290 0 FrameStrobe[18]
rlabel metal2 32522 3132 32522 3132 0 FrameStrobe[19]
rlabel metal2 14582 3332 14582 3332 0 FrameStrobe[1]
rlabel metal2 16606 3196 16606 3196 0 FrameStrobe[2]
rlabel metal1 8464 3570 8464 3570 0 FrameStrobe[3]
rlabel metal2 9062 123 9062 123 0 FrameStrobe[4]
rlabel via2 10626 55 10626 55 0 FrameStrobe[5]
rlabel metal1 25852 3502 25852 3502 0 FrameStrobe[6]
rlabel metal2 23506 3553 23506 3553 0 FrameStrobe[7]
rlabel metal2 23782 4301 23782 4301 0 FrameStrobe[8]
rlabel metal2 16882 1143 16882 1143 0 FrameStrobe[9]
rlabel metal1 24518 8602 24518 8602 0 FrameStrobe_O[0]
rlabel metal2 27370 8755 27370 8755 0 FrameStrobe_O[10]
rlabel metal1 27876 8602 27876 8602 0 FrameStrobe_O[11]
rlabel metal2 28658 8840 28658 8840 0 FrameStrobe_O[12]
rlabel metal1 29026 8568 29026 8568 0 FrameStrobe_O[13]
rlabel metal1 28336 8058 28336 8058 0 FrameStrobe_O[14]
rlabel metal1 28704 8058 28704 8058 0 FrameStrobe_O[15]
rlabel metal1 29256 8330 29256 8330 0 FrameStrobe_O[16]
rlabel metal1 30130 8364 30130 8364 0 FrameStrobe_O[17]
rlabel metal1 29532 8058 29532 8058 0 FrameStrobe_O[18]
rlabel metal1 29992 8602 29992 8602 0 FrameStrobe_O[19]
rlabel metal1 24840 8602 24840 8602 0 FrameStrobe_O[1]
rlabel metal1 25208 8330 25208 8330 0 FrameStrobe_O[2]
rlabel metal1 25438 8602 25438 8602 0 FrameStrobe_O[3]
rlabel metal1 25760 8330 25760 8330 0 FrameStrobe_O[4]
rlabel metal2 25714 10414 25714 10414 0 FrameStrobe_O[5]
rlabel metal1 26036 8058 26036 8058 0 FrameStrobe_O[6]
rlabel metal1 26726 8602 26726 8602 0 FrameStrobe_O[7]
rlabel metal1 27094 8330 27094 8330 0 FrameStrobe_O[8]
rlabel metal1 27876 8330 27876 8330 0 FrameStrobe_O[9]
rlabel metal1 4278 8058 4278 8058 0 N1BEG[0]
rlabel metal1 4324 8602 4324 8602 0 N1BEG[1]
rlabel metal1 4646 8602 4646 8602 0 N1BEG[2]
rlabel metal1 4968 8602 4968 8602 0 N1BEG[3]
rlabel metal1 5428 8058 5428 8058 0 N2BEG[0]
rlabel metal1 5474 8602 5474 8602 0 N2BEG[1]
rlabel metal1 5750 8602 5750 8602 0 N2BEG[2]
rlabel metal1 6210 8058 6210 8058 0 N2BEG[3]
rlabel metal1 6210 8602 6210 8602 0 N2BEG[4]
rlabel metal1 6762 8058 6762 8058 0 N2BEG[5]
rlabel metal1 6854 8602 6854 8602 0 N2BEG[6]
rlabel metal1 7176 8602 7176 8602 0 N2BEG[7]
rlabel metal1 7636 8058 7636 8058 0 N2BEGb[0]
rlabel metal1 7682 8602 7682 8602 0 N2BEGb[1]
rlabel metal1 8004 8602 8004 8602 0 N2BEGb[2]
rlabel metal1 8418 8058 8418 8058 0 N2BEGb[3]
rlabel metal1 8372 8602 8372 8602 0 N2BEGb[4]
rlabel metal1 8694 8602 8694 8602 0 N2BEGb[5]
rlabel metal1 9108 8058 9108 8058 0 N2BEGb[6]
rlabel metal1 9384 8602 9384 8602 0 N2BEGb[7]
rlabel metal1 9798 8058 9798 8058 0 N4BEG[0]
rlabel metal2 12466 9904 12466 9904 0 N4BEG[10]
rlabel metal2 12742 9904 12742 9904 0 N4BEG[11]
rlabel metal1 13064 8602 13064 8602 0 N4BEG[12]
rlabel metal1 13386 8602 13386 8602 0 N4BEG[13]
rlabel metal1 13708 8602 13708 8602 0 N4BEG[14]
rlabel metal1 14122 8602 14122 8602 0 N4BEG[15]
rlabel metal1 9844 8602 9844 8602 0 N4BEG[1]
rlabel metal1 10166 8602 10166 8602 0 N4BEG[2]
rlabel metal1 10488 8602 10488 8602 0 N4BEG[3]
rlabel metal1 10902 8058 10902 8058 0 N4BEG[4]
rlabel metal1 10948 8602 10948 8602 0 N4BEG[5]
rlabel metal1 11454 8058 11454 8058 0 N4BEG[6]
rlabel metal1 11408 8602 11408 8602 0 N4BEG[7]
rlabel metal1 12006 8058 12006 8058 0 N4BEG[8]
rlabel metal1 12098 8602 12098 8602 0 N4BEG[9]
rlabel metal2 14122 10465 14122 10465 0 S1END[0]
rlabel metal2 14398 10465 14398 10465 0 S1END[1]
rlabel metal2 14674 10601 14674 10601 0 S1END[2]
rlabel metal2 14950 11009 14950 11009 0 S1END[3]
rlabel metal2 17434 9224 17434 9224 0 S2END[0]
rlabel metal2 17710 9190 17710 9190 0 S2END[1]
rlabel metal2 17986 10210 17986 10210 0 S2END[2]
rlabel metal2 18262 10261 18262 10261 0 S2END[3]
rlabel metal2 18538 9649 18538 9649 0 S2END[4]
rlabel metal2 18814 10312 18814 10312 0 S2END[5]
rlabel metal2 19090 10805 19090 10805 0 S2END[6]
rlabel metal2 19366 10618 19366 10618 0 S2END[7]
rlabel metal2 15226 10057 15226 10057 0 S2MID[0]
rlabel metal2 15502 10193 15502 10193 0 S2MID[1]
rlabel metal2 15778 9989 15778 9989 0 S2MID[2]
rlabel metal2 16054 8697 16054 8697 0 S2MID[3]
rlabel metal2 16330 9853 16330 9853 0 S2MID[4]
rlabel metal2 16606 9802 16606 9802 0 S2MID[5]
rlabel metal2 16882 9853 16882 9853 0 S2MID[6]
rlabel metal2 17158 8442 17158 8442 0 S2MID[7]
rlabel metal2 19642 8748 19642 8748 0 S4END[0]
rlabel metal2 22126 6357 22126 6357 0 S4END[10]
rlabel metal2 22678 10125 22678 10125 0 S4END[11]
rlabel metal1 22586 6630 22586 6630 0 S4END[12]
rlabel metal2 23230 8680 23230 8680 0 S4END[13]
rlabel metal2 23552 6732 23552 6732 0 S4END[14]
rlabel metal1 23506 6766 23506 6766 0 S4END[15]
rlabel metal2 19918 10193 19918 10193 0 S4END[1]
rlabel metal2 20194 10125 20194 10125 0 S4END[2]
rlabel metal2 20470 10057 20470 10057 0 S4END[3]
rlabel metal2 20746 10397 20746 10397 0 S4END[4]
rlabel metal2 21022 10244 21022 10244 0 S4END[5]
rlabel metal2 21298 10006 21298 10006 0 S4END[6]
rlabel metal2 21574 10125 21574 10125 0 S4END[7]
rlabel metal2 21850 9088 21850 9088 0 S4END[8]
rlabel metal2 22126 11162 22126 11162 0 S4END[9]
rlabel metal2 1242 55 1242 55 0 UserCLK
rlabel metal2 24058 9904 24058 9904 0 UserCLKo
rlabel metal1 26726 2380 26726 2380 0 net1
rlabel metal2 31418 5542 31418 5542 0 net10
rlabel metal1 22770 4556 22770 4556 0 net11
rlabel metal2 11546 2924 11546 2924 0 net12
rlabel metal2 31694 6188 31694 6188 0 net13
rlabel metal1 31050 7242 31050 7242 0 net14
rlabel metal1 27002 6630 27002 6630 0 net15
rlabel metal1 24610 7480 24610 7480 0 net16
rlabel metal2 27462 7752 27462 7752 0 net17
rlabel metal2 26266 7480 26266 7480 0 net18
rlabel metal1 27738 7242 27738 7242 0 net19
rlabel metal2 29026 4080 29026 4080 0 net2
rlabel metal2 22862 6783 22862 6783 0 net20
rlabel metal1 30774 7854 30774 7854 0 net21
rlabel metal1 31326 7344 31326 7344 0 net22
rlabel metal2 12190 2958 12190 2958 0 net23
rlabel metal2 30498 7038 30498 7038 0 net24
rlabel metal1 31142 6834 31142 6834 0 net25
rlabel metal2 12466 2992 12466 2992 0 net26
rlabel metal1 30866 3026 30866 3026 0 net27
rlabel metal2 31694 3247 31694 3247 0 net28
rlabel metal2 31602 3298 31602 3298 0 net29
rlabel metal2 31970 4420 31970 4420 0 net3
rlabel metal2 31970 3332 31970 3332 0 net30
rlabel metal2 26910 3570 26910 3570 0 net31
rlabel metal2 31418 3502 31418 3502 0 net32
rlabel metal1 23414 8398 23414 8398 0 net33
rlabel metal1 27186 7820 27186 7820 0 net34
rlabel metal2 28106 8738 28106 8738 0 net35
rlabel metal2 22310 5950 22310 5950 0 net36
rlabel metal1 22954 7174 22954 7174 0 net37
rlabel metal2 23598 6392 23598 6392 0 net38
rlabel metal2 23874 6358 23874 6358 0 net39
rlabel metal1 26220 5236 26220 5236 0 net4
rlabel metal1 25254 6834 25254 6834 0 net40
rlabel metal1 26680 6970 26680 6970 0 net41
rlabel metal1 28934 6426 28934 6426 0 net42
rlabel metal1 30728 6426 30728 6426 0 net43
rlabel metal1 24150 8568 24150 8568 0 net44
rlabel metal2 25070 8738 25070 8738 0 net45
rlabel metal2 25530 6256 25530 6256 0 net46
rlabel metal1 23046 3366 23046 3366 0 net47
rlabel metal1 26082 3366 26082 3366 0 net48
rlabel metal1 26036 3706 26036 3706 0 net49
rlabel metal2 31694 4964 31694 4964 0 net5
rlabel metal2 25530 3808 25530 3808 0 net50
rlabel metal1 24380 4454 24380 4454 0 net51
rlabel metal1 22862 4488 22862 4488 0 net52
rlabel metal2 6302 7378 6302 7378 0 net53
rlabel metal1 6118 6630 6118 6630 0 net54
rlabel metal1 6348 6154 6348 6154 0 net55
rlabel metal1 9062 6154 9062 6154 0 net56
rlabel metal1 4922 6970 4922 6970 0 net57
rlabel metal1 5244 6426 5244 6426 0 net58
rlabel metal1 6256 6426 6256 6426 0 net59
rlabel metal2 31234 4828 31234 4828 0 net6
rlabel metal1 7314 6426 7314 6426 0 net60
rlabel metal1 7590 5542 7590 5542 0 net61
rlabel metal1 9752 6426 9752 6426 0 net62
rlabel metal2 11086 6137 11086 6137 0 net63
rlabel metal1 7912 5338 7912 5338 0 net64
rlabel metal1 6992 5882 6992 5882 0 net65
rlabel metal2 7406 7174 7406 7174 0 net66
rlabel metal1 7728 5882 7728 5882 0 net67
rlabel metal2 8694 7140 8694 7140 0 net68
rlabel metal1 9016 6426 9016 6426 0 net69
rlabel metal2 31326 4556 31326 4556 0 net7
rlabel metal2 10304 6426 10304 6426 0 net70
rlabel metal1 9752 6630 9752 6630 0 net71
rlabel metal1 10764 6154 10764 6154 0 net72
rlabel metal1 20792 6970 20792 6970 0 net73
rlabel metal2 12190 7310 12190 7310 0 net74
rlabel metal2 12558 8874 12558 8874 0 net75
rlabel metal1 12926 8432 12926 8432 0 net76
rlabel metal1 13294 8500 13294 8500 0 net77
rlabel metal2 13386 7582 13386 7582 0 net78
rlabel metal2 14122 8738 14122 8738 0 net79
rlabel metal2 31878 4658 31878 4658 0 net8
rlabel metal1 19550 6970 19550 6970 0 net80
rlabel metal2 18262 7854 18262 7854 0 net81
rlabel metal2 17526 7480 17526 7480 0 net82
rlabel metal1 17158 6664 17158 6664 0 net83
rlabel metal2 15594 7752 15594 7752 0 net84
rlabel metal2 14398 7378 14398 7378 0 net85
rlabel metal2 13478 7718 13478 7718 0 net86
rlabel metal2 12650 7412 12650 7412 0 net87
rlabel metal2 11546 7548 11546 7548 0 net88
rlabel metal2 24242 6088 24242 6088 0 net89
rlabel metal2 31326 6086 31326 6086 0 net9
<< properties >>
string FIXED_BBOX 0 0 33750 11250
<< end >>
