magic
tech sky130A
magscale 1 2
timestamp 1740383397
<< viali >>
rect 2421 8585 2455 8619
rect 2697 8585 2731 8619
rect 3433 8585 3467 8619
rect 4261 8585 4295 8619
rect 4629 8585 4663 8619
rect 4997 8585 5031 8619
rect 5273 8585 5307 8619
rect 5641 8585 5675 8619
rect 6009 8585 6043 8619
rect 6745 8585 6779 8619
rect 7113 8585 7147 8619
rect 7481 8585 7515 8619
rect 7849 8585 7883 8619
rect 8217 8585 8251 8619
rect 8585 8585 8619 8619
rect 9321 8585 9355 8619
rect 9689 8585 9723 8619
rect 10057 8585 10091 8619
rect 10425 8585 10459 8619
rect 10793 8585 10827 8619
rect 11253 8585 11287 8619
rect 11713 8585 11747 8619
rect 12081 8585 12115 8619
rect 12817 8585 12851 8619
rect 13829 8585 13863 8619
rect 14473 8585 14507 8619
rect 14841 8585 14875 8619
rect 15209 8585 15243 8619
rect 15669 8585 15703 8619
rect 15945 8585 15979 8619
rect 16313 8585 16347 8619
rect 17049 8585 17083 8619
rect 17601 8585 17635 8619
rect 18797 8585 18831 8619
rect 19349 8585 19383 8619
rect 19625 8585 19659 8619
rect 21833 8585 21867 8619
rect 23765 8585 23799 8619
rect 25513 8585 25547 8619
rect 30481 8585 30515 8619
rect 32321 8585 32355 8619
rect 32781 8585 32815 8619
rect 33149 8585 33183 8619
rect 33517 8585 33551 8619
rect 34253 8585 34287 8619
rect 35541 8585 35575 8619
rect 36737 8585 36771 8619
rect 37841 8585 37875 8619
rect 38577 8585 38611 8619
rect 1409 8449 1443 8483
rect 1685 8449 1719 8483
rect 1961 8449 1995 8483
rect 2237 8449 2271 8483
rect 2513 8449 2547 8483
rect 3249 8449 3283 8483
rect 3617 8449 3651 8483
rect 4077 8449 4111 8483
rect 4445 8449 4479 8483
rect 4813 8449 4847 8483
rect 5457 8449 5491 8483
rect 5825 8449 5859 8483
rect 6193 8449 6227 8483
rect 6929 8449 6963 8483
rect 7297 8449 7331 8483
rect 7665 8449 7699 8483
rect 8033 8449 8067 8483
rect 8401 8449 8435 8483
rect 8769 8449 8803 8483
rect 9505 8449 9539 8483
rect 9873 8449 9907 8483
rect 10241 8449 10275 8483
rect 10609 8449 10643 8483
rect 10977 8449 11011 8483
rect 11069 8449 11103 8483
rect 11897 8449 11931 8483
rect 12265 8449 12299 8483
rect 12633 8449 12667 8483
rect 13001 8449 13035 8483
rect 13369 8449 13403 8483
rect 13461 8449 13495 8483
rect 13645 8449 13679 8483
rect 14657 8449 14691 8483
rect 15025 8449 15059 8483
rect 15393 8449 15427 8483
rect 15485 8449 15519 8483
rect 16129 8449 16163 8483
rect 16497 8449 16531 8483
rect 16865 8449 16899 8483
rect 17417 8449 17451 8483
rect 17785 8449 17819 8483
rect 18521 8449 18555 8483
rect 18613 8449 18647 8483
rect 18889 8449 18923 8483
rect 19533 8449 19567 8483
rect 19809 8449 19843 8483
rect 19901 8449 19935 8483
rect 21465 8449 21499 8483
rect 22017 8449 22051 8483
rect 22293 8449 22327 8483
rect 22385 8449 22419 8483
rect 22845 8449 22879 8483
rect 23121 8449 23155 8483
rect 23397 8449 23431 8483
rect 23489 8449 23523 8483
rect 23949 8449 23983 8483
rect 24225 8449 24259 8483
rect 24593 8449 24627 8483
rect 24869 8449 24903 8483
rect 25145 8449 25179 8483
rect 25421 8449 25455 8483
rect 25697 8449 25731 8483
rect 25789 8449 25823 8483
rect 28089 8449 28123 8483
rect 28181 8449 28215 8483
rect 29285 8449 29319 8483
rect 30665 8449 30699 8483
rect 32505 8449 32539 8483
rect 32597 8449 32631 8483
rect 32953 8449 32987 8483
rect 33333 8449 33367 8483
rect 33701 8449 33735 8483
rect 34069 8449 34103 8483
rect 34713 8449 34747 8483
rect 35081 8449 35115 8483
rect 35725 8449 35759 8483
rect 35817 8449 35851 8483
rect 36185 8449 36219 8483
rect 36553 8449 36587 8483
rect 37289 8449 37323 8483
rect 37657 8449 37691 8483
rect 38025 8449 38059 8483
rect 38393 8449 38427 8483
rect 39129 8449 39163 8483
rect 39221 8449 39255 8483
rect 28457 8381 28491 8415
rect 29561 8381 29595 8415
rect 29837 8381 29871 8415
rect 2145 8313 2179 8347
rect 3065 8313 3099 8347
rect 12449 8313 12483 8347
rect 13185 8313 13219 8347
rect 17969 8313 18003 8347
rect 18337 8313 18371 8347
rect 19073 8313 19107 8347
rect 20085 8313 20119 8347
rect 21281 8313 21315 8347
rect 22109 8313 22143 8347
rect 22569 8313 22603 8347
rect 23213 8313 23247 8347
rect 24041 8313 24075 8347
rect 24685 8313 24719 8347
rect 24961 8313 24995 8347
rect 25237 8313 25271 8347
rect 25973 8313 26007 8347
rect 27905 8313 27939 8347
rect 29101 8313 29135 8347
rect 33885 8313 33919 8347
rect 34897 8313 34931 8347
rect 35265 8313 35299 8347
rect 36001 8313 36035 8347
rect 38209 8313 38243 8347
rect 39037 8313 39071 8347
rect 39405 8313 39439 8347
rect 1593 8245 1627 8279
rect 1869 8245 1903 8279
rect 22661 8245 22695 8279
rect 22937 8245 22971 8279
rect 23673 8245 23707 8279
rect 24409 8245 24443 8279
rect 36369 8245 36403 8279
rect 37473 8245 37507 8279
rect 3433 8041 3467 8075
rect 4261 8041 4295 8075
rect 5181 8041 5215 8075
rect 6193 8041 6227 8075
rect 6745 8041 6779 8075
rect 7297 8041 7331 8075
rect 8493 8041 8527 8075
rect 9045 8041 9079 8075
rect 9505 8041 9539 8075
rect 10609 8041 10643 8075
rect 11437 8041 11471 8075
rect 11989 8041 12023 8075
rect 12909 8041 12943 8075
rect 13645 8041 13679 8075
rect 14473 8041 14507 8075
rect 15025 8041 15059 8075
rect 16221 8041 16255 8075
rect 17693 8041 17727 8075
rect 34897 8041 34931 8075
rect 35817 8041 35851 8075
rect 36369 8041 36403 8075
rect 36921 8041 36955 8075
rect 37933 8041 37967 8075
rect 38669 8041 38703 8075
rect 1869 7973 1903 8007
rect 18153 7973 18187 8007
rect 1409 7837 1443 7871
rect 1685 7837 1719 7871
rect 1961 7837 1995 7871
rect 2237 7837 2271 7871
rect 3617 7837 3651 7871
rect 4445 7837 4479 7871
rect 4997 7837 5031 7871
rect 6377 7837 6411 7871
rect 6929 7837 6963 7871
rect 7481 7837 7515 7871
rect 8309 7837 8343 7871
rect 9229 7837 9263 7871
rect 9689 7837 9723 7871
rect 10793 7837 10827 7871
rect 11621 7837 11655 7871
rect 12173 7837 12207 7871
rect 12725 7837 12759 7871
rect 13829 7837 13863 7871
rect 14657 7837 14691 7871
rect 15209 7837 15243 7871
rect 16037 7837 16071 7871
rect 17969 7837 18003 7871
rect 18429 7837 18463 7871
rect 28917 7837 28951 7871
rect 29193 7837 29227 7871
rect 29745 7837 29779 7871
rect 34713 7837 34747 7871
rect 35633 7837 35667 7871
rect 36185 7837 36219 7871
rect 36737 7837 36771 7871
rect 38117 7837 38151 7871
rect 38485 7837 38519 7871
rect 38853 7837 38887 7871
rect 39221 7837 39255 7871
rect 1593 7701 1627 7735
rect 2145 7701 2179 7735
rect 2421 7701 2455 7735
rect 18245 7701 18279 7735
rect 28733 7701 28767 7735
rect 29009 7701 29043 7735
rect 29561 7701 29595 7735
rect 39037 7701 39071 7735
rect 39405 7701 39439 7735
rect 1869 7497 1903 7531
rect 4077 7497 4111 7531
rect 4721 7497 4755 7531
rect 19165 7497 19199 7531
rect 21557 7497 21591 7531
rect 34437 7497 34471 7531
rect 38301 7497 38335 7531
rect 38669 7497 38703 7531
rect 39037 7497 39071 7531
rect 39405 7497 39439 7531
rect 22293 7429 22327 7463
rect 22385 7429 22419 7463
rect 1409 7361 1443 7395
rect 1685 7361 1719 7395
rect 1961 7361 1995 7395
rect 2881 7361 2915 7395
rect 3249 7361 3283 7395
rect 3709 7361 3743 7395
rect 3893 7361 3927 7395
rect 4261 7361 4295 7395
rect 4537 7361 4571 7395
rect 14105 7361 14139 7395
rect 19349 7361 19383 7395
rect 20821 7361 20855 7395
rect 21925 7361 21959 7395
rect 22109 7361 22143 7395
rect 22569 7361 22603 7395
rect 22845 7361 22879 7395
rect 23029 7361 23063 7395
rect 31217 7361 31251 7395
rect 31493 7361 31527 7395
rect 31769 7361 31803 7395
rect 32321 7361 32355 7395
rect 32597 7361 32631 7395
rect 32873 7361 32907 7395
rect 33517 7361 33551 7395
rect 34253 7361 34287 7395
rect 37381 7361 37415 7395
rect 37473 7361 37507 7395
rect 37749 7361 37783 7395
rect 38117 7361 38151 7395
rect 38485 7361 38519 7395
rect 38853 7361 38887 7395
rect 39221 7361 39255 7395
rect 14381 7293 14415 7327
rect 20545 7293 20579 7327
rect 21833 7293 21867 7327
rect 1593 7225 1627 7259
rect 3065 7225 3099 7259
rect 4445 7225 4479 7259
rect 32689 7225 32723 7259
rect 33701 7225 33735 7259
rect 37657 7225 37691 7259
rect 37933 7225 37967 7259
rect 2145 7157 2179 7191
rect 3341 7157 3375 7191
rect 13369 7157 13403 7191
rect 31033 7157 31067 7191
rect 31309 7157 31343 7191
rect 31585 7157 31619 7191
rect 32137 7157 32171 7191
rect 32413 7157 32447 7191
rect 9873 6953 9907 6987
rect 13737 6953 13771 6987
rect 21281 6953 21315 6987
rect 16497 6885 16531 6919
rect 16589 6885 16623 6919
rect 22385 6885 22419 6919
rect 27721 6885 27755 6919
rect 15117 6817 15151 6851
rect 15485 6817 15519 6851
rect 23489 6817 23523 6851
rect 37749 6817 37783 6851
rect 3433 6749 3467 6783
rect 3801 6749 3835 6783
rect 9137 6749 9171 6783
rect 9230 6749 9264 6783
rect 9643 6749 9677 6783
rect 10057 6749 10091 6783
rect 11989 6749 12023 6783
rect 13921 6749 13955 6783
rect 14841 6749 14875 6783
rect 15761 6749 15795 6783
rect 17325 6749 17359 6783
rect 17601 6749 17635 6783
rect 19993 6749 20027 6783
rect 20269 6749 20303 6783
rect 20545 6749 20579 6783
rect 21373 6749 21407 6783
rect 21649 6749 21683 6783
rect 23213 6749 23247 6783
rect 24869 6749 24903 6783
rect 25329 6749 25363 6783
rect 27353 6749 27387 6783
rect 27629 6749 27663 6783
rect 27905 6749 27939 6783
rect 28181 6749 28215 6783
rect 28457 6749 28491 6783
rect 28733 6749 28767 6783
rect 29009 6749 29043 6783
rect 29285 6749 29319 6783
rect 29745 6749 29779 6783
rect 30021 6749 30055 6783
rect 31953 6749 31987 6783
rect 32229 6749 32263 6783
rect 32413 6749 32447 6783
rect 32689 6749 32723 6783
rect 37841 6749 37875 6783
rect 37933 6749 37967 6783
rect 38485 6749 38519 6783
rect 38853 6749 38887 6783
rect 39221 6749 39255 6783
rect 2881 6681 2915 6715
rect 3065 6681 3099 6715
rect 9413 6681 9447 6715
rect 9505 6681 9539 6715
rect 3617 6613 3651 6647
rect 3985 6613 4019 6647
rect 9781 6613 9815 6647
rect 11805 6613 11839 6647
rect 14105 6613 14139 6647
rect 20177 6613 20211 6647
rect 21281 6613 21315 6647
rect 22477 6613 22511 6647
rect 24685 6613 24719 6647
rect 25145 6613 25179 6647
rect 27169 6613 27203 6647
rect 27445 6613 27479 6647
rect 27997 6613 28031 6647
rect 28273 6613 28307 6647
rect 28549 6613 28583 6647
rect 28825 6613 28859 6647
rect 29101 6613 29135 6647
rect 29561 6613 29595 6647
rect 29837 6613 29871 6647
rect 31769 6613 31803 6647
rect 32045 6613 32079 6647
rect 32597 6613 32631 6647
rect 32873 6613 32907 6647
rect 38117 6613 38151 6647
rect 38669 6613 38703 6647
rect 39037 6613 39071 6647
rect 39405 6613 39439 6647
rect 7573 6409 7607 6443
rect 11805 6409 11839 6443
rect 12817 6409 12851 6443
rect 15945 6409 15979 6443
rect 20453 6409 20487 6443
rect 39405 6409 39439 6443
rect 14841 6341 14875 6375
rect 7389 6273 7423 6307
rect 10057 6273 10091 6307
rect 11621 6273 11655 6307
rect 13001 6273 13035 6307
rect 14473 6273 14507 6307
rect 14566 6273 14600 6307
rect 14749 6273 14783 6307
rect 14979 6273 15013 6307
rect 16129 6273 16163 6307
rect 17417 6273 17451 6307
rect 17693 6273 17727 6307
rect 17969 6273 18003 6307
rect 19165 6273 19199 6307
rect 19717 6273 19751 6307
rect 21281 6273 21315 6307
rect 21833 6273 21867 6307
rect 21926 6273 21960 6307
rect 22109 6273 22143 6307
rect 22201 6273 22235 6307
rect 22339 6273 22373 6307
rect 22845 6273 22879 6307
rect 34989 6273 35023 6307
rect 37749 6273 37783 6307
rect 37933 6273 37967 6307
rect 38853 6273 38887 6307
rect 39221 6273 39255 6307
rect 9781 6205 9815 6239
rect 19441 6205 19475 6239
rect 21557 6205 21591 6239
rect 23121 6205 23155 6239
rect 10241 6137 10275 6171
rect 19349 6137 19383 6171
rect 22477 6137 22511 6171
rect 35173 6137 35207 6171
rect 9873 6069 9907 6103
rect 15117 6069 15151 6103
rect 16681 6069 16715 6103
rect 17785 6069 17819 6103
rect 20545 6069 20579 6103
rect 22661 6069 22695 6103
rect 23029 6069 23063 6103
rect 38117 6069 38151 6103
rect 39037 6069 39071 6103
rect 7665 5865 7699 5899
rect 8953 5865 8987 5899
rect 14841 5865 14875 5899
rect 15945 5865 15979 5899
rect 17049 5865 17083 5899
rect 18521 5865 18555 5899
rect 20545 5865 20579 5899
rect 24041 5865 24075 5899
rect 36093 5865 36127 5899
rect 36921 5865 36955 5899
rect 37749 5865 37783 5899
rect 39405 5865 39439 5899
rect 6745 5797 6779 5831
rect 13369 5797 13403 5831
rect 13829 5797 13863 5831
rect 17141 5797 17175 5831
rect 32229 5797 32263 5831
rect 10333 5729 10367 5763
rect 3801 5661 3835 5695
rect 6561 5661 6595 5695
rect 7481 5661 7515 5695
rect 9137 5661 9171 5695
rect 9781 5661 9815 5695
rect 10149 5661 10183 5695
rect 13185 5661 13219 5695
rect 13645 5661 13679 5695
rect 14381 5661 14415 5695
rect 14473 5661 14507 5695
rect 14657 5661 14691 5695
rect 16129 5661 16163 5695
rect 16865 5661 16899 5695
rect 17325 5661 17359 5695
rect 18705 5661 18739 5695
rect 20361 5661 20395 5695
rect 21097 5661 21131 5695
rect 21251 5661 21285 5695
rect 24225 5661 24259 5695
rect 24593 5661 24627 5695
rect 24869 5661 24903 5695
rect 31953 5661 31987 5695
rect 32045 5661 32079 5695
rect 35909 5661 35943 5695
rect 36737 5661 36771 5695
rect 37841 5661 37875 5695
rect 37933 5661 37967 5695
rect 38853 5661 38887 5695
rect 39221 5661 39255 5695
rect 2973 5593 3007 5627
rect 3157 5593 3191 5627
rect 9965 5593 9999 5627
rect 3985 5525 4019 5559
rect 21465 5525 21499 5559
rect 24409 5525 24443 5559
rect 24685 5525 24719 5559
rect 31861 5525 31895 5559
rect 38117 5525 38151 5559
rect 39037 5525 39071 5559
rect 15485 5321 15519 5355
rect 32321 5321 32355 5355
rect 37657 5321 37691 5355
rect 38117 5321 38151 5355
rect 39405 5321 39439 5355
rect 9413 5253 9447 5287
rect 2973 5185 3007 5219
rect 3341 5185 3375 5219
rect 14013 5185 14047 5219
rect 15301 5185 15335 5219
rect 17049 5185 17083 5219
rect 17693 5185 17727 5219
rect 19809 5185 19843 5219
rect 26801 5185 26835 5219
rect 31493 5185 31527 5219
rect 32137 5185 32171 5219
rect 37473 5185 37507 5219
rect 37933 5185 37967 5219
rect 38853 5185 38887 5219
rect 39221 5185 39255 5219
rect 9597 5117 9631 5151
rect 19533 5117 19567 5151
rect 3525 5049 3559 5083
rect 17509 5049 17543 5083
rect 26617 5049 26651 5083
rect 31677 5049 31711 5083
rect 3065 4981 3099 5015
rect 14197 4981 14231 5015
rect 16865 4981 16899 5015
rect 20545 4981 20579 5015
rect 39037 4981 39071 5015
rect 10793 4777 10827 4811
rect 12265 4777 12299 4811
rect 13369 4777 13403 4811
rect 13553 4777 13587 4811
rect 14289 4777 14323 4811
rect 16221 4777 16255 4811
rect 21741 4777 21775 4811
rect 32045 4777 32079 4811
rect 37933 4777 37967 4811
rect 39405 4777 39439 4811
rect 3157 4641 3191 4675
rect 3433 4573 3467 4607
rect 10977 4573 11011 4607
rect 11253 4573 11287 4607
rect 11437 4573 11471 4607
rect 12081 4573 12115 4607
rect 13737 4573 13771 4607
rect 14105 4573 14139 4607
rect 16405 4573 16439 4607
rect 16681 4573 16715 4607
rect 16865 4573 16899 4607
rect 21925 4573 21959 4607
rect 31493 4573 31527 4607
rect 31585 4573 31619 4607
rect 31861 4573 31895 4607
rect 38117 4573 38151 4607
rect 38853 4573 38887 4607
rect 39221 4573 39255 4607
rect 2973 4505 3007 4539
rect 13277 4505 13311 4539
rect 31217 4505 31251 4539
rect 3617 4437 3651 4471
rect 31125 4437 31159 4471
rect 31401 4437 31435 4471
rect 31769 4437 31803 4471
rect 39037 4437 39071 4471
rect 8677 4233 8711 4267
rect 23857 4233 23891 4267
rect 2513 4165 2547 4199
rect 3249 4165 3283 4199
rect 3617 4165 3651 4199
rect 2881 4097 2915 4131
rect 6377 4097 6411 4131
rect 7297 4097 7331 4131
rect 7414 4097 7448 4131
rect 7573 4097 7607 4131
rect 8585 4097 8619 4131
rect 9873 4097 9907 4131
rect 10148 4097 10182 4131
rect 10241 4097 10275 4131
rect 15209 4097 15243 4131
rect 17866 4097 17900 4131
rect 18025 4097 18059 4131
rect 18153 4097 18187 4131
rect 18245 4097 18279 4131
rect 18383 4097 18417 4131
rect 20269 4097 20303 4131
rect 24041 4097 24075 4131
rect 24310 4097 24344 4131
rect 24501 4097 24535 4131
rect 30665 4097 30699 4131
rect 30757 4097 30791 4131
rect 38853 4097 38887 4131
rect 39221 4097 39255 4131
rect 2697 4029 2731 4063
rect 6561 4029 6595 4063
rect 8217 4029 8251 4063
rect 8493 4029 8527 4063
rect 15301 4029 15335 4063
rect 15485 4029 15519 4063
rect 3065 3961 3099 3995
rect 3801 3961 3835 3995
rect 7021 3961 7055 3995
rect 9045 3961 9079 3995
rect 14841 3961 14875 3995
rect 18521 3961 18555 3995
rect 20453 3961 20487 3995
rect 30941 3961 30975 3995
rect 39405 3961 39439 3995
rect 3341 3893 3375 3927
rect 30573 3893 30607 3927
rect 39037 3893 39071 3927
rect 9229 3689 9263 3723
rect 10701 3689 10735 3723
rect 14197 3689 14231 3723
rect 15393 3689 15427 3723
rect 15945 3689 15979 3723
rect 20729 3689 20763 3723
rect 22293 3689 22327 3723
rect 22385 3689 22419 3723
rect 30113 3689 30147 3723
rect 30665 3689 30699 3723
rect 31401 3689 31435 3723
rect 35541 3689 35575 3723
rect 39405 3689 39439 3723
rect 19717 3621 19751 3655
rect 23581 3621 23615 3655
rect 26157 3621 26191 3655
rect 38117 3621 38151 3655
rect 11345 3553 11379 3587
rect 11504 3553 11538 3587
rect 11621 3553 11655 3587
rect 11897 3553 11931 3587
rect 12357 3553 12391 3587
rect 12541 3553 12575 3587
rect 16589 3553 16623 3587
rect 16748 3553 16782 3587
rect 16865 3553 16899 3587
rect 17141 3553 17175 3587
rect 17785 3553 17819 3587
rect 21281 3553 21315 3587
rect 21741 3553 21775 3587
rect 23029 3553 23063 3587
rect 23188 3553 23222 3587
rect 24041 3553 24075 3587
rect 9137 3485 9171 3519
rect 14289 3485 14323 3519
rect 15484 3485 15518 3519
rect 15577 3485 15611 3519
rect 17601 3485 17635 3519
rect 19533 3485 19567 3519
rect 19625 3485 19659 3519
rect 21097 3485 21131 3519
rect 23305 3485 23339 3519
rect 24225 3485 24259 3519
rect 29929 3485 29963 3519
rect 30481 3485 30515 3519
rect 31217 3485 31251 3519
rect 35449 3485 35483 3519
rect 35725 3485 35759 3519
rect 37657 3485 37691 3519
rect 37841 3485 37875 3519
rect 37933 3485 37967 3519
rect 38393 3485 38427 3519
rect 38485 3485 38519 3519
rect 38945 3485 38979 3519
rect 39221 3485 39255 3519
rect 21189 3417 21223 3451
rect 21925 3417 21959 3451
rect 26341 3417 26375 3451
rect 38761 3417 38795 3451
rect 19349 3349 19383 3383
rect 21833 3349 21867 3383
rect 35357 3349 35391 3383
rect 37473 3349 37507 3383
rect 37749 3349 37783 3383
rect 38209 3349 38243 3383
rect 38669 3349 38703 3383
rect 22477 3145 22511 3179
rect 39037 3145 39071 3179
rect 21557 3077 21591 3111
rect 21465 3009 21499 3043
rect 22691 3009 22725 3043
rect 22845 3009 22879 3043
rect 38485 3009 38519 3043
rect 38853 3009 38887 3043
rect 39221 3009 39255 3043
rect 39405 2873 39439 2907
rect 38669 2805 38703 2839
rect 39405 2601 39439 2635
rect 37565 2533 37599 2567
rect 39037 2533 39071 2567
rect 1685 2397 1719 2431
rect 2053 2397 2087 2431
rect 3617 2397 3651 2431
rect 5181 2397 5215 2431
rect 6745 2397 6779 2431
rect 9597 2397 9631 2431
rect 9873 2397 9907 2431
rect 37381 2397 37415 2431
rect 38025 2397 38059 2431
rect 38117 2397 38151 2431
rect 38485 2397 38519 2431
rect 38853 2397 38887 2431
rect 39221 2397 39255 2431
rect 1869 2261 1903 2295
rect 3433 2261 3467 2295
rect 4997 2261 5031 2295
rect 6561 2261 6595 2295
rect 37841 2261 37875 2295
rect 38301 2261 38335 2295
rect 38669 2261 38703 2295
<< metal1 >>
rect 3878 11160 3884 11212
rect 3936 11200 3942 11212
rect 20070 11200 20076 11212
rect 3936 11172 20076 11200
rect 3936 11160 3942 11172
rect 20070 11160 20076 11172
rect 20128 11160 20134 11212
rect 7834 11092 7840 11144
rect 7892 11132 7898 11144
rect 20898 11132 20904 11144
rect 7892 11104 20904 11132
rect 7892 11092 7898 11104
rect 20898 11092 20904 11104
rect 20956 11092 20962 11144
rect 9766 11024 9772 11076
rect 9824 11064 9830 11076
rect 20622 11064 20628 11076
rect 9824 11036 20628 11064
rect 9824 11024 9830 11036
rect 20622 11024 20628 11036
rect 20680 11024 20686 11076
rect 7190 10072 7196 10124
rect 7248 10112 7254 10124
rect 26786 10112 26792 10124
rect 7248 10084 26792 10112
rect 7248 10072 7254 10084
rect 26786 10072 26792 10084
rect 26844 10072 26850 10124
rect 10594 10004 10600 10056
rect 10652 10044 10658 10056
rect 24118 10044 24124 10056
rect 10652 10016 24124 10044
rect 10652 10004 10658 10016
rect 24118 10004 24124 10016
rect 24176 10004 24182 10056
rect 14642 9936 14648 9988
rect 14700 9976 14706 9988
rect 29914 9976 29920 9988
rect 14700 9948 29920 9976
rect 14700 9936 14706 9948
rect 29914 9936 29920 9948
rect 29972 9936 29978 9988
rect 10870 9868 10876 9920
rect 10928 9908 10934 9920
rect 26602 9908 26608 9920
rect 10928 9880 26608 9908
rect 10928 9868 10934 9880
rect 26602 9868 26608 9880
rect 26660 9868 26666 9920
rect 10042 9800 10048 9852
rect 10100 9840 10106 9852
rect 28534 9840 28540 9852
rect 10100 9812 28540 9840
rect 10100 9800 10106 9812
rect 28534 9800 28540 9812
rect 28592 9800 28598 9852
rect 9490 9732 9496 9784
rect 9548 9772 9554 9784
rect 28718 9772 28724 9784
rect 9548 9744 28724 9772
rect 9548 9732 9554 9744
rect 28718 9732 28724 9744
rect 28776 9732 28782 9784
rect 7742 9664 7748 9716
rect 7800 9704 7806 9716
rect 17126 9704 17132 9716
rect 7800 9676 17132 9704
rect 7800 9664 7806 9676
rect 17126 9664 17132 9676
rect 17184 9664 17190 9716
rect 5810 9596 5816 9648
rect 5868 9636 5874 9648
rect 15562 9636 15568 9648
rect 5868 9608 15568 9636
rect 5868 9596 5874 9608
rect 15562 9596 15568 9608
rect 15620 9596 15626 9648
rect 10318 9528 10324 9580
rect 10376 9568 10382 9580
rect 19334 9568 19340 9580
rect 10376 9540 19340 9568
rect 10376 9528 10382 9540
rect 19334 9528 19340 9540
rect 19392 9528 19398 9580
rect 2682 9460 2688 9512
rect 2740 9500 2746 9512
rect 14458 9500 14464 9512
rect 2740 9472 14464 9500
rect 2740 9460 2746 9472
rect 14458 9460 14464 9472
rect 14516 9460 14522 9512
rect 16666 9460 16672 9512
rect 16724 9500 16730 9512
rect 24394 9500 24400 9512
rect 16724 9472 24400 9500
rect 16724 9460 16730 9472
rect 24394 9460 24400 9472
rect 24452 9460 24458 9512
rect 16022 9392 16028 9444
rect 16080 9432 16086 9444
rect 22094 9432 22100 9444
rect 16080 9404 22100 9432
rect 16080 9392 16086 9404
rect 22094 9392 22100 9404
rect 22152 9392 22158 9444
rect 15470 9324 15476 9376
rect 15528 9364 15534 9376
rect 23474 9364 23480 9376
rect 15528 9336 23480 9364
rect 15528 9324 15534 9336
rect 23474 9324 23480 9336
rect 23532 9324 23538 9376
rect 6914 9256 6920 9308
rect 6972 9296 6978 9308
rect 17494 9296 17500 9308
rect 6972 9268 17500 9296
rect 6972 9256 6978 9268
rect 17494 9256 17500 9268
rect 17552 9256 17558 9308
rect 19058 9256 19064 9308
rect 19116 9296 19122 9308
rect 32582 9296 32588 9308
rect 19116 9268 32588 9296
rect 19116 9256 19122 9268
rect 32582 9256 32588 9268
rect 32640 9256 32646 9308
rect 7558 9188 7564 9240
rect 7616 9228 7622 9240
rect 25222 9228 25228 9240
rect 7616 9200 25228 9228
rect 7616 9188 7622 9200
rect 25222 9188 25228 9200
rect 25280 9188 25286 9240
rect 2130 9120 2136 9172
rect 2188 9160 2194 9172
rect 20438 9160 20444 9172
rect 2188 9132 20444 9160
rect 2188 9120 2194 9132
rect 20438 9120 20444 9132
rect 20496 9120 20502 9172
rect 22646 9120 22652 9172
rect 22704 9160 22710 9172
rect 23842 9160 23848 9172
rect 22704 9132 23848 9160
rect 22704 9120 22710 9132
rect 23842 9120 23848 9132
rect 23900 9120 23906 9172
rect 12434 9092 12440 9104
rect 2746 9064 12440 9092
rect 2038 8984 2044 9036
rect 2096 9024 2102 9036
rect 2746 9024 2774 9064
rect 12434 9052 12440 9064
rect 12492 9052 12498 9104
rect 13814 9052 13820 9104
rect 13872 9092 13878 9104
rect 13872 9064 16712 9092
rect 13872 9052 13878 9064
rect 2096 8996 2774 9024
rect 2096 8984 2102 8996
rect 8386 8984 8392 9036
rect 8444 9024 8450 9036
rect 16574 9024 16580 9036
rect 8444 8996 16580 9024
rect 8444 8984 8450 8996
rect 16574 8984 16580 8996
rect 16632 8984 16638 9036
rect 658 8916 664 8968
rect 716 8956 722 8968
rect 16390 8956 16396 8968
rect 716 8928 16396 8956
rect 716 8916 722 8928
rect 16390 8916 16396 8928
rect 16448 8916 16454 8968
rect 2406 8848 2412 8900
rect 2464 8888 2470 8900
rect 6730 8888 6736 8900
rect 2464 8860 6736 8888
rect 2464 8848 2470 8860
rect 6730 8848 6736 8860
rect 6788 8848 6794 8900
rect 7282 8848 7288 8900
rect 7340 8888 7346 8900
rect 15746 8888 15752 8900
rect 7340 8860 15752 8888
rect 7340 8848 7346 8860
rect 15746 8848 15752 8860
rect 15804 8848 15810 8900
rect 16684 8888 16712 9064
rect 17954 9052 17960 9104
rect 18012 9092 18018 9104
rect 23198 9092 23204 9104
rect 18012 9064 23204 9092
rect 18012 9052 18018 9064
rect 23198 9052 23204 9064
rect 23256 9052 23262 9104
rect 17218 8984 17224 9036
rect 17276 9024 17282 9036
rect 17276 8996 25820 9024
rect 17276 8984 17282 8996
rect 18782 8916 18788 8968
rect 18840 8956 18846 8968
rect 22646 8956 22652 8968
rect 18840 8928 22652 8956
rect 18840 8916 18846 8928
rect 22646 8916 22652 8928
rect 22704 8916 22710 8968
rect 25792 8956 25820 8996
rect 25866 8984 25872 9036
rect 25924 9024 25930 9036
rect 27890 9024 27896 9036
rect 25924 8996 27896 9024
rect 25924 8984 25930 8996
rect 27890 8984 27896 8996
rect 27948 8984 27954 9036
rect 30466 8956 30472 8968
rect 25792 8928 30472 8956
rect 30466 8916 30472 8928
rect 30524 8916 30530 8968
rect 30650 8916 30656 8968
rect 30708 8956 30714 8968
rect 33778 8956 33784 8968
rect 30708 8928 33784 8956
rect 30708 8916 30714 8928
rect 33778 8916 33784 8928
rect 33836 8916 33842 8968
rect 25498 8888 25504 8900
rect 16684 8860 25504 8888
rect 25498 8848 25504 8860
rect 25556 8848 25562 8900
rect 32398 8848 32404 8900
rect 32456 8888 32462 8900
rect 35066 8888 35072 8900
rect 32456 8860 35072 8888
rect 32456 8848 32462 8860
rect 35066 8848 35072 8860
rect 35124 8848 35130 8900
rect 1578 8780 1584 8832
rect 1636 8820 1642 8832
rect 8570 8820 8576 8832
rect 1636 8792 8576 8820
rect 1636 8780 1642 8792
rect 8570 8780 8576 8792
rect 8628 8780 8634 8832
rect 12526 8780 12532 8832
rect 12584 8820 12590 8832
rect 14734 8820 14740 8832
rect 12584 8792 14740 8820
rect 12584 8780 12590 8792
rect 14734 8780 14740 8792
rect 14792 8780 14798 8832
rect 19702 8780 19708 8832
rect 19760 8820 19766 8832
rect 23750 8820 23756 8832
rect 19760 8792 23756 8820
rect 19760 8780 19766 8792
rect 23750 8780 23756 8792
rect 23808 8780 23814 8832
rect 26142 8780 26148 8832
rect 26200 8820 26206 8832
rect 28442 8820 28448 8832
rect 26200 8792 28448 8820
rect 26200 8780 26206 8792
rect 28442 8780 28448 8792
rect 28500 8780 28506 8832
rect 33042 8780 33048 8832
rect 33100 8820 33106 8832
rect 33502 8820 33508 8832
rect 33100 8792 33508 8820
rect 33100 8780 33106 8792
rect 33502 8780 33508 8792
rect 33560 8780 33566 8832
rect 34974 8780 34980 8832
rect 35032 8820 35038 8832
rect 35618 8820 35624 8832
rect 35032 8792 35624 8820
rect 35032 8780 35038 8792
rect 35618 8780 35624 8792
rect 35676 8780 35682 8832
rect 1104 8730 39836 8752
rect 1104 8678 3010 8730
rect 3062 8678 3074 8730
rect 3126 8678 3138 8730
rect 3190 8678 3202 8730
rect 3254 8678 3266 8730
rect 3318 8678 9010 8730
rect 9062 8678 9074 8730
rect 9126 8678 9138 8730
rect 9190 8678 9202 8730
rect 9254 8678 9266 8730
rect 9318 8678 15010 8730
rect 15062 8678 15074 8730
rect 15126 8678 15138 8730
rect 15190 8678 15202 8730
rect 15254 8678 15266 8730
rect 15318 8678 21010 8730
rect 21062 8678 21074 8730
rect 21126 8678 21138 8730
rect 21190 8678 21202 8730
rect 21254 8678 21266 8730
rect 21318 8678 27010 8730
rect 27062 8678 27074 8730
rect 27126 8678 27138 8730
rect 27190 8678 27202 8730
rect 27254 8678 27266 8730
rect 27318 8678 33010 8730
rect 33062 8678 33074 8730
rect 33126 8678 33138 8730
rect 33190 8678 33202 8730
rect 33254 8678 33266 8730
rect 33318 8678 39010 8730
rect 39062 8678 39074 8730
rect 39126 8678 39138 8730
rect 39190 8678 39202 8730
rect 39254 8678 39266 8730
rect 39318 8678 39836 8730
rect 1104 8656 39836 8678
rect 1118 8576 1124 8628
rect 1176 8616 1182 8628
rect 1176 8588 2268 8616
rect 1176 8576 1182 8588
rect 1302 8508 1308 8560
rect 1360 8548 1366 8560
rect 1360 8520 2084 8548
rect 1360 8508 1366 8520
rect 566 8440 572 8492
rect 624 8480 630 8492
rect 1397 8483 1455 8489
rect 1397 8480 1409 8483
rect 624 8452 1409 8480
rect 624 8440 630 8452
rect 1397 8449 1409 8452
rect 1443 8449 1455 8483
rect 1397 8443 1455 8449
rect 1673 8483 1731 8489
rect 1673 8449 1685 8483
rect 1719 8449 1731 8483
rect 1673 8443 1731 8449
rect 1949 8483 2007 8489
rect 1949 8449 1961 8483
rect 1995 8449 2007 8483
rect 1949 8443 2007 8449
rect 842 8372 848 8424
rect 900 8412 906 8424
rect 1688 8412 1716 8443
rect 900 8384 1716 8412
rect 900 8372 906 8384
rect 1026 8304 1032 8356
rect 1084 8344 1090 8356
rect 1964 8344 1992 8443
rect 2056 8412 2084 8520
rect 2240 8489 2268 8588
rect 2406 8576 2412 8628
rect 2464 8576 2470 8628
rect 2682 8576 2688 8628
rect 2740 8576 2746 8628
rect 3421 8619 3479 8625
rect 3421 8585 3433 8619
rect 3467 8616 3479 8619
rect 3786 8616 3792 8628
rect 3467 8588 3792 8616
rect 3467 8585 3479 8588
rect 3421 8579 3479 8585
rect 3786 8576 3792 8588
rect 3844 8576 3850 8628
rect 4249 8619 4307 8625
rect 4249 8585 4261 8619
rect 4295 8616 4307 8619
rect 4338 8616 4344 8628
rect 4295 8588 4344 8616
rect 4295 8585 4307 8588
rect 4249 8579 4307 8585
rect 4338 8576 4344 8588
rect 4396 8576 4402 8628
rect 4614 8576 4620 8628
rect 4672 8576 4678 8628
rect 4985 8619 5043 8625
rect 4985 8585 4997 8619
rect 5031 8616 5043 8619
rect 5166 8616 5172 8628
rect 5031 8588 5172 8616
rect 5031 8585 5043 8588
rect 4985 8579 5043 8585
rect 5166 8576 5172 8588
rect 5224 8576 5230 8628
rect 5261 8619 5319 8625
rect 5261 8585 5273 8619
rect 5307 8616 5319 8619
rect 5442 8616 5448 8628
rect 5307 8588 5448 8616
rect 5307 8585 5319 8588
rect 5261 8579 5319 8585
rect 5442 8576 5448 8588
rect 5500 8576 5506 8628
rect 5629 8619 5687 8625
rect 5629 8585 5641 8619
rect 5675 8616 5687 8619
rect 5718 8616 5724 8628
rect 5675 8588 5724 8616
rect 5675 8585 5687 8588
rect 5629 8579 5687 8585
rect 5718 8576 5724 8588
rect 5776 8576 5782 8628
rect 5997 8619 6055 8625
rect 5997 8585 6009 8619
rect 6043 8616 6055 8619
rect 6270 8616 6276 8628
rect 6043 8588 6276 8616
rect 6043 8585 6055 8588
rect 5997 8579 6055 8585
rect 6270 8576 6276 8588
rect 6328 8576 6334 8628
rect 6733 8619 6791 8625
rect 6733 8585 6745 8619
rect 6779 8616 6791 8619
rect 6822 8616 6828 8628
rect 6779 8588 6828 8616
rect 6779 8585 6791 8588
rect 6733 8579 6791 8585
rect 6822 8576 6828 8588
rect 6880 8576 6886 8628
rect 7101 8619 7159 8625
rect 7101 8585 7113 8619
rect 7147 8616 7159 8619
rect 7374 8616 7380 8628
rect 7147 8588 7380 8616
rect 7147 8585 7159 8588
rect 7101 8579 7159 8585
rect 7374 8576 7380 8588
rect 7432 8576 7438 8628
rect 7469 8619 7527 8625
rect 7469 8585 7481 8619
rect 7515 8616 7527 8619
rect 7650 8616 7656 8628
rect 7515 8588 7656 8616
rect 7515 8585 7527 8588
rect 7469 8579 7527 8585
rect 7650 8576 7656 8588
rect 7708 8576 7714 8628
rect 7837 8619 7895 8625
rect 7837 8585 7849 8619
rect 7883 8616 7895 8619
rect 7926 8616 7932 8628
rect 7883 8588 7932 8616
rect 7883 8585 7895 8588
rect 7837 8579 7895 8585
rect 7926 8576 7932 8588
rect 7984 8576 7990 8628
rect 8205 8619 8263 8625
rect 8205 8585 8217 8619
rect 8251 8616 8263 8619
rect 8478 8616 8484 8628
rect 8251 8588 8484 8616
rect 8251 8585 8263 8588
rect 8205 8579 8263 8585
rect 8478 8576 8484 8588
rect 8536 8576 8542 8628
rect 8573 8619 8631 8625
rect 8573 8585 8585 8619
rect 8619 8616 8631 8619
rect 8846 8616 8852 8628
rect 8619 8588 8852 8616
rect 8619 8585 8631 8588
rect 8573 8579 8631 8585
rect 8846 8576 8852 8588
rect 8904 8576 8910 8628
rect 9309 8619 9367 8625
rect 9309 8585 9321 8619
rect 9355 8616 9367 8619
rect 9582 8616 9588 8628
rect 9355 8588 9588 8616
rect 9355 8585 9367 8588
rect 9309 8579 9367 8585
rect 9582 8576 9588 8588
rect 9640 8576 9646 8628
rect 9677 8619 9735 8625
rect 9677 8585 9689 8619
rect 9723 8616 9735 8619
rect 9858 8616 9864 8628
rect 9723 8588 9864 8616
rect 9723 8585 9735 8588
rect 9677 8579 9735 8585
rect 9858 8576 9864 8588
rect 9916 8576 9922 8628
rect 10045 8619 10103 8625
rect 10045 8585 10057 8619
rect 10091 8616 10103 8619
rect 10134 8616 10140 8628
rect 10091 8588 10140 8616
rect 10091 8585 10103 8588
rect 10045 8579 10103 8585
rect 10134 8576 10140 8588
rect 10192 8576 10198 8628
rect 10413 8619 10471 8625
rect 10413 8585 10425 8619
rect 10459 8616 10471 8619
rect 10686 8616 10692 8628
rect 10459 8588 10692 8616
rect 10459 8585 10471 8588
rect 10413 8579 10471 8585
rect 10686 8576 10692 8588
rect 10744 8576 10750 8628
rect 10781 8619 10839 8625
rect 10781 8585 10793 8619
rect 10827 8616 10839 8619
rect 10962 8616 10968 8628
rect 10827 8588 10968 8616
rect 10827 8585 10839 8588
rect 10781 8579 10839 8585
rect 10962 8576 10968 8588
rect 11020 8576 11026 8628
rect 11241 8619 11299 8625
rect 11241 8585 11253 8619
rect 11287 8616 11299 8619
rect 11514 8616 11520 8628
rect 11287 8588 11520 8616
rect 11287 8585 11299 8588
rect 11241 8579 11299 8585
rect 11514 8576 11520 8588
rect 11572 8576 11578 8628
rect 11701 8619 11759 8625
rect 11701 8585 11713 8619
rect 11747 8616 11759 8619
rect 11974 8616 11980 8628
rect 11747 8588 11980 8616
rect 11747 8585 11759 8588
rect 11701 8579 11759 8585
rect 11974 8576 11980 8588
rect 12032 8576 12038 8628
rect 12069 8619 12127 8625
rect 12069 8585 12081 8619
rect 12115 8616 12127 8619
rect 12342 8616 12348 8628
rect 12115 8588 12348 8616
rect 12115 8585 12127 8588
rect 12069 8579 12127 8585
rect 12342 8576 12348 8588
rect 12400 8576 12406 8628
rect 12805 8619 12863 8625
rect 12805 8585 12817 8619
rect 12851 8616 12863 8619
rect 13170 8616 13176 8628
rect 12851 8588 13176 8616
rect 12851 8585 12863 8588
rect 12805 8579 12863 8585
rect 13170 8576 13176 8588
rect 13228 8576 13234 8628
rect 13817 8619 13875 8625
rect 13817 8585 13829 8619
rect 13863 8616 13875 8619
rect 13998 8616 14004 8628
rect 13863 8588 14004 8616
rect 13863 8585 13875 8588
rect 13817 8579 13875 8585
rect 13998 8576 14004 8588
rect 14056 8576 14062 8628
rect 14461 8619 14519 8625
rect 14461 8585 14473 8619
rect 14507 8616 14519 8619
rect 14550 8616 14556 8628
rect 14507 8588 14556 8616
rect 14507 8585 14519 8588
rect 14461 8579 14519 8585
rect 14550 8576 14556 8588
rect 14608 8576 14614 8628
rect 14829 8619 14887 8625
rect 14829 8585 14841 8619
rect 14875 8616 14887 8619
rect 14918 8616 14924 8628
rect 14875 8588 14924 8616
rect 14875 8585 14887 8588
rect 14829 8579 14887 8585
rect 14918 8576 14924 8588
rect 14976 8576 14982 8628
rect 15197 8619 15255 8625
rect 15197 8585 15209 8619
rect 15243 8616 15255 8619
rect 15378 8616 15384 8628
rect 15243 8588 15384 8616
rect 15243 8585 15255 8588
rect 15197 8579 15255 8585
rect 15378 8576 15384 8588
rect 15436 8576 15442 8628
rect 15654 8576 15660 8628
rect 15712 8576 15718 8628
rect 15933 8619 15991 8625
rect 15933 8585 15945 8619
rect 15979 8616 15991 8619
rect 16206 8616 16212 8628
rect 15979 8588 16212 8616
rect 15979 8585 15991 8588
rect 15933 8579 15991 8585
rect 16206 8576 16212 8588
rect 16264 8576 16270 8628
rect 16301 8619 16359 8625
rect 16301 8585 16313 8619
rect 16347 8616 16359 8619
rect 16482 8616 16488 8628
rect 16347 8588 16488 8616
rect 16347 8585 16359 8588
rect 16301 8579 16359 8585
rect 16482 8576 16488 8588
rect 16540 8576 16546 8628
rect 16758 8576 16764 8628
rect 16816 8616 16822 8628
rect 17037 8619 17095 8625
rect 17037 8616 17049 8619
rect 16816 8588 17049 8616
rect 16816 8576 16822 8588
rect 17037 8585 17049 8588
rect 17083 8585 17095 8619
rect 17037 8579 17095 8585
rect 17310 8576 17316 8628
rect 17368 8616 17374 8628
rect 17589 8619 17647 8625
rect 17589 8616 17601 8619
rect 17368 8588 17601 8616
rect 17368 8576 17374 8588
rect 17589 8585 17601 8588
rect 17635 8585 17647 8619
rect 17589 8579 17647 8585
rect 18782 8576 18788 8628
rect 18840 8576 18846 8628
rect 19334 8576 19340 8628
rect 19392 8576 19398 8628
rect 19518 8576 19524 8628
rect 19576 8576 19582 8628
rect 19610 8576 19616 8628
rect 19668 8576 19674 8628
rect 20530 8576 20536 8628
rect 20588 8616 20594 8628
rect 21821 8619 21879 8625
rect 21821 8616 21833 8619
rect 20588 8588 21833 8616
rect 20588 8576 20594 8588
rect 21821 8585 21833 8588
rect 21867 8585 21879 8619
rect 21821 8579 21879 8585
rect 22002 8576 22008 8628
rect 22060 8616 22066 8628
rect 22060 8588 22416 8616
rect 22060 8576 22066 8588
rect 7742 8548 7748 8560
rect 3252 8520 7748 8548
rect 3252 8489 3280 8520
rect 7742 8508 7748 8520
rect 7800 8508 7806 8560
rect 11606 8548 11612 8560
rect 7944 8520 11612 8548
rect 2225 8483 2283 8489
rect 2225 8449 2237 8483
rect 2271 8449 2283 8483
rect 2225 8443 2283 8449
rect 2501 8483 2559 8489
rect 2501 8449 2513 8483
rect 2547 8449 2559 8483
rect 2501 8443 2559 8449
rect 3237 8483 3295 8489
rect 3237 8449 3249 8483
rect 3283 8449 3295 8483
rect 3237 8443 3295 8449
rect 3605 8483 3663 8489
rect 3605 8449 3617 8483
rect 3651 8449 3663 8483
rect 3605 8443 3663 8449
rect 2516 8412 2544 8443
rect 2056 8384 2544 8412
rect 1084 8316 1992 8344
rect 1084 8304 1090 8316
rect 2038 8304 2044 8356
rect 2096 8304 2102 8356
rect 2130 8304 2136 8356
rect 2188 8304 2194 8356
rect 3053 8347 3111 8353
rect 3053 8313 3065 8347
rect 3099 8344 3111 8347
rect 3510 8344 3516 8356
rect 3099 8316 3516 8344
rect 3099 8313 3111 8316
rect 3053 8307 3111 8313
rect 3510 8304 3516 8316
rect 3568 8304 3574 8356
rect 3620 8344 3648 8443
rect 3694 8440 3700 8492
rect 3752 8480 3758 8492
rect 4065 8483 4123 8489
rect 4065 8480 4077 8483
rect 3752 8452 4077 8480
rect 3752 8440 3758 8452
rect 4065 8449 4077 8452
rect 4111 8449 4123 8483
rect 4065 8443 4123 8449
rect 4433 8483 4491 8489
rect 4433 8449 4445 8483
rect 4479 8449 4491 8483
rect 4433 8443 4491 8449
rect 3970 8372 3976 8424
rect 4028 8412 4034 8424
rect 4448 8412 4476 8443
rect 4522 8440 4528 8492
rect 4580 8480 4586 8492
rect 4801 8483 4859 8489
rect 4801 8480 4813 8483
rect 4580 8452 4813 8480
rect 4580 8440 4586 8452
rect 4801 8449 4813 8452
rect 4847 8449 4859 8483
rect 4801 8443 4859 8449
rect 5445 8483 5503 8489
rect 5445 8449 5457 8483
rect 5491 8480 5503 8483
rect 5626 8480 5632 8492
rect 5491 8452 5632 8480
rect 5491 8449 5503 8452
rect 5445 8443 5503 8449
rect 5626 8440 5632 8452
rect 5684 8440 5690 8492
rect 5810 8440 5816 8492
rect 5868 8440 5874 8492
rect 6181 8483 6239 8489
rect 6181 8449 6193 8483
rect 6227 8449 6239 8483
rect 6181 8443 6239 8449
rect 4028 8384 4476 8412
rect 6196 8412 6224 8443
rect 6914 8440 6920 8492
rect 6972 8440 6978 8492
rect 7282 8440 7288 8492
rect 7340 8440 7346 8492
rect 7650 8440 7656 8492
rect 7708 8440 7714 8492
rect 7006 8412 7012 8424
rect 6196 8384 7012 8412
rect 4028 8372 4034 8384
rect 7006 8372 7012 8384
rect 7064 8372 7070 8424
rect 7944 8344 7972 8520
rect 11606 8508 11612 8520
rect 11664 8508 11670 8560
rect 12526 8548 12532 8560
rect 11900 8520 12532 8548
rect 8021 8483 8079 8489
rect 8021 8449 8033 8483
rect 8067 8449 8079 8483
rect 8021 8443 8079 8449
rect 3620 8316 7972 8344
rect 8036 8344 8064 8443
rect 8386 8440 8392 8492
rect 8444 8440 8450 8492
rect 8662 8440 8668 8492
rect 8720 8480 8726 8492
rect 8757 8483 8815 8489
rect 8757 8480 8769 8483
rect 8720 8452 8769 8480
rect 8720 8440 8726 8452
rect 8757 8449 8769 8452
rect 8803 8449 8815 8483
rect 8757 8443 8815 8449
rect 9490 8440 9496 8492
rect 9548 8440 9554 8492
rect 9861 8483 9919 8489
rect 9861 8449 9873 8483
rect 9907 8480 9919 8483
rect 10042 8480 10048 8492
rect 9907 8452 10048 8480
rect 9907 8449 9919 8452
rect 9861 8443 9919 8449
rect 10042 8440 10048 8452
rect 10100 8440 10106 8492
rect 10226 8440 10232 8492
rect 10284 8440 10290 8492
rect 10594 8440 10600 8492
rect 10652 8440 10658 8492
rect 10870 8440 10876 8492
rect 10928 8480 10934 8492
rect 11900 8489 11928 8520
rect 12526 8508 12532 8520
rect 12584 8508 12590 8560
rect 14734 8548 14740 8560
rect 12636 8520 14740 8548
rect 12636 8489 12664 8520
rect 14734 8508 14740 8520
rect 14792 8508 14798 8560
rect 17218 8548 17224 8560
rect 15021 8520 17224 8548
rect 10965 8483 11023 8489
rect 10965 8480 10977 8483
rect 10928 8452 10977 8480
rect 10928 8440 10934 8452
rect 10965 8449 10977 8452
rect 11011 8449 11023 8483
rect 10965 8443 11023 8449
rect 11057 8483 11115 8489
rect 11057 8449 11069 8483
rect 11103 8449 11115 8483
rect 11057 8443 11115 8449
rect 11885 8483 11943 8489
rect 11885 8449 11897 8483
rect 11931 8449 11943 8483
rect 11885 8443 11943 8449
rect 12253 8483 12311 8489
rect 12253 8449 12265 8483
rect 12299 8480 12311 8483
rect 12621 8483 12679 8489
rect 12299 8452 12572 8480
rect 12299 8449 12311 8452
rect 12253 8443 12311 8449
rect 8478 8372 8484 8424
rect 8536 8412 8542 8424
rect 11072 8412 11100 8443
rect 8536 8384 11100 8412
rect 12544 8412 12572 8452
rect 12621 8449 12633 8483
rect 12667 8449 12679 8483
rect 12621 8443 12679 8449
rect 12986 8440 12992 8492
rect 13044 8440 13050 8492
rect 13354 8440 13360 8492
rect 13412 8440 13418 8492
rect 13449 8483 13507 8489
rect 13449 8449 13461 8483
rect 13495 8480 13507 8483
rect 13633 8483 13691 8489
rect 13633 8480 13645 8483
rect 13495 8452 13645 8480
rect 13495 8449 13507 8452
rect 13449 8443 13507 8449
rect 13633 8449 13645 8452
rect 13679 8449 13691 8483
rect 13633 8443 13691 8449
rect 13538 8412 13544 8424
rect 12544 8384 13544 8412
rect 8536 8372 8542 8384
rect 13538 8372 13544 8384
rect 13596 8372 13602 8424
rect 13648 8412 13676 8443
rect 14642 8440 14648 8492
rect 14700 8440 14706 8492
rect 15021 8489 15049 8520
rect 17218 8508 17224 8520
rect 17276 8508 17282 8560
rect 19536 8548 19564 8576
rect 19536 8520 19840 8548
rect 15013 8483 15071 8489
rect 15013 8449 15025 8483
rect 15059 8449 15071 8483
rect 15013 8443 15071 8449
rect 15378 8440 15384 8492
rect 15436 8440 15442 8492
rect 15473 8483 15531 8489
rect 15473 8449 15485 8483
rect 15519 8480 15531 8483
rect 15838 8480 15844 8492
rect 15519 8452 15844 8480
rect 15519 8449 15531 8452
rect 15473 8443 15531 8449
rect 15838 8440 15844 8452
rect 15896 8440 15902 8492
rect 16114 8440 16120 8492
rect 16172 8440 16178 8492
rect 16485 8483 16543 8489
rect 16485 8449 16497 8483
rect 16531 8480 16543 8483
rect 16666 8480 16672 8492
rect 16531 8452 16672 8480
rect 16531 8449 16543 8452
rect 16485 8443 16543 8449
rect 16666 8440 16672 8452
rect 16724 8440 16730 8492
rect 16850 8440 16856 8492
rect 16908 8440 16914 8492
rect 17402 8440 17408 8492
rect 17460 8440 17466 8492
rect 17773 8483 17831 8489
rect 17773 8449 17785 8483
rect 17819 8480 17831 8483
rect 18046 8480 18052 8492
rect 17819 8452 18052 8480
rect 17819 8449 17831 8452
rect 17773 8443 17831 8449
rect 18046 8440 18052 8452
rect 18104 8440 18110 8492
rect 18414 8440 18420 8492
rect 18472 8480 18478 8492
rect 18509 8483 18567 8489
rect 18509 8480 18521 8483
rect 18472 8452 18521 8480
rect 18472 8440 18478 8452
rect 18509 8449 18521 8452
rect 18555 8449 18567 8483
rect 18509 8443 18567 8449
rect 18601 8483 18659 8489
rect 18601 8449 18613 8483
rect 18647 8480 18659 8483
rect 18690 8480 18696 8492
rect 18647 8452 18696 8480
rect 18647 8449 18659 8452
rect 18601 8443 18659 8449
rect 18690 8440 18696 8452
rect 18748 8440 18754 8492
rect 18877 8483 18935 8489
rect 18877 8449 18889 8483
rect 18923 8480 18935 8483
rect 18966 8480 18972 8492
rect 18923 8452 18972 8480
rect 18923 8449 18935 8452
rect 18877 8443 18935 8449
rect 18966 8440 18972 8452
rect 19024 8440 19030 8492
rect 19242 8440 19248 8492
rect 19300 8480 19306 8492
rect 19812 8489 19840 8520
rect 21726 8508 21732 8560
rect 21784 8548 21790 8560
rect 21784 8520 22324 8548
rect 21784 8508 21790 8520
rect 19521 8483 19579 8489
rect 19521 8480 19533 8483
rect 19300 8452 19533 8480
rect 19300 8440 19306 8452
rect 19521 8449 19533 8452
rect 19567 8449 19579 8483
rect 19521 8443 19579 8449
rect 19797 8483 19855 8489
rect 19797 8449 19809 8483
rect 19843 8449 19855 8483
rect 19797 8443 19855 8449
rect 19886 8440 19892 8492
rect 19944 8440 19950 8492
rect 21358 8440 21364 8492
rect 21416 8480 21422 8492
rect 21453 8483 21511 8489
rect 21453 8480 21465 8483
rect 21416 8452 21465 8480
rect 21416 8440 21422 8452
rect 21453 8449 21465 8452
rect 21499 8449 21511 8483
rect 21453 8443 21511 8449
rect 21542 8440 21548 8492
rect 21600 8480 21606 8492
rect 22296 8489 22324 8520
rect 22388 8489 22416 8588
rect 23106 8576 23112 8628
rect 23164 8616 23170 8628
rect 23164 8588 23520 8616
rect 23164 8576 23170 8588
rect 22554 8508 22560 8560
rect 22612 8548 22618 8560
rect 22612 8520 23152 8548
rect 22612 8508 22618 8520
rect 22005 8483 22063 8489
rect 22005 8480 22017 8483
rect 21600 8452 22017 8480
rect 21600 8440 21606 8452
rect 22005 8449 22017 8452
rect 22051 8449 22063 8483
rect 22005 8443 22063 8449
rect 22281 8483 22339 8489
rect 22281 8449 22293 8483
rect 22327 8449 22339 8483
rect 22281 8443 22339 8449
rect 22373 8483 22431 8489
rect 22373 8449 22385 8483
rect 22419 8449 22431 8483
rect 22373 8443 22431 8449
rect 22462 8440 22468 8492
rect 22520 8480 22526 8492
rect 23124 8489 23152 8520
rect 23492 8489 23520 8588
rect 23750 8576 23756 8628
rect 23808 8576 23814 8628
rect 23934 8576 23940 8628
rect 23992 8616 23998 8628
rect 23992 8588 24624 8616
rect 23992 8576 23998 8588
rect 23658 8508 23664 8560
rect 23716 8548 23722 8560
rect 23716 8520 24256 8548
rect 23716 8508 23722 8520
rect 24228 8489 24256 8520
rect 24596 8489 24624 8588
rect 24762 8576 24768 8628
rect 24820 8616 24826 8628
rect 24820 8588 25268 8616
rect 24820 8576 24826 8588
rect 24670 8508 24676 8560
rect 24728 8548 24734 8560
rect 24728 8520 25176 8548
rect 24728 8508 24734 8520
rect 25148 8489 25176 8520
rect 22833 8483 22891 8489
rect 22833 8480 22845 8483
rect 22520 8452 22845 8480
rect 22520 8440 22526 8452
rect 22833 8449 22845 8452
rect 22879 8449 22891 8483
rect 22833 8443 22891 8449
rect 23109 8483 23167 8489
rect 23109 8449 23121 8483
rect 23155 8449 23167 8483
rect 23109 8443 23167 8449
rect 23385 8483 23443 8489
rect 23385 8449 23397 8483
rect 23431 8449 23443 8483
rect 23385 8443 23443 8449
rect 23477 8483 23535 8489
rect 23477 8449 23489 8483
rect 23523 8449 23535 8483
rect 23477 8443 23535 8449
rect 23937 8483 23995 8489
rect 23937 8449 23949 8483
rect 23983 8449 23995 8483
rect 23937 8443 23995 8449
rect 24213 8483 24271 8489
rect 24213 8449 24225 8483
rect 24259 8449 24271 8483
rect 24213 8443 24271 8449
rect 24581 8483 24639 8489
rect 24581 8449 24593 8483
rect 24627 8449 24639 8483
rect 24581 8443 24639 8449
rect 24857 8483 24915 8489
rect 24857 8449 24869 8483
rect 24903 8449 24915 8483
rect 24857 8443 24915 8449
rect 25133 8483 25191 8489
rect 25133 8449 25145 8483
rect 25179 8449 25191 8483
rect 25240 8480 25268 8588
rect 25498 8576 25504 8628
rect 25556 8576 25562 8628
rect 25682 8576 25688 8628
rect 25740 8616 25746 8628
rect 30469 8619 30527 8625
rect 30469 8616 30481 8619
rect 25740 8588 30481 8616
rect 25740 8576 25746 8588
rect 30469 8585 30481 8588
rect 30515 8585 30527 8619
rect 30469 8579 30527 8585
rect 32214 8576 32220 8628
rect 32272 8616 32278 8628
rect 32309 8619 32367 8625
rect 32309 8616 32321 8619
rect 32272 8588 32321 8616
rect 32272 8576 32278 8588
rect 32309 8585 32321 8588
rect 32355 8585 32367 8619
rect 32309 8579 32367 8585
rect 32490 8576 32496 8628
rect 32548 8616 32554 8628
rect 32769 8619 32827 8625
rect 32769 8616 32781 8619
rect 32548 8588 32781 8616
rect 32548 8576 32554 8588
rect 32769 8585 32781 8588
rect 32815 8585 32827 8619
rect 32769 8579 32827 8585
rect 32858 8576 32864 8628
rect 32916 8616 32922 8628
rect 33137 8619 33195 8625
rect 33137 8616 33149 8619
rect 32916 8588 33149 8616
rect 32916 8576 32922 8588
rect 33137 8585 33149 8588
rect 33183 8585 33195 8619
rect 33137 8579 33195 8585
rect 33502 8576 33508 8628
rect 33560 8576 33566 8628
rect 33594 8576 33600 8628
rect 33652 8616 33658 8628
rect 34241 8619 34299 8625
rect 34241 8616 34253 8619
rect 33652 8588 34253 8616
rect 33652 8576 33658 8588
rect 34241 8585 34253 8588
rect 34287 8585 34299 8619
rect 34241 8579 34299 8585
rect 34698 8576 34704 8628
rect 34756 8616 34762 8628
rect 35529 8619 35587 8625
rect 35529 8616 35541 8619
rect 34756 8588 35541 8616
rect 34756 8576 34762 8588
rect 35529 8585 35541 8588
rect 35575 8585 35587 8619
rect 35529 8579 35587 8585
rect 35802 8576 35808 8628
rect 35860 8616 35866 8628
rect 36725 8619 36783 8625
rect 36725 8616 36737 8619
rect 35860 8588 36737 8616
rect 35860 8576 35866 8588
rect 36725 8585 36737 8588
rect 36771 8585 36783 8619
rect 36725 8579 36783 8585
rect 36906 8576 36912 8628
rect 36964 8616 36970 8628
rect 37829 8619 37887 8625
rect 37829 8616 37841 8619
rect 36964 8588 37841 8616
rect 36964 8576 36970 8588
rect 37829 8585 37841 8588
rect 37875 8585 37887 8619
rect 37829 8579 37887 8585
rect 38565 8619 38623 8625
rect 38565 8585 38577 8619
rect 38611 8585 38623 8619
rect 38565 8579 38623 8585
rect 25314 8508 25320 8560
rect 25372 8548 25378 8560
rect 25372 8520 25820 8548
rect 25372 8508 25378 8520
rect 25792 8489 25820 8520
rect 26510 8508 26516 8560
rect 26568 8548 26574 8560
rect 26568 8520 29684 8548
rect 26568 8508 26574 8520
rect 25409 8483 25467 8489
rect 25409 8480 25421 8483
rect 25240 8452 25421 8480
rect 25133 8443 25191 8449
rect 25409 8449 25421 8452
rect 25455 8449 25467 8483
rect 25409 8443 25467 8449
rect 25685 8483 25743 8489
rect 25685 8449 25697 8483
rect 25731 8449 25743 8483
rect 25685 8443 25743 8449
rect 25777 8483 25835 8489
rect 25777 8449 25789 8483
rect 25823 8449 25835 8483
rect 25777 8443 25835 8449
rect 15102 8412 15108 8424
rect 13648 8384 15108 8412
rect 15102 8372 15108 8384
rect 15160 8372 15166 8424
rect 17678 8372 17684 8424
rect 17736 8412 17742 8424
rect 17736 8384 18368 8412
rect 17736 8372 17742 8384
rect 11974 8344 11980 8356
rect 8036 8316 11980 8344
rect 11974 8304 11980 8316
rect 12032 8304 12038 8356
rect 12437 8347 12495 8353
rect 12437 8313 12449 8347
rect 12483 8344 12495 8347
rect 12894 8344 12900 8356
rect 12483 8316 12900 8344
rect 12483 8313 12495 8316
rect 12437 8307 12495 8313
rect 12894 8304 12900 8316
rect 12952 8304 12958 8356
rect 13173 8347 13231 8353
rect 13173 8313 13185 8347
rect 13219 8344 13231 8347
rect 13722 8344 13728 8356
rect 13219 8316 13728 8344
rect 13219 8313 13231 8316
rect 13173 8307 13231 8313
rect 13722 8304 13728 8316
rect 13780 8304 13786 8356
rect 17034 8304 17040 8356
rect 17092 8344 17098 8356
rect 18340 8353 18368 8384
rect 20088 8384 22508 8412
rect 17957 8347 18015 8353
rect 17957 8344 17969 8347
rect 17092 8316 17969 8344
rect 17092 8304 17098 8316
rect 17957 8313 17969 8316
rect 18003 8313 18015 8347
rect 17957 8307 18015 8313
rect 18325 8347 18383 8353
rect 18325 8313 18337 8347
rect 18371 8313 18383 8347
rect 18325 8307 18383 8313
rect 19061 8347 19119 8353
rect 19061 8313 19073 8347
rect 19107 8344 19119 8347
rect 19794 8344 19800 8356
rect 19107 8316 19800 8344
rect 19107 8313 19119 8316
rect 19061 8307 19119 8313
rect 19794 8304 19800 8316
rect 19852 8304 19858 8356
rect 20088 8353 20116 8384
rect 22480 8356 22508 8384
rect 22572 8384 22876 8412
rect 20073 8347 20131 8353
rect 20073 8313 20085 8347
rect 20119 8313 20131 8347
rect 20073 8307 20131 8313
rect 21269 8347 21327 8353
rect 21269 8313 21281 8347
rect 21315 8344 21327 8347
rect 21634 8344 21640 8356
rect 21315 8316 21640 8344
rect 21315 8313 21327 8316
rect 21269 8307 21327 8313
rect 21634 8304 21640 8316
rect 21692 8304 21698 8356
rect 22094 8304 22100 8356
rect 22152 8304 22158 8356
rect 22462 8304 22468 8356
rect 22520 8304 22526 8356
rect 22572 8353 22600 8384
rect 22848 8356 22876 8384
rect 22922 8372 22928 8424
rect 22980 8412 22986 8424
rect 23400 8412 23428 8443
rect 22980 8384 23428 8412
rect 22980 8372 22986 8384
rect 22557 8347 22615 8353
rect 22557 8313 22569 8347
rect 22603 8313 22615 8347
rect 22557 8307 22615 8313
rect 22830 8304 22836 8356
rect 22888 8304 22894 8356
rect 23198 8304 23204 8356
rect 23256 8304 23262 8356
rect 23382 8304 23388 8356
rect 23440 8344 23446 8356
rect 23952 8344 23980 8443
rect 24302 8372 24308 8424
rect 24360 8412 24366 8424
rect 24872 8412 24900 8443
rect 24360 8384 24900 8412
rect 24360 8372 24366 8384
rect 25038 8372 25044 8424
rect 25096 8412 25102 8424
rect 25700 8412 25728 8443
rect 27798 8440 27804 8492
rect 27856 8480 27862 8492
rect 28077 8483 28135 8489
rect 28077 8480 28089 8483
rect 27856 8452 28089 8480
rect 27856 8440 27862 8452
rect 28077 8449 28089 8452
rect 28123 8449 28135 8483
rect 28077 8443 28135 8449
rect 28166 8440 28172 8492
rect 28224 8440 28230 8492
rect 28350 8440 28356 8492
rect 28408 8480 28414 8492
rect 29273 8483 29331 8489
rect 29273 8480 29285 8483
rect 28408 8452 29285 8480
rect 28408 8440 28414 8452
rect 29273 8449 29285 8452
rect 29319 8449 29331 8483
rect 29273 8443 29331 8449
rect 28445 8415 28503 8421
rect 28445 8412 28457 8415
rect 25096 8384 25728 8412
rect 25792 8384 28457 8412
rect 25096 8372 25102 8384
rect 23440 8316 23980 8344
rect 23440 8304 23446 8316
rect 24026 8304 24032 8356
rect 24084 8304 24090 8356
rect 24210 8304 24216 8356
rect 24268 8344 24274 8356
rect 24673 8347 24731 8353
rect 24673 8344 24685 8347
rect 24268 8316 24685 8344
rect 24268 8304 24274 8316
rect 24673 8313 24685 8316
rect 24719 8313 24731 8347
rect 24673 8307 24731 8313
rect 24762 8304 24768 8356
rect 24820 8344 24826 8356
rect 24949 8347 25007 8353
rect 24949 8344 24961 8347
rect 24820 8316 24961 8344
rect 24820 8304 24826 8316
rect 24949 8313 24961 8316
rect 24995 8313 25007 8347
rect 24949 8307 25007 8313
rect 25222 8304 25228 8356
rect 25280 8304 25286 8356
rect 25314 8304 25320 8356
rect 25372 8344 25378 8356
rect 25792 8344 25820 8384
rect 28445 8381 28457 8384
rect 28491 8381 28503 8415
rect 28445 8375 28503 8381
rect 29178 8372 29184 8424
rect 29236 8412 29242 8424
rect 29549 8415 29607 8421
rect 29549 8412 29561 8415
rect 29236 8384 29561 8412
rect 29236 8372 29242 8384
rect 29549 8381 29561 8384
rect 29595 8381 29607 8415
rect 29656 8412 29684 8520
rect 30926 8508 30932 8560
rect 30984 8548 30990 8560
rect 30984 8520 32720 8548
rect 30984 8508 30990 8520
rect 29730 8440 29736 8492
rect 29788 8480 29794 8492
rect 30653 8483 30711 8489
rect 30653 8480 30665 8483
rect 29788 8452 30665 8480
rect 29788 8440 29794 8452
rect 30653 8449 30665 8452
rect 30699 8449 30711 8483
rect 32493 8483 32551 8489
rect 32493 8480 32505 8483
rect 30653 8443 30711 8449
rect 31726 8452 32505 8480
rect 29825 8415 29883 8421
rect 29825 8412 29837 8415
rect 29656 8384 29837 8412
rect 29549 8375 29607 8381
rect 29825 8381 29837 8384
rect 29871 8381 29883 8415
rect 29825 8375 29883 8381
rect 30098 8372 30104 8424
rect 30156 8412 30162 8424
rect 31726 8412 31754 8452
rect 32493 8449 32505 8452
rect 32539 8449 32551 8483
rect 32493 8443 32551 8449
rect 32582 8440 32588 8492
rect 32640 8440 32646 8492
rect 32692 8480 32720 8520
rect 33042 8508 33048 8560
rect 33100 8548 33106 8560
rect 33100 8520 33732 8548
rect 33100 8508 33106 8520
rect 32941 8483 32999 8489
rect 32941 8480 32953 8483
rect 32692 8452 32953 8480
rect 32941 8449 32953 8452
rect 32987 8449 32999 8483
rect 32941 8443 32999 8449
rect 33321 8483 33379 8489
rect 33321 8449 33333 8483
rect 33367 8480 33379 8483
rect 33502 8480 33508 8492
rect 33367 8452 33508 8480
rect 33367 8449 33379 8452
rect 33321 8443 33379 8449
rect 33502 8440 33508 8452
rect 33560 8440 33566 8492
rect 33704 8489 33732 8520
rect 33778 8508 33784 8560
rect 33836 8548 33842 8560
rect 33836 8520 35848 8548
rect 33836 8508 33842 8520
rect 33689 8483 33747 8489
rect 33689 8449 33701 8483
rect 33735 8449 33747 8483
rect 33689 8443 33747 8449
rect 34054 8440 34060 8492
rect 34112 8440 34118 8492
rect 34698 8440 34704 8492
rect 34756 8440 34762 8492
rect 35066 8440 35072 8492
rect 35124 8440 35130 8492
rect 35250 8440 35256 8492
rect 35308 8480 35314 8492
rect 35308 8452 35664 8480
rect 35308 8440 35314 8452
rect 30156 8384 31754 8412
rect 30156 8372 30162 8384
rect 34146 8372 34152 8424
rect 34204 8412 34210 8424
rect 35636 8412 35664 8452
rect 35710 8440 35716 8492
rect 35768 8440 35774 8492
rect 35820 8489 35848 8520
rect 35894 8508 35900 8560
rect 35952 8548 35958 8560
rect 35952 8520 37320 8548
rect 35952 8508 35958 8520
rect 35805 8483 35863 8489
rect 35805 8449 35817 8483
rect 35851 8449 35863 8483
rect 35805 8443 35863 8449
rect 36170 8440 36176 8492
rect 36228 8440 36234 8492
rect 36538 8440 36544 8492
rect 36596 8440 36602 8492
rect 37292 8489 37320 8520
rect 37458 8508 37464 8560
rect 37516 8548 37522 8560
rect 38580 8548 38608 8579
rect 37516 8520 38608 8548
rect 37516 8508 37522 8520
rect 37277 8483 37335 8489
rect 37277 8449 37289 8483
rect 37323 8449 37335 8483
rect 37277 8443 37335 8449
rect 37645 8483 37703 8489
rect 37645 8449 37657 8483
rect 37691 8449 37703 8483
rect 37645 8443 37703 8449
rect 34204 8384 35296 8412
rect 35636 8384 36308 8412
rect 34204 8372 34210 8384
rect 25961 8347 26019 8353
rect 25961 8344 25973 8347
rect 25372 8316 25820 8344
rect 25884 8316 25973 8344
rect 25372 8304 25378 8316
rect 1578 8236 1584 8288
rect 1636 8236 1642 8288
rect 1857 8279 1915 8285
rect 1857 8245 1869 8279
rect 1903 8276 1915 8279
rect 2056 8276 2084 8304
rect 1903 8248 2084 8276
rect 1903 8245 1915 8248
rect 1857 8239 1915 8245
rect 2314 8236 2320 8288
rect 2372 8276 2378 8288
rect 12802 8276 12808 8288
rect 2372 8248 12808 8276
rect 2372 8236 2378 8248
rect 12802 8236 12808 8248
rect 12860 8236 12866 8288
rect 14550 8236 14556 8288
rect 14608 8276 14614 8288
rect 20346 8276 20352 8288
rect 14608 8248 20352 8276
rect 14608 8236 14614 8248
rect 20346 8236 20352 8248
rect 20404 8236 20410 8288
rect 21726 8236 21732 8288
rect 21784 8276 21790 8288
rect 22649 8279 22707 8285
rect 22649 8276 22661 8279
rect 21784 8248 22661 8276
rect 21784 8236 21790 8248
rect 22649 8245 22661 8248
rect 22695 8245 22707 8279
rect 22649 8239 22707 8245
rect 22922 8236 22928 8288
rect 22980 8236 22986 8288
rect 23566 8236 23572 8288
rect 23624 8276 23630 8288
rect 23661 8279 23719 8285
rect 23661 8276 23673 8279
rect 23624 8248 23673 8276
rect 23624 8236 23630 8248
rect 23661 8245 23673 8248
rect 23707 8245 23719 8279
rect 23661 8239 23719 8245
rect 23750 8236 23756 8288
rect 23808 8276 23814 8288
rect 24397 8279 24455 8285
rect 24397 8276 24409 8279
rect 23808 8248 24409 8276
rect 23808 8236 23814 8248
rect 24397 8245 24409 8248
rect 24443 8245 24455 8279
rect 24397 8239 24455 8245
rect 25774 8236 25780 8288
rect 25832 8276 25838 8288
rect 25884 8276 25912 8316
rect 25961 8313 25973 8316
rect 26007 8313 26019 8347
rect 25961 8307 26019 8313
rect 26326 8304 26332 8356
rect 26384 8344 26390 8356
rect 27893 8347 27951 8353
rect 27893 8344 27905 8347
rect 26384 8316 27905 8344
rect 26384 8304 26390 8316
rect 27893 8313 27905 8316
rect 27939 8313 27951 8347
rect 29089 8347 29147 8353
rect 29089 8344 29101 8347
rect 27893 8307 27951 8313
rect 28000 8316 29101 8344
rect 25832 8248 25912 8276
rect 25832 8236 25838 8248
rect 26878 8236 26884 8288
rect 26936 8276 26942 8288
rect 28000 8276 28028 8316
rect 29089 8313 29101 8316
rect 29135 8313 29147 8347
rect 29089 8307 29147 8313
rect 33410 8304 33416 8356
rect 33468 8344 33474 8356
rect 33873 8347 33931 8353
rect 33873 8344 33885 8347
rect 33468 8316 33885 8344
rect 33468 8304 33474 8316
rect 33873 8313 33885 8316
rect 33919 8313 33931 8347
rect 33873 8307 33931 8313
rect 33962 8304 33968 8356
rect 34020 8344 34026 8356
rect 35268 8353 35296 8384
rect 34885 8347 34943 8353
rect 34885 8344 34897 8347
rect 34020 8316 34897 8344
rect 34020 8304 34026 8316
rect 34885 8313 34897 8316
rect 34931 8313 34943 8347
rect 34885 8307 34943 8313
rect 35253 8347 35311 8353
rect 35253 8313 35265 8347
rect 35299 8313 35311 8347
rect 35253 8307 35311 8313
rect 35618 8304 35624 8356
rect 35676 8344 35682 8356
rect 35989 8347 36047 8353
rect 35989 8344 36001 8347
rect 35676 8316 36001 8344
rect 35676 8304 35682 8316
rect 35989 8313 36001 8316
rect 36035 8313 36047 8347
rect 35989 8307 36047 8313
rect 26936 8248 28028 8276
rect 36280 8276 36308 8384
rect 36354 8372 36360 8424
rect 36412 8372 36418 8424
rect 36906 8372 36912 8424
rect 36964 8412 36970 8424
rect 37660 8412 37688 8443
rect 37826 8440 37832 8492
rect 37884 8480 37890 8492
rect 38013 8483 38071 8489
rect 38013 8480 38025 8483
rect 37884 8452 38025 8480
rect 37884 8440 37890 8452
rect 38013 8449 38025 8452
rect 38059 8449 38071 8483
rect 38013 8443 38071 8449
rect 38378 8440 38384 8492
rect 38436 8440 38442 8492
rect 39117 8483 39175 8489
rect 39117 8449 39129 8483
rect 39163 8480 39175 8483
rect 39209 8483 39267 8489
rect 39209 8480 39221 8483
rect 39163 8452 39221 8480
rect 39163 8449 39175 8452
rect 39117 8443 39175 8449
rect 39209 8449 39221 8452
rect 39255 8449 39267 8483
rect 39209 8443 39267 8449
rect 36964 8384 37688 8412
rect 36964 8372 36970 8384
rect 36372 8344 36400 8372
rect 36372 8316 37136 8344
rect 36357 8279 36415 8285
rect 36357 8276 36369 8279
rect 36280 8248 36369 8276
rect 26936 8236 26942 8248
rect 36357 8245 36369 8248
rect 36403 8245 36415 8279
rect 37108 8276 37136 8316
rect 37182 8304 37188 8356
rect 37240 8344 37246 8356
rect 38197 8347 38255 8353
rect 38197 8344 38209 8347
rect 37240 8316 38209 8344
rect 37240 8304 37246 8316
rect 38197 8313 38209 8316
rect 38243 8313 38255 8347
rect 38197 8307 38255 8313
rect 39022 8304 39028 8356
rect 39080 8304 39086 8356
rect 39390 8304 39396 8356
rect 39448 8304 39454 8356
rect 37461 8279 37519 8285
rect 37461 8276 37473 8279
rect 37108 8248 37473 8276
rect 36357 8239 36415 8245
rect 37461 8245 37473 8248
rect 37507 8245 37519 8279
rect 37461 8239 37519 8245
rect 1104 8186 39836 8208
rect 1104 8134 1950 8186
rect 2002 8134 2014 8186
rect 2066 8134 2078 8186
rect 2130 8134 2142 8186
rect 2194 8134 2206 8186
rect 2258 8134 7950 8186
rect 8002 8134 8014 8186
rect 8066 8134 8078 8186
rect 8130 8134 8142 8186
rect 8194 8134 8206 8186
rect 8258 8134 13950 8186
rect 14002 8134 14014 8186
rect 14066 8134 14078 8186
rect 14130 8134 14142 8186
rect 14194 8134 14206 8186
rect 14258 8134 19950 8186
rect 20002 8134 20014 8186
rect 20066 8134 20078 8186
rect 20130 8134 20142 8186
rect 20194 8134 20206 8186
rect 20258 8134 25950 8186
rect 26002 8134 26014 8186
rect 26066 8134 26078 8186
rect 26130 8134 26142 8186
rect 26194 8134 26206 8186
rect 26258 8134 31950 8186
rect 32002 8134 32014 8186
rect 32066 8134 32078 8186
rect 32130 8134 32142 8186
rect 32194 8134 32206 8186
rect 32258 8134 37950 8186
rect 38002 8134 38014 8186
rect 38066 8134 38078 8186
rect 38130 8134 38142 8186
rect 38194 8134 38206 8186
rect 38258 8134 39836 8186
rect 1104 8112 39836 8134
rect 1210 8032 1216 8084
rect 1268 8072 1274 8084
rect 1268 8044 2084 8072
rect 1268 8032 1274 8044
rect 1857 8007 1915 8013
rect 1857 7973 1869 8007
rect 1903 8004 1915 8007
rect 1946 8004 1952 8016
rect 1903 7976 1952 8004
rect 1903 7973 1915 7976
rect 1857 7967 1915 7973
rect 1946 7964 1952 7976
rect 2004 7964 2010 8016
rect 1026 7896 1032 7948
rect 1084 7936 1090 7948
rect 1084 7908 1992 7936
rect 1084 7896 1090 7908
rect 750 7828 756 7880
rect 808 7868 814 7880
rect 1964 7877 1992 7908
rect 1397 7871 1455 7877
rect 1397 7868 1409 7871
rect 808 7840 1409 7868
rect 808 7828 814 7840
rect 1397 7837 1409 7840
rect 1443 7837 1455 7871
rect 1397 7831 1455 7837
rect 1673 7871 1731 7877
rect 1673 7837 1685 7871
rect 1719 7837 1731 7871
rect 1673 7831 1731 7837
rect 1949 7871 2007 7877
rect 1949 7837 1961 7871
rect 1995 7837 2007 7871
rect 2056 7868 2084 8044
rect 3418 8032 3424 8084
rect 3476 8032 3482 8084
rect 3510 8032 3516 8084
rect 3568 8072 3574 8084
rect 3878 8072 3884 8084
rect 3568 8044 3884 8072
rect 3568 8032 3574 8044
rect 3878 8032 3884 8044
rect 3936 8032 3942 8084
rect 4062 8032 4068 8084
rect 4120 8072 4126 8084
rect 4249 8075 4307 8081
rect 4249 8072 4261 8075
rect 4120 8044 4261 8072
rect 4120 8032 4126 8044
rect 4249 8041 4261 8044
rect 4295 8041 4307 8075
rect 4249 8035 4307 8041
rect 4890 8032 4896 8084
rect 4948 8072 4954 8084
rect 5169 8075 5227 8081
rect 5169 8072 5181 8075
rect 4948 8044 5181 8072
rect 4948 8032 4954 8044
rect 5169 8041 5181 8044
rect 5215 8041 5227 8075
rect 5169 8035 5227 8041
rect 5994 8032 6000 8084
rect 6052 8072 6058 8084
rect 6181 8075 6239 8081
rect 6181 8072 6193 8075
rect 6052 8044 6193 8072
rect 6052 8032 6058 8044
rect 6181 8041 6193 8044
rect 6227 8041 6239 8075
rect 6181 8035 6239 8041
rect 6546 8032 6552 8084
rect 6604 8072 6610 8084
rect 6733 8075 6791 8081
rect 6733 8072 6745 8075
rect 6604 8044 6745 8072
rect 6604 8032 6610 8044
rect 6733 8041 6745 8044
rect 6779 8041 6791 8075
rect 6733 8035 6791 8041
rect 7098 8032 7104 8084
rect 7156 8072 7162 8084
rect 7285 8075 7343 8081
rect 7285 8072 7297 8075
rect 7156 8044 7297 8072
rect 7156 8032 7162 8044
rect 7285 8041 7297 8044
rect 7331 8041 7343 8075
rect 7285 8035 7343 8041
rect 8294 8032 8300 8084
rect 8352 8072 8358 8084
rect 8481 8075 8539 8081
rect 8481 8072 8493 8075
rect 8352 8044 8493 8072
rect 8352 8032 8358 8044
rect 8481 8041 8493 8044
rect 8527 8041 8539 8075
rect 8481 8035 8539 8041
rect 8754 8032 8760 8084
rect 8812 8072 8818 8084
rect 9033 8075 9091 8081
rect 9033 8072 9045 8075
rect 8812 8044 9045 8072
rect 8812 8032 8818 8044
rect 9033 8041 9045 8044
rect 9079 8041 9091 8075
rect 9033 8035 9091 8041
rect 9398 8032 9404 8084
rect 9456 8072 9462 8084
rect 9493 8075 9551 8081
rect 9493 8072 9505 8075
rect 9456 8044 9505 8072
rect 9456 8032 9462 8044
rect 9493 8041 9505 8044
rect 9539 8041 9551 8075
rect 9493 8035 9551 8041
rect 10410 8032 10416 8084
rect 10468 8072 10474 8084
rect 10597 8075 10655 8081
rect 10597 8072 10609 8075
rect 10468 8044 10609 8072
rect 10468 8032 10474 8044
rect 10597 8041 10609 8044
rect 10643 8041 10655 8075
rect 10597 8035 10655 8041
rect 11238 8032 11244 8084
rect 11296 8072 11302 8084
rect 11425 8075 11483 8081
rect 11425 8072 11437 8075
rect 11296 8044 11437 8072
rect 11296 8032 11302 8044
rect 11425 8041 11437 8044
rect 11471 8041 11483 8075
rect 11425 8035 11483 8041
rect 11790 8032 11796 8084
rect 11848 8072 11854 8084
rect 11977 8075 12035 8081
rect 11977 8072 11989 8075
rect 11848 8044 11989 8072
rect 11848 8032 11854 8044
rect 11977 8041 11989 8044
rect 12023 8041 12035 8075
rect 11977 8035 12035 8041
rect 12618 8032 12624 8084
rect 12676 8072 12682 8084
rect 12897 8075 12955 8081
rect 12897 8072 12909 8075
rect 12676 8044 12909 8072
rect 12676 8032 12682 8044
rect 12897 8041 12909 8044
rect 12943 8041 12955 8075
rect 12897 8035 12955 8041
rect 13446 8032 13452 8084
rect 13504 8072 13510 8084
rect 13633 8075 13691 8081
rect 13633 8072 13645 8075
rect 13504 8044 13645 8072
rect 13504 8032 13510 8044
rect 13633 8041 13645 8044
rect 13679 8041 13691 8075
rect 13633 8035 13691 8041
rect 14274 8032 14280 8084
rect 14332 8072 14338 8084
rect 14461 8075 14519 8081
rect 14461 8072 14473 8075
rect 14332 8044 14473 8072
rect 14332 8032 14338 8044
rect 14461 8041 14473 8044
rect 14507 8041 14519 8075
rect 14461 8035 14519 8041
rect 14826 8032 14832 8084
rect 14884 8072 14890 8084
rect 15013 8075 15071 8081
rect 15013 8072 15025 8075
rect 14884 8044 15025 8072
rect 14884 8032 14890 8044
rect 15013 8041 15025 8044
rect 15059 8041 15071 8075
rect 15013 8035 15071 8041
rect 15930 8032 15936 8084
rect 15988 8072 15994 8084
rect 16209 8075 16267 8081
rect 16209 8072 16221 8075
rect 15988 8044 16221 8072
rect 15988 8032 15994 8044
rect 16209 8041 16221 8044
rect 16255 8041 16267 8075
rect 16209 8035 16267 8041
rect 17586 8032 17592 8084
rect 17644 8072 17650 8084
rect 17681 8075 17739 8081
rect 17681 8072 17693 8075
rect 17644 8044 17693 8072
rect 17644 8032 17650 8044
rect 17681 8041 17693 8044
rect 17727 8041 17739 8075
rect 17681 8035 17739 8041
rect 18046 8032 18052 8084
rect 18104 8072 18110 8084
rect 20530 8072 20536 8084
rect 18104 8044 20536 8072
rect 18104 8032 18110 8044
rect 20530 8032 20536 8044
rect 20588 8032 20594 8084
rect 23382 8032 23388 8084
rect 23440 8072 23446 8084
rect 23440 8044 31754 8072
rect 23440 8032 23446 8044
rect 6914 7964 6920 8016
rect 6972 8004 6978 8016
rect 6972 7976 8340 8004
rect 6972 7964 6978 7976
rect 2130 7896 2136 7948
rect 2188 7936 2194 7948
rect 3878 7936 3884 7948
rect 2188 7908 3884 7936
rect 2188 7896 2194 7908
rect 3878 7896 3884 7908
rect 3936 7896 3942 7948
rect 8202 7936 8208 7948
rect 4448 7908 8208 7936
rect 2225 7871 2283 7877
rect 2225 7868 2237 7871
rect 2056 7840 2237 7868
rect 1949 7831 2007 7837
rect 2225 7837 2237 7840
rect 2271 7837 2283 7871
rect 2225 7831 2283 7837
rect 566 7760 572 7812
rect 624 7800 630 7812
rect 1688 7800 1716 7831
rect 3602 7828 3608 7880
rect 3660 7828 3666 7880
rect 4448 7877 4476 7908
rect 8202 7896 8208 7908
rect 8260 7896 8266 7948
rect 8312 7936 8340 7976
rect 11882 7964 11888 8016
rect 11940 8004 11946 8016
rect 16850 8004 16856 8016
rect 11940 7976 16856 8004
rect 11940 7964 11946 7976
rect 16850 7964 16856 7976
rect 16908 7964 16914 8016
rect 18141 8007 18199 8013
rect 18141 7973 18153 8007
rect 18187 8004 18199 8007
rect 20622 8004 20628 8016
rect 18187 7976 20628 8004
rect 18187 7973 18199 7976
rect 18141 7967 18199 7973
rect 20622 7964 20628 7976
rect 20680 8004 20686 8016
rect 23014 8004 23020 8016
rect 20680 7976 23020 8004
rect 20680 7964 20686 7976
rect 23014 7964 23020 7976
rect 23072 7964 23078 8016
rect 23198 7964 23204 8016
rect 23256 8004 23262 8016
rect 23750 8004 23756 8016
rect 23256 7976 23756 8004
rect 23256 7964 23262 7976
rect 23750 7964 23756 7976
rect 23808 7964 23814 8016
rect 28902 7964 28908 8016
rect 28960 8004 28966 8016
rect 31726 8004 31754 8044
rect 34422 8032 34428 8084
rect 34480 8072 34486 8084
rect 34885 8075 34943 8081
rect 34885 8072 34897 8075
rect 34480 8044 34897 8072
rect 34480 8032 34486 8044
rect 34885 8041 34897 8044
rect 34931 8041 34943 8075
rect 34885 8035 34943 8041
rect 35526 8032 35532 8084
rect 35584 8072 35590 8084
rect 35805 8075 35863 8081
rect 35805 8072 35817 8075
rect 35584 8044 35817 8072
rect 35584 8032 35590 8044
rect 35805 8041 35817 8044
rect 35851 8041 35863 8075
rect 35805 8035 35863 8041
rect 36078 8032 36084 8084
rect 36136 8072 36142 8084
rect 36357 8075 36415 8081
rect 36357 8072 36369 8075
rect 36136 8044 36369 8072
rect 36136 8032 36142 8044
rect 36357 8041 36369 8044
rect 36403 8041 36415 8075
rect 36357 8035 36415 8041
rect 36630 8032 36636 8084
rect 36688 8072 36694 8084
rect 36909 8075 36967 8081
rect 36909 8072 36921 8075
rect 36688 8044 36921 8072
rect 36688 8032 36694 8044
rect 36909 8041 36921 8044
rect 36955 8041 36967 8075
rect 36909 8035 36967 8041
rect 37734 8032 37740 8084
rect 37792 8072 37798 8084
rect 37921 8075 37979 8081
rect 37921 8072 37933 8075
rect 37792 8044 37933 8072
rect 37792 8032 37798 8044
rect 37921 8041 37933 8044
rect 37967 8041 37979 8075
rect 37921 8035 37979 8041
rect 38654 8032 38660 8084
rect 38712 8032 38718 8084
rect 37458 8004 37464 8016
rect 28960 7976 29224 8004
rect 31726 7976 37464 8004
rect 28960 7964 28966 7976
rect 8312 7908 12434 7936
rect 4433 7871 4491 7877
rect 4433 7837 4445 7871
rect 4479 7837 4491 7871
rect 4433 7831 4491 7837
rect 4706 7828 4712 7880
rect 4764 7868 4770 7880
rect 4985 7871 5043 7877
rect 4985 7868 4997 7871
rect 4764 7840 4997 7868
rect 4764 7828 4770 7840
rect 4985 7837 4997 7840
rect 5031 7837 5043 7871
rect 4985 7831 5043 7837
rect 6365 7871 6423 7877
rect 6365 7837 6377 7871
rect 6411 7837 6423 7871
rect 6365 7831 6423 7837
rect 6917 7871 6975 7877
rect 6917 7837 6929 7871
rect 6963 7868 6975 7871
rect 7190 7868 7196 7880
rect 6963 7840 7196 7868
rect 6963 7837 6975 7840
rect 6917 7831 6975 7837
rect 6178 7800 6184 7812
rect 624 7772 1716 7800
rect 2056 7772 6184 7800
rect 624 7760 630 7772
rect 1581 7735 1639 7741
rect 1581 7701 1593 7735
rect 1627 7732 1639 7735
rect 2056 7732 2084 7772
rect 6178 7760 6184 7772
rect 6236 7760 6242 7812
rect 1627 7704 2084 7732
rect 1627 7701 1639 7704
rect 1581 7695 1639 7701
rect 2130 7692 2136 7744
rect 2188 7692 2194 7744
rect 2409 7735 2467 7741
rect 2409 7701 2421 7735
rect 2455 7732 2467 7735
rect 6270 7732 6276 7744
rect 2455 7704 6276 7732
rect 2455 7701 2467 7704
rect 2409 7695 2467 7701
rect 6270 7692 6276 7704
rect 6328 7692 6334 7744
rect 6380 7732 6408 7831
rect 7190 7828 7196 7840
rect 7248 7828 7254 7880
rect 7469 7871 7527 7877
rect 7469 7837 7481 7871
rect 7515 7837 7527 7871
rect 7469 7831 7527 7837
rect 7484 7800 7512 7831
rect 8294 7828 8300 7880
rect 8352 7828 8358 7880
rect 9214 7828 9220 7880
rect 9272 7828 9278 7880
rect 9674 7828 9680 7880
rect 9732 7828 9738 7880
rect 10778 7828 10784 7880
rect 10836 7828 10842 7880
rect 11609 7871 11667 7877
rect 11609 7837 11621 7871
rect 11655 7837 11667 7871
rect 11609 7831 11667 7837
rect 8846 7800 8852 7812
rect 7484 7772 8852 7800
rect 8846 7760 8852 7772
rect 8904 7760 8910 7812
rect 11624 7800 11652 7831
rect 12158 7828 12164 7880
rect 12216 7828 12222 7880
rect 12406 7868 12434 7908
rect 13170 7896 13176 7948
rect 13228 7936 13234 7948
rect 13228 7908 16068 7936
rect 13228 7896 13234 7908
rect 12713 7871 12771 7877
rect 12713 7868 12725 7871
rect 12406 7840 12725 7868
rect 12713 7837 12725 7840
rect 12759 7837 12771 7871
rect 12713 7831 12771 7837
rect 13814 7828 13820 7880
rect 13872 7828 13878 7880
rect 14642 7828 14648 7880
rect 14700 7828 14706 7880
rect 16040 7877 16068 7908
rect 16206 7896 16212 7948
rect 16264 7936 16270 7948
rect 22922 7936 22928 7948
rect 16264 7908 22928 7936
rect 16264 7896 16270 7908
rect 22922 7896 22928 7908
rect 22980 7896 22986 7948
rect 28994 7936 29000 7948
rect 26896 7908 29000 7936
rect 15197 7871 15255 7877
rect 15197 7837 15209 7871
rect 15243 7837 15255 7871
rect 15197 7831 15255 7837
rect 16025 7871 16083 7877
rect 16025 7837 16037 7871
rect 16071 7837 16083 7871
rect 16025 7831 16083 7837
rect 16132 7840 17264 7868
rect 13722 7800 13728 7812
rect 11624 7772 13728 7800
rect 13722 7760 13728 7772
rect 13780 7760 13786 7812
rect 15212 7800 15240 7831
rect 16132 7800 16160 7840
rect 15212 7772 16160 7800
rect 17236 7800 17264 7840
rect 17862 7828 17868 7880
rect 17920 7868 17926 7880
rect 17957 7871 18015 7877
rect 17957 7868 17969 7871
rect 17920 7840 17969 7868
rect 17920 7828 17926 7840
rect 17957 7837 17969 7840
rect 18003 7837 18015 7871
rect 17957 7831 18015 7837
rect 18138 7828 18144 7880
rect 18196 7868 18202 7880
rect 18417 7871 18475 7877
rect 18417 7868 18429 7871
rect 18196 7840 18429 7868
rect 18196 7828 18202 7840
rect 18417 7837 18429 7840
rect 18463 7837 18475 7871
rect 18417 7831 18475 7837
rect 19518 7828 19524 7880
rect 19576 7868 19582 7880
rect 20530 7868 20536 7880
rect 19576 7840 20536 7868
rect 19576 7828 19582 7840
rect 20530 7828 20536 7840
rect 20588 7828 20594 7880
rect 20714 7828 20720 7880
rect 20772 7868 20778 7880
rect 26896 7868 26924 7908
rect 28994 7896 29000 7908
rect 29052 7896 29058 7948
rect 20772 7840 26924 7868
rect 20772 7828 20778 7840
rect 28626 7828 28632 7880
rect 28684 7868 28690 7880
rect 29196 7877 29224 7976
rect 37458 7964 37464 7976
rect 37516 7964 37522 8016
rect 30742 7896 30748 7948
rect 30800 7936 30806 7948
rect 30800 7908 38884 7936
rect 30800 7896 30806 7908
rect 28905 7871 28963 7877
rect 28905 7868 28917 7871
rect 28684 7840 28917 7868
rect 28684 7828 28690 7840
rect 28905 7837 28917 7840
rect 28951 7837 28963 7871
rect 28905 7831 28963 7837
rect 29181 7871 29239 7877
rect 29181 7837 29193 7871
rect 29227 7837 29239 7871
rect 29181 7831 29239 7837
rect 29454 7828 29460 7880
rect 29512 7868 29518 7880
rect 29733 7871 29791 7877
rect 29733 7868 29745 7871
rect 29512 7840 29745 7868
rect 29512 7828 29518 7840
rect 29733 7837 29745 7840
rect 29779 7837 29791 7871
rect 29733 7831 29791 7837
rect 29914 7828 29920 7880
rect 29972 7868 29978 7880
rect 31570 7868 31576 7880
rect 29972 7840 31576 7868
rect 29972 7828 29978 7840
rect 31570 7828 31576 7840
rect 31628 7828 31634 7880
rect 33410 7828 33416 7880
rect 33468 7868 33474 7880
rect 34701 7871 34759 7877
rect 34701 7868 34713 7871
rect 33468 7840 34713 7868
rect 33468 7828 33474 7840
rect 34701 7837 34713 7840
rect 34747 7837 34759 7871
rect 34701 7831 34759 7837
rect 35618 7828 35624 7880
rect 35676 7828 35682 7880
rect 36170 7828 36176 7880
rect 36228 7828 36234 7880
rect 36722 7828 36728 7880
rect 36780 7828 36786 7880
rect 37826 7828 37832 7880
rect 37884 7868 37890 7880
rect 38856 7877 38884 7908
rect 38105 7871 38163 7877
rect 38105 7868 38117 7871
rect 37884 7840 38117 7868
rect 37884 7828 37890 7840
rect 38105 7837 38117 7840
rect 38151 7837 38163 7871
rect 38105 7831 38163 7837
rect 38473 7871 38531 7877
rect 38473 7837 38485 7871
rect 38519 7837 38531 7871
rect 38473 7831 38531 7837
rect 38841 7871 38899 7877
rect 38841 7837 38853 7871
rect 38887 7837 38899 7871
rect 38841 7831 38899 7837
rect 39209 7871 39267 7877
rect 39209 7837 39221 7871
rect 39255 7837 39267 7871
rect 39209 7831 39267 7837
rect 31294 7800 31300 7812
rect 17236 7772 31300 7800
rect 31294 7760 31300 7772
rect 31352 7760 31358 7812
rect 37274 7760 37280 7812
rect 37332 7800 37338 7812
rect 38488 7800 38516 7831
rect 39224 7800 39252 7831
rect 37332 7772 38516 7800
rect 38580 7772 39252 7800
rect 37332 7760 37338 7772
rect 9858 7732 9864 7744
rect 6380 7704 9864 7732
rect 9858 7692 9864 7704
rect 9916 7692 9922 7744
rect 13354 7692 13360 7744
rect 13412 7732 13418 7744
rect 14550 7732 14556 7744
rect 13412 7704 14556 7732
rect 13412 7692 13418 7704
rect 14550 7692 14556 7704
rect 14608 7692 14614 7744
rect 14642 7692 14648 7744
rect 14700 7732 14706 7744
rect 16206 7732 16212 7744
rect 14700 7704 16212 7732
rect 14700 7692 14706 7704
rect 16206 7692 16212 7704
rect 16264 7692 16270 7744
rect 18230 7692 18236 7744
rect 18288 7692 18294 7744
rect 18874 7692 18880 7744
rect 18932 7732 18938 7744
rect 22370 7732 22376 7744
rect 18932 7704 22376 7732
rect 18932 7692 18938 7704
rect 22370 7692 22376 7704
rect 22428 7692 22434 7744
rect 24578 7692 24584 7744
rect 24636 7732 24642 7744
rect 28721 7735 28779 7741
rect 28721 7732 28733 7735
rect 24636 7704 28733 7732
rect 24636 7692 24642 7704
rect 28721 7701 28733 7704
rect 28767 7701 28779 7735
rect 28721 7695 28779 7701
rect 28810 7692 28816 7744
rect 28868 7732 28874 7744
rect 28997 7735 29055 7741
rect 28997 7732 29009 7735
rect 28868 7704 29009 7732
rect 28868 7692 28874 7704
rect 28997 7701 29009 7704
rect 29043 7701 29055 7735
rect 28997 7695 29055 7701
rect 29546 7692 29552 7744
rect 29604 7692 29610 7744
rect 31110 7692 31116 7744
rect 31168 7732 31174 7744
rect 32582 7732 32588 7744
rect 31168 7704 32588 7732
rect 31168 7692 31174 7704
rect 32582 7692 32588 7704
rect 32640 7692 32646 7744
rect 32766 7692 32772 7744
rect 32824 7732 32830 7744
rect 38580 7732 38608 7772
rect 32824 7704 38608 7732
rect 32824 7692 32830 7704
rect 38930 7692 38936 7744
rect 38988 7732 38994 7744
rect 39025 7735 39083 7741
rect 39025 7732 39037 7735
rect 38988 7704 39037 7732
rect 38988 7692 38994 7704
rect 39025 7701 39037 7704
rect 39071 7701 39083 7735
rect 39025 7695 39083 7701
rect 39390 7692 39396 7744
rect 39448 7692 39454 7744
rect 1104 7642 39836 7664
rect 1104 7590 3010 7642
rect 3062 7590 3074 7642
rect 3126 7590 3138 7642
rect 3190 7590 3202 7642
rect 3254 7590 3266 7642
rect 3318 7590 9010 7642
rect 9062 7590 9074 7642
rect 9126 7590 9138 7642
rect 9190 7590 9202 7642
rect 9254 7590 9266 7642
rect 9318 7590 15010 7642
rect 15062 7590 15074 7642
rect 15126 7590 15138 7642
rect 15190 7590 15202 7642
rect 15254 7590 15266 7642
rect 15318 7590 21010 7642
rect 21062 7590 21074 7642
rect 21126 7590 21138 7642
rect 21190 7590 21202 7642
rect 21254 7590 21266 7642
rect 21318 7590 27010 7642
rect 27062 7590 27074 7642
rect 27126 7590 27138 7642
rect 27190 7590 27202 7642
rect 27254 7590 27266 7642
rect 27318 7590 33010 7642
rect 33062 7590 33074 7642
rect 33126 7590 33138 7642
rect 33190 7590 33202 7642
rect 33254 7590 33266 7642
rect 33318 7590 39010 7642
rect 39062 7590 39074 7642
rect 39126 7590 39138 7642
rect 39190 7590 39202 7642
rect 39254 7590 39266 7642
rect 39318 7590 39836 7642
rect 1104 7568 39836 7590
rect 1857 7531 1915 7537
rect 1857 7497 1869 7531
rect 1903 7528 1915 7531
rect 4065 7531 4123 7537
rect 1903 7500 4016 7528
rect 1903 7497 1915 7500
rect 1857 7491 1915 7497
rect 934 7420 940 7472
rect 992 7460 998 7472
rect 992 7432 1716 7460
rect 992 7420 998 7432
rect 750 7352 756 7404
rect 808 7392 814 7404
rect 1688 7401 1716 7432
rect 2130 7420 2136 7472
rect 2188 7460 2194 7472
rect 3786 7460 3792 7472
rect 2188 7432 3792 7460
rect 2188 7420 2194 7432
rect 3786 7420 3792 7432
rect 3844 7420 3850 7472
rect 1397 7395 1455 7401
rect 1397 7392 1409 7395
rect 808 7364 1409 7392
rect 808 7352 814 7364
rect 1397 7361 1409 7364
rect 1443 7361 1455 7395
rect 1397 7355 1455 7361
rect 1673 7395 1731 7401
rect 1673 7361 1685 7395
rect 1719 7361 1731 7395
rect 1673 7355 1731 7361
rect 1949 7395 2007 7401
rect 1949 7361 1961 7395
rect 1995 7361 2007 7395
rect 1949 7355 2007 7361
rect 934 7284 940 7336
rect 992 7324 998 7336
rect 1964 7324 1992 7355
rect 2866 7352 2872 7404
rect 2924 7352 2930 7404
rect 3237 7395 3295 7401
rect 3237 7361 3249 7395
rect 3283 7392 3295 7395
rect 3418 7392 3424 7404
rect 3283 7364 3424 7392
rect 3283 7361 3295 7364
rect 3237 7355 3295 7361
rect 3418 7352 3424 7364
rect 3476 7352 3482 7404
rect 3510 7352 3516 7404
rect 3568 7392 3574 7404
rect 3697 7395 3755 7401
rect 3697 7392 3709 7395
rect 3568 7364 3709 7392
rect 3568 7352 3574 7364
rect 3697 7361 3709 7364
rect 3743 7392 3755 7395
rect 3881 7395 3939 7401
rect 3881 7392 3893 7395
rect 3743 7364 3893 7392
rect 3743 7361 3755 7364
rect 3697 7355 3755 7361
rect 3881 7361 3893 7364
rect 3927 7361 3939 7395
rect 3881 7355 3939 7361
rect 3988 7324 4016 7500
rect 4065 7497 4077 7531
rect 4111 7528 4123 7531
rect 4522 7528 4528 7540
rect 4111 7500 4528 7528
rect 4111 7497 4123 7500
rect 4065 7491 4123 7497
rect 4522 7488 4528 7500
rect 4580 7488 4586 7540
rect 4706 7488 4712 7540
rect 4764 7488 4770 7540
rect 6178 7488 6184 7540
rect 6236 7528 6242 7540
rect 10134 7528 10140 7540
rect 6236 7500 10140 7528
rect 6236 7488 6242 7500
rect 10134 7488 10140 7500
rect 10192 7488 10198 7540
rect 12158 7488 12164 7540
rect 12216 7528 12222 7540
rect 19153 7531 19211 7537
rect 19153 7528 19165 7531
rect 12216 7500 19165 7528
rect 12216 7488 12222 7500
rect 19153 7497 19165 7500
rect 19199 7497 19211 7531
rect 19153 7491 19211 7497
rect 19334 7488 19340 7540
rect 19392 7528 19398 7540
rect 21545 7531 21603 7537
rect 19392 7500 21282 7528
rect 19392 7488 19398 7500
rect 21254 7472 21282 7500
rect 21545 7497 21557 7531
rect 21591 7528 21603 7531
rect 21910 7528 21916 7540
rect 21591 7500 21916 7528
rect 21591 7497 21603 7500
rect 21545 7491 21603 7497
rect 21910 7488 21916 7500
rect 21968 7528 21974 7540
rect 21968 7500 22692 7528
rect 21968 7488 21974 7500
rect 13354 7460 13360 7472
rect 4540 7432 13360 7460
rect 4062 7352 4068 7404
rect 4120 7392 4126 7404
rect 4540 7401 4568 7432
rect 13354 7420 13360 7432
rect 13412 7420 13418 7472
rect 13814 7420 13820 7472
rect 13872 7460 13878 7472
rect 13872 7432 21220 7460
rect 21254 7432 21272 7472
rect 13872 7420 13878 7432
rect 4249 7395 4307 7401
rect 4249 7392 4261 7395
rect 4120 7364 4261 7392
rect 4120 7352 4126 7364
rect 4249 7361 4261 7364
rect 4295 7361 4307 7395
rect 4249 7355 4307 7361
rect 4525 7395 4583 7401
rect 4525 7361 4537 7395
rect 4571 7361 4583 7395
rect 4525 7355 4583 7361
rect 6270 7352 6276 7404
rect 6328 7392 6334 7404
rect 13078 7392 13084 7404
rect 6328 7364 13084 7392
rect 6328 7352 6334 7364
rect 13078 7352 13084 7364
rect 13136 7352 13142 7404
rect 14093 7395 14151 7401
rect 14093 7392 14105 7395
rect 13280 7364 14105 7392
rect 7466 7324 7472 7336
rect 992 7296 1992 7324
rect 2746 7296 3188 7324
rect 3988 7296 7472 7324
rect 992 7284 998 7296
rect 1581 7259 1639 7265
rect 1581 7225 1593 7259
rect 1627 7256 1639 7259
rect 2746 7256 2774 7296
rect 1627 7228 2774 7256
rect 1627 7225 1639 7228
rect 1581 7219 1639 7225
rect 3050 7216 3056 7268
rect 3108 7216 3114 7268
rect 3160 7256 3188 7296
rect 7466 7284 7472 7296
rect 7524 7284 7530 7336
rect 10134 7284 10140 7336
rect 10192 7324 10198 7336
rect 13280 7324 13308 7364
rect 14093 7361 14105 7364
rect 14139 7361 14151 7395
rect 14093 7355 14151 7361
rect 14182 7352 14188 7404
rect 14240 7392 14246 7404
rect 15470 7392 15476 7404
rect 14240 7364 15476 7392
rect 14240 7352 14246 7364
rect 15470 7352 15476 7364
rect 15528 7352 15534 7404
rect 19242 7352 19248 7404
rect 19300 7392 19306 7404
rect 19337 7395 19395 7401
rect 19337 7392 19349 7395
rect 19300 7364 19349 7392
rect 19300 7352 19306 7364
rect 19337 7361 19349 7364
rect 19383 7361 19395 7395
rect 20809 7395 20867 7401
rect 20809 7392 20821 7395
rect 19337 7355 19395 7361
rect 19444 7364 20821 7392
rect 10192 7296 13308 7324
rect 14369 7327 14427 7333
rect 10192 7284 10198 7296
rect 14369 7293 14381 7327
rect 14415 7324 14427 7327
rect 15102 7324 15108 7336
rect 14415 7296 15108 7324
rect 14415 7293 14427 7296
rect 14369 7287 14427 7293
rect 15102 7284 15108 7296
rect 15160 7284 15166 7336
rect 19168 7296 19334 7324
rect 3160 7228 4384 7256
rect 2133 7191 2191 7197
rect 2133 7157 2145 7191
rect 2179 7188 2191 7191
rect 2314 7188 2320 7200
rect 2179 7160 2320 7188
rect 2179 7157 2191 7160
rect 2133 7151 2191 7157
rect 2314 7148 2320 7160
rect 2372 7148 2378 7200
rect 3329 7191 3387 7197
rect 3329 7157 3341 7191
rect 3375 7188 3387 7191
rect 3602 7188 3608 7200
rect 3375 7160 3608 7188
rect 3375 7157 3387 7160
rect 3329 7151 3387 7157
rect 3602 7148 3608 7160
rect 3660 7148 3666 7200
rect 4356 7188 4384 7228
rect 4430 7216 4436 7268
rect 4488 7216 4494 7268
rect 12802 7216 12808 7268
rect 12860 7256 12866 7268
rect 19168 7256 19196 7296
rect 12860 7228 13768 7256
rect 12860 7216 12866 7228
rect 7558 7188 7564 7200
rect 4356 7160 7564 7188
rect 7558 7148 7564 7160
rect 7616 7148 7622 7200
rect 12710 7148 12716 7200
rect 12768 7188 12774 7200
rect 13357 7191 13415 7197
rect 13357 7188 13369 7191
rect 12768 7160 13369 7188
rect 12768 7148 12774 7160
rect 13357 7157 13369 7160
rect 13403 7157 13415 7191
rect 13740 7188 13768 7228
rect 14292 7228 19196 7256
rect 19306 7256 19334 7296
rect 19444 7256 19472 7364
rect 20809 7361 20821 7364
rect 20855 7361 20867 7395
rect 20809 7355 20867 7361
rect 20438 7284 20444 7336
rect 20496 7324 20502 7336
rect 20533 7327 20591 7333
rect 20533 7324 20545 7327
rect 20496 7296 20545 7324
rect 20496 7284 20502 7296
rect 20533 7293 20545 7296
rect 20579 7293 20591 7327
rect 20533 7287 20591 7293
rect 19306 7228 19472 7256
rect 21192 7256 21220 7432
rect 21266 7420 21272 7432
rect 21324 7460 21330 7472
rect 21726 7460 21732 7472
rect 21324 7432 21732 7460
rect 21324 7420 21330 7432
rect 21726 7420 21732 7432
rect 21784 7420 21790 7472
rect 21818 7420 21824 7472
rect 21876 7460 21882 7472
rect 21876 7432 21956 7460
rect 21876 7420 21882 7432
rect 21928 7401 21956 7432
rect 22278 7420 22284 7472
rect 22336 7420 22342 7472
rect 22370 7420 22376 7472
rect 22428 7420 22434 7472
rect 21913 7395 21971 7401
rect 21913 7361 21925 7395
rect 21959 7361 21971 7395
rect 21913 7355 21971 7361
rect 22094 7352 22100 7404
rect 22152 7352 22158 7404
rect 22557 7395 22615 7401
rect 22557 7361 22569 7395
rect 22603 7361 22615 7395
rect 22664 7392 22692 7500
rect 30834 7488 30840 7540
rect 30892 7528 30898 7540
rect 34425 7531 34483 7537
rect 30892 7500 32352 7528
rect 30892 7488 30898 7500
rect 25498 7420 25504 7472
rect 25556 7460 25562 7472
rect 29546 7460 29552 7472
rect 25556 7432 29552 7460
rect 25556 7420 25562 7432
rect 29546 7420 29552 7432
rect 29604 7420 29610 7472
rect 30282 7420 30288 7472
rect 30340 7460 30346 7472
rect 30340 7432 31524 7460
rect 30340 7420 30346 7432
rect 22833 7395 22891 7401
rect 22833 7392 22845 7395
rect 22664 7364 22845 7392
rect 22557 7355 22615 7361
rect 22833 7361 22845 7364
rect 22879 7361 22891 7395
rect 22833 7355 22891 7361
rect 21358 7284 21364 7336
rect 21416 7324 21422 7336
rect 21821 7327 21879 7333
rect 21821 7324 21833 7327
rect 21416 7296 21833 7324
rect 21416 7284 21422 7296
rect 21821 7293 21833 7296
rect 21867 7293 21879 7327
rect 21821 7287 21879 7293
rect 22002 7284 22008 7336
rect 22060 7324 22066 7336
rect 22572 7324 22600 7355
rect 23014 7352 23020 7404
rect 23072 7352 23078 7404
rect 24118 7352 24124 7404
rect 24176 7392 24182 7404
rect 27246 7392 27252 7404
rect 24176 7364 27252 7392
rect 24176 7352 24182 7364
rect 27246 7352 27252 7364
rect 27304 7352 27310 7404
rect 30006 7352 30012 7404
rect 30064 7392 30070 7404
rect 31496 7401 31524 7432
rect 31588 7432 31800 7460
rect 31205 7395 31263 7401
rect 31205 7392 31217 7395
rect 30064 7364 31217 7392
rect 30064 7352 30070 7364
rect 31205 7361 31217 7364
rect 31251 7361 31263 7395
rect 31205 7355 31263 7361
rect 31481 7395 31539 7401
rect 31481 7361 31493 7395
rect 31527 7361 31539 7395
rect 31481 7355 31539 7361
rect 22060 7296 22600 7324
rect 22060 7284 22066 7296
rect 22738 7284 22744 7336
rect 22796 7324 22802 7336
rect 28810 7324 28816 7336
rect 22796 7296 28816 7324
rect 22796 7284 22802 7296
rect 28810 7284 28816 7296
rect 28868 7284 28874 7336
rect 30558 7284 30564 7336
rect 30616 7324 30622 7336
rect 31588 7324 31616 7432
rect 31772 7401 31800 7432
rect 32324 7401 32352 7500
rect 34425 7497 34437 7531
rect 34471 7528 34483 7531
rect 36170 7528 36176 7540
rect 34471 7500 36176 7528
rect 34471 7497 34483 7500
rect 34425 7491 34483 7497
rect 36170 7488 36176 7500
rect 36228 7488 36234 7540
rect 36262 7488 36268 7540
rect 36320 7528 36326 7540
rect 36320 7500 38240 7528
rect 36320 7488 36326 7500
rect 35894 7420 35900 7472
rect 35952 7460 35958 7472
rect 35952 7432 38148 7460
rect 35952 7420 35958 7432
rect 31757 7395 31815 7401
rect 31757 7361 31769 7395
rect 31803 7361 31815 7395
rect 31757 7355 31815 7361
rect 32309 7395 32367 7401
rect 32309 7361 32321 7395
rect 32355 7361 32367 7395
rect 32309 7355 32367 7361
rect 32582 7352 32588 7404
rect 32640 7352 32646 7404
rect 32861 7395 32919 7401
rect 32861 7361 32873 7395
rect 32907 7361 32919 7395
rect 32861 7355 32919 7361
rect 33505 7395 33563 7401
rect 33505 7361 33517 7395
rect 33551 7361 33563 7395
rect 33505 7355 33563 7361
rect 30616 7296 31616 7324
rect 30616 7284 30622 7296
rect 31662 7284 31668 7336
rect 31720 7324 31726 7336
rect 32876 7324 32904 7355
rect 31720 7296 32904 7324
rect 31720 7284 31726 7296
rect 32677 7259 32735 7265
rect 32677 7256 32689 7259
rect 21192 7228 32689 7256
rect 14292 7188 14320 7228
rect 32677 7225 32689 7228
rect 32723 7225 32735 7259
rect 32677 7219 32735 7225
rect 13740 7160 14320 7188
rect 13357 7151 13415 7157
rect 14458 7148 14464 7200
rect 14516 7188 14522 7200
rect 15378 7188 15384 7200
rect 14516 7160 15384 7188
rect 14516 7148 14522 7160
rect 15378 7148 15384 7160
rect 15436 7148 15442 7200
rect 15562 7148 15568 7200
rect 15620 7188 15626 7200
rect 15838 7188 15844 7200
rect 15620 7160 15844 7188
rect 15620 7148 15626 7160
rect 15838 7148 15844 7160
rect 15896 7148 15902 7200
rect 17770 7148 17776 7200
rect 17828 7188 17834 7200
rect 19242 7188 19248 7200
rect 17828 7160 19248 7188
rect 17828 7148 17834 7160
rect 19242 7148 19248 7160
rect 19300 7188 19306 7200
rect 24762 7188 24768 7200
rect 19300 7160 24768 7188
rect 19300 7148 19306 7160
rect 24762 7148 24768 7160
rect 24820 7148 24826 7200
rect 30466 7148 30472 7200
rect 30524 7188 30530 7200
rect 31021 7191 31079 7197
rect 31021 7188 31033 7191
rect 30524 7160 31033 7188
rect 30524 7148 30530 7160
rect 31021 7157 31033 7160
rect 31067 7157 31079 7191
rect 31021 7151 31079 7157
rect 31294 7148 31300 7200
rect 31352 7148 31358 7200
rect 31570 7148 31576 7200
rect 31628 7148 31634 7200
rect 32122 7148 32128 7200
rect 32180 7148 32186 7200
rect 32398 7148 32404 7200
rect 32456 7148 32462 7200
rect 32582 7148 32588 7200
rect 32640 7188 32646 7200
rect 33520 7188 33548 7355
rect 34238 7352 34244 7404
rect 34296 7352 34302 7404
rect 37366 7352 37372 7404
rect 37424 7392 37430 7404
rect 37461 7395 37519 7401
rect 37461 7392 37473 7395
rect 37424 7364 37473 7392
rect 37424 7352 37430 7364
rect 37461 7361 37473 7364
rect 37507 7361 37519 7395
rect 37461 7355 37519 7361
rect 37550 7352 37556 7404
rect 37608 7392 37614 7404
rect 38120 7401 38148 7432
rect 37737 7395 37795 7401
rect 37737 7392 37749 7395
rect 37608 7364 37749 7392
rect 37608 7352 37614 7364
rect 37737 7361 37749 7364
rect 37783 7361 37795 7395
rect 37737 7355 37795 7361
rect 38105 7395 38163 7401
rect 38105 7361 38117 7395
rect 38151 7361 38163 7395
rect 38212 7392 38240 7500
rect 38286 7488 38292 7540
rect 38344 7488 38350 7540
rect 38657 7531 38715 7537
rect 38657 7497 38669 7531
rect 38703 7528 38715 7531
rect 38746 7528 38752 7540
rect 38703 7500 38752 7528
rect 38703 7497 38715 7500
rect 38657 7491 38715 7497
rect 38746 7488 38752 7500
rect 38804 7488 38810 7540
rect 39025 7531 39083 7537
rect 39025 7497 39037 7531
rect 39071 7497 39083 7531
rect 39025 7491 39083 7497
rect 39393 7531 39451 7537
rect 39393 7497 39405 7531
rect 39439 7528 39451 7531
rect 39482 7528 39488 7540
rect 39439 7500 39488 7528
rect 39439 7497 39451 7500
rect 39393 7491 39451 7497
rect 39040 7460 39068 7491
rect 39482 7488 39488 7500
rect 39540 7488 39546 7540
rect 39850 7460 39856 7472
rect 39040 7432 39856 7460
rect 39850 7420 39856 7432
rect 39908 7420 39914 7472
rect 38473 7395 38531 7401
rect 38473 7392 38485 7395
rect 38212 7364 38485 7392
rect 38105 7355 38163 7361
rect 38473 7361 38485 7364
rect 38519 7361 38531 7395
rect 38473 7355 38531 7361
rect 38838 7352 38844 7404
rect 38896 7352 38902 7404
rect 39022 7352 39028 7404
rect 39080 7392 39086 7404
rect 39209 7395 39267 7401
rect 39209 7392 39221 7395
rect 39080 7364 39221 7392
rect 39080 7352 39086 7364
rect 39209 7361 39221 7364
rect 39255 7361 39267 7395
rect 39209 7355 39267 7361
rect 38930 7324 38936 7336
rect 37660 7296 38936 7324
rect 33689 7259 33747 7265
rect 33689 7225 33701 7259
rect 33735 7256 33747 7259
rect 36538 7256 36544 7268
rect 33735 7228 36544 7256
rect 33735 7225 33747 7228
rect 33689 7219 33747 7225
rect 36538 7216 36544 7228
rect 36596 7216 36602 7268
rect 37660 7265 37688 7296
rect 38930 7284 38936 7296
rect 38988 7284 38994 7336
rect 37645 7259 37703 7265
rect 37645 7225 37657 7259
rect 37691 7225 37703 7259
rect 37645 7219 37703 7225
rect 37921 7259 37979 7265
rect 37921 7225 37933 7259
rect 37967 7256 37979 7259
rect 39482 7256 39488 7268
rect 37967 7228 39488 7256
rect 37967 7225 37979 7228
rect 37921 7219 37979 7225
rect 39482 7216 39488 7228
rect 39540 7216 39546 7268
rect 32640 7160 33548 7188
rect 32640 7148 32646 7160
rect 35986 7148 35992 7200
rect 36044 7188 36050 7200
rect 38838 7188 38844 7200
rect 36044 7160 38844 7188
rect 36044 7148 36050 7160
rect 38838 7148 38844 7160
rect 38896 7148 38902 7200
rect 1104 7098 39836 7120
rect 1104 7046 1950 7098
rect 2002 7046 2014 7098
rect 2066 7046 2078 7098
rect 2130 7046 2142 7098
rect 2194 7046 2206 7098
rect 2258 7046 7950 7098
rect 8002 7046 8014 7098
rect 8066 7046 8078 7098
rect 8130 7046 8142 7098
rect 8194 7046 8206 7098
rect 8258 7046 13950 7098
rect 14002 7046 14014 7098
rect 14066 7046 14078 7098
rect 14130 7046 14142 7098
rect 14194 7046 14206 7098
rect 14258 7046 19950 7098
rect 20002 7046 20014 7098
rect 20066 7046 20078 7098
rect 20130 7046 20142 7098
rect 20194 7046 20206 7098
rect 20258 7046 25950 7098
rect 26002 7046 26014 7098
rect 26066 7046 26078 7098
rect 26130 7046 26142 7098
rect 26194 7046 26206 7098
rect 26258 7046 31950 7098
rect 32002 7046 32014 7098
rect 32066 7046 32078 7098
rect 32130 7046 32142 7098
rect 32194 7046 32206 7098
rect 32258 7046 37950 7098
rect 38002 7046 38014 7098
rect 38066 7046 38078 7098
rect 38130 7046 38142 7098
rect 38194 7046 38206 7098
rect 38258 7046 39836 7098
rect 1104 7024 39836 7046
rect 3786 6944 3792 6996
rect 3844 6984 3850 6996
rect 9674 6984 9680 6996
rect 3844 6956 9680 6984
rect 3844 6944 3850 6956
rect 9674 6944 9680 6956
rect 9732 6944 9738 6996
rect 9858 6944 9864 6996
rect 9916 6944 9922 6996
rect 13722 6944 13728 6996
rect 13780 6944 13786 6996
rect 18230 6984 18236 6996
rect 14476 6956 18236 6984
rect 12250 6876 12256 6928
rect 12308 6916 12314 6928
rect 14476 6916 14504 6956
rect 18230 6944 18236 6956
rect 18288 6944 18294 6996
rect 18322 6944 18328 6996
rect 18380 6984 18386 6996
rect 20622 6984 20628 6996
rect 18380 6956 20628 6984
rect 18380 6944 18386 6956
rect 20622 6944 20628 6956
rect 20680 6944 20686 6996
rect 21269 6987 21327 6993
rect 21269 6953 21281 6987
rect 21315 6984 21327 6987
rect 22002 6984 22008 6996
rect 21315 6956 22008 6984
rect 21315 6953 21327 6956
rect 21269 6947 21327 6953
rect 22002 6944 22008 6956
rect 22060 6944 22066 6996
rect 22462 6944 22468 6996
rect 22520 6984 22526 6996
rect 23014 6984 23020 6996
rect 22520 6956 23020 6984
rect 22520 6944 22526 6956
rect 23014 6944 23020 6956
rect 23072 6984 23078 6996
rect 23072 6956 24992 6984
rect 23072 6944 23078 6956
rect 12308 6888 14504 6916
rect 12308 6876 12314 6888
rect 16482 6876 16488 6928
rect 16540 6876 16546 6928
rect 16577 6919 16635 6925
rect 16577 6885 16589 6919
rect 16623 6885 16635 6919
rect 16577 6879 16635 6885
rect 22373 6919 22431 6925
rect 22373 6885 22385 6919
rect 22419 6916 22431 6919
rect 22554 6916 22560 6928
rect 22419 6888 22560 6916
rect 22419 6885 22431 6888
rect 22373 6879 22431 6885
rect 9766 6848 9772 6860
rect 3804 6820 9772 6848
rect 3804 6789 3832 6820
rect 9766 6808 9772 6820
rect 9824 6808 9830 6860
rect 15102 6808 15108 6860
rect 15160 6848 15166 6860
rect 15473 6851 15531 6857
rect 15473 6848 15485 6851
rect 15160 6820 15485 6848
rect 15160 6808 15166 6820
rect 15473 6817 15485 6820
rect 15519 6817 15531 6851
rect 15473 6811 15531 6817
rect 16298 6808 16304 6860
rect 16356 6848 16362 6860
rect 16592 6848 16620 6879
rect 22554 6876 22560 6888
rect 22612 6876 22618 6928
rect 24964 6916 24992 6956
rect 27338 6944 27344 6996
rect 27396 6984 27402 6996
rect 27396 6956 28856 6984
rect 27396 6944 27402 6956
rect 24964 6888 25084 6916
rect 16356 6820 16620 6848
rect 23477 6851 23535 6857
rect 16356 6808 16362 6820
rect 23477 6817 23489 6851
rect 23523 6848 23535 6851
rect 23658 6848 23664 6860
rect 23523 6820 23664 6848
rect 23523 6817 23535 6820
rect 23477 6811 23535 6817
rect 23658 6808 23664 6820
rect 23716 6848 23722 6860
rect 24486 6848 24492 6860
rect 23716 6820 24492 6848
rect 23716 6808 23722 6820
rect 24486 6808 24492 6820
rect 24544 6808 24550 6860
rect 3421 6783 3479 6789
rect 3421 6749 3433 6783
rect 3467 6780 3479 6783
rect 3789 6783 3847 6789
rect 3467 6752 3740 6780
rect 3467 6749 3479 6752
rect 3421 6743 3479 6749
rect 2774 6672 2780 6724
rect 2832 6712 2838 6724
rect 2869 6715 2927 6721
rect 2869 6712 2881 6715
rect 2832 6684 2881 6712
rect 2832 6672 2838 6684
rect 2869 6681 2881 6684
rect 2915 6681 2927 6715
rect 2869 6675 2927 6681
rect 3053 6715 3111 6721
rect 3053 6681 3065 6715
rect 3099 6712 3111 6715
rect 3510 6712 3516 6724
rect 3099 6684 3516 6712
rect 3099 6681 3111 6684
rect 3053 6675 3111 6681
rect 3510 6672 3516 6684
rect 3568 6672 3574 6724
rect 3712 6712 3740 6752
rect 3789 6749 3801 6783
rect 3835 6749 3847 6783
rect 3789 6743 3847 6749
rect 8570 6740 8576 6792
rect 8628 6780 8634 6792
rect 9125 6783 9183 6789
rect 9125 6780 9137 6783
rect 8628 6752 9137 6780
rect 8628 6740 8634 6752
rect 9125 6749 9137 6752
rect 9171 6749 9183 6783
rect 9125 6743 9183 6749
rect 9218 6783 9276 6789
rect 9218 6749 9230 6783
rect 9264 6749 9276 6783
rect 9218 6743 9276 6749
rect 9631 6783 9689 6789
rect 9631 6749 9643 6783
rect 9677 6780 9689 6783
rect 9858 6780 9864 6792
rect 9677 6752 9864 6780
rect 9677 6749 9689 6752
rect 9631 6743 9689 6749
rect 7834 6712 7840 6724
rect 3712 6684 7840 6712
rect 7834 6672 7840 6684
rect 7892 6672 7898 6724
rect 8754 6672 8760 6724
rect 8812 6712 8818 6724
rect 9232 6712 9260 6743
rect 9858 6740 9864 6752
rect 9916 6740 9922 6792
rect 10045 6783 10103 6789
rect 10045 6749 10057 6783
rect 10091 6780 10103 6783
rect 10318 6780 10324 6792
rect 10091 6752 10324 6780
rect 10091 6749 10103 6752
rect 10045 6743 10103 6749
rect 10318 6740 10324 6752
rect 10376 6740 10382 6792
rect 11422 6740 11428 6792
rect 11480 6780 11486 6792
rect 11977 6783 12035 6789
rect 11977 6780 11989 6783
rect 11480 6752 11989 6780
rect 11480 6740 11486 6752
rect 11977 6749 11989 6752
rect 12023 6780 12035 6783
rect 12250 6780 12256 6792
rect 12023 6752 12256 6780
rect 12023 6749 12035 6752
rect 11977 6743 12035 6749
rect 12250 6740 12256 6752
rect 12308 6740 12314 6792
rect 12986 6740 12992 6792
rect 13044 6780 13050 6792
rect 13814 6780 13820 6792
rect 13044 6752 13820 6780
rect 13044 6740 13050 6752
rect 13814 6740 13820 6752
rect 13872 6780 13878 6792
rect 13909 6783 13967 6789
rect 13909 6780 13921 6783
rect 13872 6752 13921 6780
rect 13872 6740 13878 6752
rect 13909 6749 13921 6752
rect 13955 6749 13967 6783
rect 14829 6783 14887 6789
rect 14829 6750 14841 6783
rect 13909 6743 13967 6749
rect 14752 6749 14841 6750
rect 14875 6749 14887 6783
rect 14752 6743 14887 6749
rect 8812 6684 9260 6712
rect 8812 6672 8818 6684
rect 9398 6672 9404 6724
rect 9456 6672 9462 6724
rect 9493 6715 9551 6721
rect 9493 6681 9505 6715
rect 9539 6681 9551 6715
rect 9493 6675 9551 6681
rect 3605 6647 3663 6653
rect 3605 6613 3617 6647
rect 3651 6644 3663 6647
rect 3694 6644 3700 6656
rect 3651 6616 3700 6644
rect 3651 6613 3663 6616
rect 3605 6607 3663 6613
rect 3694 6604 3700 6616
rect 3752 6604 3758 6656
rect 3970 6604 3976 6656
rect 4028 6604 4034 6656
rect 9508 6644 9536 6675
rect 12158 6672 12164 6724
rect 12216 6712 12222 6724
rect 14752 6722 14872 6743
rect 15378 6740 15384 6792
rect 15436 6780 15442 6792
rect 15749 6783 15807 6789
rect 15749 6780 15761 6783
rect 15436 6752 15761 6780
rect 15436 6740 15442 6752
rect 15749 6749 15761 6752
rect 15795 6749 15807 6783
rect 15749 6743 15807 6749
rect 15838 6740 15844 6792
rect 15896 6780 15902 6792
rect 17313 6783 17371 6789
rect 17313 6780 17325 6783
rect 15896 6752 17325 6780
rect 15896 6740 15902 6752
rect 17313 6749 17325 6752
rect 17359 6749 17371 6783
rect 17313 6743 17371 6749
rect 17589 6783 17647 6789
rect 17589 6749 17601 6783
rect 17635 6749 17647 6783
rect 17589 6743 17647 6749
rect 19981 6783 20039 6789
rect 19981 6749 19993 6783
rect 20027 6780 20039 6783
rect 20162 6780 20168 6792
rect 20027 6752 20168 6780
rect 20027 6749 20039 6752
rect 19981 6743 20039 6749
rect 14752 6712 14780 6722
rect 12216 6684 14780 6712
rect 12216 6672 12222 6684
rect 15102 6672 15108 6724
rect 15160 6712 15166 6724
rect 17604 6712 17632 6743
rect 20162 6740 20168 6752
rect 20220 6740 20226 6792
rect 20257 6783 20315 6789
rect 20257 6749 20269 6783
rect 20303 6749 20315 6783
rect 20257 6743 20315 6749
rect 17678 6712 17684 6724
rect 15160 6684 17684 6712
rect 15160 6672 15166 6684
rect 17678 6672 17684 6684
rect 17736 6712 17742 6724
rect 20272 6712 20300 6743
rect 20530 6740 20536 6792
rect 20588 6740 20594 6792
rect 21361 6783 21419 6789
rect 21361 6749 21373 6783
rect 21407 6749 21419 6783
rect 21361 6743 21419 6749
rect 21637 6783 21695 6789
rect 21637 6749 21649 6783
rect 21683 6780 21695 6783
rect 21726 6780 21732 6792
rect 21683 6752 21732 6780
rect 21683 6749 21695 6752
rect 21637 6743 21695 6749
rect 20438 6712 20444 6724
rect 17736 6684 20444 6712
rect 17736 6672 17742 6684
rect 20438 6672 20444 6684
rect 20496 6712 20502 6724
rect 21376 6712 21404 6743
rect 21726 6740 21732 6752
rect 21784 6740 21790 6792
rect 23106 6740 23112 6792
rect 23164 6780 23170 6792
rect 23201 6783 23259 6789
rect 23201 6780 23213 6783
rect 23164 6752 23213 6780
rect 23164 6740 23170 6752
rect 23201 6749 23213 6752
rect 23247 6749 23259 6783
rect 24857 6783 24915 6789
rect 24857 6780 24869 6783
rect 23201 6743 23259 6749
rect 23308 6752 24869 6780
rect 22646 6712 22652 6724
rect 20496 6684 22652 6712
rect 20496 6672 20502 6684
rect 22646 6672 22652 6684
rect 22704 6672 22710 6724
rect 9582 6644 9588 6656
rect 9508 6616 9588 6644
rect 9582 6604 9588 6616
rect 9640 6604 9646 6656
rect 9769 6647 9827 6653
rect 9769 6613 9781 6647
rect 9815 6644 9827 6647
rect 10042 6644 10048 6656
rect 9815 6616 10048 6644
rect 9815 6613 9827 6616
rect 9769 6607 9827 6613
rect 10042 6604 10048 6616
rect 10100 6604 10106 6656
rect 11606 6604 11612 6656
rect 11664 6644 11670 6656
rect 11793 6647 11851 6653
rect 11793 6644 11805 6647
rect 11664 6616 11805 6644
rect 11664 6604 11670 6616
rect 11793 6613 11805 6616
rect 11839 6613 11851 6647
rect 11793 6607 11851 6613
rect 13814 6604 13820 6656
rect 13872 6644 13878 6656
rect 14093 6647 14151 6653
rect 14093 6644 14105 6647
rect 13872 6616 14105 6644
rect 13872 6604 13878 6616
rect 14093 6613 14105 6616
rect 14139 6613 14151 6647
rect 14093 6607 14151 6613
rect 14182 6604 14188 6656
rect 14240 6644 14246 6656
rect 15470 6644 15476 6656
rect 14240 6616 15476 6644
rect 14240 6604 14246 6616
rect 15470 6604 15476 6616
rect 15528 6644 15534 6656
rect 16022 6644 16028 6656
rect 15528 6616 16028 6644
rect 15528 6604 15534 6616
rect 16022 6604 16028 6616
rect 16080 6604 16086 6656
rect 16206 6604 16212 6656
rect 16264 6644 16270 6656
rect 19334 6644 19340 6656
rect 16264 6616 19340 6644
rect 16264 6604 16270 6616
rect 19334 6604 19340 6616
rect 19392 6604 19398 6656
rect 20165 6647 20223 6653
rect 20165 6613 20177 6647
rect 20211 6644 20223 6647
rect 20898 6644 20904 6656
rect 20211 6616 20904 6644
rect 20211 6613 20223 6616
rect 20165 6607 20223 6613
rect 20898 6604 20904 6616
rect 20956 6604 20962 6656
rect 21269 6647 21327 6653
rect 21269 6613 21281 6647
rect 21315 6644 21327 6647
rect 21450 6644 21456 6656
rect 21315 6616 21456 6644
rect 21315 6613 21327 6616
rect 21269 6607 21327 6613
rect 21450 6604 21456 6616
rect 21508 6604 21514 6656
rect 22462 6604 22468 6656
rect 22520 6604 22526 6656
rect 22830 6604 22836 6656
rect 22888 6644 22894 6656
rect 23308 6644 23336 6752
rect 24857 6749 24869 6752
rect 24903 6749 24915 6783
rect 25056 6780 25084 6888
rect 25590 6876 25596 6928
rect 25648 6916 25654 6928
rect 25648 6888 27568 6916
rect 25648 6876 25654 6888
rect 26418 6808 26424 6860
rect 26476 6848 26482 6860
rect 26476 6820 27476 6848
rect 26476 6808 26482 6820
rect 25317 6783 25375 6789
rect 25317 6780 25329 6783
rect 25056 6752 25329 6780
rect 24857 6743 24915 6749
rect 25317 6749 25329 6752
rect 25363 6749 25375 6783
rect 25317 6743 25375 6749
rect 27341 6783 27399 6789
rect 27341 6749 27353 6783
rect 27387 6749 27399 6783
rect 27341 6743 27399 6749
rect 23566 6672 23572 6724
rect 23624 6712 23630 6724
rect 27356 6712 27384 6743
rect 23624 6684 27384 6712
rect 27448 6712 27476 6820
rect 27540 6780 27568 6888
rect 27706 6876 27712 6928
rect 27764 6876 27770 6928
rect 28828 6848 28856 6956
rect 30374 6944 30380 6996
rect 30432 6984 30438 6996
rect 37550 6984 37556 6996
rect 30432 6956 37556 6984
rect 30432 6944 30438 6956
rect 37550 6944 37556 6956
rect 37608 6944 37614 6996
rect 28994 6876 29000 6928
rect 29052 6916 29058 6928
rect 37642 6916 37648 6928
rect 29052 6888 37648 6916
rect 29052 6876 29058 6888
rect 37642 6876 37648 6888
rect 37700 6876 37706 6928
rect 28828 6820 29316 6848
rect 27617 6783 27675 6789
rect 27617 6780 27629 6783
rect 27540 6752 27629 6780
rect 27617 6749 27629 6752
rect 27663 6749 27675 6783
rect 27617 6743 27675 6749
rect 27890 6740 27896 6792
rect 27948 6740 27954 6792
rect 28166 6740 28172 6792
rect 28224 6740 28230 6792
rect 28442 6740 28448 6792
rect 28500 6740 28506 6792
rect 28721 6783 28779 6789
rect 28721 6749 28733 6783
rect 28767 6749 28779 6783
rect 28721 6743 28779 6749
rect 28736 6712 28764 6743
rect 28994 6740 29000 6792
rect 29052 6740 29058 6792
rect 29288 6789 29316 6820
rect 31846 6808 31852 6860
rect 31904 6848 31910 6860
rect 31904 6820 32260 6848
rect 31904 6808 31910 6820
rect 29273 6783 29331 6789
rect 29273 6749 29285 6783
rect 29319 6749 29331 6783
rect 29273 6743 29331 6749
rect 29730 6740 29736 6792
rect 29788 6740 29794 6792
rect 30006 6740 30012 6792
rect 30064 6740 30070 6792
rect 31386 6740 31392 6792
rect 31444 6780 31450 6792
rect 32232 6789 32260 6820
rect 37090 6808 37096 6860
rect 37148 6848 37154 6860
rect 37737 6851 37795 6857
rect 37737 6848 37749 6851
rect 37148 6820 37749 6848
rect 37148 6808 37154 6820
rect 37737 6817 37749 6820
rect 37783 6817 37795 6851
rect 37737 6811 37795 6817
rect 38286 6808 38292 6860
rect 38344 6848 38350 6860
rect 39022 6848 39028 6860
rect 38344 6820 39028 6848
rect 38344 6808 38350 6820
rect 39022 6808 39028 6820
rect 39080 6808 39086 6860
rect 31941 6783 31999 6789
rect 31941 6780 31953 6783
rect 31444 6752 31953 6780
rect 31444 6740 31450 6752
rect 31941 6749 31953 6752
rect 31987 6749 31999 6783
rect 31941 6743 31999 6749
rect 32217 6783 32275 6789
rect 32217 6749 32229 6783
rect 32263 6749 32275 6783
rect 32217 6743 32275 6749
rect 32398 6740 32404 6792
rect 32456 6740 32462 6792
rect 32677 6783 32735 6789
rect 32677 6749 32689 6783
rect 32723 6749 32735 6783
rect 32677 6743 32735 6749
rect 37829 6783 37887 6789
rect 37829 6749 37841 6783
rect 37875 6780 37887 6783
rect 37921 6783 37979 6789
rect 37921 6780 37933 6783
rect 37875 6752 37933 6780
rect 37875 6749 37887 6752
rect 37829 6743 37887 6749
rect 37921 6749 37933 6752
rect 37967 6749 37979 6783
rect 37921 6743 37979 6749
rect 27448 6684 28764 6712
rect 23624 6672 23630 6684
rect 29178 6672 29184 6724
rect 29236 6712 29242 6724
rect 32692 6712 32720 6743
rect 38470 6740 38476 6792
rect 38528 6740 38534 6792
rect 38746 6740 38752 6792
rect 38804 6780 38810 6792
rect 38841 6783 38899 6789
rect 38841 6780 38853 6783
rect 38804 6752 38853 6780
rect 38804 6740 38810 6752
rect 38841 6749 38853 6752
rect 38887 6749 38899 6783
rect 39209 6783 39267 6789
rect 39209 6780 39221 6783
rect 38841 6743 38899 6749
rect 38948 6752 39221 6780
rect 35618 6712 35624 6724
rect 29236 6684 32720 6712
rect 32784 6684 35624 6712
rect 29236 6672 29242 6684
rect 22888 6616 23336 6644
rect 22888 6604 22894 6616
rect 24670 6604 24676 6656
rect 24728 6604 24734 6656
rect 25130 6604 25136 6656
rect 25188 6604 25194 6656
rect 26786 6604 26792 6656
rect 26844 6644 26850 6656
rect 27157 6647 27215 6653
rect 27157 6644 27169 6647
rect 26844 6616 27169 6644
rect 26844 6604 26850 6616
rect 27157 6613 27169 6616
rect 27203 6613 27215 6647
rect 27157 6607 27215 6613
rect 27246 6604 27252 6656
rect 27304 6644 27310 6656
rect 27433 6647 27491 6653
rect 27433 6644 27445 6647
rect 27304 6616 27445 6644
rect 27304 6604 27310 6616
rect 27433 6613 27445 6616
rect 27479 6613 27491 6647
rect 27433 6607 27491 6613
rect 27982 6604 27988 6656
rect 28040 6604 28046 6656
rect 28258 6604 28264 6656
rect 28316 6604 28322 6656
rect 28534 6604 28540 6656
rect 28592 6604 28598 6656
rect 28718 6604 28724 6656
rect 28776 6644 28782 6656
rect 28813 6647 28871 6653
rect 28813 6644 28825 6647
rect 28776 6616 28825 6644
rect 28776 6604 28782 6616
rect 28813 6613 28825 6616
rect 28859 6613 28871 6647
rect 28813 6607 28871 6613
rect 28902 6604 28908 6656
rect 28960 6644 28966 6656
rect 29089 6647 29147 6653
rect 29089 6644 29101 6647
rect 28960 6616 29101 6644
rect 28960 6604 28966 6616
rect 29089 6613 29101 6616
rect 29135 6613 29147 6647
rect 29089 6607 29147 6613
rect 29362 6604 29368 6656
rect 29420 6644 29426 6656
rect 29549 6647 29607 6653
rect 29549 6644 29561 6647
rect 29420 6616 29561 6644
rect 29420 6604 29426 6616
rect 29549 6613 29561 6616
rect 29595 6613 29607 6647
rect 29549 6607 29607 6613
rect 29822 6604 29828 6656
rect 29880 6604 29886 6656
rect 31478 6604 31484 6656
rect 31536 6644 31542 6656
rect 31757 6647 31815 6653
rect 31757 6644 31769 6647
rect 31536 6616 31769 6644
rect 31536 6604 31542 6616
rect 31757 6613 31769 6616
rect 31803 6613 31815 6647
rect 31757 6607 31815 6613
rect 31846 6604 31852 6656
rect 31904 6644 31910 6656
rect 32033 6647 32091 6653
rect 32033 6644 32045 6647
rect 31904 6616 32045 6644
rect 31904 6604 31910 6616
rect 32033 6613 32045 6616
rect 32079 6613 32091 6647
rect 32033 6607 32091 6613
rect 32585 6647 32643 6653
rect 32585 6613 32597 6647
rect 32631 6644 32643 6647
rect 32784 6644 32812 6684
rect 35618 6672 35624 6684
rect 35676 6672 35682 6724
rect 32631 6616 32812 6644
rect 32861 6647 32919 6653
rect 32631 6613 32643 6616
rect 32585 6607 32643 6613
rect 32861 6613 32873 6647
rect 32907 6644 32919 6647
rect 34698 6644 34704 6656
rect 32907 6616 34704 6644
rect 32907 6613 32919 6616
rect 32861 6607 32919 6613
rect 34698 6604 34704 6616
rect 34756 6604 34762 6656
rect 38105 6647 38163 6653
rect 38105 6613 38117 6647
rect 38151 6644 38163 6647
rect 38562 6644 38568 6656
rect 38151 6616 38568 6644
rect 38151 6613 38163 6616
rect 38105 6607 38163 6613
rect 38562 6604 38568 6616
rect 38620 6604 38626 6656
rect 38654 6604 38660 6656
rect 38712 6604 38718 6656
rect 38838 6604 38844 6656
rect 38896 6644 38902 6656
rect 38948 6644 38976 6752
rect 39209 6749 39221 6752
rect 39255 6749 39267 6783
rect 39209 6743 39267 6749
rect 39574 6712 39580 6724
rect 39040 6684 39580 6712
rect 39040 6653 39068 6684
rect 39574 6672 39580 6684
rect 39632 6672 39638 6724
rect 38896 6616 38976 6644
rect 39025 6647 39083 6653
rect 38896 6604 38902 6616
rect 39025 6613 39037 6647
rect 39071 6613 39083 6647
rect 39025 6607 39083 6613
rect 39390 6604 39396 6656
rect 39448 6604 39454 6656
rect 1104 6554 39836 6576
rect 1104 6502 3010 6554
rect 3062 6502 3074 6554
rect 3126 6502 3138 6554
rect 3190 6502 3202 6554
rect 3254 6502 3266 6554
rect 3318 6502 9010 6554
rect 9062 6502 9074 6554
rect 9126 6502 9138 6554
rect 9190 6502 9202 6554
rect 9254 6502 9266 6554
rect 9318 6502 15010 6554
rect 15062 6502 15074 6554
rect 15126 6502 15138 6554
rect 15190 6502 15202 6554
rect 15254 6502 15266 6554
rect 15318 6502 21010 6554
rect 21062 6502 21074 6554
rect 21126 6502 21138 6554
rect 21190 6502 21202 6554
rect 21254 6502 21266 6554
rect 21318 6502 27010 6554
rect 27062 6502 27074 6554
rect 27126 6502 27138 6554
rect 27190 6502 27202 6554
rect 27254 6502 27266 6554
rect 27318 6502 33010 6554
rect 33062 6502 33074 6554
rect 33126 6502 33138 6554
rect 33190 6502 33202 6554
rect 33254 6502 33266 6554
rect 33318 6502 39010 6554
rect 39062 6502 39074 6554
rect 39126 6502 39138 6554
rect 39190 6502 39202 6554
rect 39254 6502 39266 6554
rect 39318 6502 39836 6554
rect 1104 6480 39836 6502
rect 7561 6443 7619 6449
rect 7561 6409 7573 6443
rect 7607 6440 7619 6443
rect 8294 6440 8300 6452
rect 7607 6412 8300 6440
rect 7607 6409 7619 6412
rect 7561 6403 7619 6409
rect 8294 6400 8300 6412
rect 8352 6400 8358 6452
rect 8662 6400 8668 6452
rect 8720 6440 8726 6452
rect 8938 6440 8944 6452
rect 8720 6412 8944 6440
rect 8720 6400 8726 6412
rect 8938 6400 8944 6412
rect 8996 6400 9002 6452
rect 9122 6400 9128 6452
rect 9180 6440 9186 6452
rect 11793 6443 11851 6449
rect 9180 6412 9674 6440
rect 9180 6400 9186 6412
rect 9646 6372 9674 6412
rect 11793 6409 11805 6443
rect 11839 6440 11851 6443
rect 11882 6440 11888 6452
rect 11839 6412 11888 6440
rect 11839 6409 11851 6412
rect 11793 6403 11851 6409
rect 11882 6400 11888 6412
rect 11940 6400 11946 6452
rect 11974 6400 11980 6452
rect 12032 6440 12038 6452
rect 12805 6443 12863 6449
rect 12805 6440 12817 6443
rect 12032 6412 12817 6440
rect 12032 6400 12038 6412
rect 12805 6409 12817 6412
rect 12851 6409 12863 6443
rect 12805 6403 12863 6409
rect 13262 6400 13268 6452
rect 13320 6440 13326 6452
rect 13320 6412 15700 6440
rect 13320 6400 13326 6412
rect 14642 6372 14648 6384
rect 9646 6344 14648 6372
rect 14642 6332 14648 6344
rect 14700 6332 14706 6384
rect 14829 6375 14887 6381
rect 14829 6341 14841 6375
rect 14875 6372 14887 6375
rect 15378 6372 15384 6384
rect 14875 6344 15384 6372
rect 14875 6341 14887 6344
rect 14829 6335 14887 6341
rect 15378 6332 15384 6344
rect 15436 6332 15442 6384
rect 15672 6372 15700 6412
rect 15746 6400 15752 6452
rect 15804 6440 15810 6452
rect 15933 6443 15991 6449
rect 15933 6440 15945 6443
rect 15804 6412 15945 6440
rect 15804 6400 15810 6412
rect 15933 6409 15945 6412
rect 15979 6409 15991 6443
rect 20441 6443 20499 6449
rect 15933 6403 15991 6409
rect 16592 6412 20024 6440
rect 16592 6372 16620 6412
rect 15672 6344 16620 6372
rect 7377 6307 7435 6313
rect 7377 6273 7389 6307
rect 7423 6304 7435 6307
rect 8662 6304 8668 6316
rect 7423 6276 8668 6304
rect 7423 6273 7435 6276
rect 7377 6267 7435 6273
rect 8662 6264 8668 6276
rect 8720 6264 8726 6316
rect 8938 6264 8944 6316
rect 8996 6304 9002 6316
rect 8996 6276 9996 6304
rect 8996 6264 9002 6276
rect 3878 6196 3884 6248
rect 3936 6236 3942 6248
rect 9214 6236 9220 6248
rect 3936 6208 9220 6236
rect 3936 6196 3942 6208
rect 9214 6196 9220 6208
rect 9272 6196 9278 6248
rect 9490 6196 9496 6248
rect 9548 6236 9554 6248
rect 9769 6239 9827 6245
rect 9769 6236 9781 6239
rect 9548 6208 9781 6236
rect 9548 6196 9554 6208
rect 9769 6205 9781 6208
rect 9815 6205 9827 6239
rect 9968 6236 9996 6276
rect 10042 6264 10048 6316
rect 10100 6264 10106 6316
rect 11514 6264 11520 6316
rect 11572 6304 11578 6316
rect 11609 6307 11667 6313
rect 11609 6304 11621 6307
rect 11572 6276 11621 6304
rect 11572 6264 11578 6276
rect 11609 6273 11621 6276
rect 11655 6304 11667 6307
rect 12526 6304 12532 6316
rect 11655 6276 12532 6304
rect 11655 6273 11667 6276
rect 11609 6267 11667 6273
rect 12526 6264 12532 6276
rect 12584 6264 12590 6316
rect 12989 6307 13047 6313
rect 12989 6273 13001 6307
rect 13035 6273 13047 6307
rect 12989 6267 13047 6273
rect 12158 6236 12164 6248
rect 9968 6208 12164 6236
rect 9769 6199 9827 6205
rect 12158 6196 12164 6208
rect 12216 6196 12222 6248
rect 13004 6236 13032 6267
rect 14090 6264 14096 6316
rect 14148 6304 14154 6316
rect 14461 6307 14519 6313
rect 14461 6304 14473 6307
rect 14148 6276 14473 6304
rect 14148 6264 14154 6276
rect 14461 6273 14473 6276
rect 14507 6273 14519 6307
rect 14461 6267 14519 6273
rect 14550 6264 14556 6316
rect 14608 6304 14614 6316
rect 14608 6276 14653 6304
rect 14608 6264 14614 6276
rect 14734 6264 14740 6316
rect 14792 6264 14798 6316
rect 14967 6307 15025 6313
rect 14967 6273 14979 6307
rect 15013 6304 15025 6307
rect 16022 6304 16028 6316
rect 15013 6276 16028 6304
rect 15013 6273 15025 6276
rect 14967 6267 15025 6273
rect 16022 6264 16028 6276
rect 16080 6264 16086 6316
rect 16117 6307 16175 6313
rect 16117 6273 16129 6307
rect 16163 6304 16175 6307
rect 16206 6304 16212 6316
rect 16163 6276 16212 6304
rect 16163 6273 16175 6276
rect 16117 6267 16175 6273
rect 16206 6264 16212 6276
rect 16264 6264 16270 6316
rect 17405 6307 17463 6313
rect 17405 6304 17417 6307
rect 16316 6276 17417 6304
rect 14182 6236 14188 6248
rect 13004 6208 14188 6236
rect 14182 6196 14188 6208
rect 14240 6196 14246 6248
rect 14274 6196 14280 6248
rect 14332 6236 14338 6248
rect 16316 6236 16344 6276
rect 17405 6273 17417 6276
rect 17451 6273 17463 6307
rect 17405 6267 17463 6273
rect 17678 6264 17684 6316
rect 17736 6264 17742 6316
rect 17954 6264 17960 6316
rect 18012 6264 18018 6316
rect 19153 6307 19211 6313
rect 19153 6273 19165 6307
rect 19199 6273 19211 6307
rect 19153 6267 19211 6273
rect 14332 6208 16344 6236
rect 19168 6236 19196 6267
rect 19242 6264 19248 6316
rect 19300 6304 19306 6316
rect 19610 6304 19616 6316
rect 19300 6276 19616 6304
rect 19300 6264 19306 6276
rect 19610 6264 19616 6276
rect 19668 6304 19674 6316
rect 19705 6307 19763 6313
rect 19705 6304 19717 6307
rect 19668 6276 19717 6304
rect 19668 6264 19674 6276
rect 19705 6273 19717 6276
rect 19751 6273 19763 6307
rect 19996 6304 20024 6412
rect 20441 6409 20453 6443
rect 20487 6440 20499 6443
rect 20990 6440 20996 6452
rect 20487 6412 20996 6440
rect 20487 6409 20499 6412
rect 20441 6403 20499 6409
rect 20990 6400 20996 6412
rect 21048 6400 21054 6452
rect 22094 6400 22100 6452
rect 22152 6440 22158 6452
rect 38470 6440 38476 6452
rect 22152 6412 38476 6440
rect 22152 6400 22158 6412
rect 38470 6400 38476 6412
rect 38528 6400 38534 6452
rect 39393 6443 39451 6449
rect 39393 6409 39405 6443
rect 39439 6440 39451 6443
rect 40034 6440 40040 6452
rect 39439 6412 40040 6440
rect 39439 6409 39451 6412
rect 39393 6403 39451 6409
rect 40034 6400 40040 6412
rect 40092 6400 40098 6452
rect 21008 6372 21036 6400
rect 23842 6372 23848 6384
rect 21008 6344 21772 6372
rect 21744 6334 21772 6344
rect 22342 6344 23848 6372
rect 20438 6304 20444 6316
rect 19996 6276 20444 6304
rect 19705 6267 19763 6273
rect 20438 6264 20444 6276
rect 20496 6304 20502 6316
rect 21744 6313 21864 6334
rect 21269 6307 21327 6313
rect 21269 6304 21281 6307
rect 20496 6276 21281 6304
rect 20496 6264 20502 6276
rect 21269 6273 21281 6276
rect 21315 6273 21327 6307
rect 21744 6307 21879 6313
rect 21744 6306 21833 6307
rect 21269 6267 21327 6273
rect 21821 6273 21833 6306
rect 21867 6273 21879 6307
rect 21821 6267 21879 6273
rect 21910 6264 21916 6316
rect 21968 6304 21974 6316
rect 21968 6276 22013 6304
rect 21968 6264 21974 6276
rect 22094 6264 22100 6316
rect 22152 6264 22158 6316
rect 22186 6264 22192 6316
rect 22244 6264 22250 6316
rect 22342 6313 22370 6344
rect 23842 6332 23848 6344
rect 23900 6332 23906 6384
rect 26694 6332 26700 6384
rect 26752 6372 26758 6384
rect 28994 6372 29000 6384
rect 26752 6344 29000 6372
rect 26752 6332 26758 6344
rect 28994 6332 29000 6344
rect 29052 6332 29058 6384
rect 31846 6332 31852 6384
rect 31904 6372 31910 6384
rect 38746 6372 38752 6384
rect 31904 6344 38752 6372
rect 31904 6332 31910 6344
rect 38746 6332 38752 6344
rect 38804 6332 38810 6384
rect 22327 6307 22385 6313
rect 22327 6273 22339 6307
rect 22373 6273 22385 6307
rect 22327 6267 22385 6273
rect 22833 6307 22891 6313
rect 22833 6273 22845 6307
rect 22879 6273 22891 6307
rect 22833 6267 22891 6273
rect 19426 6236 19432 6248
rect 19168 6208 19432 6236
rect 14332 6196 14338 6208
rect 19426 6196 19432 6208
rect 19484 6196 19490 6248
rect 20530 6236 20536 6248
rect 20088 6208 20536 6236
rect 5534 6128 5540 6180
rect 5592 6168 5598 6180
rect 10229 6171 10287 6177
rect 10229 6168 10241 6171
rect 5592 6140 10241 6168
rect 5592 6128 5598 6140
rect 10229 6137 10241 6140
rect 10275 6137 10287 6171
rect 15838 6168 15844 6180
rect 10229 6131 10287 6137
rect 12406 6140 15844 6168
rect 7742 6060 7748 6112
rect 7800 6100 7806 6112
rect 9861 6103 9919 6109
rect 9861 6100 9873 6103
rect 7800 6072 9873 6100
rect 7800 6060 7806 6072
rect 9861 6069 9873 6072
rect 9907 6069 9919 6103
rect 9861 6063 9919 6069
rect 10042 6060 10048 6112
rect 10100 6100 10106 6112
rect 12406 6100 12434 6140
rect 15838 6128 15844 6140
rect 15896 6128 15902 6180
rect 18966 6128 18972 6180
rect 19024 6168 19030 6180
rect 19337 6171 19395 6177
rect 19337 6168 19349 6171
rect 19024 6140 19349 6168
rect 19024 6128 19030 6140
rect 19337 6137 19349 6140
rect 19383 6137 19395 6171
rect 19337 6131 19395 6137
rect 10100 6072 12434 6100
rect 10100 6060 10106 6072
rect 12526 6060 12532 6112
rect 12584 6100 12590 6112
rect 13722 6100 13728 6112
rect 12584 6072 13728 6100
rect 12584 6060 12590 6072
rect 13722 6060 13728 6072
rect 13780 6060 13786 6112
rect 14642 6060 14648 6112
rect 14700 6100 14706 6112
rect 15105 6103 15163 6109
rect 15105 6100 15117 6103
rect 14700 6072 15117 6100
rect 14700 6060 14706 6072
rect 15105 6069 15117 6072
rect 15151 6069 15163 6103
rect 15105 6063 15163 6069
rect 16390 6060 16396 6112
rect 16448 6100 16454 6112
rect 16669 6103 16727 6109
rect 16669 6100 16681 6103
rect 16448 6072 16681 6100
rect 16448 6060 16454 6072
rect 16669 6069 16681 6072
rect 16715 6069 16727 6103
rect 16669 6063 16727 6069
rect 17678 6060 17684 6112
rect 17736 6100 17742 6112
rect 17773 6103 17831 6109
rect 17773 6100 17785 6103
rect 17736 6072 17785 6100
rect 17736 6060 17742 6072
rect 17773 6069 17785 6072
rect 17819 6069 17831 6103
rect 17773 6063 17831 6069
rect 17862 6060 17868 6112
rect 17920 6100 17926 6112
rect 20088 6100 20116 6208
rect 20530 6196 20536 6208
rect 20588 6196 20594 6248
rect 21545 6239 21603 6245
rect 21545 6205 21557 6239
rect 21591 6236 21603 6239
rect 22646 6236 22652 6248
rect 21591 6208 22652 6236
rect 21591 6205 21603 6208
rect 21545 6199 21603 6205
rect 22646 6196 22652 6208
rect 22704 6196 22710 6248
rect 22465 6171 22523 6177
rect 22465 6137 22477 6171
rect 22511 6168 22523 6171
rect 22848 6168 22876 6267
rect 23750 6264 23756 6316
rect 23808 6304 23814 6316
rect 26510 6304 26516 6316
rect 23808 6276 26516 6304
rect 23808 6264 23814 6276
rect 26510 6264 26516 6276
rect 26568 6264 26574 6316
rect 27430 6264 27436 6316
rect 27488 6304 27494 6316
rect 29730 6304 29736 6316
rect 27488 6276 29736 6304
rect 27488 6264 27494 6276
rect 29730 6264 29736 6276
rect 29788 6264 29794 6316
rect 31386 6264 31392 6316
rect 31444 6304 31450 6316
rect 34977 6307 35035 6313
rect 34977 6304 34989 6307
rect 31444 6276 34989 6304
rect 31444 6264 31450 6276
rect 34977 6273 34989 6276
rect 35023 6273 35035 6307
rect 34977 6267 35035 6273
rect 37458 6264 37464 6316
rect 37516 6304 37522 6316
rect 37737 6307 37795 6313
rect 37737 6304 37749 6307
rect 37516 6276 37749 6304
rect 37516 6264 37522 6276
rect 37737 6273 37749 6276
rect 37783 6304 37795 6307
rect 37921 6307 37979 6313
rect 37921 6304 37933 6307
rect 37783 6276 37933 6304
rect 37783 6273 37795 6276
rect 37737 6267 37795 6273
rect 37921 6273 37933 6276
rect 37967 6273 37979 6307
rect 37921 6267 37979 6273
rect 38841 6307 38899 6313
rect 38841 6273 38853 6307
rect 38887 6273 38899 6307
rect 38841 6267 38899 6273
rect 23106 6196 23112 6248
rect 23164 6196 23170 6248
rect 23934 6196 23940 6248
rect 23992 6236 23998 6248
rect 24762 6236 24768 6248
rect 23992 6208 24768 6236
rect 23992 6196 23998 6208
rect 24762 6196 24768 6208
rect 24820 6236 24826 6248
rect 24820 6208 27476 6236
rect 24820 6196 24826 6208
rect 22511 6140 22876 6168
rect 27448 6168 27476 6208
rect 27522 6196 27528 6248
rect 27580 6236 27586 6248
rect 30006 6236 30012 6248
rect 27580 6208 30012 6236
rect 27580 6196 27586 6208
rect 30006 6196 30012 6208
rect 30064 6196 30070 6248
rect 35250 6196 35256 6248
rect 35308 6236 35314 6248
rect 38856 6236 38884 6267
rect 39206 6264 39212 6316
rect 39264 6264 39270 6316
rect 35308 6208 38884 6236
rect 35308 6196 35314 6208
rect 28166 6168 28172 6180
rect 27448 6140 28172 6168
rect 22511 6137 22523 6140
rect 22465 6131 22523 6137
rect 28166 6128 28172 6140
rect 28224 6128 28230 6180
rect 35161 6171 35219 6177
rect 35161 6137 35173 6171
rect 35207 6168 35219 6171
rect 35802 6168 35808 6180
rect 35207 6140 35808 6168
rect 35207 6137 35219 6140
rect 35161 6131 35219 6137
rect 35802 6128 35808 6140
rect 35860 6128 35866 6180
rect 17920 6072 20116 6100
rect 17920 6060 17926 6072
rect 20530 6060 20536 6112
rect 20588 6060 20594 6112
rect 22278 6060 22284 6112
rect 22336 6100 22342 6112
rect 22649 6103 22707 6109
rect 22649 6100 22661 6103
rect 22336 6072 22661 6100
rect 22336 6060 22342 6072
rect 22649 6069 22661 6072
rect 22695 6069 22707 6103
rect 22649 6063 22707 6069
rect 23014 6060 23020 6112
rect 23072 6060 23078 6112
rect 23474 6060 23480 6112
rect 23532 6100 23538 6112
rect 24670 6100 24676 6112
rect 23532 6072 24676 6100
rect 23532 6060 23538 6072
rect 24670 6060 24676 6072
rect 24728 6060 24734 6112
rect 30374 6060 30380 6112
rect 30432 6100 30438 6112
rect 37274 6100 37280 6112
rect 30432 6072 37280 6100
rect 30432 6060 30438 6072
rect 37274 6060 37280 6072
rect 37332 6060 37338 6112
rect 38105 6103 38163 6109
rect 38105 6069 38117 6103
rect 38151 6100 38163 6103
rect 38654 6100 38660 6112
rect 38151 6072 38660 6100
rect 38151 6069 38163 6072
rect 38105 6063 38163 6069
rect 38654 6060 38660 6072
rect 38712 6060 38718 6112
rect 39022 6060 39028 6112
rect 39080 6060 39086 6112
rect 1104 6010 39836 6032
rect 1104 5958 1950 6010
rect 2002 5958 2014 6010
rect 2066 5958 2078 6010
rect 2130 5958 2142 6010
rect 2194 5958 2206 6010
rect 2258 5958 7950 6010
rect 8002 5958 8014 6010
rect 8066 5958 8078 6010
rect 8130 5958 8142 6010
rect 8194 5958 8206 6010
rect 8258 5958 13950 6010
rect 14002 5958 14014 6010
rect 14066 5958 14078 6010
rect 14130 5958 14142 6010
rect 14194 5958 14206 6010
rect 14258 5958 19950 6010
rect 20002 5958 20014 6010
rect 20066 5958 20078 6010
rect 20130 5958 20142 6010
rect 20194 5958 20206 6010
rect 20258 5958 25950 6010
rect 26002 5958 26014 6010
rect 26066 5958 26078 6010
rect 26130 5958 26142 6010
rect 26194 5958 26206 6010
rect 26258 5958 31950 6010
rect 32002 5958 32014 6010
rect 32066 5958 32078 6010
rect 32130 5958 32142 6010
rect 32194 5958 32206 6010
rect 32258 5958 37950 6010
rect 38002 5958 38014 6010
rect 38066 5958 38078 6010
rect 38130 5958 38142 6010
rect 38194 5958 38206 6010
rect 38258 5958 39836 6010
rect 1104 5936 39836 5958
rect 7374 5896 7380 5908
rect 3896 5868 7380 5896
rect 3789 5695 3847 5701
rect 3789 5661 3801 5695
rect 3835 5692 3847 5695
rect 3896 5692 3924 5868
rect 7374 5856 7380 5868
rect 7432 5856 7438 5908
rect 7653 5899 7711 5905
rect 7653 5865 7665 5899
rect 7699 5896 7711 5899
rect 8478 5896 8484 5908
rect 7699 5868 8484 5896
rect 7699 5865 7711 5868
rect 7653 5859 7711 5865
rect 8478 5856 8484 5868
rect 8536 5856 8542 5908
rect 8846 5856 8852 5908
rect 8904 5896 8910 5908
rect 8941 5899 8999 5905
rect 8941 5896 8953 5899
rect 8904 5868 8953 5896
rect 8904 5856 8910 5868
rect 8941 5865 8953 5868
rect 8987 5865 8999 5899
rect 14090 5896 14096 5908
rect 8941 5859 8999 5865
rect 9048 5868 14096 5896
rect 6733 5831 6791 5837
rect 6733 5797 6745 5831
rect 6779 5828 6791 5831
rect 6914 5828 6920 5840
rect 6779 5800 6920 5828
rect 6779 5797 6791 5800
rect 6733 5791 6791 5797
rect 6914 5788 6920 5800
rect 6972 5788 6978 5840
rect 7466 5788 7472 5840
rect 7524 5828 7530 5840
rect 9048 5828 9076 5868
rect 14090 5856 14096 5868
rect 14148 5856 14154 5908
rect 14366 5896 14372 5908
rect 14292 5868 14372 5896
rect 7524 5800 9076 5828
rect 7524 5788 7530 5800
rect 9214 5788 9220 5840
rect 9272 5828 9278 5840
rect 13262 5828 13268 5840
rect 9272 5800 13268 5828
rect 9272 5788 9278 5800
rect 13262 5788 13268 5800
rect 13320 5788 13326 5840
rect 13354 5788 13360 5840
rect 13412 5788 13418 5840
rect 13817 5831 13875 5837
rect 13817 5797 13829 5831
rect 13863 5828 13875 5831
rect 14292 5828 14320 5868
rect 14366 5856 14372 5868
rect 14424 5856 14430 5908
rect 14826 5856 14832 5908
rect 14884 5856 14890 5908
rect 15654 5856 15660 5908
rect 15712 5896 15718 5908
rect 15933 5899 15991 5905
rect 15933 5896 15945 5899
rect 15712 5868 15945 5896
rect 15712 5856 15718 5868
rect 15933 5865 15945 5868
rect 15979 5865 15991 5899
rect 15933 5859 15991 5865
rect 17037 5899 17095 5905
rect 17037 5865 17049 5899
rect 17083 5896 17095 5899
rect 17402 5896 17408 5908
rect 17083 5868 17408 5896
rect 17083 5865 17095 5868
rect 17037 5859 17095 5865
rect 17402 5856 17408 5868
rect 17460 5856 17466 5908
rect 17494 5856 17500 5908
rect 17552 5896 17558 5908
rect 17678 5896 17684 5908
rect 17552 5868 17684 5896
rect 17552 5856 17558 5868
rect 17678 5856 17684 5868
rect 17736 5856 17742 5908
rect 18506 5856 18512 5908
rect 18564 5856 18570 5908
rect 19610 5856 19616 5908
rect 19668 5896 19674 5908
rect 20346 5896 20352 5908
rect 19668 5868 20352 5896
rect 19668 5856 19674 5868
rect 20346 5856 20352 5868
rect 20404 5856 20410 5908
rect 20533 5899 20591 5905
rect 20533 5865 20545 5899
rect 20579 5896 20591 5899
rect 20622 5896 20628 5908
rect 20579 5868 20628 5896
rect 20579 5865 20591 5868
rect 20533 5859 20591 5865
rect 20622 5856 20628 5868
rect 20680 5856 20686 5908
rect 21174 5856 21180 5908
rect 21232 5896 21238 5908
rect 21450 5896 21456 5908
rect 21232 5868 21456 5896
rect 21232 5856 21238 5868
rect 21450 5856 21456 5868
rect 21508 5856 21514 5908
rect 21542 5856 21548 5908
rect 21600 5896 21606 5908
rect 24029 5899 24087 5905
rect 24029 5896 24041 5899
rect 21600 5868 24041 5896
rect 21600 5856 21606 5868
rect 24029 5865 24041 5868
rect 24075 5865 24087 5899
rect 24029 5859 24087 5865
rect 24302 5856 24308 5908
rect 24360 5896 24366 5908
rect 35250 5896 35256 5908
rect 24360 5868 35256 5896
rect 24360 5856 24366 5868
rect 35250 5856 35256 5868
rect 35308 5856 35314 5908
rect 36081 5899 36139 5905
rect 36081 5865 36093 5899
rect 36127 5896 36139 5899
rect 36722 5896 36728 5908
rect 36127 5868 36728 5896
rect 36127 5865 36139 5868
rect 36081 5859 36139 5865
rect 36722 5856 36728 5868
rect 36780 5856 36786 5908
rect 36906 5856 36912 5908
rect 36964 5856 36970 5908
rect 37642 5856 37648 5908
rect 37700 5896 37706 5908
rect 37737 5899 37795 5905
rect 37737 5896 37749 5899
rect 37700 5868 37749 5896
rect 37700 5856 37706 5868
rect 37737 5865 37749 5868
rect 37783 5865 37795 5899
rect 37737 5859 37795 5865
rect 39393 5899 39451 5905
rect 39393 5865 39405 5899
rect 39439 5896 39451 5899
rect 39574 5896 39580 5908
rect 39439 5868 39580 5896
rect 39439 5865 39451 5868
rect 39393 5859 39451 5865
rect 39574 5856 39580 5868
rect 39632 5856 39638 5908
rect 13863 5800 14320 5828
rect 13863 5797 13875 5800
rect 13817 5791 13875 5797
rect 17126 5788 17132 5840
rect 17184 5788 17190 5840
rect 21726 5828 21732 5840
rect 17236 5800 21732 5828
rect 10318 5720 10324 5772
rect 10376 5720 10382 5772
rect 12802 5720 12808 5772
rect 12860 5760 12866 5772
rect 12860 5732 13584 5760
rect 12860 5720 12866 5732
rect 3835 5664 3924 5692
rect 6549 5695 6607 5701
rect 3835 5661 3847 5664
rect 3789 5655 3847 5661
rect 6549 5661 6561 5695
rect 6595 5692 6607 5695
rect 6638 5692 6644 5704
rect 6595 5664 6644 5692
rect 6595 5661 6607 5664
rect 6549 5655 6607 5661
rect 6638 5652 6644 5664
rect 6696 5652 6702 5704
rect 7098 5652 7104 5704
rect 7156 5692 7162 5704
rect 7469 5695 7527 5701
rect 7469 5692 7481 5695
rect 7156 5664 7481 5692
rect 7156 5652 7162 5664
rect 7469 5661 7481 5664
rect 7515 5692 7527 5695
rect 7650 5692 7656 5704
rect 7515 5664 7656 5692
rect 7515 5661 7527 5664
rect 7469 5655 7527 5661
rect 7650 5652 7656 5664
rect 7708 5652 7714 5704
rect 8570 5652 8576 5704
rect 8628 5692 8634 5704
rect 9122 5692 9128 5704
rect 8628 5664 9128 5692
rect 8628 5652 8634 5664
rect 9122 5652 9128 5664
rect 9180 5652 9186 5704
rect 9674 5652 9680 5704
rect 9732 5692 9738 5704
rect 9769 5695 9827 5701
rect 9769 5692 9781 5695
rect 9732 5664 9781 5692
rect 9732 5652 9738 5664
rect 9769 5661 9781 5664
rect 9815 5692 9827 5695
rect 10042 5692 10048 5704
rect 9815 5664 10048 5692
rect 9815 5661 9827 5664
rect 9769 5655 9827 5661
rect 10042 5652 10048 5664
rect 10100 5652 10106 5704
rect 10134 5652 10140 5704
rect 10192 5652 10198 5704
rect 13078 5652 13084 5704
rect 13136 5692 13142 5704
rect 13173 5695 13231 5701
rect 13173 5692 13185 5695
rect 13136 5664 13185 5692
rect 13136 5652 13142 5664
rect 13173 5661 13185 5664
rect 13219 5692 13231 5695
rect 13262 5692 13268 5704
rect 13219 5664 13268 5692
rect 13219 5661 13231 5664
rect 13173 5655 13231 5661
rect 13262 5652 13268 5664
rect 13320 5652 13326 5704
rect 13556 5688 13584 5732
rect 13722 5720 13728 5772
rect 13780 5760 13786 5772
rect 13780 5732 14596 5760
rect 13780 5720 13786 5732
rect 13633 5695 13691 5701
rect 13633 5688 13645 5695
rect 13556 5661 13645 5688
rect 13679 5661 13691 5695
rect 13556 5660 13691 5661
rect 13633 5655 13691 5660
rect 14366 5652 14372 5704
rect 14424 5652 14430 5704
rect 14461 5695 14519 5701
rect 14461 5661 14473 5695
rect 14507 5661 14519 5695
rect 14461 5655 14519 5661
rect 2866 5584 2872 5636
rect 2924 5624 2930 5636
rect 2961 5627 3019 5633
rect 2961 5624 2973 5627
rect 2924 5596 2973 5624
rect 2924 5584 2930 5596
rect 2961 5593 2973 5596
rect 3007 5593 3019 5627
rect 2961 5587 3019 5593
rect 3145 5627 3203 5633
rect 3145 5593 3157 5627
rect 3191 5624 3203 5627
rect 6914 5624 6920 5636
rect 3191 5596 6920 5624
rect 3191 5593 3203 5596
rect 3145 5587 3203 5593
rect 6914 5584 6920 5596
rect 6972 5584 6978 5636
rect 9950 5584 9956 5636
rect 10008 5584 10014 5636
rect 13722 5584 13728 5636
rect 13780 5624 13786 5636
rect 14476 5624 14504 5655
rect 13780 5596 14504 5624
rect 14568 5624 14596 5732
rect 14642 5652 14648 5704
rect 14700 5652 14706 5704
rect 15654 5652 15660 5704
rect 15712 5692 15718 5704
rect 16117 5695 16175 5701
rect 16117 5692 16129 5695
rect 15712 5664 16129 5692
rect 15712 5652 15718 5664
rect 16117 5661 16129 5664
rect 16163 5692 16175 5695
rect 16666 5692 16672 5704
rect 16163 5664 16672 5692
rect 16163 5661 16175 5664
rect 16117 5655 16175 5661
rect 16666 5652 16672 5664
rect 16724 5652 16730 5704
rect 16758 5652 16764 5704
rect 16816 5692 16822 5704
rect 16853 5695 16911 5701
rect 16853 5692 16865 5695
rect 16816 5664 16865 5692
rect 16816 5652 16822 5664
rect 16853 5661 16865 5664
rect 16899 5692 16911 5695
rect 17236 5692 17264 5800
rect 21726 5788 21732 5800
rect 21784 5788 21790 5840
rect 31846 5828 31852 5840
rect 22066 5800 31852 5828
rect 19794 5720 19800 5772
rect 19852 5760 19858 5772
rect 19852 5732 20484 5760
rect 19852 5720 19858 5732
rect 16899 5664 17264 5692
rect 17313 5695 17371 5701
rect 16899 5661 16911 5664
rect 16853 5655 16911 5661
rect 17313 5661 17325 5695
rect 17359 5692 17371 5695
rect 17586 5692 17592 5704
rect 17359 5664 17592 5692
rect 17359 5661 17371 5664
rect 17313 5655 17371 5661
rect 17586 5652 17592 5664
rect 17644 5652 17650 5704
rect 18690 5652 18696 5704
rect 18748 5692 18754 5704
rect 19702 5692 19708 5704
rect 18748 5664 19708 5692
rect 18748 5652 18754 5664
rect 19702 5652 19708 5664
rect 19760 5652 19766 5704
rect 20346 5652 20352 5704
rect 20404 5652 20410 5704
rect 20456 5692 20484 5732
rect 20898 5720 20904 5772
rect 20956 5760 20962 5772
rect 22066 5760 22094 5800
rect 31846 5788 31852 5800
rect 31904 5788 31910 5840
rect 32217 5831 32275 5837
rect 32217 5797 32229 5831
rect 32263 5828 32275 5831
rect 34054 5828 34060 5840
rect 32263 5800 34060 5828
rect 32263 5797 32275 5800
rect 32217 5791 32275 5797
rect 34054 5788 34060 5800
rect 34112 5788 34118 5840
rect 20956 5732 22094 5760
rect 23400 5732 25820 5760
rect 20956 5720 20962 5732
rect 21085 5695 21143 5701
rect 21085 5692 21097 5695
rect 20456 5664 21097 5692
rect 21085 5661 21097 5664
rect 21131 5661 21143 5695
rect 21085 5655 21143 5661
rect 21239 5695 21297 5701
rect 21239 5661 21251 5695
rect 21285 5692 21297 5695
rect 22002 5692 22008 5704
rect 21285 5664 22008 5692
rect 21285 5661 21297 5664
rect 21239 5655 21297 5661
rect 22002 5652 22008 5664
rect 22060 5652 22066 5704
rect 23400 5624 23428 5732
rect 24210 5652 24216 5704
rect 24268 5652 24274 5704
rect 24578 5652 24584 5704
rect 24636 5652 24642 5704
rect 24854 5652 24860 5704
rect 24912 5692 24918 5704
rect 25682 5692 25688 5704
rect 24912 5664 25688 5692
rect 24912 5652 24918 5664
rect 25682 5652 25688 5664
rect 25740 5652 25746 5704
rect 25792 5692 25820 5732
rect 26694 5720 26700 5772
rect 26752 5760 26758 5772
rect 32398 5760 32404 5772
rect 26752 5732 32404 5760
rect 26752 5720 26758 5732
rect 32398 5720 32404 5732
rect 32456 5720 32462 5772
rect 26878 5692 26884 5704
rect 25792 5664 26884 5692
rect 26878 5652 26884 5664
rect 26936 5652 26942 5704
rect 31941 5695 31999 5701
rect 31941 5661 31953 5695
rect 31987 5692 31999 5695
rect 32033 5695 32091 5701
rect 32033 5692 32045 5695
rect 31987 5664 32045 5692
rect 31987 5661 31999 5664
rect 31941 5655 31999 5661
rect 32033 5661 32045 5664
rect 32079 5661 32091 5695
rect 32033 5655 32091 5661
rect 32766 5652 32772 5704
rect 32824 5692 32830 5704
rect 35897 5695 35955 5701
rect 35897 5692 35909 5695
rect 32824 5664 35909 5692
rect 32824 5652 32830 5664
rect 35897 5661 35909 5664
rect 35943 5661 35955 5695
rect 35897 5655 35955 5661
rect 36725 5695 36783 5701
rect 36725 5661 36737 5695
rect 36771 5661 36783 5695
rect 36725 5655 36783 5661
rect 37829 5695 37887 5701
rect 37829 5661 37841 5695
rect 37875 5692 37887 5695
rect 37921 5695 37979 5701
rect 37921 5692 37933 5695
rect 37875 5664 37933 5692
rect 37875 5661 37887 5664
rect 37829 5655 37887 5661
rect 37921 5661 37933 5664
rect 37967 5661 37979 5695
rect 37921 5655 37979 5661
rect 14568 5596 23428 5624
rect 13780 5584 13786 5596
rect 23474 5584 23480 5636
rect 23532 5624 23538 5636
rect 24596 5624 24624 5652
rect 23532 5596 24624 5624
rect 23532 5584 23538 5596
rect 34606 5584 34612 5636
rect 34664 5624 34670 5636
rect 36740 5624 36768 5655
rect 38562 5652 38568 5704
rect 38620 5692 38626 5704
rect 38841 5695 38899 5701
rect 38841 5692 38853 5695
rect 38620 5664 38853 5692
rect 38620 5652 38626 5664
rect 38841 5661 38853 5664
rect 38887 5661 38899 5695
rect 38841 5655 38899 5661
rect 38930 5652 38936 5704
rect 38988 5692 38994 5704
rect 39209 5695 39267 5701
rect 39209 5692 39221 5695
rect 38988 5664 39221 5692
rect 38988 5652 38994 5664
rect 39209 5661 39221 5664
rect 39255 5661 39267 5695
rect 39209 5655 39267 5661
rect 34664 5596 36768 5624
rect 34664 5584 34670 5596
rect 3973 5559 4031 5565
rect 3973 5525 3985 5559
rect 4019 5556 4031 5559
rect 14918 5556 14924 5568
rect 4019 5528 14924 5556
rect 4019 5525 4031 5528
rect 3973 5519 4031 5525
rect 14918 5516 14924 5528
rect 14976 5516 14982 5568
rect 19426 5516 19432 5568
rect 19484 5556 19490 5568
rect 21174 5556 21180 5568
rect 19484 5528 21180 5556
rect 19484 5516 19490 5528
rect 21174 5516 21180 5528
rect 21232 5516 21238 5568
rect 21450 5516 21456 5568
rect 21508 5516 21514 5568
rect 21542 5516 21548 5568
rect 21600 5556 21606 5568
rect 24302 5556 24308 5568
rect 21600 5528 24308 5556
rect 21600 5516 21606 5528
rect 24302 5516 24308 5528
rect 24360 5516 24366 5568
rect 24394 5516 24400 5568
rect 24452 5516 24458 5568
rect 24670 5516 24676 5568
rect 24728 5516 24734 5568
rect 31662 5516 31668 5568
rect 31720 5556 31726 5568
rect 31849 5559 31907 5565
rect 31849 5556 31861 5559
rect 31720 5528 31861 5556
rect 31720 5516 31726 5528
rect 31849 5525 31861 5528
rect 31895 5525 31907 5559
rect 31849 5519 31907 5525
rect 38105 5559 38163 5565
rect 38105 5525 38117 5559
rect 38151 5556 38163 5559
rect 38746 5556 38752 5568
rect 38151 5528 38752 5556
rect 38151 5525 38163 5528
rect 38105 5519 38163 5525
rect 38746 5516 38752 5528
rect 38804 5516 38810 5568
rect 39025 5559 39083 5565
rect 39025 5525 39037 5559
rect 39071 5556 39083 5559
rect 39298 5556 39304 5568
rect 39071 5528 39304 5556
rect 39071 5525 39083 5528
rect 39025 5519 39083 5525
rect 39298 5516 39304 5528
rect 39356 5516 39362 5568
rect 1104 5466 39836 5488
rect 1104 5414 3010 5466
rect 3062 5414 3074 5466
rect 3126 5414 3138 5466
rect 3190 5414 3202 5466
rect 3254 5414 3266 5466
rect 3318 5414 9010 5466
rect 9062 5414 9074 5466
rect 9126 5414 9138 5466
rect 9190 5414 9202 5466
rect 9254 5414 9266 5466
rect 9318 5414 15010 5466
rect 15062 5414 15074 5466
rect 15126 5414 15138 5466
rect 15190 5414 15202 5466
rect 15254 5414 15266 5466
rect 15318 5414 21010 5466
rect 21062 5414 21074 5466
rect 21126 5414 21138 5466
rect 21190 5414 21202 5466
rect 21254 5414 21266 5466
rect 21318 5414 27010 5466
rect 27062 5414 27074 5466
rect 27126 5414 27138 5466
rect 27190 5414 27202 5466
rect 27254 5414 27266 5466
rect 27318 5414 33010 5466
rect 33062 5414 33074 5466
rect 33126 5414 33138 5466
rect 33190 5414 33202 5466
rect 33254 5414 33266 5466
rect 33318 5414 39010 5466
rect 39062 5414 39074 5466
rect 39126 5414 39138 5466
rect 39190 5414 39202 5466
rect 39254 5414 39266 5466
rect 39318 5414 39836 5466
rect 1104 5392 39836 5414
rect 7558 5312 7564 5364
rect 7616 5352 7622 5364
rect 15286 5352 15292 5364
rect 7616 5324 15292 5352
rect 7616 5312 7622 5324
rect 15286 5312 15292 5324
rect 15344 5312 15350 5364
rect 15473 5355 15531 5361
rect 15473 5321 15485 5355
rect 15519 5352 15531 5355
rect 32309 5355 32367 5361
rect 15519 5324 24164 5352
rect 15519 5321 15531 5324
rect 15473 5315 15531 5321
rect 8846 5244 8852 5296
rect 8904 5284 8910 5296
rect 9401 5287 9459 5293
rect 9401 5284 9413 5287
rect 8904 5256 9413 5284
rect 8904 5244 8910 5256
rect 9401 5253 9413 5256
rect 9447 5253 9459 5287
rect 9401 5247 9459 5253
rect 13262 5244 13268 5296
rect 13320 5284 13326 5296
rect 15746 5284 15752 5296
rect 13320 5256 15752 5284
rect 13320 5244 13326 5256
rect 15746 5244 15752 5256
rect 15804 5244 15810 5296
rect 17862 5284 17868 5296
rect 16960 5256 17868 5284
rect 658 5176 664 5228
rect 716 5216 722 5228
rect 2961 5219 3019 5225
rect 2961 5216 2973 5219
rect 716 5188 2973 5216
rect 716 5176 722 5188
rect 2961 5185 2973 5188
rect 3007 5185 3019 5219
rect 2961 5179 3019 5185
rect 3329 5219 3387 5225
rect 3329 5185 3341 5219
rect 3375 5216 3387 5219
rect 3418 5216 3424 5228
rect 3375 5188 3424 5216
rect 3375 5185 3387 5188
rect 3329 5179 3387 5185
rect 3418 5176 3424 5188
rect 3476 5176 3482 5228
rect 14001 5219 14059 5225
rect 14001 5185 14013 5219
rect 14047 5216 14059 5219
rect 14274 5216 14280 5228
rect 14047 5188 14280 5216
rect 14047 5185 14059 5188
rect 14001 5179 14059 5185
rect 14274 5176 14280 5188
rect 14332 5176 14338 5228
rect 15286 5176 15292 5228
rect 15344 5216 15350 5228
rect 16960 5216 16988 5256
rect 17862 5244 17868 5256
rect 17920 5244 17926 5296
rect 19306 5256 20300 5284
rect 15344 5188 16988 5216
rect 15344 5176 15350 5188
rect 17034 5176 17040 5228
rect 17092 5176 17098 5228
rect 17678 5176 17684 5228
rect 17736 5216 17742 5228
rect 19306 5216 19334 5256
rect 17736 5188 19334 5216
rect 17736 5176 17742 5188
rect 19702 5176 19708 5228
rect 19760 5216 19766 5228
rect 19797 5219 19855 5225
rect 19797 5216 19809 5219
rect 19760 5188 19809 5216
rect 19760 5176 19766 5188
rect 19797 5185 19809 5188
rect 19843 5185 19855 5219
rect 20272 5216 20300 5256
rect 20346 5244 20352 5296
rect 20404 5284 20410 5296
rect 24136 5284 24164 5324
rect 26804 5324 31754 5352
rect 26804 5284 26832 5324
rect 20404 5256 22876 5284
rect 24136 5256 26832 5284
rect 31726 5284 31754 5324
rect 32309 5321 32321 5355
rect 32355 5352 32367 5355
rect 32490 5352 32496 5364
rect 32355 5324 32496 5352
rect 32355 5321 32367 5324
rect 32309 5315 32367 5321
rect 32490 5312 32496 5324
rect 32548 5312 32554 5364
rect 37645 5355 37703 5361
rect 37645 5321 37657 5355
rect 37691 5352 37703 5355
rect 37734 5352 37740 5364
rect 37691 5324 37740 5352
rect 37691 5321 37703 5324
rect 37645 5315 37703 5321
rect 37734 5312 37740 5324
rect 37792 5312 37798 5364
rect 38105 5355 38163 5361
rect 38105 5321 38117 5355
rect 38151 5352 38163 5355
rect 38378 5352 38384 5364
rect 38151 5324 38384 5352
rect 38151 5321 38163 5324
rect 38105 5315 38163 5321
rect 38378 5312 38384 5324
rect 38436 5312 38442 5364
rect 38838 5312 38844 5364
rect 38896 5312 38902 5364
rect 39393 5355 39451 5361
rect 39393 5321 39405 5355
rect 39439 5352 39451 5355
rect 39482 5352 39488 5364
rect 39439 5324 39488 5352
rect 39439 5321 39451 5324
rect 39393 5315 39451 5321
rect 39482 5312 39488 5324
rect 39540 5312 39546 5364
rect 38856 5284 38884 5312
rect 31726 5256 38884 5284
rect 20404 5244 20410 5256
rect 22738 5216 22744 5228
rect 20272 5188 22744 5216
rect 19797 5179 19855 5185
rect 22738 5176 22744 5188
rect 22796 5176 22802 5228
rect 9582 5108 9588 5160
rect 9640 5108 9646 5160
rect 13354 5108 13360 5160
rect 13412 5148 13418 5160
rect 13412 5120 17632 5148
rect 13412 5108 13418 5120
rect 3513 5083 3571 5089
rect 3513 5049 3525 5083
rect 3559 5080 3571 5083
rect 4062 5080 4068 5092
rect 3559 5052 4068 5080
rect 3559 5049 3571 5052
rect 3513 5043 3571 5049
rect 4062 5040 4068 5052
rect 4120 5040 4126 5092
rect 12250 5040 12256 5092
rect 12308 5080 12314 5092
rect 15562 5080 15568 5092
rect 12308 5052 15568 5080
rect 12308 5040 12314 5052
rect 15562 5040 15568 5052
rect 15620 5040 15626 5092
rect 16114 5040 16120 5092
rect 16172 5080 16178 5092
rect 17497 5083 17555 5089
rect 17497 5080 17509 5083
rect 16172 5052 17509 5080
rect 16172 5040 16178 5052
rect 17497 5049 17509 5052
rect 17543 5049 17555 5083
rect 17497 5043 17555 5049
rect 3053 5015 3111 5021
rect 3053 4981 3065 5015
rect 3099 5012 3111 5015
rect 3970 5012 3976 5024
rect 3099 4984 3976 5012
rect 3099 4981 3111 4984
rect 3053 4975 3111 4981
rect 3970 4972 3976 4984
rect 4028 4972 4034 5024
rect 14185 5015 14243 5021
rect 14185 4981 14197 5015
rect 14231 5012 14243 5015
rect 15286 5012 15292 5024
rect 14231 4984 15292 5012
rect 14231 4981 14243 4984
rect 14185 4975 14243 4981
rect 15286 4972 15292 4984
rect 15344 4972 15350 5024
rect 16574 4972 16580 5024
rect 16632 5012 16638 5024
rect 16853 5015 16911 5021
rect 16853 5012 16865 5015
rect 16632 4984 16865 5012
rect 16632 4972 16638 4984
rect 16853 4981 16865 4984
rect 16899 4981 16911 5015
rect 17604 5012 17632 5120
rect 19242 5108 19248 5160
rect 19300 5148 19306 5160
rect 19521 5151 19579 5157
rect 19521 5148 19533 5151
rect 19300 5120 19533 5148
rect 19300 5108 19306 5120
rect 19521 5117 19533 5120
rect 19567 5117 19579 5151
rect 22848 5148 22876 5256
rect 25866 5176 25872 5228
rect 25924 5216 25930 5228
rect 26789 5219 26847 5225
rect 26789 5216 26801 5219
rect 25924 5188 26801 5216
rect 25924 5176 25930 5188
rect 26789 5185 26801 5188
rect 26835 5185 26847 5219
rect 26789 5179 26847 5185
rect 26878 5176 26884 5228
rect 26936 5216 26942 5228
rect 31481 5219 31539 5225
rect 31481 5216 31493 5219
rect 26936 5188 31493 5216
rect 26936 5176 26942 5188
rect 31481 5185 31493 5188
rect 31527 5185 31539 5219
rect 31481 5179 31539 5185
rect 31570 5176 31576 5228
rect 31628 5216 31634 5228
rect 32125 5219 32183 5225
rect 32125 5216 32137 5219
rect 31628 5188 32137 5216
rect 31628 5176 31634 5188
rect 32125 5185 32137 5188
rect 32171 5185 32183 5219
rect 32125 5179 32183 5185
rect 36078 5176 36084 5228
rect 36136 5216 36142 5228
rect 37461 5219 37519 5225
rect 37461 5216 37473 5219
rect 36136 5188 37473 5216
rect 36136 5176 36142 5188
rect 37461 5185 37473 5188
rect 37507 5185 37519 5219
rect 37461 5179 37519 5185
rect 37642 5176 37648 5228
rect 37700 5216 37706 5228
rect 37921 5219 37979 5225
rect 37921 5216 37933 5219
rect 37700 5188 37933 5216
rect 37700 5176 37706 5188
rect 37921 5185 37933 5188
rect 37967 5185 37979 5219
rect 37921 5179 37979 5185
rect 38838 5176 38844 5228
rect 38896 5176 38902 5228
rect 39206 5176 39212 5228
rect 39264 5176 39270 5228
rect 36262 5148 36268 5160
rect 22848 5120 36268 5148
rect 19521 5111 19579 5117
rect 36262 5108 36268 5120
rect 36320 5108 36326 5160
rect 26602 5040 26608 5092
rect 26660 5040 26666 5092
rect 31665 5083 31723 5089
rect 31665 5049 31677 5083
rect 31711 5080 31723 5083
rect 35986 5080 35992 5092
rect 31711 5052 35992 5080
rect 31711 5049 31723 5052
rect 31665 5043 31723 5049
rect 35986 5040 35992 5052
rect 36044 5040 36050 5092
rect 20346 5012 20352 5024
rect 17604 4984 20352 5012
rect 16853 4975 16911 4981
rect 20346 4972 20352 4984
rect 20404 4972 20410 5024
rect 20533 5015 20591 5021
rect 20533 4981 20545 5015
rect 20579 5012 20591 5015
rect 21910 5012 21916 5024
rect 20579 4984 21916 5012
rect 20579 4981 20591 4984
rect 20533 4975 20591 4981
rect 21910 4972 21916 4984
rect 21968 5012 21974 5024
rect 22646 5012 22652 5024
rect 21968 4984 22652 5012
rect 21968 4972 21974 4984
rect 22646 4972 22652 4984
rect 22704 4972 22710 5024
rect 39022 4972 39028 5024
rect 39080 4972 39086 5024
rect 1104 4922 39836 4944
rect 1104 4870 1950 4922
rect 2002 4870 2014 4922
rect 2066 4870 2078 4922
rect 2130 4870 2142 4922
rect 2194 4870 2206 4922
rect 2258 4870 7950 4922
rect 8002 4870 8014 4922
rect 8066 4870 8078 4922
rect 8130 4870 8142 4922
rect 8194 4870 8206 4922
rect 8258 4870 13950 4922
rect 14002 4870 14014 4922
rect 14066 4870 14078 4922
rect 14130 4870 14142 4922
rect 14194 4870 14206 4922
rect 14258 4870 19950 4922
rect 20002 4870 20014 4922
rect 20066 4870 20078 4922
rect 20130 4870 20142 4922
rect 20194 4870 20206 4922
rect 20258 4870 25950 4922
rect 26002 4870 26014 4922
rect 26066 4870 26078 4922
rect 26130 4870 26142 4922
rect 26194 4870 26206 4922
rect 26258 4870 31950 4922
rect 32002 4870 32014 4922
rect 32066 4870 32078 4922
rect 32130 4870 32142 4922
rect 32194 4870 32206 4922
rect 32258 4870 37950 4922
rect 38002 4870 38014 4922
rect 38066 4870 38078 4922
rect 38130 4870 38142 4922
rect 38194 4870 38206 4922
rect 38258 4870 39836 4922
rect 1104 4848 39836 4870
rect 9858 4768 9864 4820
rect 9916 4808 9922 4820
rect 10781 4811 10839 4817
rect 10781 4808 10793 4811
rect 9916 4780 10793 4808
rect 9916 4768 9922 4780
rect 10781 4777 10793 4780
rect 10827 4777 10839 4811
rect 10781 4771 10839 4777
rect 12250 4768 12256 4820
rect 12308 4768 12314 4820
rect 13354 4768 13360 4820
rect 13412 4768 13418 4820
rect 13538 4768 13544 4820
rect 13596 4768 13602 4820
rect 14274 4768 14280 4820
rect 14332 4768 14338 4820
rect 16022 4768 16028 4820
rect 16080 4808 16086 4820
rect 16209 4811 16267 4817
rect 16209 4808 16221 4811
rect 16080 4780 16221 4808
rect 16080 4768 16086 4780
rect 16209 4777 16221 4780
rect 16255 4777 16267 4811
rect 16209 4771 16267 4777
rect 17034 4768 17040 4820
rect 17092 4808 17098 4820
rect 21634 4808 21640 4820
rect 17092 4780 21640 4808
rect 17092 4768 17098 4780
rect 21634 4768 21640 4780
rect 21692 4768 21698 4820
rect 21726 4768 21732 4820
rect 21784 4768 21790 4820
rect 32033 4811 32091 4817
rect 32033 4777 32045 4811
rect 32079 4808 32091 4811
rect 32858 4808 32864 4820
rect 32079 4780 32864 4808
rect 32079 4777 32091 4780
rect 32033 4771 32091 4777
rect 32858 4768 32864 4780
rect 32916 4768 32922 4820
rect 37826 4768 37832 4820
rect 37884 4808 37890 4820
rect 37921 4811 37979 4817
rect 37921 4808 37933 4811
rect 37884 4780 37933 4808
rect 37884 4768 37890 4780
rect 37921 4777 37933 4780
rect 37967 4777 37979 4811
rect 37921 4771 37979 4777
rect 39390 4768 39396 4820
rect 39448 4768 39454 4820
rect 3510 4700 3516 4752
rect 3568 4740 3574 4752
rect 38838 4740 38844 4752
rect 3568 4712 38844 4740
rect 3568 4700 3574 4712
rect 38838 4700 38844 4712
rect 38896 4700 38902 4752
rect 3145 4675 3203 4681
rect 3145 4641 3157 4675
rect 3191 4672 3203 4675
rect 3878 4672 3884 4684
rect 3191 4644 3884 4672
rect 3191 4641 3203 4644
rect 3145 4635 3203 4641
rect 3878 4632 3884 4644
rect 3936 4632 3942 4684
rect 12710 4672 12716 4684
rect 7484 4644 11100 4672
rect 3421 4607 3479 4613
rect 3421 4573 3433 4607
rect 3467 4604 3479 4607
rect 7282 4604 7288 4616
rect 3467 4576 7288 4604
rect 3467 4573 3479 4576
rect 3421 4567 3479 4573
rect 7282 4564 7288 4576
rect 7340 4564 7346 4616
rect 2774 4496 2780 4548
rect 2832 4536 2838 4548
rect 2961 4539 3019 4545
rect 2961 4536 2973 4539
rect 2832 4508 2973 4536
rect 2832 4496 2838 4508
rect 2961 4505 2973 4508
rect 3007 4505 3019 4539
rect 7484 4536 7512 4644
rect 7558 4564 7564 4616
rect 7616 4604 7622 4616
rect 8754 4604 8760 4616
rect 7616 4576 8760 4604
rect 7616 4564 7622 4576
rect 8754 4564 8760 4576
rect 8812 4604 8818 4616
rect 10965 4607 11023 4613
rect 10965 4604 10977 4607
rect 8812 4576 10977 4604
rect 8812 4564 8818 4576
rect 10965 4573 10977 4576
rect 11011 4573 11023 4607
rect 10965 4567 11023 4573
rect 2961 4499 3019 4505
rect 3620 4508 7512 4536
rect 3620 4477 3648 4508
rect 3605 4471 3663 4477
rect 3605 4437 3617 4471
rect 3651 4437 3663 4471
rect 10980 4468 11008 4567
rect 11072 4536 11100 4644
rect 11256 4644 12716 4672
rect 11256 4613 11284 4644
rect 12710 4632 12716 4644
rect 12768 4632 12774 4684
rect 13814 4672 13820 4684
rect 13280 4644 13820 4672
rect 11241 4607 11299 4613
rect 11241 4573 11253 4607
rect 11287 4573 11299 4607
rect 11241 4567 11299 4573
rect 11422 4564 11428 4616
rect 11480 4564 11486 4616
rect 11606 4564 11612 4616
rect 11664 4604 11670 4616
rect 12066 4604 12072 4616
rect 11664 4576 12072 4604
rect 11664 4564 11670 4576
rect 12066 4564 12072 4576
rect 12124 4564 12130 4616
rect 12158 4564 12164 4616
rect 12216 4604 12222 4616
rect 13280 4604 13308 4644
rect 13814 4632 13820 4644
rect 13872 4632 13878 4684
rect 15286 4632 15292 4684
rect 15344 4672 15350 4684
rect 38286 4672 38292 4684
rect 15344 4644 38292 4672
rect 15344 4632 15350 4644
rect 38286 4632 38292 4644
rect 38344 4632 38350 4684
rect 38654 4632 38660 4684
rect 38712 4672 38718 4684
rect 38712 4644 39252 4672
rect 38712 4632 38718 4644
rect 12216 4576 13308 4604
rect 12216 4564 12222 4576
rect 13722 4564 13728 4616
rect 13780 4564 13786 4616
rect 14093 4607 14151 4613
rect 14093 4573 14105 4607
rect 14139 4604 14151 4607
rect 14458 4604 14464 4616
rect 14139 4576 14464 4604
rect 14139 4573 14151 4576
rect 14093 4567 14151 4573
rect 14458 4564 14464 4576
rect 14516 4564 14522 4616
rect 14550 4564 14556 4616
rect 14608 4604 14614 4616
rect 16390 4604 16396 4616
rect 14608 4576 16396 4604
rect 14608 4564 14614 4576
rect 16390 4564 16396 4576
rect 16448 4564 16454 4616
rect 16666 4564 16672 4616
rect 16724 4564 16730 4616
rect 16853 4607 16911 4613
rect 16853 4573 16865 4607
rect 16899 4604 16911 4607
rect 17586 4604 17592 4616
rect 16899 4576 17592 4604
rect 16899 4573 16911 4576
rect 16853 4567 16911 4573
rect 17586 4564 17592 4576
rect 17644 4564 17650 4616
rect 20714 4564 20720 4616
rect 20772 4604 20778 4616
rect 21913 4607 21971 4613
rect 21913 4604 21925 4607
rect 20772 4576 21925 4604
rect 20772 4564 20778 4576
rect 21913 4573 21925 4576
rect 21959 4573 21971 4607
rect 21913 4567 21971 4573
rect 31481 4607 31539 4613
rect 31481 4573 31493 4607
rect 31527 4604 31539 4607
rect 31573 4607 31631 4613
rect 31573 4604 31585 4607
rect 31527 4576 31585 4604
rect 31527 4573 31539 4576
rect 31481 4567 31539 4573
rect 31573 4573 31585 4576
rect 31619 4573 31631 4607
rect 31849 4607 31907 4613
rect 31849 4604 31861 4607
rect 31573 4567 31631 4573
rect 31726 4576 31861 4604
rect 13170 4536 13176 4548
rect 11072 4508 12296 4536
rect 12158 4468 12164 4480
rect 10980 4440 12164 4468
rect 3605 4431 3663 4437
rect 12158 4428 12164 4440
rect 12216 4428 12222 4480
rect 12268 4468 12296 4508
rect 12406 4508 13176 4536
rect 12406 4468 12434 4508
rect 13170 4496 13176 4508
rect 13228 4496 13234 4548
rect 13265 4539 13323 4545
rect 13265 4505 13277 4539
rect 13311 4505 13323 4539
rect 13265 4499 13323 4505
rect 12268 4440 12434 4468
rect 12526 4428 12532 4480
rect 12584 4468 12590 4480
rect 13280 4468 13308 4499
rect 14274 4496 14280 4548
rect 14332 4536 14338 4548
rect 30374 4536 30380 4548
rect 14332 4508 30380 4536
rect 14332 4496 14338 4508
rect 30374 4496 30380 4508
rect 30432 4496 30438 4548
rect 31205 4539 31263 4545
rect 31205 4505 31217 4539
rect 31251 4536 31263 4539
rect 31726 4536 31754 4576
rect 31849 4573 31861 4576
rect 31895 4573 31907 4607
rect 31849 4567 31907 4573
rect 38105 4607 38163 4613
rect 38105 4573 38117 4607
rect 38151 4573 38163 4607
rect 38105 4567 38163 4573
rect 38841 4607 38899 4613
rect 38841 4573 38853 4607
rect 38887 4604 38899 4607
rect 38930 4604 38936 4616
rect 38887 4576 38936 4604
rect 38887 4573 38899 4576
rect 38841 4567 38899 4573
rect 31251 4508 31754 4536
rect 38120 4536 38148 4567
rect 38930 4564 38936 4576
rect 38988 4564 38994 4616
rect 39224 4613 39252 4644
rect 39209 4607 39267 4613
rect 39209 4573 39221 4607
rect 39255 4573 39267 4607
rect 39209 4567 39267 4573
rect 39574 4536 39580 4548
rect 38120 4508 39580 4536
rect 31251 4505 31263 4508
rect 31205 4499 31263 4505
rect 39574 4496 39580 4508
rect 39632 4496 39638 4548
rect 18322 4468 18328 4480
rect 12584 4440 18328 4468
rect 12584 4428 12590 4440
rect 18322 4428 18328 4440
rect 18380 4428 18386 4480
rect 19702 4428 19708 4480
rect 19760 4468 19766 4480
rect 22462 4468 22468 4480
rect 19760 4440 22468 4468
rect 19760 4428 19766 4440
rect 22462 4428 22468 4440
rect 22520 4428 22526 4480
rect 25038 4428 25044 4480
rect 25096 4468 25102 4480
rect 31113 4471 31171 4477
rect 31113 4468 31125 4471
rect 25096 4440 31125 4468
rect 25096 4428 25102 4440
rect 31113 4437 31125 4440
rect 31159 4437 31171 4471
rect 31113 4431 31171 4437
rect 31294 4428 31300 4480
rect 31352 4468 31358 4480
rect 31389 4471 31447 4477
rect 31389 4468 31401 4471
rect 31352 4440 31401 4468
rect 31352 4428 31358 4440
rect 31389 4437 31401 4440
rect 31435 4437 31447 4471
rect 31389 4431 31447 4437
rect 31757 4471 31815 4477
rect 31757 4437 31769 4471
rect 31803 4468 31815 4471
rect 33502 4468 33508 4480
rect 31803 4440 33508 4468
rect 31803 4437 31815 4440
rect 31757 4431 31815 4437
rect 33502 4428 33508 4440
rect 33560 4428 33566 4480
rect 39025 4471 39083 4477
rect 39025 4437 39037 4471
rect 39071 4468 39083 4471
rect 39298 4468 39304 4480
rect 39071 4440 39304 4468
rect 39071 4437 39083 4440
rect 39025 4431 39083 4437
rect 39298 4428 39304 4440
rect 39356 4428 39362 4480
rect 1104 4378 39836 4400
rect 1104 4326 3010 4378
rect 3062 4326 3074 4378
rect 3126 4326 3138 4378
rect 3190 4326 3202 4378
rect 3254 4326 3266 4378
rect 3318 4326 9010 4378
rect 9062 4326 9074 4378
rect 9126 4326 9138 4378
rect 9190 4326 9202 4378
rect 9254 4326 9266 4378
rect 9318 4326 15010 4378
rect 15062 4326 15074 4378
rect 15126 4326 15138 4378
rect 15190 4326 15202 4378
rect 15254 4326 15266 4378
rect 15318 4326 21010 4378
rect 21062 4326 21074 4378
rect 21126 4326 21138 4378
rect 21190 4326 21202 4378
rect 21254 4326 21266 4378
rect 21318 4326 27010 4378
rect 27062 4326 27074 4378
rect 27126 4326 27138 4378
rect 27190 4326 27202 4378
rect 27254 4326 27266 4378
rect 27318 4326 33010 4378
rect 33062 4326 33074 4378
rect 33126 4326 33138 4378
rect 33190 4326 33202 4378
rect 33254 4326 33266 4378
rect 33318 4326 39010 4378
rect 39062 4326 39074 4378
rect 39126 4326 39138 4378
rect 39190 4326 39202 4378
rect 39254 4326 39266 4378
rect 39318 4326 39836 4378
rect 1104 4304 39836 4326
rect 1210 4224 1216 4276
rect 1268 4264 1274 4276
rect 1268 4236 2774 4264
rect 1268 4224 1274 4236
rect 1302 4156 1308 4208
rect 1360 4196 1366 4208
rect 2501 4199 2559 4205
rect 2501 4196 2513 4199
rect 1360 4168 2513 4196
rect 1360 4156 1366 4168
rect 2501 4165 2513 4168
rect 2547 4165 2559 4199
rect 2746 4196 2774 4236
rect 7282 4224 7288 4276
rect 7340 4264 7346 4276
rect 7340 4236 8064 4264
rect 7340 4224 7346 4236
rect 3237 4199 3295 4205
rect 3237 4196 3249 4199
rect 2746 4168 3249 4196
rect 2501 4159 2559 4165
rect 3237 4165 3249 4168
rect 3283 4165 3295 4199
rect 3237 4159 3295 4165
rect 3602 4156 3608 4208
rect 3660 4156 3666 4208
rect 8036 4196 8064 4236
rect 8662 4224 8668 4276
rect 8720 4264 8726 4276
rect 18046 4264 18052 4276
rect 8720 4236 18052 4264
rect 8720 4224 8726 4236
rect 18046 4224 18052 4236
rect 18104 4224 18110 4276
rect 19518 4224 19524 4276
rect 19576 4264 19582 4276
rect 21818 4264 21824 4276
rect 19576 4236 21824 4264
rect 19576 4224 19582 4236
rect 21818 4224 21824 4236
rect 21876 4224 21882 4276
rect 23842 4224 23848 4276
rect 23900 4224 23906 4276
rect 23750 4196 23756 4208
rect 8036 4168 23756 4196
rect 23750 4156 23756 4168
rect 23808 4156 23814 4208
rect 28258 4156 28264 4208
rect 28316 4196 28322 4208
rect 32582 4196 32588 4208
rect 28316 4168 32588 4196
rect 28316 4156 28322 4168
rect 32582 4156 32588 4168
rect 32640 4156 32646 4208
rect 2866 4088 2872 4140
rect 2924 4088 2930 4140
rect 6365 4131 6423 4137
rect 6365 4097 6377 4131
rect 6411 4128 6423 4131
rect 6411 4100 6776 4128
rect 6411 4097 6423 4100
rect 6365 4091 6423 4097
rect 2685 4063 2743 4069
rect 2685 4029 2697 4063
rect 2731 4060 2743 4063
rect 4706 4060 4712 4072
rect 2731 4032 4712 4060
rect 2731 4029 2743 4032
rect 2685 4023 2743 4029
rect 4706 4020 4712 4032
rect 4764 4020 4770 4072
rect 6549 4063 6607 4069
rect 6549 4029 6561 4063
rect 6595 4060 6607 4063
rect 6638 4060 6644 4072
rect 6595 4032 6644 4060
rect 6595 4029 6607 4032
rect 6549 4023 6607 4029
rect 6638 4020 6644 4032
rect 6696 4020 6702 4072
rect 6748 4060 6776 4100
rect 7282 4088 7288 4140
rect 7340 4088 7346 4140
rect 7374 4088 7380 4140
rect 7432 4137 7438 4140
rect 7432 4131 7460 4137
rect 7448 4097 7460 4131
rect 7432 4091 7460 4097
rect 7432 4088 7438 4091
rect 7558 4088 7564 4140
rect 7616 4088 7622 4140
rect 8570 4088 8576 4140
rect 8628 4088 8634 4140
rect 9582 4088 9588 4140
rect 9640 4128 9646 4140
rect 9861 4131 9919 4137
rect 9861 4128 9873 4131
rect 9640 4100 9873 4128
rect 9640 4088 9646 4100
rect 9861 4097 9873 4100
rect 9907 4097 9919 4131
rect 9861 4091 9919 4097
rect 10136 4131 10194 4137
rect 10136 4097 10148 4131
rect 10182 4097 10194 4131
rect 10136 4091 10194 4097
rect 7098 4060 7104 4072
rect 6748 4032 7104 4060
rect 7098 4020 7104 4032
rect 7156 4020 7162 4072
rect 7742 4020 7748 4072
rect 7800 4060 7806 4072
rect 8205 4063 8263 4069
rect 8205 4060 8217 4063
rect 7800 4032 8217 4060
rect 7800 4020 7806 4032
rect 8205 4029 8217 4032
rect 8251 4029 8263 4063
rect 8205 4023 8263 4029
rect 8481 4063 8539 4069
rect 8481 4029 8493 4063
rect 8527 4029 8539 4063
rect 10152 4060 10180 4091
rect 10226 4088 10232 4140
rect 10284 4088 10290 4140
rect 11330 4088 11336 4140
rect 11388 4128 11394 4140
rect 14550 4128 14556 4140
rect 11388 4100 14556 4128
rect 11388 4088 11394 4100
rect 14550 4088 14556 4100
rect 14608 4088 14614 4140
rect 15197 4131 15255 4137
rect 15197 4097 15209 4131
rect 15243 4128 15255 4131
rect 15562 4128 15568 4140
rect 15243 4100 15568 4128
rect 15243 4097 15255 4100
rect 15197 4091 15255 4097
rect 15562 4088 15568 4100
rect 15620 4088 15626 4140
rect 18046 4137 18052 4140
rect 17854 4132 17912 4137
rect 17788 4131 17912 4132
rect 17788 4104 17866 4131
rect 12710 4060 12716 4072
rect 8481 4023 8539 4029
rect 8680 4032 12716 4060
rect 3050 3952 3056 4004
rect 3108 3952 3114 4004
rect 3786 3952 3792 4004
rect 3844 3952 3850 4004
rect 7009 3995 7067 4001
rect 7009 3961 7021 3995
rect 7055 3961 7067 3995
rect 8496 3992 8524 4023
rect 8680 3992 8708 4032
rect 12710 4020 12716 4032
rect 12768 4020 12774 4072
rect 15289 4063 15347 4069
rect 15289 4029 15301 4063
rect 15335 4029 15347 4063
rect 15289 4023 15347 4029
rect 7009 3955 7067 3961
rect 7944 3964 8708 3992
rect 9033 3995 9091 4001
rect 3329 3927 3387 3933
rect 3329 3893 3341 3927
rect 3375 3924 3387 3927
rect 3510 3924 3516 3936
rect 3375 3896 3516 3924
rect 3375 3893 3387 3896
rect 3329 3887 3387 3893
rect 3510 3884 3516 3896
rect 3568 3884 3574 3936
rect 7024 3924 7052 3955
rect 7944 3924 7972 3964
rect 9033 3961 9045 3995
rect 9079 3992 9091 3995
rect 9398 3992 9404 4004
rect 9079 3964 9404 3992
rect 9079 3961 9091 3964
rect 9033 3955 9091 3961
rect 9398 3952 9404 3964
rect 9456 3952 9462 4004
rect 14734 3952 14740 4004
rect 14792 3992 14798 4004
rect 14829 3995 14887 4001
rect 14829 3992 14841 3995
rect 14792 3964 14841 3992
rect 14792 3952 14798 3964
rect 14829 3961 14841 3964
rect 14875 3961 14887 3995
rect 15304 3992 15332 4023
rect 15470 4020 15476 4072
rect 15528 4060 15534 4072
rect 16666 4060 16672 4072
rect 15528 4032 16672 4060
rect 15528 4020 15534 4032
rect 16666 4020 16672 4032
rect 16724 4020 16730 4072
rect 17788 4060 17816 4104
rect 17854 4097 17866 4104
rect 17900 4097 17912 4131
rect 17854 4091 17912 4097
rect 18013 4131 18052 4137
rect 18013 4097 18025 4131
rect 18013 4091 18052 4097
rect 18046 4088 18052 4091
rect 18104 4088 18110 4140
rect 18138 4088 18144 4140
rect 18196 4088 18202 4140
rect 18233 4131 18291 4137
rect 18233 4097 18245 4131
rect 18279 4097 18291 4131
rect 18233 4091 18291 4097
rect 18371 4131 18429 4137
rect 18371 4097 18383 4131
rect 18417 4128 18429 4131
rect 18874 4128 18880 4140
rect 18417 4100 18880 4128
rect 18417 4097 18429 4100
rect 18371 4091 18429 4097
rect 18248 4060 18276 4091
rect 18874 4088 18880 4100
rect 18932 4088 18938 4140
rect 20254 4088 20260 4140
rect 20312 4088 20318 4140
rect 21450 4128 21456 4140
rect 20364 4100 21456 4128
rect 20364 4060 20392 4100
rect 21450 4088 21456 4100
rect 21508 4088 21514 4140
rect 22646 4088 22652 4140
rect 22704 4128 22710 4140
rect 24029 4131 24087 4137
rect 24298 4132 24356 4137
rect 24029 4128 24041 4131
rect 22704 4100 24041 4128
rect 22704 4088 22710 4100
rect 24029 4097 24041 4100
rect 24075 4097 24087 4131
rect 24228 4131 24356 4132
rect 24228 4128 24310 4131
rect 24029 4091 24087 4097
rect 24136 4104 24310 4128
rect 24136 4100 24256 4104
rect 17788 4032 18000 4060
rect 18248 4032 20392 4060
rect 17862 3992 17868 4004
rect 15304 3964 17868 3992
rect 14829 3955 14887 3961
rect 17862 3952 17868 3964
rect 17920 3952 17926 4004
rect 7024 3896 7972 3924
rect 17972 3924 18000 4032
rect 22278 4020 22284 4072
rect 22336 4060 22342 4072
rect 22830 4060 22836 4072
rect 22336 4032 22836 4060
rect 22336 4020 22342 4032
rect 22830 4020 22836 4032
rect 22888 4020 22894 4072
rect 23290 4020 23296 4072
rect 23348 4060 23354 4072
rect 24136 4060 24164 4100
rect 24298 4097 24310 4104
rect 24344 4097 24356 4131
rect 24298 4091 24356 4097
rect 24489 4131 24547 4137
rect 24489 4097 24501 4131
rect 24535 4128 24547 4131
rect 24762 4128 24768 4140
rect 24535 4100 24768 4128
rect 24535 4097 24547 4100
rect 24489 4091 24547 4097
rect 24762 4088 24768 4100
rect 24820 4088 24826 4140
rect 30653 4131 30711 4137
rect 30653 4097 30665 4131
rect 30699 4128 30711 4131
rect 30745 4131 30803 4137
rect 30745 4128 30757 4131
rect 30699 4100 30757 4128
rect 30699 4097 30711 4100
rect 30653 4091 30711 4097
rect 30745 4097 30757 4100
rect 30791 4097 30803 4131
rect 30745 4091 30803 4097
rect 38838 4088 38844 4140
rect 38896 4088 38902 4140
rect 39209 4131 39267 4137
rect 39209 4097 39221 4131
rect 39255 4097 39267 4131
rect 39209 4091 39267 4097
rect 23348 4032 24164 4060
rect 23348 4020 23354 4032
rect 38746 4020 38752 4072
rect 38804 4060 38810 4072
rect 39224 4060 39252 4091
rect 38804 4032 39252 4060
rect 38804 4020 38810 4032
rect 18509 3995 18567 4001
rect 18509 3961 18521 3995
rect 18555 3992 18567 3995
rect 20346 3992 20352 4004
rect 18555 3964 20352 3992
rect 18555 3961 18567 3964
rect 18509 3955 18567 3961
rect 20346 3952 20352 3964
rect 20404 3952 20410 4004
rect 20441 3995 20499 4001
rect 20441 3961 20453 3995
rect 20487 3992 20499 3995
rect 30742 3992 30748 4004
rect 20487 3964 30748 3992
rect 20487 3961 20499 3964
rect 20441 3955 20499 3961
rect 30742 3952 30748 3964
rect 30800 3952 30806 4004
rect 30926 3952 30932 4004
rect 30984 3952 30990 4004
rect 39393 3995 39451 4001
rect 39393 3961 39405 3995
rect 39439 3992 39451 3995
rect 39482 3992 39488 4004
rect 39439 3964 39488 3992
rect 39439 3961 39451 3964
rect 39393 3955 39451 3961
rect 39482 3952 39488 3964
rect 39540 3952 39546 4004
rect 19610 3924 19616 3936
rect 17972 3896 19616 3924
rect 19610 3884 19616 3896
rect 19668 3884 19674 3936
rect 22554 3884 22560 3936
rect 22612 3924 22618 3936
rect 23290 3924 23296 3936
rect 22612 3896 23296 3924
rect 22612 3884 22618 3896
rect 23290 3884 23296 3896
rect 23348 3884 23354 3936
rect 23382 3884 23388 3936
rect 23440 3924 23446 3936
rect 24854 3924 24860 3936
rect 23440 3896 24860 3924
rect 23440 3884 23446 3896
rect 24854 3884 24860 3896
rect 24912 3884 24918 3936
rect 30282 3884 30288 3936
rect 30340 3924 30346 3936
rect 30561 3927 30619 3933
rect 30561 3924 30573 3927
rect 30340 3896 30573 3924
rect 30340 3884 30346 3896
rect 30561 3893 30573 3896
rect 30607 3893 30619 3927
rect 30561 3887 30619 3893
rect 39022 3884 39028 3936
rect 39080 3884 39086 3936
rect 1104 3834 39836 3856
rect 1104 3782 1950 3834
rect 2002 3782 2014 3834
rect 2066 3782 2078 3834
rect 2130 3782 2142 3834
rect 2194 3782 2206 3834
rect 2258 3782 7950 3834
rect 8002 3782 8014 3834
rect 8066 3782 8078 3834
rect 8130 3782 8142 3834
rect 8194 3782 8206 3834
rect 8258 3782 13950 3834
rect 14002 3782 14014 3834
rect 14066 3782 14078 3834
rect 14130 3782 14142 3834
rect 14194 3782 14206 3834
rect 14258 3782 19950 3834
rect 20002 3782 20014 3834
rect 20066 3782 20078 3834
rect 20130 3782 20142 3834
rect 20194 3782 20206 3834
rect 20258 3782 25950 3834
rect 26002 3782 26014 3834
rect 26066 3782 26078 3834
rect 26130 3782 26142 3834
rect 26194 3782 26206 3834
rect 26258 3782 31950 3834
rect 32002 3782 32014 3834
rect 32066 3782 32078 3834
rect 32130 3782 32142 3834
rect 32194 3782 32206 3834
rect 32258 3782 37950 3834
rect 38002 3782 38014 3834
rect 38066 3782 38078 3834
rect 38130 3782 38142 3834
rect 38194 3782 38206 3834
rect 38258 3782 39836 3834
rect 1104 3760 39836 3782
rect 9217 3723 9275 3729
rect 9217 3689 9229 3723
rect 9263 3720 9275 3723
rect 9490 3720 9496 3732
rect 9263 3692 9496 3720
rect 9263 3689 9275 3692
rect 9217 3683 9275 3689
rect 9490 3680 9496 3692
rect 9548 3680 9554 3732
rect 10689 3723 10747 3729
rect 10689 3689 10701 3723
rect 10735 3720 10747 3723
rect 13630 3720 13636 3732
rect 10735 3692 13636 3720
rect 10735 3689 10747 3692
rect 10689 3683 10747 3689
rect 13630 3680 13636 3692
rect 13688 3680 13694 3732
rect 14185 3723 14243 3729
rect 14185 3689 14197 3723
rect 14231 3720 14243 3723
rect 14366 3720 14372 3732
rect 14231 3692 14372 3720
rect 14231 3689 14243 3692
rect 14185 3683 14243 3689
rect 14366 3680 14372 3692
rect 14424 3680 14430 3732
rect 15378 3680 15384 3732
rect 15436 3680 15442 3732
rect 15933 3723 15991 3729
rect 15933 3689 15945 3723
rect 15979 3720 15991 3723
rect 15979 3692 18092 3720
rect 15979 3689 15991 3692
rect 15933 3683 15991 3689
rect 13722 3652 13728 3664
rect 12360 3624 13728 3652
rect 11330 3544 11336 3596
rect 11388 3544 11394 3596
rect 11514 3593 11520 3596
rect 11492 3587 11520 3593
rect 11492 3553 11504 3587
rect 11492 3547 11520 3553
rect 11514 3544 11520 3547
rect 11572 3544 11578 3596
rect 11606 3544 11612 3596
rect 11664 3544 11670 3596
rect 12360 3593 12388 3624
rect 13722 3612 13728 3624
rect 13780 3612 13786 3664
rect 17678 3652 17684 3664
rect 17052 3624 17684 3652
rect 11885 3587 11943 3593
rect 11885 3553 11897 3587
rect 11931 3584 11943 3587
rect 12345 3587 12403 3593
rect 11931 3556 12296 3584
rect 11931 3553 11943 3556
rect 11885 3547 11943 3553
rect 8478 3476 8484 3528
rect 8536 3516 8542 3528
rect 9125 3519 9183 3525
rect 9125 3516 9137 3519
rect 8536 3488 9137 3516
rect 8536 3476 8542 3488
rect 9125 3485 9137 3488
rect 9171 3485 9183 3519
rect 12268 3516 12296 3556
rect 12345 3553 12357 3587
rect 12391 3553 12403 3587
rect 12345 3547 12403 3553
rect 12529 3587 12587 3593
rect 12529 3553 12541 3587
rect 12575 3584 12587 3587
rect 12986 3584 12992 3596
rect 12575 3556 12992 3584
rect 12575 3553 12587 3556
rect 12529 3547 12587 3553
rect 12986 3544 12992 3556
rect 13044 3544 13050 3596
rect 16574 3544 16580 3596
rect 16632 3544 16638 3596
rect 16758 3593 16764 3596
rect 16736 3587 16764 3593
rect 16736 3553 16748 3587
rect 16736 3547 16764 3553
rect 16758 3544 16764 3547
rect 16816 3544 16822 3596
rect 16853 3587 16911 3593
rect 16853 3553 16865 3587
rect 16899 3584 16911 3587
rect 17052 3584 17080 3624
rect 17678 3612 17684 3624
rect 17736 3612 17742 3664
rect 18064 3652 18092 3692
rect 18138 3680 18144 3732
rect 18196 3720 18202 3732
rect 20717 3723 20775 3729
rect 20717 3720 20729 3723
rect 18196 3692 20729 3720
rect 18196 3680 18202 3692
rect 20717 3689 20729 3692
rect 20763 3689 20775 3723
rect 22002 3720 22008 3732
rect 20717 3683 20775 3689
rect 21652 3692 22008 3720
rect 19518 3652 19524 3664
rect 18064 3624 19524 3652
rect 19518 3612 19524 3624
rect 19576 3612 19582 3664
rect 19705 3655 19763 3661
rect 19705 3621 19717 3655
rect 19751 3652 19763 3655
rect 21358 3652 21364 3664
rect 19751 3624 21364 3652
rect 19751 3621 19763 3624
rect 19705 3615 19763 3621
rect 21358 3612 21364 3624
rect 21416 3612 21422 3664
rect 16899 3556 17080 3584
rect 17129 3587 17187 3593
rect 16899 3553 16911 3556
rect 16853 3547 16911 3553
rect 17129 3553 17141 3587
rect 17175 3584 17187 3587
rect 17175 3556 17724 3584
rect 17175 3553 17187 3556
rect 17129 3547 17187 3553
rect 14277 3519 14335 3525
rect 12268 3488 14228 3516
rect 9125 3479 9183 3485
rect 9140 3380 9168 3479
rect 14200 3448 14228 3488
rect 14277 3485 14289 3519
rect 14323 3516 14335 3519
rect 14458 3516 14464 3528
rect 14323 3488 14464 3516
rect 14323 3485 14335 3488
rect 14277 3479 14335 3485
rect 14458 3476 14464 3488
rect 14516 3476 14522 3528
rect 15212 3510 15424 3516
rect 15470 3510 15476 3528
rect 15212 3488 15476 3510
rect 15212 3448 15240 3488
rect 15396 3482 15476 3488
rect 15470 3476 15476 3482
rect 15528 3476 15534 3528
rect 15565 3519 15623 3525
rect 15565 3485 15577 3519
rect 15611 3516 15623 3519
rect 15654 3516 15660 3528
rect 15611 3488 15660 3516
rect 15611 3485 15623 3488
rect 15565 3479 15623 3485
rect 15654 3476 15660 3488
rect 15712 3476 15718 3528
rect 17589 3519 17647 3525
rect 17589 3485 17601 3519
rect 17635 3485 17647 3519
rect 17589 3479 17647 3485
rect 14200 3420 15240 3448
rect 15396 3420 16068 3448
rect 15396 3380 15424 3420
rect 9140 3352 15424 3380
rect 16040 3380 16068 3420
rect 16298 3380 16304 3392
rect 16040 3352 16304 3380
rect 16298 3340 16304 3352
rect 16356 3340 16362 3392
rect 17604 3380 17632 3479
rect 17696 3448 17724 3556
rect 17770 3544 17776 3596
rect 17828 3544 17834 3596
rect 19794 3584 19800 3596
rect 19536 3556 19800 3584
rect 18046 3476 18052 3528
rect 18104 3516 18110 3528
rect 19426 3516 19432 3528
rect 18104 3488 19432 3516
rect 18104 3476 18110 3488
rect 19426 3476 19432 3488
rect 19484 3476 19490 3528
rect 19536 3525 19564 3556
rect 19794 3544 19800 3556
rect 19852 3544 19858 3596
rect 21269 3587 21327 3593
rect 21269 3584 21281 3587
rect 20732 3556 21281 3584
rect 19521 3519 19579 3525
rect 19521 3485 19533 3519
rect 19567 3485 19579 3519
rect 19521 3479 19579 3485
rect 19610 3476 19616 3528
rect 19668 3516 19674 3528
rect 20530 3516 20536 3528
rect 19668 3488 20536 3516
rect 19668 3476 19674 3488
rect 20530 3476 20536 3488
rect 20588 3476 20594 3528
rect 20732 3448 20760 3556
rect 21269 3553 21281 3556
rect 21315 3584 21327 3587
rect 21652 3584 21680 3692
rect 22002 3680 22008 3692
rect 22060 3680 22066 3732
rect 22094 3680 22100 3732
rect 22152 3720 22158 3732
rect 22281 3723 22339 3729
rect 22281 3720 22293 3723
rect 22152 3692 22293 3720
rect 22152 3680 22158 3692
rect 22281 3689 22293 3692
rect 22327 3689 22339 3723
rect 22281 3683 22339 3689
rect 22373 3723 22431 3729
rect 22373 3689 22385 3723
rect 22419 3720 22431 3723
rect 23014 3720 23020 3732
rect 22419 3692 23020 3720
rect 22419 3689 22431 3692
rect 22373 3683 22431 3689
rect 23014 3680 23020 3692
rect 23072 3680 23078 3732
rect 23290 3680 23296 3732
rect 23348 3720 23354 3732
rect 25866 3720 25872 3732
rect 23348 3692 23612 3720
rect 23348 3680 23354 3692
rect 22554 3652 22560 3664
rect 21744 3624 22560 3652
rect 21744 3593 21772 3624
rect 22554 3612 22560 3624
rect 22612 3612 22618 3664
rect 23584 3661 23612 3692
rect 23952 3692 25872 3720
rect 23569 3655 23627 3661
rect 23569 3621 23581 3655
rect 23615 3621 23627 3655
rect 23569 3615 23627 3621
rect 21315 3556 21680 3584
rect 21729 3587 21787 3593
rect 21315 3553 21327 3556
rect 21269 3547 21327 3553
rect 21729 3553 21741 3587
rect 21775 3553 21787 3587
rect 21729 3547 21787 3553
rect 22646 3544 22652 3596
rect 22704 3584 22710 3596
rect 23017 3587 23075 3593
rect 23017 3584 23029 3587
rect 22704 3556 23029 3584
rect 22704 3544 22710 3556
rect 23017 3553 23029 3556
rect 23063 3553 23075 3587
rect 23017 3547 23075 3553
rect 23176 3587 23234 3593
rect 23176 3553 23188 3587
rect 23222 3584 23234 3587
rect 23474 3584 23480 3596
rect 23222 3556 23480 3584
rect 23222 3553 23234 3556
rect 23176 3547 23234 3553
rect 23474 3544 23480 3556
rect 23532 3544 23538 3596
rect 21085 3519 21143 3525
rect 21085 3485 21097 3519
rect 21131 3516 21143 3519
rect 21634 3516 21640 3528
rect 21131 3488 21640 3516
rect 21131 3485 21143 3488
rect 21085 3479 21143 3485
rect 21634 3476 21640 3488
rect 21692 3476 21698 3528
rect 23290 3476 23296 3528
rect 23348 3476 23354 3528
rect 23952 3516 23980 3692
rect 25866 3680 25872 3692
rect 25924 3680 25930 3732
rect 30098 3680 30104 3732
rect 30156 3680 30162 3732
rect 30650 3680 30656 3732
rect 30708 3680 30714 3732
rect 31389 3723 31447 3729
rect 31389 3689 31401 3723
rect 31435 3720 31447 3723
rect 33410 3720 33416 3732
rect 31435 3692 33416 3720
rect 31435 3689 31447 3692
rect 31389 3683 31447 3689
rect 33410 3680 33416 3692
rect 33468 3680 33474 3732
rect 35529 3723 35587 3729
rect 35529 3689 35541 3723
rect 35575 3720 35587 3723
rect 35710 3720 35716 3732
rect 35575 3692 35716 3720
rect 35575 3689 35587 3692
rect 35529 3683 35587 3689
rect 35710 3680 35716 3692
rect 35768 3680 35774 3732
rect 39390 3680 39396 3732
rect 39448 3680 39454 3732
rect 24210 3612 24216 3664
rect 24268 3612 24274 3664
rect 24486 3612 24492 3664
rect 24544 3652 24550 3664
rect 26145 3655 26203 3661
rect 26145 3652 26157 3655
rect 24544 3624 26157 3652
rect 24544 3612 24550 3624
rect 26145 3621 26157 3624
rect 26191 3621 26203 3655
rect 26145 3615 26203 3621
rect 38105 3655 38163 3661
rect 38105 3621 38117 3655
rect 38151 3652 38163 3655
rect 38378 3652 38384 3664
rect 38151 3624 38384 3652
rect 38151 3621 38163 3624
rect 38105 3615 38163 3621
rect 38378 3612 38384 3624
rect 38436 3612 38442 3664
rect 24029 3587 24087 3593
rect 24029 3553 24041 3587
rect 24075 3584 24087 3587
rect 24228 3584 24256 3612
rect 24075 3556 24256 3584
rect 24320 3556 30512 3584
rect 24075 3553 24087 3556
rect 24029 3547 24087 3553
rect 24213 3519 24271 3525
rect 24213 3516 24225 3519
rect 23952 3488 24225 3516
rect 24213 3485 24225 3488
rect 24259 3485 24271 3519
rect 24213 3479 24271 3485
rect 17696 3420 20760 3448
rect 20806 3408 20812 3460
rect 20864 3448 20870 3460
rect 21177 3451 21235 3457
rect 21177 3448 21189 3451
rect 20864 3420 21189 3448
rect 20864 3408 20870 3420
rect 21177 3417 21189 3420
rect 21223 3417 21235 3451
rect 21177 3411 21235 3417
rect 21913 3451 21971 3457
rect 21913 3417 21925 3451
rect 21959 3448 21971 3451
rect 22278 3448 22284 3460
rect 21959 3420 22284 3448
rect 21959 3417 21971 3420
rect 21913 3411 21971 3417
rect 22278 3408 22284 3420
rect 22336 3408 22342 3460
rect 18690 3380 18696 3392
rect 17604 3352 18696 3380
rect 18690 3340 18696 3352
rect 18748 3340 18754 3392
rect 19334 3340 19340 3392
rect 19392 3340 19398 3392
rect 21821 3383 21879 3389
rect 21821 3349 21833 3383
rect 21867 3380 21879 3383
rect 23474 3380 23480 3392
rect 21867 3352 23480 3380
rect 21867 3349 21879 3352
rect 21821 3343 21879 3349
rect 23474 3340 23480 3352
rect 23532 3340 23538 3392
rect 23566 3340 23572 3392
rect 23624 3380 23630 3392
rect 24320 3380 24348 3556
rect 29914 3476 29920 3528
rect 29972 3476 29978 3528
rect 30484 3525 30512 3556
rect 37458 3544 37464 3596
rect 37516 3584 37522 3596
rect 37516 3556 38516 3584
rect 37516 3544 37522 3556
rect 30469 3519 30527 3525
rect 30469 3485 30481 3519
rect 30515 3485 30527 3519
rect 30469 3479 30527 3485
rect 31202 3476 31208 3528
rect 31260 3476 31266 3528
rect 35437 3519 35495 3525
rect 35437 3485 35449 3519
rect 35483 3516 35495 3519
rect 35713 3519 35771 3525
rect 35713 3516 35725 3519
rect 35483 3488 35725 3516
rect 35483 3485 35495 3488
rect 35437 3479 35495 3485
rect 35713 3485 35725 3488
rect 35759 3485 35771 3519
rect 35713 3479 35771 3485
rect 35802 3476 35808 3528
rect 35860 3516 35866 3528
rect 38488 3525 38516 3556
rect 37645 3519 37703 3525
rect 37645 3516 37657 3519
rect 35860 3488 37657 3516
rect 35860 3476 35866 3488
rect 37645 3485 37657 3488
rect 37691 3485 37703 3519
rect 37645 3479 37703 3485
rect 37829 3519 37887 3525
rect 37829 3485 37841 3519
rect 37875 3516 37887 3519
rect 37921 3519 37979 3525
rect 37921 3516 37933 3519
rect 37875 3488 37933 3516
rect 37875 3485 37887 3488
rect 37829 3479 37887 3485
rect 37921 3485 37933 3488
rect 37967 3485 37979 3519
rect 37921 3479 37979 3485
rect 38381 3519 38439 3525
rect 38381 3485 38393 3519
rect 38427 3485 38439 3519
rect 38381 3479 38439 3485
rect 38473 3519 38531 3525
rect 38473 3485 38485 3519
rect 38519 3516 38531 3519
rect 38933 3519 38991 3525
rect 38933 3516 38945 3519
rect 38519 3488 38945 3516
rect 38519 3485 38531 3488
rect 38473 3479 38531 3485
rect 38933 3485 38945 3488
rect 38979 3485 38991 3519
rect 38933 3479 38991 3485
rect 26326 3408 26332 3460
rect 26384 3408 26390 3460
rect 34514 3408 34520 3460
rect 34572 3448 34578 3460
rect 38396 3448 38424 3479
rect 39206 3476 39212 3528
rect 39264 3476 39270 3528
rect 38749 3451 38807 3457
rect 38749 3448 38761 3451
rect 34572 3420 38761 3448
rect 34572 3408 34578 3420
rect 38749 3417 38761 3420
rect 38795 3417 38807 3451
rect 38749 3411 38807 3417
rect 23624 3352 24348 3380
rect 23624 3340 23630 3352
rect 35342 3340 35348 3392
rect 35400 3340 35406 3392
rect 37366 3340 37372 3392
rect 37424 3380 37430 3392
rect 37461 3383 37519 3389
rect 37461 3380 37473 3383
rect 37424 3352 37473 3380
rect 37424 3340 37430 3352
rect 37461 3349 37473 3352
rect 37507 3349 37519 3383
rect 37461 3343 37519 3349
rect 37734 3340 37740 3392
rect 37792 3340 37798 3392
rect 38197 3383 38255 3389
rect 38197 3349 38209 3383
rect 38243 3380 38255 3383
rect 38286 3380 38292 3392
rect 38243 3352 38292 3380
rect 38243 3349 38255 3352
rect 38197 3343 38255 3349
rect 38286 3340 38292 3352
rect 38344 3340 38350 3392
rect 38654 3340 38660 3392
rect 38712 3340 38718 3392
rect 1104 3290 39836 3312
rect 1104 3238 3010 3290
rect 3062 3238 3074 3290
rect 3126 3238 3138 3290
rect 3190 3238 3202 3290
rect 3254 3238 3266 3290
rect 3318 3238 9010 3290
rect 9062 3238 9074 3290
rect 9126 3238 9138 3290
rect 9190 3238 9202 3290
rect 9254 3238 9266 3290
rect 9318 3238 15010 3290
rect 15062 3238 15074 3290
rect 15126 3238 15138 3290
rect 15190 3238 15202 3290
rect 15254 3238 15266 3290
rect 15318 3238 21010 3290
rect 21062 3238 21074 3290
rect 21126 3238 21138 3290
rect 21190 3238 21202 3290
rect 21254 3238 21266 3290
rect 21318 3238 27010 3290
rect 27062 3238 27074 3290
rect 27126 3238 27138 3290
rect 27190 3238 27202 3290
rect 27254 3238 27266 3290
rect 27318 3238 33010 3290
rect 33062 3238 33074 3290
rect 33126 3238 33138 3290
rect 33190 3238 33202 3290
rect 33254 3238 33266 3290
rect 33318 3238 39010 3290
rect 39062 3238 39074 3290
rect 39126 3238 39138 3290
rect 39190 3238 39202 3290
rect 39254 3238 39266 3290
rect 39318 3238 39836 3290
rect 1104 3216 39836 3238
rect 3510 3136 3516 3188
rect 3568 3176 3574 3188
rect 15194 3176 15200 3188
rect 3568 3148 15200 3176
rect 3568 3136 3574 3148
rect 15194 3136 15200 3148
rect 15252 3136 15258 3188
rect 22186 3136 22192 3188
rect 22244 3176 22250 3188
rect 22465 3179 22523 3185
rect 22465 3176 22477 3179
rect 22244 3148 22477 3176
rect 22244 3136 22250 3148
rect 22465 3145 22477 3148
rect 22511 3145 22523 3179
rect 22465 3139 22523 3145
rect 39025 3179 39083 3185
rect 39025 3145 39037 3179
rect 39071 3176 39083 3179
rect 39390 3176 39396 3188
rect 39071 3148 39396 3176
rect 39071 3145 39083 3148
rect 39025 3139 39083 3145
rect 39390 3136 39396 3148
rect 39448 3136 39454 3188
rect 7006 3068 7012 3120
rect 7064 3108 7070 3120
rect 19334 3108 19340 3120
rect 7064 3080 19340 3108
rect 7064 3068 7070 3080
rect 19334 3068 19340 3080
rect 19392 3068 19398 3120
rect 21545 3111 21603 3117
rect 21545 3077 21557 3111
rect 21591 3108 21603 3111
rect 23106 3108 23112 3120
rect 21591 3080 23112 3108
rect 21591 3077 21603 3080
rect 21545 3071 21603 3077
rect 23106 3068 23112 3080
rect 23164 3068 23170 3120
rect 20898 3000 20904 3052
rect 20956 3040 20962 3052
rect 21453 3043 21511 3049
rect 21453 3040 21465 3043
rect 20956 3012 21465 3040
rect 20956 3000 20962 3012
rect 21453 3009 21465 3012
rect 21499 3009 21511 3043
rect 21453 3003 21511 3009
rect 22554 3000 22560 3052
rect 22612 3040 22618 3052
rect 22679 3043 22737 3049
rect 22679 3040 22691 3043
rect 22612 3012 22691 3040
rect 22612 3000 22618 3012
rect 22679 3009 22691 3012
rect 22725 3009 22737 3043
rect 22679 3003 22737 3009
rect 22833 3043 22891 3049
rect 22833 3009 22845 3043
rect 22879 3040 22891 3043
rect 22922 3040 22928 3052
rect 22879 3012 22928 3040
rect 22879 3009 22891 3012
rect 22833 3003 22891 3009
rect 22922 3000 22928 3012
rect 22980 3000 22986 3052
rect 38470 3000 38476 3052
rect 38528 3000 38534 3052
rect 38838 3000 38844 3052
rect 38896 3000 38902 3052
rect 39206 3000 39212 3052
rect 39264 3000 39270 3052
rect 22002 2932 22008 2984
rect 22060 2972 22066 2984
rect 35342 2972 35348 2984
rect 22060 2944 35348 2972
rect 22060 2932 22066 2944
rect 35342 2932 35348 2944
rect 35400 2932 35406 2984
rect 13722 2864 13728 2916
rect 13780 2904 13786 2916
rect 23198 2904 23204 2916
rect 13780 2876 23204 2904
rect 13780 2864 13786 2876
rect 23198 2864 23204 2876
rect 23256 2864 23262 2916
rect 39393 2907 39451 2913
rect 39393 2873 39405 2907
rect 39439 2904 39451 2907
rect 39482 2904 39488 2916
rect 39439 2876 39488 2904
rect 39439 2873 39451 2876
rect 39393 2867 39451 2873
rect 39482 2864 39488 2876
rect 39540 2864 39546 2916
rect 9858 2796 9864 2848
rect 9916 2836 9922 2848
rect 19242 2836 19248 2848
rect 9916 2808 19248 2836
rect 9916 2796 9922 2808
rect 19242 2796 19248 2808
rect 19300 2836 19306 2848
rect 26326 2836 26332 2848
rect 19300 2808 26332 2836
rect 19300 2796 19306 2808
rect 26326 2796 26332 2808
rect 26384 2796 26390 2848
rect 38657 2839 38715 2845
rect 38657 2805 38669 2839
rect 38703 2836 38715 2839
rect 38838 2836 38844 2848
rect 38703 2808 38844 2836
rect 38703 2805 38715 2808
rect 38657 2799 38715 2805
rect 38838 2796 38844 2808
rect 38896 2796 38902 2848
rect 1104 2746 39836 2768
rect 1104 2694 1950 2746
rect 2002 2694 2014 2746
rect 2066 2694 2078 2746
rect 2130 2694 2142 2746
rect 2194 2694 2206 2746
rect 2258 2694 7950 2746
rect 8002 2694 8014 2746
rect 8066 2694 8078 2746
rect 8130 2694 8142 2746
rect 8194 2694 8206 2746
rect 8258 2694 13950 2746
rect 14002 2694 14014 2746
rect 14066 2694 14078 2746
rect 14130 2694 14142 2746
rect 14194 2694 14206 2746
rect 14258 2694 19950 2746
rect 20002 2694 20014 2746
rect 20066 2694 20078 2746
rect 20130 2694 20142 2746
rect 20194 2694 20206 2746
rect 20258 2694 25950 2746
rect 26002 2694 26014 2746
rect 26066 2694 26078 2746
rect 26130 2694 26142 2746
rect 26194 2694 26206 2746
rect 26258 2694 31950 2746
rect 32002 2694 32014 2746
rect 32066 2694 32078 2746
rect 32130 2694 32142 2746
rect 32194 2694 32206 2746
rect 32258 2694 37950 2746
rect 38002 2694 38014 2746
rect 38066 2694 38078 2746
rect 38130 2694 38142 2746
rect 38194 2694 38206 2746
rect 38258 2694 39836 2746
rect 1104 2672 39836 2694
rect 6914 2592 6920 2644
rect 6972 2632 6978 2644
rect 38930 2632 38936 2644
rect 6972 2604 38936 2632
rect 6972 2592 6978 2604
rect 38930 2592 38936 2604
rect 38988 2592 38994 2644
rect 39390 2592 39396 2644
rect 39448 2592 39454 2644
rect 1302 2524 1308 2576
rect 1360 2564 1366 2576
rect 35802 2564 35808 2576
rect 1360 2536 35808 2564
rect 1360 2524 1366 2536
rect 35802 2524 35808 2536
rect 35860 2524 35866 2576
rect 37550 2524 37556 2576
rect 37608 2524 37614 2576
rect 39025 2567 39083 2573
rect 39025 2533 39037 2567
rect 39071 2564 39083 2567
rect 39942 2564 39948 2576
rect 39071 2536 39948 2564
rect 39071 2533 39083 2536
rect 39025 2527 39083 2533
rect 39942 2524 39948 2536
rect 40000 2524 40006 2576
rect 14826 2496 14832 2508
rect 5184 2468 14832 2496
rect 1673 2431 1731 2437
rect 1673 2397 1685 2431
rect 1719 2428 1731 2431
rect 2038 2428 2044 2440
rect 1719 2400 2044 2428
rect 1719 2397 1731 2400
rect 1673 2391 1731 2397
rect 2038 2388 2044 2400
rect 2096 2388 2102 2440
rect 5184 2437 5212 2468
rect 14826 2456 14832 2468
rect 14884 2456 14890 2508
rect 15194 2456 15200 2508
rect 15252 2496 15258 2508
rect 38286 2496 38292 2508
rect 15252 2468 22094 2496
rect 15252 2456 15258 2468
rect 3605 2431 3663 2437
rect 3605 2397 3617 2431
rect 3651 2397 3663 2431
rect 3605 2391 3663 2397
rect 5169 2431 5227 2437
rect 5169 2397 5181 2431
rect 5215 2397 5227 2431
rect 5169 2391 5227 2397
rect 3620 2360 3648 2391
rect 6730 2388 6736 2440
rect 6788 2388 6794 2440
rect 9490 2388 9496 2440
rect 9548 2428 9554 2440
rect 9585 2431 9643 2437
rect 9585 2428 9597 2431
rect 9548 2400 9597 2428
rect 9548 2388 9554 2400
rect 9585 2397 9597 2400
rect 9631 2397 9643 2431
rect 9585 2391 9643 2397
rect 9858 2388 9864 2440
rect 9916 2388 9922 2440
rect 5534 2360 5540 2372
rect 3620 2332 5540 2360
rect 5534 2320 5540 2332
rect 5592 2320 5598 2372
rect 22066 2360 22094 2468
rect 38028 2468 38292 2496
rect 37366 2388 37372 2440
rect 37424 2388 37430 2440
rect 38028 2437 38056 2468
rect 38286 2456 38292 2468
rect 38344 2456 38350 2508
rect 38013 2431 38071 2437
rect 38013 2397 38025 2431
rect 38059 2397 38071 2431
rect 38013 2391 38071 2397
rect 38105 2431 38163 2437
rect 38105 2397 38117 2431
rect 38151 2397 38163 2431
rect 38105 2391 38163 2397
rect 38120 2360 38148 2391
rect 38378 2388 38384 2440
rect 38436 2428 38442 2440
rect 38473 2431 38531 2437
rect 38473 2428 38485 2431
rect 38436 2400 38485 2428
rect 38436 2388 38442 2400
rect 38473 2397 38485 2400
rect 38519 2397 38531 2431
rect 38473 2391 38531 2397
rect 38746 2388 38752 2440
rect 38804 2428 38810 2440
rect 38841 2431 38899 2437
rect 38841 2428 38853 2431
rect 38804 2400 38853 2428
rect 38804 2388 38810 2400
rect 38841 2397 38853 2400
rect 38887 2397 38899 2431
rect 38841 2391 38899 2397
rect 39209 2431 39267 2437
rect 39209 2397 39221 2431
rect 39255 2428 39267 2431
rect 39255 2400 39896 2428
rect 39255 2397 39267 2400
rect 39209 2391 39267 2397
rect 22066 2332 38148 2360
rect 1670 2252 1676 2304
rect 1728 2292 1734 2304
rect 1857 2295 1915 2301
rect 1857 2292 1869 2295
rect 1728 2264 1869 2292
rect 1728 2252 1734 2264
rect 1857 2261 1869 2264
rect 1903 2261 1915 2295
rect 1857 2255 1915 2261
rect 3418 2252 3424 2304
rect 3476 2252 3482 2304
rect 4798 2252 4804 2304
rect 4856 2292 4862 2304
rect 4985 2295 5043 2301
rect 4985 2292 4997 2295
rect 4856 2264 4997 2292
rect 4856 2252 4862 2264
rect 4985 2261 4997 2264
rect 5031 2261 5043 2295
rect 4985 2255 5043 2261
rect 6362 2252 6368 2304
rect 6420 2292 6426 2304
rect 6549 2295 6607 2301
rect 6549 2292 6561 2295
rect 6420 2264 6561 2292
rect 6420 2252 6426 2264
rect 6549 2261 6561 2264
rect 6595 2261 6607 2295
rect 6549 2255 6607 2261
rect 37826 2252 37832 2304
rect 37884 2252 37890 2304
rect 38286 2252 38292 2304
rect 38344 2252 38350 2304
rect 38654 2252 38660 2304
rect 38712 2252 38718 2304
rect 1104 2202 39836 2224
rect 1104 2150 3010 2202
rect 3062 2150 3074 2202
rect 3126 2150 3138 2202
rect 3190 2150 3202 2202
rect 3254 2150 3266 2202
rect 3318 2150 9010 2202
rect 9062 2150 9074 2202
rect 9126 2150 9138 2202
rect 9190 2150 9202 2202
rect 9254 2150 9266 2202
rect 9318 2150 15010 2202
rect 15062 2150 15074 2202
rect 15126 2150 15138 2202
rect 15190 2150 15202 2202
rect 15254 2150 15266 2202
rect 15318 2150 21010 2202
rect 21062 2150 21074 2202
rect 21126 2150 21138 2202
rect 21190 2150 21202 2202
rect 21254 2150 21266 2202
rect 21318 2150 27010 2202
rect 27062 2150 27074 2202
rect 27126 2150 27138 2202
rect 27190 2150 27202 2202
rect 27254 2150 27266 2202
rect 27318 2150 33010 2202
rect 33062 2150 33074 2202
rect 33126 2150 33138 2202
rect 33190 2150 33202 2202
rect 33254 2150 33266 2202
rect 33318 2150 39010 2202
rect 39062 2150 39074 2202
rect 39126 2150 39138 2202
rect 39190 2150 39202 2202
rect 39254 2150 39266 2202
rect 39318 2150 39836 2202
rect 1104 2128 39836 2150
rect 6730 2048 6736 2100
rect 6788 2088 6794 2100
rect 17494 2088 17500 2100
rect 6788 2060 17500 2088
rect 6788 2048 6794 2060
rect 17494 2048 17500 2060
rect 17552 2048 17558 2100
rect 20438 2048 20444 2100
rect 20496 2088 20502 2100
rect 31202 2088 31208 2100
rect 20496 2060 31208 2088
rect 20496 2048 20502 2060
rect 31202 2048 31208 2060
rect 31260 2048 31266 2100
rect 4706 1980 4712 2032
rect 4764 2020 4770 2032
rect 39868 2020 39896 2400
rect 4764 1992 39896 2020
rect 4764 1980 4770 1992
rect 25130 824 25136 876
rect 25188 864 25194 876
rect 26878 864 26884 876
rect 25188 836 26884 864
rect 25188 824 25194 836
rect 26878 824 26884 836
rect 26936 824 26942 876
rect 14182 144 14188 196
rect 14240 184 14246 196
rect 25038 184 25044 196
rect 14240 156 25044 184
rect 14240 144 14246 156
rect 25038 144 25044 156
rect 25096 144 25102 196
rect 18966 76 18972 128
rect 19024 116 19030 128
rect 31570 116 31576 128
rect 19024 88 31576 116
rect 19024 76 19030 88
rect 31570 76 31576 88
rect 31628 76 31634 128
rect 8018 8 8024 60
rect 8076 48 8082 60
rect 29914 48 29920 60
rect 8076 20 29920 48
rect 8076 8 8082 20
rect 29914 8 29920 20
rect 29972 8 29978 60
<< via1 >>
rect 3884 11160 3936 11212
rect 20076 11160 20128 11212
rect 7840 11092 7892 11144
rect 20904 11092 20956 11144
rect 9772 11024 9824 11076
rect 20628 11024 20680 11076
rect 7196 10072 7248 10124
rect 26792 10072 26844 10124
rect 10600 10004 10652 10056
rect 24124 10004 24176 10056
rect 14648 9936 14700 9988
rect 29920 9936 29972 9988
rect 10876 9868 10928 9920
rect 26608 9868 26660 9920
rect 10048 9800 10100 9852
rect 28540 9800 28592 9852
rect 9496 9732 9548 9784
rect 28724 9732 28776 9784
rect 7748 9664 7800 9716
rect 17132 9664 17184 9716
rect 5816 9596 5868 9648
rect 15568 9596 15620 9648
rect 10324 9528 10376 9580
rect 19340 9528 19392 9580
rect 2688 9460 2740 9512
rect 14464 9460 14516 9512
rect 16672 9460 16724 9512
rect 24400 9460 24452 9512
rect 16028 9392 16080 9444
rect 22100 9392 22152 9444
rect 15476 9324 15528 9376
rect 23480 9324 23532 9376
rect 6920 9256 6972 9308
rect 17500 9256 17552 9308
rect 19064 9256 19116 9308
rect 32588 9256 32640 9308
rect 7564 9188 7616 9240
rect 25228 9188 25280 9240
rect 2136 9120 2188 9172
rect 20444 9120 20496 9172
rect 22652 9120 22704 9172
rect 23848 9120 23900 9172
rect 2044 8984 2096 9036
rect 12440 9052 12492 9104
rect 13820 9052 13872 9104
rect 8392 8984 8444 9036
rect 16580 8984 16632 9036
rect 664 8916 716 8968
rect 16396 8916 16448 8968
rect 2412 8848 2464 8900
rect 6736 8848 6788 8900
rect 7288 8848 7340 8900
rect 15752 8848 15804 8900
rect 17960 9052 18012 9104
rect 23204 9052 23256 9104
rect 17224 8984 17276 9036
rect 18788 8916 18840 8968
rect 22652 8916 22704 8968
rect 25872 8984 25924 9036
rect 27896 8984 27948 9036
rect 30472 8916 30524 8968
rect 30656 8916 30708 8968
rect 33784 8916 33836 8968
rect 25504 8848 25556 8900
rect 32404 8848 32456 8900
rect 35072 8848 35124 8900
rect 1584 8780 1636 8832
rect 8576 8780 8628 8832
rect 12532 8780 12584 8832
rect 14740 8780 14792 8832
rect 19708 8780 19760 8832
rect 23756 8780 23808 8832
rect 26148 8780 26200 8832
rect 28448 8780 28500 8832
rect 33048 8780 33100 8832
rect 33508 8780 33560 8832
rect 34980 8780 35032 8832
rect 35624 8780 35676 8832
rect 3010 8678 3062 8730
rect 3074 8678 3126 8730
rect 3138 8678 3190 8730
rect 3202 8678 3254 8730
rect 3266 8678 3318 8730
rect 9010 8678 9062 8730
rect 9074 8678 9126 8730
rect 9138 8678 9190 8730
rect 9202 8678 9254 8730
rect 9266 8678 9318 8730
rect 15010 8678 15062 8730
rect 15074 8678 15126 8730
rect 15138 8678 15190 8730
rect 15202 8678 15254 8730
rect 15266 8678 15318 8730
rect 21010 8678 21062 8730
rect 21074 8678 21126 8730
rect 21138 8678 21190 8730
rect 21202 8678 21254 8730
rect 21266 8678 21318 8730
rect 27010 8678 27062 8730
rect 27074 8678 27126 8730
rect 27138 8678 27190 8730
rect 27202 8678 27254 8730
rect 27266 8678 27318 8730
rect 33010 8678 33062 8730
rect 33074 8678 33126 8730
rect 33138 8678 33190 8730
rect 33202 8678 33254 8730
rect 33266 8678 33318 8730
rect 39010 8678 39062 8730
rect 39074 8678 39126 8730
rect 39138 8678 39190 8730
rect 39202 8678 39254 8730
rect 39266 8678 39318 8730
rect 1124 8576 1176 8628
rect 1308 8508 1360 8560
rect 572 8440 624 8492
rect 848 8372 900 8424
rect 1032 8304 1084 8356
rect 2412 8619 2464 8628
rect 2412 8585 2421 8619
rect 2421 8585 2455 8619
rect 2455 8585 2464 8619
rect 2412 8576 2464 8585
rect 2688 8619 2740 8628
rect 2688 8585 2697 8619
rect 2697 8585 2731 8619
rect 2731 8585 2740 8619
rect 2688 8576 2740 8585
rect 3792 8576 3844 8628
rect 4344 8576 4396 8628
rect 4620 8619 4672 8628
rect 4620 8585 4629 8619
rect 4629 8585 4663 8619
rect 4663 8585 4672 8619
rect 4620 8576 4672 8585
rect 5172 8576 5224 8628
rect 5448 8576 5500 8628
rect 5724 8576 5776 8628
rect 6276 8576 6328 8628
rect 6828 8576 6880 8628
rect 7380 8576 7432 8628
rect 7656 8576 7708 8628
rect 7932 8576 7984 8628
rect 8484 8576 8536 8628
rect 8852 8576 8904 8628
rect 9588 8576 9640 8628
rect 9864 8576 9916 8628
rect 10140 8576 10192 8628
rect 10692 8576 10744 8628
rect 10968 8576 11020 8628
rect 11520 8576 11572 8628
rect 11980 8576 12032 8628
rect 12348 8576 12400 8628
rect 13176 8576 13228 8628
rect 14004 8576 14056 8628
rect 14556 8576 14608 8628
rect 14924 8576 14976 8628
rect 15384 8576 15436 8628
rect 15660 8619 15712 8628
rect 15660 8585 15669 8619
rect 15669 8585 15703 8619
rect 15703 8585 15712 8619
rect 15660 8576 15712 8585
rect 16212 8576 16264 8628
rect 16488 8576 16540 8628
rect 16764 8576 16816 8628
rect 17316 8576 17368 8628
rect 18788 8619 18840 8628
rect 18788 8585 18797 8619
rect 18797 8585 18831 8619
rect 18831 8585 18840 8619
rect 18788 8576 18840 8585
rect 19340 8619 19392 8628
rect 19340 8585 19349 8619
rect 19349 8585 19383 8619
rect 19383 8585 19392 8619
rect 19340 8576 19392 8585
rect 19524 8576 19576 8628
rect 19616 8619 19668 8628
rect 19616 8585 19625 8619
rect 19625 8585 19659 8619
rect 19659 8585 19668 8619
rect 19616 8576 19668 8585
rect 20536 8576 20588 8628
rect 22008 8576 22060 8628
rect 7748 8508 7800 8560
rect 2044 8304 2096 8356
rect 2136 8347 2188 8356
rect 2136 8313 2145 8347
rect 2145 8313 2179 8347
rect 2179 8313 2188 8347
rect 2136 8304 2188 8313
rect 3516 8304 3568 8356
rect 3700 8440 3752 8492
rect 3976 8372 4028 8424
rect 4528 8440 4580 8492
rect 5632 8440 5684 8492
rect 5816 8483 5868 8492
rect 5816 8449 5825 8483
rect 5825 8449 5859 8483
rect 5859 8449 5868 8483
rect 5816 8440 5868 8449
rect 6920 8483 6972 8492
rect 6920 8449 6929 8483
rect 6929 8449 6963 8483
rect 6963 8449 6972 8483
rect 6920 8440 6972 8449
rect 7288 8483 7340 8492
rect 7288 8449 7297 8483
rect 7297 8449 7331 8483
rect 7331 8449 7340 8483
rect 7288 8440 7340 8449
rect 7656 8483 7708 8492
rect 7656 8449 7665 8483
rect 7665 8449 7699 8483
rect 7699 8449 7708 8483
rect 7656 8440 7708 8449
rect 7012 8372 7064 8424
rect 11612 8508 11664 8560
rect 8392 8483 8444 8492
rect 8392 8449 8401 8483
rect 8401 8449 8435 8483
rect 8435 8449 8444 8483
rect 8392 8440 8444 8449
rect 8668 8440 8720 8492
rect 9496 8483 9548 8492
rect 9496 8449 9505 8483
rect 9505 8449 9539 8483
rect 9539 8449 9548 8483
rect 9496 8440 9548 8449
rect 10048 8440 10100 8492
rect 10232 8483 10284 8492
rect 10232 8449 10241 8483
rect 10241 8449 10275 8483
rect 10275 8449 10284 8483
rect 10232 8440 10284 8449
rect 10600 8483 10652 8492
rect 10600 8449 10609 8483
rect 10609 8449 10643 8483
rect 10643 8449 10652 8483
rect 10600 8440 10652 8449
rect 10876 8440 10928 8492
rect 12532 8508 12584 8560
rect 14740 8508 14792 8560
rect 8484 8372 8536 8424
rect 12992 8483 13044 8492
rect 12992 8449 13001 8483
rect 13001 8449 13035 8483
rect 13035 8449 13044 8483
rect 12992 8440 13044 8449
rect 13360 8483 13412 8492
rect 13360 8449 13369 8483
rect 13369 8449 13403 8483
rect 13403 8449 13412 8483
rect 13360 8440 13412 8449
rect 13544 8372 13596 8424
rect 14648 8483 14700 8492
rect 14648 8449 14657 8483
rect 14657 8449 14691 8483
rect 14691 8449 14700 8483
rect 14648 8440 14700 8449
rect 17224 8508 17276 8560
rect 15384 8483 15436 8492
rect 15384 8449 15393 8483
rect 15393 8449 15427 8483
rect 15427 8449 15436 8483
rect 15384 8440 15436 8449
rect 15844 8440 15896 8492
rect 16120 8483 16172 8492
rect 16120 8449 16129 8483
rect 16129 8449 16163 8483
rect 16163 8449 16172 8483
rect 16120 8440 16172 8449
rect 16672 8440 16724 8492
rect 16856 8483 16908 8492
rect 16856 8449 16865 8483
rect 16865 8449 16899 8483
rect 16899 8449 16908 8483
rect 16856 8440 16908 8449
rect 17408 8483 17460 8492
rect 17408 8449 17417 8483
rect 17417 8449 17451 8483
rect 17451 8449 17460 8483
rect 17408 8440 17460 8449
rect 18052 8440 18104 8492
rect 18420 8440 18472 8492
rect 18696 8440 18748 8492
rect 18972 8440 19024 8492
rect 19248 8440 19300 8492
rect 21732 8508 21784 8560
rect 19892 8483 19944 8492
rect 19892 8449 19901 8483
rect 19901 8449 19935 8483
rect 19935 8449 19944 8483
rect 19892 8440 19944 8449
rect 21364 8440 21416 8492
rect 21548 8440 21600 8492
rect 23112 8576 23164 8628
rect 22560 8508 22612 8560
rect 22468 8440 22520 8492
rect 23756 8619 23808 8628
rect 23756 8585 23765 8619
rect 23765 8585 23799 8619
rect 23799 8585 23808 8619
rect 23756 8576 23808 8585
rect 23940 8576 23992 8628
rect 23664 8508 23716 8560
rect 24768 8576 24820 8628
rect 24676 8508 24728 8560
rect 25504 8619 25556 8628
rect 25504 8585 25513 8619
rect 25513 8585 25547 8619
rect 25547 8585 25556 8619
rect 25504 8576 25556 8585
rect 25688 8576 25740 8628
rect 32220 8576 32272 8628
rect 32496 8576 32548 8628
rect 32864 8576 32916 8628
rect 33508 8619 33560 8628
rect 33508 8585 33517 8619
rect 33517 8585 33551 8619
rect 33551 8585 33560 8619
rect 33508 8576 33560 8585
rect 33600 8576 33652 8628
rect 34704 8576 34756 8628
rect 35808 8576 35860 8628
rect 36912 8576 36964 8628
rect 25320 8508 25372 8560
rect 26516 8508 26568 8560
rect 15108 8372 15160 8424
rect 17684 8372 17736 8424
rect 11980 8304 12032 8356
rect 12900 8304 12952 8356
rect 13728 8304 13780 8356
rect 17040 8304 17092 8356
rect 19800 8304 19852 8356
rect 21640 8304 21692 8356
rect 22100 8347 22152 8356
rect 22100 8313 22109 8347
rect 22109 8313 22143 8347
rect 22143 8313 22152 8347
rect 22100 8304 22152 8313
rect 22468 8304 22520 8356
rect 22928 8372 22980 8424
rect 22836 8304 22888 8356
rect 23204 8347 23256 8356
rect 23204 8313 23213 8347
rect 23213 8313 23247 8347
rect 23247 8313 23256 8347
rect 23204 8304 23256 8313
rect 23388 8304 23440 8356
rect 24308 8372 24360 8424
rect 25044 8372 25096 8424
rect 27804 8440 27856 8492
rect 28172 8483 28224 8492
rect 28172 8449 28181 8483
rect 28181 8449 28215 8483
rect 28215 8449 28224 8483
rect 28172 8440 28224 8449
rect 28356 8440 28408 8492
rect 24032 8347 24084 8356
rect 24032 8313 24041 8347
rect 24041 8313 24075 8347
rect 24075 8313 24084 8347
rect 24032 8304 24084 8313
rect 24216 8304 24268 8356
rect 24768 8304 24820 8356
rect 25228 8347 25280 8356
rect 25228 8313 25237 8347
rect 25237 8313 25271 8347
rect 25271 8313 25280 8347
rect 25228 8304 25280 8313
rect 25320 8304 25372 8356
rect 29184 8372 29236 8424
rect 30932 8508 30984 8560
rect 29736 8440 29788 8492
rect 30104 8372 30156 8424
rect 32588 8483 32640 8492
rect 32588 8449 32597 8483
rect 32597 8449 32631 8483
rect 32631 8449 32640 8483
rect 32588 8440 32640 8449
rect 33048 8508 33100 8560
rect 33508 8440 33560 8492
rect 33784 8508 33836 8560
rect 34060 8483 34112 8492
rect 34060 8449 34069 8483
rect 34069 8449 34103 8483
rect 34103 8449 34112 8483
rect 34060 8440 34112 8449
rect 34704 8483 34756 8492
rect 34704 8449 34713 8483
rect 34713 8449 34747 8483
rect 34747 8449 34756 8483
rect 34704 8440 34756 8449
rect 35072 8483 35124 8492
rect 35072 8449 35081 8483
rect 35081 8449 35115 8483
rect 35115 8449 35124 8483
rect 35072 8440 35124 8449
rect 35256 8440 35308 8492
rect 34152 8372 34204 8424
rect 35716 8483 35768 8492
rect 35716 8449 35725 8483
rect 35725 8449 35759 8483
rect 35759 8449 35768 8483
rect 35716 8440 35768 8449
rect 35900 8508 35952 8560
rect 36176 8483 36228 8492
rect 36176 8449 36185 8483
rect 36185 8449 36219 8483
rect 36219 8449 36228 8483
rect 36176 8440 36228 8449
rect 36544 8483 36596 8492
rect 36544 8449 36553 8483
rect 36553 8449 36587 8483
rect 36587 8449 36596 8483
rect 36544 8440 36596 8449
rect 37464 8508 37516 8560
rect 1584 8279 1636 8288
rect 1584 8245 1593 8279
rect 1593 8245 1627 8279
rect 1627 8245 1636 8279
rect 1584 8236 1636 8245
rect 2320 8236 2372 8288
rect 12808 8236 12860 8288
rect 14556 8236 14608 8288
rect 20352 8236 20404 8288
rect 21732 8236 21784 8288
rect 22928 8279 22980 8288
rect 22928 8245 22937 8279
rect 22937 8245 22971 8279
rect 22971 8245 22980 8279
rect 22928 8236 22980 8245
rect 23572 8236 23624 8288
rect 23756 8236 23808 8288
rect 25780 8236 25832 8288
rect 26332 8304 26384 8356
rect 26884 8236 26936 8288
rect 33416 8304 33468 8356
rect 33968 8304 34020 8356
rect 35624 8304 35676 8356
rect 36360 8372 36412 8424
rect 36912 8372 36964 8424
rect 37832 8440 37884 8492
rect 38384 8483 38436 8492
rect 38384 8449 38393 8483
rect 38393 8449 38427 8483
rect 38427 8449 38436 8483
rect 38384 8440 38436 8449
rect 37188 8304 37240 8356
rect 39028 8347 39080 8356
rect 39028 8313 39037 8347
rect 39037 8313 39071 8347
rect 39071 8313 39080 8347
rect 39028 8304 39080 8313
rect 39396 8347 39448 8356
rect 39396 8313 39405 8347
rect 39405 8313 39439 8347
rect 39439 8313 39448 8347
rect 39396 8304 39448 8313
rect 1950 8134 2002 8186
rect 2014 8134 2066 8186
rect 2078 8134 2130 8186
rect 2142 8134 2194 8186
rect 2206 8134 2258 8186
rect 7950 8134 8002 8186
rect 8014 8134 8066 8186
rect 8078 8134 8130 8186
rect 8142 8134 8194 8186
rect 8206 8134 8258 8186
rect 13950 8134 14002 8186
rect 14014 8134 14066 8186
rect 14078 8134 14130 8186
rect 14142 8134 14194 8186
rect 14206 8134 14258 8186
rect 19950 8134 20002 8186
rect 20014 8134 20066 8186
rect 20078 8134 20130 8186
rect 20142 8134 20194 8186
rect 20206 8134 20258 8186
rect 25950 8134 26002 8186
rect 26014 8134 26066 8186
rect 26078 8134 26130 8186
rect 26142 8134 26194 8186
rect 26206 8134 26258 8186
rect 31950 8134 32002 8186
rect 32014 8134 32066 8186
rect 32078 8134 32130 8186
rect 32142 8134 32194 8186
rect 32206 8134 32258 8186
rect 37950 8134 38002 8186
rect 38014 8134 38066 8186
rect 38078 8134 38130 8186
rect 38142 8134 38194 8186
rect 38206 8134 38258 8186
rect 1216 8032 1268 8084
rect 1952 7964 2004 8016
rect 1032 7896 1084 7948
rect 756 7828 808 7880
rect 3424 8075 3476 8084
rect 3424 8041 3433 8075
rect 3433 8041 3467 8075
rect 3467 8041 3476 8075
rect 3424 8032 3476 8041
rect 3516 8032 3568 8084
rect 3884 8032 3936 8084
rect 4068 8032 4120 8084
rect 4896 8032 4948 8084
rect 6000 8032 6052 8084
rect 6552 8032 6604 8084
rect 7104 8032 7156 8084
rect 8300 8032 8352 8084
rect 8760 8032 8812 8084
rect 9404 8032 9456 8084
rect 10416 8032 10468 8084
rect 11244 8032 11296 8084
rect 11796 8032 11848 8084
rect 12624 8032 12676 8084
rect 13452 8032 13504 8084
rect 14280 8032 14332 8084
rect 14832 8032 14884 8084
rect 15936 8032 15988 8084
rect 17592 8032 17644 8084
rect 18052 8032 18104 8084
rect 20536 8032 20588 8084
rect 23388 8032 23440 8084
rect 6920 7964 6972 8016
rect 2136 7896 2188 7948
rect 3884 7896 3936 7948
rect 572 7760 624 7812
rect 3608 7871 3660 7880
rect 3608 7837 3617 7871
rect 3617 7837 3651 7871
rect 3651 7837 3660 7871
rect 3608 7828 3660 7837
rect 8208 7896 8260 7948
rect 11888 7964 11940 8016
rect 16856 7964 16908 8016
rect 20628 7964 20680 8016
rect 23020 7964 23072 8016
rect 23204 7964 23256 8016
rect 23756 7964 23808 8016
rect 28908 7964 28960 8016
rect 34428 8032 34480 8084
rect 35532 8032 35584 8084
rect 36084 8032 36136 8084
rect 36636 8032 36688 8084
rect 37740 8032 37792 8084
rect 38660 8075 38712 8084
rect 38660 8041 38669 8075
rect 38669 8041 38703 8075
rect 38703 8041 38712 8075
rect 38660 8032 38712 8041
rect 4712 7828 4764 7880
rect 6184 7760 6236 7812
rect 2136 7735 2188 7744
rect 2136 7701 2145 7735
rect 2145 7701 2179 7735
rect 2179 7701 2188 7735
rect 2136 7692 2188 7701
rect 6276 7692 6328 7744
rect 7196 7828 7248 7880
rect 8300 7871 8352 7880
rect 8300 7837 8309 7871
rect 8309 7837 8343 7871
rect 8343 7837 8352 7871
rect 8300 7828 8352 7837
rect 9220 7871 9272 7880
rect 9220 7837 9229 7871
rect 9229 7837 9263 7871
rect 9263 7837 9272 7871
rect 9220 7828 9272 7837
rect 9680 7871 9732 7880
rect 9680 7837 9689 7871
rect 9689 7837 9723 7871
rect 9723 7837 9732 7871
rect 9680 7828 9732 7837
rect 10784 7871 10836 7880
rect 10784 7837 10793 7871
rect 10793 7837 10827 7871
rect 10827 7837 10836 7871
rect 10784 7828 10836 7837
rect 8852 7760 8904 7812
rect 12164 7871 12216 7880
rect 12164 7837 12173 7871
rect 12173 7837 12207 7871
rect 12207 7837 12216 7871
rect 12164 7828 12216 7837
rect 13176 7896 13228 7948
rect 13820 7871 13872 7880
rect 13820 7837 13829 7871
rect 13829 7837 13863 7871
rect 13863 7837 13872 7871
rect 13820 7828 13872 7837
rect 14648 7871 14700 7880
rect 14648 7837 14657 7871
rect 14657 7837 14691 7871
rect 14691 7837 14700 7871
rect 14648 7828 14700 7837
rect 16212 7896 16264 7948
rect 22928 7896 22980 7948
rect 13728 7760 13780 7812
rect 17868 7828 17920 7880
rect 18144 7828 18196 7880
rect 19524 7828 19576 7880
rect 20536 7828 20588 7880
rect 20720 7828 20772 7880
rect 29000 7896 29052 7948
rect 28632 7828 28684 7880
rect 37464 7964 37516 8016
rect 30748 7896 30800 7948
rect 29460 7828 29512 7880
rect 29920 7828 29972 7880
rect 31576 7828 31628 7880
rect 33416 7828 33468 7880
rect 35624 7871 35676 7880
rect 35624 7837 35633 7871
rect 35633 7837 35667 7871
rect 35667 7837 35676 7871
rect 35624 7828 35676 7837
rect 36176 7871 36228 7880
rect 36176 7837 36185 7871
rect 36185 7837 36219 7871
rect 36219 7837 36228 7871
rect 36176 7828 36228 7837
rect 36728 7871 36780 7880
rect 36728 7837 36737 7871
rect 36737 7837 36771 7871
rect 36771 7837 36780 7871
rect 36728 7828 36780 7837
rect 37832 7828 37884 7880
rect 31300 7760 31352 7812
rect 37280 7760 37332 7812
rect 9864 7692 9916 7744
rect 13360 7692 13412 7744
rect 14556 7692 14608 7744
rect 14648 7692 14700 7744
rect 16212 7692 16264 7744
rect 18236 7735 18288 7744
rect 18236 7701 18245 7735
rect 18245 7701 18279 7735
rect 18279 7701 18288 7735
rect 18236 7692 18288 7701
rect 18880 7692 18932 7744
rect 22376 7692 22428 7744
rect 24584 7692 24636 7744
rect 28816 7692 28868 7744
rect 29552 7735 29604 7744
rect 29552 7701 29561 7735
rect 29561 7701 29595 7735
rect 29595 7701 29604 7735
rect 29552 7692 29604 7701
rect 31116 7692 31168 7744
rect 32588 7692 32640 7744
rect 32772 7692 32824 7744
rect 38936 7692 38988 7744
rect 39396 7735 39448 7744
rect 39396 7701 39405 7735
rect 39405 7701 39439 7735
rect 39439 7701 39448 7735
rect 39396 7692 39448 7701
rect 3010 7590 3062 7642
rect 3074 7590 3126 7642
rect 3138 7590 3190 7642
rect 3202 7590 3254 7642
rect 3266 7590 3318 7642
rect 9010 7590 9062 7642
rect 9074 7590 9126 7642
rect 9138 7590 9190 7642
rect 9202 7590 9254 7642
rect 9266 7590 9318 7642
rect 15010 7590 15062 7642
rect 15074 7590 15126 7642
rect 15138 7590 15190 7642
rect 15202 7590 15254 7642
rect 15266 7590 15318 7642
rect 21010 7590 21062 7642
rect 21074 7590 21126 7642
rect 21138 7590 21190 7642
rect 21202 7590 21254 7642
rect 21266 7590 21318 7642
rect 27010 7590 27062 7642
rect 27074 7590 27126 7642
rect 27138 7590 27190 7642
rect 27202 7590 27254 7642
rect 27266 7590 27318 7642
rect 33010 7590 33062 7642
rect 33074 7590 33126 7642
rect 33138 7590 33190 7642
rect 33202 7590 33254 7642
rect 33266 7590 33318 7642
rect 39010 7590 39062 7642
rect 39074 7590 39126 7642
rect 39138 7590 39190 7642
rect 39202 7590 39254 7642
rect 39266 7590 39318 7642
rect 940 7420 992 7472
rect 756 7352 808 7404
rect 2136 7420 2188 7472
rect 3792 7420 3844 7472
rect 940 7284 992 7336
rect 2872 7395 2924 7404
rect 2872 7361 2881 7395
rect 2881 7361 2915 7395
rect 2915 7361 2924 7395
rect 2872 7352 2924 7361
rect 3424 7352 3476 7404
rect 3516 7352 3568 7404
rect 4528 7488 4580 7540
rect 4712 7531 4764 7540
rect 4712 7497 4721 7531
rect 4721 7497 4755 7531
rect 4755 7497 4764 7531
rect 4712 7488 4764 7497
rect 6184 7488 6236 7540
rect 10140 7488 10192 7540
rect 12164 7488 12216 7540
rect 19340 7488 19392 7540
rect 21916 7488 21968 7540
rect 4068 7352 4120 7404
rect 13360 7420 13412 7472
rect 13820 7420 13872 7472
rect 6276 7352 6328 7404
rect 13084 7352 13136 7404
rect 3056 7259 3108 7268
rect 3056 7225 3065 7259
rect 3065 7225 3099 7259
rect 3099 7225 3108 7259
rect 3056 7216 3108 7225
rect 7472 7284 7524 7336
rect 10140 7284 10192 7336
rect 14188 7352 14240 7404
rect 15476 7352 15528 7404
rect 19248 7352 19300 7404
rect 15108 7284 15160 7336
rect 2320 7148 2372 7200
rect 3608 7148 3660 7200
rect 4436 7259 4488 7268
rect 4436 7225 4445 7259
rect 4445 7225 4479 7259
rect 4479 7225 4488 7259
rect 4436 7216 4488 7225
rect 12808 7216 12860 7268
rect 7564 7148 7616 7200
rect 12716 7148 12768 7200
rect 20444 7284 20496 7336
rect 21272 7420 21324 7472
rect 21732 7420 21784 7472
rect 21824 7420 21876 7472
rect 22284 7463 22336 7472
rect 22284 7429 22293 7463
rect 22293 7429 22327 7463
rect 22327 7429 22336 7463
rect 22284 7420 22336 7429
rect 22376 7463 22428 7472
rect 22376 7429 22385 7463
rect 22385 7429 22419 7463
rect 22419 7429 22428 7463
rect 22376 7420 22428 7429
rect 22100 7395 22152 7404
rect 22100 7361 22109 7395
rect 22109 7361 22143 7395
rect 22143 7361 22152 7395
rect 22100 7352 22152 7361
rect 30840 7488 30892 7540
rect 25504 7420 25556 7472
rect 29552 7420 29604 7472
rect 30288 7420 30340 7472
rect 21364 7284 21416 7336
rect 22008 7284 22060 7336
rect 23020 7395 23072 7404
rect 23020 7361 23029 7395
rect 23029 7361 23063 7395
rect 23063 7361 23072 7395
rect 23020 7352 23072 7361
rect 24124 7352 24176 7404
rect 27252 7352 27304 7404
rect 30012 7352 30064 7404
rect 22744 7284 22796 7336
rect 28816 7284 28868 7336
rect 30564 7284 30616 7336
rect 36176 7488 36228 7540
rect 36268 7488 36320 7540
rect 35900 7420 35952 7472
rect 32588 7395 32640 7404
rect 32588 7361 32597 7395
rect 32597 7361 32631 7395
rect 32631 7361 32640 7395
rect 32588 7352 32640 7361
rect 31668 7284 31720 7336
rect 14464 7148 14516 7200
rect 15384 7148 15436 7200
rect 15568 7148 15620 7200
rect 15844 7148 15896 7200
rect 17776 7148 17828 7200
rect 19248 7148 19300 7200
rect 24768 7148 24820 7200
rect 30472 7148 30524 7200
rect 31300 7191 31352 7200
rect 31300 7157 31309 7191
rect 31309 7157 31343 7191
rect 31343 7157 31352 7191
rect 31300 7148 31352 7157
rect 31576 7191 31628 7200
rect 31576 7157 31585 7191
rect 31585 7157 31619 7191
rect 31619 7157 31628 7191
rect 31576 7148 31628 7157
rect 32128 7191 32180 7200
rect 32128 7157 32137 7191
rect 32137 7157 32171 7191
rect 32171 7157 32180 7191
rect 32128 7148 32180 7157
rect 32404 7191 32456 7200
rect 32404 7157 32413 7191
rect 32413 7157 32447 7191
rect 32447 7157 32456 7191
rect 32404 7148 32456 7157
rect 32588 7148 32640 7200
rect 34244 7395 34296 7404
rect 34244 7361 34253 7395
rect 34253 7361 34287 7395
rect 34287 7361 34296 7395
rect 34244 7352 34296 7361
rect 37372 7395 37424 7404
rect 37372 7361 37381 7395
rect 37381 7361 37415 7395
rect 37415 7361 37424 7395
rect 37372 7352 37424 7361
rect 37556 7352 37608 7404
rect 38292 7531 38344 7540
rect 38292 7497 38301 7531
rect 38301 7497 38335 7531
rect 38335 7497 38344 7531
rect 38292 7488 38344 7497
rect 38752 7488 38804 7540
rect 39488 7488 39540 7540
rect 39856 7420 39908 7472
rect 38844 7395 38896 7404
rect 38844 7361 38853 7395
rect 38853 7361 38887 7395
rect 38887 7361 38896 7395
rect 38844 7352 38896 7361
rect 39028 7352 39080 7404
rect 36544 7216 36596 7268
rect 38936 7284 38988 7336
rect 39488 7216 39540 7268
rect 35992 7148 36044 7200
rect 38844 7148 38896 7200
rect 1950 7046 2002 7098
rect 2014 7046 2066 7098
rect 2078 7046 2130 7098
rect 2142 7046 2194 7098
rect 2206 7046 2258 7098
rect 7950 7046 8002 7098
rect 8014 7046 8066 7098
rect 8078 7046 8130 7098
rect 8142 7046 8194 7098
rect 8206 7046 8258 7098
rect 13950 7046 14002 7098
rect 14014 7046 14066 7098
rect 14078 7046 14130 7098
rect 14142 7046 14194 7098
rect 14206 7046 14258 7098
rect 19950 7046 20002 7098
rect 20014 7046 20066 7098
rect 20078 7046 20130 7098
rect 20142 7046 20194 7098
rect 20206 7046 20258 7098
rect 25950 7046 26002 7098
rect 26014 7046 26066 7098
rect 26078 7046 26130 7098
rect 26142 7046 26194 7098
rect 26206 7046 26258 7098
rect 31950 7046 32002 7098
rect 32014 7046 32066 7098
rect 32078 7046 32130 7098
rect 32142 7046 32194 7098
rect 32206 7046 32258 7098
rect 37950 7046 38002 7098
rect 38014 7046 38066 7098
rect 38078 7046 38130 7098
rect 38142 7046 38194 7098
rect 38206 7046 38258 7098
rect 3792 6944 3844 6996
rect 9680 6944 9732 6996
rect 9864 6987 9916 6996
rect 9864 6953 9873 6987
rect 9873 6953 9907 6987
rect 9907 6953 9916 6987
rect 9864 6944 9916 6953
rect 13728 6987 13780 6996
rect 13728 6953 13737 6987
rect 13737 6953 13771 6987
rect 13771 6953 13780 6987
rect 13728 6944 13780 6953
rect 12256 6876 12308 6928
rect 18236 6944 18288 6996
rect 18328 6944 18380 6996
rect 20628 6944 20680 6996
rect 22008 6944 22060 6996
rect 22468 6944 22520 6996
rect 23020 6944 23072 6996
rect 16488 6919 16540 6928
rect 16488 6885 16497 6919
rect 16497 6885 16531 6919
rect 16531 6885 16540 6919
rect 16488 6876 16540 6885
rect 9772 6808 9824 6860
rect 15108 6851 15160 6860
rect 15108 6817 15117 6851
rect 15117 6817 15151 6851
rect 15151 6817 15160 6851
rect 15108 6808 15160 6817
rect 16304 6808 16356 6860
rect 22560 6876 22612 6928
rect 27344 6944 27396 6996
rect 23664 6808 23716 6860
rect 24492 6808 24544 6860
rect 2780 6672 2832 6724
rect 3516 6672 3568 6724
rect 8576 6740 8628 6792
rect 7840 6672 7892 6724
rect 8760 6672 8812 6724
rect 9864 6740 9916 6792
rect 10324 6740 10376 6792
rect 11428 6740 11480 6792
rect 12256 6740 12308 6792
rect 12992 6740 13044 6792
rect 13820 6740 13872 6792
rect 9404 6715 9456 6724
rect 9404 6681 9413 6715
rect 9413 6681 9447 6715
rect 9447 6681 9456 6715
rect 9404 6672 9456 6681
rect 3700 6604 3752 6656
rect 3976 6647 4028 6656
rect 3976 6613 3985 6647
rect 3985 6613 4019 6647
rect 4019 6613 4028 6647
rect 3976 6604 4028 6613
rect 12164 6672 12216 6724
rect 15384 6740 15436 6792
rect 15844 6740 15896 6792
rect 15108 6672 15160 6724
rect 20168 6740 20220 6792
rect 17684 6672 17736 6724
rect 20536 6783 20588 6792
rect 20536 6749 20545 6783
rect 20545 6749 20579 6783
rect 20579 6749 20588 6783
rect 20536 6740 20588 6749
rect 20444 6672 20496 6724
rect 21732 6740 21784 6792
rect 23112 6740 23164 6792
rect 22652 6672 22704 6724
rect 9588 6604 9640 6656
rect 10048 6604 10100 6656
rect 11612 6604 11664 6656
rect 13820 6604 13872 6656
rect 14188 6604 14240 6656
rect 15476 6604 15528 6656
rect 16028 6604 16080 6656
rect 16212 6604 16264 6656
rect 19340 6604 19392 6656
rect 20904 6604 20956 6656
rect 21456 6604 21508 6656
rect 22468 6647 22520 6656
rect 22468 6613 22477 6647
rect 22477 6613 22511 6647
rect 22511 6613 22520 6647
rect 22468 6604 22520 6613
rect 22836 6604 22888 6656
rect 25596 6876 25648 6928
rect 26424 6808 26476 6860
rect 23572 6672 23624 6724
rect 27712 6919 27764 6928
rect 27712 6885 27721 6919
rect 27721 6885 27755 6919
rect 27755 6885 27764 6919
rect 27712 6876 27764 6885
rect 30380 6944 30432 6996
rect 37556 6944 37608 6996
rect 29000 6876 29052 6928
rect 37648 6876 37700 6928
rect 27896 6783 27948 6792
rect 27896 6749 27905 6783
rect 27905 6749 27939 6783
rect 27939 6749 27948 6783
rect 27896 6740 27948 6749
rect 28172 6783 28224 6792
rect 28172 6749 28181 6783
rect 28181 6749 28215 6783
rect 28215 6749 28224 6783
rect 28172 6740 28224 6749
rect 28448 6783 28500 6792
rect 28448 6749 28457 6783
rect 28457 6749 28491 6783
rect 28491 6749 28500 6783
rect 28448 6740 28500 6749
rect 29000 6783 29052 6792
rect 29000 6749 29009 6783
rect 29009 6749 29043 6783
rect 29043 6749 29052 6783
rect 29000 6740 29052 6749
rect 31852 6808 31904 6860
rect 29736 6783 29788 6792
rect 29736 6749 29745 6783
rect 29745 6749 29779 6783
rect 29779 6749 29788 6783
rect 29736 6740 29788 6749
rect 30012 6783 30064 6792
rect 30012 6749 30021 6783
rect 30021 6749 30055 6783
rect 30055 6749 30064 6783
rect 30012 6740 30064 6749
rect 31392 6740 31444 6792
rect 37096 6808 37148 6860
rect 38292 6808 38344 6860
rect 39028 6808 39080 6860
rect 32404 6783 32456 6792
rect 32404 6749 32413 6783
rect 32413 6749 32447 6783
rect 32447 6749 32456 6783
rect 32404 6740 32456 6749
rect 29184 6672 29236 6724
rect 38476 6783 38528 6792
rect 38476 6749 38485 6783
rect 38485 6749 38519 6783
rect 38519 6749 38528 6783
rect 38476 6740 38528 6749
rect 38752 6740 38804 6792
rect 24676 6647 24728 6656
rect 24676 6613 24685 6647
rect 24685 6613 24719 6647
rect 24719 6613 24728 6647
rect 24676 6604 24728 6613
rect 25136 6647 25188 6656
rect 25136 6613 25145 6647
rect 25145 6613 25179 6647
rect 25179 6613 25188 6647
rect 25136 6604 25188 6613
rect 26792 6604 26844 6656
rect 27252 6604 27304 6656
rect 27988 6647 28040 6656
rect 27988 6613 27997 6647
rect 27997 6613 28031 6647
rect 28031 6613 28040 6647
rect 27988 6604 28040 6613
rect 28264 6647 28316 6656
rect 28264 6613 28273 6647
rect 28273 6613 28307 6647
rect 28307 6613 28316 6647
rect 28264 6604 28316 6613
rect 28540 6647 28592 6656
rect 28540 6613 28549 6647
rect 28549 6613 28583 6647
rect 28583 6613 28592 6647
rect 28540 6604 28592 6613
rect 28724 6604 28776 6656
rect 28908 6604 28960 6656
rect 29368 6604 29420 6656
rect 29828 6647 29880 6656
rect 29828 6613 29837 6647
rect 29837 6613 29871 6647
rect 29871 6613 29880 6647
rect 29828 6604 29880 6613
rect 31484 6604 31536 6656
rect 31852 6604 31904 6656
rect 35624 6672 35676 6724
rect 34704 6604 34756 6656
rect 38568 6604 38620 6656
rect 38660 6647 38712 6656
rect 38660 6613 38669 6647
rect 38669 6613 38703 6647
rect 38703 6613 38712 6647
rect 38660 6604 38712 6613
rect 38844 6604 38896 6656
rect 39580 6672 39632 6724
rect 39396 6647 39448 6656
rect 39396 6613 39405 6647
rect 39405 6613 39439 6647
rect 39439 6613 39448 6647
rect 39396 6604 39448 6613
rect 3010 6502 3062 6554
rect 3074 6502 3126 6554
rect 3138 6502 3190 6554
rect 3202 6502 3254 6554
rect 3266 6502 3318 6554
rect 9010 6502 9062 6554
rect 9074 6502 9126 6554
rect 9138 6502 9190 6554
rect 9202 6502 9254 6554
rect 9266 6502 9318 6554
rect 15010 6502 15062 6554
rect 15074 6502 15126 6554
rect 15138 6502 15190 6554
rect 15202 6502 15254 6554
rect 15266 6502 15318 6554
rect 21010 6502 21062 6554
rect 21074 6502 21126 6554
rect 21138 6502 21190 6554
rect 21202 6502 21254 6554
rect 21266 6502 21318 6554
rect 27010 6502 27062 6554
rect 27074 6502 27126 6554
rect 27138 6502 27190 6554
rect 27202 6502 27254 6554
rect 27266 6502 27318 6554
rect 33010 6502 33062 6554
rect 33074 6502 33126 6554
rect 33138 6502 33190 6554
rect 33202 6502 33254 6554
rect 33266 6502 33318 6554
rect 39010 6502 39062 6554
rect 39074 6502 39126 6554
rect 39138 6502 39190 6554
rect 39202 6502 39254 6554
rect 39266 6502 39318 6554
rect 8300 6400 8352 6452
rect 8668 6400 8720 6452
rect 8944 6400 8996 6452
rect 9128 6400 9180 6452
rect 11888 6400 11940 6452
rect 11980 6400 12032 6452
rect 13268 6400 13320 6452
rect 14648 6332 14700 6384
rect 15384 6332 15436 6384
rect 15752 6400 15804 6452
rect 8668 6264 8720 6316
rect 8944 6264 8996 6316
rect 3884 6196 3936 6248
rect 9220 6196 9272 6248
rect 9496 6196 9548 6248
rect 10048 6307 10100 6316
rect 10048 6273 10057 6307
rect 10057 6273 10091 6307
rect 10091 6273 10100 6307
rect 10048 6264 10100 6273
rect 11520 6264 11572 6316
rect 12532 6264 12584 6316
rect 12164 6196 12216 6248
rect 14096 6264 14148 6316
rect 14556 6307 14608 6316
rect 14556 6273 14566 6307
rect 14566 6273 14600 6307
rect 14600 6273 14608 6307
rect 14556 6264 14608 6273
rect 14740 6307 14792 6316
rect 14740 6273 14749 6307
rect 14749 6273 14783 6307
rect 14783 6273 14792 6307
rect 14740 6264 14792 6273
rect 16028 6264 16080 6316
rect 16212 6264 16264 6316
rect 14188 6196 14240 6248
rect 14280 6196 14332 6248
rect 17684 6307 17736 6316
rect 17684 6273 17693 6307
rect 17693 6273 17727 6307
rect 17727 6273 17736 6307
rect 17684 6264 17736 6273
rect 17960 6307 18012 6316
rect 17960 6273 17969 6307
rect 17969 6273 18003 6307
rect 18003 6273 18012 6307
rect 17960 6264 18012 6273
rect 19248 6264 19300 6316
rect 19616 6264 19668 6316
rect 20996 6400 21048 6452
rect 22100 6400 22152 6452
rect 38476 6400 38528 6452
rect 40040 6400 40092 6452
rect 20444 6264 20496 6316
rect 21916 6307 21968 6316
rect 21916 6273 21926 6307
rect 21926 6273 21960 6307
rect 21960 6273 21968 6307
rect 21916 6264 21968 6273
rect 22100 6307 22152 6316
rect 22100 6273 22109 6307
rect 22109 6273 22143 6307
rect 22143 6273 22152 6307
rect 22100 6264 22152 6273
rect 22192 6307 22244 6316
rect 22192 6273 22201 6307
rect 22201 6273 22235 6307
rect 22235 6273 22244 6307
rect 22192 6264 22244 6273
rect 23848 6332 23900 6384
rect 26700 6332 26752 6384
rect 29000 6332 29052 6384
rect 31852 6332 31904 6384
rect 38752 6332 38804 6384
rect 19432 6239 19484 6248
rect 19432 6205 19441 6239
rect 19441 6205 19475 6239
rect 19475 6205 19484 6239
rect 19432 6196 19484 6205
rect 5540 6128 5592 6180
rect 7748 6060 7800 6112
rect 10048 6060 10100 6112
rect 15844 6128 15896 6180
rect 18972 6128 19024 6180
rect 12532 6060 12584 6112
rect 13728 6060 13780 6112
rect 14648 6060 14700 6112
rect 16396 6060 16448 6112
rect 17684 6060 17736 6112
rect 17868 6060 17920 6112
rect 20536 6196 20588 6248
rect 22652 6196 22704 6248
rect 23756 6264 23808 6316
rect 26516 6264 26568 6316
rect 27436 6264 27488 6316
rect 29736 6264 29788 6316
rect 31392 6264 31444 6316
rect 37464 6264 37516 6316
rect 23112 6239 23164 6248
rect 23112 6205 23121 6239
rect 23121 6205 23155 6239
rect 23155 6205 23164 6239
rect 23112 6196 23164 6205
rect 23940 6196 23992 6248
rect 24768 6196 24820 6248
rect 27528 6196 27580 6248
rect 30012 6196 30064 6248
rect 35256 6196 35308 6248
rect 39212 6307 39264 6316
rect 39212 6273 39221 6307
rect 39221 6273 39255 6307
rect 39255 6273 39264 6307
rect 39212 6264 39264 6273
rect 28172 6128 28224 6180
rect 35808 6128 35860 6180
rect 20536 6103 20588 6112
rect 20536 6069 20545 6103
rect 20545 6069 20579 6103
rect 20579 6069 20588 6103
rect 20536 6060 20588 6069
rect 22284 6060 22336 6112
rect 23020 6103 23072 6112
rect 23020 6069 23029 6103
rect 23029 6069 23063 6103
rect 23063 6069 23072 6103
rect 23020 6060 23072 6069
rect 23480 6060 23532 6112
rect 24676 6060 24728 6112
rect 30380 6060 30432 6112
rect 37280 6060 37332 6112
rect 38660 6060 38712 6112
rect 39028 6103 39080 6112
rect 39028 6069 39037 6103
rect 39037 6069 39071 6103
rect 39071 6069 39080 6103
rect 39028 6060 39080 6069
rect 1950 5958 2002 6010
rect 2014 5958 2066 6010
rect 2078 5958 2130 6010
rect 2142 5958 2194 6010
rect 2206 5958 2258 6010
rect 7950 5958 8002 6010
rect 8014 5958 8066 6010
rect 8078 5958 8130 6010
rect 8142 5958 8194 6010
rect 8206 5958 8258 6010
rect 13950 5958 14002 6010
rect 14014 5958 14066 6010
rect 14078 5958 14130 6010
rect 14142 5958 14194 6010
rect 14206 5958 14258 6010
rect 19950 5958 20002 6010
rect 20014 5958 20066 6010
rect 20078 5958 20130 6010
rect 20142 5958 20194 6010
rect 20206 5958 20258 6010
rect 25950 5958 26002 6010
rect 26014 5958 26066 6010
rect 26078 5958 26130 6010
rect 26142 5958 26194 6010
rect 26206 5958 26258 6010
rect 31950 5958 32002 6010
rect 32014 5958 32066 6010
rect 32078 5958 32130 6010
rect 32142 5958 32194 6010
rect 32206 5958 32258 6010
rect 37950 5958 38002 6010
rect 38014 5958 38066 6010
rect 38078 5958 38130 6010
rect 38142 5958 38194 6010
rect 38206 5958 38258 6010
rect 7380 5856 7432 5908
rect 8484 5856 8536 5908
rect 8852 5856 8904 5908
rect 6920 5788 6972 5840
rect 7472 5788 7524 5840
rect 14096 5856 14148 5908
rect 9220 5788 9272 5840
rect 13268 5788 13320 5840
rect 13360 5831 13412 5840
rect 13360 5797 13369 5831
rect 13369 5797 13403 5831
rect 13403 5797 13412 5831
rect 13360 5788 13412 5797
rect 14372 5856 14424 5908
rect 14832 5899 14884 5908
rect 14832 5865 14841 5899
rect 14841 5865 14875 5899
rect 14875 5865 14884 5899
rect 14832 5856 14884 5865
rect 15660 5856 15712 5908
rect 17408 5856 17460 5908
rect 17500 5856 17552 5908
rect 17684 5856 17736 5908
rect 18512 5899 18564 5908
rect 18512 5865 18521 5899
rect 18521 5865 18555 5899
rect 18555 5865 18564 5899
rect 18512 5856 18564 5865
rect 19616 5856 19668 5908
rect 20352 5856 20404 5908
rect 20628 5856 20680 5908
rect 21180 5856 21232 5908
rect 21456 5856 21508 5908
rect 21548 5856 21600 5908
rect 24308 5856 24360 5908
rect 35256 5856 35308 5908
rect 36728 5856 36780 5908
rect 36912 5899 36964 5908
rect 36912 5865 36921 5899
rect 36921 5865 36955 5899
rect 36955 5865 36964 5899
rect 36912 5856 36964 5865
rect 37648 5856 37700 5908
rect 39580 5856 39632 5908
rect 17132 5831 17184 5840
rect 17132 5797 17141 5831
rect 17141 5797 17175 5831
rect 17175 5797 17184 5831
rect 17132 5788 17184 5797
rect 10324 5763 10376 5772
rect 10324 5729 10333 5763
rect 10333 5729 10367 5763
rect 10367 5729 10376 5763
rect 10324 5720 10376 5729
rect 12808 5720 12860 5772
rect 6644 5652 6696 5704
rect 7104 5652 7156 5704
rect 7656 5652 7708 5704
rect 8576 5652 8628 5704
rect 9128 5695 9180 5704
rect 9128 5661 9137 5695
rect 9137 5661 9171 5695
rect 9171 5661 9180 5695
rect 9128 5652 9180 5661
rect 9680 5652 9732 5704
rect 10048 5652 10100 5704
rect 10140 5695 10192 5704
rect 10140 5661 10149 5695
rect 10149 5661 10183 5695
rect 10183 5661 10192 5695
rect 10140 5652 10192 5661
rect 13084 5652 13136 5704
rect 13268 5652 13320 5704
rect 13728 5720 13780 5772
rect 14372 5695 14424 5704
rect 14372 5661 14381 5695
rect 14381 5661 14415 5695
rect 14415 5661 14424 5695
rect 14372 5652 14424 5661
rect 2872 5584 2924 5636
rect 6920 5584 6972 5636
rect 9956 5627 10008 5636
rect 9956 5593 9965 5627
rect 9965 5593 9999 5627
rect 9999 5593 10008 5627
rect 9956 5584 10008 5593
rect 13728 5584 13780 5636
rect 14648 5695 14700 5704
rect 14648 5661 14657 5695
rect 14657 5661 14691 5695
rect 14691 5661 14700 5695
rect 14648 5652 14700 5661
rect 15660 5652 15712 5704
rect 16672 5652 16724 5704
rect 16764 5652 16816 5704
rect 21732 5788 21784 5840
rect 19800 5720 19852 5772
rect 17592 5652 17644 5704
rect 18696 5695 18748 5704
rect 18696 5661 18705 5695
rect 18705 5661 18739 5695
rect 18739 5661 18748 5695
rect 18696 5652 18748 5661
rect 19708 5652 19760 5704
rect 20352 5695 20404 5704
rect 20352 5661 20361 5695
rect 20361 5661 20395 5695
rect 20395 5661 20404 5695
rect 20352 5652 20404 5661
rect 20904 5720 20956 5772
rect 31852 5788 31904 5840
rect 34060 5788 34112 5840
rect 22008 5652 22060 5704
rect 24216 5695 24268 5704
rect 24216 5661 24225 5695
rect 24225 5661 24259 5695
rect 24259 5661 24268 5695
rect 24216 5652 24268 5661
rect 24584 5695 24636 5704
rect 24584 5661 24593 5695
rect 24593 5661 24627 5695
rect 24627 5661 24636 5695
rect 24584 5652 24636 5661
rect 24860 5695 24912 5704
rect 24860 5661 24869 5695
rect 24869 5661 24903 5695
rect 24903 5661 24912 5695
rect 24860 5652 24912 5661
rect 25688 5652 25740 5704
rect 26700 5720 26752 5772
rect 32404 5720 32456 5772
rect 26884 5652 26936 5704
rect 32772 5652 32824 5704
rect 23480 5584 23532 5636
rect 34612 5584 34664 5636
rect 38568 5652 38620 5704
rect 38936 5652 38988 5704
rect 14924 5516 14976 5568
rect 19432 5516 19484 5568
rect 21180 5516 21232 5568
rect 21456 5559 21508 5568
rect 21456 5525 21465 5559
rect 21465 5525 21499 5559
rect 21499 5525 21508 5559
rect 21456 5516 21508 5525
rect 21548 5516 21600 5568
rect 24308 5516 24360 5568
rect 24400 5559 24452 5568
rect 24400 5525 24409 5559
rect 24409 5525 24443 5559
rect 24443 5525 24452 5559
rect 24400 5516 24452 5525
rect 24676 5559 24728 5568
rect 24676 5525 24685 5559
rect 24685 5525 24719 5559
rect 24719 5525 24728 5559
rect 24676 5516 24728 5525
rect 31668 5516 31720 5568
rect 38752 5516 38804 5568
rect 39304 5516 39356 5568
rect 3010 5414 3062 5466
rect 3074 5414 3126 5466
rect 3138 5414 3190 5466
rect 3202 5414 3254 5466
rect 3266 5414 3318 5466
rect 9010 5414 9062 5466
rect 9074 5414 9126 5466
rect 9138 5414 9190 5466
rect 9202 5414 9254 5466
rect 9266 5414 9318 5466
rect 15010 5414 15062 5466
rect 15074 5414 15126 5466
rect 15138 5414 15190 5466
rect 15202 5414 15254 5466
rect 15266 5414 15318 5466
rect 21010 5414 21062 5466
rect 21074 5414 21126 5466
rect 21138 5414 21190 5466
rect 21202 5414 21254 5466
rect 21266 5414 21318 5466
rect 27010 5414 27062 5466
rect 27074 5414 27126 5466
rect 27138 5414 27190 5466
rect 27202 5414 27254 5466
rect 27266 5414 27318 5466
rect 33010 5414 33062 5466
rect 33074 5414 33126 5466
rect 33138 5414 33190 5466
rect 33202 5414 33254 5466
rect 33266 5414 33318 5466
rect 39010 5414 39062 5466
rect 39074 5414 39126 5466
rect 39138 5414 39190 5466
rect 39202 5414 39254 5466
rect 39266 5414 39318 5466
rect 7564 5312 7616 5364
rect 15292 5312 15344 5364
rect 8852 5244 8904 5296
rect 13268 5244 13320 5296
rect 15752 5244 15804 5296
rect 664 5176 716 5228
rect 3424 5176 3476 5228
rect 14280 5176 14332 5228
rect 15292 5219 15344 5228
rect 15292 5185 15301 5219
rect 15301 5185 15335 5219
rect 15335 5185 15344 5219
rect 17868 5244 17920 5296
rect 15292 5176 15344 5185
rect 17040 5219 17092 5228
rect 17040 5185 17049 5219
rect 17049 5185 17083 5219
rect 17083 5185 17092 5219
rect 17040 5176 17092 5185
rect 17684 5219 17736 5228
rect 17684 5185 17693 5219
rect 17693 5185 17727 5219
rect 17727 5185 17736 5219
rect 17684 5176 17736 5185
rect 19708 5176 19760 5228
rect 20352 5244 20404 5296
rect 32496 5312 32548 5364
rect 37740 5312 37792 5364
rect 38384 5312 38436 5364
rect 38844 5312 38896 5364
rect 39488 5312 39540 5364
rect 22744 5176 22796 5228
rect 9588 5151 9640 5160
rect 9588 5117 9597 5151
rect 9597 5117 9631 5151
rect 9631 5117 9640 5151
rect 9588 5108 9640 5117
rect 13360 5108 13412 5160
rect 4068 5040 4120 5092
rect 12256 5040 12308 5092
rect 15568 5040 15620 5092
rect 16120 5040 16172 5092
rect 3976 4972 4028 5024
rect 15292 4972 15344 5024
rect 16580 4972 16632 5024
rect 19248 5108 19300 5160
rect 25872 5176 25924 5228
rect 26884 5176 26936 5228
rect 31576 5176 31628 5228
rect 36084 5176 36136 5228
rect 37648 5176 37700 5228
rect 38844 5219 38896 5228
rect 38844 5185 38853 5219
rect 38853 5185 38887 5219
rect 38887 5185 38896 5219
rect 38844 5176 38896 5185
rect 39212 5219 39264 5228
rect 39212 5185 39221 5219
rect 39221 5185 39255 5219
rect 39255 5185 39264 5219
rect 39212 5176 39264 5185
rect 36268 5108 36320 5160
rect 26608 5083 26660 5092
rect 26608 5049 26617 5083
rect 26617 5049 26651 5083
rect 26651 5049 26660 5083
rect 26608 5040 26660 5049
rect 35992 5040 36044 5092
rect 20352 4972 20404 5024
rect 21916 4972 21968 5024
rect 22652 4972 22704 5024
rect 39028 5015 39080 5024
rect 39028 4981 39037 5015
rect 39037 4981 39071 5015
rect 39071 4981 39080 5015
rect 39028 4972 39080 4981
rect 1950 4870 2002 4922
rect 2014 4870 2066 4922
rect 2078 4870 2130 4922
rect 2142 4870 2194 4922
rect 2206 4870 2258 4922
rect 7950 4870 8002 4922
rect 8014 4870 8066 4922
rect 8078 4870 8130 4922
rect 8142 4870 8194 4922
rect 8206 4870 8258 4922
rect 13950 4870 14002 4922
rect 14014 4870 14066 4922
rect 14078 4870 14130 4922
rect 14142 4870 14194 4922
rect 14206 4870 14258 4922
rect 19950 4870 20002 4922
rect 20014 4870 20066 4922
rect 20078 4870 20130 4922
rect 20142 4870 20194 4922
rect 20206 4870 20258 4922
rect 25950 4870 26002 4922
rect 26014 4870 26066 4922
rect 26078 4870 26130 4922
rect 26142 4870 26194 4922
rect 26206 4870 26258 4922
rect 31950 4870 32002 4922
rect 32014 4870 32066 4922
rect 32078 4870 32130 4922
rect 32142 4870 32194 4922
rect 32206 4870 32258 4922
rect 37950 4870 38002 4922
rect 38014 4870 38066 4922
rect 38078 4870 38130 4922
rect 38142 4870 38194 4922
rect 38206 4870 38258 4922
rect 9864 4768 9916 4820
rect 12256 4811 12308 4820
rect 12256 4777 12265 4811
rect 12265 4777 12299 4811
rect 12299 4777 12308 4811
rect 12256 4768 12308 4777
rect 13360 4811 13412 4820
rect 13360 4777 13369 4811
rect 13369 4777 13403 4811
rect 13403 4777 13412 4811
rect 13360 4768 13412 4777
rect 13544 4811 13596 4820
rect 13544 4777 13553 4811
rect 13553 4777 13587 4811
rect 13587 4777 13596 4811
rect 13544 4768 13596 4777
rect 14280 4811 14332 4820
rect 14280 4777 14289 4811
rect 14289 4777 14323 4811
rect 14323 4777 14332 4811
rect 14280 4768 14332 4777
rect 16028 4768 16080 4820
rect 17040 4768 17092 4820
rect 21640 4768 21692 4820
rect 21732 4811 21784 4820
rect 21732 4777 21741 4811
rect 21741 4777 21775 4811
rect 21775 4777 21784 4811
rect 21732 4768 21784 4777
rect 32864 4768 32916 4820
rect 37832 4768 37884 4820
rect 39396 4811 39448 4820
rect 39396 4777 39405 4811
rect 39405 4777 39439 4811
rect 39439 4777 39448 4811
rect 39396 4768 39448 4777
rect 3516 4700 3568 4752
rect 38844 4700 38896 4752
rect 3884 4632 3936 4684
rect 7288 4564 7340 4616
rect 2780 4496 2832 4548
rect 7564 4564 7616 4616
rect 8760 4564 8812 4616
rect 12716 4632 12768 4684
rect 11428 4607 11480 4616
rect 11428 4573 11437 4607
rect 11437 4573 11471 4607
rect 11471 4573 11480 4607
rect 11428 4564 11480 4573
rect 11612 4564 11664 4616
rect 12072 4607 12124 4616
rect 12072 4573 12081 4607
rect 12081 4573 12115 4607
rect 12115 4573 12124 4607
rect 12072 4564 12124 4573
rect 12164 4564 12216 4616
rect 13820 4632 13872 4684
rect 15292 4632 15344 4684
rect 38292 4632 38344 4684
rect 38660 4632 38712 4684
rect 13728 4607 13780 4616
rect 13728 4573 13737 4607
rect 13737 4573 13771 4607
rect 13771 4573 13780 4607
rect 13728 4564 13780 4573
rect 14464 4564 14516 4616
rect 14556 4564 14608 4616
rect 16396 4607 16448 4616
rect 16396 4573 16405 4607
rect 16405 4573 16439 4607
rect 16439 4573 16448 4607
rect 16396 4564 16448 4573
rect 16672 4607 16724 4616
rect 16672 4573 16681 4607
rect 16681 4573 16715 4607
rect 16715 4573 16724 4607
rect 16672 4564 16724 4573
rect 17592 4564 17644 4616
rect 20720 4564 20772 4616
rect 12164 4428 12216 4480
rect 13176 4496 13228 4548
rect 12532 4428 12584 4480
rect 14280 4496 14332 4548
rect 30380 4496 30432 4548
rect 38936 4564 38988 4616
rect 39580 4496 39632 4548
rect 18328 4428 18380 4480
rect 19708 4428 19760 4480
rect 22468 4428 22520 4480
rect 25044 4428 25096 4480
rect 31300 4428 31352 4480
rect 33508 4428 33560 4480
rect 39304 4428 39356 4480
rect 3010 4326 3062 4378
rect 3074 4326 3126 4378
rect 3138 4326 3190 4378
rect 3202 4326 3254 4378
rect 3266 4326 3318 4378
rect 9010 4326 9062 4378
rect 9074 4326 9126 4378
rect 9138 4326 9190 4378
rect 9202 4326 9254 4378
rect 9266 4326 9318 4378
rect 15010 4326 15062 4378
rect 15074 4326 15126 4378
rect 15138 4326 15190 4378
rect 15202 4326 15254 4378
rect 15266 4326 15318 4378
rect 21010 4326 21062 4378
rect 21074 4326 21126 4378
rect 21138 4326 21190 4378
rect 21202 4326 21254 4378
rect 21266 4326 21318 4378
rect 27010 4326 27062 4378
rect 27074 4326 27126 4378
rect 27138 4326 27190 4378
rect 27202 4326 27254 4378
rect 27266 4326 27318 4378
rect 33010 4326 33062 4378
rect 33074 4326 33126 4378
rect 33138 4326 33190 4378
rect 33202 4326 33254 4378
rect 33266 4326 33318 4378
rect 39010 4326 39062 4378
rect 39074 4326 39126 4378
rect 39138 4326 39190 4378
rect 39202 4326 39254 4378
rect 39266 4326 39318 4378
rect 1216 4224 1268 4276
rect 1308 4156 1360 4208
rect 7288 4224 7340 4276
rect 3608 4199 3660 4208
rect 3608 4165 3617 4199
rect 3617 4165 3651 4199
rect 3651 4165 3660 4199
rect 3608 4156 3660 4165
rect 8668 4267 8720 4276
rect 8668 4233 8677 4267
rect 8677 4233 8711 4267
rect 8711 4233 8720 4267
rect 8668 4224 8720 4233
rect 18052 4224 18104 4276
rect 19524 4224 19576 4276
rect 21824 4224 21876 4276
rect 23848 4267 23900 4276
rect 23848 4233 23857 4267
rect 23857 4233 23891 4267
rect 23891 4233 23900 4267
rect 23848 4224 23900 4233
rect 23756 4156 23808 4208
rect 28264 4156 28316 4208
rect 32588 4156 32640 4208
rect 2872 4131 2924 4140
rect 2872 4097 2881 4131
rect 2881 4097 2915 4131
rect 2915 4097 2924 4131
rect 2872 4088 2924 4097
rect 4712 4020 4764 4072
rect 6644 4020 6696 4072
rect 7288 4131 7340 4140
rect 7288 4097 7297 4131
rect 7297 4097 7331 4131
rect 7331 4097 7340 4131
rect 7288 4088 7340 4097
rect 7380 4131 7432 4140
rect 7380 4097 7414 4131
rect 7414 4097 7432 4131
rect 7380 4088 7432 4097
rect 7564 4131 7616 4140
rect 7564 4097 7573 4131
rect 7573 4097 7607 4131
rect 7607 4097 7616 4131
rect 7564 4088 7616 4097
rect 8576 4131 8628 4140
rect 8576 4097 8585 4131
rect 8585 4097 8619 4131
rect 8619 4097 8628 4131
rect 8576 4088 8628 4097
rect 9588 4088 9640 4140
rect 7104 4020 7156 4072
rect 7748 4020 7800 4072
rect 10232 4131 10284 4140
rect 10232 4097 10241 4131
rect 10241 4097 10275 4131
rect 10275 4097 10284 4131
rect 10232 4088 10284 4097
rect 11336 4088 11388 4140
rect 14556 4088 14608 4140
rect 15568 4088 15620 4140
rect 3056 3995 3108 4004
rect 3056 3961 3065 3995
rect 3065 3961 3099 3995
rect 3099 3961 3108 3995
rect 3056 3952 3108 3961
rect 3792 3995 3844 4004
rect 3792 3961 3801 3995
rect 3801 3961 3835 3995
rect 3835 3961 3844 3995
rect 3792 3952 3844 3961
rect 12716 4020 12768 4072
rect 3516 3884 3568 3936
rect 9404 3952 9456 4004
rect 14740 3952 14792 4004
rect 15476 4063 15528 4072
rect 15476 4029 15485 4063
rect 15485 4029 15519 4063
rect 15519 4029 15528 4063
rect 15476 4020 15528 4029
rect 16672 4020 16724 4072
rect 18052 4131 18104 4140
rect 18052 4097 18059 4131
rect 18059 4097 18104 4131
rect 18052 4088 18104 4097
rect 18144 4131 18196 4140
rect 18144 4097 18153 4131
rect 18153 4097 18187 4131
rect 18187 4097 18196 4131
rect 18144 4088 18196 4097
rect 18880 4088 18932 4140
rect 20260 4131 20312 4140
rect 20260 4097 20269 4131
rect 20269 4097 20303 4131
rect 20303 4097 20312 4131
rect 20260 4088 20312 4097
rect 21456 4088 21508 4140
rect 22652 4088 22704 4140
rect 17868 3952 17920 4004
rect 22284 4020 22336 4072
rect 22836 4020 22888 4072
rect 23296 4020 23348 4072
rect 24768 4088 24820 4140
rect 38844 4131 38896 4140
rect 38844 4097 38853 4131
rect 38853 4097 38887 4131
rect 38887 4097 38896 4131
rect 38844 4088 38896 4097
rect 38752 4020 38804 4072
rect 20352 3952 20404 4004
rect 30748 3952 30800 4004
rect 30932 3995 30984 4004
rect 30932 3961 30941 3995
rect 30941 3961 30975 3995
rect 30975 3961 30984 3995
rect 30932 3952 30984 3961
rect 39488 3952 39540 4004
rect 19616 3884 19668 3936
rect 22560 3884 22612 3936
rect 23296 3884 23348 3936
rect 23388 3884 23440 3936
rect 24860 3884 24912 3936
rect 30288 3884 30340 3936
rect 39028 3927 39080 3936
rect 39028 3893 39037 3927
rect 39037 3893 39071 3927
rect 39071 3893 39080 3927
rect 39028 3884 39080 3893
rect 1950 3782 2002 3834
rect 2014 3782 2066 3834
rect 2078 3782 2130 3834
rect 2142 3782 2194 3834
rect 2206 3782 2258 3834
rect 7950 3782 8002 3834
rect 8014 3782 8066 3834
rect 8078 3782 8130 3834
rect 8142 3782 8194 3834
rect 8206 3782 8258 3834
rect 13950 3782 14002 3834
rect 14014 3782 14066 3834
rect 14078 3782 14130 3834
rect 14142 3782 14194 3834
rect 14206 3782 14258 3834
rect 19950 3782 20002 3834
rect 20014 3782 20066 3834
rect 20078 3782 20130 3834
rect 20142 3782 20194 3834
rect 20206 3782 20258 3834
rect 25950 3782 26002 3834
rect 26014 3782 26066 3834
rect 26078 3782 26130 3834
rect 26142 3782 26194 3834
rect 26206 3782 26258 3834
rect 31950 3782 32002 3834
rect 32014 3782 32066 3834
rect 32078 3782 32130 3834
rect 32142 3782 32194 3834
rect 32206 3782 32258 3834
rect 37950 3782 38002 3834
rect 38014 3782 38066 3834
rect 38078 3782 38130 3834
rect 38142 3782 38194 3834
rect 38206 3782 38258 3834
rect 9496 3680 9548 3732
rect 13636 3680 13688 3732
rect 14372 3680 14424 3732
rect 15384 3723 15436 3732
rect 15384 3689 15393 3723
rect 15393 3689 15427 3723
rect 15427 3689 15436 3723
rect 15384 3680 15436 3689
rect 11336 3587 11388 3596
rect 11336 3553 11345 3587
rect 11345 3553 11379 3587
rect 11379 3553 11388 3587
rect 11336 3544 11388 3553
rect 11520 3587 11572 3596
rect 11520 3553 11538 3587
rect 11538 3553 11572 3587
rect 11520 3544 11572 3553
rect 11612 3587 11664 3596
rect 11612 3553 11621 3587
rect 11621 3553 11655 3587
rect 11655 3553 11664 3587
rect 11612 3544 11664 3553
rect 13728 3612 13780 3664
rect 8484 3476 8536 3528
rect 12992 3544 13044 3596
rect 16580 3587 16632 3596
rect 16580 3553 16589 3587
rect 16589 3553 16623 3587
rect 16623 3553 16632 3587
rect 16580 3544 16632 3553
rect 16764 3587 16816 3596
rect 16764 3553 16782 3587
rect 16782 3553 16816 3587
rect 16764 3544 16816 3553
rect 17684 3612 17736 3664
rect 18144 3680 18196 3732
rect 19524 3612 19576 3664
rect 21364 3612 21416 3664
rect 14464 3476 14516 3528
rect 15476 3519 15528 3528
rect 15476 3485 15484 3519
rect 15484 3485 15518 3519
rect 15518 3485 15528 3519
rect 15476 3476 15528 3485
rect 15660 3476 15712 3528
rect 16304 3340 16356 3392
rect 17776 3587 17828 3596
rect 17776 3553 17785 3587
rect 17785 3553 17819 3587
rect 17819 3553 17828 3587
rect 17776 3544 17828 3553
rect 18052 3476 18104 3528
rect 19432 3476 19484 3528
rect 19800 3544 19852 3596
rect 19616 3519 19668 3528
rect 19616 3485 19625 3519
rect 19625 3485 19659 3519
rect 19659 3485 19668 3519
rect 19616 3476 19668 3485
rect 20536 3476 20588 3528
rect 22008 3680 22060 3732
rect 22100 3680 22152 3732
rect 23020 3680 23072 3732
rect 23296 3680 23348 3732
rect 22560 3612 22612 3664
rect 22652 3544 22704 3596
rect 23480 3544 23532 3596
rect 21640 3476 21692 3528
rect 23296 3519 23348 3528
rect 23296 3485 23305 3519
rect 23305 3485 23339 3519
rect 23339 3485 23348 3519
rect 23296 3476 23348 3485
rect 25872 3680 25924 3732
rect 30104 3723 30156 3732
rect 30104 3689 30113 3723
rect 30113 3689 30147 3723
rect 30147 3689 30156 3723
rect 30104 3680 30156 3689
rect 30656 3723 30708 3732
rect 30656 3689 30665 3723
rect 30665 3689 30699 3723
rect 30699 3689 30708 3723
rect 30656 3680 30708 3689
rect 33416 3680 33468 3732
rect 35716 3680 35768 3732
rect 39396 3723 39448 3732
rect 39396 3689 39405 3723
rect 39405 3689 39439 3723
rect 39439 3689 39448 3723
rect 39396 3680 39448 3689
rect 24216 3612 24268 3664
rect 24492 3612 24544 3664
rect 38384 3612 38436 3664
rect 20812 3408 20864 3460
rect 22284 3408 22336 3460
rect 18696 3340 18748 3392
rect 19340 3383 19392 3392
rect 19340 3349 19349 3383
rect 19349 3349 19383 3383
rect 19383 3349 19392 3383
rect 19340 3340 19392 3349
rect 23480 3340 23532 3392
rect 23572 3340 23624 3392
rect 29920 3519 29972 3528
rect 29920 3485 29929 3519
rect 29929 3485 29963 3519
rect 29963 3485 29972 3519
rect 29920 3476 29972 3485
rect 37464 3544 37516 3596
rect 31208 3519 31260 3528
rect 31208 3485 31217 3519
rect 31217 3485 31251 3519
rect 31251 3485 31260 3519
rect 31208 3476 31260 3485
rect 35808 3476 35860 3528
rect 26332 3451 26384 3460
rect 26332 3417 26341 3451
rect 26341 3417 26375 3451
rect 26375 3417 26384 3451
rect 26332 3408 26384 3417
rect 34520 3408 34572 3460
rect 39212 3519 39264 3528
rect 39212 3485 39221 3519
rect 39221 3485 39255 3519
rect 39255 3485 39264 3519
rect 39212 3476 39264 3485
rect 35348 3383 35400 3392
rect 35348 3349 35357 3383
rect 35357 3349 35391 3383
rect 35391 3349 35400 3383
rect 35348 3340 35400 3349
rect 37372 3340 37424 3392
rect 37740 3383 37792 3392
rect 37740 3349 37749 3383
rect 37749 3349 37783 3383
rect 37783 3349 37792 3383
rect 37740 3340 37792 3349
rect 38292 3340 38344 3392
rect 38660 3383 38712 3392
rect 38660 3349 38669 3383
rect 38669 3349 38703 3383
rect 38703 3349 38712 3383
rect 38660 3340 38712 3349
rect 3010 3238 3062 3290
rect 3074 3238 3126 3290
rect 3138 3238 3190 3290
rect 3202 3238 3254 3290
rect 3266 3238 3318 3290
rect 9010 3238 9062 3290
rect 9074 3238 9126 3290
rect 9138 3238 9190 3290
rect 9202 3238 9254 3290
rect 9266 3238 9318 3290
rect 15010 3238 15062 3290
rect 15074 3238 15126 3290
rect 15138 3238 15190 3290
rect 15202 3238 15254 3290
rect 15266 3238 15318 3290
rect 21010 3238 21062 3290
rect 21074 3238 21126 3290
rect 21138 3238 21190 3290
rect 21202 3238 21254 3290
rect 21266 3238 21318 3290
rect 27010 3238 27062 3290
rect 27074 3238 27126 3290
rect 27138 3238 27190 3290
rect 27202 3238 27254 3290
rect 27266 3238 27318 3290
rect 33010 3238 33062 3290
rect 33074 3238 33126 3290
rect 33138 3238 33190 3290
rect 33202 3238 33254 3290
rect 33266 3238 33318 3290
rect 39010 3238 39062 3290
rect 39074 3238 39126 3290
rect 39138 3238 39190 3290
rect 39202 3238 39254 3290
rect 39266 3238 39318 3290
rect 3516 3136 3568 3188
rect 15200 3136 15252 3188
rect 22192 3136 22244 3188
rect 39396 3136 39448 3188
rect 7012 3068 7064 3120
rect 19340 3068 19392 3120
rect 23112 3068 23164 3120
rect 20904 3000 20956 3052
rect 22560 3000 22612 3052
rect 22928 3000 22980 3052
rect 38476 3043 38528 3052
rect 38476 3009 38485 3043
rect 38485 3009 38519 3043
rect 38519 3009 38528 3043
rect 38476 3000 38528 3009
rect 38844 3043 38896 3052
rect 38844 3009 38853 3043
rect 38853 3009 38887 3043
rect 38887 3009 38896 3043
rect 38844 3000 38896 3009
rect 39212 3043 39264 3052
rect 39212 3009 39221 3043
rect 39221 3009 39255 3043
rect 39255 3009 39264 3043
rect 39212 3000 39264 3009
rect 22008 2932 22060 2984
rect 35348 2932 35400 2984
rect 13728 2864 13780 2916
rect 23204 2864 23256 2916
rect 39488 2864 39540 2916
rect 9864 2796 9916 2848
rect 19248 2796 19300 2848
rect 26332 2796 26384 2848
rect 38844 2796 38896 2848
rect 1950 2694 2002 2746
rect 2014 2694 2066 2746
rect 2078 2694 2130 2746
rect 2142 2694 2194 2746
rect 2206 2694 2258 2746
rect 7950 2694 8002 2746
rect 8014 2694 8066 2746
rect 8078 2694 8130 2746
rect 8142 2694 8194 2746
rect 8206 2694 8258 2746
rect 13950 2694 14002 2746
rect 14014 2694 14066 2746
rect 14078 2694 14130 2746
rect 14142 2694 14194 2746
rect 14206 2694 14258 2746
rect 19950 2694 20002 2746
rect 20014 2694 20066 2746
rect 20078 2694 20130 2746
rect 20142 2694 20194 2746
rect 20206 2694 20258 2746
rect 25950 2694 26002 2746
rect 26014 2694 26066 2746
rect 26078 2694 26130 2746
rect 26142 2694 26194 2746
rect 26206 2694 26258 2746
rect 31950 2694 32002 2746
rect 32014 2694 32066 2746
rect 32078 2694 32130 2746
rect 32142 2694 32194 2746
rect 32206 2694 32258 2746
rect 37950 2694 38002 2746
rect 38014 2694 38066 2746
rect 38078 2694 38130 2746
rect 38142 2694 38194 2746
rect 38206 2694 38258 2746
rect 6920 2592 6972 2644
rect 38936 2592 38988 2644
rect 39396 2635 39448 2644
rect 39396 2601 39405 2635
rect 39405 2601 39439 2635
rect 39439 2601 39448 2635
rect 39396 2592 39448 2601
rect 1308 2524 1360 2576
rect 35808 2524 35860 2576
rect 37556 2567 37608 2576
rect 37556 2533 37565 2567
rect 37565 2533 37599 2567
rect 37599 2533 37608 2567
rect 37556 2524 37608 2533
rect 39948 2524 40000 2576
rect 2044 2431 2096 2440
rect 2044 2397 2053 2431
rect 2053 2397 2087 2431
rect 2087 2397 2096 2431
rect 2044 2388 2096 2397
rect 14832 2456 14884 2508
rect 15200 2456 15252 2508
rect 6736 2431 6788 2440
rect 6736 2397 6745 2431
rect 6745 2397 6779 2431
rect 6779 2397 6788 2431
rect 6736 2388 6788 2397
rect 9496 2388 9548 2440
rect 9864 2431 9916 2440
rect 9864 2397 9873 2431
rect 9873 2397 9907 2431
rect 9907 2397 9916 2431
rect 9864 2388 9916 2397
rect 5540 2320 5592 2372
rect 37372 2431 37424 2440
rect 37372 2397 37381 2431
rect 37381 2397 37415 2431
rect 37415 2397 37424 2431
rect 37372 2388 37424 2397
rect 38292 2456 38344 2508
rect 38384 2388 38436 2440
rect 38752 2388 38804 2440
rect 1676 2252 1728 2304
rect 3424 2295 3476 2304
rect 3424 2261 3433 2295
rect 3433 2261 3467 2295
rect 3467 2261 3476 2295
rect 3424 2252 3476 2261
rect 4804 2252 4856 2304
rect 6368 2252 6420 2304
rect 37832 2295 37884 2304
rect 37832 2261 37841 2295
rect 37841 2261 37875 2295
rect 37875 2261 37884 2295
rect 37832 2252 37884 2261
rect 38292 2295 38344 2304
rect 38292 2261 38301 2295
rect 38301 2261 38335 2295
rect 38335 2261 38344 2295
rect 38292 2252 38344 2261
rect 38660 2295 38712 2304
rect 38660 2261 38669 2295
rect 38669 2261 38703 2295
rect 38703 2261 38712 2295
rect 38660 2252 38712 2261
rect 3010 2150 3062 2202
rect 3074 2150 3126 2202
rect 3138 2150 3190 2202
rect 3202 2150 3254 2202
rect 3266 2150 3318 2202
rect 9010 2150 9062 2202
rect 9074 2150 9126 2202
rect 9138 2150 9190 2202
rect 9202 2150 9254 2202
rect 9266 2150 9318 2202
rect 15010 2150 15062 2202
rect 15074 2150 15126 2202
rect 15138 2150 15190 2202
rect 15202 2150 15254 2202
rect 15266 2150 15318 2202
rect 21010 2150 21062 2202
rect 21074 2150 21126 2202
rect 21138 2150 21190 2202
rect 21202 2150 21254 2202
rect 21266 2150 21318 2202
rect 27010 2150 27062 2202
rect 27074 2150 27126 2202
rect 27138 2150 27190 2202
rect 27202 2150 27254 2202
rect 27266 2150 27318 2202
rect 33010 2150 33062 2202
rect 33074 2150 33126 2202
rect 33138 2150 33190 2202
rect 33202 2150 33254 2202
rect 33266 2150 33318 2202
rect 39010 2150 39062 2202
rect 39074 2150 39126 2202
rect 39138 2150 39190 2202
rect 39202 2150 39254 2202
rect 39266 2150 39318 2202
rect 6736 2048 6788 2100
rect 17500 2048 17552 2100
rect 20444 2048 20496 2100
rect 31208 2048 31260 2100
rect 4712 1980 4764 2032
rect 25136 824 25188 876
rect 26884 824 26936 876
rect 14188 144 14240 196
rect 25044 144 25096 196
rect 18972 76 19024 128
rect 31576 76 31628 128
rect 8024 8 8076 60
rect 29920 8 29972 60
<< metal2 >>
rect 3238 11194 3294 11250
rect 3514 11194 3570 11250
rect 3790 11194 3846 11250
rect 3884 11212 3936 11218
rect 1122 9888 1178 9897
rect 1122 9823 1178 9832
rect 1030 9616 1086 9625
rect 1030 9551 1086 9560
rect 846 9344 902 9353
rect 846 9279 902 9288
rect 664 8968 716 8974
rect 664 8910 716 8916
rect 572 8492 624 8498
rect 572 8434 624 8440
rect 584 7993 612 8434
rect 570 7984 626 7993
rect 570 7919 626 7928
rect 572 7812 624 7818
rect 572 7754 624 7760
rect 584 7449 612 7754
rect 570 7440 626 7449
rect 570 7375 626 7384
rect 676 6914 704 8910
rect 860 8430 888 9279
rect 938 8800 994 8809
rect 938 8735 994 8744
rect 848 8424 900 8430
rect 848 8366 900 8372
rect 756 7880 808 7886
rect 756 7822 808 7828
rect 768 7721 796 7822
rect 754 7712 810 7721
rect 754 7647 810 7656
rect 952 7478 980 8735
rect 1044 8362 1072 9551
rect 1136 8634 1164 9823
rect 2688 9512 2740 9518
rect 2688 9454 2740 9460
rect 3252 9466 3280 11194
rect 2136 9172 2188 9178
rect 2136 9114 2188 9120
rect 1214 9072 1270 9081
rect 1214 9007 1270 9016
rect 2044 9036 2096 9042
rect 1124 8628 1176 8634
rect 1124 8570 1176 8576
rect 1122 8392 1178 8401
rect 1032 8356 1084 8362
rect 1122 8327 1178 8336
rect 1032 8298 1084 8304
rect 1030 8256 1086 8265
rect 1030 8191 1086 8200
rect 1044 7954 1072 8191
rect 1032 7948 1084 7954
rect 1032 7890 1084 7896
rect 940 7472 992 7478
rect 940 7414 992 7420
rect 756 7404 808 7410
rect 756 7346 808 7352
rect 768 7177 796 7346
rect 940 7336 992 7342
rect 940 7278 992 7284
rect 754 7168 810 7177
rect 754 7103 810 7112
rect 584 6886 704 6914
rect 952 6905 980 7278
rect 1136 6914 1164 8327
rect 1228 8090 1256 9007
rect 2044 8978 2096 8984
rect 1584 8832 1636 8838
rect 1584 8774 1636 8780
rect 1308 8560 1360 8566
rect 1306 8528 1308 8537
rect 1360 8528 1362 8537
rect 1306 8463 1362 8472
rect 1596 8294 1624 8774
rect 2056 8362 2084 8978
rect 2148 8362 2176 9114
rect 2412 8900 2464 8906
rect 2412 8842 2464 8848
rect 2424 8634 2452 8842
rect 2700 8634 2728 9454
rect 3252 9438 3464 9466
rect 3010 8732 3318 8741
rect 3010 8730 3016 8732
rect 3072 8730 3096 8732
rect 3152 8730 3176 8732
rect 3232 8730 3256 8732
rect 3312 8730 3318 8732
rect 3072 8678 3074 8730
rect 3254 8678 3256 8730
rect 3010 8676 3016 8678
rect 3072 8676 3096 8678
rect 3152 8676 3176 8678
rect 3232 8676 3256 8678
rect 3312 8676 3318 8678
rect 3010 8667 3318 8676
rect 2412 8628 2464 8634
rect 2412 8570 2464 8576
rect 2688 8628 2740 8634
rect 2688 8570 2740 8576
rect 2044 8356 2096 8362
rect 2044 8298 2096 8304
rect 2136 8356 2188 8362
rect 2136 8298 2188 8304
rect 1584 8288 1636 8294
rect 1584 8230 1636 8236
rect 2320 8288 2372 8294
rect 2320 8230 2372 8236
rect 1950 8188 2258 8197
rect 1950 8186 1956 8188
rect 2012 8186 2036 8188
rect 2092 8186 2116 8188
rect 2172 8186 2196 8188
rect 2252 8186 2258 8188
rect 2012 8134 2014 8186
rect 2194 8134 2196 8186
rect 1950 8132 1956 8134
rect 2012 8132 2036 8134
rect 2092 8132 2116 8134
rect 2172 8132 2196 8134
rect 2252 8132 2258 8134
rect 1950 8123 2258 8132
rect 1216 8084 1268 8090
rect 1216 8026 1268 8032
rect 1952 8016 2004 8022
rect 1306 7984 1362 7993
rect 2004 7964 2176 7970
rect 1952 7958 2176 7964
rect 1964 7954 2176 7958
rect 1964 7948 2188 7954
rect 1964 7942 2136 7948
rect 1306 7919 1362 7928
rect 938 6896 994 6905
rect 584 6633 612 6886
rect 1136 6886 1256 6914
rect 938 6831 994 6840
rect 570 6624 626 6633
rect 570 6559 626 6568
rect 1228 5545 1256 6886
rect 1214 5536 1270 5545
rect 1214 5471 1270 5480
rect 664 5228 716 5234
rect 664 5170 716 5176
rect 676 4185 704 5170
rect 1320 4729 1348 7919
rect 2136 7890 2188 7896
rect 2136 7744 2188 7750
rect 2136 7686 2188 7692
rect 2148 7478 2176 7686
rect 2136 7472 2188 7478
rect 2136 7414 2188 7420
rect 2332 7206 2360 8230
rect 3436 8090 3464 9438
rect 3528 8362 3556 11194
rect 3606 9208 3662 9217
rect 3606 9143 3662 9152
rect 3516 8356 3568 8362
rect 3516 8298 3568 8304
rect 3424 8084 3476 8090
rect 3424 8026 3476 8032
rect 3516 8084 3568 8090
rect 3516 8026 3568 8032
rect 3010 7644 3318 7653
rect 3010 7642 3016 7644
rect 3072 7642 3096 7644
rect 3152 7642 3176 7644
rect 3232 7642 3256 7644
rect 3312 7642 3318 7644
rect 3072 7590 3074 7642
rect 3254 7590 3256 7642
rect 3010 7588 3016 7590
rect 3072 7588 3096 7590
rect 3152 7588 3176 7590
rect 3232 7588 3256 7590
rect 3312 7588 3318 7590
rect 3010 7579 3318 7588
rect 3528 7410 3556 8026
rect 3620 7886 3648 9143
rect 3804 8634 3832 11194
rect 4066 11194 4122 11250
rect 4342 11194 4398 11250
rect 4618 11194 4674 11250
rect 4894 11194 4950 11250
rect 5170 11194 5226 11250
rect 5446 11194 5502 11250
rect 5722 11194 5778 11250
rect 5998 11194 6054 11250
rect 6274 11194 6330 11250
rect 6550 11194 6606 11250
rect 6826 11194 6882 11250
rect 7102 11194 7158 11250
rect 7378 11194 7434 11250
rect 7654 11194 7710 11250
rect 7930 11194 7986 11250
rect 8206 11194 8262 11250
rect 8482 11194 8538 11250
rect 8758 11194 8814 11250
rect 9034 11194 9090 11250
rect 9310 11194 9366 11250
rect 9586 11194 9642 11250
rect 9862 11194 9918 11250
rect 10138 11194 10194 11250
rect 10414 11194 10470 11250
rect 10690 11194 10746 11250
rect 10966 11194 11022 11250
rect 11242 11194 11298 11250
rect 11518 11194 11574 11250
rect 11794 11194 11850 11250
rect 12070 11194 12126 11250
rect 12346 11194 12402 11250
rect 12622 11194 12678 11250
rect 12898 11194 12954 11250
rect 13174 11194 13230 11250
rect 13450 11194 13506 11250
rect 13726 11194 13782 11250
rect 14002 11194 14058 11250
rect 14278 11194 14334 11250
rect 14554 11194 14610 11250
rect 14830 11194 14886 11250
rect 15106 11194 15162 11250
rect 15382 11194 15438 11250
rect 15658 11194 15714 11250
rect 15934 11194 15990 11250
rect 16210 11194 16266 11250
rect 16486 11194 16542 11250
rect 16762 11194 16818 11250
rect 17038 11194 17094 11250
rect 17314 11194 17370 11250
rect 17590 11194 17646 11250
rect 17866 11194 17922 11250
rect 18142 11194 18198 11250
rect 18418 11194 18474 11250
rect 18694 11194 18750 11250
rect 18970 11194 19026 11250
rect 19246 11194 19302 11250
rect 19522 11194 19578 11250
rect 19798 11194 19854 11250
rect 20074 11212 20130 11250
rect 20074 11194 20076 11212
rect 3884 11154 3936 11160
rect 3792 8628 3844 8634
rect 3792 8570 3844 8576
rect 3700 8492 3752 8498
rect 3700 8434 3752 8440
rect 3608 7880 3660 7886
rect 3608 7822 3660 7828
rect 2872 7404 2924 7410
rect 2872 7346 2924 7352
rect 3424 7404 3476 7410
rect 3424 7346 3476 7352
rect 3516 7404 3568 7410
rect 3516 7346 3568 7352
rect 2320 7200 2372 7206
rect 2320 7142 2372 7148
rect 1950 7100 2258 7109
rect 1950 7098 1956 7100
rect 2012 7098 2036 7100
rect 2092 7098 2116 7100
rect 2172 7098 2196 7100
rect 2252 7098 2258 7100
rect 2012 7046 2014 7098
rect 2194 7046 2196 7098
rect 1950 7044 1956 7046
rect 2012 7044 2036 7046
rect 2092 7044 2116 7046
rect 2172 7044 2196 7046
rect 2252 7044 2258 7046
rect 1950 7035 2258 7044
rect 2780 6724 2832 6730
rect 2780 6666 2832 6672
rect 1950 6012 2258 6021
rect 1950 6010 1956 6012
rect 2012 6010 2036 6012
rect 2092 6010 2116 6012
rect 2172 6010 2196 6012
rect 2252 6010 2258 6012
rect 2012 5958 2014 6010
rect 2194 5958 2196 6010
rect 1950 5956 1956 5958
rect 2012 5956 2036 5958
rect 2092 5956 2116 5958
rect 2172 5956 2196 5958
rect 2252 5956 2258 5958
rect 1950 5947 2258 5956
rect 2792 5137 2820 6666
rect 2884 6361 2912 7346
rect 3056 7268 3108 7274
rect 3056 7210 3108 7216
rect 3068 6905 3096 7210
rect 3054 6896 3110 6905
rect 3054 6831 3110 6840
rect 3010 6556 3318 6565
rect 3010 6554 3016 6556
rect 3072 6554 3096 6556
rect 3152 6554 3176 6556
rect 3232 6554 3256 6556
rect 3312 6554 3318 6556
rect 3072 6502 3074 6554
rect 3254 6502 3256 6554
rect 3010 6500 3016 6502
rect 3072 6500 3096 6502
rect 3152 6500 3176 6502
rect 3232 6500 3256 6502
rect 3312 6500 3318 6502
rect 3010 6491 3318 6500
rect 2870 6352 2926 6361
rect 2870 6287 2926 6296
rect 3436 6225 3464 7346
rect 3608 7200 3660 7206
rect 3608 7142 3660 7148
rect 3516 6724 3568 6730
rect 3516 6666 3568 6672
rect 3422 6216 3478 6225
rect 3422 6151 3478 6160
rect 2872 5636 2924 5642
rect 2872 5578 2924 5584
rect 2778 5128 2834 5137
rect 2778 5063 2834 5072
rect 1950 4924 2258 4933
rect 1950 4922 1956 4924
rect 2012 4922 2036 4924
rect 2092 4922 2116 4924
rect 2172 4922 2196 4924
rect 2252 4922 2258 4924
rect 2012 4870 2014 4922
rect 2194 4870 2196 4922
rect 1950 4868 1956 4870
rect 2012 4868 2036 4870
rect 2092 4868 2116 4870
rect 2172 4868 2196 4870
rect 2252 4868 2258 4870
rect 1950 4859 2258 4868
rect 1306 4720 1362 4729
rect 1306 4655 1362 4664
rect 2780 4548 2832 4554
rect 2780 4490 2832 4496
rect 1216 4276 1268 4282
rect 1216 4218 1268 4224
rect 662 4176 718 4185
rect 662 4111 718 4120
rect 1228 1737 1256 4218
rect 1308 4208 1360 4214
rect 1308 4150 1360 4156
rect 1320 3097 1348 4150
rect 1950 3836 2258 3845
rect 1950 3834 1956 3836
rect 2012 3834 2036 3836
rect 2092 3834 2116 3836
rect 2172 3834 2196 3836
rect 2252 3834 2258 3836
rect 2012 3782 2014 3834
rect 2194 3782 2196 3834
rect 1950 3780 1956 3782
rect 2012 3780 2036 3782
rect 2092 3780 2116 3782
rect 2172 3780 2196 3782
rect 2252 3780 2258 3782
rect 1950 3771 2258 3780
rect 2792 3641 2820 4490
rect 2884 4457 2912 5578
rect 3010 5468 3318 5477
rect 3010 5466 3016 5468
rect 3072 5466 3096 5468
rect 3152 5466 3176 5468
rect 3232 5466 3256 5468
rect 3312 5466 3318 5468
rect 3072 5414 3074 5466
rect 3254 5414 3256 5466
rect 3010 5412 3016 5414
rect 3072 5412 3096 5414
rect 3152 5412 3176 5414
rect 3232 5412 3256 5414
rect 3312 5412 3318 5414
rect 3010 5403 3318 5412
rect 3424 5228 3476 5234
rect 3424 5170 3476 5176
rect 2870 4448 2926 4457
rect 2870 4383 2926 4392
rect 3010 4380 3318 4389
rect 3010 4378 3016 4380
rect 3072 4378 3096 4380
rect 3152 4378 3176 4380
rect 3232 4378 3256 4380
rect 3312 4378 3318 4380
rect 3072 4326 3074 4378
rect 3254 4326 3256 4378
rect 3010 4324 3016 4326
rect 3072 4324 3096 4326
rect 3152 4324 3176 4326
rect 3232 4324 3256 4326
rect 3312 4324 3318 4326
rect 3010 4315 3318 4324
rect 2872 4140 2924 4146
rect 2872 4082 2924 4088
rect 2778 3632 2834 3641
rect 2778 3567 2834 3576
rect 2884 3369 2912 4082
rect 3436 4049 3464 5170
rect 3528 4758 3556 6666
rect 3516 4752 3568 4758
rect 3516 4694 3568 4700
rect 3620 4298 3648 7142
rect 3712 6662 3740 8434
rect 3896 8090 3924 11154
rect 3976 8424 4028 8430
rect 3976 8366 4028 8372
rect 3884 8084 3936 8090
rect 3884 8026 3936 8032
rect 3884 7948 3936 7954
rect 3884 7890 3936 7896
rect 3792 7472 3844 7478
rect 3792 7414 3844 7420
rect 3804 7002 3832 7414
rect 3792 6996 3844 7002
rect 3792 6938 3844 6944
rect 3700 6656 3752 6662
rect 3700 6598 3752 6604
rect 3896 6254 3924 7890
rect 3988 6662 4016 8366
rect 4080 8090 4108 11194
rect 4356 8634 4384 11194
rect 4632 8634 4660 11194
rect 4344 8628 4396 8634
rect 4344 8570 4396 8576
rect 4620 8628 4672 8634
rect 4620 8570 4672 8576
rect 4528 8492 4580 8498
rect 4528 8434 4580 8440
rect 4068 8084 4120 8090
rect 4068 8026 4120 8032
rect 4540 7546 4568 8434
rect 4908 8090 4936 11194
rect 5184 8634 5212 11194
rect 5460 8634 5488 11194
rect 5630 10432 5686 10441
rect 5630 10367 5686 10376
rect 5172 8628 5224 8634
rect 5172 8570 5224 8576
rect 5448 8628 5500 8634
rect 5448 8570 5500 8576
rect 5644 8498 5672 10367
rect 5736 8634 5764 11194
rect 5816 9648 5868 9654
rect 5816 9590 5868 9596
rect 5724 8628 5776 8634
rect 5724 8570 5776 8576
rect 5828 8498 5856 9590
rect 5632 8492 5684 8498
rect 5632 8434 5684 8440
rect 5816 8492 5868 8498
rect 5816 8434 5868 8440
rect 6012 8090 6040 11194
rect 6288 8634 6316 11194
rect 6276 8628 6328 8634
rect 6276 8570 6328 8576
rect 6564 8090 6592 11194
rect 6642 10296 6698 10305
rect 6642 10231 6698 10240
rect 4896 8084 4948 8090
rect 4896 8026 4948 8032
rect 6000 8084 6052 8090
rect 6000 8026 6052 8032
rect 6552 8084 6604 8090
rect 6552 8026 6604 8032
rect 4712 7880 4764 7886
rect 4712 7822 4764 7828
rect 4724 7546 4752 7822
rect 6184 7812 6236 7818
rect 6184 7754 6236 7760
rect 6196 7546 6224 7754
rect 6276 7744 6328 7750
rect 6276 7686 6328 7692
rect 4528 7540 4580 7546
rect 4528 7482 4580 7488
rect 4712 7540 4764 7546
rect 4712 7482 4764 7488
rect 6184 7540 6236 7546
rect 6184 7482 6236 7488
rect 6288 7410 6316 7686
rect 4068 7404 4120 7410
rect 4068 7346 4120 7352
rect 6276 7404 6328 7410
rect 6276 7346 6328 7352
rect 3976 6656 4028 6662
rect 3976 6598 4028 6604
rect 3884 6248 3936 6254
rect 3884 6190 3936 6196
rect 4080 5817 4108 7346
rect 4436 7268 4488 7274
rect 4436 7210 4488 7216
rect 4066 5808 4122 5817
rect 4066 5743 4122 5752
rect 4448 5273 4476 7210
rect 5540 6180 5592 6186
rect 5540 6122 5592 6128
rect 4434 5264 4490 5273
rect 4434 5199 4490 5208
rect 4068 5092 4120 5098
rect 4068 5034 4120 5040
rect 3976 5024 4028 5030
rect 3976 4966 4028 4972
rect 3884 4684 3936 4690
rect 3884 4626 3936 4632
rect 3620 4270 3740 4298
rect 3608 4208 3660 4214
rect 3712 4185 3740 4270
rect 3608 4150 3660 4156
rect 3698 4176 3754 4185
rect 3422 4040 3478 4049
rect 3056 4004 3108 4010
rect 3422 3975 3478 3984
rect 3056 3946 3108 3952
rect 3068 3505 3096 3946
rect 3516 3936 3568 3942
rect 3516 3878 3568 3884
rect 3054 3496 3110 3505
rect 3054 3431 3110 3440
rect 2870 3360 2926 3369
rect 2870 3295 2926 3304
rect 3010 3292 3318 3301
rect 3010 3290 3016 3292
rect 3072 3290 3096 3292
rect 3152 3290 3176 3292
rect 3232 3290 3256 3292
rect 3312 3290 3318 3292
rect 3072 3238 3074 3290
rect 3254 3238 3256 3290
rect 3010 3236 3016 3238
rect 3072 3236 3096 3238
rect 3152 3236 3176 3238
rect 3232 3236 3256 3238
rect 3312 3236 3318 3238
rect 3010 3227 3318 3236
rect 3528 3194 3556 3878
rect 3516 3188 3568 3194
rect 3516 3130 3568 3136
rect 1306 3088 1362 3097
rect 1306 3023 1362 3032
rect 3620 2961 3648 4150
rect 3698 4111 3754 4120
rect 3792 4004 3844 4010
rect 3792 3946 3844 3952
rect 3804 3097 3832 3946
rect 3790 3088 3846 3097
rect 3790 3023 3846 3032
rect 3896 2961 3924 4626
rect 3988 3641 4016 4966
rect 4080 4049 4108 5034
rect 4712 4072 4764 4078
rect 4066 4040 4122 4049
rect 4712 4014 4764 4020
rect 4066 3975 4122 3984
rect 3974 3632 4030 3641
rect 3974 3567 4030 3576
rect 3606 2952 3662 2961
rect 3606 2887 3662 2896
rect 3882 2952 3938 2961
rect 3882 2887 3938 2896
rect 1950 2748 2258 2757
rect 1950 2746 1956 2748
rect 2012 2746 2036 2748
rect 2092 2746 2116 2748
rect 2172 2746 2196 2748
rect 2252 2746 2258 2748
rect 2012 2694 2014 2746
rect 2194 2694 2196 2746
rect 1950 2692 1956 2694
rect 2012 2692 2036 2694
rect 2092 2692 2116 2694
rect 2172 2692 2196 2694
rect 2252 2692 2258 2694
rect 1950 2683 2258 2692
rect 1308 2576 1360 2582
rect 1306 2544 1308 2553
rect 1360 2544 1362 2553
rect 1306 2479 1362 2488
rect 2044 2440 2096 2446
rect 2042 2408 2044 2417
rect 2096 2408 2098 2417
rect 2042 2343 2098 2352
rect 1676 2304 1728 2310
rect 3424 2304 3476 2310
rect 1676 2246 1728 2252
rect 2870 2272 2926 2281
rect 1214 1728 1270 1737
rect 1214 1663 1270 1672
rect 1688 56 1716 2246
rect 3424 2246 3476 2252
rect 2870 2207 2926 2216
rect 2884 1737 2912 2207
rect 3010 2204 3318 2213
rect 3010 2202 3016 2204
rect 3072 2202 3096 2204
rect 3152 2202 3176 2204
rect 3232 2202 3256 2204
rect 3312 2202 3318 2204
rect 3072 2150 3074 2202
rect 3254 2150 3256 2202
rect 3010 2148 3016 2150
rect 3072 2148 3096 2150
rect 3152 2148 3176 2150
rect 3232 2148 3256 2150
rect 3312 2148 3318 2150
rect 3010 2139 3318 2148
rect 2870 1728 2926 1737
rect 2870 1663 2926 1672
rect 3252 56 3372 82
rect 1674 0 1730 56
rect 3238 54 3372 56
rect 3238 0 3294 54
rect 3344 42 3372 54
rect 3436 42 3464 2246
rect 4724 2038 4752 4014
rect 5552 2378 5580 6122
rect 6656 5710 6684 10231
rect 6734 10024 6790 10033
rect 6734 9959 6790 9968
rect 6748 8906 6776 9959
rect 6736 8900 6788 8906
rect 6736 8842 6788 8848
rect 6840 8634 6868 11194
rect 6920 9308 6972 9314
rect 6920 9250 6972 9256
rect 6828 8628 6880 8634
rect 6828 8570 6880 8576
rect 6932 8498 6960 9250
rect 6920 8492 6972 8498
rect 6920 8434 6972 8440
rect 7012 8424 7064 8430
rect 7012 8366 7064 8372
rect 6920 8016 6972 8022
rect 6920 7958 6972 7964
rect 6932 5846 6960 7958
rect 6920 5840 6972 5846
rect 6920 5782 6972 5788
rect 6644 5704 6696 5710
rect 6644 5646 6696 5652
rect 6656 4078 6684 5646
rect 6920 5636 6972 5642
rect 6920 5578 6972 5584
rect 6644 4072 6696 4078
rect 6644 4014 6696 4020
rect 6932 2650 6960 5578
rect 7024 3126 7052 8366
rect 7116 8090 7144 11194
rect 7196 10124 7248 10130
rect 7196 10066 7248 10072
rect 7104 8084 7156 8090
rect 7104 8026 7156 8032
rect 7208 7886 7236 10066
rect 7288 8900 7340 8906
rect 7288 8842 7340 8848
rect 7300 8498 7328 8842
rect 7392 8634 7420 11194
rect 7564 9240 7616 9246
rect 7564 9182 7616 9188
rect 7380 8628 7432 8634
rect 7380 8570 7432 8576
rect 7288 8492 7340 8498
rect 7288 8434 7340 8440
rect 7196 7880 7248 7886
rect 7196 7822 7248 7828
rect 7472 7336 7524 7342
rect 7472 7278 7524 7284
rect 7576 7290 7604 9182
rect 7668 8634 7696 11194
rect 7840 11144 7892 11150
rect 7840 11086 7892 11092
rect 7748 9716 7800 9722
rect 7748 9658 7800 9664
rect 7656 8628 7708 8634
rect 7656 8570 7708 8576
rect 7760 8566 7788 9658
rect 7748 8560 7800 8566
rect 7748 8502 7800 8508
rect 7656 8492 7708 8498
rect 7656 8434 7708 8440
rect 7668 8401 7696 8434
rect 7654 8392 7710 8401
rect 7654 8327 7710 8336
rect 7378 6352 7434 6361
rect 7378 6287 7434 6296
rect 7392 5914 7420 6287
rect 7380 5908 7432 5914
rect 7380 5850 7432 5856
rect 7104 5704 7156 5710
rect 7104 5646 7156 5652
rect 7116 4078 7144 5646
rect 7288 4616 7340 4622
rect 7288 4558 7340 4564
rect 7300 4282 7328 4558
rect 7288 4276 7340 4282
rect 7288 4218 7340 4224
rect 7300 4146 7328 4218
rect 7392 4146 7420 5850
rect 7484 5846 7512 7278
rect 7576 7262 7696 7290
rect 7564 7200 7616 7206
rect 7564 7142 7616 7148
rect 7472 5840 7524 5846
rect 7472 5782 7524 5788
rect 7576 5370 7604 7142
rect 7668 5710 7696 7262
rect 7852 6730 7880 11086
rect 7944 8634 7972 11194
rect 7932 8628 7984 8634
rect 7932 8570 7984 8576
rect 8220 8276 8248 11194
rect 8392 9036 8444 9042
rect 8392 8978 8444 8984
rect 8404 8498 8432 8978
rect 8496 8634 8524 11194
rect 8666 9752 8722 9761
rect 8666 9687 8722 9696
rect 8576 8832 8628 8838
rect 8576 8774 8628 8780
rect 8484 8628 8536 8634
rect 8484 8570 8536 8576
rect 8392 8492 8444 8498
rect 8392 8434 8444 8440
rect 8484 8424 8536 8430
rect 8484 8366 8536 8372
rect 8220 8248 8340 8276
rect 7950 8188 8258 8197
rect 7950 8186 7956 8188
rect 8012 8186 8036 8188
rect 8092 8186 8116 8188
rect 8172 8186 8196 8188
rect 8252 8186 8258 8188
rect 8012 8134 8014 8186
rect 8194 8134 8196 8186
rect 7950 8132 7956 8134
rect 8012 8132 8036 8134
rect 8092 8132 8116 8134
rect 8172 8132 8196 8134
rect 8252 8132 8258 8134
rect 7950 8123 8258 8132
rect 8312 8090 8340 8248
rect 8300 8084 8352 8090
rect 8300 8026 8352 8032
rect 8208 7948 8260 7954
rect 8208 7890 8260 7896
rect 8220 7313 8248 7890
rect 8300 7880 8352 7886
rect 8300 7822 8352 7828
rect 8206 7304 8262 7313
rect 8206 7239 8262 7248
rect 7950 7100 8258 7109
rect 7950 7098 7956 7100
rect 8012 7098 8036 7100
rect 8092 7098 8116 7100
rect 8172 7098 8196 7100
rect 8252 7098 8258 7100
rect 8012 7046 8014 7098
rect 8194 7046 8196 7098
rect 7950 7044 7956 7046
rect 8012 7044 8036 7046
rect 8092 7044 8116 7046
rect 8172 7044 8196 7046
rect 8252 7044 8258 7046
rect 7950 7035 8258 7044
rect 7840 6724 7892 6730
rect 7840 6666 7892 6672
rect 8312 6458 8340 7822
rect 8390 7168 8446 7177
rect 8390 7103 8446 7112
rect 8300 6452 8352 6458
rect 8300 6394 8352 6400
rect 7748 6112 7800 6118
rect 7748 6054 7800 6060
rect 7656 5704 7708 5710
rect 7656 5646 7708 5652
rect 7564 5364 7616 5370
rect 7564 5306 7616 5312
rect 7564 4616 7616 4622
rect 7564 4558 7616 4564
rect 7576 4146 7604 4558
rect 7288 4140 7340 4146
rect 7288 4082 7340 4088
rect 7380 4140 7432 4146
rect 7380 4082 7432 4088
rect 7564 4140 7616 4146
rect 7564 4082 7616 4088
rect 7760 4078 7788 6054
rect 7950 6012 8258 6021
rect 7950 6010 7956 6012
rect 8012 6010 8036 6012
rect 8092 6010 8116 6012
rect 8172 6010 8196 6012
rect 8252 6010 8258 6012
rect 8012 5958 8014 6010
rect 8194 5958 8196 6010
rect 7950 5956 7956 5958
rect 8012 5956 8036 5958
rect 8092 5956 8116 5958
rect 8172 5956 8196 5958
rect 8252 5956 8258 5958
rect 7950 5947 8258 5956
rect 8404 5409 8432 7103
rect 8496 5914 8524 8366
rect 8588 6882 8616 8774
rect 8680 8498 8708 9687
rect 8668 8492 8720 8498
rect 8668 8434 8720 8440
rect 8772 8090 8800 11194
rect 9048 8922 9076 11194
rect 8864 8894 9076 8922
rect 8864 8634 8892 8894
rect 9324 8820 9352 11194
rect 9496 9784 9548 9790
rect 9496 9726 9548 9732
rect 9324 8792 9444 8820
rect 9010 8732 9318 8741
rect 9010 8730 9016 8732
rect 9072 8730 9096 8732
rect 9152 8730 9176 8732
rect 9232 8730 9256 8732
rect 9312 8730 9318 8732
rect 9072 8678 9074 8730
rect 9254 8678 9256 8730
rect 9010 8676 9016 8678
rect 9072 8676 9096 8678
rect 9152 8676 9176 8678
rect 9232 8676 9256 8678
rect 9312 8676 9318 8678
rect 9010 8667 9318 8676
rect 8852 8628 8904 8634
rect 8852 8570 8904 8576
rect 9416 8090 9444 8792
rect 9508 8498 9536 9726
rect 9600 8634 9628 11194
rect 9772 11076 9824 11082
rect 9772 11018 9824 11024
rect 9678 10160 9734 10169
rect 9678 10095 9734 10104
rect 9588 8628 9640 8634
rect 9588 8570 9640 8576
rect 9496 8492 9548 8498
rect 9496 8434 9548 8440
rect 8760 8084 8812 8090
rect 8760 8026 8812 8032
rect 9404 8084 9456 8090
rect 9404 8026 9456 8032
rect 9692 7886 9720 10095
rect 9220 7880 9272 7886
rect 9218 7848 9220 7857
rect 9680 7880 9732 7886
rect 9272 7848 9274 7857
rect 8852 7812 8904 7818
rect 9680 7822 9732 7828
rect 9218 7783 9274 7792
rect 8852 7754 8904 7760
rect 8588 6854 8708 6882
rect 8576 6792 8628 6798
rect 8576 6734 8628 6740
rect 8484 5908 8536 5914
rect 8484 5850 8536 5856
rect 8588 5794 8616 6734
rect 8680 6458 8708 6854
rect 8760 6724 8812 6730
rect 8760 6666 8812 6672
rect 8668 6452 8720 6458
rect 8668 6394 8720 6400
rect 8668 6316 8720 6322
rect 8668 6258 8720 6264
rect 8496 5766 8616 5794
rect 8390 5400 8446 5409
rect 8390 5335 8446 5344
rect 7950 4924 8258 4933
rect 7950 4922 7956 4924
rect 8012 4922 8036 4924
rect 8092 4922 8116 4924
rect 8172 4922 8196 4924
rect 8252 4922 8258 4924
rect 8012 4870 8014 4922
rect 8194 4870 8196 4922
rect 7950 4868 7956 4870
rect 8012 4868 8036 4870
rect 8092 4868 8116 4870
rect 8172 4868 8196 4870
rect 8252 4868 8258 4870
rect 7950 4859 8258 4868
rect 7104 4072 7156 4078
rect 7104 4014 7156 4020
rect 7748 4072 7800 4078
rect 7748 4014 7800 4020
rect 7950 3836 8258 3845
rect 7950 3834 7956 3836
rect 8012 3834 8036 3836
rect 8092 3834 8116 3836
rect 8172 3834 8196 3836
rect 8252 3834 8258 3836
rect 8012 3782 8014 3834
rect 8194 3782 8196 3834
rect 7950 3780 7956 3782
rect 8012 3780 8036 3782
rect 8092 3780 8116 3782
rect 8172 3780 8196 3782
rect 8252 3780 8258 3782
rect 7950 3771 8258 3780
rect 8496 3534 8524 5766
rect 8576 5704 8628 5710
rect 8576 5646 8628 5652
rect 8588 4146 8616 5646
rect 8680 4282 8708 6258
rect 8772 4622 8800 6666
rect 8864 5914 8892 7754
rect 9010 7644 9318 7653
rect 9010 7642 9016 7644
rect 9072 7642 9096 7644
rect 9152 7642 9176 7644
rect 9232 7642 9256 7644
rect 9312 7642 9318 7644
rect 9072 7590 9074 7642
rect 9254 7590 9256 7642
rect 9010 7588 9016 7590
rect 9072 7588 9096 7590
rect 9152 7588 9176 7590
rect 9232 7588 9256 7590
rect 9312 7588 9318 7590
rect 9010 7579 9318 7588
rect 9680 6996 9732 7002
rect 9680 6938 9732 6944
rect 9404 6724 9456 6730
rect 9404 6666 9456 6672
rect 9010 6556 9318 6565
rect 9010 6554 9016 6556
rect 9072 6554 9096 6556
rect 9152 6554 9176 6556
rect 9232 6554 9256 6556
rect 9312 6554 9318 6556
rect 9072 6502 9074 6554
rect 9254 6502 9256 6554
rect 9010 6500 9016 6502
rect 9072 6500 9096 6502
rect 9152 6500 9176 6502
rect 9232 6500 9256 6502
rect 9312 6500 9318 6502
rect 9010 6491 9318 6500
rect 8944 6452 8996 6458
rect 8944 6394 8996 6400
rect 9128 6452 9180 6458
rect 9128 6394 9180 6400
rect 8956 6322 8984 6394
rect 8944 6316 8996 6322
rect 8944 6258 8996 6264
rect 8852 5908 8904 5914
rect 8852 5850 8904 5856
rect 8956 5522 8984 6258
rect 9140 5710 9168 6394
rect 9220 6248 9272 6254
rect 9220 6190 9272 6196
rect 9232 5846 9260 6190
rect 9220 5840 9272 5846
rect 9220 5782 9272 5788
rect 9128 5704 9180 5710
rect 9128 5646 9180 5652
rect 8864 5494 8984 5522
rect 8864 5302 8892 5494
rect 9010 5468 9318 5477
rect 9010 5466 9016 5468
rect 9072 5466 9096 5468
rect 9152 5466 9176 5468
rect 9232 5466 9256 5468
rect 9312 5466 9318 5468
rect 9072 5414 9074 5466
rect 9254 5414 9256 5466
rect 9010 5412 9016 5414
rect 9072 5412 9096 5414
rect 9152 5412 9176 5414
rect 9232 5412 9256 5414
rect 9312 5412 9318 5414
rect 9010 5403 9318 5412
rect 8852 5296 8904 5302
rect 8852 5238 8904 5244
rect 8760 4616 8812 4622
rect 8760 4558 8812 4564
rect 9010 4380 9318 4389
rect 9010 4378 9016 4380
rect 9072 4378 9096 4380
rect 9152 4378 9176 4380
rect 9232 4378 9256 4380
rect 9312 4378 9318 4380
rect 9072 4326 9074 4378
rect 9254 4326 9256 4378
rect 9010 4324 9016 4326
rect 9072 4324 9096 4326
rect 9152 4324 9176 4326
rect 9232 4324 9256 4326
rect 9312 4324 9318 4326
rect 9010 4315 9318 4324
rect 8668 4276 8720 4282
rect 8668 4218 8720 4224
rect 8576 4140 8628 4146
rect 8576 4082 8628 4088
rect 9416 4010 9444 6666
rect 9588 6656 9640 6662
rect 9588 6598 9640 6604
rect 9496 6248 9548 6254
rect 9496 6190 9548 6196
rect 9404 4004 9456 4010
rect 9404 3946 9456 3952
rect 9508 3738 9536 6190
rect 9600 5250 9628 6598
rect 9692 5710 9720 6938
rect 9784 6866 9812 11018
rect 9876 8634 9904 11194
rect 10048 9852 10100 9858
rect 10048 9794 10100 9800
rect 9864 8628 9916 8634
rect 9864 8570 9916 8576
rect 10060 8498 10088 9794
rect 10152 8634 10180 11194
rect 10324 9580 10376 9586
rect 10324 9522 10376 9528
rect 10230 9480 10286 9489
rect 10230 9415 10286 9424
rect 10140 8628 10192 8634
rect 10140 8570 10192 8576
rect 10244 8498 10272 9415
rect 10048 8492 10100 8498
rect 10048 8434 10100 8440
rect 10232 8492 10284 8498
rect 10232 8434 10284 8440
rect 9864 7744 9916 7750
rect 9864 7686 9916 7692
rect 9876 7002 9904 7686
rect 10140 7540 10192 7546
rect 10140 7482 10192 7488
rect 10152 7342 10180 7482
rect 10140 7336 10192 7342
rect 10140 7278 10192 7284
rect 9864 6996 9916 7002
rect 9864 6938 9916 6944
rect 9772 6860 9824 6866
rect 9772 6802 9824 6808
rect 9864 6792 9916 6798
rect 9864 6734 9916 6740
rect 9680 5704 9732 5710
rect 9680 5646 9732 5652
rect 9600 5222 9720 5250
rect 9588 5160 9640 5166
rect 9586 5128 9588 5137
rect 9640 5128 9642 5137
rect 9586 5063 9642 5072
rect 9692 4978 9720 5222
rect 9600 4950 9720 4978
rect 9600 4146 9628 4950
rect 9876 4826 9904 6734
rect 10048 6656 10100 6662
rect 10048 6598 10100 6604
rect 10060 6322 10088 6598
rect 10048 6316 10100 6322
rect 10048 6258 10100 6264
rect 10048 6112 10100 6118
rect 10048 6054 10100 6060
rect 10060 5710 10088 6054
rect 10152 5710 10180 7278
rect 10336 6798 10364 9522
rect 10428 8090 10456 11194
rect 10600 10056 10652 10062
rect 10600 9998 10652 10004
rect 10612 8498 10640 9998
rect 10704 8634 10732 11194
rect 10876 9920 10928 9926
rect 10876 9862 10928 9868
rect 10692 8628 10744 8634
rect 10692 8570 10744 8576
rect 10888 8498 10916 9862
rect 10980 8634 11008 11194
rect 10968 8628 11020 8634
rect 10968 8570 11020 8576
rect 10600 8492 10652 8498
rect 10600 8434 10652 8440
rect 10876 8492 10928 8498
rect 10876 8434 10928 8440
rect 11256 8090 11284 11194
rect 11532 8634 11560 11194
rect 11520 8628 11572 8634
rect 11520 8570 11572 8576
rect 11612 8560 11664 8566
rect 11612 8502 11664 8508
rect 10416 8084 10468 8090
rect 10416 8026 10468 8032
rect 11244 8084 11296 8090
rect 11244 8026 11296 8032
rect 10784 7880 10836 7886
rect 10784 7822 10836 7828
rect 10796 7449 10824 7822
rect 10782 7440 10838 7449
rect 10782 7375 10838 7384
rect 10324 6792 10376 6798
rect 10244 6740 10324 6746
rect 10244 6734 10376 6740
rect 11428 6792 11480 6798
rect 11428 6734 11480 6740
rect 10244 6718 10364 6734
rect 10048 5704 10100 5710
rect 9954 5672 10010 5681
rect 10048 5646 10100 5652
rect 10140 5704 10192 5710
rect 10140 5646 10192 5652
rect 9954 5607 9956 5616
rect 10008 5607 10010 5616
rect 9956 5578 10008 5584
rect 9864 4820 9916 4826
rect 9864 4762 9916 4768
rect 10244 4146 10272 6718
rect 10322 6216 10378 6225
rect 10322 6151 10378 6160
rect 10336 5778 10364 6151
rect 10324 5772 10376 5778
rect 10324 5714 10376 5720
rect 11440 4622 11468 6734
rect 11624 6662 11652 8502
rect 11808 8090 11836 11194
rect 11980 8628 12032 8634
rect 12084 8616 12112 11194
rect 12360 8634 12388 11194
rect 12440 9104 12492 9110
rect 12440 9046 12492 9052
rect 12032 8588 12112 8616
rect 12348 8628 12400 8634
rect 11980 8570 12032 8576
rect 12348 8570 12400 8576
rect 11980 8356 12032 8362
rect 11980 8298 12032 8304
rect 11796 8084 11848 8090
rect 11796 8026 11848 8032
rect 11888 8016 11940 8022
rect 11888 7958 11940 7964
rect 11612 6656 11664 6662
rect 11612 6598 11664 6604
rect 11900 6458 11928 7958
rect 11992 6458 12020 8298
rect 12164 7880 12216 7886
rect 12164 7822 12216 7828
rect 12176 7546 12204 7822
rect 12164 7540 12216 7546
rect 12164 7482 12216 7488
rect 12256 6928 12308 6934
rect 12256 6870 12308 6876
rect 12268 6798 12296 6870
rect 12256 6792 12308 6798
rect 12256 6734 12308 6740
rect 12164 6724 12216 6730
rect 12164 6666 12216 6672
rect 11888 6452 11940 6458
rect 11888 6394 11940 6400
rect 11980 6452 12032 6458
rect 11980 6394 12032 6400
rect 11520 6316 11572 6322
rect 11520 6258 11572 6264
rect 11428 4616 11480 4622
rect 11428 4558 11480 4564
rect 9588 4140 9640 4146
rect 9588 4082 9640 4088
rect 10232 4140 10284 4146
rect 10232 4082 10284 4088
rect 11336 4140 11388 4146
rect 11336 4082 11388 4088
rect 9496 3732 9548 3738
rect 9496 3674 9548 3680
rect 11348 3602 11376 4082
rect 11532 3602 11560 6258
rect 12176 6254 12204 6666
rect 12164 6248 12216 6254
rect 12164 6190 12216 6196
rect 12256 5092 12308 5098
rect 12256 5034 12308 5040
rect 12268 4826 12296 5034
rect 12256 4820 12308 4826
rect 12256 4762 12308 4768
rect 11612 4616 11664 4622
rect 12072 4616 12124 4622
rect 11612 4558 11664 4564
rect 12070 4584 12072 4593
rect 12164 4616 12216 4622
rect 12124 4584 12126 4593
rect 11624 3602 11652 4558
rect 12164 4558 12216 4564
rect 12070 4519 12126 4528
rect 12176 4486 12204 4558
rect 12164 4480 12216 4486
rect 12452 4468 12480 9046
rect 12532 8832 12584 8838
rect 12532 8774 12584 8780
rect 12544 8566 12572 8774
rect 12532 8560 12584 8566
rect 12532 8502 12584 8508
rect 12636 8090 12664 11194
rect 12912 8362 12940 11194
rect 13188 8634 13216 11194
rect 13358 9344 13414 9353
rect 13358 9279 13414 9288
rect 13176 8628 13228 8634
rect 13176 8570 13228 8576
rect 12990 8528 13046 8537
rect 13372 8498 13400 9279
rect 12990 8463 12992 8472
rect 13044 8463 13046 8472
rect 13360 8492 13412 8498
rect 12992 8434 13044 8440
rect 13360 8434 13412 8440
rect 12900 8356 12952 8362
rect 12900 8298 12952 8304
rect 12808 8288 12860 8294
rect 12808 8230 12860 8236
rect 12624 8084 12676 8090
rect 12624 8026 12676 8032
rect 12820 7274 12848 8230
rect 13464 8090 13492 11194
rect 13544 8424 13596 8430
rect 13544 8366 13596 8372
rect 13452 8084 13504 8090
rect 13452 8026 13504 8032
rect 13176 7948 13228 7954
rect 13176 7890 13228 7896
rect 13084 7404 13136 7410
rect 13084 7346 13136 7352
rect 12808 7268 12860 7274
rect 12808 7210 12860 7216
rect 12716 7200 12768 7206
rect 12716 7142 12768 7148
rect 12532 6316 12584 6322
rect 12532 6258 12584 6264
rect 12544 6118 12572 6258
rect 12532 6112 12584 6118
rect 12532 6054 12584 6060
rect 12728 4690 12756 7142
rect 12820 5778 12848 7210
rect 12992 6792 13044 6798
rect 12992 6734 13044 6740
rect 12808 5772 12860 5778
rect 12808 5714 12860 5720
rect 12716 4684 12768 4690
rect 12716 4626 12768 4632
rect 12532 4480 12584 4486
rect 12452 4440 12532 4468
rect 12164 4422 12216 4428
rect 12532 4422 12584 4428
rect 12728 4078 12756 4626
rect 12716 4072 12768 4078
rect 12716 4014 12768 4020
rect 13004 3602 13032 6734
rect 13096 5710 13124 7346
rect 13084 5704 13136 5710
rect 13084 5646 13136 5652
rect 13188 4554 13216 7890
rect 13360 7744 13412 7750
rect 13360 7686 13412 7692
rect 13372 7478 13400 7686
rect 13450 7576 13506 7585
rect 13450 7511 13506 7520
rect 13360 7472 13412 7478
rect 13360 7414 13412 7420
rect 13464 7313 13492 7511
rect 13450 7304 13506 7313
rect 13450 7239 13506 7248
rect 13268 6452 13320 6458
rect 13268 6394 13320 6400
rect 13280 5846 13308 6394
rect 13268 5840 13320 5846
rect 13360 5840 13412 5846
rect 13268 5782 13320 5788
rect 13358 5808 13360 5817
rect 13412 5808 13414 5817
rect 13358 5743 13414 5752
rect 13268 5704 13320 5710
rect 13268 5646 13320 5652
rect 13280 5302 13308 5646
rect 13268 5296 13320 5302
rect 13268 5238 13320 5244
rect 13360 5160 13412 5166
rect 13360 5102 13412 5108
rect 13372 4826 13400 5102
rect 13556 4826 13584 8366
rect 13740 8362 13768 11194
rect 13820 9104 13872 9110
rect 13820 9046 13872 9052
rect 13728 8356 13780 8362
rect 13728 8298 13780 8304
rect 13832 7970 13860 9046
rect 14016 8634 14044 11194
rect 14004 8628 14056 8634
rect 14004 8570 14056 8576
rect 13950 8188 14258 8197
rect 13950 8186 13956 8188
rect 14012 8186 14036 8188
rect 14092 8186 14116 8188
rect 14172 8186 14196 8188
rect 14252 8186 14258 8188
rect 14012 8134 14014 8186
rect 14194 8134 14196 8186
rect 13950 8132 13956 8134
rect 14012 8132 14036 8134
rect 14092 8132 14116 8134
rect 14172 8132 14196 8134
rect 14252 8132 14258 8134
rect 13950 8123 14258 8132
rect 14292 8090 14320 11194
rect 14464 9512 14516 9518
rect 14464 9454 14516 9460
rect 14280 8084 14332 8090
rect 14280 8026 14332 8032
rect 13832 7942 13952 7970
rect 13820 7880 13872 7886
rect 13820 7822 13872 7828
rect 13728 7812 13780 7818
rect 13728 7754 13780 7760
rect 13740 7002 13768 7754
rect 13832 7478 13860 7822
rect 13820 7472 13872 7478
rect 13820 7414 13872 7420
rect 13924 7290 13952 7942
rect 14186 7576 14242 7585
rect 14186 7511 14242 7520
rect 14200 7410 14228 7511
rect 14278 7440 14334 7449
rect 14188 7404 14240 7410
rect 14334 7398 14412 7426
rect 14278 7375 14334 7384
rect 14188 7346 14240 7352
rect 13832 7262 13952 7290
rect 13728 6996 13780 7002
rect 13728 6938 13780 6944
rect 13832 6798 13860 7262
rect 13950 7100 14258 7109
rect 13950 7098 13956 7100
rect 14012 7098 14036 7100
rect 14092 7098 14116 7100
rect 14172 7098 14196 7100
rect 14252 7098 14258 7100
rect 14012 7046 14014 7098
rect 14194 7046 14196 7098
rect 13950 7044 13956 7046
rect 14012 7044 14036 7046
rect 14092 7044 14116 7046
rect 14172 7044 14196 7046
rect 14252 7044 14258 7046
rect 13950 7035 14258 7044
rect 14384 7041 14412 7398
rect 14476 7206 14504 9454
rect 14568 8634 14596 11194
rect 14648 9988 14700 9994
rect 14648 9930 14700 9936
rect 14556 8628 14608 8634
rect 14556 8570 14608 8576
rect 14660 8498 14688 9930
rect 14738 9888 14794 9897
rect 14738 9823 14794 9832
rect 14752 8838 14780 9823
rect 14740 8832 14792 8838
rect 14740 8774 14792 8780
rect 14740 8560 14792 8566
rect 14740 8502 14792 8508
rect 14648 8492 14700 8498
rect 14648 8434 14700 8440
rect 14556 8288 14608 8294
rect 14556 8230 14608 8236
rect 14568 7750 14596 8230
rect 14648 7880 14700 7886
rect 14646 7848 14648 7857
rect 14700 7848 14702 7857
rect 14646 7783 14702 7792
rect 14556 7744 14608 7750
rect 14556 7686 14608 7692
rect 14648 7744 14700 7750
rect 14648 7686 14700 7692
rect 14464 7200 14516 7206
rect 14464 7142 14516 7148
rect 14370 7032 14426 7041
rect 14370 6967 14426 6976
rect 13820 6792 13872 6798
rect 13820 6734 13872 6740
rect 14370 6760 14426 6769
rect 14370 6695 14426 6704
rect 13820 6656 13872 6662
rect 13820 6598 13872 6604
rect 14188 6656 14240 6662
rect 14188 6598 14240 6604
rect 13728 6112 13780 6118
rect 13728 6054 13780 6060
rect 13740 5778 13768 6054
rect 13728 5772 13780 5778
rect 13728 5714 13780 5720
rect 13728 5636 13780 5642
rect 13648 5596 13728 5624
rect 13360 4820 13412 4826
rect 13360 4762 13412 4768
rect 13544 4820 13596 4826
rect 13544 4762 13596 4768
rect 13176 4548 13228 4554
rect 13176 4490 13228 4496
rect 13648 3738 13676 5596
rect 13728 5578 13780 5584
rect 13832 4690 13860 6598
rect 14094 6488 14150 6497
rect 14094 6423 14150 6432
rect 14108 6322 14136 6423
rect 14096 6316 14148 6322
rect 14096 6258 14148 6264
rect 14200 6254 14228 6598
rect 14188 6248 14240 6254
rect 14188 6190 14240 6196
rect 14280 6248 14332 6254
rect 14280 6190 14332 6196
rect 13950 6012 14258 6021
rect 13950 6010 13956 6012
rect 14012 6010 14036 6012
rect 14092 6010 14116 6012
rect 14172 6010 14196 6012
rect 14252 6010 14258 6012
rect 14012 5958 14014 6010
rect 14194 5958 14196 6010
rect 13950 5956 13956 5958
rect 14012 5956 14036 5958
rect 14092 5956 14116 5958
rect 14172 5956 14196 5958
rect 14252 5956 14258 5958
rect 13950 5947 14258 5956
rect 14096 5908 14148 5914
rect 14292 5896 14320 6190
rect 14384 5914 14412 6695
rect 14148 5868 14320 5896
rect 14096 5850 14148 5856
rect 14292 5234 14320 5868
rect 14372 5908 14424 5914
rect 14372 5850 14424 5856
rect 14372 5704 14424 5710
rect 14372 5646 14424 5652
rect 14280 5228 14332 5234
rect 14280 5170 14332 5176
rect 13950 4924 14258 4933
rect 13950 4922 13956 4924
rect 14012 4922 14036 4924
rect 14092 4922 14116 4924
rect 14172 4922 14196 4924
rect 14252 4922 14258 4924
rect 14012 4870 14014 4922
rect 14194 4870 14196 4922
rect 13950 4868 13956 4870
rect 14012 4868 14036 4870
rect 14092 4868 14116 4870
rect 14172 4868 14196 4870
rect 14252 4868 14258 4870
rect 13950 4859 14258 4868
rect 14280 4820 14332 4826
rect 14280 4762 14332 4768
rect 13820 4684 13872 4690
rect 13820 4626 13872 4632
rect 13728 4616 13780 4622
rect 13728 4558 13780 4564
rect 13636 3732 13688 3738
rect 13636 3674 13688 3680
rect 13740 3670 13768 4558
rect 14292 4554 14320 4762
rect 14280 4548 14332 4554
rect 14280 4490 14332 4496
rect 13950 3836 14258 3845
rect 13950 3834 13956 3836
rect 14012 3834 14036 3836
rect 14092 3834 14116 3836
rect 14172 3834 14196 3836
rect 14252 3834 14258 3836
rect 14012 3782 14014 3834
rect 14194 3782 14196 3834
rect 13950 3780 13956 3782
rect 14012 3780 14036 3782
rect 14092 3780 14116 3782
rect 14172 3780 14196 3782
rect 14252 3780 14258 3782
rect 13950 3771 14258 3780
rect 14384 3738 14412 5646
rect 14476 4622 14504 7142
rect 14660 6390 14688 7686
rect 14752 7177 14780 8502
rect 14844 8090 14872 11194
rect 15120 8922 15148 11194
rect 14936 8894 15148 8922
rect 14936 8634 14964 8894
rect 15010 8732 15318 8741
rect 15010 8730 15016 8732
rect 15072 8730 15096 8732
rect 15152 8730 15176 8732
rect 15232 8730 15256 8732
rect 15312 8730 15318 8732
rect 15072 8678 15074 8730
rect 15254 8678 15256 8730
rect 15010 8676 15016 8678
rect 15072 8676 15096 8678
rect 15152 8676 15176 8678
rect 15232 8676 15256 8678
rect 15312 8676 15318 8678
rect 15010 8667 15318 8676
rect 15396 8634 15424 11194
rect 15568 9648 15620 9654
rect 15568 9590 15620 9596
rect 15476 9376 15528 9382
rect 15476 9318 15528 9324
rect 14924 8628 14976 8634
rect 14924 8570 14976 8576
rect 15384 8628 15436 8634
rect 15384 8570 15436 8576
rect 15488 8514 15516 9318
rect 15396 8498 15516 8514
rect 15384 8492 15516 8498
rect 15436 8486 15516 8492
rect 15384 8434 15436 8440
rect 15108 8424 15160 8430
rect 15108 8366 15160 8372
rect 14922 8256 14978 8265
rect 14922 8191 14978 8200
rect 14832 8084 14884 8090
rect 14832 8026 14884 8032
rect 14738 7168 14794 7177
rect 14738 7103 14794 7112
rect 14648 6384 14700 6390
rect 14648 6326 14700 6332
rect 14556 6316 14608 6322
rect 14556 6258 14608 6264
rect 14740 6316 14792 6322
rect 14740 6258 14792 6264
rect 14568 4622 14596 6258
rect 14648 6112 14700 6118
rect 14648 6054 14700 6060
rect 14660 5710 14688 6054
rect 14648 5704 14700 5710
rect 14648 5646 14700 5652
rect 14464 4616 14516 4622
rect 14464 4558 14516 4564
rect 14556 4616 14608 4622
rect 14556 4558 14608 4564
rect 14568 4146 14596 4558
rect 14556 4140 14608 4146
rect 14556 4082 14608 4088
rect 14752 4010 14780 6258
rect 14832 5908 14884 5914
rect 14832 5850 14884 5856
rect 14740 4004 14792 4010
rect 14740 3946 14792 3952
rect 14462 3904 14518 3913
rect 14462 3839 14518 3848
rect 14372 3732 14424 3738
rect 14372 3674 14424 3680
rect 13728 3664 13780 3670
rect 13728 3606 13780 3612
rect 11336 3596 11388 3602
rect 11336 3538 11388 3544
rect 11520 3596 11572 3602
rect 11520 3538 11572 3544
rect 11612 3596 11664 3602
rect 11612 3538 11664 3544
rect 12992 3596 13044 3602
rect 12992 3538 13044 3544
rect 8484 3528 8536 3534
rect 8484 3470 8536 3476
rect 9010 3292 9318 3301
rect 9010 3290 9016 3292
rect 9072 3290 9096 3292
rect 9152 3290 9176 3292
rect 9232 3290 9256 3292
rect 9312 3290 9318 3292
rect 9072 3238 9074 3290
rect 9254 3238 9256 3290
rect 9010 3236 9016 3238
rect 9072 3236 9096 3238
rect 9152 3236 9176 3238
rect 9232 3236 9256 3238
rect 9312 3236 9318 3238
rect 9010 3227 9318 3236
rect 7012 3120 7064 3126
rect 7012 3062 7064 3068
rect 13740 2922 13768 3606
rect 14476 3534 14504 3839
rect 14464 3528 14516 3534
rect 14464 3470 14516 3476
rect 13728 2916 13780 2922
rect 13728 2858 13780 2864
rect 9864 2848 9916 2854
rect 9864 2790 9916 2796
rect 7950 2748 8258 2757
rect 7950 2746 7956 2748
rect 8012 2746 8036 2748
rect 8092 2746 8116 2748
rect 8172 2746 8196 2748
rect 8252 2746 8258 2748
rect 8012 2694 8014 2746
rect 8194 2694 8196 2746
rect 7950 2692 7956 2694
rect 8012 2692 8036 2694
rect 8092 2692 8116 2694
rect 8172 2692 8196 2694
rect 8252 2692 8258 2694
rect 7950 2683 8258 2692
rect 6920 2644 6972 2650
rect 6920 2586 6972 2592
rect 9876 2446 9904 2790
rect 13950 2748 14258 2757
rect 13950 2746 13956 2748
rect 14012 2746 14036 2748
rect 14092 2746 14116 2748
rect 14172 2746 14196 2748
rect 14252 2746 14258 2748
rect 14012 2694 14014 2746
rect 14194 2694 14196 2746
rect 13950 2692 13956 2694
rect 14012 2692 14036 2694
rect 14092 2692 14116 2694
rect 14172 2692 14196 2694
rect 14252 2692 14258 2694
rect 13950 2683 14258 2692
rect 12622 2544 12678 2553
rect 14844 2514 14872 5850
rect 14936 5574 14964 8191
rect 15120 7732 15148 8366
rect 15120 7721 15516 7732
rect 15120 7712 15530 7721
rect 15120 7704 15474 7712
rect 15010 7644 15318 7653
rect 15474 7647 15530 7656
rect 15010 7642 15016 7644
rect 15072 7642 15096 7644
rect 15152 7642 15176 7644
rect 15232 7642 15256 7644
rect 15312 7642 15318 7644
rect 15072 7590 15074 7642
rect 15254 7590 15256 7642
rect 15010 7588 15016 7590
rect 15072 7588 15096 7590
rect 15152 7588 15176 7590
rect 15232 7588 15256 7590
rect 15312 7588 15318 7590
rect 15010 7579 15318 7588
rect 15474 7576 15530 7585
rect 15474 7511 15530 7520
rect 15488 7410 15516 7511
rect 15476 7404 15528 7410
rect 15476 7346 15528 7352
rect 15108 7336 15160 7342
rect 15108 7278 15160 7284
rect 15580 7290 15608 9590
rect 15672 8634 15700 11194
rect 15752 8900 15804 8906
rect 15752 8842 15804 8848
rect 15660 8628 15712 8634
rect 15660 8570 15712 8576
rect 15120 6866 15148 7278
rect 15580 7262 15700 7290
rect 15384 7200 15436 7206
rect 15384 7142 15436 7148
rect 15568 7200 15620 7206
rect 15568 7142 15620 7148
rect 15108 6860 15160 6866
rect 15108 6802 15160 6808
rect 15120 6730 15148 6802
rect 15396 6798 15424 7142
rect 15384 6792 15436 6798
rect 15384 6734 15436 6740
rect 15108 6724 15160 6730
rect 15108 6666 15160 6672
rect 15476 6656 15528 6662
rect 15476 6598 15528 6604
rect 15010 6556 15318 6565
rect 15010 6554 15016 6556
rect 15072 6554 15096 6556
rect 15152 6554 15176 6556
rect 15232 6554 15256 6556
rect 15312 6554 15318 6556
rect 15072 6502 15074 6554
rect 15254 6502 15256 6554
rect 15010 6500 15016 6502
rect 15072 6500 15096 6502
rect 15152 6500 15176 6502
rect 15232 6500 15256 6502
rect 15312 6500 15318 6502
rect 15010 6491 15318 6500
rect 15384 6384 15436 6390
rect 15384 6326 15436 6332
rect 14924 5568 14976 5574
rect 14924 5510 14976 5516
rect 15010 5468 15318 5477
rect 15010 5466 15016 5468
rect 15072 5466 15096 5468
rect 15152 5466 15176 5468
rect 15232 5466 15256 5468
rect 15312 5466 15318 5468
rect 15072 5414 15074 5466
rect 15254 5414 15256 5466
rect 15010 5412 15016 5414
rect 15072 5412 15096 5414
rect 15152 5412 15176 5414
rect 15232 5412 15256 5414
rect 15312 5412 15318 5414
rect 15010 5403 15318 5412
rect 15292 5364 15344 5370
rect 15292 5306 15344 5312
rect 15304 5234 15332 5306
rect 15292 5228 15344 5234
rect 15292 5170 15344 5176
rect 15292 5024 15344 5030
rect 15292 4966 15344 4972
rect 15304 4690 15332 4966
rect 15292 4684 15344 4690
rect 15292 4626 15344 4632
rect 15010 4380 15318 4389
rect 15010 4378 15016 4380
rect 15072 4378 15096 4380
rect 15152 4378 15176 4380
rect 15232 4378 15256 4380
rect 15312 4378 15318 4380
rect 15072 4326 15074 4378
rect 15254 4326 15256 4378
rect 15010 4324 15016 4326
rect 15072 4324 15096 4326
rect 15152 4324 15176 4326
rect 15232 4324 15256 4326
rect 15312 4324 15318 4326
rect 15010 4315 15318 4324
rect 15396 3738 15424 6326
rect 15488 4298 15516 6598
rect 15580 5098 15608 7142
rect 15672 5914 15700 7262
rect 15764 6458 15792 8842
rect 15844 8492 15896 8498
rect 15844 8434 15896 8440
rect 15856 7206 15884 8434
rect 15948 8090 15976 11194
rect 16028 9444 16080 9450
rect 16028 9386 16080 9392
rect 15936 8084 15988 8090
rect 15936 8026 15988 8032
rect 15844 7200 15896 7206
rect 15844 7142 15896 7148
rect 15844 6792 15896 6798
rect 15844 6734 15896 6740
rect 15752 6452 15804 6458
rect 15752 6394 15804 6400
rect 15856 6186 15884 6734
rect 16040 6662 16068 9386
rect 16224 8634 16252 11194
rect 16394 9072 16450 9081
rect 16394 9007 16450 9016
rect 16408 8974 16436 9007
rect 16396 8968 16448 8974
rect 16396 8910 16448 8916
rect 16500 8634 16528 11194
rect 16672 9512 16724 9518
rect 16672 9454 16724 9460
rect 16580 9036 16632 9042
rect 16580 8978 16632 8984
rect 16212 8628 16264 8634
rect 16212 8570 16264 8576
rect 16488 8628 16540 8634
rect 16488 8570 16540 8576
rect 16120 8492 16172 8498
rect 16120 8434 16172 8440
rect 16028 6656 16080 6662
rect 16028 6598 16080 6604
rect 16028 6316 16080 6322
rect 16028 6258 16080 6264
rect 15844 6180 15896 6186
rect 15844 6122 15896 6128
rect 15660 5908 15712 5914
rect 15660 5850 15712 5856
rect 15660 5704 15712 5710
rect 15660 5646 15712 5652
rect 15568 5092 15620 5098
rect 15568 5034 15620 5040
rect 15488 4270 15608 4298
rect 15580 4146 15608 4270
rect 15568 4140 15620 4146
rect 15568 4082 15620 4088
rect 15476 4072 15528 4078
rect 15476 4014 15528 4020
rect 15384 3732 15436 3738
rect 15384 3674 15436 3680
rect 15488 3534 15516 4014
rect 15672 3534 15700 5646
rect 15750 5536 15806 5545
rect 15750 5471 15806 5480
rect 15764 5302 15792 5471
rect 15752 5296 15804 5302
rect 15752 5238 15804 5244
rect 16040 4826 16068 6258
rect 16132 5098 16160 8434
rect 16212 7948 16264 7954
rect 16212 7890 16264 7896
rect 16224 7750 16252 7890
rect 16212 7744 16264 7750
rect 16212 7686 16264 7692
rect 16488 6928 16540 6934
rect 16488 6870 16540 6876
rect 16304 6860 16356 6866
rect 16304 6802 16356 6808
rect 16212 6656 16264 6662
rect 16212 6598 16264 6604
rect 16224 6322 16252 6598
rect 16212 6316 16264 6322
rect 16212 6258 16264 6264
rect 16120 5092 16172 5098
rect 16120 5034 16172 5040
rect 16028 4820 16080 4826
rect 16028 4762 16080 4768
rect 15476 3528 15528 3534
rect 15476 3470 15528 3476
rect 15660 3528 15712 3534
rect 15660 3470 15712 3476
rect 16316 3398 16344 6802
rect 16396 6112 16448 6118
rect 16396 6054 16448 6060
rect 16408 4622 16436 6054
rect 16396 4616 16448 4622
rect 16500 4604 16528 6870
rect 16592 5030 16620 8978
rect 16684 8498 16712 9454
rect 16776 8634 16804 11194
rect 16764 8628 16816 8634
rect 16764 8570 16816 8576
rect 16672 8492 16724 8498
rect 16672 8434 16724 8440
rect 16856 8492 16908 8498
rect 16856 8434 16908 8440
rect 16868 8022 16896 8434
rect 17052 8362 17080 11194
rect 17132 9716 17184 9722
rect 17132 9658 17184 9664
rect 17040 8356 17092 8362
rect 17040 8298 17092 8304
rect 16856 8016 16908 8022
rect 16856 7958 16908 7964
rect 16670 6488 16726 6497
rect 16670 6423 16726 6432
rect 16684 5710 16712 6423
rect 17144 5846 17172 9658
rect 17224 9036 17276 9042
rect 17224 8978 17276 8984
rect 17236 8566 17264 8978
rect 17328 8634 17356 11194
rect 17500 9308 17552 9314
rect 17500 9250 17552 9256
rect 17316 8628 17368 8634
rect 17316 8570 17368 8576
rect 17224 8560 17276 8566
rect 17224 8502 17276 8508
rect 17408 8492 17460 8498
rect 17408 8434 17460 8440
rect 17420 5914 17448 8434
rect 17512 5914 17540 9250
rect 17604 8090 17632 11194
rect 17684 8424 17736 8430
rect 17684 8366 17736 8372
rect 17592 8084 17644 8090
rect 17592 8026 17644 8032
rect 17696 6882 17724 8366
rect 17880 7886 17908 11194
rect 17960 9104 18012 9110
rect 17960 9046 18012 9052
rect 17868 7880 17920 7886
rect 17868 7822 17920 7828
rect 17776 7200 17828 7206
rect 17776 7142 17828 7148
rect 17604 6854 17724 6882
rect 17408 5908 17460 5914
rect 17408 5850 17460 5856
rect 17500 5908 17552 5914
rect 17500 5850 17552 5856
rect 17132 5840 17184 5846
rect 17132 5782 17184 5788
rect 17604 5710 17632 6854
rect 17684 6724 17736 6730
rect 17684 6666 17736 6672
rect 17696 6322 17724 6666
rect 17684 6316 17736 6322
rect 17684 6258 17736 6264
rect 17684 6112 17736 6118
rect 17684 6054 17736 6060
rect 17696 5914 17724 6054
rect 17684 5908 17736 5914
rect 17684 5850 17736 5856
rect 16672 5704 16724 5710
rect 16672 5646 16724 5652
rect 16764 5704 16816 5710
rect 16764 5646 16816 5652
rect 17592 5704 17644 5710
rect 17592 5646 17644 5652
rect 16580 5024 16632 5030
rect 16580 4966 16632 4972
rect 16672 4616 16724 4622
rect 16500 4576 16672 4604
rect 16396 4558 16448 4564
rect 16672 4558 16724 4564
rect 16684 4078 16712 4558
rect 16672 4072 16724 4078
rect 16672 4014 16724 4020
rect 16578 3768 16634 3777
rect 16578 3703 16634 3712
rect 16592 3602 16620 3703
rect 16776 3602 16804 5646
rect 17040 5228 17092 5234
rect 17040 5170 17092 5176
rect 17052 4826 17080 5170
rect 17040 4820 17092 4826
rect 17040 4762 17092 4768
rect 17498 4720 17554 4729
rect 17498 4655 17554 4664
rect 16580 3596 16632 3602
rect 16580 3538 16632 3544
rect 16764 3596 16816 3602
rect 16764 3538 16816 3544
rect 17130 3496 17186 3505
rect 17130 3431 17186 3440
rect 16304 3392 16356 3398
rect 16304 3334 16356 3340
rect 15010 3292 15318 3301
rect 15010 3290 15016 3292
rect 15072 3290 15096 3292
rect 15152 3290 15176 3292
rect 15232 3290 15256 3292
rect 15312 3290 15318 3292
rect 15072 3238 15074 3290
rect 15254 3238 15256 3290
rect 15010 3236 15016 3238
rect 15072 3236 15096 3238
rect 15152 3236 15176 3238
rect 15232 3236 15256 3238
rect 15312 3236 15318 3238
rect 15010 3227 15318 3236
rect 15200 3188 15252 3194
rect 15200 3130 15252 3136
rect 15212 2514 15240 3130
rect 17144 3097 17172 3431
rect 17130 3088 17186 3097
rect 17130 3023 17186 3032
rect 17314 3088 17370 3097
rect 17314 3023 17370 3032
rect 12622 2479 12678 2488
rect 14832 2508 14884 2514
rect 6736 2440 6788 2446
rect 6736 2382 6788 2388
rect 9496 2440 9548 2446
rect 9496 2382 9548 2388
rect 9864 2440 9916 2446
rect 9864 2382 9916 2388
rect 5540 2372 5592 2378
rect 5540 2314 5592 2320
rect 4804 2304 4856 2310
rect 4804 2246 4856 2252
rect 6368 2304 6420 2310
rect 6368 2246 6420 2252
rect 4712 2032 4764 2038
rect 4712 1974 4764 1980
rect 4816 56 4844 2246
rect 6380 56 6408 2246
rect 6748 2106 6776 2382
rect 9010 2204 9318 2213
rect 9010 2202 9016 2204
rect 9072 2202 9096 2204
rect 9152 2202 9176 2204
rect 9232 2202 9256 2204
rect 9312 2202 9318 2204
rect 9072 2150 9074 2202
rect 9254 2150 9256 2202
rect 9010 2148 9016 2150
rect 9072 2148 9096 2150
rect 9152 2148 9176 2150
rect 9232 2148 9256 2150
rect 9312 2148 9318 2150
rect 9010 2139 9318 2148
rect 6736 2100 6788 2106
rect 6736 2042 6788 2048
rect 7944 66 8064 82
rect 7944 60 8076 66
rect 7944 56 8024 60
rect 3344 14 3464 42
rect 4802 0 4858 56
rect 6366 0 6422 56
rect 7930 54 8024 56
rect 7930 0 7986 54
rect 9508 56 9536 2382
rect 11058 1864 11114 1873
rect 11058 1799 11114 1808
rect 11072 56 11100 1799
rect 12636 56 12664 2479
rect 14832 2450 14884 2456
rect 15200 2508 15252 2514
rect 15200 2450 15252 2456
rect 15010 2204 15318 2213
rect 15010 2202 15016 2204
rect 15072 2202 15096 2204
rect 15152 2202 15176 2204
rect 15232 2202 15256 2204
rect 15312 2202 15318 2204
rect 15072 2150 15074 2202
rect 15254 2150 15256 2202
rect 15010 2148 15016 2150
rect 15072 2148 15096 2150
rect 15152 2148 15176 2150
rect 15232 2148 15256 2150
rect 15312 2148 15318 2150
rect 15010 2139 15318 2148
rect 14188 196 14240 202
rect 14188 138 14240 144
rect 14200 56 14228 138
rect 15750 96 15806 105
rect 8024 2 8076 8
rect 9494 0 9550 56
rect 11058 0 11114 56
rect 12622 0 12678 56
rect 14186 0 14242 56
rect 17328 56 17356 3023
rect 17512 2106 17540 4655
rect 17604 4622 17632 5646
rect 17684 5228 17736 5234
rect 17684 5170 17736 5176
rect 17592 4616 17644 4622
rect 17592 4558 17644 4564
rect 17696 3670 17724 5170
rect 17684 3664 17736 3670
rect 17684 3606 17736 3612
rect 17788 3602 17816 7142
rect 17972 6322 18000 9046
rect 18052 8492 18104 8498
rect 18052 8434 18104 8440
rect 18064 8265 18092 8434
rect 18050 8256 18106 8265
rect 18050 8191 18106 8200
rect 18052 8084 18104 8090
rect 18052 8026 18104 8032
rect 17960 6316 18012 6322
rect 17960 6258 18012 6264
rect 17868 6112 17920 6118
rect 17868 6054 17920 6060
rect 17880 5302 17908 6054
rect 17868 5296 17920 5302
rect 17868 5238 17920 5244
rect 17972 4298 18000 6258
rect 17880 4270 18000 4298
rect 18064 4282 18092 8026
rect 18156 7886 18184 11194
rect 18432 8498 18460 11194
rect 18708 8498 18736 11194
rect 18788 8968 18840 8974
rect 18788 8910 18840 8916
rect 18800 8634 18828 8910
rect 18788 8628 18840 8634
rect 18788 8570 18840 8576
rect 18984 8498 19012 11194
rect 19154 10024 19210 10033
rect 19154 9959 19210 9968
rect 19064 9308 19116 9314
rect 19064 9250 19116 9256
rect 18420 8492 18472 8498
rect 18420 8434 18472 8440
rect 18696 8492 18748 8498
rect 18696 8434 18748 8440
rect 18972 8492 19024 8498
rect 18972 8434 19024 8440
rect 18144 7880 18196 7886
rect 18144 7822 18196 7828
rect 18236 7744 18288 7750
rect 18236 7686 18288 7692
rect 18880 7744 18932 7750
rect 18880 7686 18932 7692
rect 18248 7002 18276 7686
rect 18510 7168 18566 7177
rect 18510 7103 18566 7112
rect 18236 6996 18288 7002
rect 18236 6938 18288 6944
rect 18328 6996 18380 7002
rect 18328 6938 18380 6944
rect 18340 4486 18368 6938
rect 18524 5914 18552 7103
rect 18512 5908 18564 5914
rect 18512 5850 18564 5856
rect 18696 5704 18748 5710
rect 18696 5646 18748 5652
rect 18328 4480 18380 4486
rect 18328 4422 18380 4428
rect 18052 4276 18104 4282
rect 17880 4010 17908 4270
rect 18052 4218 18104 4224
rect 18052 4140 18104 4146
rect 18052 4082 18104 4088
rect 18144 4140 18196 4146
rect 18144 4082 18196 4088
rect 17868 4004 17920 4010
rect 17868 3946 17920 3952
rect 18064 3777 18092 4082
rect 18050 3768 18106 3777
rect 18156 3738 18184 4082
rect 18050 3703 18106 3712
rect 18144 3732 18196 3738
rect 17776 3596 17828 3602
rect 17776 3538 17828 3544
rect 18064 3534 18092 3703
rect 18144 3674 18196 3680
rect 18052 3528 18104 3534
rect 18052 3470 18104 3476
rect 18708 3398 18736 5646
rect 18892 4146 18920 7686
rect 19076 6610 19104 9250
rect 18984 6582 19104 6610
rect 18984 6186 19012 6582
rect 19168 6304 19196 9959
rect 19260 8498 19288 11194
rect 19340 9580 19392 9586
rect 19340 9522 19392 9528
rect 19352 8634 19380 9522
rect 19536 8634 19564 11194
rect 19708 8832 19760 8838
rect 19708 8774 19760 8780
rect 19340 8628 19392 8634
rect 19340 8570 19392 8576
rect 19524 8628 19576 8634
rect 19524 8570 19576 8576
rect 19616 8628 19668 8634
rect 19616 8570 19668 8576
rect 19248 8492 19300 8498
rect 19248 8434 19300 8440
rect 19524 7880 19576 7886
rect 19524 7822 19576 7828
rect 19340 7540 19392 7546
rect 19340 7482 19392 7488
rect 19248 7404 19300 7410
rect 19248 7346 19300 7352
rect 19260 7206 19288 7346
rect 19248 7200 19300 7206
rect 19248 7142 19300 7148
rect 19352 6662 19380 7482
rect 19536 7041 19564 7822
rect 19522 7032 19578 7041
rect 19522 6967 19578 6976
rect 19340 6656 19392 6662
rect 19340 6598 19392 6604
rect 19628 6497 19656 8570
rect 19614 6488 19670 6497
rect 19614 6423 19670 6432
rect 19248 6316 19300 6322
rect 19168 6276 19248 6304
rect 19248 6258 19300 6264
rect 19616 6316 19668 6322
rect 19616 6258 19668 6264
rect 19432 6248 19484 6254
rect 19352 6208 19432 6236
rect 18972 6180 19024 6186
rect 18972 6122 19024 6128
rect 19248 5160 19300 5166
rect 19352 5148 19380 6208
rect 19432 6190 19484 6196
rect 19628 5914 19656 6258
rect 19616 5908 19668 5914
rect 19616 5850 19668 5856
rect 19720 5710 19748 8774
rect 19812 8480 19840 11194
rect 20128 11194 20130 11212
rect 20350 11194 20406 11250
rect 20626 11194 20682 11250
rect 20902 11194 20958 11250
rect 21178 11194 21234 11250
rect 21454 11194 21510 11250
rect 21730 11194 21786 11250
rect 22006 11194 22062 11250
rect 22282 11194 22338 11250
rect 22558 11194 22614 11250
rect 22834 11194 22890 11250
rect 23110 11194 23166 11250
rect 23386 11194 23442 11250
rect 23662 11194 23718 11250
rect 23938 11194 23994 11250
rect 24214 11194 24270 11250
rect 24490 11194 24546 11250
rect 24766 11194 24822 11250
rect 25042 11194 25098 11250
rect 25318 11194 25374 11250
rect 25594 11194 25650 11250
rect 25870 11194 25926 11250
rect 26146 11194 26202 11250
rect 26422 11194 26478 11250
rect 26698 11194 26754 11250
rect 26974 11194 27030 11250
rect 27250 11194 27306 11250
rect 27526 11194 27582 11250
rect 27802 11194 27858 11250
rect 28078 11194 28134 11250
rect 28354 11194 28410 11250
rect 28630 11194 28686 11250
rect 28906 11194 28962 11250
rect 29182 11194 29238 11250
rect 29458 11194 29514 11250
rect 29734 11194 29790 11250
rect 30010 11194 30066 11250
rect 30286 11194 30342 11250
rect 30562 11194 30618 11250
rect 30838 11194 30894 11250
rect 31114 11194 31170 11250
rect 31390 11194 31446 11250
rect 31666 11194 31722 11250
rect 31942 11194 31998 11250
rect 32218 11194 32274 11250
rect 32494 11194 32550 11250
rect 32770 11194 32826 11250
rect 33046 11194 33102 11250
rect 33322 11194 33378 11250
rect 33598 11194 33654 11250
rect 33874 11194 33930 11250
rect 34150 11194 34206 11250
rect 34426 11194 34482 11250
rect 34702 11194 34758 11250
rect 34978 11194 35034 11250
rect 35254 11194 35310 11250
rect 35530 11194 35586 11250
rect 35806 11194 35862 11250
rect 36082 11194 36138 11250
rect 36358 11194 36414 11250
rect 36634 11194 36690 11250
rect 36910 11194 36966 11250
rect 37186 11194 37242 11250
rect 37462 11194 37518 11250
rect 37738 11194 37794 11250
rect 20076 11154 20128 11160
rect 19892 8492 19944 8498
rect 19812 8452 19892 8480
rect 19892 8434 19944 8440
rect 19800 8356 19852 8362
rect 19800 8298 19852 8304
rect 19812 5778 19840 8298
rect 20364 8294 20392 11194
rect 20640 11082 20668 11194
rect 20916 11150 20944 11194
rect 20904 11144 20956 11150
rect 20904 11086 20956 11092
rect 20628 11076 20680 11082
rect 20628 11018 20680 11024
rect 20902 9888 20958 9897
rect 21192 9874 21220 11194
rect 21192 9846 21404 9874
rect 20902 9823 20958 9832
rect 20444 9172 20496 9178
rect 20444 9114 20496 9120
rect 20352 8288 20404 8294
rect 20352 8230 20404 8236
rect 19950 8188 20258 8197
rect 19950 8186 19956 8188
rect 20012 8186 20036 8188
rect 20092 8186 20116 8188
rect 20172 8186 20196 8188
rect 20252 8186 20258 8188
rect 20012 8134 20014 8186
rect 20194 8134 20196 8186
rect 19950 8132 19956 8134
rect 20012 8132 20036 8134
rect 20092 8132 20116 8134
rect 20172 8132 20196 8134
rect 20252 8132 20258 8134
rect 19950 8123 20258 8132
rect 20456 7426 20484 9114
rect 20536 8628 20588 8634
rect 20536 8570 20588 8576
rect 20548 8090 20576 8570
rect 20916 8344 20944 9823
rect 21010 8732 21318 8741
rect 21010 8730 21016 8732
rect 21072 8730 21096 8732
rect 21152 8730 21176 8732
rect 21232 8730 21256 8732
rect 21312 8730 21318 8732
rect 21072 8678 21074 8730
rect 21254 8678 21256 8730
rect 21010 8676 21016 8678
rect 21072 8676 21096 8678
rect 21152 8676 21176 8678
rect 21232 8676 21256 8678
rect 21312 8676 21318 8678
rect 21010 8667 21318 8676
rect 21376 8498 21404 9846
rect 21364 8492 21416 8498
rect 21468 8480 21496 11194
rect 21744 8566 21772 11194
rect 22020 8634 22048 11194
rect 22296 9874 22324 11194
rect 22296 9846 22508 9874
rect 22100 9444 22152 9450
rect 22100 9386 22152 9392
rect 22008 8628 22060 8634
rect 22008 8570 22060 8576
rect 21732 8560 21784 8566
rect 21732 8502 21784 8508
rect 21548 8492 21600 8498
rect 21468 8452 21548 8480
rect 21364 8434 21416 8440
rect 21548 8434 21600 8440
rect 22112 8362 22140 9386
rect 22480 8498 22508 9846
rect 22572 8566 22600 11194
rect 22848 9874 22876 11194
rect 22848 9846 22968 9874
rect 22652 9172 22704 9178
rect 22652 9114 22704 9120
rect 22664 8974 22692 9114
rect 22652 8968 22704 8974
rect 22652 8910 22704 8916
rect 22560 8560 22612 8566
rect 22560 8502 22612 8508
rect 22468 8492 22520 8498
rect 22468 8434 22520 8440
rect 22940 8430 22968 9846
rect 23124 8634 23152 11194
rect 23204 9104 23256 9110
rect 23204 9046 23256 9052
rect 23112 8628 23164 8634
rect 23112 8570 23164 8576
rect 22928 8424 22980 8430
rect 22928 8366 22980 8372
rect 23216 8362 23244 9046
rect 23400 8362 23428 11194
rect 23480 9376 23532 9382
rect 23480 9318 23532 9324
rect 21640 8356 21692 8362
rect 20916 8316 21588 8344
rect 20536 8084 20588 8090
rect 20536 8026 20588 8032
rect 20628 8016 20680 8022
rect 20628 7958 20680 7964
rect 20718 7984 20774 7993
rect 20536 7880 20588 7886
rect 20536 7822 20588 7828
rect 20364 7398 20484 7426
rect 19950 7100 20258 7109
rect 19950 7098 19956 7100
rect 20012 7098 20036 7100
rect 20092 7098 20116 7100
rect 20172 7098 20196 7100
rect 20252 7098 20258 7100
rect 20012 7046 20014 7098
rect 20194 7046 20196 7098
rect 19950 7044 19956 7046
rect 20012 7044 20036 7046
rect 20092 7044 20116 7046
rect 20172 7044 20196 7046
rect 20252 7044 20258 7046
rect 19950 7035 20258 7044
rect 20364 6848 20392 7398
rect 20444 7336 20496 7342
rect 20444 7278 20496 7284
rect 20272 6820 20392 6848
rect 20168 6792 20220 6798
rect 20272 6780 20300 6820
rect 20220 6752 20300 6780
rect 20168 6734 20220 6740
rect 20180 6497 20208 6734
rect 20456 6730 20484 7278
rect 20548 7041 20576 7822
rect 20640 7732 20668 7958
rect 20718 7919 20774 7928
rect 20902 7984 20958 7993
rect 20902 7919 20958 7928
rect 20732 7886 20760 7919
rect 20720 7880 20772 7886
rect 20720 7822 20772 7828
rect 20640 7704 20760 7732
rect 20626 7168 20682 7177
rect 20626 7103 20682 7112
rect 20534 7032 20590 7041
rect 20640 7002 20668 7103
rect 20534 6967 20590 6976
rect 20628 6996 20680 7002
rect 20628 6938 20680 6944
rect 20536 6792 20588 6798
rect 20536 6734 20588 6740
rect 20626 6760 20682 6769
rect 20444 6724 20496 6730
rect 20444 6666 20496 6672
rect 20166 6488 20222 6497
rect 20166 6423 20222 6432
rect 20350 6352 20406 6361
rect 20350 6287 20406 6296
rect 20444 6316 20496 6322
rect 20364 6089 20392 6287
rect 20444 6258 20496 6264
rect 20350 6080 20406 6089
rect 19950 6012 20258 6021
rect 20350 6015 20406 6024
rect 19950 6010 19956 6012
rect 20012 6010 20036 6012
rect 20092 6010 20116 6012
rect 20172 6010 20196 6012
rect 20252 6010 20258 6012
rect 20012 5958 20014 6010
rect 20194 5958 20196 6010
rect 19950 5956 19956 5958
rect 20012 5956 20036 5958
rect 20092 5956 20116 5958
rect 20172 5956 20196 5958
rect 20252 5956 20258 5958
rect 19950 5947 20258 5956
rect 20352 5908 20404 5914
rect 20352 5850 20404 5856
rect 19800 5772 19852 5778
rect 19800 5714 19852 5720
rect 19708 5704 19760 5710
rect 19708 5646 19760 5652
rect 19432 5568 19484 5574
rect 19432 5510 19484 5516
rect 19300 5120 19380 5148
rect 19248 5102 19300 5108
rect 18880 4140 18932 4146
rect 18880 4082 18932 4088
rect 18696 3392 18748 3398
rect 18696 3334 18748 3340
rect 19260 2854 19288 5102
rect 19444 3534 19472 5510
rect 19706 5400 19762 5409
rect 19706 5335 19762 5344
rect 19720 5234 19748 5335
rect 19708 5228 19760 5234
rect 19708 5170 19760 5176
rect 19708 4480 19760 4486
rect 19708 4422 19760 4428
rect 19524 4276 19576 4282
rect 19524 4218 19576 4224
rect 19536 3670 19564 4218
rect 19616 3936 19668 3942
rect 19720 3913 19748 4422
rect 19616 3878 19668 3884
rect 19706 3904 19762 3913
rect 19524 3664 19576 3670
rect 19524 3606 19576 3612
rect 19628 3534 19656 3878
rect 19706 3839 19762 3848
rect 19812 3602 19840 5714
rect 20364 5710 20392 5850
rect 20352 5704 20404 5710
rect 20352 5646 20404 5652
rect 20352 5296 20404 5302
rect 20352 5238 20404 5244
rect 20364 5030 20392 5238
rect 20352 5024 20404 5030
rect 20352 4966 20404 4972
rect 19950 4924 20258 4933
rect 19950 4922 19956 4924
rect 20012 4922 20036 4924
rect 20092 4922 20116 4924
rect 20172 4922 20196 4924
rect 20252 4922 20258 4924
rect 20012 4870 20014 4922
rect 20194 4870 20196 4922
rect 19950 4868 19956 4870
rect 20012 4868 20036 4870
rect 20092 4868 20116 4870
rect 20172 4868 20196 4870
rect 20252 4868 20258 4870
rect 19950 4859 20258 4868
rect 20260 4140 20312 4146
rect 20456 4128 20484 6258
rect 20548 6254 20576 6734
rect 20626 6695 20682 6704
rect 20536 6248 20588 6254
rect 20536 6190 20588 6196
rect 20536 6112 20588 6118
rect 20536 6054 20588 6060
rect 20312 4100 20484 4128
rect 20260 4082 20312 4088
rect 20352 4004 20404 4010
rect 20352 3946 20404 3952
rect 20364 3913 20392 3946
rect 20350 3904 20406 3913
rect 19950 3836 20258 3845
rect 20350 3839 20406 3848
rect 19950 3834 19956 3836
rect 20012 3834 20036 3836
rect 20092 3834 20116 3836
rect 20172 3834 20196 3836
rect 20252 3834 20258 3836
rect 20012 3782 20014 3834
rect 20194 3782 20196 3834
rect 19950 3780 19956 3782
rect 20012 3780 20036 3782
rect 20092 3780 20116 3782
rect 20172 3780 20196 3782
rect 20252 3780 20258 3782
rect 19950 3771 20258 3780
rect 19800 3596 19852 3602
rect 19800 3538 19852 3544
rect 20548 3534 20576 6054
rect 20640 5914 20668 6695
rect 20628 5908 20680 5914
rect 20628 5850 20680 5856
rect 20732 4622 20760 7704
rect 20810 7712 20866 7721
rect 20810 7647 20866 7656
rect 20824 7290 20852 7647
rect 20916 7449 20944 7919
rect 21010 7644 21318 7653
rect 21010 7642 21016 7644
rect 21072 7642 21096 7644
rect 21152 7642 21176 7644
rect 21232 7642 21256 7644
rect 21312 7642 21318 7644
rect 21072 7590 21074 7642
rect 21254 7590 21256 7642
rect 21010 7588 21016 7590
rect 21072 7588 21096 7590
rect 21152 7588 21176 7590
rect 21232 7588 21256 7590
rect 21312 7588 21318 7590
rect 21010 7579 21318 7588
rect 21272 7472 21324 7478
rect 20902 7440 20958 7449
rect 21272 7414 21324 7420
rect 20902 7375 20958 7384
rect 21178 7304 21234 7313
rect 20824 7262 21178 7290
rect 21178 7239 21234 7248
rect 21284 6746 21312 7414
rect 21364 7336 21416 7342
rect 21364 7278 21416 7284
rect 20824 6718 21312 6746
rect 20720 4616 20772 4622
rect 20720 4558 20772 4564
rect 19432 3528 19484 3534
rect 19432 3470 19484 3476
rect 19616 3528 19668 3534
rect 19616 3470 19668 3476
rect 20536 3528 20588 3534
rect 20536 3470 20588 3476
rect 20824 3466 20852 6718
rect 20904 6656 20956 6662
rect 20904 6598 20956 6604
rect 20916 5778 20944 6598
rect 21010 6556 21318 6565
rect 21010 6554 21016 6556
rect 21072 6554 21096 6556
rect 21152 6554 21176 6556
rect 21232 6554 21256 6556
rect 21312 6554 21318 6556
rect 21072 6502 21074 6554
rect 21254 6502 21256 6554
rect 21010 6500 21016 6502
rect 21072 6500 21096 6502
rect 21152 6500 21176 6502
rect 21232 6500 21256 6502
rect 21312 6500 21318 6502
rect 21010 6491 21318 6500
rect 20996 6452 21048 6458
rect 20996 6394 21048 6400
rect 20904 5772 20956 5778
rect 20904 5714 20956 5720
rect 21008 5658 21036 6394
rect 21180 5908 21232 5914
rect 21180 5850 21232 5856
rect 20916 5630 21036 5658
rect 20812 3460 20864 3466
rect 20812 3402 20864 3408
rect 19340 3392 19392 3398
rect 19340 3334 19392 3340
rect 19352 3126 19380 3334
rect 19340 3120 19392 3126
rect 19340 3062 19392 3068
rect 20350 3088 20406 3097
rect 20916 3058 20944 5630
rect 21192 5574 21220 5850
rect 21180 5568 21232 5574
rect 21180 5510 21232 5516
rect 21010 5468 21318 5477
rect 21010 5466 21016 5468
rect 21072 5466 21096 5468
rect 21152 5466 21176 5468
rect 21232 5466 21256 5468
rect 21312 5466 21318 5468
rect 21072 5414 21074 5466
rect 21254 5414 21256 5466
rect 21010 5412 21016 5414
rect 21072 5412 21096 5414
rect 21152 5412 21176 5414
rect 21232 5412 21256 5414
rect 21312 5412 21318 5414
rect 21010 5403 21318 5412
rect 21010 4380 21318 4389
rect 21010 4378 21016 4380
rect 21072 4378 21096 4380
rect 21152 4378 21176 4380
rect 21232 4378 21256 4380
rect 21312 4378 21318 4380
rect 21072 4326 21074 4378
rect 21254 4326 21256 4378
rect 21010 4324 21016 4326
rect 21072 4324 21096 4326
rect 21152 4324 21176 4326
rect 21232 4324 21256 4326
rect 21312 4324 21318 4326
rect 21010 4315 21318 4324
rect 21376 3670 21404 7278
rect 21456 6656 21508 6662
rect 21456 6598 21508 6604
rect 21468 5914 21496 6598
rect 21560 5914 21588 8316
rect 21640 8298 21692 8304
rect 22100 8356 22152 8362
rect 22100 8298 22152 8304
rect 22468 8356 22520 8362
rect 22468 8298 22520 8304
rect 22836 8356 22888 8362
rect 22836 8298 22888 8304
rect 23204 8356 23256 8362
rect 23204 8298 23256 8304
rect 23388 8356 23440 8362
rect 23388 8298 23440 8304
rect 21456 5908 21508 5914
rect 21456 5850 21508 5856
rect 21548 5908 21600 5914
rect 21548 5850 21600 5856
rect 21456 5568 21508 5574
rect 21456 5510 21508 5516
rect 21548 5568 21600 5574
rect 21548 5510 21600 5516
rect 21468 4146 21496 5510
rect 21560 4185 21588 5510
rect 21652 4826 21680 8298
rect 21732 8288 21784 8294
rect 21732 8230 21784 8236
rect 21744 7478 21772 8230
rect 22376 7744 22428 7750
rect 22376 7686 22428 7692
rect 22282 7576 22338 7585
rect 21916 7540 21968 7546
rect 22282 7511 22338 7520
rect 21916 7482 21968 7488
rect 21732 7472 21784 7478
rect 21732 7414 21784 7420
rect 21824 7472 21876 7478
rect 21824 7414 21876 7420
rect 21730 7168 21786 7177
rect 21730 7103 21786 7112
rect 21744 6798 21772 7103
rect 21732 6792 21784 6798
rect 21732 6734 21784 6740
rect 21730 6624 21786 6633
rect 21730 6559 21786 6568
rect 21744 5953 21772 6559
rect 21730 5944 21786 5953
rect 21730 5879 21786 5888
rect 21732 5840 21784 5846
rect 21732 5782 21784 5788
rect 21744 5545 21772 5782
rect 21730 5536 21786 5545
rect 21730 5471 21786 5480
rect 21730 4856 21786 4865
rect 21640 4820 21692 4826
rect 21730 4791 21732 4800
rect 21640 4762 21692 4768
rect 21784 4791 21786 4800
rect 21732 4762 21784 4768
rect 21546 4176 21602 4185
rect 21456 4140 21508 4146
rect 21546 4111 21602 4120
rect 21456 4082 21508 4088
rect 21364 3664 21416 3670
rect 21364 3606 21416 3612
rect 21652 3534 21680 4762
rect 21836 4282 21864 7414
rect 21928 6610 21956 7482
rect 22296 7478 22324 7511
rect 22388 7478 22416 7686
rect 22284 7472 22336 7478
rect 22284 7414 22336 7420
rect 22376 7472 22428 7478
rect 22376 7414 22428 7420
rect 22100 7404 22152 7410
rect 22100 7346 22152 7352
rect 22008 7336 22060 7342
rect 22008 7278 22060 7284
rect 22020 7002 22048 7278
rect 22008 6996 22060 7002
rect 22008 6938 22060 6944
rect 22006 6896 22062 6905
rect 22006 6831 22062 6840
rect 22020 6712 22048 6831
rect 22112 6780 22140 7346
rect 22480 7002 22508 8298
rect 22744 7336 22796 7342
rect 22744 7278 22796 7284
rect 22468 6996 22520 7002
rect 22468 6938 22520 6944
rect 22560 6928 22612 6934
rect 22560 6870 22612 6876
rect 22112 6752 22416 6780
rect 22020 6684 22140 6712
rect 21928 6582 22048 6610
rect 21916 6316 21968 6322
rect 21916 6258 21968 6264
rect 21928 5030 21956 6258
rect 22020 5710 22048 6582
rect 22112 6458 22140 6684
rect 22100 6452 22152 6458
rect 22100 6394 22152 6400
rect 22100 6316 22152 6322
rect 22100 6258 22152 6264
rect 22192 6316 22244 6322
rect 22192 6258 22244 6264
rect 22008 5704 22060 5710
rect 22008 5646 22060 5652
rect 21916 5024 21968 5030
rect 21916 4966 21968 4972
rect 21824 4276 21876 4282
rect 21824 4218 21876 4224
rect 22020 3738 22048 5646
rect 22112 3738 22140 6258
rect 22008 3732 22060 3738
rect 22008 3674 22060 3680
rect 22100 3732 22152 3738
rect 22100 3674 22152 3680
rect 21640 3528 21692 3534
rect 21640 3470 21692 3476
rect 21010 3292 21318 3301
rect 21010 3290 21016 3292
rect 21072 3290 21096 3292
rect 21152 3290 21176 3292
rect 21232 3290 21256 3292
rect 21312 3290 21318 3292
rect 21072 3238 21074 3290
rect 21254 3238 21256 3290
rect 21010 3236 21016 3238
rect 21072 3236 21096 3238
rect 21152 3236 21176 3238
rect 21232 3236 21256 3238
rect 21312 3236 21318 3238
rect 21010 3227 21318 3236
rect 22204 3194 22232 6258
rect 22284 6112 22336 6118
rect 22284 6054 22336 6060
rect 22296 4729 22324 6054
rect 22282 4720 22338 4729
rect 22282 4655 22338 4664
rect 22284 4072 22336 4078
rect 22284 4014 22336 4020
rect 22296 3466 22324 4014
rect 22388 3913 22416 6752
rect 22468 6656 22520 6662
rect 22468 6598 22520 6604
rect 22480 4486 22508 6598
rect 22468 4480 22520 4486
rect 22468 4422 22520 4428
rect 22572 3942 22600 6870
rect 22652 6724 22704 6730
rect 22652 6666 22704 6672
rect 22664 6497 22692 6666
rect 22650 6488 22706 6497
rect 22650 6423 22706 6432
rect 22664 6254 22692 6423
rect 22652 6248 22704 6254
rect 22652 6190 22704 6196
rect 22756 5234 22784 7278
rect 22848 6662 22876 8298
rect 22928 8288 22980 8294
rect 22928 8230 22980 8236
rect 22940 7954 22968 8230
rect 23388 8084 23440 8090
rect 23388 8026 23440 8032
rect 23020 8016 23072 8022
rect 23020 7958 23072 7964
rect 23204 8016 23256 8022
rect 23204 7958 23256 7964
rect 22928 7948 22980 7954
rect 22928 7890 22980 7896
rect 23032 7410 23060 7958
rect 23020 7404 23072 7410
rect 23020 7346 23072 7352
rect 23020 6996 23072 7002
rect 22940 6956 23020 6984
rect 22836 6656 22888 6662
rect 22836 6598 22888 6604
rect 22744 5228 22796 5234
rect 22744 5170 22796 5176
rect 22652 5024 22704 5030
rect 22652 4966 22704 4972
rect 22664 4146 22692 4966
rect 22652 4140 22704 4146
rect 22652 4082 22704 4088
rect 22560 3936 22612 3942
rect 22374 3904 22430 3913
rect 22560 3878 22612 3884
rect 22374 3839 22430 3848
rect 22572 3670 22600 3878
rect 22560 3664 22612 3670
rect 22560 3606 22612 3612
rect 22284 3460 22336 3466
rect 22284 3402 22336 3408
rect 22192 3188 22244 3194
rect 22192 3130 22244 3136
rect 22572 3058 22600 3606
rect 22664 3602 22692 4082
rect 22848 4078 22876 6598
rect 22836 4072 22888 4078
rect 22836 4014 22888 4020
rect 22652 3596 22704 3602
rect 22652 3538 22704 3544
rect 22940 3058 22968 6956
rect 23020 6938 23072 6944
rect 23112 6792 23164 6798
rect 23112 6734 23164 6740
rect 23124 6633 23152 6734
rect 23110 6624 23166 6633
rect 23110 6559 23166 6568
rect 23112 6248 23164 6254
rect 23112 6190 23164 6196
rect 23020 6112 23072 6118
rect 23020 6054 23072 6060
rect 23032 3738 23060 6054
rect 23020 3732 23072 3738
rect 23020 3674 23072 3680
rect 23124 3126 23152 6190
rect 23112 3120 23164 3126
rect 23112 3062 23164 3068
rect 20350 3023 20406 3032
rect 20904 3052 20956 3058
rect 19248 2848 19300 2854
rect 20364 2825 20392 3023
rect 20904 2994 20956 3000
rect 22560 3052 22612 3058
rect 22560 2994 22612 3000
rect 22928 3052 22980 3058
rect 22928 2994 22980 3000
rect 22008 2984 22060 2990
rect 22008 2926 22060 2932
rect 19248 2790 19300 2796
rect 20350 2816 20406 2825
rect 19950 2748 20258 2757
rect 20350 2751 20406 2760
rect 19950 2746 19956 2748
rect 20012 2746 20036 2748
rect 20092 2746 20116 2748
rect 20172 2746 20196 2748
rect 20252 2746 20258 2748
rect 20012 2694 20014 2746
rect 20194 2694 20196 2746
rect 19950 2692 19956 2694
rect 20012 2692 20036 2694
rect 20092 2692 20116 2694
rect 20172 2692 20196 2694
rect 20252 2692 20258 2694
rect 19950 2683 20258 2692
rect 21010 2204 21318 2213
rect 21010 2202 21016 2204
rect 21072 2202 21096 2204
rect 21152 2202 21176 2204
rect 21232 2202 21256 2204
rect 21312 2202 21318 2204
rect 21072 2150 21074 2202
rect 21254 2150 21256 2202
rect 21010 2148 21016 2150
rect 21072 2148 21096 2150
rect 21152 2148 21176 2150
rect 21232 2148 21256 2150
rect 21312 2148 21318 2150
rect 21010 2139 21318 2148
rect 17500 2100 17552 2106
rect 17500 2042 17552 2048
rect 20444 2100 20496 2106
rect 20444 2042 20496 2048
rect 18892 190 19012 218
rect 18892 56 18920 190
rect 18984 134 19012 190
rect 18972 128 19024 134
rect 18972 70 19024 76
rect 20456 56 20484 2042
rect 22020 56 22048 2926
rect 23216 2922 23244 7958
rect 23400 7449 23428 8026
rect 23386 7440 23442 7449
rect 23386 7375 23442 7384
rect 23492 6118 23520 9318
rect 23676 8566 23704 11194
rect 23848 9172 23900 9178
rect 23848 9114 23900 9120
rect 23756 8832 23808 8838
rect 23756 8774 23808 8780
rect 23768 8634 23796 8774
rect 23756 8628 23808 8634
rect 23756 8570 23808 8576
rect 23664 8560 23716 8566
rect 23664 8502 23716 8508
rect 23572 8288 23624 8294
rect 23572 8230 23624 8236
rect 23756 8288 23808 8294
rect 23756 8230 23808 8236
rect 23584 6730 23612 8230
rect 23768 8022 23796 8230
rect 23756 8016 23808 8022
rect 23756 7958 23808 7964
rect 23664 6860 23716 6866
rect 23664 6802 23716 6808
rect 23572 6724 23624 6730
rect 23572 6666 23624 6672
rect 23480 6112 23532 6118
rect 23480 6054 23532 6060
rect 23480 5636 23532 5642
rect 23480 5578 23532 5584
rect 23296 4072 23348 4078
rect 23296 4014 23348 4020
rect 23308 3942 23336 4014
rect 23296 3936 23348 3942
rect 23296 3878 23348 3884
rect 23388 3936 23440 3942
rect 23388 3878 23440 3884
rect 23308 3738 23336 3878
rect 23296 3732 23348 3738
rect 23296 3674 23348 3680
rect 23296 3528 23348 3534
rect 23400 3516 23428 3878
rect 23492 3602 23520 5578
rect 23480 3596 23532 3602
rect 23480 3538 23532 3544
rect 23348 3488 23428 3516
rect 23584 3482 23612 6666
rect 23676 6497 23704 6802
rect 23662 6488 23718 6497
rect 23860 6474 23888 9114
rect 23952 8634 23980 11194
rect 24030 10296 24086 10305
rect 24030 10231 24086 10240
rect 23940 8628 23992 8634
rect 23940 8570 23992 8576
rect 24044 8362 24072 10231
rect 24124 10056 24176 10062
rect 24124 9998 24176 10004
rect 24032 8356 24084 8362
rect 24032 8298 24084 8304
rect 24136 7410 24164 9998
rect 24228 9874 24256 11194
rect 24228 9846 24348 9874
rect 24320 8430 24348 9846
rect 24400 9512 24452 9518
rect 24400 9454 24452 9460
rect 24308 8424 24360 8430
rect 24308 8366 24360 8372
rect 24216 8356 24268 8362
rect 24216 8298 24268 8304
rect 24124 7404 24176 7410
rect 24124 7346 24176 7352
rect 23860 6446 23980 6474
rect 23662 6423 23718 6432
rect 23848 6384 23900 6390
rect 23848 6326 23900 6332
rect 23756 6316 23808 6322
rect 23756 6258 23808 6264
rect 23768 4214 23796 6258
rect 23860 4282 23888 6326
rect 23952 6254 23980 6446
rect 23940 6248 23992 6254
rect 23940 6190 23992 6196
rect 24228 5710 24256 8298
rect 24308 5908 24360 5914
rect 24308 5850 24360 5856
rect 24216 5704 24268 5710
rect 24216 5646 24268 5652
rect 23848 4276 23900 4282
rect 23848 4218 23900 4224
rect 23756 4208 23808 4214
rect 23756 4150 23808 4156
rect 24228 3670 24256 5646
rect 24320 5574 24348 5850
rect 24412 5574 24440 9454
rect 24504 8548 24532 11194
rect 24780 8634 24808 11194
rect 24768 8628 24820 8634
rect 24768 8570 24820 8576
rect 24676 8560 24728 8566
rect 24504 8520 24676 8548
rect 24676 8502 24728 8508
rect 25056 8430 25084 11194
rect 25134 10432 25190 10441
rect 25134 10367 25190 10376
rect 25044 8424 25096 8430
rect 25044 8366 25096 8372
rect 24768 8356 24820 8362
rect 24768 8298 24820 8304
rect 24674 8256 24730 8265
rect 24674 8191 24730 8200
rect 24584 7744 24636 7750
rect 24584 7686 24636 7692
rect 24492 6860 24544 6866
rect 24492 6802 24544 6808
rect 24308 5568 24360 5574
rect 24308 5510 24360 5516
rect 24400 5568 24452 5574
rect 24400 5510 24452 5516
rect 24504 3670 24532 6802
rect 24596 5710 24624 7686
rect 24688 6662 24716 8191
rect 24780 7206 24808 8298
rect 24768 7200 24820 7206
rect 24768 7142 24820 7148
rect 25148 6662 25176 10367
rect 25228 9240 25280 9246
rect 25228 9182 25280 9188
rect 25240 8362 25268 9182
rect 25332 8566 25360 11194
rect 25504 8900 25556 8906
rect 25504 8842 25556 8848
rect 25516 8634 25544 8842
rect 25504 8628 25556 8634
rect 25504 8570 25556 8576
rect 25320 8560 25372 8566
rect 25320 8502 25372 8508
rect 25228 8356 25280 8362
rect 25228 8298 25280 8304
rect 25320 8356 25372 8362
rect 25320 8298 25372 8304
rect 24676 6656 24728 6662
rect 24676 6598 24728 6604
rect 25136 6656 25188 6662
rect 25136 6598 25188 6604
rect 24768 6248 24820 6254
rect 24768 6190 24820 6196
rect 24676 6112 24728 6118
rect 24676 6054 24728 6060
rect 24584 5704 24636 5710
rect 24584 5646 24636 5652
rect 24688 5574 24716 6054
rect 24676 5568 24728 5574
rect 24676 5510 24728 5516
rect 24780 4146 24808 6190
rect 25332 6089 25360 8298
rect 25504 7472 25556 7478
rect 25504 7414 25556 7420
rect 25318 6080 25374 6089
rect 25318 6015 25374 6024
rect 24860 5704 24912 5710
rect 24860 5646 24912 5652
rect 24768 4140 24820 4146
rect 24768 4082 24820 4088
rect 24872 3942 24900 5646
rect 25516 4593 25544 7414
rect 25608 6934 25636 11194
rect 25884 9042 25912 11194
rect 25872 9036 25924 9042
rect 25872 8978 25924 8984
rect 26160 8838 26188 11194
rect 26148 8832 26200 8838
rect 26148 8774 26200 8780
rect 25688 8628 25740 8634
rect 25688 8570 25740 8576
rect 25596 6928 25648 6934
rect 25596 6870 25648 6876
rect 25700 5710 25728 8570
rect 26332 8356 26384 8362
rect 26332 8298 26384 8304
rect 25780 8288 25832 8294
rect 25780 8230 25832 8236
rect 25792 6610 25820 8230
rect 25950 8188 26258 8197
rect 25950 8186 25956 8188
rect 26012 8186 26036 8188
rect 26092 8186 26116 8188
rect 26172 8186 26196 8188
rect 26252 8186 26258 8188
rect 26012 8134 26014 8186
rect 26194 8134 26196 8186
rect 25950 8132 25956 8134
rect 26012 8132 26036 8134
rect 26092 8132 26116 8134
rect 26172 8132 26196 8134
rect 26252 8132 26258 8134
rect 25950 8123 26258 8132
rect 25950 7100 26258 7109
rect 25950 7098 25956 7100
rect 26012 7098 26036 7100
rect 26092 7098 26116 7100
rect 26172 7098 26196 7100
rect 26252 7098 26258 7100
rect 26012 7046 26014 7098
rect 26194 7046 26196 7098
rect 25950 7044 25956 7046
rect 26012 7044 26036 7046
rect 26092 7044 26116 7046
rect 26172 7044 26196 7046
rect 26252 7044 26258 7046
rect 25950 7035 26258 7044
rect 25792 6582 25912 6610
rect 25688 5704 25740 5710
rect 25688 5646 25740 5652
rect 25884 5234 25912 6582
rect 25950 6012 26258 6021
rect 25950 6010 25956 6012
rect 26012 6010 26036 6012
rect 26092 6010 26116 6012
rect 26172 6010 26196 6012
rect 26252 6010 26258 6012
rect 26012 5958 26014 6010
rect 26194 5958 26196 6010
rect 25950 5956 25956 5958
rect 26012 5956 26036 5958
rect 26092 5956 26116 5958
rect 26172 5956 26196 5958
rect 26252 5956 26258 5958
rect 25950 5947 26258 5956
rect 26344 5545 26372 8298
rect 26436 6866 26464 11194
rect 26608 9920 26660 9926
rect 26608 9862 26660 9868
rect 26516 8560 26568 8566
rect 26516 8502 26568 8508
rect 26424 6860 26476 6866
rect 26424 6802 26476 6808
rect 26528 6322 26556 8502
rect 26516 6316 26568 6322
rect 26516 6258 26568 6264
rect 26330 5536 26386 5545
rect 26330 5471 26386 5480
rect 25872 5228 25924 5234
rect 25872 5170 25924 5176
rect 25502 4584 25558 4593
rect 25502 4519 25558 4528
rect 25044 4480 25096 4486
rect 25044 4422 25096 4428
rect 24860 3936 24912 3942
rect 24860 3878 24912 3884
rect 24216 3664 24268 3670
rect 24216 3606 24268 3612
rect 24492 3664 24544 3670
rect 24492 3606 24544 3612
rect 23296 3470 23348 3476
rect 23492 3454 23612 3482
rect 23492 3398 23520 3454
rect 23480 3392 23532 3398
rect 23480 3334 23532 3340
rect 23572 3392 23624 3398
rect 23572 3334 23624 3340
rect 23204 2916 23256 2922
rect 23204 2858 23256 2864
rect 23584 56 23612 3334
rect 25056 202 25084 4422
rect 25884 3738 25912 5170
rect 26620 5098 26648 9862
rect 26712 6390 26740 11194
rect 26792 10124 26844 10130
rect 26792 10066 26844 10072
rect 26804 6662 26832 10066
rect 26988 9058 27016 11194
rect 27264 9194 27292 11194
rect 27264 9166 27476 9194
rect 26988 9030 27384 9058
rect 27010 8732 27318 8741
rect 27010 8730 27016 8732
rect 27072 8730 27096 8732
rect 27152 8730 27176 8732
rect 27232 8730 27256 8732
rect 27312 8730 27318 8732
rect 27072 8678 27074 8730
rect 27254 8678 27256 8730
rect 27010 8676 27016 8678
rect 27072 8676 27096 8678
rect 27152 8676 27176 8678
rect 27232 8676 27256 8678
rect 27312 8676 27318 8678
rect 27010 8667 27318 8676
rect 26884 8288 26936 8294
rect 26884 8230 26936 8236
rect 26792 6656 26844 6662
rect 26792 6598 26844 6604
rect 26700 6384 26752 6390
rect 26700 6326 26752 6332
rect 26700 5772 26752 5778
rect 26700 5714 26752 5720
rect 26608 5092 26660 5098
rect 26608 5034 26660 5040
rect 25950 4924 26258 4933
rect 25950 4922 25956 4924
rect 26012 4922 26036 4924
rect 26092 4922 26116 4924
rect 26172 4922 26196 4924
rect 26252 4922 26258 4924
rect 26012 4870 26014 4922
rect 26194 4870 26196 4922
rect 25950 4868 25956 4870
rect 26012 4868 26036 4870
rect 26092 4868 26116 4870
rect 26172 4868 26196 4870
rect 26252 4868 26258 4870
rect 25950 4859 26258 4868
rect 25950 3836 26258 3845
rect 25950 3834 25956 3836
rect 26012 3834 26036 3836
rect 26092 3834 26116 3836
rect 26172 3834 26196 3836
rect 26252 3834 26258 3836
rect 26012 3782 26014 3834
rect 26194 3782 26196 3834
rect 25950 3780 25956 3782
rect 26012 3780 26036 3782
rect 26092 3780 26116 3782
rect 26172 3780 26196 3782
rect 26252 3780 26258 3782
rect 25950 3771 26258 3780
rect 26514 3768 26570 3777
rect 25872 3732 25924 3738
rect 26514 3703 26570 3712
rect 25872 3674 25924 3680
rect 26332 3460 26384 3466
rect 26332 3402 26384 3408
rect 25778 3224 25834 3233
rect 25778 3159 25834 3168
rect 25792 2825 25820 3159
rect 26344 2854 26372 3402
rect 26528 3233 26556 3703
rect 26606 3496 26662 3505
rect 26606 3431 26662 3440
rect 26514 3224 26570 3233
rect 26514 3159 26570 3168
rect 26332 2848 26384 2854
rect 25778 2816 25834 2825
rect 26620 2825 26648 3431
rect 26332 2790 26384 2796
rect 26606 2816 26662 2825
rect 25778 2751 25834 2760
rect 25950 2748 26258 2757
rect 26606 2751 26662 2760
rect 25950 2746 25956 2748
rect 26012 2746 26036 2748
rect 26092 2746 26116 2748
rect 26172 2746 26196 2748
rect 26252 2746 26258 2748
rect 26012 2694 26014 2746
rect 26194 2694 26196 2746
rect 25950 2692 25956 2694
rect 26012 2692 26036 2694
rect 26092 2692 26116 2694
rect 26172 2692 26196 2694
rect 26252 2692 26258 2694
rect 25950 2683 26258 2692
rect 25136 876 25188 882
rect 25136 818 25188 824
rect 25044 196 25096 202
rect 25044 138 25096 144
rect 25148 56 25176 818
rect 26712 56 26740 5714
rect 26896 5710 26924 8230
rect 27010 7644 27318 7653
rect 27010 7642 27016 7644
rect 27072 7642 27096 7644
rect 27152 7642 27176 7644
rect 27232 7642 27256 7644
rect 27312 7642 27318 7644
rect 27072 7590 27074 7642
rect 27254 7590 27256 7642
rect 27010 7588 27016 7590
rect 27072 7588 27096 7590
rect 27152 7588 27176 7590
rect 27232 7588 27256 7590
rect 27312 7588 27318 7590
rect 27010 7579 27318 7588
rect 27252 7404 27304 7410
rect 27252 7346 27304 7352
rect 27264 6662 27292 7346
rect 27356 7002 27384 9030
rect 27344 6996 27396 7002
rect 27344 6938 27396 6944
rect 27252 6656 27304 6662
rect 27252 6598 27304 6604
rect 27010 6556 27318 6565
rect 27010 6554 27016 6556
rect 27072 6554 27096 6556
rect 27152 6554 27176 6556
rect 27232 6554 27256 6556
rect 27312 6554 27318 6556
rect 27072 6502 27074 6554
rect 27254 6502 27256 6554
rect 27010 6500 27016 6502
rect 27072 6500 27096 6502
rect 27152 6500 27176 6502
rect 27232 6500 27256 6502
rect 27312 6500 27318 6502
rect 27010 6491 27318 6500
rect 27448 6322 27476 9166
rect 27436 6316 27488 6322
rect 27436 6258 27488 6264
rect 27540 6254 27568 11194
rect 27816 8498 27844 11194
rect 28092 9874 28120 11194
rect 28092 9846 28212 9874
rect 27986 9208 28042 9217
rect 27986 9143 28042 9152
rect 27896 9036 27948 9042
rect 27896 8978 27948 8984
rect 27804 8492 27856 8498
rect 27804 8434 27856 8440
rect 27712 6928 27764 6934
rect 27710 6896 27712 6905
rect 27764 6896 27766 6905
rect 27710 6831 27766 6840
rect 27908 6798 27936 8978
rect 27896 6792 27948 6798
rect 27896 6734 27948 6740
rect 28000 6662 28028 9143
rect 28184 8498 28212 9846
rect 28262 9480 28318 9489
rect 28262 9415 28318 9424
rect 28172 8492 28224 8498
rect 28172 8434 28224 8440
rect 28172 6792 28224 6798
rect 28172 6734 28224 6740
rect 27988 6656 28040 6662
rect 27988 6598 28040 6604
rect 27528 6248 27580 6254
rect 27528 6190 27580 6196
rect 28184 6186 28212 6734
rect 28276 6662 28304 9415
rect 28368 8498 28396 11194
rect 28540 9852 28592 9858
rect 28540 9794 28592 9800
rect 28448 8832 28500 8838
rect 28448 8774 28500 8780
rect 28356 8492 28408 8498
rect 28356 8434 28408 8440
rect 28460 6798 28488 8774
rect 28448 6792 28500 6798
rect 28448 6734 28500 6740
rect 28552 6662 28580 9794
rect 28644 7886 28672 11194
rect 28814 10160 28870 10169
rect 28814 10095 28870 10104
rect 28724 9784 28776 9790
rect 28724 9726 28776 9732
rect 28632 7880 28684 7886
rect 28632 7822 28684 7828
rect 28736 6662 28764 9726
rect 28828 7834 28856 10095
rect 28920 8022 28948 11194
rect 29196 8430 29224 11194
rect 29366 9752 29422 9761
rect 29366 9687 29422 9696
rect 29184 8424 29236 8430
rect 29184 8366 29236 8372
rect 28908 8016 28960 8022
rect 28908 7958 28960 7964
rect 29000 7948 29052 7954
rect 29000 7890 29052 7896
rect 28828 7806 28948 7834
rect 28816 7744 28868 7750
rect 28816 7686 28868 7692
rect 28828 7342 28856 7686
rect 28816 7336 28868 7342
rect 28816 7278 28868 7284
rect 28920 6662 28948 7806
rect 29012 6934 29040 7890
rect 29000 6928 29052 6934
rect 29000 6870 29052 6876
rect 29000 6792 29052 6798
rect 29000 6734 29052 6740
rect 28264 6656 28316 6662
rect 28264 6598 28316 6604
rect 28540 6656 28592 6662
rect 28540 6598 28592 6604
rect 28724 6656 28776 6662
rect 28724 6598 28776 6604
rect 28908 6656 28960 6662
rect 28908 6598 28960 6604
rect 29012 6390 29040 6734
rect 29184 6724 29236 6730
rect 29184 6666 29236 6672
rect 29000 6384 29052 6390
rect 29000 6326 29052 6332
rect 28172 6180 28224 6186
rect 28172 6122 28224 6128
rect 26884 5704 26936 5710
rect 26884 5646 26936 5652
rect 27010 5468 27318 5477
rect 27010 5466 27016 5468
rect 27072 5466 27096 5468
rect 27152 5466 27176 5468
rect 27232 5466 27256 5468
rect 27312 5466 27318 5468
rect 27072 5414 27074 5466
rect 27254 5414 27256 5466
rect 27010 5412 27016 5414
rect 27072 5412 27096 5414
rect 27152 5412 27176 5414
rect 27232 5412 27256 5414
rect 27312 5412 27318 5414
rect 27010 5403 27318 5412
rect 26884 5228 26936 5234
rect 26884 5170 26936 5176
rect 26896 882 26924 5170
rect 27010 4380 27318 4389
rect 27010 4378 27016 4380
rect 27072 4378 27096 4380
rect 27152 4378 27176 4380
rect 27232 4378 27256 4380
rect 27312 4378 27318 4380
rect 27072 4326 27074 4378
rect 27254 4326 27256 4378
rect 27010 4324 27016 4326
rect 27072 4324 27096 4326
rect 27152 4324 27176 4326
rect 27232 4324 27256 4326
rect 27312 4324 27318 4326
rect 27010 4315 27318 4324
rect 28264 4208 28316 4214
rect 28264 4150 28316 4156
rect 27010 3292 27318 3301
rect 27010 3290 27016 3292
rect 27072 3290 27096 3292
rect 27152 3290 27176 3292
rect 27232 3290 27256 3292
rect 27312 3290 27318 3292
rect 27072 3238 27074 3290
rect 27254 3238 27256 3290
rect 27010 3236 27016 3238
rect 27072 3236 27096 3238
rect 27152 3236 27176 3238
rect 27232 3236 27256 3238
rect 27312 3236 27318 3238
rect 27010 3227 27318 3236
rect 27010 2204 27318 2213
rect 27010 2202 27016 2204
rect 27072 2202 27096 2204
rect 27152 2202 27176 2204
rect 27232 2202 27256 2204
rect 27312 2202 27318 2204
rect 27072 2150 27074 2202
rect 27254 2150 27256 2202
rect 27010 2148 27016 2150
rect 27072 2148 27096 2150
rect 27152 2148 27176 2150
rect 27232 2148 27256 2150
rect 27312 2148 27318 2150
rect 27010 2139 27318 2148
rect 26884 876 26936 882
rect 26884 818 26936 824
rect 28276 56 28304 4150
rect 29196 3777 29224 6666
rect 29380 6662 29408 9687
rect 29472 7886 29500 11194
rect 29748 8498 29776 11194
rect 29920 9988 29972 9994
rect 29920 9930 29972 9936
rect 29736 8492 29788 8498
rect 29736 8434 29788 8440
rect 29826 7984 29882 7993
rect 29826 7919 29882 7928
rect 29460 7880 29512 7886
rect 29460 7822 29512 7828
rect 29552 7744 29604 7750
rect 29552 7686 29604 7692
rect 29564 7478 29592 7686
rect 29552 7472 29604 7478
rect 29552 7414 29604 7420
rect 29736 6792 29788 6798
rect 29736 6734 29788 6740
rect 29368 6656 29420 6662
rect 29368 6598 29420 6604
rect 29748 6322 29776 6734
rect 29840 6662 29868 7919
rect 29932 7886 29960 9930
rect 29920 7880 29972 7886
rect 29920 7822 29972 7828
rect 29918 7440 29974 7449
rect 30024 7410 30052 11194
rect 30104 8424 30156 8430
rect 30104 8366 30156 8372
rect 29918 7375 29974 7384
rect 30012 7404 30064 7410
rect 29828 6656 29880 6662
rect 29828 6598 29880 6604
rect 29736 6316 29788 6322
rect 29736 6258 29788 6264
rect 29182 3768 29238 3777
rect 29182 3703 29238 3712
rect 29932 3618 29960 7375
rect 30012 7346 30064 7352
rect 30012 6792 30064 6798
rect 30012 6734 30064 6740
rect 30024 6254 30052 6734
rect 30012 6248 30064 6254
rect 30012 6190 30064 6196
rect 30116 3738 30144 8366
rect 30300 7478 30328 11194
rect 30472 8968 30524 8974
rect 30472 8910 30524 8916
rect 30288 7472 30340 7478
rect 30288 7414 30340 7420
rect 30484 7206 30512 8910
rect 30576 7342 30604 11194
rect 30656 8968 30708 8974
rect 30656 8910 30708 8916
rect 30564 7336 30616 7342
rect 30564 7278 30616 7284
rect 30472 7200 30524 7206
rect 30472 7142 30524 7148
rect 30380 6996 30432 7002
rect 30380 6938 30432 6944
rect 30392 6361 30420 6938
rect 30378 6352 30434 6361
rect 30378 6287 30434 6296
rect 30380 6112 30432 6118
rect 30380 6054 30432 6060
rect 30392 4554 30420 6054
rect 30380 4548 30432 4554
rect 30380 4490 30432 4496
rect 30288 3936 30340 3942
rect 30288 3878 30340 3884
rect 30104 3732 30156 3738
rect 30104 3674 30156 3680
rect 29840 3590 29960 3618
rect 29840 56 29868 3590
rect 29920 3528 29972 3534
rect 29920 3470 29972 3476
rect 29932 66 29960 3470
rect 30300 1873 30328 3878
rect 30668 3738 30696 8910
rect 30748 7948 30800 7954
rect 30748 7890 30800 7896
rect 30760 4010 30788 7890
rect 30852 7546 30880 11194
rect 30932 8560 30984 8566
rect 30932 8502 30984 8508
rect 30840 7540 30892 7546
rect 30840 7482 30892 7488
rect 30944 4010 30972 8502
rect 31128 7750 31156 11194
rect 31300 7812 31352 7818
rect 31300 7754 31352 7760
rect 31116 7744 31168 7750
rect 31116 7686 31168 7692
rect 31312 7206 31340 7754
rect 31300 7200 31352 7206
rect 31300 7142 31352 7148
rect 31404 6798 31432 11194
rect 31482 9344 31538 9353
rect 31482 9279 31538 9288
rect 31392 6792 31444 6798
rect 31392 6734 31444 6740
rect 31496 6662 31524 9279
rect 31576 7880 31628 7886
rect 31576 7822 31628 7828
rect 31588 7206 31616 7822
rect 31680 7342 31708 11194
rect 31956 9058 31984 11194
rect 31864 9030 31984 9058
rect 31758 8528 31814 8537
rect 31758 8463 31814 8472
rect 31668 7336 31720 7342
rect 31668 7278 31720 7284
rect 31576 7200 31628 7206
rect 31576 7142 31628 7148
rect 31484 6656 31536 6662
rect 31772 6644 31800 8463
rect 31864 6866 31892 9030
rect 32232 8634 32260 11194
rect 32404 8900 32456 8906
rect 32404 8842 32456 8848
rect 32220 8628 32272 8634
rect 32220 8570 32272 8576
rect 31950 8188 32258 8197
rect 31950 8186 31956 8188
rect 32012 8186 32036 8188
rect 32092 8186 32116 8188
rect 32172 8186 32196 8188
rect 32252 8186 32258 8188
rect 32012 8134 32014 8186
rect 32194 8134 32196 8186
rect 31950 8132 31956 8134
rect 32012 8132 32036 8134
rect 32092 8132 32116 8134
rect 32172 8132 32196 8134
rect 32252 8132 32258 8134
rect 31950 8123 32258 8132
rect 32126 7848 32182 7857
rect 32126 7783 32182 7792
rect 32140 7206 32168 7783
rect 32416 7426 32444 8842
rect 32508 8634 32536 11194
rect 32588 9308 32640 9314
rect 32588 9250 32640 9256
rect 32496 8628 32548 8634
rect 32496 8570 32548 8576
rect 32600 8498 32628 9250
rect 32784 8650 32812 11194
rect 33060 8838 33088 11194
rect 33336 9466 33364 11194
rect 33336 9438 33456 9466
rect 33048 8832 33100 8838
rect 33048 8774 33100 8780
rect 33010 8732 33318 8741
rect 33010 8730 33016 8732
rect 33072 8730 33096 8732
rect 33152 8730 33176 8732
rect 33232 8730 33256 8732
rect 33312 8730 33318 8732
rect 33072 8678 33074 8730
rect 33254 8678 33256 8730
rect 33010 8676 33016 8678
rect 33072 8676 33096 8678
rect 33152 8676 33176 8678
rect 33232 8676 33256 8678
rect 33312 8676 33318 8678
rect 33010 8667 33318 8676
rect 32784 8634 32904 8650
rect 32784 8628 32916 8634
rect 32784 8622 32864 8628
rect 32864 8570 32916 8576
rect 33048 8560 33100 8566
rect 33048 8502 33100 8508
rect 32588 8492 32640 8498
rect 32588 8434 32640 8440
rect 33060 7800 33088 8502
rect 33428 8362 33456 9438
rect 33508 8832 33560 8838
rect 33508 8774 33560 8780
rect 33520 8634 33548 8774
rect 33612 8634 33640 11194
rect 33784 8968 33836 8974
rect 33784 8910 33836 8916
rect 33508 8628 33560 8634
rect 33508 8570 33560 8576
rect 33600 8628 33652 8634
rect 33600 8570 33652 8576
rect 33796 8566 33824 8910
rect 33784 8560 33836 8566
rect 33784 8502 33836 8508
rect 33508 8492 33560 8498
rect 33508 8434 33560 8440
rect 33416 8356 33468 8362
rect 33416 8298 33468 8304
rect 33416 7880 33468 7886
rect 33416 7822 33468 7828
rect 32876 7772 33088 7800
rect 32588 7744 32640 7750
rect 32588 7686 32640 7692
rect 32772 7744 32824 7750
rect 32772 7686 32824 7692
rect 32416 7398 32536 7426
rect 32600 7410 32628 7686
rect 32402 7304 32458 7313
rect 32402 7239 32458 7248
rect 32416 7206 32444 7239
rect 32128 7200 32180 7206
rect 32128 7142 32180 7148
rect 32404 7200 32456 7206
rect 32404 7142 32456 7148
rect 31950 7100 32258 7109
rect 31950 7098 31956 7100
rect 32012 7098 32036 7100
rect 32092 7098 32116 7100
rect 32172 7098 32196 7100
rect 32252 7098 32258 7100
rect 32012 7046 32014 7098
rect 32194 7046 32196 7098
rect 31950 7044 31956 7046
rect 32012 7044 32036 7046
rect 32092 7044 32116 7046
rect 32172 7044 32196 7046
rect 32252 7044 32258 7046
rect 31950 7035 32258 7044
rect 31852 6860 31904 6866
rect 31852 6802 31904 6808
rect 32404 6792 32456 6798
rect 32404 6734 32456 6740
rect 31852 6656 31904 6662
rect 31772 6616 31852 6644
rect 31484 6598 31536 6604
rect 31852 6598 31904 6604
rect 31852 6384 31904 6390
rect 31852 6326 31904 6332
rect 31392 6316 31444 6322
rect 31392 6258 31444 6264
rect 31300 4480 31352 4486
rect 31300 4422 31352 4428
rect 30748 4004 30800 4010
rect 30748 3946 30800 3952
rect 30932 4004 30984 4010
rect 30932 3946 30984 3952
rect 30656 3732 30708 3738
rect 30656 3674 30708 3680
rect 31208 3528 31260 3534
rect 31208 3470 31260 3476
rect 31220 2106 31248 3470
rect 31312 2553 31340 4422
rect 31298 2544 31354 2553
rect 31298 2479 31354 2488
rect 31208 2100 31260 2106
rect 31208 2042 31260 2048
rect 30286 1864 30342 1873
rect 30286 1799 30342 1808
rect 29920 60 29972 66
rect 15750 0 15806 40
rect 17314 0 17370 56
rect 18878 0 18934 56
rect 20442 0 20498 56
rect 22006 0 22062 56
rect 23570 0 23626 56
rect 25134 0 25190 56
rect 26698 0 26754 56
rect 28262 0 28318 56
rect 29826 0 29882 56
rect 31404 56 31432 6258
rect 31864 5846 31892 6326
rect 31950 6012 32258 6021
rect 31950 6010 31956 6012
rect 32012 6010 32036 6012
rect 32092 6010 32116 6012
rect 32172 6010 32196 6012
rect 32252 6010 32258 6012
rect 32012 5958 32014 6010
rect 32194 5958 32196 6010
rect 31950 5956 31956 5958
rect 32012 5956 32036 5958
rect 32092 5956 32116 5958
rect 32172 5956 32196 5958
rect 32252 5956 32258 5958
rect 31950 5947 32258 5956
rect 31852 5840 31904 5846
rect 31852 5782 31904 5788
rect 32416 5778 32444 6734
rect 32404 5772 32456 5778
rect 32404 5714 32456 5720
rect 31668 5568 31720 5574
rect 31668 5510 31720 5516
rect 31576 5228 31628 5234
rect 31576 5170 31628 5176
rect 31588 134 31616 5170
rect 31576 128 31628 134
rect 31680 105 31708 5510
rect 32508 5370 32536 7398
rect 32588 7404 32640 7410
rect 32588 7346 32640 7352
rect 32588 7200 32640 7206
rect 32588 7142 32640 7148
rect 32496 5364 32548 5370
rect 32496 5306 32548 5312
rect 31950 4924 32258 4933
rect 31950 4922 31956 4924
rect 32012 4922 32036 4924
rect 32092 4922 32116 4924
rect 32172 4922 32196 4924
rect 32252 4922 32258 4924
rect 32012 4870 32014 4922
rect 32194 4870 32196 4922
rect 31950 4868 31956 4870
rect 32012 4868 32036 4870
rect 32092 4868 32116 4870
rect 32172 4868 32196 4870
rect 32252 4868 32258 4870
rect 31950 4859 32258 4868
rect 32600 4214 32628 7142
rect 32784 6225 32812 7686
rect 32770 6216 32826 6225
rect 32770 6151 32826 6160
rect 32772 5704 32824 5710
rect 32772 5646 32824 5652
rect 32588 4208 32640 4214
rect 32588 4150 32640 4156
rect 31950 3836 32258 3845
rect 31950 3834 31956 3836
rect 32012 3834 32036 3836
rect 32092 3834 32116 3836
rect 32172 3834 32196 3836
rect 32252 3834 32258 3836
rect 32012 3782 32014 3834
rect 32194 3782 32196 3834
rect 31950 3780 31956 3782
rect 32012 3780 32036 3782
rect 32092 3780 32116 3782
rect 32172 3780 32196 3782
rect 32252 3780 32258 3782
rect 31950 3771 32258 3780
rect 31950 2748 32258 2757
rect 31950 2746 31956 2748
rect 32012 2746 32036 2748
rect 32092 2746 32116 2748
rect 32172 2746 32196 2748
rect 32252 2746 32258 2748
rect 32012 2694 32014 2746
rect 32194 2694 32196 2746
rect 31950 2692 31956 2694
rect 32012 2692 32036 2694
rect 32092 2692 32116 2694
rect 32172 2692 32196 2694
rect 32252 2692 32258 2694
rect 31950 2683 32258 2692
rect 31576 70 31628 76
rect 31666 96 31722 105
rect 29920 2 29972 8
rect 31390 0 31446 56
rect 31666 31 31722 40
rect 32784 42 32812 5646
rect 32876 4826 32904 7772
rect 33010 7644 33318 7653
rect 33010 7642 33016 7644
rect 33072 7642 33096 7644
rect 33152 7642 33176 7644
rect 33232 7642 33256 7644
rect 33312 7642 33318 7644
rect 33072 7590 33074 7642
rect 33254 7590 33256 7642
rect 33010 7588 33016 7590
rect 33072 7588 33096 7590
rect 33152 7588 33176 7590
rect 33232 7588 33256 7590
rect 33312 7588 33318 7590
rect 33010 7579 33318 7588
rect 33010 6556 33318 6565
rect 33010 6554 33016 6556
rect 33072 6554 33096 6556
rect 33152 6554 33176 6556
rect 33232 6554 33256 6556
rect 33312 6554 33318 6556
rect 33072 6502 33074 6554
rect 33254 6502 33256 6554
rect 33010 6500 33016 6502
rect 33072 6500 33096 6502
rect 33152 6500 33176 6502
rect 33232 6500 33256 6502
rect 33312 6500 33318 6502
rect 33010 6491 33318 6500
rect 33010 5468 33318 5477
rect 33010 5466 33016 5468
rect 33072 5466 33096 5468
rect 33152 5466 33176 5468
rect 33232 5466 33256 5468
rect 33312 5466 33318 5468
rect 33072 5414 33074 5466
rect 33254 5414 33256 5466
rect 33010 5412 33016 5414
rect 33072 5412 33096 5414
rect 33152 5412 33176 5414
rect 33232 5412 33256 5414
rect 33312 5412 33318 5414
rect 33010 5403 33318 5412
rect 32864 4820 32916 4826
rect 32864 4762 32916 4768
rect 33010 4380 33318 4389
rect 33010 4378 33016 4380
rect 33072 4378 33096 4380
rect 33152 4378 33176 4380
rect 33232 4378 33256 4380
rect 33312 4378 33318 4380
rect 33072 4326 33074 4378
rect 33254 4326 33256 4378
rect 33010 4324 33016 4326
rect 33072 4324 33096 4326
rect 33152 4324 33176 4326
rect 33232 4324 33256 4326
rect 33312 4324 33318 4326
rect 33010 4315 33318 4324
rect 33428 3738 33456 7822
rect 33520 4486 33548 8434
rect 33888 8378 33916 11194
rect 34060 8492 34112 8498
rect 34060 8434 34112 8440
rect 33888 8362 34008 8378
rect 33888 8356 34020 8362
rect 33888 8350 33968 8356
rect 33968 8298 34020 8304
rect 34072 5846 34100 8434
rect 34164 8430 34192 11194
rect 34152 8424 34204 8430
rect 34152 8366 34204 8372
rect 34440 8090 34468 11194
rect 34716 8634 34744 11194
rect 34992 8838 35020 11194
rect 35072 8900 35124 8906
rect 35072 8842 35124 8848
rect 34980 8832 35032 8838
rect 34980 8774 35032 8780
rect 34704 8628 34756 8634
rect 34704 8570 34756 8576
rect 35084 8498 35112 8842
rect 35268 8498 35296 11194
rect 34704 8492 34756 8498
rect 34704 8434 34756 8440
rect 35072 8492 35124 8498
rect 35072 8434 35124 8440
rect 35256 8492 35308 8498
rect 35256 8434 35308 8440
rect 34428 8084 34480 8090
rect 34428 8026 34480 8032
rect 34242 7440 34298 7449
rect 34242 7375 34244 7384
rect 34296 7375 34298 7384
rect 34244 7346 34296 7352
rect 34716 6662 34744 8434
rect 35544 8090 35572 11194
rect 35624 8832 35676 8838
rect 35624 8774 35676 8780
rect 35636 8362 35664 8774
rect 35820 8634 35848 11194
rect 35808 8628 35860 8634
rect 35808 8570 35860 8576
rect 35900 8560 35952 8566
rect 35820 8508 35900 8514
rect 35820 8502 35952 8508
rect 35716 8492 35768 8498
rect 35716 8434 35768 8440
rect 35820 8486 35940 8502
rect 35624 8356 35676 8362
rect 35624 8298 35676 8304
rect 35532 8084 35584 8090
rect 35532 8026 35584 8032
rect 35624 7880 35676 7886
rect 35624 7822 35676 7828
rect 35636 6730 35664 7822
rect 35624 6724 35676 6730
rect 35624 6666 35676 6672
rect 34704 6656 34756 6662
rect 34704 6598 34756 6604
rect 35256 6248 35308 6254
rect 35256 6190 35308 6196
rect 35268 5914 35296 6190
rect 35256 5908 35308 5914
rect 35256 5850 35308 5856
rect 34060 5840 34112 5846
rect 34060 5782 34112 5788
rect 34612 5636 34664 5642
rect 34612 5578 34664 5584
rect 33508 4480 33560 4486
rect 33508 4422 33560 4428
rect 33416 3732 33468 3738
rect 33416 3674 33468 3680
rect 34520 3460 34572 3466
rect 34520 3402 34572 3408
rect 33010 3292 33318 3301
rect 33010 3290 33016 3292
rect 33072 3290 33096 3292
rect 33152 3290 33176 3292
rect 33232 3290 33256 3292
rect 33312 3290 33318 3292
rect 33072 3238 33074 3290
rect 33254 3238 33256 3290
rect 33010 3236 33016 3238
rect 33072 3236 33096 3238
rect 33152 3236 33176 3238
rect 33232 3236 33256 3238
rect 33312 3236 33318 3238
rect 33010 3227 33318 3236
rect 33010 2204 33318 2213
rect 33010 2202 33016 2204
rect 33072 2202 33096 2204
rect 33152 2202 33176 2204
rect 33232 2202 33256 2204
rect 33312 2202 33318 2204
rect 33072 2150 33074 2202
rect 33254 2150 33256 2202
rect 33010 2148 33016 2150
rect 33072 2148 33096 2150
rect 33152 2148 33176 2150
rect 33232 2148 33256 2150
rect 33312 2148 33318 2150
rect 33010 2139 33318 2148
rect 34532 2009 34560 3402
rect 34518 2000 34574 2009
rect 34518 1935 34574 1944
rect 34624 1850 34652 5578
rect 35728 3738 35756 8434
rect 35820 6186 35848 8486
rect 36096 8090 36124 11194
rect 36176 8492 36228 8498
rect 36176 8434 36228 8440
rect 36084 8084 36136 8090
rect 36084 8026 36136 8032
rect 36188 7970 36216 8434
rect 36372 8430 36400 11194
rect 36544 8492 36596 8498
rect 36544 8434 36596 8440
rect 36360 8424 36412 8430
rect 36360 8366 36412 8372
rect 36096 7942 36216 7970
rect 35900 7472 35952 7478
rect 35900 7414 35952 7420
rect 35912 6769 35940 7414
rect 35992 7200 36044 7206
rect 35992 7142 36044 7148
rect 35898 6760 35954 6769
rect 35898 6695 35954 6704
rect 35808 6180 35860 6186
rect 35808 6122 35860 6128
rect 36004 5681 36032 7142
rect 35990 5672 36046 5681
rect 35990 5607 36046 5616
rect 36096 5386 36124 7942
rect 36176 7880 36228 7886
rect 36176 7822 36228 7828
rect 36188 7546 36216 7822
rect 36176 7540 36228 7546
rect 36176 7482 36228 7488
rect 36268 7540 36320 7546
rect 36268 7482 36320 7488
rect 36004 5358 36124 5386
rect 36004 5098 36032 5358
rect 36084 5228 36136 5234
rect 36084 5170 36136 5176
rect 35992 5092 36044 5098
rect 35992 5034 36044 5040
rect 35716 3732 35768 3738
rect 35716 3674 35768 3680
rect 35808 3528 35860 3534
rect 35808 3470 35860 3476
rect 35348 3392 35400 3398
rect 35348 3334 35400 3340
rect 35360 2990 35388 3334
rect 35348 2984 35400 2990
rect 35348 2926 35400 2932
rect 35820 2582 35848 3470
rect 35808 2576 35860 2582
rect 35808 2518 35860 2524
rect 34532 1822 34652 1850
rect 32876 56 32996 82
rect 34532 56 34560 1822
rect 36096 56 36124 5170
rect 36280 5166 36308 7482
rect 36556 7274 36584 8434
rect 36648 8090 36676 11194
rect 36924 8634 36952 11194
rect 37094 8936 37150 8945
rect 37094 8871 37150 8880
rect 36912 8628 36964 8634
rect 36912 8570 36964 8576
rect 36912 8424 36964 8430
rect 36912 8366 36964 8372
rect 36636 8084 36688 8090
rect 36636 8026 36688 8032
rect 36728 7880 36780 7886
rect 36728 7822 36780 7828
rect 36544 7268 36596 7274
rect 36544 7210 36596 7216
rect 36740 5914 36768 7822
rect 36924 5914 36952 8366
rect 37108 6866 37136 8871
rect 37200 8362 37228 11194
rect 37370 9072 37426 9081
rect 37370 9007 37426 9016
rect 37188 8356 37240 8362
rect 37188 8298 37240 8304
rect 37280 7812 37332 7818
rect 37280 7754 37332 7760
rect 37096 6860 37148 6866
rect 37096 6802 37148 6808
rect 37292 6118 37320 7754
rect 37384 7410 37412 9007
rect 37476 8566 37504 11194
rect 37464 8560 37516 8566
rect 37464 8502 37516 8508
rect 37752 8090 37780 11194
rect 38290 9888 38346 9897
rect 38290 9823 38346 9832
rect 37832 8492 37884 8498
rect 37832 8434 37884 8440
rect 37740 8084 37792 8090
rect 37740 8026 37792 8032
rect 37464 8016 37516 8022
rect 37844 7970 37872 8434
rect 37950 8188 38258 8197
rect 37950 8186 37956 8188
rect 38012 8186 38036 8188
rect 38092 8186 38116 8188
rect 38172 8186 38196 8188
rect 38252 8186 38258 8188
rect 38012 8134 38014 8186
rect 38194 8134 38196 8186
rect 37950 8132 37956 8134
rect 38012 8132 38036 8134
rect 38092 8132 38116 8134
rect 38172 8132 38196 8134
rect 38252 8132 38258 8134
rect 37950 8123 38258 8132
rect 37464 7958 37516 7964
rect 37372 7404 37424 7410
rect 37372 7346 37424 7352
rect 37476 6322 37504 7958
rect 37752 7942 37872 7970
rect 37556 7404 37608 7410
rect 37556 7346 37608 7352
rect 37568 7002 37596 7346
rect 37556 6996 37608 7002
rect 37556 6938 37608 6944
rect 37648 6928 37700 6934
rect 37648 6870 37700 6876
rect 37464 6316 37516 6322
rect 37464 6258 37516 6264
rect 37280 6112 37332 6118
rect 37280 6054 37332 6060
rect 37660 5914 37688 6870
rect 36728 5908 36780 5914
rect 36728 5850 36780 5856
rect 36912 5908 36964 5914
rect 36912 5850 36964 5856
rect 37648 5908 37700 5914
rect 37648 5850 37700 5856
rect 37752 5370 37780 7942
rect 37832 7880 37884 7886
rect 37832 7822 37884 7828
rect 37740 5364 37792 5370
rect 37740 5306 37792 5312
rect 37648 5228 37700 5234
rect 37648 5170 37700 5176
rect 36268 5160 36320 5166
rect 36268 5102 36320 5108
rect 37464 3596 37516 3602
rect 37464 3538 37516 3544
rect 37372 3392 37424 3398
rect 37372 3334 37424 3340
rect 37384 2446 37412 3334
rect 37372 2440 37424 2446
rect 37372 2382 37424 2388
rect 37476 1737 37504 3538
rect 37556 2576 37608 2582
rect 37554 2544 37556 2553
rect 37608 2544 37610 2553
rect 37554 2479 37610 2488
rect 37462 1728 37518 1737
rect 37462 1663 37518 1672
rect 37660 56 37688 5170
rect 37844 4826 37872 7822
rect 38304 7546 38332 9823
rect 39578 9616 39634 9625
rect 39578 9551 39634 9560
rect 38750 9344 38806 9353
rect 38750 9279 38806 9288
rect 38658 8528 38714 8537
rect 38384 8492 38436 8498
rect 38658 8463 38714 8472
rect 38384 8434 38436 8440
rect 38292 7540 38344 7546
rect 38292 7482 38344 7488
rect 37950 7100 38258 7109
rect 37950 7098 37956 7100
rect 38012 7098 38036 7100
rect 38092 7098 38116 7100
rect 38172 7098 38196 7100
rect 38252 7098 38258 7100
rect 38012 7046 38014 7098
rect 38194 7046 38196 7098
rect 37950 7044 37956 7046
rect 38012 7044 38036 7046
rect 38092 7044 38116 7046
rect 38172 7044 38196 7046
rect 38252 7044 38258 7046
rect 37950 7035 38258 7044
rect 38292 6860 38344 6866
rect 38292 6802 38344 6808
rect 37950 6012 38258 6021
rect 37950 6010 37956 6012
rect 38012 6010 38036 6012
rect 38092 6010 38116 6012
rect 38172 6010 38196 6012
rect 38252 6010 38258 6012
rect 38012 5958 38014 6010
rect 38194 5958 38196 6010
rect 37950 5956 37956 5958
rect 38012 5956 38036 5958
rect 38092 5956 38116 5958
rect 38172 5956 38196 5958
rect 38252 5956 38258 5958
rect 37950 5947 38258 5956
rect 37950 4924 38258 4933
rect 37950 4922 37956 4924
rect 38012 4922 38036 4924
rect 38092 4922 38116 4924
rect 38172 4922 38196 4924
rect 38252 4922 38258 4924
rect 38012 4870 38014 4922
rect 38194 4870 38196 4922
rect 37950 4868 37956 4870
rect 38012 4868 38036 4870
rect 38092 4868 38116 4870
rect 38172 4868 38196 4870
rect 38252 4868 38258 4870
rect 37950 4859 38258 4868
rect 37832 4820 37884 4826
rect 37832 4762 37884 4768
rect 38304 4690 38332 6802
rect 38396 5370 38424 8434
rect 38672 8090 38700 8463
rect 38660 8084 38712 8090
rect 38660 8026 38712 8032
rect 38764 7546 38792 9279
rect 39486 8800 39542 8809
rect 39010 8732 39318 8741
rect 39486 8735 39542 8744
rect 39010 8730 39016 8732
rect 39072 8730 39096 8732
rect 39152 8730 39176 8732
rect 39232 8730 39256 8732
rect 39312 8730 39318 8732
rect 39072 8678 39074 8730
rect 39254 8678 39256 8730
rect 39010 8676 39016 8678
rect 39072 8676 39096 8678
rect 39152 8676 39176 8678
rect 39232 8676 39256 8678
rect 39312 8676 39318 8678
rect 39010 8667 39318 8676
rect 39026 8392 39082 8401
rect 39026 8327 39028 8336
rect 39080 8327 39082 8336
rect 39396 8356 39448 8362
rect 39028 8298 39080 8304
rect 39396 8298 39448 8304
rect 39408 7993 39436 8298
rect 39394 7984 39450 7993
rect 39394 7919 39450 7928
rect 38936 7744 38988 7750
rect 39396 7744 39448 7750
rect 38936 7686 38988 7692
rect 39394 7712 39396 7721
rect 39448 7712 39450 7721
rect 38752 7540 38804 7546
rect 38752 7482 38804 7488
rect 38948 7449 38976 7686
rect 39010 7644 39318 7653
rect 39394 7647 39450 7656
rect 39010 7642 39016 7644
rect 39072 7642 39096 7644
rect 39152 7642 39176 7644
rect 39232 7642 39256 7644
rect 39312 7642 39318 7644
rect 39072 7590 39074 7642
rect 39254 7590 39256 7642
rect 39010 7588 39016 7590
rect 39072 7588 39096 7590
rect 39152 7588 39176 7590
rect 39232 7588 39256 7590
rect 39312 7588 39318 7590
rect 39010 7579 39318 7588
rect 39500 7546 39528 8735
rect 39488 7540 39540 7546
rect 39488 7482 39540 7488
rect 38934 7440 38990 7449
rect 38844 7404 38896 7410
rect 38934 7375 38990 7384
rect 39028 7404 39080 7410
rect 38844 7346 38896 7352
rect 39028 7346 39080 7352
rect 38856 7206 38884 7346
rect 38936 7336 38988 7342
rect 38936 7278 38988 7284
rect 38844 7200 38896 7206
rect 38844 7142 38896 7148
rect 38476 6792 38528 6798
rect 38476 6734 38528 6740
rect 38752 6792 38804 6798
rect 38752 6734 38804 6740
rect 38488 6458 38516 6734
rect 38568 6656 38620 6662
rect 38568 6598 38620 6604
rect 38660 6656 38712 6662
rect 38660 6598 38712 6604
rect 38476 6452 38528 6458
rect 38476 6394 38528 6400
rect 38580 5710 38608 6598
rect 38672 6361 38700 6598
rect 38764 6390 38792 6734
rect 38844 6656 38896 6662
rect 38844 6598 38896 6604
rect 38752 6384 38804 6390
rect 38658 6352 38714 6361
rect 38752 6326 38804 6332
rect 38658 6287 38714 6296
rect 38660 6112 38712 6118
rect 38660 6054 38712 6060
rect 38568 5704 38620 5710
rect 38568 5646 38620 5652
rect 38384 5364 38436 5370
rect 38384 5306 38436 5312
rect 38672 4690 38700 6054
rect 38752 5568 38804 5574
rect 38752 5510 38804 5516
rect 38292 4684 38344 4690
rect 38292 4626 38344 4632
rect 38660 4684 38712 4690
rect 38660 4626 38712 4632
rect 38764 4078 38792 5510
rect 38856 5370 38884 6598
rect 38948 5710 38976 7278
rect 39040 6866 39068 7346
rect 39488 7268 39540 7274
rect 39488 7210 39540 7216
rect 39394 7168 39450 7177
rect 39394 7103 39450 7112
rect 39028 6860 39080 6866
rect 39028 6802 39080 6808
rect 39408 6662 39436 7103
rect 39500 6905 39528 7210
rect 39486 6896 39542 6905
rect 39486 6831 39542 6840
rect 39592 6730 39620 9551
rect 40038 9072 40094 9081
rect 40038 9007 40094 9016
rect 39854 8256 39910 8265
rect 39854 8191 39910 8200
rect 39868 7478 39896 8191
rect 39856 7472 39908 7478
rect 39856 7414 39908 7420
rect 39580 6724 39632 6730
rect 39580 6666 39632 6672
rect 39396 6656 39448 6662
rect 39396 6598 39448 6604
rect 39578 6624 39634 6633
rect 39010 6556 39318 6565
rect 39578 6559 39634 6568
rect 39010 6554 39016 6556
rect 39072 6554 39096 6556
rect 39152 6554 39176 6556
rect 39232 6554 39256 6556
rect 39312 6554 39318 6556
rect 39072 6502 39074 6554
rect 39254 6502 39256 6554
rect 39010 6500 39016 6502
rect 39072 6500 39096 6502
rect 39152 6500 39176 6502
rect 39232 6500 39256 6502
rect 39312 6500 39318 6502
rect 39010 6491 39318 6500
rect 39212 6316 39264 6322
rect 39212 6258 39264 6264
rect 39028 6112 39080 6118
rect 39026 6080 39028 6089
rect 39080 6080 39082 6089
rect 39026 6015 39082 6024
rect 39224 5817 39252 6258
rect 39592 5914 39620 6559
rect 40052 6458 40080 9007
rect 40040 6452 40092 6458
rect 40040 6394 40092 6400
rect 39580 5908 39632 5914
rect 39580 5850 39632 5856
rect 39210 5808 39266 5817
rect 39210 5743 39266 5752
rect 39486 5808 39542 5817
rect 39486 5743 39542 5752
rect 38936 5704 38988 5710
rect 38936 5646 38988 5652
rect 39304 5568 39356 5574
rect 39356 5545 39436 5556
rect 39356 5536 39450 5545
rect 39356 5528 39394 5536
rect 39304 5510 39356 5516
rect 39010 5468 39318 5477
rect 39394 5471 39450 5480
rect 39010 5466 39016 5468
rect 39072 5466 39096 5468
rect 39152 5466 39176 5468
rect 39232 5466 39256 5468
rect 39312 5466 39318 5468
rect 39072 5414 39074 5466
rect 39254 5414 39256 5466
rect 39010 5412 39016 5414
rect 39072 5412 39096 5414
rect 39152 5412 39176 5414
rect 39232 5412 39256 5414
rect 39312 5412 39318 5414
rect 39010 5403 39318 5412
rect 39500 5370 39528 5743
rect 38844 5364 38896 5370
rect 38844 5306 38896 5312
rect 39488 5364 39540 5370
rect 39488 5306 39540 5312
rect 39210 5264 39266 5273
rect 38844 5228 38896 5234
rect 39210 5199 39212 5208
rect 38844 5170 38896 5176
rect 39264 5199 39266 5208
rect 39394 5264 39450 5273
rect 39394 5199 39450 5208
rect 39212 5170 39264 5176
rect 38856 4758 38884 5170
rect 39028 5024 39080 5030
rect 39026 4992 39028 5001
rect 39080 4992 39082 5001
rect 39026 4927 39082 4936
rect 39408 4826 39436 5199
rect 39396 4820 39448 4826
rect 39396 4762 39448 4768
rect 38844 4752 38896 4758
rect 38844 4694 38896 4700
rect 39486 4720 39542 4729
rect 39486 4655 39542 4664
rect 38936 4616 38988 4622
rect 38936 4558 38988 4564
rect 38844 4140 38896 4146
rect 38844 4082 38896 4088
rect 38752 4072 38804 4078
rect 38856 4049 38884 4082
rect 38752 4014 38804 4020
rect 38842 4040 38898 4049
rect 38842 3975 38898 3984
rect 37950 3836 38258 3845
rect 37950 3834 37956 3836
rect 38012 3834 38036 3836
rect 38092 3834 38116 3836
rect 38172 3834 38196 3836
rect 38252 3834 38258 3836
rect 38012 3782 38014 3834
rect 38194 3782 38196 3834
rect 37950 3780 37956 3782
rect 38012 3780 38036 3782
rect 38092 3780 38116 3782
rect 38172 3780 38196 3782
rect 38252 3780 38258 3782
rect 37950 3771 38258 3780
rect 38384 3664 38436 3670
rect 38384 3606 38436 3612
rect 37740 3392 37792 3398
rect 37740 3334 37792 3340
rect 38292 3392 38344 3398
rect 38292 3334 38344 3340
rect 37752 1465 37780 3334
rect 37950 2748 38258 2757
rect 37950 2746 37956 2748
rect 38012 2746 38036 2748
rect 38092 2746 38116 2748
rect 38172 2746 38196 2748
rect 38252 2746 38258 2748
rect 38012 2694 38014 2746
rect 38194 2694 38196 2746
rect 37950 2692 37956 2694
rect 38012 2692 38036 2694
rect 38092 2692 38116 2694
rect 38172 2692 38196 2694
rect 38252 2692 38258 2694
rect 37950 2683 38258 2692
rect 38304 2514 38332 3334
rect 38292 2508 38344 2514
rect 38292 2450 38344 2456
rect 38396 2446 38424 3606
rect 38842 3496 38898 3505
rect 38842 3431 38898 3440
rect 38660 3392 38712 3398
rect 38660 3334 38712 3340
rect 38476 3052 38528 3058
rect 38476 2994 38528 3000
rect 38488 2961 38516 2994
rect 38474 2952 38530 2961
rect 38474 2887 38530 2896
rect 38672 2774 38700 3334
rect 38856 3058 38884 3431
rect 38844 3052 38896 3058
rect 38844 2994 38896 3000
rect 38844 2848 38896 2854
rect 38842 2816 38844 2825
rect 38896 2816 38898 2825
rect 38672 2746 38792 2774
rect 38842 2751 38898 2760
rect 38764 2446 38792 2746
rect 38948 2650 38976 4558
rect 39304 4480 39356 4486
rect 39356 4457 39436 4468
rect 39356 4448 39450 4457
rect 39356 4440 39394 4448
rect 39304 4422 39356 4428
rect 39010 4380 39318 4389
rect 39394 4383 39450 4392
rect 39010 4378 39016 4380
rect 39072 4378 39096 4380
rect 39152 4378 39176 4380
rect 39232 4378 39256 4380
rect 39312 4378 39318 4380
rect 39072 4326 39074 4378
rect 39254 4326 39256 4378
rect 39010 4324 39016 4326
rect 39072 4324 39096 4326
rect 39152 4324 39176 4326
rect 39232 4324 39256 4326
rect 39312 4324 39318 4326
rect 39010 4315 39318 4324
rect 39394 4176 39450 4185
rect 39394 4111 39450 4120
rect 39028 3936 39080 3942
rect 39026 3904 39028 3913
rect 39080 3904 39082 3913
rect 39026 3839 39082 3848
rect 39408 3738 39436 4111
rect 39500 4010 39528 4655
rect 39580 4548 39632 4554
rect 39580 4490 39632 4496
rect 39488 4004 39540 4010
rect 39488 3946 39540 3952
rect 39396 3732 39448 3738
rect 39396 3674 39448 3680
rect 39210 3632 39266 3641
rect 39210 3567 39266 3576
rect 39486 3632 39542 3641
rect 39486 3567 39542 3576
rect 39224 3534 39252 3567
rect 39212 3528 39264 3534
rect 39212 3470 39264 3476
rect 39394 3360 39450 3369
rect 39010 3292 39318 3301
rect 39394 3295 39450 3304
rect 39010 3290 39016 3292
rect 39072 3290 39096 3292
rect 39152 3290 39176 3292
rect 39232 3290 39256 3292
rect 39312 3290 39318 3292
rect 39072 3238 39074 3290
rect 39254 3238 39256 3290
rect 39010 3236 39016 3238
rect 39072 3236 39096 3238
rect 39152 3236 39176 3238
rect 39232 3236 39256 3238
rect 39312 3236 39318 3238
rect 39010 3227 39318 3236
rect 39408 3194 39436 3295
rect 39396 3188 39448 3194
rect 39396 3130 39448 3136
rect 39210 3088 39266 3097
rect 39210 3023 39212 3032
rect 39264 3023 39266 3032
rect 39394 3088 39450 3097
rect 39394 3023 39450 3032
rect 39212 2994 39264 3000
rect 39408 2650 39436 3023
rect 39500 2922 39528 3567
rect 39488 2916 39540 2922
rect 39488 2858 39540 2864
rect 38936 2644 38988 2650
rect 38936 2586 38988 2592
rect 39396 2644 39448 2650
rect 39396 2586 39448 2592
rect 38384 2440 38436 2446
rect 38384 2382 38436 2388
rect 38752 2440 38804 2446
rect 38752 2382 38804 2388
rect 37832 2304 37884 2310
rect 37832 2246 37884 2252
rect 38292 2304 38344 2310
rect 38292 2246 38344 2252
rect 38660 2304 38712 2310
rect 38660 2246 38712 2252
rect 37844 2009 37872 2246
rect 37830 2000 37886 2009
rect 37830 1935 37886 1944
rect 38304 1737 38332 2246
rect 38290 1728 38346 1737
rect 38290 1663 38346 1672
rect 38672 1465 38700 2246
rect 39010 2204 39318 2213
rect 39010 2202 39016 2204
rect 39072 2202 39096 2204
rect 39152 2202 39176 2204
rect 39232 2202 39256 2204
rect 39312 2202 39318 2204
rect 39072 2150 39074 2202
rect 39254 2150 39256 2202
rect 39010 2148 39016 2150
rect 39072 2148 39096 2150
rect 39152 2148 39176 2150
rect 39232 2148 39256 2150
rect 39312 2148 39318 2150
rect 39010 2139 39318 2148
rect 37738 1456 37794 1465
rect 37738 1391 37794 1400
rect 38658 1456 38714 1465
rect 38658 1391 38714 1400
rect 39224 56 39344 82
rect 32876 54 33010 56
rect 32876 42 32904 54
rect 32784 14 32904 42
rect 32954 0 33010 54
rect 34518 0 34574 56
rect 36082 0 36138 56
rect 37646 0 37702 56
rect 39210 54 39344 56
rect 39210 0 39266 54
rect 39316 42 39344 54
rect 39592 42 39620 4490
rect 39948 2576 40000 2582
rect 39948 2518 40000 2524
rect 39960 2281 39988 2518
rect 39946 2272 40002 2281
rect 39946 2207 40002 2216
rect 39316 14 39620 42
<< via2 >>
rect 1122 9832 1178 9888
rect 1030 9560 1086 9616
rect 846 9288 902 9344
rect 570 7928 626 7984
rect 570 7384 626 7440
rect 938 8744 994 8800
rect 754 7656 810 7712
rect 1214 9016 1270 9072
rect 1122 8336 1178 8392
rect 1030 8200 1086 8256
rect 754 7112 810 7168
rect 1306 8508 1308 8528
rect 1308 8508 1360 8528
rect 1360 8508 1362 8528
rect 1306 8472 1362 8508
rect 3016 8730 3072 8732
rect 3096 8730 3152 8732
rect 3176 8730 3232 8732
rect 3256 8730 3312 8732
rect 3016 8678 3062 8730
rect 3062 8678 3072 8730
rect 3096 8678 3126 8730
rect 3126 8678 3138 8730
rect 3138 8678 3152 8730
rect 3176 8678 3190 8730
rect 3190 8678 3202 8730
rect 3202 8678 3232 8730
rect 3256 8678 3266 8730
rect 3266 8678 3312 8730
rect 3016 8676 3072 8678
rect 3096 8676 3152 8678
rect 3176 8676 3232 8678
rect 3256 8676 3312 8678
rect 1956 8186 2012 8188
rect 2036 8186 2092 8188
rect 2116 8186 2172 8188
rect 2196 8186 2252 8188
rect 1956 8134 2002 8186
rect 2002 8134 2012 8186
rect 2036 8134 2066 8186
rect 2066 8134 2078 8186
rect 2078 8134 2092 8186
rect 2116 8134 2130 8186
rect 2130 8134 2142 8186
rect 2142 8134 2172 8186
rect 2196 8134 2206 8186
rect 2206 8134 2252 8186
rect 1956 8132 2012 8134
rect 2036 8132 2092 8134
rect 2116 8132 2172 8134
rect 2196 8132 2252 8134
rect 1306 7928 1362 7984
rect 938 6840 994 6896
rect 570 6568 626 6624
rect 1214 5480 1270 5536
rect 3606 9152 3662 9208
rect 3016 7642 3072 7644
rect 3096 7642 3152 7644
rect 3176 7642 3232 7644
rect 3256 7642 3312 7644
rect 3016 7590 3062 7642
rect 3062 7590 3072 7642
rect 3096 7590 3126 7642
rect 3126 7590 3138 7642
rect 3138 7590 3152 7642
rect 3176 7590 3190 7642
rect 3190 7590 3202 7642
rect 3202 7590 3232 7642
rect 3256 7590 3266 7642
rect 3266 7590 3312 7642
rect 3016 7588 3072 7590
rect 3096 7588 3152 7590
rect 3176 7588 3232 7590
rect 3256 7588 3312 7590
rect 1956 7098 2012 7100
rect 2036 7098 2092 7100
rect 2116 7098 2172 7100
rect 2196 7098 2252 7100
rect 1956 7046 2002 7098
rect 2002 7046 2012 7098
rect 2036 7046 2066 7098
rect 2066 7046 2078 7098
rect 2078 7046 2092 7098
rect 2116 7046 2130 7098
rect 2130 7046 2142 7098
rect 2142 7046 2172 7098
rect 2196 7046 2206 7098
rect 2206 7046 2252 7098
rect 1956 7044 2012 7046
rect 2036 7044 2092 7046
rect 2116 7044 2172 7046
rect 2196 7044 2252 7046
rect 1956 6010 2012 6012
rect 2036 6010 2092 6012
rect 2116 6010 2172 6012
rect 2196 6010 2252 6012
rect 1956 5958 2002 6010
rect 2002 5958 2012 6010
rect 2036 5958 2066 6010
rect 2066 5958 2078 6010
rect 2078 5958 2092 6010
rect 2116 5958 2130 6010
rect 2130 5958 2142 6010
rect 2142 5958 2172 6010
rect 2196 5958 2206 6010
rect 2206 5958 2252 6010
rect 1956 5956 2012 5958
rect 2036 5956 2092 5958
rect 2116 5956 2172 5958
rect 2196 5956 2252 5958
rect 3054 6840 3110 6896
rect 3016 6554 3072 6556
rect 3096 6554 3152 6556
rect 3176 6554 3232 6556
rect 3256 6554 3312 6556
rect 3016 6502 3062 6554
rect 3062 6502 3072 6554
rect 3096 6502 3126 6554
rect 3126 6502 3138 6554
rect 3138 6502 3152 6554
rect 3176 6502 3190 6554
rect 3190 6502 3202 6554
rect 3202 6502 3232 6554
rect 3256 6502 3266 6554
rect 3266 6502 3312 6554
rect 3016 6500 3072 6502
rect 3096 6500 3152 6502
rect 3176 6500 3232 6502
rect 3256 6500 3312 6502
rect 2870 6296 2926 6352
rect 3422 6160 3478 6216
rect 2778 5072 2834 5128
rect 1956 4922 2012 4924
rect 2036 4922 2092 4924
rect 2116 4922 2172 4924
rect 2196 4922 2252 4924
rect 1956 4870 2002 4922
rect 2002 4870 2012 4922
rect 2036 4870 2066 4922
rect 2066 4870 2078 4922
rect 2078 4870 2092 4922
rect 2116 4870 2130 4922
rect 2130 4870 2142 4922
rect 2142 4870 2172 4922
rect 2196 4870 2206 4922
rect 2206 4870 2252 4922
rect 1956 4868 2012 4870
rect 2036 4868 2092 4870
rect 2116 4868 2172 4870
rect 2196 4868 2252 4870
rect 1306 4664 1362 4720
rect 662 4120 718 4176
rect 1956 3834 2012 3836
rect 2036 3834 2092 3836
rect 2116 3834 2172 3836
rect 2196 3834 2252 3836
rect 1956 3782 2002 3834
rect 2002 3782 2012 3834
rect 2036 3782 2066 3834
rect 2066 3782 2078 3834
rect 2078 3782 2092 3834
rect 2116 3782 2130 3834
rect 2130 3782 2142 3834
rect 2142 3782 2172 3834
rect 2196 3782 2206 3834
rect 2206 3782 2252 3834
rect 1956 3780 2012 3782
rect 2036 3780 2092 3782
rect 2116 3780 2172 3782
rect 2196 3780 2252 3782
rect 3016 5466 3072 5468
rect 3096 5466 3152 5468
rect 3176 5466 3232 5468
rect 3256 5466 3312 5468
rect 3016 5414 3062 5466
rect 3062 5414 3072 5466
rect 3096 5414 3126 5466
rect 3126 5414 3138 5466
rect 3138 5414 3152 5466
rect 3176 5414 3190 5466
rect 3190 5414 3202 5466
rect 3202 5414 3232 5466
rect 3256 5414 3266 5466
rect 3266 5414 3312 5466
rect 3016 5412 3072 5414
rect 3096 5412 3152 5414
rect 3176 5412 3232 5414
rect 3256 5412 3312 5414
rect 2870 4392 2926 4448
rect 3016 4378 3072 4380
rect 3096 4378 3152 4380
rect 3176 4378 3232 4380
rect 3256 4378 3312 4380
rect 3016 4326 3062 4378
rect 3062 4326 3072 4378
rect 3096 4326 3126 4378
rect 3126 4326 3138 4378
rect 3138 4326 3152 4378
rect 3176 4326 3190 4378
rect 3190 4326 3202 4378
rect 3202 4326 3232 4378
rect 3256 4326 3266 4378
rect 3266 4326 3312 4378
rect 3016 4324 3072 4326
rect 3096 4324 3152 4326
rect 3176 4324 3232 4326
rect 3256 4324 3312 4326
rect 2778 3576 2834 3632
rect 5630 10376 5686 10432
rect 6642 10240 6698 10296
rect 4066 5752 4122 5808
rect 4434 5208 4490 5264
rect 3422 3984 3478 4040
rect 3054 3440 3110 3496
rect 2870 3304 2926 3360
rect 3016 3290 3072 3292
rect 3096 3290 3152 3292
rect 3176 3290 3232 3292
rect 3256 3290 3312 3292
rect 3016 3238 3062 3290
rect 3062 3238 3072 3290
rect 3096 3238 3126 3290
rect 3126 3238 3138 3290
rect 3138 3238 3152 3290
rect 3176 3238 3190 3290
rect 3190 3238 3202 3290
rect 3202 3238 3232 3290
rect 3256 3238 3266 3290
rect 3266 3238 3312 3290
rect 3016 3236 3072 3238
rect 3096 3236 3152 3238
rect 3176 3236 3232 3238
rect 3256 3236 3312 3238
rect 1306 3032 1362 3088
rect 3698 4120 3754 4176
rect 3790 3032 3846 3088
rect 4066 3984 4122 4040
rect 3974 3576 4030 3632
rect 3606 2896 3662 2952
rect 3882 2896 3938 2952
rect 1956 2746 2012 2748
rect 2036 2746 2092 2748
rect 2116 2746 2172 2748
rect 2196 2746 2252 2748
rect 1956 2694 2002 2746
rect 2002 2694 2012 2746
rect 2036 2694 2066 2746
rect 2066 2694 2078 2746
rect 2078 2694 2092 2746
rect 2116 2694 2130 2746
rect 2130 2694 2142 2746
rect 2142 2694 2172 2746
rect 2196 2694 2206 2746
rect 2206 2694 2252 2746
rect 1956 2692 2012 2694
rect 2036 2692 2092 2694
rect 2116 2692 2172 2694
rect 2196 2692 2252 2694
rect 1306 2524 1308 2544
rect 1308 2524 1360 2544
rect 1360 2524 1362 2544
rect 1306 2488 1362 2524
rect 2042 2388 2044 2408
rect 2044 2388 2096 2408
rect 2096 2388 2098 2408
rect 2042 2352 2098 2388
rect 1214 1672 1270 1728
rect 2870 2216 2926 2272
rect 3016 2202 3072 2204
rect 3096 2202 3152 2204
rect 3176 2202 3232 2204
rect 3256 2202 3312 2204
rect 3016 2150 3062 2202
rect 3062 2150 3072 2202
rect 3096 2150 3126 2202
rect 3126 2150 3138 2202
rect 3138 2150 3152 2202
rect 3176 2150 3190 2202
rect 3190 2150 3202 2202
rect 3202 2150 3232 2202
rect 3256 2150 3266 2202
rect 3266 2150 3312 2202
rect 3016 2148 3072 2150
rect 3096 2148 3152 2150
rect 3176 2148 3232 2150
rect 3256 2148 3312 2150
rect 2870 1672 2926 1728
rect 6734 9968 6790 10024
rect 7654 8336 7710 8392
rect 7378 6296 7434 6352
rect 8666 9696 8722 9752
rect 7956 8186 8012 8188
rect 8036 8186 8092 8188
rect 8116 8186 8172 8188
rect 8196 8186 8252 8188
rect 7956 8134 8002 8186
rect 8002 8134 8012 8186
rect 8036 8134 8066 8186
rect 8066 8134 8078 8186
rect 8078 8134 8092 8186
rect 8116 8134 8130 8186
rect 8130 8134 8142 8186
rect 8142 8134 8172 8186
rect 8196 8134 8206 8186
rect 8206 8134 8252 8186
rect 7956 8132 8012 8134
rect 8036 8132 8092 8134
rect 8116 8132 8172 8134
rect 8196 8132 8252 8134
rect 8206 7248 8262 7304
rect 7956 7098 8012 7100
rect 8036 7098 8092 7100
rect 8116 7098 8172 7100
rect 8196 7098 8252 7100
rect 7956 7046 8002 7098
rect 8002 7046 8012 7098
rect 8036 7046 8066 7098
rect 8066 7046 8078 7098
rect 8078 7046 8092 7098
rect 8116 7046 8130 7098
rect 8130 7046 8142 7098
rect 8142 7046 8172 7098
rect 8196 7046 8206 7098
rect 8206 7046 8252 7098
rect 7956 7044 8012 7046
rect 8036 7044 8092 7046
rect 8116 7044 8172 7046
rect 8196 7044 8252 7046
rect 8390 7112 8446 7168
rect 7956 6010 8012 6012
rect 8036 6010 8092 6012
rect 8116 6010 8172 6012
rect 8196 6010 8252 6012
rect 7956 5958 8002 6010
rect 8002 5958 8012 6010
rect 8036 5958 8066 6010
rect 8066 5958 8078 6010
rect 8078 5958 8092 6010
rect 8116 5958 8130 6010
rect 8130 5958 8142 6010
rect 8142 5958 8172 6010
rect 8196 5958 8206 6010
rect 8206 5958 8252 6010
rect 7956 5956 8012 5958
rect 8036 5956 8092 5958
rect 8116 5956 8172 5958
rect 8196 5956 8252 5958
rect 9016 8730 9072 8732
rect 9096 8730 9152 8732
rect 9176 8730 9232 8732
rect 9256 8730 9312 8732
rect 9016 8678 9062 8730
rect 9062 8678 9072 8730
rect 9096 8678 9126 8730
rect 9126 8678 9138 8730
rect 9138 8678 9152 8730
rect 9176 8678 9190 8730
rect 9190 8678 9202 8730
rect 9202 8678 9232 8730
rect 9256 8678 9266 8730
rect 9266 8678 9312 8730
rect 9016 8676 9072 8678
rect 9096 8676 9152 8678
rect 9176 8676 9232 8678
rect 9256 8676 9312 8678
rect 9678 10104 9734 10160
rect 9218 7828 9220 7848
rect 9220 7828 9272 7848
rect 9272 7828 9274 7848
rect 9218 7792 9274 7828
rect 8390 5344 8446 5400
rect 7956 4922 8012 4924
rect 8036 4922 8092 4924
rect 8116 4922 8172 4924
rect 8196 4922 8252 4924
rect 7956 4870 8002 4922
rect 8002 4870 8012 4922
rect 8036 4870 8066 4922
rect 8066 4870 8078 4922
rect 8078 4870 8092 4922
rect 8116 4870 8130 4922
rect 8130 4870 8142 4922
rect 8142 4870 8172 4922
rect 8196 4870 8206 4922
rect 8206 4870 8252 4922
rect 7956 4868 8012 4870
rect 8036 4868 8092 4870
rect 8116 4868 8172 4870
rect 8196 4868 8252 4870
rect 7956 3834 8012 3836
rect 8036 3834 8092 3836
rect 8116 3834 8172 3836
rect 8196 3834 8252 3836
rect 7956 3782 8002 3834
rect 8002 3782 8012 3834
rect 8036 3782 8066 3834
rect 8066 3782 8078 3834
rect 8078 3782 8092 3834
rect 8116 3782 8130 3834
rect 8130 3782 8142 3834
rect 8142 3782 8172 3834
rect 8196 3782 8206 3834
rect 8206 3782 8252 3834
rect 7956 3780 8012 3782
rect 8036 3780 8092 3782
rect 8116 3780 8172 3782
rect 8196 3780 8252 3782
rect 9016 7642 9072 7644
rect 9096 7642 9152 7644
rect 9176 7642 9232 7644
rect 9256 7642 9312 7644
rect 9016 7590 9062 7642
rect 9062 7590 9072 7642
rect 9096 7590 9126 7642
rect 9126 7590 9138 7642
rect 9138 7590 9152 7642
rect 9176 7590 9190 7642
rect 9190 7590 9202 7642
rect 9202 7590 9232 7642
rect 9256 7590 9266 7642
rect 9266 7590 9312 7642
rect 9016 7588 9072 7590
rect 9096 7588 9152 7590
rect 9176 7588 9232 7590
rect 9256 7588 9312 7590
rect 9016 6554 9072 6556
rect 9096 6554 9152 6556
rect 9176 6554 9232 6556
rect 9256 6554 9312 6556
rect 9016 6502 9062 6554
rect 9062 6502 9072 6554
rect 9096 6502 9126 6554
rect 9126 6502 9138 6554
rect 9138 6502 9152 6554
rect 9176 6502 9190 6554
rect 9190 6502 9202 6554
rect 9202 6502 9232 6554
rect 9256 6502 9266 6554
rect 9266 6502 9312 6554
rect 9016 6500 9072 6502
rect 9096 6500 9152 6502
rect 9176 6500 9232 6502
rect 9256 6500 9312 6502
rect 9016 5466 9072 5468
rect 9096 5466 9152 5468
rect 9176 5466 9232 5468
rect 9256 5466 9312 5468
rect 9016 5414 9062 5466
rect 9062 5414 9072 5466
rect 9096 5414 9126 5466
rect 9126 5414 9138 5466
rect 9138 5414 9152 5466
rect 9176 5414 9190 5466
rect 9190 5414 9202 5466
rect 9202 5414 9232 5466
rect 9256 5414 9266 5466
rect 9266 5414 9312 5466
rect 9016 5412 9072 5414
rect 9096 5412 9152 5414
rect 9176 5412 9232 5414
rect 9256 5412 9312 5414
rect 9016 4378 9072 4380
rect 9096 4378 9152 4380
rect 9176 4378 9232 4380
rect 9256 4378 9312 4380
rect 9016 4326 9062 4378
rect 9062 4326 9072 4378
rect 9096 4326 9126 4378
rect 9126 4326 9138 4378
rect 9138 4326 9152 4378
rect 9176 4326 9190 4378
rect 9190 4326 9202 4378
rect 9202 4326 9232 4378
rect 9256 4326 9266 4378
rect 9266 4326 9312 4378
rect 9016 4324 9072 4326
rect 9096 4324 9152 4326
rect 9176 4324 9232 4326
rect 9256 4324 9312 4326
rect 10230 9424 10286 9480
rect 9586 5108 9588 5128
rect 9588 5108 9640 5128
rect 9640 5108 9642 5128
rect 9586 5072 9642 5108
rect 10782 7384 10838 7440
rect 9954 5636 10010 5672
rect 9954 5616 9956 5636
rect 9956 5616 10008 5636
rect 10008 5616 10010 5636
rect 10322 6160 10378 6216
rect 12070 4564 12072 4584
rect 12072 4564 12124 4584
rect 12124 4564 12126 4584
rect 12070 4528 12126 4564
rect 13358 9288 13414 9344
rect 12990 8492 13046 8528
rect 12990 8472 12992 8492
rect 12992 8472 13044 8492
rect 13044 8472 13046 8492
rect 13450 7520 13506 7576
rect 13450 7248 13506 7304
rect 13358 5788 13360 5808
rect 13360 5788 13412 5808
rect 13412 5788 13414 5808
rect 13358 5752 13414 5788
rect 13956 8186 14012 8188
rect 14036 8186 14092 8188
rect 14116 8186 14172 8188
rect 14196 8186 14252 8188
rect 13956 8134 14002 8186
rect 14002 8134 14012 8186
rect 14036 8134 14066 8186
rect 14066 8134 14078 8186
rect 14078 8134 14092 8186
rect 14116 8134 14130 8186
rect 14130 8134 14142 8186
rect 14142 8134 14172 8186
rect 14196 8134 14206 8186
rect 14206 8134 14252 8186
rect 13956 8132 14012 8134
rect 14036 8132 14092 8134
rect 14116 8132 14172 8134
rect 14196 8132 14252 8134
rect 14186 7520 14242 7576
rect 14278 7384 14334 7440
rect 13956 7098 14012 7100
rect 14036 7098 14092 7100
rect 14116 7098 14172 7100
rect 14196 7098 14252 7100
rect 13956 7046 14002 7098
rect 14002 7046 14012 7098
rect 14036 7046 14066 7098
rect 14066 7046 14078 7098
rect 14078 7046 14092 7098
rect 14116 7046 14130 7098
rect 14130 7046 14142 7098
rect 14142 7046 14172 7098
rect 14196 7046 14206 7098
rect 14206 7046 14252 7098
rect 13956 7044 14012 7046
rect 14036 7044 14092 7046
rect 14116 7044 14172 7046
rect 14196 7044 14252 7046
rect 14738 9832 14794 9888
rect 14646 7828 14648 7848
rect 14648 7828 14700 7848
rect 14700 7828 14702 7848
rect 14646 7792 14702 7828
rect 14370 6976 14426 7032
rect 14370 6704 14426 6760
rect 14094 6432 14150 6488
rect 13956 6010 14012 6012
rect 14036 6010 14092 6012
rect 14116 6010 14172 6012
rect 14196 6010 14252 6012
rect 13956 5958 14002 6010
rect 14002 5958 14012 6010
rect 14036 5958 14066 6010
rect 14066 5958 14078 6010
rect 14078 5958 14092 6010
rect 14116 5958 14130 6010
rect 14130 5958 14142 6010
rect 14142 5958 14172 6010
rect 14196 5958 14206 6010
rect 14206 5958 14252 6010
rect 13956 5956 14012 5958
rect 14036 5956 14092 5958
rect 14116 5956 14172 5958
rect 14196 5956 14252 5958
rect 13956 4922 14012 4924
rect 14036 4922 14092 4924
rect 14116 4922 14172 4924
rect 14196 4922 14252 4924
rect 13956 4870 14002 4922
rect 14002 4870 14012 4922
rect 14036 4870 14066 4922
rect 14066 4870 14078 4922
rect 14078 4870 14092 4922
rect 14116 4870 14130 4922
rect 14130 4870 14142 4922
rect 14142 4870 14172 4922
rect 14196 4870 14206 4922
rect 14206 4870 14252 4922
rect 13956 4868 14012 4870
rect 14036 4868 14092 4870
rect 14116 4868 14172 4870
rect 14196 4868 14252 4870
rect 13956 3834 14012 3836
rect 14036 3834 14092 3836
rect 14116 3834 14172 3836
rect 14196 3834 14252 3836
rect 13956 3782 14002 3834
rect 14002 3782 14012 3834
rect 14036 3782 14066 3834
rect 14066 3782 14078 3834
rect 14078 3782 14092 3834
rect 14116 3782 14130 3834
rect 14130 3782 14142 3834
rect 14142 3782 14172 3834
rect 14196 3782 14206 3834
rect 14206 3782 14252 3834
rect 13956 3780 14012 3782
rect 14036 3780 14092 3782
rect 14116 3780 14172 3782
rect 14196 3780 14252 3782
rect 15016 8730 15072 8732
rect 15096 8730 15152 8732
rect 15176 8730 15232 8732
rect 15256 8730 15312 8732
rect 15016 8678 15062 8730
rect 15062 8678 15072 8730
rect 15096 8678 15126 8730
rect 15126 8678 15138 8730
rect 15138 8678 15152 8730
rect 15176 8678 15190 8730
rect 15190 8678 15202 8730
rect 15202 8678 15232 8730
rect 15256 8678 15266 8730
rect 15266 8678 15312 8730
rect 15016 8676 15072 8678
rect 15096 8676 15152 8678
rect 15176 8676 15232 8678
rect 15256 8676 15312 8678
rect 14922 8200 14978 8256
rect 14738 7112 14794 7168
rect 14462 3848 14518 3904
rect 9016 3290 9072 3292
rect 9096 3290 9152 3292
rect 9176 3290 9232 3292
rect 9256 3290 9312 3292
rect 9016 3238 9062 3290
rect 9062 3238 9072 3290
rect 9096 3238 9126 3290
rect 9126 3238 9138 3290
rect 9138 3238 9152 3290
rect 9176 3238 9190 3290
rect 9190 3238 9202 3290
rect 9202 3238 9232 3290
rect 9256 3238 9266 3290
rect 9266 3238 9312 3290
rect 9016 3236 9072 3238
rect 9096 3236 9152 3238
rect 9176 3236 9232 3238
rect 9256 3236 9312 3238
rect 7956 2746 8012 2748
rect 8036 2746 8092 2748
rect 8116 2746 8172 2748
rect 8196 2746 8252 2748
rect 7956 2694 8002 2746
rect 8002 2694 8012 2746
rect 8036 2694 8066 2746
rect 8066 2694 8078 2746
rect 8078 2694 8092 2746
rect 8116 2694 8130 2746
rect 8130 2694 8142 2746
rect 8142 2694 8172 2746
rect 8196 2694 8206 2746
rect 8206 2694 8252 2746
rect 7956 2692 8012 2694
rect 8036 2692 8092 2694
rect 8116 2692 8172 2694
rect 8196 2692 8252 2694
rect 13956 2746 14012 2748
rect 14036 2746 14092 2748
rect 14116 2746 14172 2748
rect 14196 2746 14252 2748
rect 13956 2694 14002 2746
rect 14002 2694 14012 2746
rect 14036 2694 14066 2746
rect 14066 2694 14078 2746
rect 14078 2694 14092 2746
rect 14116 2694 14130 2746
rect 14130 2694 14142 2746
rect 14142 2694 14172 2746
rect 14196 2694 14206 2746
rect 14206 2694 14252 2746
rect 13956 2692 14012 2694
rect 14036 2692 14092 2694
rect 14116 2692 14172 2694
rect 14196 2692 14252 2694
rect 12622 2488 12678 2544
rect 15474 7656 15530 7712
rect 15016 7642 15072 7644
rect 15096 7642 15152 7644
rect 15176 7642 15232 7644
rect 15256 7642 15312 7644
rect 15016 7590 15062 7642
rect 15062 7590 15072 7642
rect 15096 7590 15126 7642
rect 15126 7590 15138 7642
rect 15138 7590 15152 7642
rect 15176 7590 15190 7642
rect 15190 7590 15202 7642
rect 15202 7590 15232 7642
rect 15256 7590 15266 7642
rect 15266 7590 15312 7642
rect 15016 7588 15072 7590
rect 15096 7588 15152 7590
rect 15176 7588 15232 7590
rect 15256 7588 15312 7590
rect 15474 7520 15530 7576
rect 15016 6554 15072 6556
rect 15096 6554 15152 6556
rect 15176 6554 15232 6556
rect 15256 6554 15312 6556
rect 15016 6502 15062 6554
rect 15062 6502 15072 6554
rect 15096 6502 15126 6554
rect 15126 6502 15138 6554
rect 15138 6502 15152 6554
rect 15176 6502 15190 6554
rect 15190 6502 15202 6554
rect 15202 6502 15232 6554
rect 15256 6502 15266 6554
rect 15266 6502 15312 6554
rect 15016 6500 15072 6502
rect 15096 6500 15152 6502
rect 15176 6500 15232 6502
rect 15256 6500 15312 6502
rect 15016 5466 15072 5468
rect 15096 5466 15152 5468
rect 15176 5466 15232 5468
rect 15256 5466 15312 5468
rect 15016 5414 15062 5466
rect 15062 5414 15072 5466
rect 15096 5414 15126 5466
rect 15126 5414 15138 5466
rect 15138 5414 15152 5466
rect 15176 5414 15190 5466
rect 15190 5414 15202 5466
rect 15202 5414 15232 5466
rect 15256 5414 15266 5466
rect 15266 5414 15312 5466
rect 15016 5412 15072 5414
rect 15096 5412 15152 5414
rect 15176 5412 15232 5414
rect 15256 5412 15312 5414
rect 15016 4378 15072 4380
rect 15096 4378 15152 4380
rect 15176 4378 15232 4380
rect 15256 4378 15312 4380
rect 15016 4326 15062 4378
rect 15062 4326 15072 4378
rect 15096 4326 15126 4378
rect 15126 4326 15138 4378
rect 15138 4326 15152 4378
rect 15176 4326 15190 4378
rect 15190 4326 15202 4378
rect 15202 4326 15232 4378
rect 15256 4326 15266 4378
rect 15266 4326 15312 4378
rect 15016 4324 15072 4326
rect 15096 4324 15152 4326
rect 15176 4324 15232 4326
rect 15256 4324 15312 4326
rect 16394 9016 16450 9072
rect 15750 5480 15806 5536
rect 16670 6432 16726 6488
rect 16578 3712 16634 3768
rect 17498 4664 17554 4720
rect 17130 3440 17186 3496
rect 15016 3290 15072 3292
rect 15096 3290 15152 3292
rect 15176 3290 15232 3292
rect 15256 3290 15312 3292
rect 15016 3238 15062 3290
rect 15062 3238 15072 3290
rect 15096 3238 15126 3290
rect 15126 3238 15138 3290
rect 15138 3238 15152 3290
rect 15176 3238 15190 3290
rect 15190 3238 15202 3290
rect 15202 3238 15232 3290
rect 15256 3238 15266 3290
rect 15266 3238 15312 3290
rect 15016 3236 15072 3238
rect 15096 3236 15152 3238
rect 15176 3236 15232 3238
rect 15256 3236 15312 3238
rect 17130 3032 17186 3088
rect 17314 3032 17370 3088
rect 9016 2202 9072 2204
rect 9096 2202 9152 2204
rect 9176 2202 9232 2204
rect 9256 2202 9312 2204
rect 9016 2150 9062 2202
rect 9062 2150 9072 2202
rect 9096 2150 9126 2202
rect 9126 2150 9138 2202
rect 9138 2150 9152 2202
rect 9176 2150 9190 2202
rect 9190 2150 9202 2202
rect 9202 2150 9232 2202
rect 9256 2150 9266 2202
rect 9266 2150 9312 2202
rect 9016 2148 9072 2150
rect 9096 2148 9152 2150
rect 9176 2148 9232 2150
rect 9256 2148 9312 2150
rect 11058 1808 11114 1864
rect 15016 2202 15072 2204
rect 15096 2202 15152 2204
rect 15176 2202 15232 2204
rect 15256 2202 15312 2204
rect 15016 2150 15062 2202
rect 15062 2150 15072 2202
rect 15096 2150 15126 2202
rect 15126 2150 15138 2202
rect 15138 2150 15152 2202
rect 15176 2150 15190 2202
rect 15190 2150 15202 2202
rect 15202 2150 15232 2202
rect 15256 2150 15266 2202
rect 15266 2150 15312 2202
rect 15016 2148 15072 2150
rect 15096 2148 15152 2150
rect 15176 2148 15232 2150
rect 15256 2148 15312 2150
rect 15750 40 15806 96
rect 18050 8200 18106 8256
rect 19154 9968 19210 10024
rect 18510 7112 18566 7168
rect 18050 3712 18106 3768
rect 19522 6976 19578 7032
rect 19614 6432 19670 6488
rect 20902 9832 20958 9888
rect 19956 8186 20012 8188
rect 20036 8186 20092 8188
rect 20116 8186 20172 8188
rect 20196 8186 20252 8188
rect 19956 8134 20002 8186
rect 20002 8134 20012 8186
rect 20036 8134 20066 8186
rect 20066 8134 20078 8186
rect 20078 8134 20092 8186
rect 20116 8134 20130 8186
rect 20130 8134 20142 8186
rect 20142 8134 20172 8186
rect 20196 8134 20206 8186
rect 20206 8134 20252 8186
rect 19956 8132 20012 8134
rect 20036 8132 20092 8134
rect 20116 8132 20172 8134
rect 20196 8132 20252 8134
rect 21016 8730 21072 8732
rect 21096 8730 21152 8732
rect 21176 8730 21232 8732
rect 21256 8730 21312 8732
rect 21016 8678 21062 8730
rect 21062 8678 21072 8730
rect 21096 8678 21126 8730
rect 21126 8678 21138 8730
rect 21138 8678 21152 8730
rect 21176 8678 21190 8730
rect 21190 8678 21202 8730
rect 21202 8678 21232 8730
rect 21256 8678 21266 8730
rect 21266 8678 21312 8730
rect 21016 8676 21072 8678
rect 21096 8676 21152 8678
rect 21176 8676 21232 8678
rect 21256 8676 21312 8678
rect 19956 7098 20012 7100
rect 20036 7098 20092 7100
rect 20116 7098 20172 7100
rect 20196 7098 20252 7100
rect 19956 7046 20002 7098
rect 20002 7046 20012 7098
rect 20036 7046 20066 7098
rect 20066 7046 20078 7098
rect 20078 7046 20092 7098
rect 20116 7046 20130 7098
rect 20130 7046 20142 7098
rect 20142 7046 20172 7098
rect 20196 7046 20206 7098
rect 20206 7046 20252 7098
rect 19956 7044 20012 7046
rect 20036 7044 20092 7046
rect 20116 7044 20172 7046
rect 20196 7044 20252 7046
rect 20718 7928 20774 7984
rect 20902 7928 20958 7984
rect 20626 7112 20682 7168
rect 20534 6976 20590 7032
rect 20166 6432 20222 6488
rect 20350 6296 20406 6352
rect 20350 6024 20406 6080
rect 19956 6010 20012 6012
rect 20036 6010 20092 6012
rect 20116 6010 20172 6012
rect 20196 6010 20252 6012
rect 19956 5958 20002 6010
rect 20002 5958 20012 6010
rect 20036 5958 20066 6010
rect 20066 5958 20078 6010
rect 20078 5958 20092 6010
rect 20116 5958 20130 6010
rect 20130 5958 20142 6010
rect 20142 5958 20172 6010
rect 20196 5958 20206 6010
rect 20206 5958 20252 6010
rect 19956 5956 20012 5958
rect 20036 5956 20092 5958
rect 20116 5956 20172 5958
rect 20196 5956 20252 5958
rect 19706 5344 19762 5400
rect 19706 3848 19762 3904
rect 19956 4922 20012 4924
rect 20036 4922 20092 4924
rect 20116 4922 20172 4924
rect 20196 4922 20252 4924
rect 19956 4870 20002 4922
rect 20002 4870 20012 4922
rect 20036 4870 20066 4922
rect 20066 4870 20078 4922
rect 20078 4870 20092 4922
rect 20116 4870 20130 4922
rect 20130 4870 20142 4922
rect 20142 4870 20172 4922
rect 20196 4870 20206 4922
rect 20206 4870 20252 4922
rect 19956 4868 20012 4870
rect 20036 4868 20092 4870
rect 20116 4868 20172 4870
rect 20196 4868 20252 4870
rect 20626 6704 20682 6760
rect 20350 3848 20406 3904
rect 19956 3834 20012 3836
rect 20036 3834 20092 3836
rect 20116 3834 20172 3836
rect 20196 3834 20252 3836
rect 19956 3782 20002 3834
rect 20002 3782 20012 3834
rect 20036 3782 20066 3834
rect 20066 3782 20078 3834
rect 20078 3782 20092 3834
rect 20116 3782 20130 3834
rect 20130 3782 20142 3834
rect 20142 3782 20172 3834
rect 20196 3782 20206 3834
rect 20206 3782 20252 3834
rect 19956 3780 20012 3782
rect 20036 3780 20092 3782
rect 20116 3780 20172 3782
rect 20196 3780 20252 3782
rect 20810 7656 20866 7712
rect 21016 7642 21072 7644
rect 21096 7642 21152 7644
rect 21176 7642 21232 7644
rect 21256 7642 21312 7644
rect 21016 7590 21062 7642
rect 21062 7590 21072 7642
rect 21096 7590 21126 7642
rect 21126 7590 21138 7642
rect 21138 7590 21152 7642
rect 21176 7590 21190 7642
rect 21190 7590 21202 7642
rect 21202 7590 21232 7642
rect 21256 7590 21266 7642
rect 21266 7590 21312 7642
rect 21016 7588 21072 7590
rect 21096 7588 21152 7590
rect 21176 7588 21232 7590
rect 21256 7588 21312 7590
rect 20902 7384 20958 7440
rect 21178 7248 21234 7304
rect 21016 6554 21072 6556
rect 21096 6554 21152 6556
rect 21176 6554 21232 6556
rect 21256 6554 21312 6556
rect 21016 6502 21062 6554
rect 21062 6502 21072 6554
rect 21096 6502 21126 6554
rect 21126 6502 21138 6554
rect 21138 6502 21152 6554
rect 21176 6502 21190 6554
rect 21190 6502 21202 6554
rect 21202 6502 21232 6554
rect 21256 6502 21266 6554
rect 21266 6502 21312 6554
rect 21016 6500 21072 6502
rect 21096 6500 21152 6502
rect 21176 6500 21232 6502
rect 21256 6500 21312 6502
rect 20350 3032 20406 3088
rect 21016 5466 21072 5468
rect 21096 5466 21152 5468
rect 21176 5466 21232 5468
rect 21256 5466 21312 5468
rect 21016 5414 21062 5466
rect 21062 5414 21072 5466
rect 21096 5414 21126 5466
rect 21126 5414 21138 5466
rect 21138 5414 21152 5466
rect 21176 5414 21190 5466
rect 21190 5414 21202 5466
rect 21202 5414 21232 5466
rect 21256 5414 21266 5466
rect 21266 5414 21312 5466
rect 21016 5412 21072 5414
rect 21096 5412 21152 5414
rect 21176 5412 21232 5414
rect 21256 5412 21312 5414
rect 21016 4378 21072 4380
rect 21096 4378 21152 4380
rect 21176 4378 21232 4380
rect 21256 4378 21312 4380
rect 21016 4326 21062 4378
rect 21062 4326 21072 4378
rect 21096 4326 21126 4378
rect 21126 4326 21138 4378
rect 21138 4326 21152 4378
rect 21176 4326 21190 4378
rect 21190 4326 21202 4378
rect 21202 4326 21232 4378
rect 21256 4326 21266 4378
rect 21266 4326 21312 4378
rect 21016 4324 21072 4326
rect 21096 4324 21152 4326
rect 21176 4324 21232 4326
rect 21256 4324 21312 4326
rect 22282 7520 22338 7576
rect 21730 7112 21786 7168
rect 21730 6568 21786 6624
rect 21730 5888 21786 5944
rect 21730 5480 21786 5536
rect 21730 4820 21786 4856
rect 21730 4800 21732 4820
rect 21732 4800 21784 4820
rect 21784 4800 21786 4820
rect 21546 4120 21602 4176
rect 22006 6840 22062 6896
rect 21016 3290 21072 3292
rect 21096 3290 21152 3292
rect 21176 3290 21232 3292
rect 21256 3290 21312 3292
rect 21016 3238 21062 3290
rect 21062 3238 21072 3290
rect 21096 3238 21126 3290
rect 21126 3238 21138 3290
rect 21138 3238 21152 3290
rect 21176 3238 21190 3290
rect 21190 3238 21202 3290
rect 21202 3238 21232 3290
rect 21256 3238 21266 3290
rect 21266 3238 21312 3290
rect 21016 3236 21072 3238
rect 21096 3236 21152 3238
rect 21176 3236 21232 3238
rect 21256 3236 21312 3238
rect 22282 4664 22338 4720
rect 22650 6432 22706 6488
rect 22374 3848 22430 3904
rect 23110 6568 23166 6624
rect 20350 2760 20406 2816
rect 19956 2746 20012 2748
rect 20036 2746 20092 2748
rect 20116 2746 20172 2748
rect 20196 2746 20252 2748
rect 19956 2694 20002 2746
rect 20002 2694 20012 2746
rect 20036 2694 20066 2746
rect 20066 2694 20078 2746
rect 20078 2694 20092 2746
rect 20116 2694 20130 2746
rect 20130 2694 20142 2746
rect 20142 2694 20172 2746
rect 20196 2694 20206 2746
rect 20206 2694 20252 2746
rect 19956 2692 20012 2694
rect 20036 2692 20092 2694
rect 20116 2692 20172 2694
rect 20196 2692 20252 2694
rect 21016 2202 21072 2204
rect 21096 2202 21152 2204
rect 21176 2202 21232 2204
rect 21256 2202 21312 2204
rect 21016 2150 21062 2202
rect 21062 2150 21072 2202
rect 21096 2150 21126 2202
rect 21126 2150 21138 2202
rect 21138 2150 21152 2202
rect 21176 2150 21190 2202
rect 21190 2150 21202 2202
rect 21202 2150 21232 2202
rect 21256 2150 21266 2202
rect 21266 2150 21312 2202
rect 21016 2148 21072 2150
rect 21096 2148 21152 2150
rect 21176 2148 21232 2150
rect 21256 2148 21312 2150
rect 23386 7384 23442 7440
rect 23662 6432 23718 6488
rect 24030 10240 24086 10296
rect 25134 10376 25190 10432
rect 24674 8200 24730 8256
rect 25318 6024 25374 6080
rect 25956 8186 26012 8188
rect 26036 8186 26092 8188
rect 26116 8186 26172 8188
rect 26196 8186 26252 8188
rect 25956 8134 26002 8186
rect 26002 8134 26012 8186
rect 26036 8134 26066 8186
rect 26066 8134 26078 8186
rect 26078 8134 26092 8186
rect 26116 8134 26130 8186
rect 26130 8134 26142 8186
rect 26142 8134 26172 8186
rect 26196 8134 26206 8186
rect 26206 8134 26252 8186
rect 25956 8132 26012 8134
rect 26036 8132 26092 8134
rect 26116 8132 26172 8134
rect 26196 8132 26252 8134
rect 25956 7098 26012 7100
rect 26036 7098 26092 7100
rect 26116 7098 26172 7100
rect 26196 7098 26252 7100
rect 25956 7046 26002 7098
rect 26002 7046 26012 7098
rect 26036 7046 26066 7098
rect 26066 7046 26078 7098
rect 26078 7046 26092 7098
rect 26116 7046 26130 7098
rect 26130 7046 26142 7098
rect 26142 7046 26172 7098
rect 26196 7046 26206 7098
rect 26206 7046 26252 7098
rect 25956 7044 26012 7046
rect 26036 7044 26092 7046
rect 26116 7044 26172 7046
rect 26196 7044 26252 7046
rect 25956 6010 26012 6012
rect 26036 6010 26092 6012
rect 26116 6010 26172 6012
rect 26196 6010 26252 6012
rect 25956 5958 26002 6010
rect 26002 5958 26012 6010
rect 26036 5958 26066 6010
rect 26066 5958 26078 6010
rect 26078 5958 26092 6010
rect 26116 5958 26130 6010
rect 26130 5958 26142 6010
rect 26142 5958 26172 6010
rect 26196 5958 26206 6010
rect 26206 5958 26252 6010
rect 25956 5956 26012 5958
rect 26036 5956 26092 5958
rect 26116 5956 26172 5958
rect 26196 5956 26252 5958
rect 26330 5480 26386 5536
rect 25502 4528 25558 4584
rect 27016 8730 27072 8732
rect 27096 8730 27152 8732
rect 27176 8730 27232 8732
rect 27256 8730 27312 8732
rect 27016 8678 27062 8730
rect 27062 8678 27072 8730
rect 27096 8678 27126 8730
rect 27126 8678 27138 8730
rect 27138 8678 27152 8730
rect 27176 8678 27190 8730
rect 27190 8678 27202 8730
rect 27202 8678 27232 8730
rect 27256 8678 27266 8730
rect 27266 8678 27312 8730
rect 27016 8676 27072 8678
rect 27096 8676 27152 8678
rect 27176 8676 27232 8678
rect 27256 8676 27312 8678
rect 25956 4922 26012 4924
rect 26036 4922 26092 4924
rect 26116 4922 26172 4924
rect 26196 4922 26252 4924
rect 25956 4870 26002 4922
rect 26002 4870 26012 4922
rect 26036 4870 26066 4922
rect 26066 4870 26078 4922
rect 26078 4870 26092 4922
rect 26116 4870 26130 4922
rect 26130 4870 26142 4922
rect 26142 4870 26172 4922
rect 26196 4870 26206 4922
rect 26206 4870 26252 4922
rect 25956 4868 26012 4870
rect 26036 4868 26092 4870
rect 26116 4868 26172 4870
rect 26196 4868 26252 4870
rect 25956 3834 26012 3836
rect 26036 3834 26092 3836
rect 26116 3834 26172 3836
rect 26196 3834 26252 3836
rect 25956 3782 26002 3834
rect 26002 3782 26012 3834
rect 26036 3782 26066 3834
rect 26066 3782 26078 3834
rect 26078 3782 26092 3834
rect 26116 3782 26130 3834
rect 26130 3782 26142 3834
rect 26142 3782 26172 3834
rect 26196 3782 26206 3834
rect 26206 3782 26252 3834
rect 25956 3780 26012 3782
rect 26036 3780 26092 3782
rect 26116 3780 26172 3782
rect 26196 3780 26252 3782
rect 26514 3712 26570 3768
rect 25778 3168 25834 3224
rect 26606 3440 26662 3496
rect 26514 3168 26570 3224
rect 25778 2760 25834 2816
rect 26606 2760 26662 2816
rect 25956 2746 26012 2748
rect 26036 2746 26092 2748
rect 26116 2746 26172 2748
rect 26196 2746 26252 2748
rect 25956 2694 26002 2746
rect 26002 2694 26012 2746
rect 26036 2694 26066 2746
rect 26066 2694 26078 2746
rect 26078 2694 26092 2746
rect 26116 2694 26130 2746
rect 26130 2694 26142 2746
rect 26142 2694 26172 2746
rect 26196 2694 26206 2746
rect 26206 2694 26252 2746
rect 25956 2692 26012 2694
rect 26036 2692 26092 2694
rect 26116 2692 26172 2694
rect 26196 2692 26252 2694
rect 27016 7642 27072 7644
rect 27096 7642 27152 7644
rect 27176 7642 27232 7644
rect 27256 7642 27312 7644
rect 27016 7590 27062 7642
rect 27062 7590 27072 7642
rect 27096 7590 27126 7642
rect 27126 7590 27138 7642
rect 27138 7590 27152 7642
rect 27176 7590 27190 7642
rect 27190 7590 27202 7642
rect 27202 7590 27232 7642
rect 27256 7590 27266 7642
rect 27266 7590 27312 7642
rect 27016 7588 27072 7590
rect 27096 7588 27152 7590
rect 27176 7588 27232 7590
rect 27256 7588 27312 7590
rect 27016 6554 27072 6556
rect 27096 6554 27152 6556
rect 27176 6554 27232 6556
rect 27256 6554 27312 6556
rect 27016 6502 27062 6554
rect 27062 6502 27072 6554
rect 27096 6502 27126 6554
rect 27126 6502 27138 6554
rect 27138 6502 27152 6554
rect 27176 6502 27190 6554
rect 27190 6502 27202 6554
rect 27202 6502 27232 6554
rect 27256 6502 27266 6554
rect 27266 6502 27312 6554
rect 27016 6500 27072 6502
rect 27096 6500 27152 6502
rect 27176 6500 27232 6502
rect 27256 6500 27312 6502
rect 27986 9152 28042 9208
rect 27710 6876 27712 6896
rect 27712 6876 27764 6896
rect 27764 6876 27766 6896
rect 27710 6840 27766 6876
rect 28262 9424 28318 9480
rect 28814 10104 28870 10160
rect 29366 9696 29422 9752
rect 27016 5466 27072 5468
rect 27096 5466 27152 5468
rect 27176 5466 27232 5468
rect 27256 5466 27312 5468
rect 27016 5414 27062 5466
rect 27062 5414 27072 5466
rect 27096 5414 27126 5466
rect 27126 5414 27138 5466
rect 27138 5414 27152 5466
rect 27176 5414 27190 5466
rect 27190 5414 27202 5466
rect 27202 5414 27232 5466
rect 27256 5414 27266 5466
rect 27266 5414 27312 5466
rect 27016 5412 27072 5414
rect 27096 5412 27152 5414
rect 27176 5412 27232 5414
rect 27256 5412 27312 5414
rect 27016 4378 27072 4380
rect 27096 4378 27152 4380
rect 27176 4378 27232 4380
rect 27256 4378 27312 4380
rect 27016 4326 27062 4378
rect 27062 4326 27072 4378
rect 27096 4326 27126 4378
rect 27126 4326 27138 4378
rect 27138 4326 27152 4378
rect 27176 4326 27190 4378
rect 27190 4326 27202 4378
rect 27202 4326 27232 4378
rect 27256 4326 27266 4378
rect 27266 4326 27312 4378
rect 27016 4324 27072 4326
rect 27096 4324 27152 4326
rect 27176 4324 27232 4326
rect 27256 4324 27312 4326
rect 27016 3290 27072 3292
rect 27096 3290 27152 3292
rect 27176 3290 27232 3292
rect 27256 3290 27312 3292
rect 27016 3238 27062 3290
rect 27062 3238 27072 3290
rect 27096 3238 27126 3290
rect 27126 3238 27138 3290
rect 27138 3238 27152 3290
rect 27176 3238 27190 3290
rect 27190 3238 27202 3290
rect 27202 3238 27232 3290
rect 27256 3238 27266 3290
rect 27266 3238 27312 3290
rect 27016 3236 27072 3238
rect 27096 3236 27152 3238
rect 27176 3236 27232 3238
rect 27256 3236 27312 3238
rect 27016 2202 27072 2204
rect 27096 2202 27152 2204
rect 27176 2202 27232 2204
rect 27256 2202 27312 2204
rect 27016 2150 27062 2202
rect 27062 2150 27072 2202
rect 27096 2150 27126 2202
rect 27126 2150 27138 2202
rect 27138 2150 27152 2202
rect 27176 2150 27190 2202
rect 27190 2150 27202 2202
rect 27202 2150 27232 2202
rect 27256 2150 27266 2202
rect 27266 2150 27312 2202
rect 27016 2148 27072 2150
rect 27096 2148 27152 2150
rect 27176 2148 27232 2150
rect 27256 2148 27312 2150
rect 29826 7928 29882 7984
rect 29918 7384 29974 7440
rect 29182 3712 29238 3768
rect 30378 6296 30434 6352
rect 31482 9288 31538 9344
rect 31758 8472 31814 8528
rect 31956 8186 32012 8188
rect 32036 8186 32092 8188
rect 32116 8186 32172 8188
rect 32196 8186 32252 8188
rect 31956 8134 32002 8186
rect 32002 8134 32012 8186
rect 32036 8134 32066 8186
rect 32066 8134 32078 8186
rect 32078 8134 32092 8186
rect 32116 8134 32130 8186
rect 32130 8134 32142 8186
rect 32142 8134 32172 8186
rect 32196 8134 32206 8186
rect 32206 8134 32252 8186
rect 31956 8132 32012 8134
rect 32036 8132 32092 8134
rect 32116 8132 32172 8134
rect 32196 8132 32252 8134
rect 32126 7792 32182 7848
rect 33016 8730 33072 8732
rect 33096 8730 33152 8732
rect 33176 8730 33232 8732
rect 33256 8730 33312 8732
rect 33016 8678 33062 8730
rect 33062 8678 33072 8730
rect 33096 8678 33126 8730
rect 33126 8678 33138 8730
rect 33138 8678 33152 8730
rect 33176 8678 33190 8730
rect 33190 8678 33202 8730
rect 33202 8678 33232 8730
rect 33256 8678 33266 8730
rect 33266 8678 33312 8730
rect 33016 8676 33072 8678
rect 33096 8676 33152 8678
rect 33176 8676 33232 8678
rect 33256 8676 33312 8678
rect 32402 7248 32458 7304
rect 31956 7098 32012 7100
rect 32036 7098 32092 7100
rect 32116 7098 32172 7100
rect 32196 7098 32252 7100
rect 31956 7046 32002 7098
rect 32002 7046 32012 7098
rect 32036 7046 32066 7098
rect 32066 7046 32078 7098
rect 32078 7046 32092 7098
rect 32116 7046 32130 7098
rect 32130 7046 32142 7098
rect 32142 7046 32172 7098
rect 32196 7046 32206 7098
rect 32206 7046 32252 7098
rect 31956 7044 32012 7046
rect 32036 7044 32092 7046
rect 32116 7044 32172 7046
rect 32196 7044 32252 7046
rect 31298 2488 31354 2544
rect 30286 1808 30342 1864
rect 31956 6010 32012 6012
rect 32036 6010 32092 6012
rect 32116 6010 32172 6012
rect 32196 6010 32252 6012
rect 31956 5958 32002 6010
rect 32002 5958 32012 6010
rect 32036 5958 32066 6010
rect 32066 5958 32078 6010
rect 32078 5958 32092 6010
rect 32116 5958 32130 6010
rect 32130 5958 32142 6010
rect 32142 5958 32172 6010
rect 32196 5958 32206 6010
rect 32206 5958 32252 6010
rect 31956 5956 32012 5958
rect 32036 5956 32092 5958
rect 32116 5956 32172 5958
rect 32196 5956 32252 5958
rect 31956 4922 32012 4924
rect 32036 4922 32092 4924
rect 32116 4922 32172 4924
rect 32196 4922 32252 4924
rect 31956 4870 32002 4922
rect 32002 4870 32012 4922
rect 32036 4870 32066 4922
rect 32066 4870 32078 4922
rect 32078 4870 32092 4922
rect 32116 4870 32130 4922
rect 32130 4870 32142 4922
rect 32142 4870 32172 4922
rect 32196 4870 32206 4922
rect 32206 4870 32252 4922
rect 31956 4868 32012 4870
rect 32036 4868 32092 4870
rect 32116 4868 32172 4870
rect 32196 4868 32252 4870
rect 32770 6160 32826 6216
rect 31956 3834 32012 3836
rect 32036 3834 32092 3836
rect 32116 3834 32172 3836
rect 32196 3834 32252 3836
rect 31956 3782 32002 3834
rect 32002 3782 32012 3834
rect 32036 3782 32066 3834
rect 32066 3782 32078 3834
rect 32078 3782 32092 3834
rect 32116 3782 32130 3834
rect 32130 3782 32142 3834
rect 32142 3782 32172 3834
rect 32196 3782 32206 3834
rect 32206 3782 32252 3834
rect 31956 3780 32012 3782
rect 32036 3780 32092 3782
rect 32116 3780 32172 3782
rect 32196 3780 32252 3782
rect 31956 2746 32012 2748
rect 32036 2746 32092 2748
rect 32116 2746 32172 2748
rect 32196 2746 32252 2748
rect 31956 2694 32002 2746
rect 32002 2694 32012 2746
rect 32036 2694 32066 2746
rect 32066 2694 32078 2746
rect 32078 2694 32092 2746
rect 32116 2694 32130 2746
rect 32130 2694 32142 2746
rect 32142 2694 32172 2746
rect 32196 2694 32206 2746
rect 32206 2694 32252 2746
rect 31956 2692 32012 2694
rect 32036 2692 32092 2694
rect 32116 2692 32172 2694
rect 32196 2692 32252 2694
rect 31666 40 31722 96
rect 33016 7642 33072 7644
rect 33096 7642 33152 7644
rect 33176 7642 33232 7644
rect 33256 7642 33312 7644
rect 33016 7590 33062 7642
rect 33062 7590 33072 7642
rect 33096 7590 33126 7642
rect 33126 7590 33138 7642
rect 33138 7590 33152 7642
rect 33176 7590 33190 7642
rect 33190 7590 33202 7642
rect 33202 7590 33232 7642
rect 33256 7590 33266 7642
rect 33266 7590 33312 7642
rect 33016 7588 33072 7590
rect 33096 7588 33152 7590
rect 33176 7588 33232 7590
rect 33256 7588 33312 7590
rect 33016 6554 33072 6556
rect 33096 6554 33152 6556
rect 33176 6554 33232 6556
rect 33256 6554 33312 6556
rect 33016 6502 33062 6554
rect 33062 6502 33072 6554
rect 33096 6502 33126 6554
rect 33126 6502 33138 6554
rect 33138 6502 33152 6554
rect 33176 6502 33190 6554
rect 33190 6502 33202 6554
rect 33202 6502 33232 6554
rect 33256 6502 33266 6554
rect 33266 6502 33312 6554
rect 33016 6500 33072 6502
rect 33096 6500 33152 6502
rect 33176 6500 33232 6502
rect 33256 6500 33312 6502
rect 33016 5466 33072 5468
rect 33096 5466 33152 5468
rect 33176 5466 33232 5468
rect 33256 5466 33312 5468
rect 33016 5414 33062 5466
rect 33062 5414 33072 5466
rect 33096 5414 33126 5466
rect 33126 5414 33138 5466
rect 33138 5414 33152 5466
rect 33176 5414 33190 5466
rect 33190 5414 33202 5466
rect 33202 5414 33232 5466
rect 33256 5414 33266 5466
rect 33266 5414 33312 5466
rect 33016 5412 33072 5414
rect 33096 5412 33152 5414
rect 33176 5412 33232 5414
rect 33256 5412 33312 5414
rect 33016 4378 33072 4380
rect 33096 4378 33152 4380
rect 33176 4378 33232 4380
rect 33256 4378 33312 4380
rect 33016 4326 33062 4378
rect 33062 4326 33072 4378
rect 33096 4326 33126 4378
rect 33126 4326 33138 4378
rect 33138 4326 33152 4378
rect 33176 4326 33190 4378
rect 33190 4326 33202 4378
rect 33202 4326 33232 4378
rect 33256 4326 33266 4378
rect 33266 4326 33312 4378
rect 33016 4324 33072 4326
rect 33096 4324 33152 4326
rect 33176 4324 33232 4326
rect 33256 4324 33312 4326
rect 34242 7404 34298 7440
rect 34242 7384 34244 7404
rect 34244 7384 34296 7404
rect 34296 7384 34298 7404
rect 33016 3290 33072 3292
rect 33096 3290 33152 3292
rect 33176 3290 33232 3292
rect 33256 3290 33312 3292
rect 33016 3238 33062 3290
rect 33062 3238 33072 3290
rect 33096 3238 33126 3290
rect 33126 3238 33138 3290
rect 33138 3238 33152 3290
rect 33176 3238 33190 3290
rect 33190 3238 33202 3290
rect 33202 3238 33232 3290
rect 33256 3238 33266 3290
rect 33266 3238 33312 3290
rect 33016 3236 33072 3238
rect 33096 3236 33152 3238
rect 33176 3236 33232 3238
rect 33256 3236 33312 3238
rect 33016 2202 33072 2204
rect 33096 2202 33152 2204
rect 33176 2202 33232 2204
rect 33256 2202 33312 2204
rect 33016 2150 33062 2202
rect 33062 2150 33072 2202
rect 33096 2150 33126 2202
rect 33126 2150 33138 2202
rect 33138 2150 33152 2202
rect 33176 2150 33190 2202
rect 33190 2150 33202 2202
rect 33202 2150 33232 2202
rect 33256 2150 33266 2202
rect 33266 2150 33312 2202
rect 33016 2148 33072 2150
rect 33096 2148 33152 2150
rect 33176 2148 33232 2150
rect 33256 2148 33312 2150
rect 34518 1944 34574 2000
rect 35898 6704 35954 6760
rect 35990 5616 36046 5672
rect 37094 8880 37150 8936
rect 37370 9016 37426 9072
rect 38290 9832 38346 9888
rect 37956 8186 38012 8188
rect 38036 8186 38092 8188
rect 38116 8186 38172 8188
rect 38196 8186 38252 8188
rect 37956 8134 38002 8186
rect 38002 8134 38012 8186
rect 38036 8134 38066 8186
rect 38066 8134 38078 8186
rect 38078 8134 38092 8186
rect 38116 8134 38130 8186
rect 38130 8134 38142 8186
rect 38142 8134 38172 8186
rect 38196 8134 38206 8186
rect 38206 8134 38252 8186
rect 37956 8132 38012 8134
rect 38036 8132 38092 8134
rect 38116 8132 38172 8134
rect 38196 8132 38252 8134
rect 37554 2524 37556 2544
rect 37556 2524 37608 2544
rect 37608 2524 37610 2544
rect 37554 2488 37610 2524
rect 37462 1672 37518 1728
rect 39578 9560 39634 9616
rect 38750 9288 38806 9344
rect 38658 8472 38714 8528
rect 37956 7098 38012 7100
rect 38036 7098 38092 7100
rect 38116 7098 38172 7100
rect 38196 7098 38252 7100
rect 37956 7046 38002 7098
rect 38002 7046 38012 7098
rect 38036 7046 38066 7098
rect 38066 7046 38078 7098
rect 38078 7046 38092 7098
rect 38116 7046 38130 7098
rect 38130 7046 38142 7098
rect 38142 7046 38172 7098
rect 38196 7046 38206 7098
rect 38206 7046 38252 7098
rect 37956 7044 38012 7046
rect 38036 7044 38092 7046
rect 38116 7044 38172 7046
rect 38196 7044 38252 7046
rect 37956 6010 38012 6012
rect 38036 6010 38092 6012
rect 38116 6010 38172 6012
rect 38196 6010 38252 6012
rect 37956 5958 38002 6010
rect 38002 5958 38012 6010
rect 38036 5958 38066 6010
rect 38066 5958 38078 6010
rect 38078 5958 38092 6010
rect 38116 5958 38130 6010
rect 38130 5958 38142 6010
rect 38142 5958 38172 6010
rect 38196 5958 38206 6010
rect 38206 5958 38252 6010
rect 37956 5956 38012 5958
rect 38036 5956 38092 5958
rect 38116 5956 38172 5958
rect 38196 5956 38252 5958
rect 37956 4922 38012 4924
rect 38036 4922 38092 4924
rect 38116 4922 38172 4924
rect 38196 4922 38252 4924
rect 37956 4870 38002 4922
rect 38002 4870 38012 4922
rect 38036 4870 38066 4922
rect 38066 4870 38078 4922
rect 38078 4870 38092 4922
rect 38116 4870 38130 4922
rect 38130 4870 38142 4922
rect 38142 4870 38172 4922
rect 38196 4870 38206 4922
rect 38206 4870 38252 4922
rect 37956 4868 38012 4870
rect 38036 4868 38092 4870
rect 38116 4868 38172 4870
rect 38196 4868 38252 4870
rect 39486 8744 39542 8800
rect 39016 8730 39072 8732
rect 39096 8730 39152 8732
rect 39176 8730 39232 8732
rect 39256 8730 39312 8732
rect 39016 8678 39062 8730
rect 39062 8678 39072 8730
rect 39096 8678 39126 8730
rect 39126 8678 39138 8730
rect 39138 8678 39152 8730
rect 39176 8678 39190 8730
rect 39190 8678 39202 8730
rect 39202 8678 39232 8730
rect 39256 8678 39266 8730
rect 39266 8678 39312 8730
rect 39016 8676 39072 8678
rect 39096 8676 39152 8678
rect 39176 8676 39232 8678
rect 39256 8676 39312 8678
rect 39026 8356 39082 8392
rect 39026 8336 39028 8356
rect 39028 8336 39080 8356
rect 39080 8336 39082 8356
rect 39394 7928 39450 7984
rect 39394 7692 39396 7712
rect 39396 7692 39448 7712
rect 39448 7692 39450 7712
rect 39394 7656 39450 7692
rect 39016 7642 39072 7644
rect 39096 7642 39152 7644
rect 39176 7642 39232 7644
rect 39256 7642 39312 7644
rect 39016 7590 39062 7642
rect 39062 7590 39072 7642
rect 39096 7590 39126 7642
rect 39126 7590 39138 7642
rect 39138 7590 39152 7642
rect 39176 7590 39190 7642
rect 39190 7590 39202 7642
rect 39202 7590 39232 7642
rect 39256 7590 39266 7642
rect 39266 7590 39312 7642
rect 39016 7588 39072 7590
rect 39096 7588 39152 7590
rect 39176 7588 39232 7590
rect 39256 7588 39312 7590
rect 38934 7384 38990 7440
rect 38658 6296 38714 6352
rect 39394 7112 39450 7168
rect 39486 6840 39542 6896
rect 40038 9016 40094 9072
rect 39854 8200 39910 8256
rect 39578 6568 39634 6624
rect 39016 6554 39072 6556
rect 39096 6554 39152 6556
rect 39176 6554 39232 6556
rect 39256 6554 39312 6556
rect 39016 6502 39062 6554
rect 39062 6502 39072 6554
rect 39096 6502 39126 6554
rect 39126 6502 39138 6554
rect 39138 6502 39152 6554
rect 39176 6502 39190 6554
rect 39190 6502 39202 6554
rect 39202 6502 39232 6554
rect 39256 6502 39266 6554
rect 39266 6502 39312 6554
rect 39016 6500 39072 6502
rect 39096 6500 39152 6502
rect 39176 6500 39232 6502
rect 39256 6500 39312 6502
rect 39026 6060 39028 6080
rect 39028 6060 39080 6080
rect 39080 6060 39082 6080
rect 39026 6024 39082 6060
rect 39210 5752 39266 5808
rect 39486 5752 39542 5808
rect 39394 5480 39450 5536
rect 39016 5466 39072 5468
rect 39096 5466 39152 5468
rect 39176 5466 39232 5468
rect 39256 5466 39312 5468
rect 39016 5414 39062 5466
rect 39062 5414 39072 5466
rect 39096 5414 39126 5466
rect 39126 5414 39138 5466
rect 39138 5414 39152 5466
rect 39176 5414 39190 5466
rect 39190 5414 39202 5466
rect 39202 5414 39232 5466
rect 39256 5414 39266 5466
rect 39266 5414 39312 5466
rect 39016 5412 39072 5414
rect 39096 5412 39152 5414
rect 39176 5412 39232 5414
rect 39256 5412 39312 5414
rect 39210 5228 39266 5264
rect 39210 5208 39212 5228
rect 39212 5208 39264 5228
rect 39264 5208 39266 5228
rect 39394 5208 39450 5264
rect 39026 4972 39028 4992
rect 39028 4972 39080 4992
rect 39080 4972 39082 4992
rect 39026 4936 39082 4972
rect 39486 4664 39542 4720
rect 38842 3984 38898 4040
rect 37956 3834 38012 3836
rect 38036 3834 38092 3836
rect 38116 3834 38172 3836
rect 38196 3834 38252 3836
rect 37956 3782 38002 3834
rect 38002 3782 38012 3834
rect 38036 3782 38066 3834
rect 38066 3782 38078 3834
rect 38078 3782 38092 3834
rect 38116 3782 38130 3834
rect 38130 3782 38142 3834
rect 38142 3782 38172 3834
rect 38196 3782 38206 3834
rect 38206 3782 38252 3834
rect 37956 3780 38012 3782
rect 38036 3780 38092 3782
rect 38116 3780 38172 3782
rect 38196 3780 38252 3782
rect 37956 2746 38012 2748
rect 38036 2746 38092 2748
rect 38116 2746 38172 2748
rect 38196 2746 38252 2748
rect 37956 2694 38002 2746
rect 38002 2694 38012 2746
rect 38036 2694 38066 2746
rect 38066 2694 38078 2746
rect 38078 2694 38092 2746
rect 38116 2694 38130 2746
rect 38130 2694 38142 2746
rect 38142 2694 38172 2746
rect 38196 2694 38206 2746
rect 38206 2694 38252 2746
rect 37956 2692 38012 2694
rect 38036 2692 38092 2694
rect 38116 2692 38172 2694
rect 38196 2692 38252 2694
rect 38842 3440 38898 3496
rect 38474 2896 38530 2952
rect 38842 2796 38844 2816
rect 38844 2796 38896 2816
rect 38896 2796 38898 2816
rect 38842 2760 38898 2796
rect 39394 4392 39450 4448
rect 39016 4378 39072 4380
rect 39096 4378 39152 4380
rect 39176 4378 39232 4380
rect 39256 4378 39312 4380
rect 39016 4326 39062 4378
rect 39062 4326 39072 4378
rect 39096 4326 39126 4378
rect 39126 4326 39138 4378
rect 39138 4326 39152 4378
rect 39176 4326 39190 4378
rect 39190 4326 39202 4378
rect 39202 4326 39232 4378
rect 39256 4326 39266 4378
rect 39266 4326 39312 4378
rect 39016 4324 39072 4326
rect 39096 4324 39152 4326
rect 39176 4324 39232 4326
rect 39256 4324 39312 4326
rect 39394 4120 39450 4176
rect 39026 3884 39028 3904
rect 39028 3884 39080 3904
rect 39080 3884 39082 3904
rect 39026 3848 39082 3884
rect 39210 3576 39266 3632
rect 39486 3576 39542 3632
rect 39394 3304 39450 3360
rect 39016 3290 39072 3292
rect 39096 3290 39152 3292
rect 39176 3290 39232 3292
rect 39256 3290 39312 3292
rect 39016 3238 39062 3290
rect 39062 3238 39072 3290
rect 39096 3238 39126 3290
rect 39126 3238 39138 3290
rect 39138 3238 39152 3290
rect 39176 3238 39190 3290
rect 39190 3238 39202 3290
rect 39202 3238 39232 3290
rect 39256 3238 39266 3290
rect 39266 3238 39312 3290
rect 39016 3236 39072 3238
rect 39096 3236 39152 3238
rect 39176 3236 39232 3238
rect 39256 3236 39312 3238
rect 39210 3052 39266 3088
rect 39210 3032 39212 3052
rect 39212 3032 39264 3052
rect 39264 3032 39266 3052
rect 39394 3032 39450 3088
rect 37830 1944 37886 2000
rect 38290 1672 38346 1728
rect 39016 2202 39072 2204
rect 39096 2202 39152 2204
rect 39176 2202 39232 2204
rect 39256 2202 39312 2204
rect 39016 2150 39062 2202
rect 39062 2150 39072 2202
rect 39096 2150 39126 2202
rect 39126 2150 39138 2202
rect 39138 2150 39152 2202
rect 39176 2150 39190 2202
rect 39190 2150 39202 2202
rect 39202 2150 39232 2202
rect 39256 2150 39266 2202
rect 39266 2150 39312 2202
rect 39016 2148 39072 2150
rect 39096 2148 39152 2150
rect 39176 2148 39232 2150
rect 39256 2148 39312 2150
rect 37738 1400 37794 1456
rect 38658 1400 38714 1456
rect 39946 2216 40002 2272
<< metal3 >>
rect 5625 10434 5691 10437
rect 25129 10434 25195 10437
rect 5625 10432 25195 10434
rect 5625 10376 5630 10432
rect 5686 10376 25134 10432
rect 25190 10376 25195 10432
rect 5625 10374 25195 10376
rect 5625 10371 5691 10374
rect 25129 10371 25195 10374
rect 6637 10298 6703 10301
rect 24025 10298 24091 10301
rect 6637 10296 24091 10298
rect 6637 10240 6642 10296
rect 6698 10240 24030 10296
rect 24086 10240 24091 10296
rect 6637 10238 24091 10240
rect 6637 10235 6703 10238
rect 24025 10235 24091 10238
rect 9673 10162 9739 10165
rect 28809 10162 28875 10165
rect 9673 10160 28875 10162
rect 9673 10104 9678 10160
rect 9734 10104 28814 10160
rect 28870 10104 28875 10160
rect 9673 10102 28875 10104
rect 9673 10099 9739 10102
rect 28809 10099 28875 10102
rect 6729 10026 6795 10029
rect 19149 10026 19215 10029
rect 6729 10024 19215 10026
rect 6729 9968 6734 10024
rect 6790 9968 19154 10024
rect 19210 9968 19215 10024
rect 6729 9966 19215 9968
rect 6729 9963 6795 9966
rect 19149 9963 19215 9966
rect 0 9890 120 9920
rect 1117 9890 1183 9893
rect 0 9888 1183 9890
rect 0 9832 1122 9888
rect 1178 9832 1183 9888
rect 0 9830 1183 9832
rect 0 9800 120 9830
rect 1117 9827 1183 9830
rect 14733 9890 14799 9893
rect 20897 9890 20963 9893
rect 14733 9888 20963 9890
rect 14733 9832 14738 9888
rect 14794 9832 20902 9888
rect 20958 9832 20963 9888
rect 14733 9830 20963 9832
rect 14733 9827 14799 9830
rect 20897 9827 20963 9830
rect 38285 9890 38351 9893
rect 40880 9890 41000 9920
rect 38285 9888 41000 9890
rect 38285 9832 38290 9888
rect 38346 9832 41000 9888
rect 38285 9830 41000 9832
rect 38285 9827 38351 9830
rect 40880 9800 41000 9830
rect 8661 9754 8727 9757
rect 29361 9754 29427 9757
rect 8661 9752 29427 9754
rect 8661 9696 8666 9752
rect 8722 9696 29366 9752
rect 29422 9696 29427 9752
rect 8661 9694 29427 9696
rect 8661 9691 8727 9694
rect 29361 9691 29427 9694
rect 0 9618 120 9648
rect 1025 9618 1091 9621
rect 0 9616 1091 9618
rect 0 9560 1030 9616
rect 1086 9560 1091 9616
rect 0 9558 1091 9560
rect 0 9528 120 9558
rect 1025 9555 1091 9558
rect 39573 9618 39639 9621
rect 40880 9618 41000 9648
rect 39573 9616 41000 9618
rect 39573 9560 39578 9616
rect 39634 9560 41000 9616
rect 39573 9558 41000 9560
rect 39573 9555 39639 9558
rect 40880 9528 41000 9558
rect 10225 9482 10291 9485
rect 28257 9482 28323 9485
rect 10225 9480 28323 9482
rect 10225 9424 10230 9480
rect 10286 9424 28262 9480
rect 28318 9424 28323 9480
rect 10225 9422 28323 9424
rect 10225 9419 10291 9422
rect 28257 9419 28323 9422
rect 0 9346 120 9376
rect 841 9346 907 9349
rect 0 9344 907 9346
rect 0 9288 846 9344
rect 902 9288 907 9344
rect 0 9286 907 9288
rect 0 9256 120 9286
rect 841 9283 907 9286
rect 13353 9346 13419 9349
rect 31477 9346 31543 9349
rect 13353 9344 31543 9346
rect 13353 9288 13358 9344
rect 13414 9288 31482 9344
rect 31538 9288 31543 9344
rect 13353 9286 31543 9288
rect 13353 9283 13419 9286
rect 31477 9283 31543 9286
rect 38745 9346 38811 9349
rect 40880 9346 41000 9376
rect 38745 9344 41000 9346
rect 38745 9288 38750 9344
rect 38806 9288 41000 9344
rect 38745 9286 41000 9288
rect 38745 9283 38811 9286
rect 40880 9256 41000 9286
rect 3601 9210 3667 9213
rect 27981 9210 28047 9213
rect 3601 9208 28047 9210
rect 3601 9152 3606 9208
rect 3662 9152 27986 9208
rect 28042 9152 28047 9208
rect 3601 9150 28047 9152
rect 3601 9147 3667 9150
rect 27981 9147 28047 9150
rect 0 9074 120 9104
rect 1209 9074 1275 9077
rect 0 9072 1275 9074
rect 0 9016 1214 9072
rect 1270 9016 1275 9072
rect 0 9014 1275 9016
rect 0 8984 120 9014
rect 1209 9011 1275 9014
rect 16389 9074 16455 9077
rect 37365 9074 37431 9077
rect 16389 9072 37431 9074
rect 16389 9016 16394 9072
rect 16450 9016 37370 9072
rect 37426 9016 37431 9072
rect 16389 9014 37431 9016
rect 16389 9011 16455 9014
rect 37365 9011 37431 9014
rect 40033 9074 40099 9077
rect 40880 9074 41000 9104
rect 40033 9072 41000 9074
rect 40033 9016 40038 9072
rect 40094 9016 41000 9072
rect 40033 9014 41000 9016
rect 40033 9011 40099 9014
rect 40880 8984 41000 9014
rect 37089 8938 37155 8941
rect 2730 8936 37155 8938
rect 2730 8880 37094 8936
rect 37150 8880 37155 8936
rect 2730 8878 37155 8880
rect 0 8802 120 8832
rect 933 8802 999 8805
rect 0 8800 999 8802
rect 0 8744 938 8800
rect 994 8744 999 8800
rect 0 8742 999 8744
rect 0 8712 120 8742
rect 933 8739 999 8742
rect 0 8530 120 8560
rect 1301 8530 1367 8533
rect 0 8528 1367 8530
rect 0 8472 1306 8528
rect 1362 8472 1367 8528
rect 0 8470 1367 8472
rect 0 8440 120 8470
rect 1301 8467 1367 8470
rect 1117 8394 1183 8397
rect 2730 8394 2790 8878
rect 37089 8875 37155 8878
rect 39481 8802 39547 8805
rect 40880 8802 41000 8832
rect 39481 8800 41000 8802
rect 39481 8744 39486 8800
rect 39542 8744 41000 8800
rect 39481 8742 41000 8744
rect 39481 8739 39547 8742
rect 3006 8736 3322 8737
rect 3006 8672 3012 8736
rect 3076 8672 3092 8736
rect 3156 8672 3172 8736
rect 3236 8672 3252 8736
rect 3316 8672 3322 8736
rect 3006 8671 3322 8672
rect 9006 8736 9322 8737
rect 9006 8672 9012 8736
rect 9076 8672 9092 8736
rect 9156 8672 9172 8736
rect 9236 8672 9252 8736
rect 9316 8672 9322 8736
rect 9006 8671 9322 8672
rect 15006 8736 15322 8737
rect 15006 8672 15012 8736
rect 15076 8672 15092 8736
rect 15156 8672 15172 8736
rect 15236 8672 15252 8736
rect 15316 8672 15322 8736
rect 15006 8671 15322 8672
rect 21006 8736 21322 8737
rect 21006 8672 21012 8736
rect 21076 8672 21092 8736
rect 21156 8672 21172 8736
rect 21236 8672 21252 8736
rect 21316 8672 21322 8736
rect 21006 8671 21322 8672
rect 27006 8736 27322 8737
rect 27006 8672 27012 8736
rect 27076 8672 27092 8736
rect 27156 8672 27172 8736
rect 27236 8672 27252 8736
rect 27316 8672 27322 8736
rect 27006 8671 27322 8672
rect 33006 8736 33322 8737
rect 33006 8672 33012 8736
rect 33076 8672 33092 8736
rect 33156 8672 33172 8736
rect 33236 8672 33252 8736
rect 33316 8672 33322 8736
rect 33006 8671 33322 8672
rect 39006 8736 39322 8737
rect 39006 8672 39012 8736
rect 39076 8672 39092 8736
rect 39156 8672 39172 8736
rect 39236 8672 39252 8736
rect 39316 8672 39322 8736
rect 40880 8712 41000 8742
rect 39006 8671 39322 8672
rect 12985 8530 13051 8533
rect 31753 8530 31819 8533
rect 12985 8528 31819 8530
rect 12985 8472 12990 8528
rect 13046 8472 31758 8528
rect 31814 8472 31819 8528
rect 12985 8470 31819 8472
rect 12985 8467 13051 8470
rect 31753 8467 31819 8470
rect 38653 8530 38719 8533
rect 40880 8530 41000 8560
rect 38653 8528 41000 8530
rect 38653 8472 38658 8528
rect 38714 8472 41000 8528
rect 38653 8470 41000 8472
rect 38653 8467 38719 8470
rect 40880 8440 41000 8470
rect 1117 8392 2790 8394
rect 1117 8336 1122 8392
rect 1178 8336 2790 8392
rect 1117 8334 2790 8336
rect 7649 8394 7715 8397
rect 7649 8392 22110 8394
rect 7649 8336 7654 8392
rect 7710 8336 22110 8392
rect 7649 8334 22110 8336
rect 1117 8331 1183 8334
rect 7649 8331 7715 8334
rect 0 8258 120 8288
rect 1025 8258 1091 8261
rect 0 8256 1091 8258
rect 0 8200 1030 8256
rect 1086 8200 1091 8256
rect 0 8198 1091 8200
rect 0 8168 120 8198
rect 1025 8195 1091 8198
rect 14917 8258 14983 8261
rect 18045 8258 18111 8261
rect 14917 8256 18111 8258
rect 14917 8200 14922 8256
rect 14978 8200 18050 8256
rect 18106 8200 18111 8256
rect 14917 8198 18111 8200
rect 22050 8258 22110 8334
rect 27654 8332 27660 8396
rect 27724 8394 27730 8396
rect 39021 8394 39087 8397
rect 27724 8392 39087 8394
rect 27724 8336 39026 8392
rect 39082 8336 39087 8392
rect 27724 8334 39087 8336
rect 27724 8332 27730 8334
rect 39021 8331 39087 8334
rect 24669 8258 24735 8261
rect 22050 8256 24735 8258
rect 22050 8200 24674 8256
rect 24730 8200 24735 8256
rect 22050 8198 24735 8200
rect 14917 8195 14983 8198
rect 18045 8195 18111 8198
rect 24669 8195 24735 8198
rect 39849 8258 39915 8261
rect 40880 8258 41000 8288
rect 39849 8256 41000 8258
rect 39849 8200 39854 8256
rect 39910 8200 41000 8256
rect 39849 8198 41000 8200
rect 39849 8195 39915 8198
rect 1946 8192 2262 8193
rect 1946 8128 1952 8192
rect 2016 8128 2032 8192
rect 2096 8128 2112 8192
rect 2176 8128 2192 8192
rect 2256 8128 2262 8192
rect 1946 8127 2262 8128
rect 7946 8192 8262 8193
rect 7946 8128 7952 8192
rect 8016 8128 8032 8192
rect 8096 8128 8112 8192
rect 8176 8128 8192 8192
rect 8256 8128 8262 8192
rect 7946 8127 8262 8128
rect 13946 8192 14262 8193
rect 13946 8128 13952 8192
rect 14016 8128 14032 8192
rect 14096 8128 14112 8192
rect 14176 8128 14192 8192
rect 14256 8128 14262 8192
rect 13946 8127 14262 8128
rect 19946 8192 20262 8193
rect 19946 8128 19952 8192
rect 20016 8128 20032 8192
rect 20096 8128 20112 8192
rect 20176 8128 20192 8192
rect 20256 8128 20262 8192
rect 19946 8127 20262 8128
rect 25946 8192 26262 8193
rect 25946 8128 25952 8192
rect 26016 8128 26032 8192
rect 26096 8128 26112 8192
rect 26176 8128 26192 8192
rect 26256 8128 26262 8192
rect 25946 8127 26262 8128
rect 31946 8192 32262 8193
rect 31946 8128 31952 8192
rect 32016 8128 32032 8192
rect 32096 8128 32112 8192
rect 32176 8128 32192 8192
rect 32256 8128 32262 8192
rect 31946 8127 32262 8128
rect 37946 8192 38262 8193
rect 37946 8128 37952 8192
rect 38016 8128 38032 8192
rect 38096 8128 38112 8192
rect 38176 8128 38192 8192
rect 38256 8128 38262 8192
rect 40880 8168 41000 8198
rect 37946 8127 38262 8128
rect 0 7986 120 8016
rect 565 7986 631 7989
rect 0 7984 631 7986
rect 0 7928 570 7984
rect 626 7928 631 7984
rect 0 7926 631 7928
rect 0 7896 120 7926
rect 565 7923 631 7926
rect 1301 7986 1367 7989
rect 20713 7986 20779 7989
rect 1301 7984 20779 7986
rect 1301 7928 1306 7984
rect 1362 7928 20718 7984
rect 20774 7928 20779 7984
rect 1301 7926 20779 7928
rect 1301 7923 1367 7926
rect 20713 7923 20779 7926
rect 20897 7986 20963 7989
rect 29821 7986 29887 7989
rect 20897 7984 29887 7986
rect 20897 7928 20902 7984
rect 20958 7928 29826 7984
rect 29882 7928 29887 7984
rect 20897 7926 29887 7928
rect 20897 7923 20963 7926
rect 29821 7923 29887 7926
rect 39389 7986 39455 7989
rect 40880 7986 41000 8016
rect 39389 7984 41000 7986
rect 39389 7928 39394 7984
rect 39450 7928 41000 7984
rect 39389 7926 41000 7928
rect 39389 7923 39455 7926
rect 40880 7896 41000 7926
rect 9213 7850 9279 7853
rect 14641 7850 14707 7853
rect 32121 7850 32187 7853
rect 9213 7848 14474 7850
rect 9213 7792 9218 7848
rect 9274 7792 14474 7848
rect 9213 7790 14474 7792
rect 9213 7787 9279 7790
rect 0 7714 120 7744
rect 749 7714 815 7717
rect 0 7712 815 7714
rect 0 7656 754 7712
rect 810 7656 815 7712
rect 0 7654 815 7656
rect 0 7624 120 7654
rect 749 7651 815 7654
rect 3006 7648 3322 7649
rect 3006 7584 3012 7648
rect 3076 7584 3092 7648
rect 3156 7584 3172 7648
rect 3236 7584 3252 7648
rect 3316 7584 3322 7648
rect 3006 7583 3322 7584
rect 9006 7648 9322 7649
rect 9006 7584 9012 7648
rect 9076 7584 9092 7648
rect 9156 7584 9172 7648
rect 9236 7584 9252 7648
rect 9316 7584 9322 7648
rect 9006 7583 9322 7584
rect 13445 7578 13511 7581
rect 14181 7578 14247 7581
rect 13445 7576 14247 7578
rect 13445 7520 13450 7576
rect 13506 7520 14186 7576
rect 14242 7520 14247 7576
rect 13445 7518 14247 7520
rect 13445 7515 13511 7518
rect 14181 7515 14247 7518
rect 0 7442 120 7472
rect 565 7442 631 7445
rect 0 7440 631 7442
rect 0 7384 570 7440
rect 626 7384 631 7440
rect 0 7382 631 7384
rect 0 7352 120 7382
rect 565 7379 631 7382
rect 10777 7442 10843 7445
rect 14273 7442 14339 7445
rect 10777 7440 14339 7442
rect 10777 7384 10782 7440
rect 10838 7384 14278 7440
rect 14334 7384 14339 7440
rect 10777 7382 14339 7384
rect 14414 7442 14474 7790
rect 14641 7848 32187 7850
rect 14641 7792 14646 7848
rect 14702 7792 32126 7848
rect 32182 7792 32187 7848
rect 14641 7790 32187 7792
rect 14641 7787 14707 7790
rect 32121 7787 32187 7790
rect 15469 7714 15535 7717
rect 20805 7714 20871 7717
rect 15469 7712 20871 7714
rect 15469 7656 15474 7712
rect 15530 7656 20810 7712
rect 20866 7656 20871 7712
rect 15469 7654 20871 7656
rect 15469 7651 15535 7654
rect 20805 7651 20871 7654
rect 39389 7714 39455 7717
rect 40880 7714 41000 7744
rect 39389 7712 41000 7714
rect 39389 7656 39394 7712
rect 39450 7656 41000 7712
rect 39389 7654 41000 7656
rect 39389 7651 39455 7654
rect 15006 7648 15322 7649
rect 15006 7584 15012 7648
rect 15076 7584 15092 7648
rect 15156 7584 15172 7648
rect 15236 7584 15252 7648
rect 15316 7584 15322 7648
rect 15006 7583 15322 7584
rect 21006 7648 21322 7649
rect 21006 7584 21012 7648
rect 21076 7584 21092 7648
rect 21156 7584 21172 7648
rect 21236 7584 21252 7648
rect 21316 7584 21322 7648
rect 21006 7583 21322 7584
rect 27006 7648 27322 7649
rect 27006 7584 27012 7648
rect 27076 7584 27092 7648
rect 27156 7584 27172 7648
rect 27236 7584 27252 7648
rect 27316 7584 27322 7648
rect 27006 7583 27322 7584
rect 33006 7648 33322 7649
rect 33006 7584 33012 7648
rect 33076 7584 33092 7648
rect 33156 7584 33172 7648
rect 33236 7584 33252 7648
rect 33316 7584 33322 7648
rect 33006 7583 33322 7584
rect 39006 7648 39322 7649
rect 39006 7584 39012 7648
rect 39076 7584 39092 7648
rect 39156 7584 39172 7648
rect 39236 7584 39252 7648
rect 39316 7584 39322 7648
rect 40880 7624 41000 7654
rect 39006 7583 39322 7584
rect 15469 7578 15535 7581
rect 20846 7578 20852 7580
rect 15469 7576 20852 7578
rect 15469 7520 15474 7576
rect 15530 7520 20852 7576
rect 15469 7518 20852 7520
rect 15469 7515 15535 7518
rect 20846 7516 20852 7518
rect 20916 7516 20922 7580
rect 22134 7516 22140 7580
rect 22204 7578 22210 7580
rect 22277 7578 22343 7581
rect 22204 7576 22343 7578
rect 22204 7520 22282 7576
rect 22338 7520 22343 7576
rect 22204 7518 22343 7520
rect 22204 7516 22210 7518
rect 22277 7515 22343 7518
rect 20897 7442 20963 7445
rect 23381 7442 23447 7445
rect 14414 7440 20963 7442
rect 14414 7384 20902 7440
rect 20958 7384 20963 7440
rect 14414 7382 20963 7384
rect 10777 7379 10843 7382
rect 14273 7379 14339 7382
rect 20897 7379 20963 7382
rect 21038 7440 23447 7442
rect 21038 7384 23386 7440
rect 23442 7384 23447 7440
rect 21038 7382 23447 7384
rect 8201 7306 8267 7309
rect 13445 7306 13511 7309
rect 21038 7306 21098 7382
rect 23381 7379 23447 7382
rect 29913 7442 29979 7445
rect 34237 7442 34303 7445
rect 29913 7440 34303 7442
rect 29913 7384 29918 7440
rect 29974 7384 34242 7440
rect 34298 7384 34303 7440
rect 29913 7382 34303 7384
rect 29913 7379 29979 7382
rect 34237 7379 34303 7382
rect 38929 7442 38995 7445
rect 40880 7442 41000 7472
rect 38929 7440 41000 7442
rect 38929 7384 38934 7440
rect 38990 7384 41000 7440
rect 38929 7382 41000 7384
rect 38929 7379 38995 7382
rect 40880 7352 41000 7382
rect 8201 7304 13511 7306
rect 8201 7248 8206 7304
rect 8262 7248 13450 7304
rect 13506 7248 13511 7304
rect 8201 7246 13511 7248
rect 8201 7243 8267 7246
rect 13445 7243 13511 7246
rect 13678 7246 21098 7306
rect 21173 7306 21239 7309
rect 32397 7306 32463 7309
rect 21173 7304 32463 7306
rect 21173 7248 21178 7304
rect 21234 7248 32402 7304
rect 32458 7248 32463 7304
rect 21173 7246 32463 7248
rect 0 7170 120 7200
rect 749 7170 815 7173
rect 0 7168 815 7170
rect 0 7112 754 7168
rect 810 7112 815 7168
rect 0 7110 815 7112
rect 0 7080 120 7110
rect 749 7107 815 7110
rect 8385 7170 8451 7173
rect 13678 7170 13738 7246
rect 21173 7243 21239 7246
rect 32397 7243 32463 7246
rect 8385 7168 13738 7170
rect 8385 7112 8390 7168
rect 8446 7112 13738 7168
rect 8385 7110 13738 7112
rect 14733 7170 14799 7173
rect 18505 7170 18571 7173
rect 14733 7168 18571 7170
rect 14733 7112 14738 7168
rect 14794 7112 18510 7168
rect 18566 7112 18571 7168
rect 14733 7110 18571 7112
rect 8385 7107 8451 7110
rect 14733 7107 14799 7110
rect 18505 7107 18571 7110
rect 20621 7170 20687 7173
rect 21725 7170 21791 7173
rect 20621 7168 21791 7170
rect 20621 7112 20626 7168
rect 20682 7112 21730 7168
rect 21786 7112 21791 7168
rect 20621 7110 21791 7112
rect 20621 7107 20687 7110
rect 21725 7107 21791 7110
rect 39389 7170 39455 7173
rect 40880 7170 41000 7200
rect 39389 7168 41000 7170
rect 39389 7112 39394 7168
rect 39450 7112 41000 7168
rect 39389 7110 41000 7112
rect 39389 7107 39455 7110
rect 1946 7104 2262 7105
rect 1946 7040 1952 7104
rect 2016 7040 2032 7104
rect 2096 7040 2112 7104
rect 2176 7040 2192 7104
rect 2256 7040 2262 7104
rect 1946 7039 2262 7040
rect 7946 7104 8262 7105
rect 7946 7040 7952 7104
rect 8016 7040 8032 7104
rect 8096 7040 8112 7104
rect 8176 7040 8192 7104
rect 8256 7040 8262 7104
rect 7946 7039 8262 7040
rect 13946 7104 14262 7105
rect 13946 7040 13952 7104
rect 14016 7040 14032 7104
rect 14096 7040 14112 7104
rect 14176 7040 14192 7104
rect 14256 7040 14262 7104
rect 13946 7039 14262 7040
rect 19946 7104 20262 7105
rect 19946 7040 19952 7104
rect 20016 7040 20032 7104
rect 20096 7040 20112 7104
rect 20176 7040 20192 7104
rect 20256 7040 20262 7104
rect 19946 7039 20262 7040
rect 25946 7104 26262 7105
rect 25946 7040 25952 7104
rect 26016 7040 26032 7104
rect 26096 7040 26112 7104
rect 26176 7040 26192 7104
rect 26256 7040 26262 7104
rect 25946 7039 26262 7040
rect 31946 7104 32262 7105
rect 31946 7040 31952 7104
rect 32016 7040 32032 7104
rect 32096 7040 32112 7104
rect 32176 7040 32192 7104
rect 32256 7040 32262 7104
rect 31946 7039 32262 7040
rect 37946 7104 38262 7105
rect 37946 7040 37952 7104
rect 38016 7040 38032 7104
rect 38096 7040 38112 7104
rect 38176 7040 38192 7104
rect 38256 7040 38262 7104
rect 40880 7080 41000 7110
rect 37946 7039 38262 7040
rect 14365 7034 14431 7037
rect 19517 7034 19583 7037
rect 14365 7032 19583 7034
rect 14365 6976 14370 7032
rect 14426 6976 19522 7032
rect 19578 6976 19583 7032
rect 14365 6974 19583 6976
rect 14365 6971 14431 6974
rect 19517 6971 19583 6974
rect 20529 7034 20595 7037
rect 20529 7032 23490 7034
rect 20529 6976 20534 7032
rect 20590 6976 23490 7032
rect 20529 6974 23490 6976
rect 20529 6971 20595 6974
rect 0 6898 120 6928
rect 933 6898 999 6901
rect 0 6896 999 6898
rect 0 6840 938 6896
rect 994 6840 999 6896
rect 0 6838 999 6840
rect 0 6808 120 6838
rect 933 6835 999 6838
rect 3049 6898 3115 6901
rect 22001 6898 22067 6901
rect 3049 6896 22067 6898
rect 3049 6840 3054 6896
rect 3110 6840 22006 6896
rect 22062 6840 22067 6896
rect 3049 6838 22067 6840
rect 23430 6898 23490 6974
rect 27705 6898 27771 6901
rect 23430 6896 27771 6898
rect 23430 6840 27710 6896
rect 27766 6840 27771 6896
rect 23430 6838 27771 6840
rect 3049 6835 3115 6838
rect 22001 6835 22067 6838
rect 27705 6835 27771 6838
rect 39481 6898 39547 6901
rect 40880 6898 41000 6928
rect 39481 6896 41000 6898
rect 39481 6840 39486 6896
rect 39542 6840 41000 6896
rect 39481 6838 41000 6840
rect 39481 6835 39547 6838
rect 40880 6808 41000 6838
rect 14365 6762 14431 6765
rect 20621 6762 20687 6765
rect 35893 6762 35959 6765
rect 14365 6760 20546 6762
rect 14365 6704 14370 6760
rect 14426 6704 20546 6760
rect 14365 6702 20546 6704
rect 14365 6699 14431 6702
rect 0 6626 120 6656
rect 565 6626 631 6629
rect 0 6624 631 6626
rect 0 6568 570 6624
rect 626 6568 631 6624
rect 0 6566 631 6568
rect 0 6536 120 6566
rect 565 6563 631 6566
rect 3006 6560 3322 6561
rect 3006 6496 3012 6560
rect 3076 6496 3092 6560
rect 3156 6496 3172 6560
rect 3236 6496 3252 6560
rect 3316 6496 3322 6560
rect 3006 6495 3322 6496
rect 9006 6560 9322 6561
rect 9006 6496 9012 6560
rect 9076 6496 9092 6560
rect 9156 6496 9172 6560
rect 9236 6496 9252 6560
rect 9316 6496 9322 6560
rect 9006 6495 9322 6496
rect 15006 6560 15322 6561
rect 15006 6496 15012 6560
rect 15076 6496 15092 6560
rect 15156 6496 15172 6560
rect 15236 6496 15252 6560
rect 15316 6496 15322 6560
rect 15006 6495 15322 6496
rect 14089 6490 14155 6493
rect 14406 6490 14412 6492
rect 14089 6488 14412 6490
rect 14089 6432 14094 6488
rect 14150 6432 14412 6488
rect 14089 6430 14412 6432
rect 14089 6427 14155 6430
rect 14406 6428 14412 6430
rect 14476 6428 14482 6492
rect 16665 6490 16731 6493
rect 19609 6490 19675 6493
rect 16665 6488 19675 6490
rect 16665 6432 16670 6488
rect 16726 6432 19614 6488
rect 19670 6432 19675 6488
rect 16665 6430 19675 6432
rect 16665 6427 16731 6430
rect 19609 6427 19675 6430
rect 19742 6428 19748 6492
rect 19812 6490 19818 6492
rect 20161 6490 20227 6493
rect 19812 6488 20227 6490
rect 19812 6432 20166 6488
rect 20222 6432 20227 6488
rect 19812 6430 20227 6432
rect 19812 6428 19818 6430
rect 20161 6427 20227 6430
rect 0 6354 120 6384
rect 2865 6354 2931 6357
rect 0 6352 2931 6354
rect 0 6296 2870 6352
rect 2926 6296 2931 6352
rect 0 6294 2931 6296
rect 0 6264 120 6294
rect 2865 6291 2931 6294
rect 7373 6354 7439 6357
rect 20345 6354 20411 6357
rect 7373 6352 20411 6354
rect 7373 6296 7378 6352
rect 7434 6296 20350 6352
rect 20406 6296 20411 6352
rect 7373 6294 20411 6296
rect 20486 6354 20546 6702
rect 20621 6760 35959 6762
rect 20621 6704 20626 6760
rect 20682 6704 35898 6760
rect 35954 6704 35959 6760
rect 20621 6702 35959 6704
rect 20621 6699 20687 6702
rect 35893 6699 35959 6702
rect 21725 6626 21791 6629
rect 23105 6626 23171 6629
rect 21725 6624 23171 6626
rect 21725 6568 21730 6624
rect 21786 6568 23110 6624
rect 23166 6568 23171 6624
rect 21725 6566 23171 6568
rect 21725 6563 21791 6566
rect 23105 6563 23171 6566
rect 39573 6626 39639 6629
rect 40880 6626 41000 6656
rect 39573 6624 41000 6626
rect 39573 6568 39578 6624
rect 39634 6568 41000 6624
rect 39573 6566 41000 6568
rect 39573 6563 39639 6566
rect 21006 6560 21322 6561
rect 21006 6496 21012 6560
rect 21076 6496 21092 6560
rect 21156 6496 21172 6560
rect 21236 6496 21252 6560
rect 21316 6496 21322 6560
rect 21006 6495 21322 6496
rect 27006 6560 27322 6561
rect 27006 6496 27012 6560
rect 27076 6496 27092 6560
rect 27156 6496 27172 6560
rect 27236 6496 27252 6560
rect 27316 6496 27322 6560
rect 27006 6495 27322 6496
rect 33006 6560 33322 6561
rect 33006 6496 33012 6560
rect 33076 6496 33092 6560
rect 33156 6496 33172 6560
rect 33236 6496 33252 6560
rect 33316 6496 33322 6560
rect 33006 6495 33322 6496
rect 39006 6560 39322 6561
rect 39006 6496 39012 6560
rect 39076 6496 39092 6560
rect 39156 6496 39172 6560
rect 39236 6496 39252 6560
rect 39316 6496 39322 6560
rect 40880 6536 41000 6566
rect 39006 6495 39322 6496
rect 22645 6490 22711 6493
rect 23657 6490 23723 6493
rect 22645 6488 23723 6490
rect 22645 6432 22650 6488
rect 22706 6432 23662 6488
rect 23718 6432 23723 6488
rect 22645 6430 23723 6432
rect 22645 6427 22711 6430
rect 23657 6427 23723 6430
rect 30373 6354 30439 6357
rect 20486 6352 30439 6354
rect 20486 6296 30378 6352
rect 30434 6296 30439 6352
rect 20486 6294 30439 6296
rect 7373 6291 7439 6294
rect 20345 6291 20411 6294
rect 30373 6291 30439 6294
rect 38653 6354 38719 6357
rect 40880 6354 41000 6384
rect 38653 6352 41000 6354
rect 38653 6296 38658 6352
rect 38714 6296 41000 6352
rect 38653 6294 41000 6296
rect 38653 6291 38719 6294
rect 40880 6264 41000 6294
rect 3417 6218 3483 6221
rect 1718 6216 3483 6218
rect 1718 6160 3422 6216
rect 3478 6160 3483 6216
rect 1718 6158 3483 6160
rect 0 6082 120 6112
rect 1718 6082 1778 6158
rect 3417 6155 3483 6158
rect 10317 6218 10383 6221
rect 32765 6218 32831 6221
rect 10317 6216 32831 6218
rect 10317 6160 10322 6216
rect 10378 6160 32770 6216
rect 32826 6160 32831 6216
rect 10317 6158 32831 6160
rect 10317 6155 10383 6158
rect 32765 6155 32831 6158
rect 0 6022 1778 6082
rect 20345 6082 20411 6085
rect 25313 6082 25379 6085
rect 20345 6080 25379 6082
rect 20345 6024 20350 6080
rect 20406 6024 25318 6080
rect 25374 6024 25379 6080
rect 20345 6022 25379 6024
rect 0 5992 120 6022
rect 20345 6019 20411 6022
rect 25313 6019 25379 6022
rect 39021 6082 39087 6085
rect 40880 6082 41000 6112
rect 39021 6080 41000 6082
rect 39021 6024 39026 6080
rect 39082 6024 41000 6080
rect 39021 6022 41000 6024
rect 39021 6019 39087 6022
rect 1946 6016 2262 6017
rect 1946 5952 1952 6016
rect 2016 5952 2032 6016
rect 2096 5952 2112 6016
rect 2176 5952 2192 6016
rect 2256 5952 2262 6016
rect 1946 5951 2262 5952
rect 7946 6016 8262 6017
rect 7946 5952 7952 6016
rect 8016 5952 8032 6016
rect 8096 5952 8112 6016
rect 8176 5952 8192 6016
rect 8256 5952 8262 6016
rect 7946 5951 8262 5952
rect 13946 6016 14262 6017
rect 13946 5952 13952 6016
rect 14016 5952 14032 6016
rect 14096 5952 14112 6016
rect 14176 5952 14192 6016
rect 14256 5952 14262 6016
rect 13946 5951 14262 5952
rect 19946 6016 20262 6017
rect 19946 5952 19952 6016
rect 20016 5952 20032 6016
rect 20096 5952 20112 6016
rect 20176 5952 20192 6016
rect 20256 5952 20262 6016
rect 19946 5951 20262 5952
rect 25946 6016 26262 6017
rect 25946 5952 25952 6016
rect 26016 5952 26032 6016
rect 26096 5952 26112 6016
rect 26176 5952 26192 6016
rect 26256 5952 26262 6016
rect 25946 5951 26262 5952
rect 31946 6016 32262 6017
rect 31946 5952 31952 6016
rect 32016 5952 32032 6016
rect 32096 5952 32112 6016
rect 32176 5952 32192 6016
rect 32256 5952 32262 6016
rect 31946 5951 32262 5952
rect 37946 6016 38262 6017
rect 37946 5952 37952 6016
rect 38016 5952 38032 6016
rect 38096 5952 38112 6016
rect 38176 5952 38192 6016
rect 38256 5952 38262 6016
rect 40880 5992 41000 6022
rect 37946 5951 38262 5952
rect 20662 5884 20668 5948
rect 20732 5946 20738 5948
rect 21725 5946 21791 5949
rect 20732 5944 21791 5946
rect 20732 5888 21730 5944
rect 21786 5888 21791 5944
rect 20732 5886 21791 5888
rect 20732 5884 20738 5886
rect 21725 5883 21791 5886
rect 0 5810 120 5840
rect 4061 5810 4127 5813
rect 0 5808 4127 5810
rect 0 5752 4066 5808
rect 4122 5752 4127 5808
rect 0 5750 4127 5752
rect 0 5720 120 5750
rect 4061 5747 4127 5750
rect 13353 5810 13419 5813
rect 39205 5810 39271 5813
rect 13353 5808 39271 5810
rect 13353 5752 13358 5808
rect 13414 5752 39210 5808
rect 39266 5752 39271 5808
rect 13353 5750 39271 5752
rect 13353 5747 13419 5750
rect 39205 5747 39271 5750
rect 39481 5810 39547 5813
rect 40880 5810 41000 5840
rect 39481 5808 41000 5810
rect 39481 5752 39486 5808
rect 39542 5752 41000 5808
rect 39481 5750 41000 5752
rect 39481 5747 39547 5750
rect 40880 5720 41000 5750
rect 9949 5674 10015 5677
rect 35985 5674 36051 5677
rect 9949 5672 36051 5674
rect 9949 5616 9954 5672
rect 10010 5616 35990 5672
rect 36046 5616 36051 5672
rect 9949 5614 36051 5616
rect 9949 5611 10015 5614
rect 35985 5611 36051 5614
rect 0 5538 120 5568
rect 1209 5538 1275 5541
rect 0 5536 1275 5538
rect 0 5480 1214 5536
rect 1270 5480 1275 5536
rect 0 5478 1275 5480
rect 0 5448 120 5478
rect 1209 5475 1275 5478
rect 15745 5538 15811 5541
rect 20662 5538 20668 5540
rect 15745 5536 20668 5538
rect 15745 5480 15750 5536
rect 15806 5480 20668 5536
rect 15745 5478 20668 5480
rect 15745 5475 15811 5478
rect 20662 5476 20668 5478
rect 20732 5476 20738 5540
rect 21725 5538 21791 5541
rect 26325 5538 26391 5541
rect 21725 5536 26391 5538
rect 21725 5480 21730 5536
rect 21786 5480 26330 5536
rect 26386 5480 26391 5536
rect 21725 5478 26391 5480
rect 21725 5475 21791 5478
rect 26325 5475 26391 5478
rect 39389 5538 39455 5541
rect 40880 5538 41000 5568
rect 39389 5536 41000 5538
rect 39389 5480 39394 5536
rect 39450 5480 41000 5536
rect 39389 5478 41000 5480
rect 39389 5475 39455 5478
rect 3006 5472 3322 5473
rect 3006 5408 3012 5472
rect 3076 5408 3092 5472
rect 3156 5408 3172 5472
rect 3236 5408 3252 5472
rect 3316 5408 3322 5472
rect 3006 5407 3322 5408
rect 9006 5472 9322 5473
rect 9006 5408 9012 5472
rect 9076 5408 9092 5472
rect 9156 5408 9172 5472
rect 9236 5408 9252 5472
rect 9316 5408 9322 5472
rect 9006 5407 9322 5408
rect 15006 5472 15322 5473
rect 15006 5408 15012 5472
rect 15076 5408 15092 5472
rect 15156 5408 15172 5472
rect 15236 5408 15252 5472
rect 15316 5408 15322 5472
rect 15006 5407 15322 5408
rect 21006 5472 21322 5473
rect 21006 5408 21012 5472
rect 21076 5408 21092 5472
rect 21156 5408 21172 5472
rect 21236 5408 21252 5472
rect 21316 5408 21322 5472
rect 21006 5407 21322 5408
rect 27006 5472 27322 5473
rect 27006 5408 27012 5472
rect 27076 5408 27092 5472
rect 27156 5408 27172 5472
rect 27236 5408 27252 5472
rect 27316 5408 27322 5472
rect 27006 5407 27322 5408
rect 33006 5472 33322 5473
rect 33006 5408 33012 5472
rect 33076 5408 33092 5472
rect 33156 5408 33172 5472
rect 33236 5408 33252 5472
rect 33316 5408 33322 5472
rect 33006 5407 33322 5408
rect 39006 5472 39322 5473
rect 39006 5408 39012 5472
rect 39076 5408 39092 5472
rect 39156 5408 39172 5472
rect 39236 5408 39252 5472
rect 39316 5408 39322 5472
rect 40880 5448 41000 5478
rect 39006 5407 39322 5408
rect 8385 5402 8451 5405
rect 19701 5404 19767 5405
rect 19701 5402 19748 5404
rect 4294 5400 8451 5402
rect 4294 5344 8390 5400
rect 8446 5344 8451 5400
rect 4294 5342 8451 5344
rect 19656 5400 19748 5402
rect 19656 5344 19706 5400
rect 19656 5342 19748 5344
rect 0 5266 120 5296
rect 4294 5266 4354 5342
rect 8385 5339 8451 5342
rect 19701 5340 19748 5342
rect 19812 5340 19818 5404
rect 19701 5339 19767 5340
rect 0 5206 4354 5266
rect 4429 5266 4495 5269
rect 39205 5266 39271 5269
rect 4429 5264 39271 5266
rect 4429 5208 4434 5264
rect 4490 5208 39210 5264
rect 39266 5208 39271 5264
rect 4429 5206 39271 5208
rect 0 5176 120 5206
rect 4429 5203 4495 5206
rect 39205 5203 39271 5206
rect 39389 5266 39455 5269
rect 40880 5266 41000 5296
rect 39389 5264 41000 5266
rect 39389 5208 39394 5264
rect 39450 5208 41000 5264
rect 39389 5206 41000 5208
rect 39389 5203 39455 5206
rect 40880 5176 41000 5206
rect 2773 5130 2839 5133
rect 1534 5128 2839 5130
rect 1534 5072 2778 5128
rect 2834 5072 2839 5128
rect 1534 5070 2839 5072
rect 0 4994 120 5024
rect 1534 4994 1594 5070
rect 2773 5067 2839 5070
rect 9581 5130 9647 5133
rect 27654 5130 27660 5132
rect 9581 5128 27660 5130
rect 9581 5072 9586 5128
rect 9642 5072 27660 5128
rect 9581 5070 27660 5072
rect 9581 5067 9647 5070
rect 27654 5068 27660 5070
rect 27724 5068 27730 5132
rect 0 4934 1594 4994
rect 39021 4994 39087 4997
rect 40880 4994 41000 5024
rect 39021 4992 41000 4994
rect 39021 4936 39026 4992
rect 39082 4936 41000 4992
rect 39021 4934 41000 4936
rect 0 4904 120 4934
rect 39021 4931 39087 4934
rect 1946 4928 2262 4929
rect 1946 4864 1952 4928
rect 2016 4864 2032 4928
rect 2096 4864 2112 4928
rect 2176 4864 2192 4928
rect 2256 4864 2262 4928
rect 1946 4863 2262 4864
rect 7946 4928 8262 4929
rect 7946 4864 7952 4928
rect 8016 4864 8032 4928
rect 8096 4864 8112 4928
rect 8176 4864 8192 4928
rect 8256 4864 8262 4928
rect 7946 4863 8262 4864
rect 13946 4928 14262 4929
rect 13946 4864 13952 4928
rect 14016 4864 14032 4928
rect 14096 4864 14112 4928
rect 14176 4864 14192 4928
rect 14256 4864 14262 4928
rect 13946 4863 14262 4864
rect 19946 4928 20262 4929
rect 19946 4864 19952 4928
rect 20016 4864 20032 4928
rect 20096 4864 20112 4928
rect 20176 4864 20192 4928
rect 20256 4864 20262 4928
rect 19946 4863 20262 4864
rect 25946 4928 26262 4929
rect 25946 4864 25952 4928
rect 26016 4864 26032 4928
rect 26096 4864 26112 4928
rect 26176 4864 26192 4928
rect 26256 4864 26262 4928
rect 25946 4863 26262 4864
rect 31946 4928 32262 4929
rect 31946 4864 31952 4928
rect 32016 4864 32032 4928
rect 32096 4864 32112 4928
rect 32176 4864 32192 4928
rect 32256 4864 32262 4928
rect 31946 4863 32262 4864
rect 37946 4928 38262 4929
rect 37946 4864 37952 4928
rect 38016 4864 38032 4928
rect 38096 4864 38112 4928
rect 38176 4864 38192 4928
rect 38256 4864 38262 4928
rect 40880 4904 41000 4934
rect 37946 4863 38262 4864
rect 20846 4796 20852 4860
rect 20916 4858 20922 4860
rect 21725 4858 21791 4861
rect 20916 4856 21791 4858
rect 20916 4800 21730 4856
rect 21786 4800 21791 4856
rect 20916 4798 21791 4800
rect 20916 4796 20922 4798
rect 21725 4795 21791 4798
rect 0 4722 120 4752
rect 1301 4722 1367 4725
rect 0 4720 1367 4722
rect 0 4664 1306 4720
rect 1362 4664 1367 4720
rect 0 4662 1367 4664
rect 0 4632 120 4662
rect 1301 4659 1367 4662
rect 17493 4722 17559 4725
rect 22277 4722 22343 4725
rect 17493 4720 22343 4722
rect 17493 4664 17498 4720
rect 17554 4664 22282 4720
rect 22338 4664 22343 4720
rect 17493 4662 22343 4664
rect 17493 4659 17559 4662
rect 22277 4659 22343 4662
rect 39481 4722 39547 4725
rect 40880 4722 41000 4752
rect 39481 4720 41000 4722
rect 39481 4664 39486 4720
rect 39542 4664 41000 4720
rect 39481 4662 41000 4664
rect 39481 4659 39547 4662
rect 40880 4632 41000 4662
rect 12065 4586 12131 4589
rect 25497 4586 25563 4589
rect 12065 4584 25563 4586
rect 12065 4528 12070 4584
rect 12126 4528 25502 4584
rect 25558 4528 25563 4584
rect 12065 4526 25563 4528
rect 12065 4523 12131 4526
rect 25497 4523 25563 4526
rect 0 4450 120 4480
rect 2865 4450 2931 4453
rect 0 4448 2931 4450
rect 0 4392 2870 4448
rect 2926 4392 2931 4448
rect 0 4390 2931 4392
rect 0 4360 120 4390
rect 2865 4387 2931 4390
rect 39389 4450 39455 4453
rect 40880 4450 41000 4480
rect 39389 4448 41000 4450
rect 39389 4392 39394 4448
rect 39450 4392 41000 4448
rect 39389 4390 41000 4392
rect 39389 4387 39455 4390
rect 3006 4384 3322 4385
rect 3006 4320 3012 4384
rect 3076 4320 3092 4384
rect 3156 4320 3172 4384
rect 3236 4320 3252 4384
rect 3316 4320 3322 4384
rect 3006 4319 3322 4320
rect 9006 4384 9322 4385
rect 9006 4320 9012 4384
rect 9076 4320 9092 4384
rect 9156 4320 9172 4384
rect 9236 4320 9252 4384
rect 9316 4320 9322 4384
rect 9006 4319 9322 4320
rect 15006 4384 15322 4385
rect 15006 4320 15012 4384
rect 15076 4320 15092 4384
rect 15156 4320 15172 4384
rect 15236 4320 15252 4384
rect 15316 4320 15322 4384
rect 15006 4319 15322 4320
rect 21006 4384 21322 4385
rect 21006 4320 21012 4384
rect 21076 4320 21092 4384
rect 21156 4320 21172 4384
rect 21236 4320 21252 4384
rect 21316 4320 21322 4384
rect 21006 4319 21322 4320
rect 27006 4384 27322 4385
rect 27006 4320 27012 4384
rect 27076 4320 27092 4384
rect 27156 4320 27172 4384
rect 27236 4320 27252 4384
rect 27316 4320 27322 4384
rect 27006 4319 27322 4320
rect 33006 4384 33322 4385
rect 33006 4320 33012 4384
rect 33076 4320 33092 4384
rect 33156 4320 33172 4384
rect 33236 4320 33252 4384
rect 33316 4320 33322 4384
rect 33006 4319 33322 4320
rect 39006 4384 39322 4385
rect 39006 4320 39012 4384
rect 39076 4320 39092 4384
rect 39156 4320 39172 4384
rect 39236 4320 39252 4384
rect 39316 4320 39322 4384
rect 40880 4360 41000 4390
rect 39006 4319 39322 4320
rect 0 4178 120 4208
rect 657 4178 723 4181
rect 0 4176 723 4178
rect 0 4120 662 4176
rect 718 4120 723 4176
rect 0 4118 723 4120
rect 0 4088 120 4118
rect 657 4115 723 4118
rect 3693 4178 3759 4181
rect 21541 4178 21607 4181
rect 3693 4176 21607 4178
rect 3693 4120 3698 4176
rect 3754 4120 21546 4176
rect 21602 4120 21607 4176
rect 3693 4118 21607 4120
rect 3693 4115 3759 4118
rect 21541 4115 21607 4118
rect 39389 4178 39455 4181
rect 40880 4178 41000 4208
rect 39389 4176 41000 4178
rect 39389 4120 39394 4176
rect 39450 4120 41000 4176
rect 39389 4118 41000 4120
rect 39389 4115 39455 4118
rect 40880 4088 41000 4118
rect 3417 4042 3483 4045
rect 1718 4040 3483 4042
rect 1718 3984 3422 4040
rect 3478 3984 3483 4040
rect 1718 3982 3483 3984
rect 0 3906 120 3936
rect 1718 3906 1778 3982
rect 3417 3979 3483 3982
rect 4061 4042 4127 4045
rect 38837 4042 38903 4045
rect 4061 4040 38903 4042
rect 4061 3984 4066 4040
rect 4122 3984 38842 4040
rect 38898 3984 38903 4040
rect 4061 3982 38903 3984
rect 4061 3979 4127 3982
rect 38837 3979 38903 3982
rect 14457 3908 14523 3909
rect 0 3846 1778 3906
rect 0 3816 120 3846
rect 14406 3844 14412 3908
rect 14476 3906 14523 3908
rect 19701 3906 19767 3909
rect 14476 3904 19767 3906
rect 14518 3848 19706 3904
rect 19762 3848 19767 3904
rect 14476 3846 19767 3848
rect 14476 3844 14523 3846
rect 14457 3843 14523 3844
rect 19701 3843 19767 3846
rect 20345 3906 20411 3909
rect 22369 3906 22435 3909
rect 20345 3904 22435 3906
rect 20345 3848 20350 3904
rect 20406 3848 22374 3904
rect 22430 3848 22435 3904
rect 20345 3846 22435 3848
rect 20345 3843 20411 3846
rect 22369 3843 22435 3846
rect 39021 3906 39087 3909
rect 40880 3906 41000 3936
rect 39021 3904 41000 3906
rect 39021 3848 39026 3904
rect 39082 3848 41000 3904
rect 39021 3846 41000 3848
rect 39021 3843 39087 3846
rect 1946 3840 2262 3841
rect 1946 3776 1952 3840
rect 2016 3776 2032 3840
rect 2096 3776 2112 3840
rect 2176 3776 2192 3840
rect 2256 3776 2262 3840
rect 1946 3775 2262 3776
rect 7946 3840 8262 3841
rect 7946 3776 7952 3840
rect 8016 3776 8032 3840
rect 8096 3776 8112 3840
rect 8176 3776 8192 3840
rect 8256 3776 8262 3840
rect 7946 3775 8262 3776
rect 13946 3840 14262 3841
rect 13946 3776 13952 3840
rect 14016 3776 14032 3840
rect 14096 3776 14112 3840
rect 14176 3776 14192 3840
rect 14256 3776 14262 3840
rect 13946 3775 14262 3776
rect 19946 3840 20262 3841
rect 19946 3776 19952 3840
rect 20016 3776 20032 3840
rect 20096 3776 20112 3840
rect 20176 3776 20192 3840
rect 20256 3776 20262 3840
rect 19946 3775 20262 3776
rect 25946 3840 26262 3841
rect 25946 3776 25952 3840
rect 26016 3776 26032 3840
rect 26096 3776 26112 3840
rect 26176 3776 26192 3840
rect 26256 3776 26262 3840
rect 25946 3775 26262 3776
rect 31946 3840 32262 3841
rect 31946 3776 31952 3840
rect 32016 3776 32032 3840
rect 32096 3776 32112 3840
rect 32176 3776 32192 3840
rect 32256 3776 32262 3840
rect 31946 3775 32262 3776
rect 37946 3840 38262 3841
rect 37946 3776 37952 3840
rect 38016 3776 38032 3840
rect 38096 3776 38112 3840
rect 38176 3776 38192 3840
rect 38256 3776 38262 3840
rect 40880 3816 41000 3846
rect 37946 3775 38262 3776
rect 16573 3770 16639 3773
rect 18045 3770 18111 3773
rect 16573 3768 18111 3770
rect 16573 3712 16578 3768
rect 16634 3712 18050 3768
rect 18106 3712 18111 3768
rect 16573 3710 18111 3712
rect 16573 3707 16639 3710
rect 18045 3707 18111 3710
rect 26509 3770 26575 3773
rect 29177 3770 29243 3773
rect 26509 3768 29243 3770
rect 26509 3712 26514 3768
rect 26570 3712 29182 3768
rect 29238 3712 29243 3768
rect 26509 3710 29243 3712
rect 26509 3707 26575 3710
rect 29177 3707 29243 3710
rect 0 3634 120 3664
rect 2773 3634 2839 3637
rect 0 3632 2839 3634
rect 0 3576 2778 3632
rect 2834 3576 2839 3632
rect 0 3574 2839 3576
rect 0 3544 120 3574
rect 2773 3571 2839 3574
rect 3969 3634 4035 3637
rect 39205 3634 39271 3637
rect 3969 3632 39271 3634
rect 3969 3576 3974 3632
rect 4030 3576 39210 3632
rect 39266 3576 39271 3632
rect 3969 3574 39271 3576
rect 3969 3571 4035 3574
rect 39205 3571 39271 3574
rect 39481 3634 39547 3637
rect 40880 3634 41000 3664
rect 39481 3632 41000 3634
rect 39481 3576 39486 3632
rect 39542 3576 41000 3632
rect 39481 3574 41000 3576
rect 39481 3571 39547 3574
rect 40880 3544 41000 3574
rect 3049 3498 3115 3501
rect 17125 3498 17191 3501
rect 26601 3498 26667 3501
rect 38837 3498 38903 3501
rect 3049 3496 17050 3498
rect 3049 3440 3054 3496
rect 3110 3440 17050 3496
rect 3049 3438 17050 3440
rect 3049 3435 3115 3438
rect 0 3362 120 3392
rect 2865 3362 2931 3365
rect 0 3360 2931 3362
rect 0 3304 2870 3360
rect 2926 3304 2931 3360
rect 0 3302 2931 3304
rect 16990 3362 17050 3438
rect 17125 3496 26667 3498
rect 17125 3440 17130 3496
rect 17186 3440 26606 3496
rect 26662 3440 26667 3496
rect 17125 3438 26667 3440
rect 17125 3435 17191 3438
rect 26601 3435 26667 3438
rect 26742 3496 38903 3498
rect 26742 3440 38842 3496
rect 38898 3440 38903 3496
rect 26742 3438 38903 3440
rect 16990 3302 20546 3362
rect 0 3272 120 3302
rect 2865 3299 2931 3302
rect 3006 3296 3322 3297
rect 3006 3232 3012 3296
rect 3076 3232 3092 3296
rect 3156 3232 3172 3296
rect 3236 3232 3252 3296
rect 3316 3232 3322 3296
rect 3006 3231 3322 3232
rect 9006 3296 9322 3297
rect 9006 3232 9012 3296
rect 9076 3232 9092 3296
rect 9156 3232 9172 3296
rect 9236 3232 9252 3296
rect 9316 3232 9322 3296
rect 9006 3231 9322 3232
rect 15006 3296 15322 3297
rect 15006 3232 15012 3296
rect 15076 3232 15092 3296
rect 15156 3232 15172 3296
rect 15236 3232 15252 3296
rect 15316 3232 15322 3296
rect 15006 3231 15322 3232
rect 0 3090 120 3120
rect 1301 3090 1367 3093
rect 0 3088 1367 3090
rect 0 3032 1306 3088
rect 1362 3032 1367 3088
rect 0 3030 1367 3032
rect 0 3000 120 3030
rect 1301 3027 1367 3030
rect 3785 3090 3851 3093
rect 17125 3090 17191 3093
rect 3785 3088 17191 3090
rect 3785 3032 3790 3088
rect 3846 3032 17130 3088
rect 17186 3032 17191 3088
rect 3785 3030 17191 3032
rect 3785 3027 3851 3030
rect 17125 3027 17191 3030
rect 17309 3090 17375 3093
rect 20345 3090 20411 3093
rect 17309 3088 20411 3090
rect 17309 3032 17314 3088
rect 17370 3032 20350 3088
rect 20406 3032 20411 3088
rect 17309 3030 20411 3032
rect 20486 3090 20546 3302
rect 21006 3296 21322 3297
rect 21006 3232 21012 3296
rect 21076 3232 21092 3296
rect 21156 3232 21172 3296
rect 21236 3232 21252 3296
rect 21316 3232 21322 3296
rect 21006 3231 21322 3232
rect 25773 3226 25839 3229
rect 26509 3226 26575 3229
rect 25773 3224 26575 3226
rect 25773 3168 25778 3224
rect 25834 3168 26514 3224
rect 26570 3168 26575 3224
rect 25773 3166 26575 3168
rect 25773 3163 25839 3166
rect 26509 3163 26575 3166
rect 26742 3090 26802 3438
rect 38837 3435 38903 3438
rect 39389 3362 39455 3365
rect 40880 3362 41000 3392
rect 39389 3360 41000 3362
rect 39389 3304 39394 3360
rect 39450 3304 41000 3360
rect 39389 3302 41000 3304
rect 39389 3299 39455 3302
rect 27006 3296 27322 3297
rect 27006 3232 27012 3296
rect 27076 3232 27092 3296
rect 27156 3232 27172 3296
rect 27236 3232 27252 3296
rect 27316 3232 27322 3296
rect 27006 3231 27322 3232
rect 33006 3296 33322 3297
rect 33006 3232 33012 3296
rect 33076 3232 33092 3296
rect 33156 3232 33172 3296
rect 33236 3232 33252 3296
rect 33316 3232 33322 3296
rect 33006 3231 33322 3232
rect 39006 3296 39322 3297
rect 39006 3232 39012 3296
rect 39076 3232 39092 3296
rect 39156 3232 39172 3296
rect 39236 3232 39252 3296
rect 39316 3232 39322 3296
rect 40880 3272 41000 3302
rect 39006 3231 39322 3232
rect 39205 3090 39271 3093
rect 20486 3030 26802 3090
rect 26926 3088 39271 3090
rect 26926 3032 39210 3088
rect 39266 3032 39271 3088
rect 26926 3030 39271 3032
rect 17309 3027 17375 3030
rect 20345 3027 20411 3030
rect 3601 2954 3667 2957
rect 1718 2952 3667 2954
rect 1718 2896 3606 2952
rect 3662 2896 3667 2952
rect 1718 2894 3667 2896
rect 0 2818 120 2848
rect 1718 2818 1778 2894
rect 3601 2891 3667 2894
rect 3877 2954 3943 2957
rect 26926 2954 26986 3030
rect 39205 3027 39271 3030
rect 39389 3090 39455 3093
rect 40880 3090 41000 3120
rect 39389 3088 41000 3090
rect 39389 3032 39394 3088
rect 39450 3032 41000 3088
rect 39389 3030 41000 3032
rect 39389 3027 39455 3030
rect 40880 3000 41000 3030
rect 38469 2954 38535 2957
rect 3877 2952 26986 2954
rect 3877 2896 3882 2952
rect 3938 2896 26986 2952
rect 3877 2894 26986 2896
rect 31710 2952 38535 2954
rect 31710 2896 38474 2952
rect 38530 2896 38535 2952
rect 31710 2894 38535 2896
rect 3877 2891 3943 2894
rect 0 2758 1778 2818
rect 20345 2818 20411 2821
rect 25773 2818 25839 2821
rect 20345 2816 25839 2818
rect 20345 2760 20350 2816
rect 20406 2760 25778 2816
rect 25834 2760 25839 2816
rect 20345 2758 25839 2760
rect 0 2728 120 2758
rect 20345 2755 20411 2758
rect 25773 2755 25839 2758
rect 26601 2818 26667 2821
rect 31710 2818 31770 2894
rect 38469 2891 38535 2894
rect 26601 2816 31770 2818
rect 26601 2760 26606 2816
rect 26662 2760 31770 2816
rect 26601 2758 31770 2760
rect 38837 2818 38903 2821
rect 40880 2818 41000 2848
rect 38837 2816 41000 2818
rect 38837 2760 38842 2816
rect 38898 2760 41000 2816
rect 38837 2758 41000 2760
rect 26601 2755 26667 2758
rect 38837 2755 38903 2758
rect 1946 2752 2262 2753
rect 1946 2688 1952 2752
rect 2016 2688 2032 2752
rect 2096 2688 2112 2752
rect 2176 2688 2192 2752
rect 2256 2688 2262 2752
rect 1946 2687 2262 2688
rect 7946 2752 8262 2753
rect 7946 2688 7952 2752
rect 8016 2688 8032 2752
rect 8096 2688 8112 2752
rect 8176 2688 8192 2752
rect 8256 2688 8262 2752
rect 7946 2687 8262 2688
rect 13946 2752 14262 2753
rect 13946 2688 13952 2752
rect 14016 2688 14032 2752
rect 14096 2688 14112 2752
rect 14176 2688 14192 2752
rect 14256 2688 14262 2752
rect 13946 2687 14262 2688
rect 19946 2752 20262 2753
rect 19946 2688 19952 2752
rect 20016 2688 20032 2752
rect 20096 2688 20112 2752
rect 20176 2688 20192 2752
rect 20256 2688 20262 2752
rect 19946 2687 20262 2688
rect 25946 2752 26262 2753
rect 25946 2688 25952 2752
rect 26016 2688 26032 2752
rect 26096 2688 26112 2752
rect 26176 2688 26192 2752
rect 26256 2688 26262 2752
rect 25946 2687 26262 2688
rect 31946 2752 32262 2753
rect 31946 2688 31952 2752
rect 32016 2688 32032 2752
rect 32096 2688 32112 2752
rect 32176 2688 32192 2752
rect 32256 2688 32262 2752
rect 31946 2687 32262 2688
rect 37946 2752 38262 2753
rect 37946 2688 37952 2752
rect 38016 2688 38032 2752
rect 38096 2688 38112 2752
rect 38176 2688 38192 2752
rect 38256 2688 38262 2752
rect 40880 2728 41000 2758
rect 37946 2687 38262 2688
rect 0 2546 120 2576
rect 1301 2546 1367 2549
rect 0 2544 1367 2546
rect 0 2488 1306 2544
rect 1362 2488 1367 2544
rect 0 2486 1367 2488
rect 0 2456 120 2486
rect 1301 2483 1367 2486
rect 12617 2546 12683 2549
rect 31293 2546 31359 2549
rect 12617 2544 31359 2546
rect 12617 2488 12622 2544
rect 12678 2488 31298 2544
rect 31354 2488 31359 2544
rect 12617 2486 31359 2488
rect 12617 2483 12683 2486
rect 31293 2483 31359 2486
rect 37549 2546 37615 2549
rect 40880 2546 41000 2576
rect 37549 2544 41000 2546
rect 37549 2488 37554 2544
rect 37610 2488 41000 2544
rect 37549 2486 41000 2488
rect 37549 2483 37615 2486
rect 40880 2456 41000 2486
rect 2037 2410 2103 2413
rect 22134 2410 22140 2412
rect 2037 2408 22140 2410
rect 2037 2352 2042 2408
rect 2098 2352 22140 2408
rect 2037 2350 22140 2352
rect 2037 2347 2103 2350
rect 22134 2348 22140 2350
rect 22204 2348 22210 2412
rect 0 2274 120 2304
rect 2865 2274 2931 2277
rect 0 2272 2931 2274
rect 0 2216 2870 2272
rect 2926 2216 2931 2272
rect 0 2214 2931 2216
rect 0 2184 120 2214
rect 2865 2211 2931 2214
rect 39941 2274 40007 2277
rect 40880 2274 41000 2304
rect 39941 2272 41000 2274
rect 39941 2216 39946 2272
rect 40002 2216 41000 2272
rect 39941 2214 41000 2216
rect 39941 2211 40007 2214
rect 3006 2208 3322 2209
rect 3006 2144 3012 2208
rect 3076 2144 3092 2208
rect 3156 2144 3172 2208
rect 3236 2144 3252 2208
rect 3316 2144 3322 2208
rect 3006 2143 3322 2144
rect 9006 2208 9322 2209
rect 9006 2144 9012 2208
rect 9076 2144 9092 2208
rect 9156 2144 9172 2208
rect 9236 2144 9252 2208
rect 9316 2144 9322 2208
rect 9006 2143 9322 2144
rect 15006 2208 15322 2209
rect 15006 2144 15012 2208
rect 15076 2144 15092 2208
rect 15156 2144 15172 2208
rect 15236 2144 15252 2208
rect 15316 2144 15322 2208
rect 15006 2143 15322 2144
rect 21006 2208 21322 2209
rect 21006 2144 21012 2208
rect 21076 2144 21092 2208
rect 21156 2144 21172 2208
rect 21236 2144 21252 2208
rect 21316 2144 21322 2208
rect 21006 2143 21322 2144
rect 27006 2208 27322 2209
rect 27006 2144 27012 2208
rect 27076 2144 27092 2208
rect 27156 2144 27172 2208
rect 27236 2144 27252 2208
rect 27316 2144 27322 2208
rect 27006 2143 27322 2144
rect 33006 2208 33322 2209
rect 33006 2144 33012 2208
rect 33076 2144 33092 2208
rect 33156 2144 33172 2208
rect 33236 2144 33252 2208
rect 33316 2144 33322 2208
rect 33006 2143 33322 2144
rect 39006 2208 39322 2209
rect 39006 2144 39012 2208
rect 39076 2144 39092 2208
rect 39156 2144 39172 2208
rect 39236 2144 39252 2208
rect 39316 2144 39322 2208
rect 40880 2184 41000 2214
rect 39006 2143 39322 2144
rect 0 2002 120 2032
rect 34513 2002 34579 2005
rect 0 2000 34579 2002
rect 0 1944 34518 2000
rect 34574 1944 34579 2000
rect 0 1942 34579 1944
rect 0 1912 120 1942
rect 34513 1939 34579 1942
rect 37825 2002 37891 2005
rect 40880 2002 41000 2032
rect 37825 2000 41000 2002
rect 37825 1944 37830 2000
rect 37886 1944 41000 2000
rect 37825 1942 41000 1944
rect 37825 1939 37891 1942
rect 40880 1912 41000 1942
rect 11053 1866 11119 1869
rect 30281 1866 30347 1869
rect 11053 1864 30347 1866
rect 11053 1808 11058 1864
rect 11114 1808 30286 1864
rect 30342 1808 30347 1864
rect 11053 1806 30347 1808
rect 11053 1803 11119 1806
rect 30281 1803 30347 1806
rect 0 1730 120 1760
rect 1209 1730 1275 1733
rect 0 1728 1275 1730
rect 0 1672 1214 1728
rect 1270 1672 1275 1728
rect 0 1670 1275 1672
rect 0 1640 120 1670
rect 1209 1667 1275 1670
rect 2865 1730 2931 1733
rect 37457 1730 37523 1733
rect 2865 1728 37523 1730
rect 2865 1672 2870 1728
rect 2926 1672 37462 1728
rect 37518 1672 37523 1728
rect 2865 1670 37523 1672
rect 2865 1667 2931 1670
rect 37457 1667 37523 1670
rect 38285 1730 38351 1733
rect 40880 1730 41000 1760
rect 38285 1728 41000 1730
rect 38285 1672 38290 1728
rect 38346 1672 41000 1728
rect 38285 1670 41000 1672
rect 38285 1667 38351 1670
rect 40880 1640 41000 1670
rect 0 1458 120 1488
rect 37733 1458 37799 1461
rect 0 1456 37799 1458
rect 0 1400 37738 1456
rect 37794 1400 37799 1456
rect 0 1398 37799 1400
rect 0 1368 120 1398
rect 37733 1395 37799 1398
rect 38653 1458 38719 1461
rect 40880 1458 41000 1488
rect 38653 1456 41000 1458
rect 38653 1400 38658 1456
rect 38714 1400 41000 1456
rect 38653 1398 41000 1400
rect 38653 1395 38719 1398
rect 40880 1368 41000 1398
rect 15745 98 15811 101
rect 31661 98 31727 101
rect 15745 96 31727 98
rect 15745 40 15750 96
rect 15806 40 31666 96
rect 31722 40 31727 96
rect 15745 38 31727 40
rect 15745 35 15811 38
rect 31661 35 31727 38
<< via3 >>
rect 3012 8732 3076 8736
rect 3012 8676 3016 8732
rect 3016 8676 3072 8732
rect 3072 8676 3076 8732
rect 3012 8672 3076 8676
rect 3092 8732 3156 8736
rect 3092 8676 3096 8732
rect 3096 8676 3152 8732
rect 3152 8676 3156 8732
rect 3092 8672 3156 8676
rect 3172 8732 3236 8736
rect 3172 8676 3176 8732
rect 3176 8676 3232 8732
rect 3232 8676 3236 8732
rect 3172 8672 3236 8676
rect 3252 8732 3316 8736
rect 3252 8676 3256 8732
rect 3256 8676 3312 8732
rect 3312 8676 3316 8732
rect 3252 8672 3316 8676
rect 9012 8732 9076 8736
rect 9012 8676 9016 8732
rect 9016 8676 9072 8732
rect 9072 8676 9076 8732
rect 9012 8672 9076 8676
rect 9092 8732 9156 8736
rect 9092 8676 9096 8732
rect 9096 8676 9152 8732
rect 9152 8676 9156 8732
rect 9092 8672 9156 8676
rect 9172 8732 9236 8736
rect 9172 8676 9176 8732
rect 9176 8676 9232 8732
rect 9232 8676 9236 8732
rect 9172 8672 9236 8676
rect 9252 8732 9316 8736
rect 9252 8676 9256 8732
rect 9256 8676 9312 8732
rect 9312 8676 9316 8732
rect 9252 8672 9316 8676
rect 15012 8732 15076 8736
rect 15012 8676 15016 8732
rect 15016 8676 15072 8732
rect 15072 8676 15076 8732
rect 15012 8672 15076 8676
rect 15092 8732 15156 8736
rect 15092 8676 15096 8732
rect 15096 8676 15152 8732
rect 15152 8676 15156 8732
rect 15092 8672 15156 8676
rect 15172 8732 15236 8736
rect 15172 8676 15176 8732
rect 15176 8676 15232 8732
rect 15232 8676 15236 8732
rect 15172 8672 15236 8676
rect 15252 8732 15316 8736
rect 15252 8676 15256 8732
rect 15256 8676 15312 8732
rect 15312 8676 15316 8732
rect 15252 8672 15316 8676
rect 21012 8732 21076 8736
rect 21012 8676 21016 8732
rect 21016 8676 21072 8732
rect 21072 8676 21076 8732
rect 21012 8672 21076 8676
rect 21092 8732 21156 8736
rect 21092 8676 21096 8732
rect 21096 8676 21152 8732
rect 21152 8676 21156 8732
rect 21092 8672 21156 8676
rect 21172 8732 21236 8736
rect 21172 8676 21176 8732
rect 21176 8676 21232 8732
rect 21232 8676 21236 8732
rect 21172 8672 21236 8676
rect 21252 8732 21316 8736
rect 21252 8676 21256 8732
rect 21256 8676 21312 8732
rect 21312 8676 21316 8732
rect 21252 8672 21316 8676
rect 27012 8732 27076 8736
rect 27012 8676 27016 8732
rect 27016 8676 27072 8732
rect 27072 8676 27076 8732
rect 27012 8672 27076 8676
rect 27092 8732 27156 8736
rect 27092 8676 27096 8732
rect 27096 8676 27152 8732
rect 27152 8676 27156 8732
rect 27092 8672 27156 8676
rect 27172 8732 27236 8736
rect 27172 8676 27176 8732
rect 27176 8676 27232 8732
rect 27232 8676 27236 8732
rect 27172 8672 27236 8676
rect 27252 8732 27316 8736
rect 27252 8676 27256 8732
rect 27256 8676 27312 8732
rect 27312 8676 27316 8732
rect 27252 8672 27316 8676
rect 33012 8732 33076 8736
rect 33012 8676 33016 8732
rect 33016 8676 33072 8732
rect 33072 8676 33076 8732
rect 33012 8672 33076 8676
rect 33092 8732 33156 8736
rect 33092 8676 33096 8732
rect 33096 8676 33152 8732
rect 33152 8676 33156 8732
rect 33092 8672 33156 8676
rect 33172 8732 33236 8736
rect 33172 8676 33176 8732
rect 33176 8676 33232 8732
rect 33232 8676 33236 8732
rect 33172 8672 33236 8676
rect 33252 8732 33316 8736
rect 33252 8676 33256 8732
rect 33256 8676 33312 8732
rect 33312 8676 33316 8732
rect 33252 8672 33316 8676
rect 39012 8732 39076 8736
rect 39012 8676 39016 8732
rect 39016 8676 39072 8732
rect 39072 8676 39076 8732
rect 39012 8672 39076 8676
rect 39092 8732 39156 8736
rect 39092 8676 39096 8732
rect 39096 8676 39152 8732
rect 39152 8676 39156 8732
rect 39092 8672 39156 8676
rect 39172 8732 39236 8736
rect 39172 8676 39176 8732
rect 39176 8676 39232 8732
rect 39232 8676 39236 8732
rect 39172 8672 39236 8676
rect 39252 8732 39316 8736
rect 39252 8676 39256 8732
rect 39256 8676 39312 8732
rect 39312 8676 39316 8732
rect 39252 8672 39316 8676
rect 27660 8332 27724 8396
rect 1952 8188 2016 8192
rect 1952 8132 1956 8188
rect 1956 8132 2012 8188
rect 2012 8132 2016 8188
rect 1952 8128 2016 8132
rect 2032 8188 2096 8192
rect 2032 8132 2036 8188
rect 2036 8132 2092 8188
rect 2092 8132 2096 8188
rect 2032 8128 2096 8132
rect 2112 8188 2176 8192
rect 2112 8132 2116 8188
rect 2116 8132 2172 8188
rect 2172 8132 2176 8188
rect 2112 8128 2176 8132
rect 2192 8188 2256 8192
rect 2192 8132 2196 8188
rect 2196 8132 2252 8188
rect 2252 8132 2256 8188
rect 2192 8128 2256 8132
rect 7952 8188 8016 8192
rect 7952 8132 7956 8188
rect 7956 8132 8012 8188
rect 8012 8132 8016 8188
rect 7952 8128 8016 8132
rect 8032 8188 8096 8192
rect 8032 8132 8036 8188
rect 8036 8132 8092 8188
rect 8092 8132 8096 8188
rect 8032 8128 8096 8132
rect 8112 8188 8176 8192
rect 8112 8132 8116 8188
rect 8116 8132 8172 8188
rect 8172 8132 8176 8188
rect 8112 8128 8176 8132
rect 8192 8188 8256 8192
rect 8192 8132 8196 8188
rect 8196 8132 8252 8188
rect 8252 8132 8256 8188
rect 8192 8128 8256 8132
rect 13952 8188 14016 8192
rect 13952 8132 13956 8188
rect 13956 8132 14012 8188
rect 14012 8132 14016 8188
rect 13952 8128 14016 8132
rect 14032 8188 14096 8192
rect 14032 8132 14036 8188
rect 14036 8132 14092 8188
rect 14092 8132 14096 8188
rect 14032 8128 14096 8132
rect 14112 8188 14176 8192
rect 14112 8132 14116 8188
rect 14116 8132 14172 8188
rect 14172 8132 14176 8188
rect 14112 8128 14176 8132
rect 14192 8188 14256 8192
rect 14192 8132 14196 8188
rect 14196 8132 14252 8188
rect 14252 8132 14256 8188
rect 14192 8128 14256 8132
rect 19952 8188 20016 8192
rect 19952 8132 19956 8188
rect 19956 8132 20012 8188
rect 20012 8132 20016 8188
rect 19952 8128 20016 8132
rect 20032 8188 20096 8192
rect 20032 8132 20036 8188
rect 20036 8132 20092 8188
rect 20092 8132 20096 8188
rect 20032 8128 20096 8132
rect 20112 8188 20176 8192
rect 20112 8132 20116 8188
rect 20116 8132 20172 8188
rect 20172 8132 20176 8188
rect 20112 8128 20176 8132
rect 20192 8188 20256 8192
rect 20192 8132 20196 8188
rect 20196 8132 20252 8188
rect 20252 8132 20256 8188
rect 20192 8128 20256 8132
rect 25952 8188 26016 8192
rect 25952 8132 25956 8188
rect 25956 8132 26012 8188
rect 26012 8132 26016 8188
rect 25952 8128 26016 8132
rect 26032 8188 26096 8192
rect 26032 8132 26036 8188
rect 26036 8132 26092 8188
rect 26092 8132 26096 8188
rect 26032 8128 26096 8132
rect 26112 8188 26176 8192
rect 26112 8132 26116 8188
rect 26116 8132 26172 8188
rect 26172 8132 26176 8188
rect 26112 8128 26176 8132
rect 26192 8188 26256 8192
rect 26192 8132 26196 8188
rect 26196 8132 26252 8188
rect 26252 8132 26256 8188
rect 26192 8128 26256 8132
rect 31952 8188 32016 8192
rect 31952 8132 31956 8188
rect 31956 8132 32012 8188
rect 32012 8132 32016 8188
rect 31952 8128 32016 8132
rect 32032 8188 32096 8192
rect 32032 8132 32036 8188
rect 32036 8132 32092 8188
rect 32092 8132 32096 8188
rect 32032 8128 32096 8132
rect 32112 8188 32176 8192
rect 32112 8132 32116 8188
rect 32116 8132 32172 8188
rect 32172 8132 32176 8188
rect 32112 8128 32176 8132
rect 32192 8188 32256 8192
rect 32192 8132 32196 8188
rect 32196 8132 32252 8188
rect 32252 8132 32256 8188
rect 32192 8128 32256 8132
rect 37952 8188 38016 8192
rect 37952 8132 37956 8188
rect 37956 8132 38012 8188
rect 38012 8132 38016 8188
rect 37952 8128 38016 8132
rect 38032 8188 38096 8192
rect 38032 8132 38036 8188
rect 38036 8132 38092 8188
rect 38092 8132 38096 8188
rect 38032 8128 38096 8132
rect 38112 8188 38176 8192
rect 38112 8132 38116 8188
rect 38116 8132 38172 8188
rect 38172 8132 38176 8188
rect 38112 8128 38176 8132
rect 38192 8188 38256 8192
rect 38192 8132 38196 8188
rect 38196 8132 38252 8188
rect 38252 8132 38256 8188
rect 38192 8128 38256 8132
rect 3012 7644 3076 7648
rect 3012 7588 3016 7644
rect 3016 7588 3072 7644
rect 3072 7588 3076 7644
rect 3012 7584 3076 7588
rect 3092 7644 3156 7648
rect 3092 7588 3096 7644
rect 3096 7588 3152 7644
rect 3152 7588 3156 7644
rect 3092 7584 3156 7588
rect 3172 7644 3236 7648
rect 3172 7588 3176 7644
rect 3176 7588 3232 7644
rect 3232 7588 3236 7644
rect 3172 7584 3236 7588
rect 3252 7644 3316 7648
rect 3252 7588 3256 7644
rect 3256 7588 3312 7644
rect 3312 7588 3316 7644
rect 3252 7584 3316 7588
rect 9012 7644 9076 7648
rect 9012 7588 9016 7644
rect 9016 7588 9072 7644
rect 9072 7588 9076 7644
rect 9012 7584 9076 7588
rect 9092 7644 9156 7648
rect 9092 7588 9096 7644
rect 9096 7588 9152 7644
rect 9152 7588 9156 7644
rect 9092 7584 9156 7588
rect 9172 7644 9236 7648
rect 9172 7588 9176 7644
rect 9176 7588 9232 7644
rect 9232 7588 9236 7644
rect 9172 7584 9236 7588
rect 9252 7644 9316 7648
rect 9252 7588 9256 7644
rect 9256 7588 9312 7644
rect 9312 7588 9316 7644
rect 9252 7584 9316 7588
rect 15012 7644 15076 7648
rect 15012 7588 15016 7644
rect 15016 7588 15072 7644
rect 15072 7588 15076 7644
rect 15012 7584 15076 7588
rect 15092 7644 15156 7648
rect 15092 7588 15096 7644
rect 15096 7588 15152 7644
rect 15152 7588 15156 7644
rect 15092 7584 15156 7588
rect 15172 7644 15236 7648
rect 15172 7588 15176 7644
rect 15176 7588 15232 7644
rect 15232 7588 15236 7644
rect 15172 7584 15236 7588
rect 15252 7644 15316 7648
rect 15252 7588 15256 7644
rect 15256 7588 15312 7644
rect 15312 7588 15316 7644
rect 15252 7584 15316 7588
rect 21012 7644 21076 7648
rect 21012 7588 21016 7644
rect 21016 7588 21072 7644
rect 21072 7588 21076 7644
rect 21012 7584 21076 7588
rect 21092 7644 21156 7648
rect 21092 7588 21096 7644
rect 21096 7588 21152 7644
rect 21152 7588 21156 7644
rect 21092 7584 21156 7588
rect 21172 7644 21236 7648
rect 21172 7588 21176 7644
rect 21176 7588 21232 7644
rect 21232 7588 21236 7644
rect 21172 7584 21236 7588
rect 21252 7644 21316 7648
rect 21252 7588 21256 7644
rect 21256 7588 21312 7644
rect 21312 7588 21316 7644
rect 21252 7584 21316 7588
rect 27012 7644 27076 7648
rect 27012 7588 27016 7644
rect 27016 7588 27072 7644
rect 27072 7588 27076 7644
rect 27012 7584 27076 7588
rect 27092 7644 27156 7648
rect 27092 7588 27096 7644
rect 27096 7588 27152 7644
rect 27152 7588 27156 7644
rect 27092 7584 27156 7588
rect 27172 7644 27236 7648
rect 27172 7588 27176 7644
rect 27176 7588 27232 7644
rect 27232 7588 27236 7644
rect 27172 7584 27236 7588
rect 27252 7644 27316 7648
rect 27252 7588 27256 7644
rect 27256 7588 27312 7644
rect 27312 7588 27316 7644
rect 27252 7584 27316 7588
rect 33012 7644 33076 7648
rect 33012 7588 33016 7644
rect 33016 7588 33072 7644
rect 33072 7588 33076 7644
rect 33012 7584 33076 7588
rect 33092 7644 33156 7648
rect 33092 7588 33096 7644
rect 33096 7588 33152 7644
rect 33152 7588 33156 7644
rect 33092 7584 33156 7588
rect 33172 7644 33236 7648
rect 33172 7588 33176 7644
rect 33176 7588 33232 7644
rect 33232 7588 33236 7644
rect 33172 7584 33236 7588
rect 33252 7644 33316 7648
rect 33252 7588 33256 7644
rect 33256 7588 33312 7644
rect 33312 7588 33316 7644
rect 33252 7584 33316 7588
rect 39012 7644 39076 7648
rect 39012 7588 39016 7644
rect 39016 7588 39072 7644
rect 39072 7588 39076 7644
rect 39012 7584 39076 7588
rect 39092 7644 39156 7648
rect 39092 7588 39096 7644
rect 39096 7588 39152 7644
rect 39152 7588 39156 7644
rect 39092 7584 39156 7588
rect 39172 7644 39236 7648
rect 39172 7588 39176 7644
rect 39176 7588 39232 7644
rect 39232 7588 39236 7644
rect 39172 7584 39236 7588
rect 39252 7644 39316 7648
rect 39252 7588 39256 7644
rect 39256 7588 39312 7644
rect 39312 7588 39316 7644
rect 39252 7584 39316 7588
rect 20852 7516 20916 7580
rect 22140 7516 22204 7580
rect 1952 7100 2016 7104
rect 1952 7044 1956 7100
rect 1956 7044 2012 7100
rect 2012 7044 2016 7100
rect 1952 7040 2016 7044
rect 2032 7100 2096 7104
rect 2032 7044 2036 7100
rect 2036 7044 2092 7100
rect 2092 7044 2096 7100
rect 2032 7040 2096 7044
rect 2112 7100 2176 7104
rect 2112 7044 2116 7100
rect 2116 7044 2172 7100
rect 2172 7044 2176 7100
rect 2112 7040 2176 7044
rect 2192 7100 2256 7104
rect 2192 7044 2196 7100
rect 2196 7044 2252 7100
rect 2252 7044 2256 7100
rect 2192 7040 2256 7044
rect 7952 7100 8016 7104
rect 7952 7044 7956 7100
rect 7956 7044 8012 7100
rect 8012 7044 8016 7100
rect 7952 7040 8016 7044
rect 8032 7100 8096 7104
rect 8032 7044 8036 7100
rect 8036 7044 8092 7100
rect 8092 7044 8096 7100
rect 8032 7040 8096 7044
rect 8112 7100 8176 7104
rect 8112 7044 8116 7100
rect 8116 7044 8172 7100
rect 8172 7044 8176 7100
rect 8112 7040 8176 7044
rect 8192 7100 8256 7104
rect 8192 7044 8196 7100
rect 8196 7044 8252 7100
rect 8252 7044 8256 7100
rect 8192 7040 8256 7044
rect 13952 7100 14016 7104
rect 13952 7044 13956 7100
rect 13956 7044 14012 7100
rect 14012 7044 14016 7100
rect 13952 7040 14016 7044
rect 14032 7100 14096 7104
rect 14032 7044 14036 7100
rect 14036 7044 14092 7100
rect 14092 7044 14096 7100
rect 14032 7040 14096 7044
rect 14112 7100 14176 7104
rect 14112 7044 14116 7100
rect 14116 7044 14172 7100
rect 14172 7044 14176 7100
rect 14112 7040 14176 7044
rect 14192 7100 14256 7104
rect 14192 7044 14196 7100
rect 14196 7044 14252 7100
rect 14252 7044 14256 7100
rect 14192 7040 14256 7044
rect 19952 7100 20016 7104
rect 19952 7044 19956 7100
rect 19956 7044 20012 7100
rect 20012 7044 20016 7100
rect 19952 7040 20016 7044
rect 20032 7100 20096 7104
rect 20032 7044 20036 7100
rect 20036 7044 20092 7100
rect 20092 7044 20096 7100
rect 20032 7040 20096 7044
rect 20112 7100 20176 7104
rect 20112 7044 20116 7100
rect 20116 7044 20172 7100
rect 20172 7044 20176 7100
rect 20112 7040 20176 7044
rect 20192 7100 20256 7104
rect 20192 7044 20196 7100
rect 20196 7044 20252 7100
rect 20252 7044 20256 7100
rect 20192 7040 20256 7044
rect 25952 7100 26016 7104
rect 25952 7044 25956 7100
rect 25956 7044 26012 7100
rect 26012 7044 26016 7100
rect 25952 7040 26016 7044
rect 26032 7100 26096 7104
rect 26032 7044 26036 7100
rect 26036 7044 26092 7100
rect 26092 7044 26096 7100
rect 26032 7040 26096 7044
rect 26112 7100 26176 7104
rect 26112 7044 26116 7100
rect 26116 7044 26172 7100
rect 26172 7044 26176 7100
rect 26112 7040 26176 7044
rect 26192 7100 26256 7104
rect 26192 7044 26196 7100
rect 26196 7044 26252 7100
rect 26252 7044 26256 7100
rect 26192 7040 26256 7044
rect 31952 7100 32016 7104
rect 31952 7044 31956 7100
rect 31956 7044 32012 7100
rect 32012 7044 32016 7100
rect 31952 7040 32016 7044
rect 32032 7100 32096 7104
rect 32032 7044 32036 7100
rect 32036 7044 32092 7100
rect 32092 7044 32096 7100
rect 32032 7040 32096 7044
rect 32112 7100 32176 7104
rect 32112 7044 32116 7100
rect 32116 7044 32172 7100
rect 32172 7044 32176 7100
rect 32112 7040 32176 7044
rect 32192 7100 32256 7104
rect 32192 7044 32196 7100
rect 32196 7044 32252 7100
rect 32252 7044 32256 7100
rect 32192 7040 32256 7044
rect 37952 7100 38016 7104
rect 37952 7044 37956 7100
rect 37956 7044 38012 7100
rect 38012 7044 38016 7100
rect 37952 7040 38016 7044
rect 38032 7100 38096 7104
rect 38032 7044 38036 7100
rect 38036 7044 38092 7100
rect 38092 7044 38096 7100
rect 38032 7040 38096 7044
rect 38112 7100 38176 7104
rect 38112 7044 38116 7100
rect 38116 7044 38172 7100
rect 38172 7044 38176 7100
rect 38112 7040 38176 7044
rect 38192 7100 38256 7104
rect 38192 7044 38196 7100
rect 38196 7044 38252 7100
rect 38252 7044 38256 7100
rect 38192 7040 38256 7044
rect 3012 6556 3076 6560
rect 3012 6500 3016 6556
rect 3016 6500 3072 6556
rect 3072 6500 3076 6556
rect 3012 6496 3076 6500
rect 3092 6556 3156 6560
rect 3092 6500 3096 6556
rect 3096 6500 3152 6556
rect 3152 6500 3156 6556
rect 3092 6496 3156 6500
rect 3172 6556 3236 6560
rect 3172 6500 3176 6556
rect 3176 6500 3232 6556
rect 3232 6500 3236 6556
rect 3172 6496 3236 6500
rect 3252 6556 3316 6560
rect 3252 6500 3256 6556
rect 3256 6500 3312 6556
rect 3312 6500 3316 6556
rect 3252 6496 3316 6500
rect 9012 6556 9076 6560
rect 9012 6500 9016 6556
rect 9016 6500 9072 6556
rect 9072 6500 9076 6556
rect 9012 6496 9076 6500
rect 9092 6556 9156 6560
rect 9092 6500 9096 6556
rect 9096 6500 9152 6556
rect 9152 6500 9156 6556
rect 9092 6496 9156 6500
rect 9172 6556 9236 6560
rect 9172 6500 9176 6556
rect 9176 6500 9232 6556
rect 9232 6500 9236 6556
rect 9172 6496 9236 6500
rect 9252 6556 9316 6560
rect 9252 6500 9256 6556
rect 9256 6500 9312 6556
rect 9312 6500 9316 6556
rect 9252 6496 9316 6500
rect 15012 6556 15076 6560
rect 15012 6500 15016 6556
rect 15016 6500 15072 6556
rect 15072 6500 15076 6556
rect 15012 6496 15076 6500
rect 15092 6556 15156 6560
rect 15092 6500 15096 6556
rect 15096 6500 15152 6556
rect 15152 6500 15156 6556
rect 15092 6496 15156 6500
rect 15172 6556 15236 6560
rect 15172 6500 15176 6556
rect 15176 6500 15232 6556
rect 15232 6500 15236 6556
rect 15172 6496 15236 6500
rect 15252 6556 15316 6560
rect 15252 6500 15256 6556
rect 15256 6500 15312 6556
rect 15312 6500 15316 6556
rect 15252 6496 15316 6500
rect 14412 6428 14476 6492
rect 19748 6428 19812 6492
rect 21012 6556 21076 6560
rect 21012 6500 21016 6556
rect 21016 6500 21072 6556
rect 21072 6500 21076 6556
rect 21012 6496 21076 6500
rect 21092 6556 21156 6560
rect 21092 6500 21096 6556
rect 21096 6500 21152 6556
rect 21152 6500 21156 6556
rect 21092 6496 21156 6500
rect 21172 6556 21236 6560
rect 21172 6500 21176 6556
rect 21176 6500 21232 6556
rect 21232 6500 21236 6556
rect 21172 6496 21236 6500
rect 21252 6556 21316 6560
rect 21252 6500 21256 6556
rect 21256 6500 21312 6556
rect 21312 6500 21316 6556
rect 21252 6496 21316 6500
rect 27012 6556 27076 6560
rect 27012 6500 27016 6556
rect 27016 6500 27072 6556
rect 27072 6500 27076 6556
rect 27012 6496 27076 6500
rect 27092 6556 27156 6560
rect 27092 6500 27096 6556
rect 27096 6500 27152 6556
rect 27152 6500 27156 6556
rect 27092 6496 27156 6500
rect 27172 6556 27236 6560
rect 27172 6500 27176 6556
rect 27176 6500 27232 6556
rect 27232 6500 27236 6556
rect 27172 6496 27236 6500
rect 27252 6556 27316 6560
rect 27252 6500 27256 6556
rect 27256 6500 27312 6556
rect 27312 6500 27316 6556
rect 27252 6496 27316 6500
rect 33012 6556 33076 6560
rect 33012 6500 33016 6556
rect 33016 6500 33072 6556
rect 33072 6500 33076 6556
rect 33012 6496 33076 6500
rect 33092 6556 33156 6560
rect 33092 6500 33096 6556
rect 33096 6500 33152 6556
rect 33152 6500 33156 6556
rect 33092 6496 33156 6500
rect 33172 6556 33236 6560
rect 33172 6500 33176 6556
rect 33176 6500 33232 6556
rect 33232 6500 33236 6556
rect 33172 6496 33236 6500
rect 33252 6556 33316 6560
rect 33252 6500 33256 6556
rect 33256 6500 33312 6556
rect 33312 6500 33316 6556
rect 33252 6496 33316 6500
rect 39012 6556 39076 6560
rect 39012 6500 39016 6556
rect 39016 6500 39072 6556
rect 39072 6500 39076 6556
rect 39012 6496 39076 6500
rect 39092 6556 39156 6560
rect 39092 6500 39096 6556
rect 39096 6500 39152 6556
rect 39152 6500 39156 6556
rect 39092 6496 39156 6500
rect 39172 6556 39236 6560
rect 39172 6500 39176 6556
rect 39176 6500 39232 6556
rect 39232 6500 39236 6556
rect 39172 6496 39236 6500
rect 39252 6556 39316 6560
rect 39252 6500 39256 6556
rect 39256 6500 39312 6556
rect 39312 6500 39316 6556
rect 39252 6496 39316 6500
rect 1952 6012 2016 6016
rect 1952 5956 1956 6012
rect 1956 5956 2012 6012
rect 2012 5956 2016 6012
rect 1952 5952 2016 5956
rect 2032 6012 2096 6016
rect 2032 5956 2036 6012
rect 2036 5956 2092 6012
rect 2092 5956 2096 6012
rect 2032 5952 2096 5956
rect 2112 6012 2176 6016
rect 2112 5956 2116 6012
rect 2116 5956 2172 6012
rect 2172 5956 2176 6012
rect 2112 5952 2176 5956
rect 2192 6012 2256 6016
rect 2192 5956 2196 6012
rect 2196 5956 2252 6012
rect 2252 5956 2256 6012
rect 2192 5952 2256 5956
rect 7952 6012 8016 6016
rect 7952 5956 7956 6012
rect 7956 5956 8012 6012
rect 8012 5956 8016 6012
rect 7952 5952 8016 5956
rect 8032 6012 8096 6016
rect 8032 5956 8036 6012
rect 8036 5956 8092 6012
rect 8092 5956 8096 6012
rect 8032 5952 8096 5956
rect 8112 6012 8176 6016
rect 8112 5956 8116 6012
rect 8116 5956 8172 6012
rect 8172 5956 8176 6012
rect 8112 5952 8176 5956
rect 8192 6012 8256 6016
rect 8192 5956 8196 6012
rect 8196 5956 8252 6012
rect 8252 5956 8256 6012
rect 8192 5952 8256 5956
rect 13952 6012 14016 6016
rect 13952 5956 13956 6012
rect 13956 5956 14012 6012
rect 14012 5956 14016 6012
rect 13952 5952 14016 5956
rect 14032 6012 14096 6016
rect 14032 5956 14036 6012
rect 14036 5956 14092 6012
rect 14092 5956 14096 6012
rect 14032 5952 14096 5956
rect 14112 6012 14176 6016
rect 14112 5956 14116 6012
rect 14116 5956 14172 6012
rect 14172 5956 14176 6012
rect 14112 5952 14176 5956
rect 14192 6012 14256 6016
rect 14192 5956 14196 6012
rect 14196 5956 14252 6012
rect 14252 5956 14256 6012
rect 14192 5952 14256 5956
rect 19952 6012 20016 6016
rect 19952 5956 19956 6012
rect 19956 5956 20012 6012
rect 20012 5956 20016 6012
rect 19952 5952 20016 5956
rect 20032 6012 20096 6016
rect 20032 5956 20036 6012
rect 20036 5956 20092 6012
rect 20092 5956 20096 6012
rect 20032 5952 20096 5956
rect 20112 6012 20176 6016
rect 20112 5956 20116 6012
rect 20116 5956 20172 6012
rect 20172 5956 20176 6012
rect 20112 5952 20176 5956
rect 20192 6012 20256 6016
rect 20192 5956 20196 6012
rect 20196 5956 20252 6012
rect 20252 5956 20256 6012
rect 20192 5952 20256 5956
rect 25952 6012 26016 6016
rect 25952 5956 25956 6012
rect 25956 5956 26012 6012
rect 26012 5956 26016 6012
rect 25952 5952 26016 5956
rect 26032 6012 26096 6016
rect 26032 5956 26036 6012
rect 26036 5956 26092 6012
rect 26092 5956 26096 6012
rect 26032 5952 26096 5956
rect 26112 6012 26176 6016
rect 26112 5956 26116 6012
rect 26116 5956 26172 6012
rect 26172 5956 26176 6012
rect 26112 5952 26176 5956
rect 26192 6012 26256 6016
rect 26192 5956 26196 6012
rect 26196 5956 26252 6012
rect 26252 5956 26256 6012
rect 26192 5952 26256 5956
rect 31952 6012 32016 6016
rect 31952 5956 31956 6012
rect 31956 5956 32012 6012
rect 32012 5956 32016 6012
rect 31952 5952 32016 5956
rect 32032 6012 32096 6016
rect 32032 5956 32036 6012
rect 32036 5956 32092 6012
rect 32092 5956 32096 6012
rect 32032 5952 32096 5956
rect 32112 6012 32176 6016
rect 32112 5956 32116 6012
rect 32116 5956 32172 6012
rect 32172 5956 32176 6012
rect 32112 5952 32176 5956
rect 32192 6012 32256 6016
rect 32192 5956 32196 6012
rect 32196 5956 32252 6012
rect 32252 5956 32256 6012
rect 32192 5952 32256 5956
rect 37952 6012 38016 6016
rect 37952 5956 37956 6012
rect 37956 5956 38012 6012
rect 38012 5956 38016 6012
rect 37952 5952 38016 5956
rect 38032 6012 38096 6016
rect 38032 5956 38036 6012
rect 38036 5956 38092 6012
rect 38092 5956 38096 6012
rect 38032 5952 38096 5956
rect 38112 6012 38176 6016
rect 38112 5956 38116 6012
rect 38116 5956 38172 6012
rect 38172 5956 38176 6012
rect 38112 5952 38176 5956
rect 38192 6012 38256 6016
rect 38192 5956 38196 6012
rect 38196 5956 38252 6012
rect 38252 5956 38256 6012
rect 38192 5952 38256 5956
rect 20668 5884 20732 5948
rect 20668 5476 20732 5540
rect 3012 5468 3076 5472
rect 3012 5412 3016 5468
rect 3016 5412 3072 5468
rect 3072 5412 3076 5468
rect 3012 5408 3076 5412
rect 3092 5468 3156 5472
rect 3092 5412 3096 5468
rect 3096 5412 3152 5468
rect 3152 5412 3156 5468
rect 3092 5408 3156 5412
rect 3172 5468 3236 5472
rect 3172 5412 3176 5468
rect 3176 5412 3232 5468
rect 3232 5412 3236 5468
rect 3172 5408 3236 5412
rect 3252 5468 3316 5472
rect 3252 5412 3256 5468
rect 3256 5412 3312 5468
rect 3312 5412 3316 5468
rect 3252 5408 3316 5412
rect 9012 5468 9076 5472
rect 9012 5412 9016 5468
rect 9016 5412 9072 5468
rect 9072 5412 9076 5468
rect 9012 5408 9076 5412
rect 9092 5468 9156 5472
rect 9092 5412 9096 5468
rect 9096 5412 9152 5468
rect 9152 5412 9156 5468
rect 9092 5408 9156 5412
rect 9172 5468 9236 5472
rect 9172 5412 9176 5468
rect 9176 5412 9232 5468
rect 9232 5412 9236 5468
rect 9172 5408 9236 5412
rect 9252 5468 9316 5472
rect 9252 5412 9256 5468
rect 9256 5412 9312 5468
rect 9312 5412 9316 5468
rect 9252 5408 9316 5412
rect 15012 5468 15076 5472
rect 15012 5412 15016 5468
rect 15016 5412 15072 5468
rect 15072 5412 15076 5468
rect 15012 5408 15076 5412
rect 15092 5468 15156 5472
rect 15092 5412 15096 5468
rect 15096 5412 15152 5468
rect 15152 5412 15156 5468
rect 15092 5408 15156 5412
rect 15172 5468 15236 5472
rect 15172 5412 15176 5468
rect 15176 5412 15232 5468
rect 15232 5412 15236 5468
rect 15172 5408 15236 5412
rect 15252 5468 15316 5472
rect 15252 5412 15256 5468
rect 15256 5412 15312 5468
rect 15312 5412 15316 5468
rect 15252 5408 15316 5412
rect 21012 5468 21076 5472
rect 21012 5412 21016 5468
rect 21016 5412 21072 5468
rect 21072 5412 21076 5468
rect 21012 5408 21076 5412
rect 21092 5468 21156 5472
rect 21092 5412 21096 5468
rect 21096 5412 21152 5468
rect 21152 5412 21156 5468
rect 21092 5408 21156 5412
rect 21172 5468 21236 5472
rect 21172 5412 21176 5468
rect 21176 5412 21232 5468
rect 21232 5412 21236 5468
rect 21172 5408 21236 5412
rect 21252 5468 21316 5472
rect 21252 5412 21256 5468
rect 21256 5412 21312 5468
rect 21312 5412 21316 5468
rect 21252 5408 21316 5412
rect 27012 5468 27076 5472
rect 27012 5412 27016 5468
rect 27016 5412 27072 5468
rect 27072 5412 27076 5468
rect 27012 5408 27076 5412
rect 27092 5468 27156 5472
rect 27092 5412 27096 5468
rect 27096 5412 27152 5468
rect 27152 5412 27156 5468
rect 27092 5408 27156 5412
rect 27172 5468 27236 5472
rect 27172 5412 27176 5468
rect 27176 5412 27232 5468
rect 27232 5412 27236 5468
rect 27172 5408 27236 5412
rect 27252 5468 27316 5472
rect 27252 5412 27256 5468
rect 27256 5412 27312 5468
rect 27312 5412 27316 5468
rect 27252 5408 27316 5412
rect 33012 5468 33076 5472
rect 33012 5412 33016 5468
rect 33016 5412 33072 5468
rect 33072 5412 33076 5468
rect 33012 5408 33076 5412
rect 33092 5468 33156 5472
rect 33092 5412 33096 5468
rect 33096 5412 33152 5468
rect 33152 5412 33156 5468
rect 33092 5408 33156 5412
rect 33172 5468 33236 5472
rect 33172 5412 33176 5468
rect 33176 5412 33232 5468
rect 33232 5412 33236 5468
rect 33172 5408 33236 5412
rect 33252 5468 33316 5472
rect 33252 5412 33256 5468
rect 33256 5412 33312 5468
rect 33312 5412 33316 5468
rect 33252 5408 33316 5412
rect 39012 5468 39076 5472
rect 39012 5412 39016 5468
rect 39016 5412 39072 5468
rect 39072 5412 39076 5468
rect 39012 5408 39076 5412
rect 39092 5468 39156 5472
rect 39092 5412 39096 5468
rect 39096 5412 39152 5468
rect 39152 5412 39156 5468
rect 39092 5408 39156 5412
rect 39172 5468 39236 5472
rect 39172 5412 39176 5468
rect 39176 5412 39232 5468
rect 39232 5412 39236 5468
rect 39172 5408 39236 5412
rect 39252 5468 39316 5472
rect 39252 5412 39256 5468
rect 39256 5412 39312 5468
rect 39312 5412 39316 5468
rect 39252 5408 39316 5412
rect 19748 5400 19812 5404
rect 19748 5344 19762 5400
rect 19762 5344 19812 5400
rect 19748 5340 19812 5344
rect 27660 5068 27724 5132
rect 1952 4924 2016 4928
rect 1952 4868 1956 4924
rect 1956 4868 2012 4924
rect 2012 4868 2016 4924
rect 1952 4864 2016 4868
rect 2032 4924 2096 4928
rect 2032 4868 2036 4924
rect 2036 4868 2092 4924
rect 2092 4868 2096 4924
rect 2032 4864 2096 4868
rect 2112 4924 2176 4928
rect 2112 4868 2116 4924
rect 2116 4868 2172 4924
rect 2172 4868 2176 4924
rect 2112 4864 2176 4868
rect 2192 4924 2256 4928
rect 2192 4868 2196 4924
rect 2196 4868 2252 4924
rect 2252 4868 2256 4924
rect 2192 4864 2256 4868
rect 7952 4924 8016 4928
rect 7952 4868 7956 4924
rect 7956 4868 8012 4924
rect 8012 4868 8016 4924
rect 7952 4864 8016 4868
rect 8032 4924 8096 4928
rect 8032 4868 8036 4924
rect 8036 4868 8092 4924
rect 8092 4868 8096 4924
rect 8032 4864 8096 4868
rect 8112 4924 8176 4928
rect 8112 4868 8116 4924
rect 8116 4868 8172 4924
rect 8172 4868 8176 4924
rect 8112 4864 8176 4868
rect 8192 4924 8256 4928
rect 8192 4868 8196 4924
rect 8196 4868 8252 4924
rect 8252 4868 8256 4924
rect 8192 4864 8256 4868
rect 13952 4924 14016 4928
rect 13952 4868 13956 4924
rect 13956 4868 14012 4924
rect 14012 4868 14016 4924
rect 13952 4864 14016 4868
rect 14032 4924 14096 4928
rect 14032 4868 14036 4924
rect 14036 4868 14092 4924
rect 14092 4868 14096 4924
rect 14032 4864 14096 4868
rect 14112 4924 14176 4928
rect 14112 4868 14116 4924
rect 14116 4868 14172 4924
rect 14172 4868 14176 4924
rect 14112 4864 14176 4868
rect 14192 4924 14256 4928
rect 14192 4868 14196 4924
rect 14196 4868 14252 4924
rect 14252 4868 14256 4924
rect 14192 4864 14256 4868
rect 19952 4924 20016 4928
rect 19952 4868 19956 4924
rect 19956 4868 20012 4924
rect 20012 4868 20016 4924
rect 19952 4864 20016 4868
rect 20032 4924 20096 4928
rect 20032 4868 20036 4924
rect 20036 4868 20092 4924
rect 20092 4868 20096 4924
rect 20032 4864 20096 4868
rect 20112 4924 20176 4928
rect 20112 4868 20116 4924
rect 20116 4868 20172 4924
rect 20172 4868 20176 4924
rect 20112 4864 20176 4868
rect 20192 4924 20256 4928
rect 20192 4868 20196 4924
rect 20196 4868 20252 4924
rect 20252 4868 20256 4924
rect 20192 4864 20256 4868
rect 25952 4924 26016 4928
rect 25952 4868 25956 4924
rect 25956 4868 26012 4924
rect 26012 4868 26016 4924
rect 25952 4864 26016 4868
rect 26032 4924 26096 4928
rect 26032 4868 26036 4924
rect 26036 4868 26092 4924
rect 26092 4868 26096 4924
rect 26032 4864 26096 4868
rect 26112 4924 26176 4928
rect 26112 4868 26116 4924
rect 26116 4868 26172 4924
rect 26172 4868 26176 4924
rect 26112 4864 26176 4868
rect 26192 4924 26256 4928
rect 26192 4868 26196 4924
rect 26196 4868 26252 4924
rect 26252 4868 26256 4924
rect 26192 4864 26256 4868
rect 31952 4924 32016 4928
rect 31952 4868 31956 4924
rect 31956 4868 32012 4924
rect 32012 4868 32016 4924
rect 31952 4864 32016 4868
rect 32032 4924 32096 4928
rect 32032 4868 32036 4924
rect 32036 4868 32092 4924
rect 32092 4868 32096 4924
rect 32032 4864 32096 4868
rect 32112 4924 32176 4928
rect 32112 4868 32116 4924
rect 32116 4868 32172 4924
rect 32172 4868 32176 4924
rect 32112 4864 32176 4868
rect 32192 4924 32256 4928
rect 32192 4868 32196 4924
rect 32196 4868 32252 4924
rect 32252 4868 32256 4924
rect 32192 4864 32256 4868
rect 37952 4924 38016 4928
rect 37952 4868 37956 4924
rect 37956 4868 38012 4924
rect 38012 4868 38016 4924
rect 37952 4864 38016 4868
rect 38032 4924 38096 4928
rect 38032 4868 38036 4924
rect 38036 4868 38092 4924
rect 38092 4868 38096 4924
rect 38032 4864 38096 4868
rect 38112 4924 38176 4928
rect 38112 4868 38116 4924
rect 38116 4868 38172 4924
rect 38172 4868 38176 4924
rect 38112 4864 38176 4868
rect 38192 4924 38256 4928
rect 38192 4868 38196 4924
rect 38196 4868 38252 4924
rect 38252 4868 38256 4924
rect 38192 4864 38256 4868
rect 20852 4796 20916 4860
rect 3012 4380 3076 4384
rect 3012 4324 3016 4380
rect 3016 4324 3072 4380
rect 3072 4324 3076 4380
rect 3012 4320 3076 4324
rect 3092 4380 3156 4384
rect 3092 4324 3096 4380
rect 3096 4324 3152 4380
rect 3152 4324 3156 4380
rect 3092 4320 3156 4324
rect 3172 4380 3236 4384
rect 3172 4324 3176 4380
rect 3176 4324 3232 4380
rect 3232 4324 3236 4380
rect 3172 4320 3236 4324
rect 3252 4380 3316 4384
rect 3252 4324 3256 4380
rect 3256 4324 3312 4380
rect 3312 4324 3316 4380
rect 3252 4320 3316 4324
rect 9012 4380 9076 4384
rect 9012 4324 9016 4380
rect 9016 4324 9072 4380
rect 9072 4324 9076 4380
rect 9012 4320 9076 4324
rect 9092 4380 9156 4384
rect 9092 4324 9096 4380
rect 9096 4324 9152 4380
rect 9152 4324 9156 4380
rect 9092 4320 9156 4324
rect 9172 4380 9236 4384
rect 9172 4324 9176 4380
rect 9176 4324 9232 4380
rect 9232 4324 9236 4380
rect 9172 4320 9236 4324
rect 9252 4380 9316 4384
rect 9252 4324 9256 4380
rect 9256 4324 9312 4380
rect 9312 4324 9316 4380
rect 9252 4320 9316 4324
rect 15012 4380 15076 4384
rect 15012 4324 15016 4380
rect 15016 4324 15072 4380
rect 15072 4324 15076 4380
rect 15012 4320 15076 4324
rect 15092 4380 15156 4384
rect 15092 4324 15096 4380
rect 15096 4324 15152 4380
rect 15152 4324 15156 4380
rect 15092 4320 15156 4324
rect 15172 4380 15236 4384
rect 15172 4324 15176 4380
rect 15176 4324 15232 4380
rect 15232 4324 15236 4380
rect 15172 4320 15236 4324
rect 15252 4380 15316 4384
rect 15252 4324 15256 4380
rect 15256 4324 15312 4380
rect 15312 4324 15316 4380
rect 15252 4320 15316 4324
rect 21012 4380 21076 4384
rect 21012 4324 21016 4380
rect 21016 4324 21072 4380
rect 21072 4324 21076 4380
rect 21012 4320 21076 4324
rect 21092 4380 21156 4384
rect 21092 4324 21096 4380
rect 21096 4324 21152 4380
rect 21152 4324 21156 4380
rect 21092 4320 21156 4324
rect 21172 4380 21236 4384
rect 21172 4324 21176 4380
rect 21176 4324 21232 4380
rect 21232 4324 21236 4380
rect 21172 4320 21236 4324
rect 21252 4380 21316 4384
rect 21252 4324 21256 4380
rect 21256 4324 21312 4380
rect 21312 4324 21316 4380
rect 21252 4320 21316 4324
rect 27012 4380 27076 4384
rect 27012 4324 27016 4380
rect 27016 4324 27072 4380
rect 27072 4324 27076 4380
rect 27012 4320 27076 4324
rect 27092 4380 27156 4384
rect 27092 4324 27096 4380
rect 27096 4324 27152 4380
rect 27152 4324 27156 4380
rect 27092 4320 27156 4324
rect 27172 4380 27236 4384
rect 27172 4324 27176 4380
rect 27176 4324 27232 4380
rect 27232 4324 27236 4380
rect 27172 4320 27236 4324
rect 27252 4380 27316 4384
rect 27252 4324 27256 4380
rect 27256 4324 27312 4380
rect 27312 4324 27316 4380
rect 27252 4320 27316 4324
rect 33012 4380 33076 4384
rect 33012 4324 33016 4380
rect 33016 4324 33072 4380
rect 33072 4324 33076 4380
rect 33012 4320 33076 4324
rect 33092 4380 33156 4384
rect 33092 4324 33096 4380
rect 33096 4324 33152 4380
rect 33152 4324 33156 4380
rect 33092 4320 33156 4324
rect 33172 4380 33236 4384
rect 33172 4324 33176 4380
rect 33176 4324 33232 4380
rect 33232 4324 33236 4380
rect 33172 4320 33236 4324
rect 33252 4380 33316 4384
rect 33252 4324 33256 4380
rect 33256 4324 33312 4380
rect 33312 4324 33316 4380
rect 33252 4320 33316 4324
rect 39012 4380 39076 4384
rect 39012 4324 39016 4380
rect 39016 4324 39072 4380
rect 39072 4324 39076 4380
rect 39012 4320 39076 4324
rect 39092 4380 39156 4384
rect 39092 4324 39096 4380
rect 39096 4324 39152 4380
rect 39152 4324 39156 4380
rect 39092 4320 39156 4324
rect 39172 4380 39236 4384
rect 39172 4324 39176 4380
rect 39176 4324 39232 4380
rect 39232 4324 39236 4380
rect 39172 4320 39236 4324
rect 39252 4380 39316 4384
rect 39252 4324 39256 4380
rect 39256 4324 39312 4380
rect 39312 4324 39316 4380
rect 39252 4320 39316 4324
rect 14412 3904 14476 3908
rect 14412 3848 14462 3904
rect 14462 3848 14476 3904
rect 14412 3844 14476 3848
rect 1952 3836 2016 3840
rect 1952 3780 1956 3836
rect 1956 3780 2012 3836
rect 2012 3780 2016 3836
rect 1952 3776 2016 3780
rect 2032 3836 2096 3840
rect 2032 3780 2036 3836
rect 2036 3780 2092 3836
rect 2092 3780 2096 3836
rect 2032 3776 2096 3780
rect 2112 3836 2176 3840
rect 2112 3780 2116 3836
rect 2116 3780 2172 3836
rect 2172 3780 2176 3836
rect 2112 3776 2176 3780
rect 2192 3836 2256 3840
rect 2192 3780 2196 3836
rect 2196 3780 2252 3836
rect 2252 3780 2256 3836
rect 2192 3776 2256 3780
rect 7952 3836 8016 3840
rect 7952 3780 7956 3836
rect 7956 3780 8012 3836
rect 8012 3780 8016 3836
rect 7952 3776 8016 3780
rect 8032 3836 8096 3840
rect 8032 3780 8036 3836
rect 8036 3780 8092 3836
rect 8092 3780 8096 3836
rect 8032 3776 8096 3780
rect 8112 3836 8176 3840
rect 8112 3780 8116 3836
rect 8116 3780 8172 3836
rect 8172 3780 8176 3836
rect 8112 3776 8176 3780
rect 8192 3836 8256 3840
rect 8192 3780 8196 3836
rect 8196 3780 8252 3836
rect 8252 3780 8256 3836
rect 8192 3776 8256 3780
rect 13952 3836 14016 3840
rect 13952 3780 13956 3836
rect 13956 3780 14012 3836
rect 14012 3780 14016 3836
rect 13952 3776 14016 3780
rect 14032 3836 14096 3840
rect 14032 3780 14036 3836
rect 14036 3780 14092 3836
rect 14092 3780 14096 3836
rect 14032 3776 14096 3780
rect 14112 3836 14176 3840
rect 14112 3780 14116 3836
rect 14116 3780 14172 3836
rect 14172 3780 14176 3836
rect 14112 3776 14176 3780
rect 14192 3836 14256 3840
rect 14192 3780 14196 3836
rect 14196 3780 14252 3836
rect 14252 3780 14256 3836
rect 14192 3776 14256 3780
rect 19952 3836 20016 3840
rect 19952 3780 19956 3836
rect 19956 3780 20012 3836
rect 20012 3780 20016 3836
rect 19952 3776 20016 3780
rect 20032 3836 20096 3840
rect 20032 3780 20036 3836
rect 20036 3780 20092 3836
rect 20092 3780 20096 3836
rect 20032 3776 20096 3780
rect 20112 3836 20176 3840
rect 20112 3780 20116 3836
rect 20116 3780 20172 3836
rect 20172 3780 20176 3836
rect 20112 3776 20176 3780
rect 20192 3836 20256 3840
rect 20192 3780 20196 3836
rect 20196 3780 20252 3836
rect 20252 3780 20256 3836
rect 20192 3776 20256 3780
rect 25952 3836 26016 3840
rect 25952 3780 25956 3836
rect 25956 3780 26012 3836
rect 26012 3780 26016 3836
rect 25952 3776 26016 3780
rect 26032 3836 26096 3840
rect 26032 3780 26036 3836
rect 26036 3780 26092 3836
rect 26092 3780 26096 3836
rect 26032 3776 26096 3780
rect 26112 3836 26176 3840
rect 26112 3780 26116 3836
rect 26116 3780 26172 3836
rect 26172 3780 26176 3836
rect 26112 3776 26176 3780
rect 26192 3836 26256 3840
rect 26192 3780 26196 3836
rect 26196 3780 26252 3836
rect 26252 3780 26256 3836
rect 26192 3776 26256 3780
rect 31952 3836 32016 3840
rect 31952 3780 31956 3836
rect 31956 3780 32012 3836
rect 32012 3780 32016 3836
rect 31952 3776 32016 3780
rect 32032 3836 32096 3840
rect 32032 3780 32036 3836
rect 32036 3780 32092 3836
rect 32092 3780 32096 3836
rect 32032 3776 32096 3780
rect 32112 3836 32176 3840
rect 32112 3780 32116 3836
rect 32116 3780 32172 3836
rect 32172 3780 32176 3836
rect 32112 3776 32176 3780
rect 32192 3836 32256 3840
rect 32192 3780 32196 3836
rect 32196 3780 32252 3836
rect 32252 3780 32256 3836
rect 32192 3776 32256 3780
rect 37952 3836 38016 3840
rect 37952 3780 37956 3836
rect 37956 3780 38012 3836
rect 38012 3780 38016 3836
rect 37952 3776 38016 3780
rect 38032 3836 38096 3840
rect 38032 3780 38036 3836
rect 38036 3780 38092 3836
rect 38092 3780 38096 3836
rect 38032 3776 38096 3780
rect 38112 3836 38176 3840
rect 38112 3780 38116 3836
rect 38116 3780 38172 3836
rect 38172 3780 38176 3836
rect 38112 3776 38176 3780
rect 38192 3836 38256 3840
rect 38192 3780 38196 3836
rect 38196 3780 38252 3836
rect 38252 3780 38256 3836
rect 38192 3776 38256 3780
rect 3012 3292 3076 3296
rect 3012 3236 3016 3292
rect 3016 3236 3072 3292
rect 3072 3236 3076 3292
rect 3012 3232 3076 3236
rect 3092 3292 3156 3296
rect 3092 3236 3096 3292
rect 3096 3236 3152 3292
rect 3152 3236 3156 3292
rect 3092 3232 3156 3236
rect 3172 3292 3236 3296
rect 3172 3236 3176 3292
rect 3176 3236 3232 3292
rect 3232 3236 3236 3292
rect 3172 3232 3236 3236
rect 3252 3292 3316 3296
rect 3252 3236 3256 3292
rect 3256 3236 3312 3292
rect 3312 3236 3316 3292
rect 3252 3232 3316 3236
rect 9012 3292 9076 3296
rect 9012 3236 9016 3292
rect 9016 3236 9072 3292
rect 9072 3236 9076 3292
rect 9012 3232 9076 3236
rect 9092 3292 9156 3296
rect 9092 3236 9096 3292
rect 9096 3236 9152 3292
rect 9152 3236 9156 3292
rect 9092 3232 9156 3236
rect 9172 3292 9236 3296
rect 9172 3236 9176 3292
rect 9176 3236 9232 3292
rect 9232 3236 9236 3292
rect 9172 3232 9236 3236
rect 9252 3292 9316 3296
rect 9252 3236 9256 3292
rect 9256 3236 9312 3292
rect 9312 3236 9316 3292
rect 9252 3232 9316 3236
rect 15012 3292 15076 3296
rect 15012 3236 15016 3292
rect 15016 3236 15072 3292
rect 15072 3236 15076 3292
rect 15012 3232 15076 3236
rect 15092 3292 15156 3296
rect 15092 3236 15096 3292
rect 15096 3236 15152 3292
rect 15152 3236 15156 3292
rect 15092 3232 15156 3236
rect 15172 3292 15236 3296
rect 15172 3236 15176 3292
rect 15176 3236 15232 3292
rect 15232 3236 15236 3292
rect 15172 3232 15236 3236
rect 15252 3292 15316 3296
rect 15252 3236 15256 3292
rect 15256 3236 15312 3292
rect 15312 3236 15316 3292
rect 15252 3232 15316 3236
rect 21012 3292 21076 3296
rect 21012 3236 21016 3292
rect 21016 3236 21072 3292
rect 21072 3236 21076 3292
rect 21012 3232 21076 3236
rect 21092 3292 21156 3296
rect 21092 3236 21096 3292
rect 21096 3236 21152 3292
rect 21152 3236 21156 3292
rect 21092 3232 21156 3236
rect 21172 3292 21236 3296
rect 21172 3236 21176 3292
rect 21176 3236 21232 3292
rect 21232 3236 21236 3292
rect 21172 3232 21236 3236
rect 21252 3292 21316 3296
rect 21252 3236 21256 3292
rect 21256 3236 21312 3292
rect 21312 3236 21316 3292
rect 21252 3232 21316 3236
rect 27012 3292 27076 3296
rect 27012 3236 27016 3292
rect 27016 3236 27072 3292
rect 27072 3236 27076 3292
rect 27012 3232 27076 3236
rect 27092 3292 27156 3296
rect 27092 3236 27096 3292
rect 27096 3236 27152 3292
rect 27152 3236 27156 3292
rect 27092 3232 27156 3236
rect 27172 3292 27236 3296
rect 27172 3236 27176 3292
rect 27176 3236 27232 3292
rect 27232 3236 27236 3292
rect 27172 3232 27236 3236
rect 27252 3292 27316 3296
rect 27252 3236 27256 3292
rect 27256 3236 27312 3292
rect 27312 3236 27316 3292
rect 27252 3232 27316 3236
rect 33012 3292 33076 3296
rect 33012 3236 33016 3292
rect 33016 3236 33072 3292
rect 33072 3236 33076 3292
rect 33012 3232 33076 3236
rect 33092 3292 33156 3296
rect 33092 3236 33096 3292
rect 33096 3236 33152 3292
rect 33152 3236 33156 3292
rect 33092 3232 33156 3236
rect 33172 3292 33236 3296
rect 33172 3236 33176 3292
rect 33176 3236 33232 3292
rect 33232 3236 33236 3292
rect 33172 3232 33236 3236
rect 33252 3292 33316 3296
rect 33252 3236 33256 3292
rect 33256 3236 33312 3292
rect 33312 3236 33316 3292
rect 33252 3232 33316 3236
rect 39012 3292 39076 3296
rect 39012 3236 39016 3292
rect 39016 3236 39072 3292
rect 39072 3236 39076 3292
rect 39012 3232 39076 3236
rect 39092 3292 39156 3296
rect 39092 3236 39096 3292
rect 39096 3236 39152 3292
rect 39152 3236 39156 3292
rect 39092 3232 39156 3236
rect 39172 3292 39236 3296
rect 39172 3236 39176 3292
rect 39176 3236 39232 3292
rect 39232 3236 39236 3292
rect 39172 3232 39236 3236
rect 39252 3292 39316 3296
rect 39252 3236 39256 3292
rect 39256 3236 39312 3292
rect 39312 3236 39316 3292
rect 39252 3232 39316 3236
rect 1952 2748 2016 2752
rect 1952 2692 1956 2748
rect 1956 2692 2012 2748
rect 2012 2692 2016 2748
rect 1952 2688 2016 2692
rect 2032 2748 2096 2752
rect 2032 2692 2036 2748
rect 2036 2692 2092 2748
rect 2092 2692 2096 2748
rect 2032 2688 2096 2692
rect 2112 2748 2176 2752
rect 2112 2692 2116 2748
rect 2116 2692 2172 2748
rect 2172 2692 2176 2748
rect 2112 2688 2176 2692
rect 2192 2748 2256 2752
rect 2192 2692 2196 2748
rect 2196 2692 2252 2748
rect 2252 2692 2256 2748
rect 2192 2688 2256 2692
rect 7952 2748 8016 2752
rect 7952 2692 7956 2748
rect 7956 2692 8012 2748
rect 8012 2692 8016 2748
rect 7952 2688 8016 2692
rect 8032 2748 8096 2752
rect 8032 2692 8036 2748
rect 8036 2692 8092 2748
rect 8092 2692 8096 2748
rect 8032 2688 8096 2692
rect 8112 2748 8176 2752
rect 8112 2692 8116 2748
rect 8116 2692 8172 2748
rect 8172 2692 8176 2748
rect 8112 2688 8176 2692
rect 8192 2748 8256 2752
rect 8192 2692 8196 2748
rect 8196 2692 8252 2748
rect 8252 2692 8256 2748
rect 8192 2688 8256 2692
rect 13952 2748 14016 2752
rect 13952 2692 13956 2748
rect 13956 2692 14012 2748
rect 14012 2692 14016 2748
rect 13952 2688 14016 2692
rect 14032 2748 14096 2752
rect 14032 2692 14036 2748
rect 14036 2692 14092 2748
rect 14092 2692 14096 2748
rect 14032 2688 14096 2692
rect 14112 2748 14176 2752
rect 14112 2692 14116 2748
rect 14116 2692 14172 2748
rect 14172 2692 14176 2748
rect 14112 2688 14176 2692
rect 14192 2748 14256 2752
rect 14192 2692 14196 2748
rect 14196 2692 14252 2748
rect 14252 2692 14256 2748
rect 14192 2688 14256 2692
rect 19952 2748 20016 2752
rect 19952 2692 19956 2748
rect 19956 2692 20012 2748
rect 20012 2692 20016 2748
rect 19952 2688 20016 2692
rect 20032 2748 20096 2752
rect 20032 2692 20036 2748
rect 20036 2692 20092 2748
rect 20092 2692 20096 2748
rect 20032 2688 20096 2692
rect 20112 2748 20176 2752
rect 20112 2692 20116 2748
rect 20116 2692 20172 2748
rect 20172 2692 20176 2748
rect 20112 2688 20176 2692
rect 20192 2748 20256 2752
rect 20192 2692 20196 2748
rect 20196 2692 20252 2748
rect 20252 2692 20256 2748
rect 20192 2688 20256 2692
rect 25952 2748 26016 2752
rect 25952 2692 25956 2748
rect 25956 2692 26012 2748
rect 26012 2692 26016 2748
rect 25952 2688 26016 2692
rect 26032 2748 26096 2752
rect 26032 2692 26036 2748
rect 26036 2692 26092 2748
rect 26092 2692 26096 2748
rect 26032 2688 26096 2692
rect 26112 2748 26176 2752
rect 26112 2692 26116 2748
rect 26116 2692 26172 2748
rect 26172 2692 26176 2748
rect 26112 2688 26176 2692
rect 26192 2748 26256 2752
rect 26192 2692 26196 2748
rect 26196 2692 26252 2748
rect 26252 2692 26256 2748
rect 26192 2688 26256 2692
rect 31952 2748 32016 2752
rect 31952 2692 31956 2748
rect 31956 2692 32012 2748
rect 32012 2692 32016 2748
rect 31952 2688 32016 2692
rect 32032 2748 32096 2752
rect 32032 2692 32036 2748
rect 32036 2692 32092 2748
rect 32092 2692 32096 2748
rect 32032 2688 32096 2692
rect 32112 2748 32176 2752
rect 32112 2692 32116 2748
rect 32116 2692 32172 2748
rect 32172 2692 32176 2748
rect 32112 2688 32176 2692
rect 32192 2748 32256 2752
rect 32192 2692 32196 2748
rect 32196 2692 32252 2748
rect 32252 2692 32256 2748
rect 32192 2688 32256 2692
rect 37952 2748 38016 2752
rect 37952 2692 37956 2748
rect 37956 2692 38012 2748
rect 38012 2692 38016 2748
rect 37952 2688 38016 2692
rect 38032 2748 38096 2752
rect 38032 2692 38036 2748
rect 38036 2692 38092 2748
rect 38092 2692 38096 2748
rect 38032 2688 38096 2692
rect 38112 2748 38176 2752
rect 38112 2692 38116 2748
rect 38116 2692 38172 2748
rect 38172 2692 38176 2748
rect 38112 2688 38176 2692
rect 38192 2748 38256 2752
rect 38192 2692 38196 2748
rect 38196 2692 38252 2748
rect 38252 2692 38256 2748
rect 38192 2688 38256 2692
rect 22140 2348 22204 2412
rect 3012 2204 3076 2208
rect 3012 2148 3016 2204
rect 3016 2148 3072 2204
rect 3072 2148 3076 2204
rect 3012 2144 3076 2148
rect 3092 2204 3156 2208
rect 3092 2148 3096 2204
rect 3096 2148 3152 2204
rect 3152 2148 3156 2204
rect 3092 2144 3156 2148
rect 3172 2204 3236 2208
rect 3172 2148 3176 2204
rect 3176 2148 3232 2204
rect 3232 2148 3236 2204
rect 3172 2144 3236 2148
rect 3252 2204 3316 2208
rect 3252 2148 3256 2204
rect 3256 2148 3312 2204
rect 3312 2148 3316 2204
rect 3252 2144 3316 2148
rect 9012 2204 9076 2208
rect 9012 2148 9016 2204
rect 9016 2148 9072 2204
rect 9072 2148 9076 2204
rect 9012 2144 9076 2148
rect 9092 2204 9156 2208
rect 9092 2148 9096 2204
rect 9096 2148 9152 2204
rect 9152 2148 9156 2204
rect 9092 2144 9156 2148
rect 9172 2204 9236 2208
rect 9172 2148 9176 2204
rect 9176 2148 9232 2204
rect 9232 2148 9236 2204
rect 9172 2144 9236 2148
rect 9252 2204 9316 2208
rect 9252 2148 9256 2204
rect 9256 2148 9312 2204
rect 9312 2148 9316 2204
rect 9252 2144 9316 2148
rect 15012 2204 15076 2208
rect 15012 2148 15016 2204
rect 15016 2148 15072 2204
rect 15072 2148 15076 2204
rect 15012 2144 15076 2148
rect 15092 2204 15156 2208
rect 15092 2148 15096 2204
rect 15096 2148 15152 2204
rect 15152 2148 15156 2204
rect 15092 2144 15156 2148
rect 15172 2204 15236 2208
rect 15172 2148 15176 2204
rect 15176 2148 15232 2204
rect 15232 2148 15236 2204
rect 15172 2144 15236 2148
rect 15252 2204 15316 2208
rect 15252 2148 15256 2204
rect 15256 2148 15312 2204
rect 15312 2148 15316 2204
rect 15252 2144 15316 2148
rect 21012 2204 21076 2208
rect 21012 2148 21016 2204
rect 21016 2148 21072 2204
rect 21072 2148 21076 2204
rect 21012 2144 21076 2148
rect 21092 2204 21156 2208
rect 21092 2148 21096 2204
rect 21096 2148 21152 2204
rect 21152 2148 21156 2204
rect 21092 2144 21156 2148
rect 21172 2204 21236 2208
rect 21172 2148 21176 2204
rect 21176 2148 21232 2204
rect 21232 2148 21236 2204
rect 21172 2144 21236 2148
rect 21252 2204 21316 2208
rect 21252 2148 21256 2204
rect 21256 2148 21312 2204
rect 21312 2148 21316 2204
rect 21252 2144 21316 2148
rect 27012 2204 27076 2208
rect 27012 2148 27016 2204
rect 27016 2148 27072 2204
rect 27072 2148 27076 2204
rect 27012 2144 27076 2148
rect 27092 2204 27156 2208
rect 27092 2148 27096 2204
rect 27096 2148 27152 2204
rect 27152 2148 27156 2204
rect 27092 2144 27156 2148
rect 27172 2204 27236 2208
rect 27172 2148 27176 2204
rect 27176 2148 27232 2204
rect 27232 2148 27236 2204
rect 27172 2144 27236 2148
rect 27252 2204 27316 2208
rect 27252 2148 27256 2204
rect 27256 2148 27312 2204
rect 27312 2148 27316 2204
rect 27252 2144 27316 2148
rect 33012 2204 33076 2208
rect 33012 2148 33016 2204
rect 33016 2148 33072 2204
rect 33072 2148 33076 2204
rect 33012 2144 33076 2148
rect 33092 2204 33156 2208
rect 33092 2148 33096 2204
rect 33096 2148 33152 2204
rect 33152 2148 33156 2204
rect 33092 2144 33156 2148
rect 33172 2204 33236 2208
rect 33172 2148 33176 2204
rect 33176 2148 33232 2204
rect 33232 2148 33236 2204
rect 33172 2144 33236 2148
rect 33252 2204 33316 2208
rect 33252 2148 33256 2204
rect 33256 2148 33312 2204
rect 33312 2148 33316 2204
rect 33252 2144 33316 2148
rect 39012 2204 39076 2208
rect 39012 2148 39016 2204
rect 39016 2148 39072 2204
rect 39072 2148 39076 2204
rect 39012 2144 39076 2148
rect 39092 2204 39156 2208
rect 39092 2148 39096 2204
rect 39096 2148 39152 2204
rect 39152 2148 39156 2204
rect 39092 2144 39156 2148
rect 39172 2204 39236 2208
rect 39172 2148 39176 2204
rect 39176 2148 39232 2204
rect 39232 2148 39236 2204
rect 39172 2144 39236 2148
rect 39252 2204 39316 2208
rect 39252 2148 39256 2204
rect 39256 2148 39312 2204
rect 39312 2148 39316 2204
rect 39252 2144 39316 2148
<< metal4 >>
rect 1944 8192 2264 11250
rect 1944 8128 1952 8192
rect 2016 8128 2032 8192
rect 2096 8128 2112 8192
rect 2176 8128 2192 8192
rect 2256 8128 2264 8192
rect 1944 7104 2264 8128
rect 1944 7040 1952 7104
rect 2016 7040 2032 7104
rect 2096 7040 2112 7104
rect 2176 7040 2192 7104
rect 2256 7040 2264 7104
rect 1944 6016 2264 7040
rect 1944 5952 1952 6016
rect 2016 5952 2032 6016
rect 2096 5952 2112 6016
rect 2176 5952 2192 6016
rect 2256 5952 2264 6016
rect 1944 4928 2264 5952
rect 1944 4864 1952 4928
rect 2016 4864 2032 4928
rect 2096 4864 2112 4928
rect 2176 4864 2192 4928
rect 2256 4864 2264 4928
rect 1944 3840 2264 4864
rect 1944 3776 1952 3840
rect 2016 3776 2032 3840
rect 2096 3776 2112 3840
rect 2176 3776 2192 3840
rect 2256 3776 2264 3840
rect 1944 2752 2264 3776
rect 1944 2688 1952 2752
rect 2016 2688 2032 2752
rect 2096 2688 2112 2752
rect 2176 2688 2192 2752
rect 2256 2688 2264 2752
rect 1944 0 2264 2688
rect 3004 8736 3324 11250
rect 3004 8672 3012 8736
rect 3076 8672 3092 8736
rect 3156 8672 3172 8736
rect 3236 8672 3252 8736
rect 3316 8672 3324 8736
rect 3004 7648 3324 8672
rect 3004 7584 3012 7648
rect 3076 7584 3092 7648
rect 3156 7584 3172 7648
rect 3236 7584 3252 7648
rect 3316 7584 3324 7648
rect 3004 6560 3324 7584
rect 3004 6496 3012 6560
rect 3076 6496 3092 6560
rect 3156 6496 3172 6560
rect 3236 6496 3252 6560
rect 3316 6496 3324 6560
rect 3004 5472 3324 6496
rect 3004 5408 3012 5472
rect 3076 5408 3092 5472
rect 3156 5408 3172 5472
rect 3236 5408 3252 5472
rect 3316 5408 3324 5472
rect 3004 4384 3324 5408
rect 3004 4320 3012 4384
rect 3076 4320 3092 4384
rect 3156 4320 3172 4384
rect 3236 4320 3252 4384
rect 3316 4320 3324 4384
rect 3004 3296 3324 4320
rect 3004 3232 3012 3296
rect 3076 3232 3092 3296
rect 3156 3232 3172 3296
rect 3236 3232 3252 3296
rect 3316 3232 3324 3296
rect 3004 2208 3324 3232
rect 3004 2144 3012 2208
rect 3076 2144 3092 2208
rect 3156 2144 3172 2208
rect 3236 2144 3252 2208
rect 3316 2144 3324 2208
rect 3004 0 3324 2144
rect 7944 8192 8264 11250
rect 7944 8128 7952 8192
rect 8016 8128 8032 8192
rect 8096 8128 8112 8192
rect 8176 8128 8192 8192
rect 8256 8128 8264 8192
rect 7944 7104 8264 8128
rect 7944 7040 7952 7104
rect 8016 7040 8032 7104
rect 8096 7040 8112 7104
rect 8176 7040 8192 7104
rect 8256 7040 8264 7104
rect 7944 6016 8264 7040
rect 7944 5952 7952 6016
rect 8016 5952 8032 6016
rect 8096 5952 8112 6016
rect 8176 5952 8192 6016
rect 8256 5952 8264 6016
rect 7944 4928 8264 5952
rect 7944 4864 7952 4928
rect 8016 4864 8032 4928
rect 8096 4864 8112 4928
rect 8176 4864 8192 4928
rect 8256 4864 8264 4928
rect 7944 3840 8264 4864
rect 7944 3776 7952 3840
rect 8016 3776 8032 3840
rect 8096 3776 8112 3840
rect 8176 3776 8192 3840
rect 8256 3776 8264 3840
rect 7944 2752 8264 3776
rect 7944 2688 7952 2752
rect 8016 2688 8032 2752
rect 8096 2688 8112 2752
rect 8176 2688 8192 2752
rect 8256 2688 8264 2752
rect 7944 0 8264 2688
rect 9004 8736 9324 11250
rect 9004 8672 9012 8736
rect 9076 8672 9092 8736
rect 9156 8672 9172 8736
rect 9236 8672 9252 8736
rect 9316 8672 9324 8736
rect 9004 7648 9324 8672
rect 9004 7584 9012 7648
rect 9076 7584 9092 7648
rect 9156 7584 9172 7648
rect 9236 7584 9252 7648
rect 9316 7584 9324 7648
rect 9004 6560 9324 7584
rect 9004 6496 9012 6560
rect 9076 6496 9092 6560
rect 9156 6496 9172 6560
rect 9236 6496 9252 6560
rect 9316 6496 9324 6560
rect 9004 5472 9324 6496
rect 9004 5408 9012 5472
rect 9076 5408 9092 5472
rect 9156 5408 9172 5472
rect 9236 5408 9252 5472
rect 9316 5408 9324 5472
rect 9004 4384 9324 5408
rect 9004 4320 9012 4384
rect 9076 4320 9092 4384
rect 9156 4320 9172 4384
rect 9236 4320 9252 4384
rect 9316 4320 9324 4384
rect 9004 3296 9324 4320
rect 9004 3232 9012 3296
rect 9076 3232 9092 3296
rect 9156 3232 9172 3296
rect 9236 3232 9252 3296
rect 9316 3232 9324 3296
rect 9004 2208 9324 3232
rect 9004 2144 9012 2208
rect 9076 2144 9092 2208
rect 9156 2144 9172 2208
rect 9236 2144 9252 2208
rect 9316 2144 9324 2208
rect 9004 0 9324 2144
rect 13944 8192 14264 11250
rect 13944 8128 13952 8192
rect 14016 8128 14032 8192
rect 14096 8128 14112 8192
rect 14176 8128 14192 8192
rect 14256 8128 14264 8192
rect 13944 7104 14264 8128
rect 13944 7040 13952 7104
rect 14016 7040 14032 7104
rect 14096 7040 14112 7104
rect 14176 7040 14192 7104
rect 14256 7040 14264 7104
rect 13944 6016 14264 7040
rect 15004 8736 15324 11250
rect 15004 8672 15012 8736
rect 15076 8672 15092 8736
rect 15156 8672 15172 8736
rect 15236 8672 15252 8736
rect 15316 8672 15324 8736
rect 15004 7648 15324 8672
rect 15004 7584 15012 7648
rect 15076 7584 15092 7648
rect 15156 7584 15172 7648
rect 15236 7584 15252 7648
rect 15316 7584 15324 7648
rect 15004 6560 15324 7584
rect 15004 6496 15012 6560
rect 15076 6496 15092 6560
rect 15156 6496 15172 6560
rect 15236 6496 15252 6560
rect 15316 6496 15324 6560
rect 14411 6492 14477 6493
rect 14411 6428 14412 6492
rect 14476 6428 14477 6492
rect 14411 6427 14477 6428
rect 13944 5952 13952 6016
rect 14016 5952 14032 6016
rect 14096 5952 14112 6016
rect 14176 5952 14192 6016
rect 14256 5952 14264 6016
rect 13944 4928 14264 5952
rect 13944 4864 13952 4928
rect 14016 4864 14032 4928
rect 14096 4864 14112 4928
rect 14176 4864 14192 4928
rect 14256 4864 14264 4928
rect 13944 3840 14264 4864
rect 14414 3909 14474 6427
rect 15004 5472 15324 6496
rect 19944 8192 20264 11250
rect 19944 8128 19952 8192
rect 20016 8128 20032 8192
rect 20096 8128 20112 8192
rect 20176 8128 20192 8192
rect 20256 8128 20264 8192
rect 19944 7104 20264 8128
rect 21004 8736 21324 11250
rect 21004 8672 21012 8736
rect 21076 8672 21092 8736
rect 21156 8672 21172 8736
rect 21236 8672 21252 8736
rect 21316 8672 21324 8736
rect 21004 7648 21324 8672
rect 21004 7584 21012 7648
rect 21076 7584 21092 7648
rect 21156 7584 21172 7648
rect 21236 7584 21252 7648
rect 21316 7584 21324 7648
rect 20851 7580 20917 7581
rect 20851 7516 20852 7580
rect 20916 7516 20917 7580
rect 20851 7515 20917 7516
rect 19944 7040 19952 7104
rect 20016 7040 20032 7104
rect 20096 7040 20112 7104
rect 20176 7040 20192 7104
rect 20256 7040 20264 7104
rect 19747 6492 19813 6493
rect 19747 6428 19748 6492
rect 19812 6428 19813 6492
rect 19747 6427 19813 6428
rect 15004 5408 15012 5472
rect 15076 5408 15092 5472
rect 15156 5408 15172 5472
rect 15236 5408 15252 5472
rect 15316 5408 15324 5472
rect 15004 4384 15324 5408
rect 19750 5405 19810 6427
rect 19944 6016 20264 7040
rect 19944 5952 19952 6016
rect 20016 5952 20032 6016
rect 20096 5952 20112 6016
rect 20176 5952 20192 6016
rect 20256 5952 20264 6016
rect 19747 5404 19813 5405
rect 19747 5340 19748 5404
rect 19812 5340 19813 5404
rect 19747 5339 19813 5340
rect 15004 4320 15012 4384
rect 15076 4320 15092 4384
rect 15156 4320 15172 4384
rect 15236 4320 15252 4384
rect 15316 4320 15324 4384
rect 14411 3908 14477 3909
rect 14411 3844 14412 3908
rect 14476 3844 14477 3908
rect 14411 3843 14477 3844
rect 13944 3776 13952 3840
rect 14016 3776 14032 3840
rect 14096 3776 14112 3840
rect 14176 3776 14192 3840
rect 14256 3776 14264 3840
rect 13944 2752 14264 3776
rect 13944 2688 13952 2752
rect 14016 2688 14032 2752
rect 14096 2688 14112 2752
rect 14176 2688 14192 2752
rect 14256 2688 14264 2752
rect 13944 0 14264 2688
rect 15004 3296 15324 4320
rect 15004 3232 15012 3296
rect 15076 3232 15092 3296
rect 15156 3232 15172 3296
rect 15236 3232 15252 3296
rect 15316 3232 15324 3296
rect 15004 2208 15324 3232
rect 15004 2144 15012 2208
rect 15076 2144 15092 2208
rect 15156 2144 15172 2208
rect 15236 2144 15252 2208
rect 15316 2144 15324 2208
rect 15004 0 15324 2144
rect 19944 4928 20264 5952
rect 20667 5948 20733 5949
rect 20667 5884 20668 5948
rect 20732 5884 20733 5948
rect 20667 5883 20733 5884
rect 20670 5541 20730 5883
rect 20667 5540 20733 5541
rect 20667 5476 20668 5540
rect 20732 5476 20733 5540
rect 20667 5475 20733 5476
rect 19944 4864 19952 4928
rect 20016 4864 20032 4928
rect 20096 4864 20112 4928
rect 20176 4864 20192 4928
rect 20256 4864 20264 4928
rect 19944 3840 20264 4864
rect 20854 4861 20914 7515
rect 21004 6560 21324 7584
rect 25944 8192 26264 11250
rect 25944 8128 25952 8192
rect 26016 8128 26032 8192
rect 26096 8128 26112 8192
rect 26176 8128 26192 8192
rect 26256 8128 26264 8192
rect 22139 7580 22205 7581
rect 22139 7516 22140 7580
rect 22204 7516 22205 7580
rect 22139 7515 22205 7516
rect 21004 6496 21012 6560
rect 21076 6496 21092 6560
rect 21156 6496 21172 6560
rect 21236 6496 21252 6560
rect 21316 6496 21324 6560
rect 21004 5472 21324 6496
rect 21004 5408 21012 5472
rect 21076 5408 21092 5472
rect 21156 5408 21172 5472
rect 21236 5408 21252 5472
rect 21316 5408 21324 5472
rect 20851 4860 20917 4861
rect 20851 4796 20852 4860
rect 20916 4796 20917 4860
rect 20851 4795 20917 4796
rect 19944 3776 19952 3840
rect 20016 3776 20032 3840
rect 20096 3776 20112 3840
rect 20176 3776 20192 3840
rect 20256 3776 20264 3840
rect 19944 2752 20264 3776
rect 19944 2688 19952 2752
rect 20016 2688 20032 2752
rect 20096 2688 20112 2752
rect 20176 2688 20192 2752
rect 20256 2688 20264 2752
rect 19944 0 20264 2688
rect 21004 4384 21324 5408
rect 21004 4320 21012 4384
rect 21076 4320 21092 4384
rect 21156 4320 21172 4384
rect 21236 4320 21252 4384
rect 21316 4320 21324 4384
rect 21004 3296 21324 4320
rect 21004 3232 21012 3296
rect 21076 3232 21092 3296
rect 21156 3232 21172 3296
rect 21236 3232 21252 3296
rect 21316 3232 21324 3296
rect 21004 2208 21324 3232
rect 22142 2413 22202 7515
rect 25944 7104 26264 8128
rect 25944 7040 25952 7104
rect 26016 7040 26032 7104
rect 26096 7040 26112 7104
rect 26176 7040 26192 7104
rect 26256 7040 26264 7104
rect 25944 6016 26264 7040
rect 25944 5952 25952 6016
rect 26016 5952 26032 6016
rect 26096 5952 26112 6016
rect 26176 5952 26192 6016
rect 26256 5952 26264 6016
rect 25944 4928 26264 5952
rect 25944 4864 25952 4928
rect 26016 4864 26032 4928
rect 26096 4864 26112 4928
rect 26176 4864 26192 4928
rect 26256 4864 26264 4928
rect 25944 3840 26264 4864
rect 25944 3776 25952 3840
rect 26016 3776 26032 3840
rect 26096 3776 26112 3840
rect 26176 3776 26192 3840
rect 26256 3776 26264 3840
rect 25944 2752 26264 3776
rect 25944 2688 25952 2752
rect 26016 2688 26032 2752
rect 26096 2688 26112 2752
rect 26176 2688 26192 2752
rect 26256 2688 26264 2752
rect 22139 2412 22205 2413
rect 22139 2348 22140 2412
rect 22204 2348 22205 2412
rect 22139 2347 22205 2348
rect 21004 2144 21012 2208
rect 21076 2144 21092 2208
rect 21156 2144 21172 2208
rect 21236 2144 21252 2208
rect 21316 2144 21324 2208
rect 21004 0 21324 2144
rect 25944 0 26264 2688
rect 27004 8736 27324 11250
rect 27004 8672 27012 8736
rect 27076 8672 27092 8736
rect 27156 8672 27172 8736
rect 27236 8672 27252 8736
rect 27316 8672 27324 8736
rect 27004 7648 27324 8672
rect 27659 8396 27725 8397
rect 27659 8332 27660 8396
rect 27724 8332 27725 8396
rect 27659 8331 27725 8332
rect 27004 7584 27012 7648
rect 27076 7584 27092 7648
rect 27156 7584 27172 7648
rect 27236 7584 27252 7648
rect 27316 7584 27324 7648
rect 27004 6560 27324 7584
rect 27004 6496 27012 6560
rect 27076 6496 27092 6560
rect 27156 6496 27172 6560
rect 27236 6496 27252 6560
rect 27316 6496 27324 6560
rect 27004 5472 27324 6496
rect 27004 5408 27012 5472
rect 27076 5408 27092 5472
rect 27156 5408 27172 5472
rect 27236 5408 27252 5472
rect 27316 5408 27324 5472
rect 27004 4384 27324 5408
rect 27662 5133 27722 8331
rect 31944 8192 32264 11250
rect 31944 8128 31952 8192
rect 32016 8128 32032 8192
rect 32096 8128 32112 8192
rect 32176 8128 32192 8192
rect 32256 8128 32264 8192
rect 31944 7104 32264 8128
rect 31944 7040 31952 7104
rect 32016 7040 32032 7104
rect 32096 7040 32112 7104
rect 32176 7040 32192 7104
rect 32256 7040 32264 7104
rect 31944 6016 32264 7040
rect 31944 5952 31952 6016
rect 32016 5952 32032 6016
rect 32096 5952 32112 6016
rect 32176 5952 32192 6016
rect 32256 5952 32264 6016
rect 27659 5132 27725 5133
rect 27659 5068 27660 5132
rect 27724 5068 27725 5132
rect 27659 5067 27725 5068
rect 27004 4320 27012 4384
rect 27076 4320 27092 4384
rect 27156 4320 27172 4384
rect 27236 4320 27252 4384
rect 27316 4320 27324 4384
rect 27004 3296 27324 4320
rect 27004 3232 27012 3296
rect 27076 3232 27092 3296
rect 27156 3232 27172 3296
rect 27236 3232 27252 3296
rect 27316 3232 27324 3296
rect 27004 2208 27324 3232
rect 27004 2144 27012 2208
rect 27076 2144 27092 2208
rect 27156 2144 27172 2208
rect 27236 2144 27252 2208
rect 27316 2144 27324 2208
rect 27004 0 27324 2144
rect 31944 4928 32264 5952
rect 31944 4864 31952 4928
rect 32016 4864 32032 4928
rect 32096 4864 32112 4928
rect 32176 4864 32192 4928
rect 32256 4864 32264 4928
rect 31944 3840 32264 4864
rect 31944 3776 31952 3840
rect 32016 3776 32032 3840
rect 32096 3776 32112 3840
rect 32176 3776 32192 3840
rect 32256 3776 32264 3840
rect 31944 2752 32264 3776
rect 31944 2688 31952 2752
rect 32016 2688 32032 2752
rect 32096 2688 32112 2752
rect 32176 2688 32192 2752
rect 32256 2688 32264 2752
rect 31944 0 32264 2688
rect 33004 8736 33324 11250
rect 33004 8672 33012 8736
rect 33076 8672 33092 8736
rect 33156 8672 33172 8736
rect 33236 8672 33252 8736
rect 33316 8672 33324 8736
rect 33004 7648 33324 8672
rect 33004 7584 33012 7648
rect 33076 7584 33092 7648
rect 33156 7584 33172 7648
rect 33236 7584 33252 7648
rect 33316 7584 33324 7648
rect 33004 6560 33324 7584
rect 33004 6496 33012 6560
rect 33076 6496 33092 6560
rect 33156 6496 33172 6560
rect 33236 6496 33252 6560
rect 33316 6496 33324 6560
rect 33004 5472 33324 6496
rect 33004 5408 33012 5472
rect 33076 5408 33092 5472
rect 33156 5408 33172 5472
rect 33236 5408 33252 5472
rect 33316 5408 33324 5472
rect 33004 4384 33324 5408
rect 33004 4320 33012 4384
rect 33076 4320 33092 4384
rect 33156 4320 33172 4384
rect 33236 4320 33252 4384
rect 33316 4320 33324 4384
rect 33004 3296 33324 4320
rect 33004 3232 33012 3296
rect 33076 3232 33092 3296
rect 33156 3232 33172 3296
rect 33236 3232 33252 3296
rect 33316 3232 33324 3296
rect 33004 2208 33324 3232
rect 33004 2144 33012 2208
rect 33076 2144 33092 2208
rect 33156 2144 33172 2208
rect 33236 2144 33252 2208
rect 33316 2144 33324 2208
rect 33004 0 33324 2144
rect 37944 8192 38264 11250
rect 37944 8128 37952 8192
rect 38016 8128 38032 8192
rect 38096 8128 38112 8192
rect 38176 8128 38192 8192
rect 38256 8128 38264 8192
rect 37944 7104 38264 8128
rect 37944 7040 37952 7104
rect 38016 7040 38032 7104
rect 38096 7040 38112 7104
rect 38176 7040 38192 7104
rect 38256 7040 38264 7104
rect 37944 6016 38264 7040
rect 37944 5952 37952 6016
rect 38016 5952 38032 6016
rect 38096 5952 38112 6016
rect 38176 5952 38192 6016
rect 38256 5952 38264 6016
rect 37944 4928 38264 5952
rect 37944 4864 37952 4928
rect 38016 4864 38032 4928
rect 38096 4864 38112 4928
rect 38176 4864 38192 4928
rect 38256 4864 38264 4928
rect 37944 3840 38264 4864
rect 37944 3776 37952 3840
rect 38016 3776 38032 3840
rect 38096 3776 38112 3840
rect 38176 3776 38192 3840
rect 38256 3776 38264 3840
rect 37944 2752 38264 3776
rect 37944 2688 37952 2752
rect 38016 2688 38032 2752
rect 38096 2688 38112 2752
rect 38176 2688 38192 2752
rect 38256 2688 38264 2752
rect 37944 0 38264 2688
rect 39004 8736 39324 11250
rect 39004 8672 39012 8736
rect 39076 8672 39092 8736
rect 39156 8672 39172 8736
rect 39236 8672 39252 8736
rect 39316 8672 39324 8736
rect 39004 7648 39324 8672
rect 39004 7584 39012 7648
rect 39076 7584 39092 7648
rect 39156 7584 39172 7648
rect 39236 7584 39252 7648
rect 39316 7584 39324 7648
rect 39004 6560 39324 7584
rect 39004 6496 39012 6560
rect 39076 6496 39092 6560
rect 39156 6496 39172 6560
rect 39236 6496 39252 6560
rect 39316 6496 39324 6560
rect 39004 5472 39324 6496
rect 39004 5408 39012 5472
rect 39076 5408 39092 5472
rect 39156 5408 39172 5472
rect 39236 5408 39252 5472
rect 39316 5408 39324 5472
rect 39004 4384 39324 5408
rect 39004 4320 39012 4384
rect 39076 4320 39092 4384
rect 39156 4320 39172 4384
rect 39236 4320 39252 4384
rect 39316 4320 39324 4384
rect 39004 3296 39324 4320
rect 39004 3232 39012 3296
rect 39076 3232 39092 3296
rect 39156 3232 39172 3296
rect 39236 3232 39252 3296
rect 39316 3232 39324 3296
rect 39004 2208 39324 3232
rect 39004 2144 39012 2208
rect 39076 2144 39092 2208
rect 39156 2144 39172 2208
rect 39236 2144 39252 2208
rect 39316 2144 39324 2208
rect 39004 0 39324 2144
use sky130_fd_sc_hd__inv_2  _024_
timestamp -3599
transform 1 0 21436 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _025_
timestamp -3599
transform -1 0 14352 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _026_
timestamp -3599
transform 1 0 9108 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _027_
timestamp -3599
transform 1 0 19596 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__mux4_1  _028_
timestamp -3599
transform -1 0 24288 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__nand2b_1  _029_
timestamp -3599
transform -1 0 22908 0 -1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__o21ba_1  _030_
timestamp -3599
transform 1 0 23828 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _031_
timestamp -3599
transform -1 0 22356 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__a221o_1  _032_
timestamp -3599
transform 1 0 21804 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _033_
timestamp -3599
transform 1 0 22632 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__mux4_1  _034_
timestamp -3599
transform -1 0 12604 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__nand2b_1  _035_
timestamp -3599
transform -1 0 15640 0 1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__o21ba_1  _036_
timestamp -3599
transform 1 0 16192 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _037_
timestamp -3599
transform 1 0 14812 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__a221o_1  _038_
timestamp -3599
transform 1 0 14444 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _039_
timestamp -3599
transform -1 0 14904 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__mux4_1  _040_
timestamp -3599
transform 1 0 6348 0 -1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__nand2b_1  _041_
timestamp -3599
transform -1 0 10304 0 -1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__o21ba_1  _042_
timestamp -3599
transform 1 0 10764 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _043_
timestamp -3599
transform -1 0 9108 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__a221o_1  _044_
timestamp -3599
transform 1 0 9108 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _045_
timestamp -3599
transform -1 0 10304 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__mux4_1  _046_
timestamp -3599
transform -1 0 17848 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__nand2b_1  _047_
timestamp -3599
transform 1 0 21068 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__o21ba_1  _048_
timestamp -3599
transform 1 0 22356 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _049_
timestamp -3599
transform 1 0 20700 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__a221o_1  _050_
timestamp -3599
transform 1 0 17848 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _051_
timestamp -3599
transform -1 0 22356 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__dlxtp_1  _052_
timestamp -3599
transform 1 0 20516 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _053_
timestamp -3599
transform 1 0 20240 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _054_
timestamp -3599
transform -1 0 21620 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _055_
timestamp -3599
transform -1 0 14444 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _056_
timestamp -3599
transform -1 0 15180 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _057_
timestamp -3599
transform -1 0 17664 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _058_
timestamp -3599
transform 1 0 15456 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _059_
timestamp -3599
transform -1 0 17756 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _060_
timestamp -3599
transform -1 0 23552 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _061_
timestamp -3599
transform 1 0 21344 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _062_
timestamp -3599
transform 1 0 19504 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _063_
timestamp -3599
transform 1 0 19412 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_1  _065_
timestamp -3599
transform -1 0 38180 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _066_
timestamp -3599
transform 1 0 3128 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _067_
timestamp -3599
transform 1 0 38180 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _068_
timestamp -3599
transform -1 0 38732 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _069_
timestamp -3599
transform 1 0 37444 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _070_
timestamp -3599
transform 1 0 3496 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _071_
timestamp -3599
transform 1 0 2392 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _072_
timestamp -3599
transform 1 0 2760 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _073_
timestamp -3599
transform 1 0 2852 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _074_
timestamp -3599
transform 1 0 3220 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _075_
timestamp -3599
transform 1 0 2852 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _076_
timestamp -3599
transform 1 0 2852 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _077_
timestamp -3599
transform -1 0 38180 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _078_
timestamp -3599
transform 1 0 2760 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _079_
timestamp -3599
transform -1 0 38180 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _080_
timestamp -3599
transform -1 0 38180 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _081_
timestamp -3599
transform 1 0 4140 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _082_
timestamp -3599
transform 1 0 3128 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _083_
timestamp -3599
transform 1 0 2760 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _084_
timestamp -3599
transform -1 0 37720 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _085_
timestamp -3599
transform 1 0 13616 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _086_
timestamp -3599
transform 1 0 15272 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _087_
timestamp -3599
transform 1 0 20240 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _088_
timestamp -3599
transform 1 0 10028 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _089_
timestamp -3599
transform 1 0 9292 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _090_
timestamp -3599
transform 1 0 9660 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  _091_
timestamp -3599
transform 1 0 14076 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _092_
timestamp -3599
transform 1 0 13984 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _093_
timestamp -3599
transform 1 0 13156 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _094_
timestamp -3599
transform 1 0 13156 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  _095_
timestamp -3599
transform 1 0 19964 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _096_
timestamp -3599
transform 1 0 20332 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _097_
timestamp -3599
transform 1 0 19136 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _098_
timestamp -3599
transform -1 0 31004 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _099_
timestamp -3599
transform -1 0 31832 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _100_
timestamp -3599
transform -1 0 32108 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _101_
timestamp -3599
transform -1 0 32292 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _102_
timestamp -3599
transform -1 0 32936 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _103_
timestamp -3599
transform -1 0 32384 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _104_
timestamp -3599
transform -1 0 31464 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _105_
timestamp -3599
transform 1 0 35512 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _106_
timestamp -3599
transform -1 0 30728 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _107_
timestamp -3599
transform -1 0 31740 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _108_
timestamp -3599
transform -1 0 32660 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _109_
timestamp -3599
transform -1 0 33764 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _110_
timestamp -3599
transform -1 0 34500 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _111_
timestamp -3599
transform -1 0 35236 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _112_
timestamp -3599
transform -1 0 36156 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _113_
timestamp -3599
transform -1 0 36984 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _114_
timestamp -3599
transform -1 0 37720 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _115_
timestamp -3599
transform -1 0 38180 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _116_
timestamp -3599
transform 1 0 37904 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _117_
timestamp -3599
transform -1 0 28244 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _118_
timestamp -3599
transform -1 0 17388 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _119_
timestamp -3599
transform 1 0 11776 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _120_
timestamp -3599
transform -1 0 21988 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _121_
timestamp -3599
transform -1 0 3680 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _122_
timestamp -3599
transform -1 0 4048 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _123_
timestamp -3599
transform -1 0 4784 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _124_
timestamp -3599
transform -1 0 4140 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _125_
timestamp -3599
transform -1 0 25392 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _126_
timestamp -3599
transform -1 0 16192 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _127_
timestamp -3599
transform 1 0 9844 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _128_
timestamp -3599
transform -1 0 19596 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _129_
timestamp -3599
transform -1 0 27416 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _130_
timestamp -3599
transform -1 0 18032 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _131_
timestamp -3599
transform 1 0 8924 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _132_
timestamp -3599
transform 1 0 15916 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _133_
timestamp -3599
transform -1 0 24932 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _134_
timestamp -3599
transform 1 0 12788 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _135_
timestamp -3599
transform -1 0 7636 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _136_
timestamp -3599
transform -1 0 17112 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _137_
timestamp -3599
transform -1 0 30084 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _138_
timestamp -3599
transform -1 0 29808 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _139_
timestamp -3599
transform -1 0 29348 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _140_
timestamp -3599
transform -1 0 29072 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _141_
timestamp -3599
transform -1 0 28796 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _142_
timestamp -3599
transform -1 0 28520 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _143_
timestamp -3599
transform -1 0 27968 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _144_
timestamp -3599
transform -1 0 27692 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _145_
timestamp -3599
transform -1 0 26864 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _146_
timestamp -3599
transform 1 0 13708 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _147_
timestamp -3599
transform -1 0 7728 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _148_
timestamp -3599
transform 1 0 19136 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _149_
timestamp -3599
transform -1 0 24288 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _150_
timestamp -3599
transform 1 0 13524 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _151_
timestamp -3599
transform -1 0 6808 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _152_
timestamp -3599
transform 1 0 18492 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _153_
timestamp -3599
transform -1 0 32292 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _154_
timestamp -3599
transform -1 0 32936 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _155_
timestamp -3599
transform -1 0 32016 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _156_
timestamp -3599
transform -1 0 32660 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _157_
timestamp -3599
transform -1 0 32384 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _158_
timestamp -3599
transform -1 0 31832 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _159_
timestamp -3599
transform -1 0 31556 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _160_
timestamp -3599
transform -1 0 31280 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _161_
timestamp -3599
transform 1 0 24656 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _162_
timestamp -3599
transform -1 0 12328 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _163_
timestamp -3599
transform 1 0 3404 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _164_
timestamp -3599
transform 1 0 17480 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _165_
timestamp -3599
transform 1 0 24380 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _166_
timestamp -3599
transform -1 0 11868 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _167_
timestamp -3599
transform 1 0 3772 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _168_
timestamp -3599
transform -1 0 17112 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _169_
timestamp -3599
transform 1 0 29900 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1
timestamp -3599
transform -1 0 37904 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_2
timestamp -3599
transform -1 0 37904 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_3
timestamp -3599
transform 1 0 37720 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_4
timestamp -3599
transform -1 0 37904 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_5
timestamp -3599
transform 1 0 37260 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_6
timestamp -3599
transform -1 0 38916 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_7
timestamp -3599
transform -1 0 39100 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_8
timestamp -3599
transform 1 0 39008 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_9
timestamp -3599
transform 1 0 30544 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_10
timestamp -3599
transform -1 0 31280 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_11
timestamp -3599
transform -1 0 32016 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_12
timestamp -3599
transform -1 0 35512 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_13
timestamp -3599
transform -1 0 1748 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_14
timestamp -3599
transform -1 0 3864 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_15
timestamp -3599
transform -1 0 31556 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_16
timestamp -3599
transform -1 0 13616 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  fanout3
timestamp -3599
transform -1 0 26496 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3
timestamp -3599
transform 1 0 1380 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11
timestamp 1636964856
transform 1 0 2116 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23
timestamp -3599
transform 1 0 3220 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29
timestamp 1636964856
transform 1 0 3772 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_45
timestamp -3599
transform 1 0 5244 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_53
timestamp -3599
transform 1 0 5980 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_57
timestamp -3599
transform 1 0 6348 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62
timestamp 1636964856
transform 1 0 6808 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_74
timestamp -3599
transform 1 0 7912 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_82
timestamp -3599
transform 1 0 8648 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_85
timestamp -3599
transform 1 0 8924 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_91
timestamp -3599
transform 1 0 9476 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_102
timestamp -3599
transform 1 0 10488 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_110
timestamp -3599
transform 1 0 11224 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_113
timestamp 1636964856
transform 1 0 11500 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_125
timestamp 1636964856
transform 1 0 12604 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_137
timestamp -3599
transform 1 0 13708 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_141
timestamp 1636964856
transform 1 0 14076 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_153
timestamp 1636964856
transform 1 0 15180 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_165
timestamp -3599
transform 1 0 16284 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_169
timestamp 1636964856
transform 1 0 16652 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_181
timestamp 1636964856
transform 1 0 17756 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_193
timestamp -3599
transform 1 0 18860 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_197
timestamp 1636964856
transform 1 0 19228 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_209
timestamp 1636964856
transform 1 0 20332 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_221
timestamp -3599
transform 1 0 21436 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_225
timestamp 1636964856
transform 1 0 21804 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_237
timestamp 1636964856
transform 1 0 22908 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_249
timestamp -3599
transform 1 0 24012 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_253
timestamp 1636964856
transform 1 0 24380 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_265
timestamp 1636964856
transform 1 0 25484 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_277
timestamp -3599
transform 1 0 26588 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_281
timestamp 1636964856
transform 1 0 26956 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_293
timestamp 1636964856
transform 1 0 28060 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_305
timestamp -3599
transform 1 0 29164 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_309
timestamp 1636964856
transform 1 0 29532 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_321
timestamp 1636964856
transform 1 0 30636 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_333
timestamp -3599
transform 1 0 31740 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_337
timestamp 1636964856
transform 1 0 32108 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_349
timestamp 1636964856
transform 1 0 33212 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_361
timestamp -3599
transform 1 0 34316 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_365
timestamp 1636964856
transform 1 0 34684 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_377
timestamp 1636964856
transform 1 0 35788 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_389
timestamp -3599
transform 1 0 36892 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_393
timestamp -3599
transform 1 0 37260 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_3
timestamp 1636964856
transform 1 0 1380 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_15
timestamp 1636964856
transform 1 0 2484 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_27
timestamp 1636964856
transform 1 0 3588 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_39
timestamp 1636964856
transform 1 0 4692 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_51
timestamp -3599
transform 1 0 5796 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_55
timestamp -3599
transform 1 0 6164 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_57
timestamp 1636964856
transform 1 0 6348 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_69
timestamp 1636964856
transform 1 0 7452 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_81
timestamp 1636964856
transform 1 0 8556 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_93
timestamp 1636964856
transform 1 0 9660 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_105
timestamp -3599
transform 1 0 10764 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_111
timestamp -3599
transform 1 0 11316 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_113
timestamp 1636964856
transform 1 0 11500 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_125
timestamp 1636964856
transform 1 0 12604 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_137
timestamp 1636964856
transform 1 0 13708 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_149
timestamp 1636964856
transform 1 0 14812 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_161
timestamp -3599
transform 1 0 15916 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_167
timestamp -3599
transform 1 0 16468 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_169
timestamp 1636964856
transform 1 0 16652 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_181
timestamp 1636964856
transform 1 0 17756 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_193
timestamp 1636964856
transform 1 0 18860 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_205
timestamp 1636964856
transform 1 0 19964 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_217
timestamp -3599
transform 1 0 21068 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_1_225
timestamp -3599
transform 1 0 21804 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_231
timestamp -3599
transform 1 0 22356 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_237
timestamp 1636964856
transform 1 0 22908 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_249
timestamp 1636964856
transform 1 0 24012 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_261
timestamp 1636964856
transform 1 0 25116 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_273
timestamp -3599
transform 1 0 26220 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_279
timestamp -3599
transform 1 0 26772 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_281
timestamp 1636964856
transform 1 0 26956 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_293
timestamp 1636964856
transform 1 0 28060 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_305
timestamp 1636964856
transform 1 0 29164 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_317
timestamp 1636964856
transform 1 0 30268 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_329
timestamp -3599
transform 1 0 31372 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_335
timestamp -3599
transform 1 0 31924 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_337
timestamp 1636964856
transform 1 0 32108 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_349
timestamp 1636964856
transform 1 0 33212 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_361
timestamp 1636964856
transform 1 0 34316 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_373
timestamp 1636964856
transform 1 0 35420 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_385
timestamp -3599
transform 1 0 36524 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_391
timestamp -3599
transform 1 0 37076 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_393
timestamp 1636964856
transform 1 0 37260 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_1_405
timestamp -3599
transform 1 0 38364 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3
timestamp 1636964856
transform 1 0 1380 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_15
timestamp 1636964856
transform 1 0 2484 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_2_27
timestamp -3599
transform 1 0 3588 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_29
timestamp 1636964856
transform 1 0 3772 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_41
timestamp 1636964856
transform 1 0 4876 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_53
timestamp 1636964856
transform 1 0 5980 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_65
timestamp 1636964856
transform 1 0 7084 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_77
timestamp -3599
transform 1 0 8188 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_83
timestamp -3599
transform 1 0 8740 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_85
timestamp -3599
transform 1 0 8924 0 1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_2_90
timestamp 1636964856
transform 1 0 9384 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_2_102
timestamp -3599
transform 1 0 10488 0 1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_2_125
timestamp 1636964856
transform 1 0 12604 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_2_137
timestamp -3599
transform 1 0 13708 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_2_144
timestamp -3599
transform 1 0 14352 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_2_152
timestamp -3599
transform 1 0 15088 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_2_158
timestamp -3599
transform 1 0 15640 0 1 3264
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_2_182
timestamp 1636964856
transform 1 0 17848 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_2_194
timestamp -3599
transform 1 0 18952 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_2_197
timestamp -3599
transform 1 0 19228 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_2_204
timestamp -3599
transform 1 0 19872 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_2_212
timestamp -3599
transform 1 0 20608 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_253
timestamp 1636964856
transform 1 0 24380 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_265
timestamp -3599
transform 1 0 25484 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_271
timestamp -3599
transform 1 0 26036 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_276
timestamp 1636964856
transform 1 0 26496 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_288
timestamp 1636964856
transform 1 0 27600 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_2_300
timestamp -3599
transform 1 0 28704 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_2_309
timestamp -3599
transform 1 0 29532 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_2_317
timestamp -3599
transform 1 0 30268 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_322
timestamp -3599
transform 1 0 30728 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_326
timestamp -3599
transform 1 0 31096 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_330
timestamp 1636964856
transform 1 0 31464 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_342
timestamp 1636964856
transform 1 0 32568 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_2_354
timestamp -3599
transform 1 0 33672 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_2_362
timestamp -3599
transform 1 0 34408 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_2_365
timestamp -3599
transform 1 0 34684 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_371
timestamp -3599
transform 1 0 35236 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_377
timestamp 1636964856
transform 1 0 35788 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_389
timestamp -3599
transform 1 0 36892 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_413
timestamp -3599
transform 1 0 39100 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_3_3
timestamp -3599
transform 1 0 1380 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_3_11
timestamp -3599
transform 1 0 2116 0 -1 4352
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_3_30
timestamp 1636964856
transform 1 0 3864 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_42
timestamp 1636964856
transform 1 0 4968 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_3_54
timestamp -3599
transform 1 0 6072 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_3_87
timestamp -3599
transform 1 0 9108 0 -1 4352
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_3_100
timestamp 1636964856
transform 1 0 10304 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_113
timestamp 1636964856
transform 1 0 11500 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_125
timestamp 1636964856
transform 1 0 12604 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_137
timestamp 1636964856
transform 1 0 13708 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_3_158
timestamp -3599
transform 1 0 15640 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_3_166
timestamp -3599
transform 1 0 16376 0 -1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_3_169
timestamp 1636964856
transform 1 0 16652 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_3_181
timestamp -3599
transform 1 0 17756 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_190
timestamp 1636964856
transform 1 0 18584 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_202
timestamp -3599
transform 1 0 19688 0 -1 4352
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_3_211
timestamp 1636964856
transform 1 0 20516 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_3_223
timestamp -3599
transform 1 0 21620 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_225
timestamp 1636964856
transform 1 0 21804 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_3_237
timestamp -3599
transform 1 0 22908 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_3_245
timestamp -3599
transform 1 0 23644 0 -1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_3_255
timestamp 1636964856
transform 1 0 24564 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_267
timestamp 1636964856
transform 1 0 25668 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_3_279
timestamp -3599
transform 1 0 26772 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_281
timestamp 1636964856
transform 1 0 26956 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_293
timestamp 1636964856
transform 1 0 28060 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_305
timestamp 1636964856
transform 1 0 29164 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_3_317
timestamp -3599
transform 1 0 30268 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_3_325
timestamp -3599
transform 1 0 31004 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_3_333
timestamp -3599
transform 1 0 31740 0 -1 4352
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_3_337
timestamp 1636964856
transform 1 0 32108 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_349
timestamp 1636964856
transform 1 0 33212 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_361
timestamp 1636964856
transform 1 0 34316 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_373
timestamp 1636964856
transform 1 0 35420 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_385
timestamp -3599
transform 1 0 36524 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_391
timestamp -3599
transform 1 0 37076 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_393
timestamp 1636964856
transform 1 0 37260 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_3_405
timestamp -3599
transform 1 0 38364 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_409
timestamp -3599
transform 1 0 38732 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3
timestamp 1636964856
transform 1 0 1380 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_4_15
timestamp -3599
transform 1 0 2484 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_4_23
timestamp -3599
transform 1 0 3220 0 1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_4_29
timestamp 1636964856
transform 1 0 3772 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_41
timestamp 1636964856
transform 1 0 4876 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_53
timestamp 1636964856
transform 1 0 5980 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_65
timestamp 1636964856
transform 1 0 7084 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_77
timestamp -3599
transform 1 0 8188 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_83
timestamp -3599
transform 1 0 8740 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_85
timestamp 1636964856
transform 1 0 8924 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_4_97
timestamp -3599
transform 1 0 10028 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_4_113
timestamp -3599
transform 1 0 11500 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_4_122
timestamp -3599
transform 1 0 12328 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_4_130
timestamp -3599
transform 1 0 13064 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_4_138
timestamp -3599
transform 1 0 13800 0 1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_4_144
timestamp 1636964856
transform 1 0 14352 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_4_156
timestamp -3599
transform 1 0 15456 0 1 4352
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_4_172
timestamp 1636964856
transform 1 0 16928 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_184
timestamp 1636964856
transform 1 0 18032 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_197
timestamp 1636964856
transform 1 0 19228 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_209
timestamp 1636964856
transform 1 0 20332 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_4_221
timestamp -3599
transform 1 0 21436 0 1 4352
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_4_227
timestamp 1636964856
transform 1 0 21988 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_239
timestamp 1636964856
transform 1 0 23092 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_4_251
timestamp -3599
transform 1 0 24196 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_253
timestamp 1636964856
transform 1 0 24380 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_265
timestamp 1636964856
transform 1 0 25484 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_277
timestamp 1636964856
transform 1 0 26588 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_289
timestamp 1636964856
transform 1 0 27692 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_301
timestamp -3599
transform 1 0 28796 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_307
timestamp -3599
transform 1 0 29348 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_309
timestamp 1636964856
transform 1 0 29532 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_4_321
timestamp -3599
transform 1 0 30636 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_325
timestamp -3599
transform 1 0 31004 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_4_328
timestamp -3599
transform 1 0 31280 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_337
timestamp 1636964856
transform 1 0 32108 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_349
timestamp 1636964856
transform 1 0 33212 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_4_361
timestamp -3599
transform 1 0 34316 0 1 4352
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_4_365
timestamp 1636964856
transform 1 0 34684 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_377
timestamp 1636964856
transform 1 0 35788 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_4_389
timestamp -3599
transform 1 0 36892 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_4_397
timestamp -3599
transform 1 0 37628 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_4_403
timestamp -3599
transform 1 0 38180 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_409
timestamp -3599
transform 1 0 38732 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3
timestamp 1636964856
transform 1 0 1380 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_5_15
timestamp -3599
transform 1 0 2484 0 -1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_5_27
timestamp 1636964856
transform 1 0 3588 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_39
timestamp 1636964856
transform 1 0 4692 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_5_51
timestamp -3599
transform 1 0 5796 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_55
timestamp -3599
transform 1 0 6164 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_57
timestamp 1636964856
transform 1 0 6348 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_69
timestamp 1636964856
transform 1 0 7452 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_5_81
timestamp -3599
transform 1 0 8556 0 -1 5440
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_5_93
timestamp 1636964856
transform 1 0 9660 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_105
timestamp -3599
transform 1 0 10764 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_111
timestamp -3599
transform 1 0 11316 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_113
timestamp 1636964856
transform 1 0 11500 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_125
timestamp 1636964856
transform 1 0 12604 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_5_137
timestamp -3599
transform 1 0 13708 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_5_143
timestamp -3599
transform 1 0 14260 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_5_151
timestamp -3599
transform 1 0 14996 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_5_157
timestamp -3599
transform 1 0 15548 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_5_165
timestamp -3599
transform 1 0 16284 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_5_169
timestamp -3599
transform 1 0 16652 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_174
timestamp -3599
transform 1 0 17112 0 -1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_5_181
timestamp 1636964856
transform 1 0 17756 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_193
timestamp -3599
transform 1 0 18860 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_199
timestamp -3599
transform 1 0 19412 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_212
timestamp 1636964856
transform 1 0 20608 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_225
timestamp 1636964856
transform 1 0 21804 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_237
timestamp 1636964856
transform 1 0 22908 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_249
timestamp 1636964856
transform 1 0 24012 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_261
timestamp 1636964856
transform 1 0 25116 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_5_273
timestamp -3599
transform 1 0 26220 0 -1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_5_281
timestamp 1636964856
transform 1 0 26956 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_293
timestamp 1636964856
transform 1 0 28060 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_305
timestamp 1636964856
transform 1 0 29164 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_317
timestamp 1636964856
transform 1 0 30268 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_5_329
timestamp -3599
transform 1 0 31372 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_5_333
timestamp -3599
transform 1 0 31740 0 -1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_5_340
timestamp 1636964856
transform 1 0 32384 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_352
timestamp 1636964856
transform 1 0 33488 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_364
timestamp 1636964856
transform 1 0 34592 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_376
timestamp 1636964856
transform 1 0 35696 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_5_388
timestamp -3599
transform 1 0 36800 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_5_393
timestamp -3599
transform 1 0 37260 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_398
timestamp -3599
transform 1 0 37720 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_5_403
timestamp -3599
transform 1 0 38180 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_409
timestamp -3599
transform 1 0 38732 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3
timestamp 1636964856
transform 1 0 1380 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_6_15
timestamp -3599
transform 1 0 2484 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_23
timestamp -3599
transform 1 0 3220 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_27
timestamp -3599
transform 1 0 3588 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_32
timestamp 1636964856
transform 1 0 4048 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_44
timestamp 1636964856
transform 1 0 5152 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_6_56
timestamp -3599
transform 1 0 6256 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_6_62
timestamp -3599
transform 1 0 6808 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_68
timestamp -3599
transform 1 0 7360 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_72
timestamp 1636964856
transform 1 0 7728 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_6_88
timestamp -3599
transform 1 0 9200 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_92
timestamp -3599
transform 1 0 9568 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_101
timestamp 1636964856
transform 1 0 10396 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_113
timestamp 1636964856
transform 1 0 11500 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_125
timestamp -3599
transform 1 0 12604 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_6_134
timestamp -3599
transform 1 0 13432 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_6_139
timestamp -3599
transform 1 0 13892 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_6_141
timestamp -3599
transform 1 0 14076 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_6_150
timestamp -3599
transform 1 0 14904 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_6_158
timestamp -3599
transform 1 0 15640 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_6_164
timestamp -3599
transform 1 0 16192 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_170
timestamp -3599
transform 1 0 16744 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_177
timestamp 1636964856
transform 1 0 17388 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_6_192
timestamp -3599
transform 1 0 18768 0 1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_6_197
timestamp 1636964856
transform 1 0 19228 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_6_212
timestamp -3599
transform 1 0 20608 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_216
timestamp -3599
transform 1 0 20976 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_222
timestamp 1636964856
transform 1 0 21528 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_234
timestamp 1636964856
transform 1 0 22632 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_6_246
timestamp -3599
transform 1 0 23736 0 1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_6_259
timestamp 1636964856
transform 1 0 24932 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_271
timestamp 1636964856
transform 1 0 26036 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_283
timestamp 1636964856
transform 1 0 27140 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_295
timestamp 1636964856
transform 1 0 28244 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_6_307
timestamp -3599
transform 1 0 29348 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_309
timestamp 1636964856
transform 1 0 29532 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_321
timestamp 1636964856
transform 1 0 30636 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_6_333
timestamp -3599
transform 1 0 31740 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_339
timestamp 1636964856
transform 1 0 32292 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_351
timestamp 1636964856
transform 1 0 33396 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_6_363
timestamp -3599
transform 1 0 34500 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_365
timestamp 1636964856
transform 1 0 34684 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_6_377
timestamp -3599
transform 1 0 35788 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_6_381
timestamp -3599
transform 1 0 36156 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_6_390
timestamp -3599
transform 1 0 36984 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_6_403
timestamp -3599
transform 1 0 38180 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_409
timestamp -3599
transform 1 0 38732 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3
timestamp 1636964856
transform 1 0 1380 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_15
timestamp 1636964856
transform 1 0 2484 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_27
timestamp 1636964856
transform 1 0 3588 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_39
timestamp 1636964856
transform 1 0 4692 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_51
timestamp -3599
transform 1 0 5796 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_55
timestamp -3599
transform 1 0 6164 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_7_57
timestamp -3599
transform 1 0 6348 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_7_65
timestamp -3599
transform 1 0 7084 0 -1 6528
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_7_71
timestamp 1636964856
transform 1 0 7636 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_7_83
timestamp -3599
transform 1 0 8740 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_7_91
timestamp -3599
transform 1 0 9476 0 -1 6528
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_7_100
timestamp 1636964856
transform 1 0 10304 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_7_113
timestamp -3599
transform 1 0 11500 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_7_117
timestamp -3599
transform 1 0 11868 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_7_125
timestamp -3599
transform 1 0 12604 0 -1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_7_130
timestamp 1636964856
transform 1 0 13064 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_7_142
timestamp -3599
transform 1 0 14168 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_7_153
timestamp -3599
transform 1 0 15180 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_7_164
timestamp -3599
transform 1 0 16192 0 -1 6528
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_7_184
timestamp 1636964856
transform 1 0 18032 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_7_223
timestamp -3599
transform 1 0 21620 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_7_233
timestamp -3599
transform 1 0 22540 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_240
timestamp 1636964856
transform 1 0 23184 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_252
timestamp 1636964856
transform 1 0 24288 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_264
timestamp 1636964856
transform 1 0 25392 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_276
timestamp -3599
transform 1 0 26496 0 -1 6528
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_7_281
timestamp 1636964856
transform 1 0 26956 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_293
timestamp 1636964856
transform 1 0 28060 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_305
timestamp 1636964856
transform 1 0 29164 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_317
timestamp 1636964856
transform 1 0 30268 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_329
timestamp -3599
transform 1 0 31372 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_335
timestamp -3599
transform 1 0 31924 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_337
timestamp 1636964856
transform 1 0 32108 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_349
timestamp 1636964856
transform 1 0 33212 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_361
timestamp -3599
transform 1 0 34316 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_367
timestamp -3599
transform 1 0 34868 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_371
timestamp 1636964856
transform 1 0 35236 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_7_383
timestamp -3599
transform 1 0 36340 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_7_391
timestamp -3599
transform 1 0 37076 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_393
timestamp -3599
transform 1 0 37260 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_397
timestamp -3599
transform 1 0 37628 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_7_403
timestamp -3599
transform 1 0 38180 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_409
timestamp -3599
transform 1 0 38732 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3
timestamp 1636964856
transform 1 0 1380 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_8_15
timestamp -3599
transform 1 0 2484 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_22
timestamp -3599
transform 1 0 3128 0 1 6528
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_8_32
timestamp 1636964856
transform 1 0 4048 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_44
timestamp 1636964856
transform 1 0 5152 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_56
timestamp 1636964856
transform 1 0 6256 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_68
timestamp 1636964856
transform 1 0 7360 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_8_80
timestamp -3599
transform 1 0 8464 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_8_85
timestamp -3599
transform 1 0 8924 0 1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_8_98
timestamp 1636964856
transform 1 0 10120 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_110
timestamp -3599
transform 1 0 11224 0 1 6528
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_8_119
timestamp 1636964856
transform 1 0 12052 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_131
timestamp -3599
transform 1 0 13156 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_8_153
timestamp -3599
transform 1 0 15180 0 1 6528
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_8_180
timestamp 1636964856
transform 1 0 17664 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_8_192
timestamp -3599
transform 1 0 18768 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_8_197
timestamp -3599
transform 1 0 19228 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_8_244
timestamp -3599
transform 1 0 23552 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_8_253
timestamp -3599
transform 1 0 24380 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_8_259
timestamp -3599
transform 1 0 24932 0 1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_8_264
timestamp 1636964856
transform 1 0 25392 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_276
timestamp -3599
transform 1 0 26496 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_282
timestamp -3599
transform 1 0 27048 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_8_307
timestamp -3599
transform 1 0 29348 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_315
timestamp 1636964856
transform 1 0 30084 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_327
timestamp -3599
transform 1 0 31188 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_339
timestamp -3599
transform 1 0 32292 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_346
timestamp 1636964856
transform 1 0 32936 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_358
timestamp -3599
transform 1 0 34040 0 1 6528
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_8_365
timestamp 1636964856
transform 1 0 34684 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_377
timestamp 1636964856
transform 1 0 35788 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_8_389
timestamp -3599
transform 1 0 36892 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_8_397
timestamp -3599
transform 1 0 37628 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_8_403
timestamp -3599
transform 1 0 38180 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_9_12
timestamp -3599
transform 1 0 2208 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_9_26
timestamp -3599
transform 1 0 3496 0 -1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_9_40
timestamp 1636964856
transform 1 0 4784 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_9_52
timestamp -3599
transform 1 0 5888 0 -1 7616
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_9_57
timestamp 1636964856
transform 1 0 6348 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_69
timestamp 1636964856
transform 1 0 7452 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_81
timestamp 1636964856
transform 1 0 8556 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_93
timestamp 1636964856
transform 1 0 9660 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_105
timestamp -3599
transform 1 0 10764 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_111
timestamp -3599
transform 1 0 11316 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_113
timestamp 1636964856
transform 1 0 11500 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_9_125
timestamp -3599
transform 1 0 12604 0 -1 7616
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_9_145
timestamp 1636964856
transform 1 0 14444 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_9_157
timestamp -3599
transform 1 0 15548 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_9_165
timestamp -3599
transform 1 0 16284 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_169
timestamp 1636964856
transform 1 0 16652 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_181
timestamp 1636964856
transform 1 0 17756 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_193
timestamp -3599
transform 1 0 18860 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_199
timestamp 1636964856
transform 1 0 19412 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_9_223
timestamp -3599
transform 1 0 21620 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_239
timestamp 1636964856
transform 1 0 23092 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_251
timestamp 1636964856
transform 1 0 24196 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_263
timestamp 1636964856
transform 1 0 25300 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_9_275
timestamp -3599
transform 1 0 26404 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_279
timestamp -3599
transform 1 0 26772 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_281
timestamp 1636964856
transform 1 0 26956 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_293
timestamp 1636964856
transform 1 0 28060 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_305
timestamp 1636964856
transform 1 0 29164 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_9_317
timestamp -3599
transform 1 0 30268 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_9_334
timestamp -3599
transform 1 0 31832 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_9_346
timestamp -3599
transform 1 0 32936 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_9_355
timestamp -3599
transform 1 0 33764 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_359
timestamp -3599
transform 1 0 34132 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_363
timestamp 1636964856
transform 1 0 34500 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_375
timestamp 1636964856
transform 1 0 35604 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_9_387
timestamp -3599
transform 1 0 36708 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_391
timestamp -3599
transform 1 0 37076 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_10_15
timestamp -3599
transform 1 0 2484 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_10_23
timestamp -3599
transform 1 0 3220 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_29
timestamp -3599
transform 1 0 3772 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_37
timestamp -3599
transform 1 0 4508 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_41
timestamp -3599
transform 1 0 4876 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_10_46
timestamp -3599
transform 1 0 5336 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_10_58
timestamp -3599
transform 1 0 6440 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_64
timestamp -3599
transform 1 0 6992 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_10_70
timestamp -3599
transform 1 0 7544 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_10_82
timestamp -3599
transform 1 0 8648 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_10_89
timestamp -3599
transform 1 0 9292 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_10_94
timestamp -3599
transform 1 0 9752 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_10_106
timestamp -3599
transform 1 0 10856 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_110
timestamp -3599
transform 1 0 11224 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_115
timestamp -3599
transform 1 0 11684 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_121
timestamp -3599
transform 1 0 12236 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_125
timestamp -3599
transform 1 0 12604 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_130
timestamp -3599
transform 1 0 13064 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_134
timestamp -3599
transform 1 0 13432 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_10_139
timestamp -3599
transform 1 0 13892 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_10_141
timestamp -3599
transform 1 0 14076 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_10_148
timestamp -3599
transform 1 0 14720 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_10_154
timestamp -3599
transform 1 0 15272 0 1 7616
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_10_166
timestamp 1636964856
transform 1 0 16376 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_10_178
timestamp -3599
transform 1 0 17480 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_10_189
timestamp -3599
transform 1 0 18492 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_195
timestamp -3599
transform 1 0 19044 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_197
timestamp 1636964856
transform 1 0 19228 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_209
timestamp 1636964856
transform 1 0 20332 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_221
timestamp 1636964856
transform 1 0 21436 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_233
timestamp 1636964856
transform 1 0 22540 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_245
timestamp -3599
transform 1 0 23644 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_251
timestamp -3599
transform 1 0 24196 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_253
timestamp 1636964856
transform 1 0 24380 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_265
timestamp 1636964856
transform 1 0 25484 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_277
timestamp 1636964856
transform 1 0 26588 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_10_289
timestamp -3599
transform 1 0 27692 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_10_297
timestamp -3599
transform 1 0 28428 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_10_306
timestamp -3599
transform 1 0 29256 0 1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_10_312
timestamp 1636964856
transform 1 0 29808 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_324
timestamp 1636964856
transform 1 0 30912 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_336
timestamp 1636964856
transform 1 0 32016 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_348
timestamp 1636964856
transform 1 0 33120 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_10_360
timestamp -3599
transform 1 0 34224 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_10_369
timestamp -3599
transform 1 0 35052 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_10_379
timestamp -3599
transform 1 0 35972 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_385
timestamp -3599
transform 1 0 36524 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_10_391
timestamp -3599
transform 1 0 37076 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_10_403
timestamp -3599
transform 1 0 38180 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_11_18
timestamp -3599
transform 1 0 2760 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_11_29
timestamp -3599
transform 1 0 3772 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_57
timestamp -3599
transform 1 0 6348 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_85
timestamp -3599
transform 1 0 8924 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_11_113
timestamp -3599
transform 1 0 11500 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_11_141
timestamp -3599
transform 1 0 14076 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_11_169
timestamp -3599
transform 1 0 16652 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_175
timestamp -3599
transform 1 0 17204 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_185
timestamp -3599
transform 1 0 18124 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_11_197
timestamp -3599
transform 1 0 19228 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_207
timestamp 1636964856
transform 1 0 20148 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_11_222
timestamp -3599
transform 1 0 21528 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_11_271
timestamp -3599
transform 1 0 26036 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_11_279
timestamp -3599
transform 1 0 26772 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_11_281
timestamp -3599
transform 1 0 26956 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_11_289
timestamp -3599
transform 1 0 27692 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_11_307
timestamp -3599
transform 1 0 29348 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_322
timestamp 1636964856
transform 1 0 30728 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_11_334
timestamp -3599
transform 1 0 31832 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_337
timestamp -3599
transform 1 0 32108 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_362
timestamp -3599
transform 1 0 34408 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_11_389
timestamp -3599
transform 1 0 36892 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_409
timestamp -3599
transform 1 0 38732 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input1
timestamp -3599
transform 1 0 1932 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input2
timestamp -3599
transform 1 0 1380 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input3
timestamp -3599
transform 1 0 1656 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input4
timestamp -3599
transform 1 0 1380 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input5
timestamp -3599
transform 1 0 1380 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input6
timestamp -3599
transform -1 0 2208 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input7
timestamp -3599
transform -1 0 2760 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input8
timestamp -3599
transform -1 0 1932 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input9
timestamp -3599
transform 1 0 2208 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input10
timestamp -3599
transform 1 0 1656 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input11
timestamp -3599
transform 1 0 1932 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input12
timestamp -3599
transform 1 0 2208 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input13
timestamp -3599
transform 1 0 9568 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__buf_1  input14
timestamp -3599
transform 1 0 17940 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input15
timestamp -3599
transform -1 0 18492 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input16
timestamp -3599
transform -1 0 18584 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input17
timestamp -3599
transform 1 0 18584 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input18
timestamp -3599
transform -1 0 21528 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input19
timestamp -3599
transform -1 0 22080 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input20
timestamp -3599
transform -1 0 22356 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input21
timestamp -3599
transform -1 0 22632 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input22
timestamp -3599
transform -1 0 22908 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input23
timestamp -3599
transform -1 0 23184 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input24
timestamp -3599
transform -1 0 23460 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input25
timestamp -3599
transform 1 0 23460 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input26
timestamp -3599
transform -1 0 19136 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input27
timestamp -3599
transform -1 0 19596 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input28
timestamp -3599
transform -1 0 19872 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input29
timestamp -3599
transform 1 0 19872 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input30
timestamp -3599
transform -1 0 24012 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input31
timestamp -3599
transform -1 0 24288 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input32
timestamp -3599
transform -1 0 24656 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input33
timestamp -3599
transform 1 0 24656 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input34
timestamp -3599
transform -1 0 25208 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input35
timestamp -3599
transform -1 0 25484 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input36
timestamp -3599
transform -1 0 25760 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input37
timestamp -3599
transform 1 0 25760 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input38
timestamp -3599
transform -1 0 28152 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input39
timestamp -3599
transform 1 0 28152 0 -1 8704
box -38 -48 958 592
use sky130_fd_sc_hd__buf_1  input40
timestamp -3599
transform -1 0 29348 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input41
timestamp -3599
transform -1 0 28980 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input42
timestamp -3599
transform -1 0 29256 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input43
timestamp -3599
transform 1 0 29532 0 -1 8704
box -38 -48 958 592
use sky130_fd_sc_hd__buf_1  input44
timestamp -3599
transform -1 0 29808 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input45
timestamp -3599
transform -1 0 30728 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output46
timestamp -3599
transform 1 0 38456 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output47
timestamp -3599
transform 1 0 39192 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output48
timestamp -3599
transform 1 0 38824 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output49
timestamp -3599
transform 1 0 39192 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output50
timestamp -3599
transform 1 0 38824 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output51
timestamp -3599
transform 1 0 39192 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output52
timestamp -3599
transform 1 0 38824 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output53
timestamp -3599
transform 1 0 39192 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output54
timestamp -3599
transform 1 0 38824 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output55
timestamp -3599
transform 1 0 38456 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output56
timestamp -3599
transform 1 0 39192 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output57
timestamp -3599
transform 1 0 38088 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output58
timestamp -3599
transform 1 0 37720 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output59
timestamp -3599
transform 1 0 39192 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output60
timestamp -3599
transform 1 0 38824 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output61
timestamp -3599
transform 1 0 39192 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output62
timestamp -3599
transform 1 0 39192 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output63
timestamp -3599
transform 1 0 38824 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output64
timestamp -3599
transform 1 0 38456 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output65
timestamp -3599
transform 1 0 39192 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output66
timestamp -3599
transform 1 0 39192 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output67
timestamp -3599
transform 1 0 38456 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output68
timestamp -3599
transform -1 0 38088 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output69
timestamp -3599
transform 1 0 38824 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output70
timestamp -3599
transform 1 0 38088 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output71
timestamp -3599
transform 1 0 38824 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output72
timestamp -3599
transform 1 0 37352 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output73
timestamp -3599
transform 1 0 38456 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output74
timestamp -3599
transform 1 0 39192 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output75
timestamp -3599
transform 1 0 38824 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output76
timestamp -3599
transform 1 0 39192 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output77
timestamp -3599
transform 1 0 38824 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output78
timestamp -3599
transform 1 0 32568 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output79
timestamp -3599
transform 1 0 36156 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output80
timestamp -3599
transform 1 0 35604 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output81
timestamp -3599
transform 1 0 36524 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output82
timestamp -3599
transform 1 0 36156 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output83
timestamp -3599
transform 1 0 37260 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output84
timestamp -3599
transform 1 0 36708 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output85
timestamp -3599
transform 1 0 37628 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output86
timestamp -3599
transform 1 0 37996 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output87
timestamp -3599
transform 1 0 38364 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output88
timestamp -3599
transform -1 0 38180 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output89
timestamp -3599
transform 1 0 32936 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output90
timestamp -3599
transform 1 0 33304 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output91
timestamp -3599
transform 1 0 33672 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output92
timestamp -3599
transform 1 0 34040 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output93
timestamp -3599
transform 1 0 34684 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output94
timestamp -3599
transform 1 0 35052 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output95
timestamp -3599
transform 1 0 34684 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output96
timestamp -3599
transform -1 0 35788 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output97
timestamp -3599
transform 1 0 35788 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output98
timestamp -3599
transform -1 0 2116 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output99
timestamp -3599
transform -1 0 3680 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output100
timestamp -3599
transform -1 0 5244 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output101
timestamp -3599
transform -1 0 6808 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output102
timestamp -3599
transform -1 0 3680 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output103
timestamp -3599
transform -1 0 3312 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output104
timestamp -3599
transform -1 0 3680 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output105
timestamp -3599
transform -1 0 4508 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output106
timestamp -3599
transform 1 0 4048 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output107
timestamp -3599
transform 1 0 4416 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output108
timestamp -3599
transform 1 0 4968 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output109
timestamp -3599
transform 1 0 4784 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output110
timestamp -3599
transform -1 0 5520 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output111
timestamp -3599
transform -1 0 5888 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output112
timestamp -3599
transform -1 0 6440 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output113
timestamp -3599
transform -1 0 6256 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output114
timestamp -3599
transform -1 0 6992 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output115
timestamp -3599
transform -1 0 6992 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output116
timestamp -3599
transform -1 0 7544 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output117
timestamp -3599
transform -1 0 7360 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output118
timestamp -3599
transform -1 0 7728 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output119
timestamp -3599
transform -1 0 8096 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output120
timestamp -3599
transform 1 0 8280 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output121
timestamp -3599
transform -1 0 8464 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output122
timestamp -3599
transform -1 0 9292 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output123
timestamp -3599
transform 1 0 11040 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output124
timestamp -3599
transform -1 0 12236 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output125
timestamp -3599
transform -1 0 11960 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output126
timestamp -3599
transform -1 0 12328 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output127
timestamp -3599
transform 1 0 12696 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output128
timestamp -3599
transform -1 0 12696 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output129
timestamp -3599
transform -1 0 8832 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output130
timestamp -3599
transform -1 0 9752 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output131
timestamp -3599
transform -1 0 9568 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output132
timestamp -3599
transform -1 0 9936 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output133
timestamp -3599
transform -1 0 10304 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output134
timestamp -3599
transform -1 0 10856 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output135
timestamp -3599
transform -1 0 10672 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output136
timestamp -3599
transform -1 0 11040 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output137
timestamp -3599
transform -1 0 11684 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output138
timestamp -3599
transform -1 0 13064 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output139
timestamp -3599
transform 1 0 16008 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output140
timestamp -3599
transform -1 0 16192 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output141
timestamp -3599
transform -1 0 16560 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output142
timestamp -3599
transform 1 0 16836 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output143
timestamp -3599
transform 1 0 17756 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output144
timestamp -3599
transform 1 0 17388 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output145
timestamp -3599
transform -1 0 13892 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output146
timestamp -3599
transform -1 0 13432 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output147
timestamp -3599
transform 1 0 13616 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output148
timestamp -3599
transform -1 0 14720 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output149
timestamp -3599
transform -1 0 14720 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output150
timestamp -3599
transform -1 0 15272 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output151
timestamp -3599
transform -1 0 15088 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output152
timestamp -3599
transform -1 0 15456 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output153
timestamp -3599
transform 1 0 15456 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  output154
timestamp -3599
transform -1 0 32568 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Left_12
timestamp -3599
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Right_0
timestamp -3599
transform -1 0 39836 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Left_13
timestamp -3599
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Right_1
timestamp -3599
transform -1 0 39836 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Left_14
timestamp -3599
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Right_2
timestamp -3599
transform -1 0 39836 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Left_15
timestamp -3599
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Right_3
timestamp -3599
transform -1 0 39836 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Left_16
timestamp -3599
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Right_4
timestamp -3599
transform -1 0 39836 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Left_17
timestamp -3599
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Right_5
timestamp -3599
transform -1 0 39836 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Left_18
timestamp -3599
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Right_6
timestamp -3599
transform -1 0 39836 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Left_19
timestamp -3599
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Right_7
timestamp -3599
transform -1 0 39836 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Left_20
timestamp -3599
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Right_8
timestamp -3599
transform -1 0 39836 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Left_21
timestamp -3599
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Right_9
timestamp -3599
transform -1 0 39836 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_Left_22
timestamp -3599
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_Right_10
timestamp -3599
transform -1 0 39836 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_Left_23
timestamp -3599
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_Right_11
timestamp -3599
transform -1 0 39836 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  S_CPU_IRQ_155
timestamp -3599
transform -1 0 17940 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_24
timestamp -3599
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_25
timestamp -3599
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_26
timestamp -3599
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_27
timestamp -3599
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_28
timestamp -3599
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_29
timestamp -3599
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_30
timestamp -3599
transform 1 0 19136 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_31
timestamp -3599
transform 1 0 21712 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_32
timestamp -3599
transform 1 0 24288 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_33
timestamp -3599
transform 1 0 26864 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_34
timestamp -3599
transform 1 0 29440 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_35
timestamp -3599
transform 1 0 32016 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_36
timestamp -3599
transform 1 0 34592 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_37
timestamp -3599
transform 1 0 37168 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_38
timestamp -3599
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_39
timestamp -3599
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_40
timestamp -3599
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_41
timestamp -3599
transform 1 0 21712 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_42
timestamp -3599
transform 1 0 26864 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_43
timestamp -3599
transform 1 0 32016 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_44
timestamp -3599
transform 1 0 37168 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_45
timestamp -3599
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_46
timestamp -3599
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_47
timestamp -3599
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_48
timestamp -3599
transform 1 0 19136 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_49
timestamp -3599
transform 1 0 24288 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_50
timestamp -3599
transform 1 0 29440 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_51
timestamp -3599
transform 1 0 34592 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_52
timestamp -3599
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_53
timestamp -3599
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_54
timestamp -3599
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_55
timestamp -3599
transform 1 0 21712 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_56
timestamp -3599
transform 1 0 26864 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_57
timestamp -3599
transform 1 0 32016 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_58
timestamp -3599
transform 1 0 37168 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_59
timestamp -3599
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_60
timestamp -3599
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_61
timestamp -3599
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_62
timestamp -3599
transform 1 0 19136 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_63
timestamp -3599
transform 1 0 24288 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_64
timestamp -3599
transform 1 0 29440 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_65
timestamp -3599
transform 1 0 34592 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_66
timestamp -3599
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_67
timestamp -3599
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_68
timestamp -3599
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_69
timestamp -3599
transform 1 0 21712 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_70
timestamp -3599
transform 1 0 26864 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_71
timestamp -3599
transform 1 0 32016 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_72
timestamp -3599
transform 1 0 37168 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_73
timestamp -3599
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_74
timestamp -3599
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_75
timestamp -3599
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_76
timestamp -3599
transform 1 0 19136 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_77
timestamp -3599
transform 1 0 24288 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_78
timestamp -3599
transform 1 0 29440 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_79
timestamp -3599
transform 1 0 34592 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_80
timestamp -3599
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_81
timestamp -3599
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_82
timestamp -3599
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_83
timestamp -3599
transform 1 0 21712 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_84
timestamp -3599
transform 1 0 26864 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_85
timestamp -3599
transform 1 0 32016 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_86
timestamp -3599
transform 1 0 37168 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_87
timestamp -3599
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_88
timestamp -3599
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_89
timestamp -3599
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_90
timestamp -3599
transform 1 0 19136 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_91
timestamp -3599
transform 1 0 24288 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_92
timestamp -3599
transform 1 0 29440 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_93
timestamp -3599
transform 1 0 34592 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_94
timestamp -3599
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_95
timestamp -3599
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_96
timestamp -3599
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_97
timestamp -3599
transform 1 0 21712 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_98
timestamp -3599
transform 1 0 26864 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_99
timestamp -3599
transform 1 0 32016 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_100
timestamp -3599
transform 1 0 37168 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_101
timestamp -3599
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_102
timestamp -3599
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_103
timestamp -3599
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_104
timestamp -3599
transform 1 0 19136 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_105
timestamp -3599
transform 1 0 24288 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_106
timestamp -3599
transform 1 0 29440 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_107
timestamp -3599
transform 1 0 34592 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_108
timestamp -3599
transform 1 0 3680 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_109
timestamp -3599
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_110
timestamp -3599
transform 1 0 8832 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_111
timestamp -3599
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_112
timestamp -3599
transform 1 0 13984 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_113
timestamp -3599
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_114
timestamp -3599
transform 1 0 19136 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_115
timestamp -3599
transform 1 0 21712 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_116
timestamp -3599
transform 1 0 24288 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_117
timestamp -3599
transform 1 0 26864 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_118
timestamp -3599
transform 1 0 29440 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_119
timestamp -3599
transform 1 0 32016 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_120
timestamp -3599
transform 1 0 34592 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_121
timestamp -3599
transform 1 0 37168 0 -1 8704
box -38 -48 130 592
<< labels >>
flabel metal2 s 17590 11194 17646 11250 0 FreeSans 224 0 0 0 Co
port 0 nsew signal output
flabel metal3 s 0 1368 120 1488 0 FreeSans 480 0 0 0 FrameData[0]
port 1 nsew signal input
flabel metal3 s 0 4088 120 4208 0 FreeSans 480 0 0 0 FrameData[10]
port 2 nsew signal input
flabel metal3 s 0 4360 120 4480 0 FreeSans 480 0 0 0 FrameData[11]
port 3 nsew signal input
flabel metal3 s 0 4632 120 4752 0 FreeSans 480 0 0 0 FrameData[12]
port 4 nsew signal input
flabel metal3 s 0 4904 120 5024 0 FreeSans 480 0 0 0 FrameData[13]
port 5 nsew signal input
flabel metal3 s 0 5176 120 5296 0 FreeSans 480 0 0 0 FrameData[14]
port 6 nsew signal input
flabel metal3 s 0 5448 120 5568 0 FreeSans 480 0 0 0 FrameData[15]
port 7 nsew signal input
flabel metal3 s 0 5720 120 5840 0 FreeSans 480 0 0 0 FrameData[16]
port 8 nsew signal input
flabel metal3 s 0 5992 120 6112 0 FreeSans 480 0 0 0 FrameData[17]
port 9 nsew signal input
flabel metal3 s 0 6264 120 6384 0 FreeSans 480 0 0 0 FrameData[18]
port 10 nsew signal input
flabel metal3 s 0 6536 120 6656 0 FreeSans 480 0 0 0 FrameData[19]
port 11 nsew signal input
flabel metal3 s 0 1640 120 1760 0 FreeSans 480 0 0 0 FrameData[1]
port 12 nsew signal input
flabel metal3 s 0 6808 120 6928 0 FreeSans 480 0 0 0 FrameData[20]
port 13 nsew signal input
flabel metal3 s 0 7080 120 7200 0 FreeSans 480 0 0 0 FrameData[21]
port 14 nsew signal input
flabel metal3 s 0 7352 120 7472 0 FreeSans 480 0 0 0 FrameData[22]
port 15 nsew signal input
flabel metal3 s 0 7624 120 7744 0 FreeSans 480 0 0 0 FrameData[23]
port 16 nsew signal input
flabel metal3 s 0 7896 120 8016 0 FreeSans 480 0 0 0 FrameData[24]
port 17 nsew signal input
flabel metal3 s 0 8168 120 8288 0 FreeSans 480 0 0 0 FrameData[25]
port 18 nsew signal input
flabel metal3 s 0 8440 120 8560 0 FreeSans 480 0 0 0 FrameData[26]
port 19 nsew signal input
flabel metal3 s 0 8712 120 8832 0 FreeSans 480 0 0 0 FrameData[27]
port 20 nsew signal input
flabel metal3 s 0 8984 120 9104 0 FreeSans 480 0 0 0 FrameData[28]
port 21 nsew signal input
flabel metal3 s 0 9256 120 9376 0 FreeSans 480 0 0 0 FrameData[29]
port 22 nsew signal input
flabel metal3 s 0 1912 120 2032 0 FreeSans 480 0 0 0 FrameData[2]
port 23 nsew signal input
flabel metal3 s 0 9528 120 9648 0 FreeSans 480 0 0 0 FrameData[30]
port 24 nsew signal input
flabel metal3 s 0 9800 120 9920 0 FreeSans 480 0 0 0 FrameData[31]
port 25 nsew signal input
flabel metal3 s 0 2184 120 2304 0 FreeSans 480 0 0 0 FrameData[3]
port 26 nsew signal input
flabel metal3 s 0 2456 120 2576 0 FreeSans 480 0 0 0 FrameData[4]
port 27 nsew signal input
flabel metal3 s 0 2728 120 2848 0 FreeSans 480 0 0 0 FrameData[5]
port 28 nsew signal input
flabel metal3 s 0 3000 120 3120 0 FreeSans 480 0 0 0 FrameData[6]
port 29 nsew signal input
flabel metal3 s 0 3272 120 3392 0 FreeSans 480 0 0 0 FrameData[7]
port 30 nsew signal input
flabel metal3 s 0 3544 120 3664 0 FreeSans 480 0 0 0 FrameData[8]
port 31 nsew signal input
flabel metal3 s 0 3816 120 3936 0 FreeSans 480 0 0 0 FrameData[9]
port 32 nsew signal input
flabel metal3 s 40880 1368 41000 1488 0 FreeSans 480 0 0 0 FrameData_O[0]
port 33 nsew signal output
flabel metal3 s 40880 4088 41000 4208 0 FreeSans 480 0 0 0 FrameData_O[10]
port 34 nsew signal output
flabel metal3 s 40880 4360 41000 4480 0 FreeSans 480 0 0 0 FrameData_O[11]
port 35 nsew signal output
flabel metal3 s 40880 4632 41000 4752 0 FreeSans 480 0 0 0 FrameData_O[12]
port 36 nsew signal output
flabel metal3 s 40880 4904 41000 5024 0 FreeSans 480 0 0 0 FrameData_O[13]
port 37 nsew signal output
flabel metal3 s 40880 5176 41000 5296 0 FreeSans 480 0 0 0 FrameData_O[14]
port 38 nsew signal output
flabel metal3 s 40880 5448 41000 5568 0 FreeSans 480 0 0 0 FrameData_O[15]
port 39 nsew signal output
flabel metal3 s 40880 5720 41000 5840 0 FreeSans 480 0 0 0 FrameData_O[16]
port 40 nsew signal output
flabel metal3 s 40880 5992 41000 6112 0 FreeSans 480 0 0 0 FrameData_O[17]
port 41 nsew signal output
flabel metal3 s 40880 6264 41000 6384 0 FreeSans 480 0 0 0 FrameData_O[18]
port 42 nsew signal output
flabel metal3 s 40880 6536 41000 6656 0 FreeSans 480 0 0 0 FrameData_O[19]
port 43 nsew signal output
flabel metal3 s 40880 1640 41000 1760 0 FreeSans 480 0 0 0 FrameData_O[1]
port 44 nsew signal output
flabel metal3 s 40880 6808 41000 6928 0 FreeSans 480 0 0 0 FrameData_O[20]
port 45 nsew signal output
flabel metal3 s 40880 7080 41000 7200 0 FreeSans 480 0 0 0 FrameData_O[21]
port 46 nsew signal output
flabel metal3 s 40880 7352 41000 7472 0 FreeSans 480 0 0 0 FrameData_O[22]
port 47 nsew signal output
flabel metal3 s 40880 7624 41000 7744 0 FreeSans 480 0 0 0 FrameData_O[23]
port 48 nsew signal output
flabel metal3 s 40880 7896 41000 8016 0 FreeSans 480 0 0 0 FrameData_O[24]
port 49 nsew signal output
flabel metal3 s 40880 8168 41000 8288 0 FreeSans 480 0 0 0 FrameData_O[25]
port 50 nsew signal output
flabel metal3 s 40880 8440 41000 8560 0 FreeSans 480 0 0 0 FrameData_O[26]
port 51 nsew signal output
flabel metal3 s 40880 8712 41000 8832 0 FreeSans 480 0 0 0 FrameData_O[27]
port 52 nsew signal output
flabel metal3 s 40880 8984 41000 9104 0 FreeSans 480 0 0 0 FrameData_O[28]
port 53 nsew signal output
flabel metal3 s 40880 9256 41000 9376 0 FreeSans 480 0 0 0 FrameData_O[29]
port 54 nsew signal output
flabel metal3 s 40880 1912 41000 2032 0 FreeSans 480 0 0 0 FrameData_O[2]
port 55 nsew signal output
flabel metal3 s 40880 9528 41000 9648 0 FreeSans 480 0 0 0 FrameData_O[30]
port 56 nsew signal output
flabel metal3 s 40880 9800 41000 9920 0 FreeSans 480 0 0 0 FrameData_O[31]
port 57 nsew signal output
flabel metal3 s 40880 2184 41000 2304 0 FreeSans 480 0 0 0 FrameData_O[3]
port 58 nsew signal output
flabel metal3 s 40880 2456 41000 2576 0 FreeSans 480 0 0 0 FrameData_O[4]
port 59 nsew signal output
flabel metal3 s 40880 2728 41000 2848 0 FreeSans 480 0 0 0 FrameData_O[5]
port 60 nsew signal output
flabel metal3 s 40880 3000 41000 3120 0 FreeSans 480 0 0 0 FrameData_O[6]
port 61 nsew signal output
flabel metal3 s 40880 3272 41000 3392 0 FreeSans 480 0 0 0 FrameData_O[7]
port 62 nsew signal output
flabel metal3 s 40880 3544 41000 3664 0 FreeSans 480 0 0 0 FrameData_O[8]
port 63 nsew signal output
flabel metal3 s 40880 3816 41000 3936 0 FreeSans 480 0 0 0 FrameData_O[9]
port 64 nsew signal output
flabel metal2 s 9494 0 9550 56 0 FreeSans 224 0 0 0 FrameStrobe[0]
port 65 nsew signal input
flabel metal2 s 25134 0 25190 56 0 FreeSans 224 0 0 0 FrameStrobe[10]
port 66 nsew signal input
flabel metal2 s 26698 0 26754 56 0 FreeSans 224 0 0 0 FrameStrobe[11]
port 67 nsew signal input
flabel metal2 s 28262 0 28318 56 0 FreeSans 224 0 0 0 FrameStrobe[12]
port 68 nsew signal input
flabel metal2 s 29826 0 29882 56 0 FreeSans 224 0 0 0 FrameStrobe[13]
port 69 nsew signal input
flabel metal2 s 31390 0 31446 56 0 FreeSans 224 0 0 0 FrameStrobe[14]
port 70 nsew signal input
flabel metal2 s 32954 0 33010 56 0 FreeSans 224 0 0 0 FrameStrobe[15]
port 71 nsew signal input
flabel metal2 s 34518 0 34574 56 0 FreeSans 224 0 0 0 FrameStrobe[16]
port 72 nsew signal input
flabel metal2 s 36082 0 36138 56 0 FreeSans 224 0 0 0 FrameStrobe[17]
port 73 nsew signal input
flabel metal2 s 37646 0 37702 56 0 FreeSans 224 0 0 0 FrameStrobe[18]
port 74 nsew signal input
flabel metal2 s 39210 0 39266 56 0 FreeSans 224 0 0 0 FrameStrobe[19]
port 75 nsew signal input
flabel metal2 s 11058 0 11114 56 0 FreeSans 224 0 0 0 FrameStrobe[1]
port 76 nsew signal input
flabel metal2 s 12622 0 12678 56 0 FreeSans 224 0 0 0 FrameStrobe[2]
port 77 nsew signal input
flabel metal2 s 14186 0 14242 56 0 FreeSans 224 0 0 0 FrameStrobe[3]
port 78 nsew signal input
flabel metal2 s 15750 0 15806 56 0 FreeSans 224 0 0 0 FrameStrobe[4]
port 79 nsew signal input
flabel metal2 s 17314 0 17370 56 0 FreeSans 224 0 0 0 FrameStrobe[5]
port 80 nsew signal input
flabel metal2 s 18878 0 18934 56 0 FreeSans 224 0 0 0 FrameStrobe[6]
port 81 nsew signal input
flabel metal2 s 20442 0 20498 56 0 FreeSans 224 0 0 0 FrameStrobe[7]
port 82 nsew signal input
flabel metal2 s 22006 0 22062 56 0 FreeSans 224 0 0 0 FrameStrobe[8]
port 83 nsew signal input
flabel metal2 s 23570 0 23626 56 0 FreeSans 224 0 0 0 FrameStrobe[9]
port 84 nsew signal input
flabel metal2 s 32494 11194 32550 11250 0 FreeSans 224 0 0 0 FrameStrobe_O[0]
port 85 nsew signal output
flabel metal2 s 35254 11194 35310 11250 0 FreeSans 224 0 0 0 FrameStrobe_O[10]
port 86 nsew signal output
flabel metal2 s 35530 11194 35586 11250 0 FreeSans 224 0 0 0 FrameStrobe_O[11]
port 87 nsew signal output
flabel metal2 s 35806 11194 35862 11250 0 FreeSans 224 0 0 0 FrameStrobe_O[12]
port 88 nsew signal output
flabel metal2 s 36082 11194 36138 11250 0 FreeSans 224 0 0 0 FrameStrobe_O[13]
port 89 nsew signal output
flabel metal2 s 36358 11194 36414 11250 0 FreeSans 224 0 0 0 FrameStrobe_O[14]
port 90 nsew signal output
flabel metal2 s 36634 11194 36690 11250 0 FreeSans 224 0 0 0 FrameStrobe_O[15]
port 91 nsew signal output
flabel metal2 s 36910 11194 36966 11250 0 FreeSans 224 0 0 0 FrameStrobe_O[16]
port 92 nsew signal output
flabel metal2 s 37186 11194 37242 11250 0 FreeSans 224 0 0 0 FrameStrobe_O[17]
port 93 nsew signal output
flabel metal2 s 37462 11194 37518 11250 0 FreeSans 224 0 0 0 FrameStrobe_O[18]
port 94 nsew signal output
flabel metal2 s 37738 11194 37794 11250 0 FreeSans 224 0 0 0 FrameStrobe_O[19]
port 95 nsew signal output
flabel metal2 s 32770 11194 32826 11250 0 FreeSans 224 0 0 0 FrameStrobe_O[1]
port 96 nsew signal output
flabel metal2 s 33046 11194 33102 11250 0 FreeSans 224 0 0 0 FrameStrobe_O[2]
port 97 nsew signal output
flabel metal2 s 33322 11194 33378 11250 0 FreeSans 224 0 0 0 FrameStrobe_O[3]
port 98 nsew signal output
flabel metal2 s 33598 11194 33654 11250 0 FreeSans 224 0 0 0 FrameStrobe_O[4]
port 99 nsew signal output
flabel metal2 s 33874 11194 33930 11250 0 FreeSans 224 0 0 0 FrameStrobe_O[5]
port 100 nsew signal output
flabel metal2 s 34150 11194 34206 11250 0 FreeSans 224 0 0 0 FrameStrobe_O[6]
port 101 nsew signal output
flabel metal2 s 34426 11194 34482 11250 0 FreeSans 224 0 0 0 FrameStrobe_O[7]
port 102 nsew signal output
flabel metal2 s 34702 11194 34758 11250 0 FreeSans 224 0 0 0 FrameStrobe_O[8]
port 103 nsew signal output
flabel metal2 s 34978 11194 35034 11250 0 FreeSans 224 0 0 0 FrameStrobe_O[9]
port 104 nsew signal output
flabel metal2 s 1674 0 1730 56 0 FreeSans 224 0 0 0 IRQ_top0
port 105 nsew signal output
flabel metal2 s 3238 0 3294 56 0 FreeSans 224 0 0 0 IRQ_top1
port 106 nsew signal output
flabel metal2 s 4802 0 4858 56 0 FreeSans 224 0 0 0 IRQ_top2
port 107 nsew signal output
flabel metal2 s 6366 0 6422 56 0 FreeSans 224 0 0 0 IRQ_top3
port 108 nsew signal output
flabel metal2 s 3238 11194 3294 11250 0 FreeSans 224 0 0 0 N1BEG[0]
port 109 nsew signal output
flabel metal2 s 3514 11194 3570 11250 0 FreeSans 224 0 0 0 N1BEG[1]
port 110 nsew signal output
flabel metal2 s 3790 11194 3846 11250 0 FreeSans 224 0 0 0 N1BEG[2]
port 111 nsew signal output
flabel metal2 s 4066 11194 4122 11250 0 FreeSans 224 0 0 0 N1BEG[3]
port 112 nsew signal output
flabel metal2 s 4342 11194 4398 11250 0 FreeSans 224 0 0 0 N2BEG[0]
port 113 nsew signal output
flabel metal2 s 4618 11194 4674 11250 0 FreeSans 224 0 0 0 N2BEG[1]
port 114 nsew signal output
flabel metal2 s 4894 11194 4950 11250 0 FreeSans 224 0 0 0 N2BEG[2]
port 115 nsew signal output
flabel metal2 s 5170 11194 5226 11250 0 FreeSans 224 0 0 0 N2BEG[3]
port 116 nsew signal output
flabel metal2 s 5446 11194 5502 11250 0 FreeSans 224 0 0 0 N2BEG[4]
port 117 nsew signal output
flabel metal2 s 5722 11194 5778 11250 0 FreeSans 224 0 0 0 N2BEG[5]
port 118 nsew signal output
flabel metal2 s 5998 11194 6054 11250 0 FreeSans 224 0 0 0 N2BEG[6]
port 119 nsew signal output
flabel metal2 s 6274 11194 6330 11250 0 FreeSans 224 0 0 0 N2BEG[7]
port 120 nsew signal output
flabel metal2 s 6550 11194 6606 11250 0 FreeSans 224 0 0 0 N2BEGb[0]
port 121 nsew signal output
flabel metal2 s 6826 11194 6882 11250 0 FreeSans 224 0 0 0 N2BEGb[1]
port 122 nsew signal output
flabel metal2 s 7102 11194 7158 11250 0 FreeSans 224 0 0 0 N2BEGb[2]
port 123 nsew signal output
flabel metal2 s 7378 11194 7434 11250 0 FreeSans 224 0 0 0 N2BEGb[3]
port 124 nsew signal output
flabel metal2 s 7654 11194 7710 11250 0 FreeSans 224 0 0 0 N2BEGb[4]
port 125 nsew signal output
flabel metal2 s 7930 11194 7986 11250 0 FreeSans 224 0 0 0 N2BEGb[5]
port 126 nsew signal output
flabel metal2 s 8206 11194 8262 11250 0 FreeSans 224 0 0 0 N2BEGb[6]
port 127 nsew signal output
flabel metal2 s 8482 11194 8538 11250 0 FreeSans 224 0 0 0 N2BEGb[7]
port 128 nsew signal output
flabel metal2 s 8758 11194 8814 11250 0 FreeSans 224 0 0 0 N4BEG[0]
port 129 nsew signal output
flabel metal2 s 11518 11194 11574 11250 0 FreeSans 224 0 0 0 N4BEG[10]
port 130 nsew signal output
flabel metal2 s 11794 11194 11850 11250 0 FreeSans 224 0 0 0 N4BEG[11]
port 131 nsew signal output
flabel metal2 s 12070 11194 12126 11250 0 FreeSans 224 0 0 0 N4BEG[12]
port 132 nsew signal output
flabel metal2 s 12346 11194 12402 11250 0 FreeSans 224 0 0 0 N4BEG[13]
port 133 nsew signal output
flabel metal2 s 12622 11194 12678 11250 0 FreeSans 224 0 0 0 N4BEG[14]
port 134 nsew signal output
flabel metal2 s 12898 11194 12954 11250 0 FreeSans 224 0 0 0 N4BEG[15]
port 135 nsew signal output
flabel metal2 s 9034 11194 9090 11250 0 FreeSans 224 0 0 0 N4BEG[1]
port 136 nsew signal output
flabel metal2 s 9310 11194 9366 11250 0 FreeSans 224 0 0 0 N4BEG[2]
port 137 nsew signal output
flabel metal2 s 9586 11194 9642 11250 0 FreeSans 224 0 0 0 N4BEG[3]
port 138 nsew signal output
flabel metal2 s 9862 11194 9918 11250 0 FreeSans 224 0 0 0 N4BEG[4]
port 139 nsew signal output
flabel metal2 s 10138 11194 10194 11250 0 FreeSans 224 0 0 0 N4BEG[5]
port 140 nsew signal output
flabel metal2 s 10414 11194 10470 11250 0 FreeSans 224 0 0 0 N4BEG[6]
port 141 nsew signal output
flabel metal2 s 10690 11194 10746 11250 0 FreeSans 224 0 0 0 N4BEG[7]
port 142 nsew signal output
flabel metal2 s 10966 11194 11022 11250 0 FreeSans 224 0 0 0 N4BEG[8]
port 143 nsew signal output
flabel metal2 s 11242 11194 11298 11250 0 FreeSans 224 0 0 0 N4BEG[9]
port 144 nsew signal output
flabel metal2 s 13174 11194 13230 11250 0 FreeSans 224 0 0 0 NN4BEG[0]
port 145 nsew signal output
flabel metal2 s 15934 11194 15990 11250 0 FreeSans 224 0 0 0 NN4BEG[10]
port 146 nsew signal output
flabel metal2 s 16210 11194 16266 11250 0 FreeSans 224 0 0 0 NN4BEG[11]
port 147 nsew signal output
flabel metal2 s 16486 11194 16542 11250 0 FreeSans 224 0 0 0 NN4BEG[12]
port 148 nsew signal output
flabel metal2 s 16762 11194 16818 11250 0 FreeSans 224 0 0 0 NN4BEG[13]
port 149 nsew signal output
flabel metal2 s 17038 11194 17094 11250 0 FreeSans 224 0 0 0 NN4BEG[14]
port 150 nsew signal output
flabel metal2 s 17314 11194 17370 11250 0 FreeSans 224 0 0 0 NN4BEG[15]
port 151 nsew signal output
flabel metal2 s 13450 11194 13506 11250 0 FreeSans 224 0 0 0 NN4BEG[1]
port 152 nsew signal output
flabel metal2 s 13726 11194 13782 11250 0 FreeSans 224 0 0 0 NN4BEG[2]
port 153 nsew signal output
flabel metal2 s 14002 11194 14058 11250 0 FreeSans 224 0 0 0 NN4BEG[3]
port 154 nsew signal output
flabel metal2 s 14278 11194 14334 11250 0 FreeSans 224 0 0 0 NN4BEG[4]
port 155 nsew signal output
flabel metal2 s 14554 11194 14610 11250 0 FreeSans 224 0 0 0 NN4BEG[5]
port 156 nsew signal output
flabel metal2 s 14830 11194 14886 11250 0 FreeSans 224 0 0 0 NN4BEG[6]
port 157 nsew signal output
flabel metal2 s 15106 11194 15162 11250 0 FreeSans 224 0 0 0 NN4BEG[7]
port 158 nsew signal output
flabel metal2 s 15382 11194 15438 11250 0 FreeSans 224 0 0 0 NN4BEG[8]
port 159 nsew signal output
flabel metal2 s 15658 11194 15714 11250 0 FreeSans 224 0 0 0 NN4BEG[9]
port 160 nsew signal output
flabel metal2 s 17866 11194 17922 11250 0 FreeSans 224 0 0 0 S1END[0]
port 161 nsew signal input
flabel metal2 s 18142 11194 18198 11250 0 FreeSans 224 0 0 0 S1END[1]
port 162 nsew signal input
flabel metal2 s 18418 11194 18474 11250 0 FreeSans 224 0 0 0 S1END[2]
port 163 nsew signal input
flabel metal2 s 18694 11194 18750 11250 0 FreeSans 224 0 0 0 S1END[3]
port 164 nsew signal input
flabel metal2 s 21178 11194 21234 11250 0 FreeSans 224 0 0 0 S2END[0]
port 165 nsew signal input
flabel metal2 s 21454 11194 21510 11250 0 FreeSans 224 0 0 0 S2END[1]
port 166 nsew signal input
flabel metal2 s 21730 11194 21786 11250 0 FreeSans 224 0 0 0 S2END[2]
port 167 nsew signal input
flabel metal2 s 22006 11194 22062 11250 0 FreeSans 224 0 0 0 S2END[3]
port 168 nsew signal input
flabel metal2 s 22282 11194 22338 11250 0 FreeSans 224 0 0 0 S2END[4]
port 169 nsew signal input
flabel metal2 s 22558 11194 22614 11250 0 FreeSans 224 0 0 0 S2END[5]
port 170 nsew signal input
flabel metal2 s 22834 11194 22890 11250 0 FreeSans 224 0 0 0 S2END[6]
port 171 nsew signal input
flabel metal2 s 23110 11194 23166 11250 0 FreeSans 224 0 0 0 S2END[7]
port 172 nsew signal input
flabel metal2 s 18970 11194 19026 11250 0 FreeSans 224 0 0 0 S2MID[0]
port 173 nsew signal input
flabel metal2 s 19246 11194 19302 11250 0 FreeSans 224 0 0 0 S2MID[1]
port 174 nsew signal input
flabel metal2 s 19522 11194 19578 11250 0 FreeSans 224 0 0 0 S2MID[2]
port 175 nsew signal input
flabel metal2 s 19798 11194 19854 11250 0 FreeSans 224 0 0 0 S2MID[3]
port 176 nsew signal input
flabel metal2 s 20074 11194 20130 11250 0 FreeSans 224 0 0 0 S2MID[4]
port 177 nsew signal input
flabel metal2 s 20350 11194 20406 11250 0 FreeSans 224 0 0 0 S2MID[5]
port 178 nsew signal input
flabel metal2 s 20626 11194 20682 11250 0 FreeSans 224 0 0 0 S2MID[6]
port 179 nsew signal input
flabel metal2 s 20902 11194 20958 11250 0 FreeSans 224 0 0 0 S2MID[7]
port 180 nsew signal input
flabel metal2 s 23386 11194 23442 11250 0 FreeSans 224 0 0 0 S4END[0]
port 181 nsew signal input
flabel metal2 s 26146 11194 26202 11250 0 FreeSans 224 0 0 0 S4END[10]
port 182 nsew signal input
flabel metal2 s 26422 11194 26478 11250 0 FreeSans 224 0 0 0 S4END[11]
port 183 nsew signal input
flabel metal2 s 26698 11194 26754 11250 0 FreeSans 224 0 0 0 S4END[12]
port 184 nsew signal input
flabel metal2 s 26974 11194 27030 11250 0 FreeSans 224 0 0 0 S4END[13]
port 185 nsew signal input
flabel metal2 s 27250 11194 27306 11250 0 FreeSans 224 0 0 0 S4END[14]
port 186 nsew signal input
flabel metal2 s 27526 11194 27582 11250 0 FreeSans 224 0 0 0 S4END[15]
port 187 nsew signal input
flabel metal2 s 23662 11194 23718 11250 0 FreeSans 224 0 0 0 S4END[1]
port 188 nsew signal input
flabel metal2 s 23938 11194 23994 11250 0 FreeSans 224 0 0 0 S4END[2]
port 189 nsew signal input
flabel metal2 s 24214 11194 24270 11250 0 FreeSans 224 0 0 0 S4END[3]
port 190 nsew signal input
flabel metal2 s 24490 11194 24546 11250 0 FreeSans 224 0 0 0 S4END[4]
port 191 nsew signal input
flabel metal2 s 24766 11194 24822 11250 0 FreeSans 224 0 0 0 S4END[5]
port 192 nsew signal input
flabel metal2 s 25042 11194 25098 11250 0 FreeSans 224 0 0 0 S4END[6]
port 193 nsew signal input
flabel metal2 s 25318 11194 25374 11250 0 FreeSans 224 0 0 0 S4END[7]
port 194 nsew signal input
flabel metal2 s 25594 11194 25650 11250 0 FreeSans 224 0 0 0 S4END[8]
port 195 nsew signal input
flabel metal2 s 25870 11194 25926 11250 0 FreeSans 224 0 0 0 S4END[9]
port 196 nsew signal input
flabel metal2 s 27802 11194 27858 11250 0 FreeSans 224 0 0 0 SS4END[0]
port 197 nsew signal input
flabel metal2 s 30562 11194 30618 11250 0 FreeSans 224 0 0 0 SS4END[10]
port 198 nsew signal input
flabel metal2 s 30838 11194 30894 11250 0 FreeSans 224 0 0 0 SS4END[11]
port 199 nsew signal input
flabel metal2 s 31114 11194 31170 11250 0 FreeSans 224 0 0 0 SS4END[12]
port 200 nsew signal input
flabel metal2 s 31390 11194 31446 11250 0 FreeSans 224 0 0 0 SS4END[13]
port 201 nsew signal input
flabel metal2 s 31666 11194 31722 11250 0 FreeSans 224 0 0 0 SS4END[14]
port 202 nsew signal input
flabel metal2 s 31942 11194 31998 11250 0 FreeSans 224 0 0 0 SS4END[15]
port 203 nsew signal input
flabel metal2 s 28078 11194 28134 11250 0 FreeSans 224 0 0 0 SS4END[1]
port 204 nsew signal input
flabel metal2 s 28354 11194 28410 11250 0 FreeSans 224 0 0 0 SS4END[2]
port 205 nsew signal input
flabel metal2 s 28630 11194 28686 11250 0 FreeSans 224 0 0 0 SS4END[3]
port 206 nsew signal input
flabel metal2 s 28906 11194 28962 11250 0 FreeSans 224 0 0 0 SS4END[4]
port 207 nsew signal input
flabel metal2 s 29182 11194 29238 11250 0 FreeSans 224 0 0 0 SS4END[5]
port 208 nsew signal input
flabel metal2 s 29458 11194 29514 11250 0 FreeSans 224 0 0 0 SS4END[6]
port 209 nsew signal input
flabel metal2 s 29734 11194 29790 11250 0 FreeSans 224 0 0 0 SS4END[7]
port 210 nsew signal input
flabel metal2 s 30010 11194 30066 11250 0 FreeSans 224 0 0 0 SS4END[8]
port 211 nsew signal input
flabel metal2 s 30286 11194 30342 11250 0 FreeSans 224 0 0 0 SS4END[9]
port 212 nsew signal input
flabel metal2 s 7930 0 7986 56 0 FreeSans 224 0 0 0 UserCLK
port 213 nsew signal input
flabel metal2 s 32218 11194 32274 11250 0 FreeSans 224 0 0 0 UserCLKo
port 214 nsew signal output
flabel metal4 s 3004 0 3324 11250 0 FreeSans 1920 90 0 0 VGND
port 215 nsew ground bidirectional
flabel metal4 s 3004 0 3324 60 0 FreeSans 480 0 0 0 VGND
port 215 nsew ground bidirectional
flabel metal4 s 3004 11190 3324 11250 0 FreeSans 480 0 0 0 VGND
port 215 nsew ground bidirectional
flabel metal4 s 9004 0 9324 11250 0 FreeSans 1920 90 0 0 VGND
port 215 nsew ground bidirectional
flabel metal4 s 9004 0 9324 60 0 FreeSans 480 0 0 0 VGND
port 215 nsew ground bidirectional
flabel metal4 s 9004 11190 9324 11250 0 FreeSans 480 0 0 0 VGND
port 215 nsew ground bidirectional
flabel metal4 s 15004 0 15324 11250 0 FreeSans 1920 90 0 0 VGND
port 215 nsew ground bidirectional
flabel metal4 s 15004 0 15324 60 0 FreeSans 480 0 0 0 VGND
port 215 nsew ground bidirectional
flabel metal4 s 15004 11190 15324 11250 0 FreeSans 480 0 0 0 VGND
port 215 nsew ground bidirectional
flabel metal4 s 21004 0 21324 11250 0 FreeSans 1920 90 0 0 VGND
port 215 nsew ground bidirectional
flabel metal4 s 21004 0 21324 60 0 FreeSans 480 0 0 0 VGND
port 215 nsew ground bidirectional
flabel metal4 s 21004 11190 21324 11250 0 FreeSans 480 0 0 0 VGND
port 215 nsew ground bidirectional
flabel metal4 s 27004 0 27324 11250 0 FreeSans 1920 90 0 0 VGND
port 215 nsew ground bidirectional
flabel metal4 s 27004 0 27324 60 0 FreeSans 480 0 0 0 VGND
port 215 nsew ground bidirectional
flabel metal4 s 27004 11190 27324 11250 0 FreeSans 480 0 0 0 VGND
port 215 nsew ground bidirectional
flabel metal4 s 33004 0 33324 11250 0 FreeSans 1920 90 0 0 VGND
port 215 nsew ground bidirectional
flabel metal4 s 33004 0 33324 60 0 FreeSans 480 0 0 0 VGND
port 215 nsew ground bidirectional
flabel metal4 s 33004 11190 33324 11250 0 FreeSans 480 0 0 0 VGND
port 215 nsew ground bidirectional
flabel metal4 s 39004 0 39324 11250 0 FreeSans 1920 90 0 0 VGND
port 215 nsew ground bidirectional
flabel metal4 s 39004 0 39324 60 0 FreeSans 480 0 0 0 VGND
port 215 nsew ground bidirectional
flabel metal4 s 39004 11190 39324 11250 0 FreeSans 480 0 0 0 VGND
port 215 nsew ground bidirectional
flabel metal4 s 1944 0 2264 11250 0 FreeSans 1920 90 0 0 VPWR
port 216 nsew power bidirectional
flabel metal4 s 1944 0 2264 60 0 FreeSans 480 0 0 0 VPWR
port 216 nsew power bidirectional
flabel metal4 s 1944 11190 2264 11250 0 FreeSans 480 0 0 0 VPWR
port 216 nsew power bidirectional
flabel metal4 s 7944 0 8264 11250 0 FreeSans 1920 90 0 0 VPWR
port 216 nsew power bidirectional
flabel metal4 s 7944 0 8264 60 0 FreeSans 480 0 0 0 VPWR
port 216 nsew power bidirectional
flabel metal4 s 7944 11190 8264 11250 0 FreeSans 480 0 0 0 VPWR
port 216 nsew power bidirectional
flabel metal4 s 13944 0 14264 11250 0 FreeSans 1920 90 0 0 VPWR
port 216 nsew power bidirectional
flabel metal4 s 13944 0 14264 60 0 FreeSans 480 0 0 0 VPWR
port 216 nsew power bidirectional
flabel metal4 s 13944 11190 14264 11250 0 FreeSans 480 0 0 0 VPWR
port 216 nsew power bidirectional
flabel metal4 s 19944 0 20264 11250 0 FreeSans 1920 90 0 0 VPWR
port 216 nsew power bidirectional
flabel metal4 s 19944 0 20264 60 0 FreeSans 480 0 0 0 VPWR
port 216 nsew power bidirectional
flabel metal4 s 19944 11190 20264 11250 0 FreeSans 480 0 0 0 VPWR
port 216 nsew power bidirectional
flabel metal4 s 25944 0 26264 11250 0 FreeSans 1920 90 0 0 VPWR
port 216 nsew power bidirectional
flabel metal4 s 25944 0 26264 60 0 FreeSans 480 0 0 0 VPWR
port 216 nsew power bidirectional
flabel metal4 s 25944 11190 26264 11250 0 FreeSans 480 0 0 0 VPWR
port 216 nsew power bidirectional
flabel metal4 s 31944 0 32264 11250 0 FreeSans 1920 90 0 0 VPWR
port 216 nsew power bidirectional
flabel metal4 s 31944 0 32264 60 0 FreeSans 480 0 0 0 VPWR
port 216 nsew power bidirectional
flabel metal4 s 31944 11190 32264 11250 0 FreeSans 480 0 0 0 VPWR
port 216 nsew power bidirectional
flabel metal4 s 37944 0 38264 11250 0 FreeSans 1920 90 0 0 VPWR
port 216 nsew power bidirectional
flabel metal4 s 37944 0 38264 60 0 FreeSans 480 0 0 0 VPWR
port 216 nsew power bidirectional
flabel metal4 s 37944 11190 38264 11250 0 FreeSans 480 0 0 0 VPWR
port 216 nsew power bidirectional
rlabel metal1 20470 8704 20470 8704 0 VGND
rlabel metal1 20470 8160 20470 8160 0 VPWR
rlabel metal1 37904 3502 37904 3502 0 FrameData[0]
rlabel metal3 390 4148 390 4148 0 FrameData[10]
rlabel metal2 2898 5015 2898 5015 0 FrameData[11]
rlabel metal3 712 4692 712 4692 0 FrameData[12]
rlabel metal3 827 4964 827 4964 0 FrameData[13]
rlabel metal3 13708 7208 13708 7208 0 FrameData[14]
rlabel metal3 666 5508 666 5508 0 FrameData[15]
rlabel metal2 4094 6579 4094 6579 0 FrameData[16]
rlabel metal3 919 6052 919 6052 0 FrameData[17]
rlabel metal2 2898 6851 2898 6851 0 FrameData[18]
rlabel metal3 344 6596 344 6596 0 FrameData[19]
rlabel metal3 666 1700 666 1700 0 FrameData[1]
rlabel metal3 528 6868 528 6868 0 FrameData[20]
rlabel metal3 436 7140 436 7140 0 FrameData[21]
rlabel metal3 344 7412 344 7412 0 FrameData[22]
rlabel metal3 436 7684 436 7684 0 FrameData[23]
rlabel metal3 344 7956 344 7956 0 FrameData[24]
rlabel metal3 574 8228 574 8228 0 FrameData[25]
rlabel metal3 712 8500 712 8500 0 FrameData[26]
rlabel metal3 528 8772 528 8772 0 FrameData[27]
rlabel metal3 666 9044 666 9044 0 FrameData[28]
rlabel metal3 482 9316 482 9316 0 FrameData[29]
rlabel metal1 38410 3468 38410 3468 0 FrameData[2]
rlabel metal3 574 9588 574 9588 0 FrameData[30]
rlabel metal3 620 9860 620 9860 0 FrameData[31]
rlabel metal3 1494 2244 1494 2244 0 FrameData[3]
rlabel metal3 712 2516 712 2516 0 FrameData[4]
rlabel metal3 919 2788 919 2788 0 FrameData[5]
rlabel metal3 712 3060 712 3060 0 FrameData[6]
rlabel metal2 2898 3723 2898 3723 0 FrameData[7]
rlabel metal2 2806 4063 2806 4063 0 FrameData[8]
rlabel metal3 919 3876 919 3876 0 FrameData[9]
rlabel metal3 39798 1428 39798 1428 0 FrameData_O[0]
rlabel metal2 39422 3927 39422 3927 0 FrameData_O[10]
rlabel metal3 40166 4420 40166 4420 0 FrameData_O[11]
rlabel metal1 39468 3978 39468 3978 0 FrameData_O[12]
rlabel metal3 39982 4964 39982 4964 0 FrameData_O[13]
rlabel metal2 39422 5015 39422 5015 0 FrameData_O[14]
rlabel metal3 40166 5508 40166 5508 0 FrameData_O[15]
rlabel metal1 39468 5338 39468 5338 0 FrameData_O[16]
rlabel metal3 39982 6052 39982 6052 0 FrameData_O[17]
rlabel metal3 39798 6324 39798 6324 0 FrameData_O[18]
rlabel metal1 39514 5882 39514 5882 0 FrameData_O[19]
rlabel metal3 39614 1700 39614 1700 0 FrameData_O[1]
rlabel metal3 40212 6868 40212 6868 0 FrameData_O[20]
rlabel metal2 39422 6885 39422 6885 0 FrameData_O[21]
rlabel metal3 39936 7412 39936 7412 0 FrameData_O[22]
rlabel metal3 40166 7684 40166 7684 0 FrameData_O[23]
rlabel metal3 40166 7956 40166 7956 0 FrameData_O[24]
rlabel metal1 39054 7480 39054 7480 0 FrameData_O[25]
rlabel metal2 38686 8279 38686 8279 0 FrameData_O[26]
rlabel metal1 39468 7514 39468 7514 0 FrameData_O[27]
rlabel metal1 39744 6426 39744 6426 0 FrameData_O[28]
rlabel metal1 38732 7514 38732 7514 0 FrameData_O[29]
rlabel metal3 39384 1972 39384 1972 0 FrameData_O[2]
rlabel metal1 39054 6664 39054 6664 0 FrameData_O[30]
rlabel metal2 38318 8687 38318 8687 0 FrameData_O[31]
rlabel metal3 40442 2244 40442 2244 0 FrameData_O[3]
rlabel metal3 39246 2516 39246 2516 0 FrameData_O[4]
rlabel metal3 39890 2788 39890 2788 0 FrameData_O[5]
rlabel metal3 40166 3060 40166 3060 0 FrameData_O[6]
rlabel metal1 39238 3162 39238 3162 0 FrameData_O[7]
rlabel metal1 39468 2890 39468 2890 0 FrameData_O[8]
rlabel metal3 39982 3876 39982 3876 0 FrameData_O[9]
rlabel metal2 9522 1228 9522 1228 0 FrameStrobe[0]
rlabel metal2 25162 446 25162 446 0 FrameStrobe[10]
rlabel metal2 32430 6256 32430 6256 0 FrameStrobe[11]
rlabel metal2 32614 5678 32614 5678 0 FrameStrobe[12]
rlabel via2 34270 7395 34270 7395 0 FrameStrobe[13]
rlabel metal2 31418 3166 31418 3166 0 FrameStrobe[14]
rlabel metal2 32982 55 32982 55 0 FrameStrobe[15]
rlabel metal2 34546 939 34546 939 0 FrameStrobe[16]
rlabel metal1 36800 5202 36800 5202 0 FrameStrobe[17]
rlabel metal1 37812 5202 37812 5202 0 FrameStrobe[18]
rlabel metal2 39238 55 39238 55 0 FrameStrobe[19]
rlabel metal2 11086 939 11086 939 0 FrameStrobe[1]
rlabel metal2 12650 1279 12650 1279 0 FrameStrobe[2]
rlabel metal2 14214 106 14214 106 0 FrameStrobe[3]
rlabel via2 15778 55 15778 55 0 FrameStrobe[4]
rlabel metal3 18860 3060 18860 3060 0 FrameStrobe[5]
rlabel metal2 18906 123 18906 123 0 FrameStrobe[6]
rlabel metal2 20470 1058 20470 1058 0 FrameStrobe[7]
rlabel metal2 22034 1500 22034 1500 0 FrameStrobe[8]
rlabel metal1 23966 3366 23966 3366 0 FrameStrobe[9]
rlabel metal1 32660 8602 32660 8602 0 FrameStrobe_O[0]
rlabel metal1 36340 8262 36340 8262 0 FrameStrobe_O[10]
rlabel metal1 35696 8058 35696 8058 0 FrameStrobe_O[11]
rlabel metal1 36294 8602 36294 8602 0 FrameStrobe_O[12]
rlabel metal1 36248 8058 36248 8058 0 FrameStrobe_O[13]
rlabel metal1 37306 8262 37306 8262 0 FrameStrobe_O[14]
rlabel metal1 36800 8058 36800 8058 0 FrameStrobe_O[15]
rlabel metal1 37398 8602 37398 8602 0 FrameStrobe_O[16]
rlabel metal1 37720 8330 37720 8330 0 FrameStrobe_O[17]
rlabel metal1 38594 8568 38594 8568 0 FrameStrobe_O[18]
rlabel metal1 37858 8058 37858 8058 0 FrameStrobe_O[19]
rlabel metal1 33028 8602 33028 8602 0 FrameStrobe_O[1]
rlabel metal2 33534 8704 33534 8704 0 FrameStrobe_O[2]
rlabel metal1 33672 8330 33672 8330 0 FrameStrobe_O[3]
rlabel metal1 33948 8602 33948 8602 0 FrameStrobe_O[4]
rlabel metal1 34454 8330 34454 8330 0 FrameStrobe_O[5]
rlabel metal1 35282 8364 35282 8364 0 FrameStrobe_O[6]
rlabel metal1 34684 8058 34684 8058 0 FrameStrobe_O[7]
rlabel metal1 35144 8602 35144 8602 0 FrameStrobe_O[8]
rlabel metal1 35834 8330 35834 8330 0 FrameStrobe_O[9]
rlabel metal2 1702 1160 1702 1160 0 IRQ_top0
rlabel metal2 3266 55 3266 55 0 IRQ_top1
rlabel metal2 4830 1160 4830 1160 0 IRQ_top2
rlabel metal2 6394 1160 6394 1160 0 IRQ_top3
rlabel metal1 17710 3502 17710 3502 0 Inst_S_CPU_IRQ_ConfigMem.Inst_frame0_bit20.Q
rlabel metal1 21390 6630 21390 6630 0 Inst_S_CPU_IRQ_ConfigMem.Inst_frame0_bit21.Q
rlabel metal1 20102 3502 20102 3502 0 Inst_S_CPU_IRQ_ConfigMem.Inst_frame0_bit22.Q
rlabel metal2 12742 5916 12742 5916 0 Inst_S_CPU_IRQ_ConfigMem.Inst_frame0_bit23.Q
rlabel metal1 13294 4624 13294 4624 0 Inst_S_CPU_IRQ_ConfigMem.Inst_frame0_bit24.Q
rlabel metal1 15410 3400 15410 3400 0 Inst_S_CPU_IRQ_ConfigMem.Inst_frame0_bit25.Q
rlabel via1 15501 3502 15501 3502 0 Inst_S_CPU_IRQ_ConfigMem.Inst_frame0_bit26.Q
rlabel via1 14582 6290 14582 6290 0 Inst_S_CPU_IRQ_ConfigMem.Inst_frame0_bit27.Q
rlabel metal2 19734 4165 19734 4165 0 Inst_S_CPU_IRQ_ConfigMem.Inst_frame0_bit28.Q
rlabel metal1 21758 3604 21758 3604 0 Inst_S_CPU_IRQ_ConfigMem.Inst_frame0_bit29.Q
rlabel metal1 22862 3570 22862 3570 0 Inst_S_CPU_IRQ_ConfigMem.Inst_frame0_bit30.Q
rlabel metal1 20746 6426 20746 6426 0 Inst_S_CPU_IRQ_ConfigMem.Inst_frame0_bit31.Q
rlabel metal2 3450 8755 3450 8755 0 N1BEG[0]
rlabel metal1 3312 8330 3312 8330 0 N1BEG[1]
rlabel metal1 3634 8602 3634 8602 0 N1BEG[2]
rlabel metal1 4186 8058 4186 8058 0 N1BEG[3]
rlabel metal1 4324 8602 4324 8602 0 N2BEG[0]
rlabel metal2 4646 9904 4646 9904 0 N2BEG[1]
rlabel metal1 5060 8058 5060 8058 0 N2BEG[2]
rlabel metal1 5106 8602 5106 8602 0 N2BEG[3]
rlabel metal1 5382 8602 5382 8602 0 N2BEG[4]
rlabel metal1 5704 8602 5704 8602 0 N2BEG[5]
rlabel metal1 6118 8058 6118 8058 0 N2BEG[6]
rlabel metal1 6164 8602 6164 8602 0 N2BEG[7]
rlabel metal1 6670 8058 6670 8058 0 N2BEGb[0]
rlabel metal1 6808 8602 6808 8602 0 N2BEGb[1]
rlabel metal1 7222 8058 7222 8058 0 N2BEGb[2]
rlabel metal1 7268 8602 7268 8602 0 N2BEGb[3]
rlabel metal1 7590 8602 7590 8602 0 N2BEGb[4]
rlabel metal1 7912 8602 7912 8602 0 N2BEGb[5]
rlabel metal1 8418 8058 8418 8058 0 N2BEGb[6]
rlabel metal1 8372 8602 8372 8602 0 N2BEGb[7]
rlabel metal1 8924 8058 8924 8058 0 N4BEG[0]
rlabel metal1 11408 8602 11408 8602 0 N4BEG[10]
rlabel metal1 11914 8058 11914 8058 0 N4BEG[11]
rlabel metal1 11868 8602 11868 8602 0 N4BEG[12]
rlabel metal1 12236 8602 12236 8602 0 N4BEG[13]
rlabel metal1 12788 8058 12788 8058 0 N4BEG[14]
rlabel metal1 12696 8330 12696 8330 0 N4BEG[15]
rlabel metal1 8740 8602 8740 8602 0 N4BEG[1]
rlabel metal1 9476 8058 9476 8058 0 N4BEG[2]
rlabel metal1 9476 8602 9476 8602 0 N4BEG[3]
rlabel metal1 9798 8602 9798 8602 0 N4BEG[4]
rlabel metal1 10120 8602 10120 8602 0 N4BEG[5]
rlabel metal1 10534 8058 10534 8058 0 N4BEG[6]
rlabel metal1 10580 8602 10580 8602 0 N4BEG[7]
rlabel metal1 10902 8602 10902 8602 0 N4BEG[8]
rlabel metal1 11362 8058 11362 8058 0 N4BEG[9]
rlabel metal1 13018 8602 13018 8602 0 NN4BEG[0]
rlabel metal1 16100 8058 16100 8058 0 NN4BEG[10]
rlabel metal1 16100 8602 16100 8602 0 NN4BEG[11]
rlabel metal1 16422 8602 16422 8602 0 NN4BEG[12]
rlabel metal1 16928 8602 16928 8602 0 NN4BEG[13]
rlabel metal1 17526 8330 17526 8330 0 NN4BEG[14]
rlabel metal1 17480 8602 17480 8602 0 NN4BEG[15]
rlabel metal1 13570 8058 13570 8058 0 NN4BEG[1]
rlabel metal1 13478 8330 13478 8330 0 NN4BEG[2]
rlabel metal1 13938 8602 13938 8602 0 NN4BEG[3]
rlabel metal1 14398 8058 14398 8058 0 NN4BEG[4]
rlabel metal1 14536 8602 14536 8602 0 NN4BEG[5]
rlabel metal1 14950 8058 14950 8058 0 NN4BEG[6]
rlabel metal1 14904 8602 14904 8602 0 NN4BEG[7]
rlabel metal1 15318 8602 15318 8602 0 NN4BEG[8]
rlabel metal2 15686 9904 15686 9904 0 NN4BEG[9]
rlabel metal2 17894 9530 17894 9530 0 S1END[0]
rlabel metal2 18170 9530 18170 9530 0 S1END[1]
rlabel metal2 18446 9836 18446 9836 0 S1END[2]
rlabel metal2 18722 9836 18722 9836 0 S1END[3]
rlabel metal2 21206 10533 21206 10533 0 S2END[0]
rlabel metal2 21482 9836 21482 9836 0 S2END[1]
rlabel metal2 21758 9870 21758 9870 0 S2END[2]
rlabel metal2 22034 9904 22034 9904 0 S2END[3]
rlabel metal2 22310 10533 22310 10533 0 S2END[4]
rlabel metal2 22586 9870 22586 9870 0 S2END[5]
rlabel metal2 22862 10533 22862 10533 0 S2END[6]
rlabel metal2 23138 9904 23138 9904 0 S2END[7]
rlabel metal2 18998 9836 18998 9836 0 S2MID[0]
rlabel metal2 19274 9836 19274 9836 0 S2MID[1]
rlabel metal2 19550 9904 19550 9904 0 S2MID[2]
rlabel metal2 19826 9836 19826 9836 0 S2MID[3]
rlabel via1 20102 11196 20102 11196 0 S2MID[4]
rlabel metal2 20378 9734 20378 9734 0 S2MID[5]
rlabel metal2 20654 11128 20654 11128 0 S2MID[6]
rlabel metal2 20930 11162 20930 11162 0 S2MID[7]
rlabel metal2 23414 9768 23414 9768 0 S4END[0]
rlabel metal1 27324 8806 27324 8806 0 S4END[10]
rlabel metal1 26956 6834 26956 6834 0 S4END[11]
rlabel metal2 26726 8782 26726 8782 0 S4END[12]
rlabel metal2 27002 10125 27002 10125 0 S4END[13]
rlabel metal2 27278 10193 27278 10193 0 S4END[14]
rlabel metal2 27554 8714 27554 8714 0 S4END[15]
rlabel metal2 23690 9870 23690 9870 0 S4END[1]
rlabel metal2 23966 9904 23966 9904 0 S4END[2]
rlabel metal2 24242 10533 24242 10533 0 S4END[3]
rlabel metal2 24518 9870 24518 9870 0 S4END[4]
rlabel metal2 24794 9904 24794 9904 0 S4END[5]
rlabel metal2 25070 9802 25070 9802 0 S4END[6]
rlabel metal2 25346 9870 25346 9870 0 S4END[7]
rlabel metal1 26588 6902 26588 6902 0 S4END[8]
rlabel metal2 25898 10108 25898 10108 0 S4END[9]
rlabel metal2 27830 9836 27830 9836 0 SS4END[0]
rlabel metal1 31786 7412 31786 7412 0 SS4END[10]
rlabel metal1 32338 7446 32338 7446 0 SS4END[11]
rlabel metal2 32614 7548 32614 7548 0 SS4END[12]
rlabel metal2 31418 8986 31418 8986 0 SS4END[13]
rlabel metal1 32890 7344 32890 7344 0 SS4END[14]
rlabel metal2 31970 10125 31970 10125 0 SS4END[15]
rlabel metal2 28106 10533 28106 10533 0 SS4END[1]
rlabel metal2 28382 9836 28382 9836 0 SS4END[2]
rlabel metal2 28658 9530 28658 9530 0 SS4END[3]
rlabel metal2 28934 9598 28934 9598 0 SS4END[4]
rlabel metal2 29210 9802 29210 9802 0 SS4END[5]
rlabel metal2 29486 9530 29486 9530 0 SS4END[6]
rlabel metal2 29762 9836 29762 9836 0 SS4END[7]
rlabel metal2 30038 9292 30038 9292 0 SS4END[8]
rlabel metal2 30314 9326 30314 9326 0 SS4END[9]
rlabel metal2 7958 55 7958 55 0 UserCLK
rlabel metal1 32292 8602 32292 8602 0 UserCLKo
rlabel metal2 23138 4658 23138 4658 0 _000_
rlabel metal1 14306 3706 14306 3706 0 _001_
rlabel metal1 9384 3706 9384 3706 0 _002_
rlabel metal1 20562 3638 20562 3638 0 _003_
rlabel metal1 22724 3706 22724 3706 0 _004_
rlabel metal1 22356 3162 22356 3162 0 _005_
rlabel metal2 23874 5304 23874 5304 0 _006_
rlabel metal1 22218 3706 22218 3706 0 _007_
rlabel metal1 22862 6222 22862 6222 0 _008_
rlabel metal1 12190 3706 12190 3706 0 _009_
rlabel metal2 15410 5032 15410 5032 0 _010_
rlabel metal1 16146 4794 16146 4794 0 _011_
rlabel metal1 14812 3978 14812 3978 0 _012_
rlabel metal2 14674 5882 14674 5882 0 _013_
rlabel metal1 8004 4046 8004 4046 0 _014_
rlabel metal1 9752 4114 9752 4114 0 _015_
rlabel metal1 10350 4794 10350 4794 0 _016_
rlabel metal1 9246 3978 9246 3978 0 _017_
rlabel metal2 10074 6460 10074 6460 0 _018_
rlabel metal1 17020 3706 17020 3706 0 _019_
rlabel metal1 18262 4080 18262 4080 0 _020_
rlabel metal2 22402 7582 22402 7582 0 _021_
rlabel metal1 19458 3706 19458 3706 0 _022_
rlabel metal2 22126 7072 22126 7072 0 _023_
rlabel metal1 2254 7174 2254 7174 0 net1
rlabel metal2 6302 7548 6302 7548 0 net10
rlabel metal1 4600 2346 4600 2346 0 net100
rlabel metal1 5198 2448 5198 2448 0 net101
rlabel metal2 6762 2244 6762 2244 0 net102
rlabel metal2 3634 8517 3634 8517 0 net103
rlabel metal2 7774 9112 7774 9112 0 net104
rlabel metal1 11730 6630 11730 6630 0 net105
rlabel via2 21758 4811 21758 4811 0 net106
rlabel metal1 3680 6630 3680 6630 0 net107
rlabel metal2 4002 7514 4002 7514 0 net108
rlabel metal2 4738 7684 4738 7684 0 net109
rlabel metal1 1978 8262 1978 8262 0 net11
rlabel metal1 4324 7514 4324 7514 0 net110
rlabel metal2 5658 9435 5658 9435 0 net111
rlabel metal1 15824 5882 15824 5882 0 net112
rlabel metal2 9890 7344 9890 7344 0 net113
rlabel metal2 19366 3230 19366 3230 0 net114
rlabel metal2 7222 8976 7222 8976 0 net115
rlabel metal1 17756 6086 17756 6086 0 net116
rlabel metal1 8924 5882 8924 5882 0 net117
rlabel metal1 15870 6426 15870 6426 0 net118
rlabel metal2 7682 8415 7682 8415 0 net119
rlabel metal2 2162 8738 2162 8738 0 net12
rlabel metal2 12006 7378 12006 7378 0 net120
rlabel metal1 7958 6426 7958 6426 0 net121
rlabel metal1 16744 4998 16744 4998 0 net122
rlabel metal3 14444 7616 14444 7616 0 net123
rlabel metal1 8096 5882 8096 5882 0 net124
rlabel metal2 12190 7684 12190 7684 0 net125
rlabel metal2 12558 8670 12558 8670 0 net126
rlabel metal2 13570 6596 13570 6596 0 net127
rlabel metal1 12581 7854 12581 7854 0 net128
rlabel metal2 18538 6511 18538 6511 0 net129
rlabel metal2 2438 8738 2438 8738 0 net13
rlabel metal2 8694 9095 8694 9095 0 net130
rlabel metal2 9706 8993 9706 8993 0 net131
rlabel metal2 9522 9112 9522 9112 0 net132
rlabel metal2 10074 9146 10074 9146 0 net133
rlabel metal2 10258 8959 10258 8959 0 net134
rlabel metal2 14352 7412 14352 7412 0 net135
rlabel metal2 10626 9248 10626 9248 0 net136
rlabel metal2 10902 9180 10902 9180 0 net137
rlabel metal2 13754 7378 13754 7378 0 net138
rlabel via2 13018 8483 13018 8483 0 net139
rlabel metal2 26358 3128 26358 3128 0 net14
rlabel metal2 13202 6222 13202 6222 0 net140
rlabel metal1 16836 5066 16836 5066 0 net141
rlabel metal2 16698 8976 16698 8976 0 net142
rlabel metal2 16882 8228 16882 8228 0 net143
rlabel metal2 14950 6885 14950 6885 0 net144
rlabel metal1 17250 5882 17250 5882 0 net145
rlabel metal1 21206 7344 21206 7344 0 net146
rlabel metal2 13386 8891 13386 8891 0 net147
rlabel metal1 13662 8432 13662 8432 0 net148
rlabel via2 14674 7837 14674 7837 0 net149
rlabel metal1 21344 4590 21344 4590 0 net15
rlabel metal2 14674 9214 14674 9214 0 net150
rlabel metal2 31326 7480 31326 7480 0 net151
rlabel metal1 30774 7174 30774 7174 0 net152
rlabel metal2 15502 8925 15502 8925 0 net153
rlabel metal2 15594 6120 15594 6120 0 net154
rlabel metal1 32131 8466 32131 8466 0 net155
rlabel metal1 17664 8058 17664 8058 0 net156
rlabel metal1 14490 6936 14490 6936 0 net16
rlabel metal1 17480 5678 17480 5678 0 net17
rlabel metal2 18814 8772 18814 8772 0 net18
rlabel metal1 21390 3502 21390 3502 0 net19
rlabel metal1 2185 7242 2185 7242 0 net2
rlabel metal2 18078 6154 18078 6154 0 net20
rlabel metal1 15410 4114 15410 4114 0 net21
rlabel metal1 22586 8364 22586 8364 0 net22
rlabel metal2 19366 7072 19366 7072 0 net23
rlabel metal2 9154 6052 9154 6052 0 net24
rlabel metal2 17986 7684 17986 7684 0 net25
rlabel metal1 23644 8262 23644 8262 0 net26
rlabel metal1 20792 5678 20792 5678 0 net27
rlabel metal2 19366 9078 19366 9078 0 net28
rlabel metal1 16422 5678 16422 5678 0 net29
rlabel metal2 15134 7072 15134 7072 0 net3
rlabel metal1 20102 8364 20102 8364 0 net30
rlabel metal1 19228 5678 19228 5678 0 net31
rlabel metal1 6624 5678 6624 5678 0 net32
rlabel metal2 13754 3740 13754 3740 0 net33
rlabel metal2 24242 7004 24242 7004 0 net34
rlabel metal2 24794 7752 24794 7752 0 net35
rlabel metal1 7590 5678 7590 5678 0 net36
rlabel metal1 13892 6766 13892 6766 0 net37
rlabel metal1 26358 5202 26358 5202 0 net38
rlabel metal2 21758 5661 21758 5661 0 net39
rlabel via1 2162 7939 2162 7939 0 net4
rlabel metal2 20378 6188 20378 6188 0 net40
rlabel metal1 23414 5678 23414 5678 0 net41
rlabel metal2 24610 6698 24610 6698 0 net42
rlabel metal1 20286 5236 20286 5236 0 net43
rlabel metal2 7314 4182 7314 4182 0 net44
rlabel metal1 11868 4590 11868 4590 0 net45
rlabel metal1 25300 5678 25300 5678 0 net46
rlabel metal1 38456 2414 38456 2414 0 net47
rlabel metal2 39238 3553 39238 3553 0 net48
rlabel metal1 38916 4590 38916 4590 0 net49
rlabel metal1 2070 7752 2070 7752 0 net5
rlabel metal1 39238 4080 39238 4080 0 net50
rlabel metal2 38870 4964 38870 4964 0 net51
rlabel metal1 39238 4624 39238 4624 0 net52
rlabel metal1 38732 5678 38732 5678 0 net53
rlabel via2 39238 5219 39238 5219 0 net54
rlabel metal2 21574 4845 21574 4845 0 net55
rlabel metal2 22034 6783 22034 6783 0 net56
rlabel metal1 39100 5678 39100 5678 0 net57
rlabel metal1 38134 2380 38134 2380 0 net58
rlabel metal3 20516 6528 20516 6528 0 net59
rlabel metal2 1610 8534 1610 8534 0 net6
rlabel metal1 38870 5304 38870 5304 0 net60
rlabel metal1 38870 7888 38870 7888 0 net61
rlabel metal2 32798 6953 32798 6953 0 net62
rlabel via2 39054 8347 39054 8347 0 net63
rlabel metal2 36018 6409 36018 6409 0 net64
rlabel metal2 37306 6936 37306 6936 0 net65
rlabel metal2 15318 4828 15318 4828 0 net66
rlabel via2 13386 5797 13386 5797 0 net67
rlabel metal2 13386 4964 13386 4964 0 net68
rlabel metal1 38042 2448 38042 2448 0 net69
rlabel metal2 2162 7582 2162 7582 0 net7
rlabel metal2 20930 6188 20930 6188 0 net70
rlabel metal1 20608 5882 20608 5882 0 net71
rlabel metal1 38824 2414 38824 2414 0 net72
rlabel metal1 37444 3366 37444 3366 0 net73
rlabel metal2 17158 3264 17158 3264 0 net74
rlabel metal1 39882 2210 39882 2210 0 net75
rlabel metal3 17020 3400 17020 3400 0 net76
rlabel via2 39238 3043 39238 3043 0 net77
rlabel metal2 38870 4063 38870 4063 0 net78
rlabel metal2 32614 8874 32614 8874 0 net79
rlabel metal2 2714 9044 2714 9044 0 net8
rlabel metal2 36018 5219 36018 5219 0 net80
rlabel metal1 32706 6630 32706 6630 0 net81
rlabel metal1 35144 7242 35144 7242 0 net82
rlabel metal1 35328 7514 35328 7514 0 net83
rlabel metal1 35512 6154 35512 6154 0 net84
rlabel metal1 36432 5882 36432 5882 0 net85
rlabel metal2 36938 7140 36938 7140 0 net86
rlabel metal1 37720 5338 37720 5338 0 net87
rlabel metal1 38272 5338 38272 5338 0 net88
rlabel metal1 37904 4794 37904 4794 0 net89
rlabel metal1 4002 7412 4002 7412 0 net9
rlabel metal1 32706 8500 32706 8500 0 net90
rlabel metal1 32660 4454 32660 4454 0 net91
rlabel metal1 32476 4794 32476 4794 0 net92
rlabel metal1 33166 5814 33166 5814 0 net93
rlabel metal1 33810 6630 33810 6630 0 net94
rlabel metal1 32430 5338 32430 5338 0 net95
rlabel metal2 33442 5780 33442 5780 0 net96
rlabel metal1 35650 3706 35650 3706 0 net97
rlabel metal2 33810 8738 33810 8738 0 net98
rlabel via2 2070 2397 2070 2397 0 net99
<< properties >>
string FIXED_BBOX 0 0 41000 11250
<< end >>
