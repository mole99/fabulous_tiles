VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO E_IO
  CLASS BLOCK ;
  FOREIGN E_IO ;
  ORIGIN 0.000 0.000 ;
  SIZE 59.200 BY 236.800 ;
  PIN A_I_top
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 58.750 9.460 59.200 9.860 ;
    END
  END A_I_top
  PIN A_O_top
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.314600 ;
    PORT
      LAYER Metal2 ;
        RECT 58.750 4.420 59.200 4.820 ;
    END
  END A_O_top
  PIN A_T_top
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 58.750 14.500 59.200 14.900 ;
    END
  END A_T_top
  PIN A_config_C_bit0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 58.750 34.660 59.200 35.060 ;
    END
  END A_config_C_bit0
  PIN A_config_C_bit1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 58.750 39.700 59.200 40.100 ;
    END
  END A_config_C_bit1
  PIN A_config_C_bit2
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 58.750 44.740 59.200 45.140 ;
    END
  END A_config_C_bit2
  PIN A_config_C_bit3
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 58.750 49.780 59.200 50.180 ;
    END
  END A_config_C_bit3
  PIN B_I_top
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 58.750 24.580 59.200 24.980 ;
    END
  END B_I_top
  PIN B_O_top
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.314600 ;
    PORT
      LAYER Metal2 ;
        RECT 58.750 19.540 59.200 19.940 ;
    END
  END B_O_top
  PIN B_T_top
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 58.750 29.620 59.200 30.020 ;
    END
  END B_T_top
  PIN B_config_C_bit0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 58.750 54.820 59.200 55.220 ;
    END
  END B_config_C_bit0
  PIN B_config_C_bit1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 58.750 59.860 59.200 60.260 ;
    END
  END B_config_C_bit1
  PIN B_config_C_bit2
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 58.750 64.900 59.200 65.300 ;
    END
  END B_config_C_bit2
  PIN B_config_C_bit3
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 58.750 69.940 59.200 70.340 ;
    END
  END B_config_C_bit3
  PIN E1END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 91.780 0.450 92.180 ;
    END
  END E1END[0]
  PIN E1END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213200 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 93.460 0.450 93.860 ;
    END
  END E1END[1]
  PIN E1END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213200 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 95.140 0.450 95.540 ;
    END
  END E1END[2]
  PIN E1END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213200 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 96.820 0.450 97.220 ;
    END
  END E1END[3]
  PIN E2END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213200 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 111.940 0.450 112.340 ;
    END
  END E2END[0]
  PIN E2END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213200 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 113.620 0.450 114.020 ;
    END
  END E2END[1]
  PIN E2END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213200 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 115.300 0.450 115.700 ;
    END
  END E2END[2]
  PIN E2END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213200 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 116.980 0.450 117.380 ;
    END
  END E2END[3]
  PIN E2END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213200 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 118.660 0.450 119.060 ;
    END
  END E2END[4]
  PIN E2END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213200 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 120.340 0.450 120.740 ;
    END
  END E2END[5]
  PIN E2END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213200 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 122.020 0.450 122.420 ;
    END
  END E2END[6]
  PIN E2END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213200 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 123.700 0.450 124.100 ;
    END
  END E2END[7]
  PIN E2MID[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213200 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 98.500 0.450 98.900 ;
    END
  END E2MID[0]
  PIN E2MID[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213200 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 100.180 0.450 100.580 ;
    END
  END E2MID[1]
  PIN E2MID[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213200 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 101.860 0.450 102.260 ;
    END
  END E2MID[2]
  PIN E2MID[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213200 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 103.540 0.450 103.940 ;
    END
  END E2MID[3]
  PIN E2MID[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213200 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 105.220 0.450 105.620 ;
    END
  END E2MID[4]
  PIN E2MID[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213200 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 106.900 0.450 107.300 ;
    END
  END E2MID[5]
  PIN E2MID[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213200 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 108.580 0.450 108.980 ;
    END
  END E2MID[6]
  PIN E2MID[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213200 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 110.260 0.450 110.660 ;
    END
  END E2MID[7]
  PIN E6END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213200 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 152.260 0.450 152.660 ;
    END
  END E6END[0]
  PIN E6END[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 169.060 0.450 169.460 ;
    END
  END E6END[10]
  PIN E6END[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 170.740 0.450 171.140 ;
    END
  END E6END[11]
  PIN E6END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.314600 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 153.940 0.450 154.340 ;
    END
  END E6END[1]
  PIN E6END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213200 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 155.620 0.450 156.020 ;
    END
  END E6END[2]
  PIN E6END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213200 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 157.300 0.450 157.700 ;
    END
  END E6END[3]
  PIN E6END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213200 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 158.980 0.450 159.380 ;
    END
  END E6END[4]
  PIN E6END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213200 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 160.660 0.450 161.060 ;
    END
  END E6END[5]
  PIN E6END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213200 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 162.340 0.450 162.740 ;
    END
  END E6END[6]
  PIN E6END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213200 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 164.020 0.450 164.420 ;
    END
  END E6END[7]
  PIN E6END[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.314600 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 165.700 0.450 166.100 ;
    END
  END E6END[8]
  PIN E6END[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213200 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 167.380 0.450 167.780 ;
    END
  END E6END[9]
  PIN EE4END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213200 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 125.380 0.450 125.780 ;
    END
  END EE4END[0]
  PIN EE4END[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213200 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 142.180 0.450 142.580 ;
    END
  END EE4END[10]
  PIN EE4END[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213200 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 143.860 0.450 144.260 ;
    END
  END EE4END[11]
  PIN EE4END[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 145.540 0.450 145.940 ;
    END
  END EE4END[12]
  PIN EE4END[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 147.220 0.450 147.620 ;
    END
  END EE4END[13]
  PIN EE4END[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 148.900 0.450 149.300 ;
    END
  END EE4END[14]
  PIN EE4END[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 150.580 0.450 150.980 ;
    END
  END EE4END[15]
  PIN EE4END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213200 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 127.060 0.450 127.460 ;
    END
  END EE4END[1]
  PIN EE4END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 128.740 0.450 129.140 ;
    END
  END EE4END[2]
  PIN EE4END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213200 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 130.420 0.450 130.820 ;
    END
  END EE4END[3]
  PIN EE4END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 132.100 0.450 132.500 ;
    END
  END EE4END[4]
  PIN EE4END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 133.780 0.450 134.180 ;
    END
  END EE4END[5]
  PIN EE4END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213200 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 135.460 0.450 135.860 ;
    END
  END EE4END[6]
  PIN EE4END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 137.140 0.450 137.540 ;
    END
  END EE4END[7]
  PIN EE4END[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213200 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 138.820 0.450 139.220 ;
    END
  END EE4END[8]
  PIN EE4END[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213200 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 140.500 0.450 140.900 ;
    END
  END EE4END[9]
  PIN FrameData[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 172.420 0.450 172.820 ;
    END
  END FrameData[0]
  PIN FrameData[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 189.220 0.450 189.620 ;
    END
  END FrameData[10]
  PIN FrameData[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 190.900 0.450 191.300 ;
    END
  END FrameData[11]
  PIN FrameData[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 192.580 0.450 192.980 ;
    END
  END FrameData[12]
  PIN FrameData[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 194.260 0.450 194.660 ;
    END
  END FrameData[13]
  PIN FrameData[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.314600 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 195.940 0.450 196.340 ;
    END
  END FrameData[14]
  PIN FrameData[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.314600 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 197.620 0.450 198.020 ;
    END
  END FrameData[15]
  PIN FrameData[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.314600 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 199.300 0.450 199.700 ;
    END
  END FrameData[16]
  PIN FrameData[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.314600 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 200.980 0.450 201.380 ;
    END
  END FrameData[17]
  PIN FrameData[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213200 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 202.660 0.450 203.060 ;
    END
  END FrameData[18]
  PIN FrameData[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.314600 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 204.340 0.450 204.740 ;
    END
  END FrameData[19]
  PIN FrameData[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 174.100 0.450 174.500 ;
    END
  END FrameData[1]
  PIN FrameData[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.314600 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 206.020 0.450 206.420 ;
    END
  END FrameData[20]
  PIN FrameData[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213200 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 207.700 0.450 208.100 ;
    END
  END FrameData[21]
  PIN FrameData[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.314600 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 209.380 0.450 209.780 ;
    END
  END FrameData[22]
  PIN FrameData[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.314600 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 211.060 0.450 211.460 ;
    END
  END FrameData[23]
  PIN FrameData[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.314600 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 212.740 0.450 213.140 ;
    END
  END FrameData[24]
  PIN FrameData[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.314600 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 214.420 0.450 214.820 ;
    END
  END FrameData[25]
  PIN FrameData[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213200 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 216.100 0.450 216.500 ;
    END
  END FrameData[26]
  PIN FrameData[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213200 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 217.780 0.450 218.180 ;
    END
  END FrameData[27]
  PIN FrameData[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 219.460 0.450 219.860 ;
    END
  END FrameData[28]
  PIN FrameData[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 221.140 0.450 221.540 ;
    END
  END FrameData[29]
  PIN FrameData[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213200 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 175.780 0.450 176.180 ;
    END
  END FrameData[2]
  PIN FrameData[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213200 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 222.820 0.450 223.220 ;
    END
  END FrameData[30]
  PIN FrameData[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213200 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 224.500 0.450 224.900 ;
    END
  END FrameData[31]
  PIN FrameData[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213200 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 177.460 0.450 177.860 ;
    END
  END FrameData[3]
  PIN FrameData[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213200 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 179.140 0.450 179.540 ;
    END
  END FrameData[4]
  PIN FrameData[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213200 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 180.820 0.450 181.220 ;
    END
  END FrameData[5]
  PIN FrameData[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213200 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 182.500 0.450 182.900 ;
    END
  END FrameData[6]
  PIN FrameData[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.314600 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 184.180 0.450 184.580 ;
    END
  END FrameData[7]
  PIN FrameData[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213200 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 185.860 0.450 186.260 ;
    END
  END FrameData[8]
  PIN FrameData[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213200 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 187.540 0.450 187.940 ;
    END
  END FrameData[9]
  PIN FrameData_O[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 58.750 74.980 59.200 75.380 ;
    END
  END FrameData_O[0]
  PIN FrameData_O[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 58.750 125.380 59.200 125.780 ;
    END
  END FrameData_O[10]
  PIN FrameData_O[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 58.750 130.420 59.200 130.820 ;
    END
  END FrameData_O[11]
  PIN FrameData_O[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 58.750 135.460 59.200 135.860 ;
    END
  END FrameData_O[12]
  PIN FrameData_O[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 58.750 140.500 59.200 140.900 ;
    END
  END FrameData_O[13]
  PIN FrameData_O[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 58.750 145.540 59.200 145.940 ;
    END
  END FrameData_O[14]
  PIN FrameData_O[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 58.750 150.580 59.200 150.980 ;
    END
  END FrameData_O[15]
  PIN FrameData_O[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 58.750 155.620 59.200 156.020 ;
    END
  END FrameData_O[16]
  PIN FrameData_O[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 58.750 160.660 59.200 161.060 ;
    END
  END FrameData_O[17]
  PIN FrameData_O[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 58.750 165.700 59.200 166.100 ;
    END
  END FrameData_O[18]
  PIN FrameData_O[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 58.750 170.740 59.200 171.140 ;
    END
  END FrameData_O[19]
  PIN FrameData_O[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 58.750 80.020 59.200 80.420 ;
    END
  END FrameData_O[1]
  PIN FrameData_O[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 58.750 175.780 59.200 176.180 ;
    END
  END FrameData_O[20]
  PIN FrameData_O[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 58.750 180.820 59.200 181.220 ;
    END
  END FrameData_O[21]
  PIN FrameData_O[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 58.750 185.860 59.200 186.260 ;
    END
  END FrameData_O[22]
  PIN FrameData_O[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 58.750 190.900 59.200 191.300 ;
    END
  END FrameData_O[23]
  PIN FrameData_O[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 58.750 195.940 59.200 196.340 ;
    END
  END FrameData_O[24]
  PIN FrameData_O[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 58.750 200.980 59.200 201.380 ;
    END
  END FrameData_O[25]
  PIN FrameData_O[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 58.750 206.020 59.200 206.420 ;
    END
  END FrameData_O[26]
  PIN FrameData_O[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 58.750 211.060 59.200 211.460 ;
    END
  END FrameData_O[27]
  PIN FrameData_O[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 58.750 216.100 59.200 216.500 ;
    END
  END FrameData_O[28]
  PIN FrameData_O[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 58.750 221.140 59.200 221.540 ;
    END
  END FrameData_O[29]
  PIN FrameData_O[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 58.750 85.060 59.200 85.460 ;
    END
  END FrameData_O[2]
  PIN FrameData_O[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 58.750 226.180 59.200 226.580 ;
    END
  END FrameData_O[30]
  PIN FrameData_O[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 58.750 231.220 59.200 231.620 ;
    END
  END FrameData_O[31]
  PIN FrameData_O[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 58.750 90.100 59.200 90.500 ;
    END
  END FrameData_O[3]
  PIN FrameData_O[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 58.750 95.140 59.200 95.540 ;
    END
  END FrameData_O[4]
  PIN FrameData_O[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 58.750 100.180 59.200 100.580 ;
    END
  END FrameData_O[5]
  PIN FrameData_O[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 58.750 105.220 59.200 105.620 ;
    END
  END FrameData_O[6]
  PIN FrameData_O[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 58.750 110.260 59.200 110.660 ;
    END
  END FrameData_O[7]
  PIN FrameData_O[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 58.750 115.300 59.200 115.700 ;
    END
  END FrameData_O[8]
  PIN FrameData_O[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 58.750 120.340 59.200 120.740 ;
    END
  END FrameData_O[9]
  PIN FrameStrobe[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426400 ;
    PORT
      LAYER Metal3 ;
        RECT 11.800 0.000 12.200 0.400 ;
    END
  END FrameStrobe[0]
  PIN FrameStrobe[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 6.264700 ;
    ANTENNADIFFAREA 20.153999 ;
    PORT
      LAYER Metal3 ;
        RECT 31.000 0.000 31.400 0.400 ;
    END
  END FrameStrobe[10]
  PIN FrameStrobe[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 5.047900 ;
    ANTENNADIFFAREA 16.123199 ;
    PORT
      LAYER Metal3 ;
        RECT 32.920 0.000 33.320 0.400 ;
    END
  END FrameStrobe[11]
  PIN FrameStrobe[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 5.047900 ;
    ANTENNADIFFAREA 16.123199 ;
    PORT
      LAYER Metal3 ;
        RECT 34.840 0.000 35.240 0.400 ;
    END
  END FrameStrobe[12]
  PIN FrameStrobe[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 36.760 0.000 37.160 0.400 ;
    END
  END FrameStrobe[13]
  PIN FrameStrobe[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.831100 ;
    ANTENNADIFFAREA 12.092400 ;
    PORT
      LAYER Metal3 ;
        RECT 38.680 0.000 39.080 0.400 ;
    END
  END FrameStrobe[14]
  PIN FrameStrobe[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 40.600 0.000 41.000 0.400 ;
    END
  END FrameStrobe[15]
  PIN FrameStrobe[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 5.656300 ;
    ANTENNADIFFAREA 18.138599 ;
    PORT
      LAYER Metal3 ;
        RECT 42.520 0.000 42.920 0.400 ;
    END
  END FrameStrobe[16]
  PIN FrameStrobe[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.005900 ;
    ANTENNADIFFAREA 6.046200 ;
    PORT
      LAYER Metal3 ;
        RECT 44.440 0.000 44.840 0.400 ;
    END
  END FrameStrobe[17]
  PIN FrameStrobe[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 6.264700 ;
    ANTENNADIFFAREA 20.153999 ;
    PORT
      LAYER Metal3 ;
        RECT 46.360 0.000 46.760 0.400 ;
    END
  END FrameStrobe[18]
  PIN FrameStrobe[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 6.264700 ;
    ANTENNADIFFAREA 20.153999 ;
    PORT
      LAYER Metal3 ;
        RECT 48.280 0.000 48.680 0.400 ;
    END
  END FrameStrobe[19]
  PIN FrameStrobe[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.639600 ;
    PORT
      LAYER Metal3 ;
        RECT 13.720 0.000 14.120 0.400 ;
    END
  END FrameStrobe[1]
  PIN FrameStrobe[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.639600 ;
    PORT
      LAYER Metal3 ;
        RECT 15.640 0.000 16.040 0.400 ;
    END
  END FrameStrobe[2]
  PIN FrameStrobe[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 5.688800 ;
    ANTENNADIFFAREA 18.138599 ;
    PORT
      LAYER Metal3 ;
        RECT 17.560 0.000 17.960 0.400 ;
    END
  END FrameStrobe[3]
  PIN FrameStrobe[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 6.264700 ;
    ANTENNADIFFAREA 20.153999 ;
    PORT
      LAYER Metal3 ;
        RECT 19.480 0.000 19.880 0.400 ;
    END
  END FrameStrobe[4]
  PIN FrameStrobe[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 21.400 0.000 21.800 0.400 ;
    END
  END FrameStrobe[5]
  PIN FrameStrobe[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 5.656300 ;
    ANTENNADIFFAREA 18.138599 ;
    PORT
      LAYER Metal3 ;
        RECT 23.320 0.000 23.720 0.400 ;
    END
  END FrameStrobe[6]
  PIN FrameStrobe[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 4.439500 ;
    ANTENNADIFFAREA 14.107800 ;
    PORT
      LAYER Metal3 ;
        RECT 25.240 0.000 25.640 0.400 ;
    END
  END FrameStrobe[7]
  PIN FrameStrobe[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.831100 ;
    ANTENNADIFFAREA 12.092400 ;
    PORT
      LAYER Metal3 ;
        RECT 27.160 0.000 27.560 0.400 ;
    END
  END FrameStrobe[8]
  PIN FrameStrobe[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 5.656300 ;
    ANTENNADIFFAREA 18.138599 ;
    PORT
      LAYER Metal3 ;
        RECT 29.080 0.000 29.480 0.400 ;
    END
  END FrameStrobe[9]
  PIN FrameStrobe_O[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 11.800 236.400 12.200 236.800 ;
    END
  END FrameStrobe_O[0]
  PIN FrameStrobe_O[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 31.000 236.400 31.400 236.800 ;
    END
  END FrameStrobe_O[10]
  PIN FrameStrobe_O[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 32.920 236.400 33.320 236.800 ;
    END
  END FrameStrobe_O[11]
  PIN FrameStrobe_O[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 34.840 236.400 35.240 236.800 ;
    END
  END FrameStrobe_O[12]
  PIN FrameStrobe_O[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 36.760 236.400 37.160 236.800 ;
    END
  END FrameStrobe_O[13]
  PIN FrameStrobe_O[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 38.680 236.400 39.080 236.800 ;
    END
  END FrameStrobe_O[14]
  PIN FrameStrobe_O[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 40.600 236.400 41.000 236.800 ;
    END
  END FrameStrobe_O[15]
  PIN FrameStrobe_O[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 42.520 236.400 42.920 236.800 ;
    END
  END FrameStrobe_O[16]
  PIN FrameStrobe_O[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 44.440 236.400 44.840 236.800 ;
    END
  END FrameStrobe_O[17]
  PIN FrameStrobe_O[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 46.360 236.400 46.760 236.800 ;
    END
  END FrameStrobe_O[18]
  PIN FrameStrobe_O[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 48.280 236.400 48.680 236.800 ;
    END
  END FrameStrobe_O[19]
  PIN FrameStrobe_O[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 13.720 236.400 14.120 236.800 ;
    END
  END FrameStrobe_O[1]
  PIN FrameStrobe_O[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 15.640 236.400 16.040 236.800 ;
    END
  END FrameStrobe_O[2]
  PIN FrameStrobe_O[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 17.560 236.400 17.960 236.800 ;
    END
  END FrameStrobe_O[3]
  PIN FrameStrobe_O[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 19.480 236.400 19.880 236.800 ;
    END
  END FrameStrobe_O[4]
  PIN FrameStrobe_O[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 21.400 236.400 21.800 236.800 ;
    END
  END FrameStrobe_O[5]
  PIN FrameStrobe_O[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 23.320 236.400 23.720 236.800 ;
    END
  END FrameStrobe_O[6]
  PIN FrameStrobe_O[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 25.240 236.400 25.640 236.800 ;
    END
  END FrameStrobe_O[7]
  PIN FrameStrobe_O[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 27.160 236.400 27.560 236.800 ;
    END
  END FrameStrobe_O[8]
  PIN FrameStrobe_O[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 29.080 236.400 29.480 236.800 ;
    END
  END FrameStrobe_O[9]
  PIN UserCLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.633100 ;
    PORT
      LAYER Metal3 ;
        RECT 9.880 0.000 10.280 0.400 ;
    END
  END UserCLK
  PIN UserCLKo
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 9.880 236.400 10.280 236.800 ;
    END
  END UserCLKo
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal5 ;
        RECT 24.460 0.000 26.660 236.800 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal5 ;
        RECT 18.260 0.000 20.460 236.800 ;
    END
  END VPWR
  PIN W1BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 11.140 0.450 11.540 ;
    END
  END W1BEG[0]
  PIN W1BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 12.820 0.450 13.220 ;
    END
  END W1BEG[1]
  PIN W1BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 14.500 0.450 14.900 ;
    END
  END W1BEG[2]
  PIN W1BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 16.180 0.450 16.580 ;
    END
  END W1BEG[3]
  PIN W2BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 17.860 0.450 18.260 ;
    END
  END W2BEG[0]
  PIN W2BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 19.540 0.450 19.940 ;
    END
  END W2BEG[1]
  PIN W2BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 21.220 0.450 21.620 ;
    END
  END W2BEG[2]
  PIN W2BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 22.900 0.450 23.300 ;
    END
  END W2BEG[3]
  PIN W2BEG[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 24.580 0.450 24.980 ;
    END
  END W2BEG[4]
  PIN W2BEG[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 26.260 0.450 26.660 ;
    END
  END W2BEG[5]
  PIN W2BEG[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 27.940 0.450 28.340 ;
    END
  END W2BEG[6]
  PIN W2BEG[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 29.620 0.450 30.020 ;
    END
  END W2BEG[7]
  PIN W2BEGb[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 31.300 0.450 31.700 ;
    END
  END W2BEGb[0]
  PIN W2BEGb[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 32.980 0.450 33.380 ;
    END
  END W2BEGb[1]
  PIN W2BEGb[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 34.660 0.450 35.060 ;
    END
  END W2BEGb[2]
  PIN W2BEGb[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 36.340 0.450 36.740 ;
    END
  END W2BEGb[3]
  PIN W2BEGb[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 38.020 0.450 38.420 ;
    END
  END W2BEGb[4]
  PIN W2BEGb[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 39.700 0.450 40.100 ;
    END
  END W2BEGb[5]
  PIN W2BEGb[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 41.380 0.450 41.780 ;
    END
  END W2BEGb[6]
  PIN W2BEGb[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 43.060 0.450 43.460 ;
    END
  END W2BEGb[7]
  PIN W6BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 71.620 0.450 72.020 ;
    END
  END W6BEG[0]
  PIN W6BEG[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 88.420 0.450 88.820 ;
    END
  END W6BEG[10]
  PIN W6BEG[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 90.100 0.450 90.500 ;
    END
  END W6BEG[11]
  PIN W6BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 73.300 0.450 73.700 ;
    END
  END W6BEG[1]
  PIN W6BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 74.980 0.450 75.380 ;
    END
  END W6BEG[2]
  PIN W6BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 76.660 0.450 77.060 ;
    END
  END W6BEG[3]
  PIN W6BEG[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 78.340 0.450 78.740 ;
    END
  END W6BEG[4]
  PIN W6BEG[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 80.020 0.450 80.420 ;
    END
  END W6BEG[5]
  PIN W6BEG[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 81.700 0.450 82.100 ;
    END
  END W6BEG[6]
  PIN W6BEG[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 83.380 0.450 83.780 ;
    END
  END W6BEG[7]
  PIN W6BEG[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 85.060 0.450 85.460 ;
    END
  END W6BEG[8]
  PIN W6BEG[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 86.740 0.450 87.140 ;
    END
  END W6BEG[9]
  PIN WW4BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 44.740 0.450 45.140 ;
    END
  END WW4BEG[0]
  PIN WW4BEG[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 61.540 0.450 61.940 ;
    END
  END WW4BEG[10]
  PIN WW4BEG[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 63.220 0.450 63.620 ;
    END
  END WW4BEG[11]
  PIN WW4BEG[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 64.900 0.450 65.300 ;
    END
  END WW4BEG[12]
  PIN WW4BEG[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 66.580 0.450 66.980 ;
    END
  END WW4BEG[13]
  PIN WW4BEG[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 68.260 0.450 68.660 ;
    END
  END WW4BEG[14]
  PIN WW4BEG[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 69.940 0.450 70.340 ;
    END
  END WW4BEG[15]
  PIN WW4BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 46.420 0.450 46.820 ;
    END
  END WW4BEG[1]
  PIN WW4BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 48.100 0.450 48.500 ;
    END
  END WW4BEG[2]
  PIN WW4BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 49.780 0.450 50.180 ;
    END
  END WW4BEG[3]
  PIN WW4BEG[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 51.460 0.450 51.860 ;
    END
  END WW4BEG[4]
  PIN WW4BEG[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 53.140 0.450 53.540 ;
    END
  END WW4BEG[5]
  PIN WW4BEG[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 54.820 0.450 55.220 ;
    END
  END WW4BEG[6]
  PIN WW4BEG[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 56.500 0.450 56.900 ;
    END
  END WW4BEG[7]
  PIN WW4BEG[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 58.180 0.450 58.580 ;
    END
  END WW4BEG[8]
  PIN WW4BEG[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 59.860 0.450 60.260 ;
    END
  END WW4BEG[9]
  OBS
      LAYER GatPoly ;
        RECT 5.760 7.410 53.280 226.950 ;
      LAYER Metal1 ;
        RECT 5.760 7.340 53.280 227.020 ;
      LAYER Metal2 ;
        RECT 0.335 231.010 58.540 231.520 ;
        RECT 0.335 226.790 59.185 231.010 ;
        RECT 0.335 225.970 58.540 226.790 ;
        RECT 0.335 225.110 59.185 225.970 ;
        RECT 0.660 224.290 59.185 225.110 ;
        RECT 0.335 223.430 59.185 224.290 ;
        RECT 0.660 222.610 59.185 223.430 ;
        RECT 0.335 221.750 59.185 222.610 ;
        RECT 0.660 220.930 58.540 221.750 ;
        RECT 0.335 220.070 59.185 220.930 ;
        RECT 0.660 219.250 59.185 220.070 ;
        RECT 0.335 218.390 59.185 219.250 ;
        RECT 0.660 217.570 59.185 218.390 ;
        RECT 0.335 216.710 59.185 217.570 ;
        RECT 0.660 215.890 58.540 216.710 ;
        RECT 0.335 215.030 59.185 215.890 ;
        RECT 0.660 214.210 59.185 215.030 ;
        RECT 0.335 213.350 59.185 214.210 ;
        RECT 0.660 212.530 59.185 213.350 ;
        RECT 0.335 211.670 59.185 212.530 ;
        RECT 0.660 210.850 58.540 211.670 ;
        RECT 0.335 209.990 59.185 210.850 ;
        RECT 0.660 209.170 59.185 209.990 ;
        RECT 0.335 208.310 59.185 209.170 ;
        RECT 0.660 207.490 59.185 208.310 ;
        RECT 0.335 206.630 59.185 207.490 ;
        RECT 0.660 205.810 58.540 206.630 ;
        RECT 0.335 204.950 59.185 205.810 ;
        RECT 0.660 204.130 59.185 204.950 ;
        RECT 0.335 203.270 59.185 204.130 ;
        RECT 0.660 202.450 59.185 203.270 ;
        RECT 0.335 201.590 59.185 202.450 ;
        RECT 0.660 200.770 58.540 201.590 ;
        RECT 0.335 199.910 59.185 200.770 ;
        RECT 0.660 199.090 59.185 199.910 ;
        RECT 0.335 198.230 59.185 199.090 ;
        RECT 0.660 197.410 59.185 198.230 ;
        RECT 0.335 196.550 59.185 197.410 ;
        RECT 0.660 195.730 58.540 196.550 ;
        RECT 0.335 194.870 59.185 195.730 ;
        RECT 0.660 194.050 59.185 194.870 ;
        RECT 0.335 193.190 59.185 194.050 ;
        RECT 0.660 192.370 59.185 193.190 ;
        RECT 0.335 191.510 59.185 192.370 ;
        RECT 0.660 190.690 58.540 191.510 ;
        RECT 0.335 189.830 59.185 190.690 ;
        RECT 0.660 189.010 59.185 189.830 ;
        RECT 0.335 188.150 59.185 189.010 ;
        RECT 0.660 187.330 59.185 188.150 ;
        RECT 0.335 186.470 59.185 187.330 ;
        RECT 0.660 185.650 58.540 186.470 ;
        RECT 0.335 184.790 59.185 185.650 ;
        RECT 0.660 183.970 59.185 184.790 ;
        RECT 0.335 183.110 59.185 183.970 ;
        RECT 0.660 182.290 59.185 183.110 ;
        RECT 0.335 181.430 59.185 182.290 ;
        RECT 0.660 180.610 58.540 181.430 ;
        RECT 0.335 179.750 59.185 180.610 ;
        RECT 0.660 178.930 59.185 179.750 ;
        RECT 0.335 178.070 59.185 178.930 ;
        RECT 0.660 177.250 59.185 178.070 ;
        RECT 0.335 176.390 59.185 177.250 ;
        RECT 0.660 175.570 58.540 176.390 ;
        RECT 0.335 174.710 59.185 175.570 ;
        RECT 0.660 173.890 59.185 174.710 ;
        RECT 0.335 173.030 59.185 173.890 ;
        RECT 0.660 172.210 59.185 173.030 ;
        RECT 0.335 171.350 59.185 172.210 ;
        RECT 0.660 170.530 58.540 171.350 ;
        RECT 0.335 169.670 59.185 170.530 ;
        RECT 0.660 168.850 59.185 169.670 ;
        RECT 0.335 167.990 59.185 168.850 ;
        RECT 0.660 167.170 59.185 167.990 ;
        RECT 0.335 166.310 59.185 167.170 ;
        RECT 0.660 165.490 58.540 166.310 ;
        RECT 0.335 164.630 59.185 165.490 ;
        RECT 0.660 163.810 59.185 164.630 ;
        RECT 0.335 162.950 59.185 163.810 ;
        RECT 0.660 162.130 59.185 162.950 ;
        RECT 0.335 161.270 59.185 162.130 ;
        RECT 0.660 160.450 58.540 161.270 ;
        RECT 0.335 159.590 59.185 160.450 ;
        RECT 0.660 158.770 59.185 159.590 ;
        RECT 0.335 157.910 59.185 158.770 ;
        RECT 0.660 157.090 59.185 157.910 ;
        RECT 0.335 156.230 59.185 157.090 ;
        RECT 0.660 155.410 58.540 156.230 ;
        RECT 0.335 154.550 59.185 155.410 ;
        RECT 0.660 153.730 59.185 154.550 ;
        RECT 0.335 152.870 59.185 153.730 ;
        RECT 0.660 152.050 59.185 152.870 ;
        RECT 0.335 151.190 59.185 152.050 ;
        RECT 0.660 150.370 58.540 151.190 ;
        RECT 0.335 149.510 59.185 150.370 ;
        RECT 0.660 148.690 59.185 149.510 ;
        RECT 0.335 147.830 59.185 148.690 ;
        RECT 0.660 147.010 59.185 147.830 ;
        RECT 0.335 146.150 59.185 147.010 ;
        RECT 0.660 145.330 58.540 146.150 ;
        RECT 0.335 144.470 59.185 145.330 ;
        RECT 0.660 143.650 59.185 144.470 ;
        RECT 0.335 142.790 59.185 143.650 ;
        RECT 0.660 141.970 59.185 142.790 ;
        RECT 0.335 141.110 59.185 141.970 ;
        RECT 0.660 140.290 58.540 141.110 ;
        RECT 0.335 139.430 59.185 140.290 ;
        RECT 0.660 138.610 59.185 139.430 ;
        RECT 0.335 137.750 59.185 138.610 ;
        RECT 0.660 136.930 59.185 137.750 ;
        RECT 0.335 136.070 59.185 136.930 ;
        RECT 0.660 135.250 58.540 136.070 ;
        RECT 0.335 134.390 59.185 135.250 ;
        RECT 0.660 133.570 59.185 134.390 ;
        RECT 0.335 132.710 59.185 133.570 ;
        RECT 0.660 131.890 59.185 132.710 ;
        RECT 0.335 131.030 59.185 131.890 ;
        RECT 0.660 130.210 58.540 131.030 ;
        RECT 0.335 129.350 59.185 130.210 ;
        RECT 0.660 128.530 59.185 129.350 ;
        RECT 0.335 127.670 59.185 128.530 ;
        RECT 0.660 126.850 59.185 127.670 ;
        RECT 0.335 125.990 59.185 126.850 ;
        RECT 0.660 125.170 58.540 125.990 ;
        RECT 0.335 124.310 59.185 125.170 ;
        RECT 0.660 123.490 59.185 124.310 ;
        RECT 0.335 122.630 59.185 123.490 ;
        RECT 0.660 121.810 59.185 122.630 ;
        RECT 0.335 120.950 59.185 121.810 ;
        RECT 0.660 120.130 58.540 120.950 ;
        RECT 0.335 119.270 59.185 120.130 ;
        RECT 0.660 118.450 59.185 119.270 ;
        RECT 0.335 117.590 59.185 118.450 ;
        RECT 0.660 116.770 59.185 117.590 ;
        RECT 0.335 115.910 59.185 116.770 ;
        RECT 0.660 115.090 58.540 115.910 ;
        RECT 0.335 114.230 59.185 115.090 ;
        RECT 0.660 113.410 59.185 114.230 ;
        RECT 0.335 112.550 59.185 113.410 ;
        RECT 0.660 111.730 59.185 112.550 ;
        RECT 0.335 110.870 59.185 111.730 ;
        RECT 0.660 110.050 58.540 110.870 ;
        RECT 0.335 109.190 59.185 110.050 ;
        RECT 0.660 108.370 59.185 109.190 ;
        RECT 0.335 107.510 59.185 108.370 ;
        RECT 0.660 106.690 59.185 107.510 ;
        RECT 0.335 105.830 59.185 106.690 ;
        RECT 0.660 105.010 58.540 105.830 ;
        RECT 0.335 104.150 59.185 105.010 ;
        RECT 0.660 103.330 59.185 104.150 ;
        RECT 0.335 102.470 59.185 103.330 ;
        RECT 0.660 101.650 59.185 102.470 ;
        RECT 0.335 100.790 59.185 101.650 ;
        RECT 0.660 99.970 58.540 100.790 ;
        RECT 0.335 99.110 59.185 99.970 ;
        RECT 0.660 98.290 59.185 99.110 ;
        RECT 0.335 97.430 59.185 98.290 ;
        RECT 0.660 96.610 59.185 97.430 ;
        RECT 0.335 95.750 59.185 96.610 ;
        RECT 0.660 94.930 58.540 95.750 ;
        RECT 0.335 94.070 59.185 94.930 ;
        RECT 0.660 93.250 59.185 94.070 ;
        RECT 0.335 92.390 59.185 93.250 ;
        RECT 0.660 91.570 59.185 92.390 ;
        RECT 0.335 90.710 59.185 91.570 ;
        RECT 0.660 89.890 58.540 90.710 ;
        RECT 0.335 89.030 59.185 89.890 ;
        RECT 0.660 88.210 59.185 89.030 ;
        RECT 0.335 87.350 59.185 88.210 ;
        RECT 0.660 86.530 59.185 87.350 ;
        RECT 0.335 85.670 59.185 86.530 ;
        RECT 0.660 84.850 58.540 85.670 ;
        RECT 0.335 83.990 59.185 84.850 ;
        RECT 0.660 83.170 59.185 83.990 ;
        RECT 0.335 82.310 59.185 83.170 ;
        RECT 0.660 81.490 59.185 82.310 ;
        RECT 0.335 80.630 59.185 81.490 ;
        RECT 0.660 79.810 58.540 80.630 ;
        RECT 0.335 78.950 59.185 79.810 ;
        RECT 0.660 78.130 59.185 78.950 ;
        RECT 0.335 77.270 59.185 78.130 ;
        RECT 0.660 76.450 59.185 77.270 ;
        RECT 0.335 75.590 59.185 76.450 ;
        RECT 0.660 74.770 58.540 75.590 ;
        RECT 0.335 73.910 59.185 74.770 ;
        RECT 0.660 73.090 59.185 73.910 ;
        RECT 0.335 72.230 59.185 73.090 ;
        RECT 0.660 71.410 59.185 72.230 ;
        RECT 0.335 70.550 59.185 71.410 ;
        RECT 0.660 69.730 58.540 70.550 ;
        RECT 0.335 68.870 59.185 69.730 ;
        RECT 0.660 68.050 59.185 68.870 ;
        RECT 0.335 67.190 59.185 68.050 ;
        RECT 0.660 66.370 59.185 67.190 ;
        RECT 0.335 65.510 59.185 66.370 ;
        RECT 0.660 64.690 58.540 65.510 ;
        RECT 0.335 63.830 59.185 64.690 ;
        RECT 0.660 63.010 59.185 63.830 ;
        RECT 0.335 62.150 59.185 63.010 ;
        RECT 0.660 61.330 59.185 62.150 ;
        RECT 0.335 60.470 59.185 61.330 ;
        RECT 0.660 59.650 58.540 60.470 ;
        RECT 0.335 58.790 59.185 59.650 ;
        RECT 0.660 57.970 59.185 58.790 ;
        RECT 0.335 57.110 59.185 57.970 ;
        RECT 0.660 56.290 59.185 57.110 ;
        RECT 0.335 55.430 59.185 56.290 ;
        RECT 0.660 54.610 58.540 55.430 ;
        RECT 0.335 53.750 59.185 54.610 ;
        RECT 0.660 52.930 59.185 53.750 ;
        RECT 0.335 52.070 59.185 52.930 ;
        RECT 0.660 51.250 59.185 52.070 ;
        RECT 0.335 50.390 59.185 51.250 ;
        RECT 0.660 49.570 58.540 50.390 ;
        RECT 0.335 48.710 59.185 49.570 ;
        RECT 0.660 47.890 59.185 48.710 ;
        RECT 0.335 47.030 59.185 47.890 ;
        RECT 0.660 46.210 59.185 47.030 ;
        RECT 0.335 45.350 59.185 46.210 ;
        RECT 0.660 44.530 58.540 45.350 ;
        RECT 0.335 43.670 59.185 44.530 ;
        RECT 0.660 42.850 59.185 43.670 ;
        RECT 0.335 41.990 59.185 42.850 ;
        RECT 0.660 41.170 59.185 41.990 ;
        RECT 0.335 40.310 59.185 41.170 ;
        RECT 0.660 39.490 58.540 40.310 ;
        RECT 0.335 38.630 59.185 39.490 ;
        RECT 0.660 37.810 59.185 38.630 ;
        RECT 0.335 36.950 59.185 37.810 ;
        RECT 0.660 36.130 59.185 36.950 ;
        RECT 0.335 35.270 59.185 36.130 ;
        RECT 0.660 34.450 58.540 35.270 ;
        RECT 0.335 33.590 59.185 34.450 ;
        RECT 0.660 32.770 59.185 33.590 ;
        RECT 0.335 31.910 59.185 32.770 ;
        RECT 0.660 31.090 59.185 31.910 ;
        RECT 0.335 30.230 59.185 31.090 ;
        RECT 0.660 29.410 58.540 30.230 ;
        RECT 0.335 28.550 59.185 29.410 ;
        RECT 0.660 27.730 59.185 28.550 ;
        RECT 0.335 26.870 59.185 27.730 ;
        RECT 0.660 26.050 59.185 26.870 ;
        RECT 0.335 25.190 59.185 26.050 ;
        RECT 0.660 24.370 58.540 25.190 ;
        RECT 0.335 23.510 59.185 24.370 ;
        RECT 0.660 22.690 59.185 23.510 ;
        RECT 0.335 21.830 59.185 22.690 ;
        RECT 0.660 21.010 59.185 21.830 ;
        RECT 0.335 20.150 59.185 21.010 ;
        RECT 0.660 19.330 58.540 20.150 ;
        RECT 0.335 18.470 59.185 19.330 ;
        RECT 0.660 17.650 59.185 18.470 ;
        RECT 0.335 16.790 59.185 17.650 ;
        RECT 0.660 15.970 59.185 16.790 ;
        RECT 0.335 15.110 59.185 15.970 ;
        RECT 0.660 14.290 58.540 15.110 ;
        RECT 0.335 13.430 59.185 14.290 ;
        RECT 0.660 12.610 59.185 13.430 ;
        RECT 0.335 11.750 59.185 12.610 ;
        RECT 0.660 10.930 59.185 11.750 ;
        RECT 0.335 10.070 59.185 10.930 ;
        RECT 0.335 9.250 58.540 10.070 ;
        RECT 0.335 5.030 59.185 9.250 ;
        RECT 0.335 4.520 58.540 5.030 ;
      LAYER Metal3 ;
        RECT 0.380 236.190 9.670 236.400 ;
        RECT 10.490 236.190 11.590 236.400 ;
        RECT 12.410 236.190 13.510 236.400 ;
        RECT 14.330 236.190 15.430 236.400 ;
        RECT 16.250 236.190 17.350 236.400 ;
        RECT 18.170 236.190 19.270 236.400 ;
        RECT 20.090 236.190 21.190 236.400 ;
        RECT 22.010 236.190 23.110 236.400 ;
        RECT 23.930 236.190 25.030 236.400 ;
        RECT 25.850 236.190 26.950 236.400 ;
        RECT 27.770 236.190 28.870 236.400 ;
        RECT 29.690 236.190 30.790 236.400 ;
        RECT 31.610 236.190 32.710 236.400 ;
        RECT 33.530 236.190 34.630 236.400 ;
        RECT 35.450 236.190 36.550 236.400 ;
        RECT 37.370 236.190 38.470 236.400 ;
        RECT 39.290 236.190 40.390 236.400 ;
        RECT 41.210 236.190 42.310 236.400 ;
        RECT 43.130 236.190 44.230 236.400 ;
        RECT 45.050 236.190 46.150 236.400 ;
        RECT 46.970 236.190 48.070 236.400 ;
        RECT 48.890 236.190 59.140 236.400 ;
        RECT 0.380 0.610 59.140 236.190 ;
        RECT 0.380 0.320 9.670 0.610 ;
        RECT 10.490 0.320 11.590 0.610 ;
        RECT 12.410 0.320 13.510 0.610 ;
        RECT 14.330 0.320 15.430 0.610 ;
        RECT 16.250 0.320 17.350 0.610 ;
        RECT 18.170 0.320 19.270 0.610 ;
        RECT 20.090 0.320 21.190 0.610 ;
        RECT 22.010 0.320 23.110 0.610 ;
        RECT 23.930 0.320 25.030 0.610 ;
        RECT 25.850 0.320 26.950 0.610 ;
        RECT 27.770 0.320 28.870 0.610 ;
        RECT 29.690 0.320 30.790 0.610 ;
        RECT 31.610 0.320 32.710 0.610 ;
        RECT 33.530 0.320 34.630 0.610 ;
        RECT 35.450 0.320 36.550 0.610 ;
        RECT 37.370 0.320 38.470 0.610 ;
        RECT 39.290 0.320 40.390 0.610 ;
        RECT 41.210 0.320 42.310 0.610 ;
        RECT 43.130 0.320 44.230 0.610 ;
        RECT 45.050 0.320 46.150 0.610 ;
        RECT 46.970 0.320 48.070 0.610 ;
        RECT 48.890 0.320 59.140 0.610 ;
      LAYER Metal4 ;
        RECT 0.335 1.160 58.705 226.900 ;
      LAYER Metal5 ;
        RECT 5.660 1.115 18.050 221.485 ;
        RECT 20.670 1.115 24.250 221.485 ;
        RECT 26.870 1.115 54.820 221.485 ;
  END
END E_IO
END LIBRARY

