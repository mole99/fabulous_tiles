magic
tech ihp-sg13g2
magscale 1 2
timestamp 1743692709
<< metal1 >>
rect 1152 9848 20448 9872
rect 1152 9808 3688 9848
rect 3728 9808 3770 9848
rect 3810 9808 3852 9848
rect 3892 9808 3934 9848
rect 3974 9808 4016 9848
rect 4056 9808 18808 9848
rect 18848 9808 18890 9848
rect 18930 9808 18972 9848
rect 19012 9808 19054 9848
rect 19094 9808 19136 9848
rect 19176 9808 20448 9848
rect 1152 9784 20448 9808
rect 1563 9680 1605 9689
rect 1563 9640 1564 9680
rect 1604 9640 1605 9680
rect 1563 9631 1605 9640
rect 2331 9680 2373 9689
rect 2331 9640 2332 9680
rect 2372 9640 2373 9680
rect 2331 9631 2373 9640
rect 3099 9680 3141 9689
rect 3099 9640 3100 9680
rect 3140 9640 3141 9680
rect 3099 9631 3141 9640
rect 3483 9680 3525 9689
rect 3483 9640 3484 9680
rect 3524 9640 3525 9680
rect 3483 9631 3525 9640
rect 3867 9680 3909 9689
rect 3867 9640 3868 9680
rect 3908 9640 3909 9680
rect 3867 9631 3909 9640
rect 5019 9680 5061 9689
rect 5019 9640 5020 9680
rect 5060 9640 5061 9680
rect 5019 9631 5061 9640
rect 5403 9680 5445 9689
rect 5403 9640 5404 9680
rect 5444 9640 5445 9680
rect 5403 9631 5445 9640
rect 5787 9680 5829 9689
rect 5787 9640 5788 9680
rect 5828 9640 5829 9680
rect 5787 9631 5829 9640
rect 6171 9680 6213 9689
rect 6171 9640 6172 9680
rect 6212 9640 6213 9680
rect 6171 9631 6213 9640
rect 6555 9680 6597 9689
rect 6555 9640 6556 9680
rect 6596 9640 6597 9680
rect 6555 9631 6597 9640
rect 6939 9680 6981 9689
rect 6939 9640 6940 9680
rect 6980 9640 6981 9680
rect 6939 9631 6981 9640
rect 7707 9680 7749 9689
rect 7707 9640 7708 9680
rect 7748 9640 7749 9680
rect 7707 9631 7749 9640
rect 8187 9680 8229 9689
rect 8187 9640 8188 9680
rect 8228 9640 8229 9680
rect 8187 9631 8229 9640
rect 8571 9680 8613 9689
rect 8571 9640 8572 9680
rect 8612 9640 8613 9680
rect 8571 9631 8613 9640
rect 8955 9680 8997 9689
rect 8955 9640 8956 9680
rect 8996 9640 8997 9680
rect 8955 9631 8997 9640
rect 16155 9680 16197 9689
rect 16155 9640 16156 9680
rect 16196 9640 16197 9680
rect 16155 9631 16197 9640
rect 16539 9680 16581 9689
rect 16539 9640 16540 9680
rect 16580 9640 16581 9680
rect 16539 9631 16581 9640
rect 16923 9680 16965 9689
rect 16923 9640 16924 9680
rect 16964 9640 16965 9680
rect 16923 9631 16965 9640
rect 17691 9680 17733 9689
rect 17691 9640 17692 9680
rect 17732 9640 17733 9680
rect 17691 9631 17733 9640
rect 18459 9680 18501 9689
rect 18459 9640 18460 9680
rect 18500 9640 18501 9680
rect 18459 9631 18501 9640
rect 19611 9680 19653 9689
rect 19611 9640 19612 9680
rect 19652 9640 19653 9680
rect 19611 9631 19653 9640
rect 1947 9596 1989 9605
rect 1947 9556 1948 9596
rect 1988 9556 1989 9596
rect 1947 9547 1989 9556
rect 2715 9596 2757 9605
rect 2715 9556 2716 9596
rect 2756 9556 2757 9596
rect 2715 9547 2757 9556
rect 4251 9596 4293 9605
rect 4251 9556 4252 9596
rect 4292 9556 4293 9596
rect 4251 9547 4293 9556
rect 7323 9596 7365 9605
rect 7323 9556 7324 9596
rect 7364 9556 7365 9596
rect 7323 9547 7365 9556
rect 7803 9596 7845 9605
rect 7803 9556 7804 9596
rect 7844 9556 7845 9596
rect 7803 9547 7845 9556
rect 15675 9596 15717 9605
rect 15675 9556 15676 9596
rect 15716 9556 15717 9596
rect 15675 9547 15717 9556
rect 17307 9596 17349 9605
rect 17307 9556 17308 9596
rect 17348 9556 17349 9596
rect 17307 9547 17349 9556
rect 19227 9596 19269 9605
rect 19227 9556 19228 9596
rect 19268 9556 19269 9596
rect 19227 9547 19269 9556
rect 1323 9512 1365 9521
rect 1323 9472 1324 9512
rect 1364 9472 1365 9512
rect 1323 9463 1365 9472
rect 1707 9512 1749 9521
rect 1707 9472 1708 9512
rect 1748 9472 1749 9512
rect 1707 9463 1749 9472
rect 2091 9512 2133 9521
rect 2091 9472 2092 9512
rect 2132 9472 2133 9512
rect 2091 9463 2133 9472
rect 2475 9512 2517 9521
rect 2475 9472 2476 9512
rect 2516 9472 2517 9512
rect 2475 9463 2517 9472
rect 2859 9512 2901 9521
rect 2859 9472 2860 9512
rect 2900 9472 2901 9512
rect 2859 9463 2901 9472
rect 3243 9512 3285 9521
rect 3243 9472 3244 9512
rect 3284 9472 3285 9512
rect 3243 9463 3285 9472
rect 3627 9512 3669 9521
rect 3627 9472 3628 9512
rect 3668 9472 3669 9512
rect 3627 9463 3669 9472
rect 4011 9512 4053 9521
rect 4011 9472 4012 9512
rect 4052 9472 4053 9512
rect 4011 9463 4053 9472
rect 4395 9512 4437 9521
rect 4395 9472 4396 9512
rect 4436 9472 4437 9512
rect 4395 9463 4437 9472
rect 4635 9512 4677 9521
rect 4635 9472 4636 9512
rect 4676 9472 4677 9512
rect 4635 9463 4677 9472
rect 4779 9512 4821 9521
rect 4779 9472 4780 9512
rect 4820 9472 4821 9512
rect 4779 9463 4821 9472
rect 5163 9512 5205 9521
rect 5163 9472 5164 9512
rect 5204 9472 5205 9512
rect 5163 9463 5205 9472
rect 5547 9512 5589 9521
rect 5547 9472 5548 9512
rect 5588 9472 5589 9512
rect 5547 9463 5589 9472
rect 5931 9512 5973 9521
rect 5931 9472 5932 9512
rect 5972 9472 5973 9512
rect 5931 9463 5973 9472
rect 6315 9512 6357 9521
rect 6315 9472 6316 9512
rect 6356 9472 6357 9512
rect 6315 9463 6357 9472
rect 6699 9512 6741 9521
rect 6699 9472 6700 9512
rect 6740 9472 6741 9512
rect 6699 9463 6741 9472
rect 7083 9512 7125 9521
rect 7083 9472 7084 9512
rect 7124 9472 7125 9512
rect 7083 9463 7125 9472
rect 7467 9512 7509 9521
rect 7467 9472 7468 9512
rect 7508 9472 7509 9512
rect 7467 9463 7509 9472
rect 8043 9512 8085 9521
rect 8043 9472 8044 9512
rect 8084 9472 8085 9512
rect 8043 9463 8085 9472
rect 8427 9512 8469 9521
rect 8427 9472 8428 9512
rect 8468 9472 8469 9512
rect 8427 9463 8469 9472
rect 8811 9512 8853 9521
rect 8811 9472 8812 9512
rect 8852 9472 8853 9512
rect 8811 9463 8853 9472
rect 9195 9512 9237 9521
rect 9195 9472 9196 9512
rect 9236 9472 9237 9512
rect 9195 9463 9237 9472
rect 11883 9512 11925 9521
rect 11883 9472 11884 9512
rect 11924 9472 11925 9512
rect 11883 9463 11925 9472
rect 12843 9512 12885 9521
rect 12843 9472 12844 9512
rect 12884 9472 12885 9512
rect 12843 9463 12885 9472
rect 14571 9512 14613 9521
rect 14571 9472 14572 9512
rect 14612 9472 14613 9512
rect 14571 9463 14613 9472
rect 15051 9512 15093 9521
rect 15051 9472 15052 9512
rect 15092 9472 15093 9512
rect 15051 9463 15093 9472
rect 15435 9512 15477 9521
rect 15435 9472 15436 9512
rect 15476 9472 15477 9512
rect 15435 9463 15477 9472
rect 15819 9512 15861 9521
rect 15819 9472 15820 9512
rect 15860 9472 15861 9512
rect 15819 9463 15861 9472
rect 16395 9512 16437 9521
rect 16395 9472 16396 9512
rect 16436 9472 16437 9512
rect 16395 9463 16437 9472
rect 16779 9512 16821 9521
rect 16779 9472 16780 9512
rect 16820 9472 16821 9512
rect 16779 9463 16821 9472
rect 17163 9512 17205 9521
rect 17163 9472 17164 9512
rect 17204 9472 17205 9512
rect 17163 9463 17205 9472
rect 17547 9512 17589 9521
rect 17547 9472 17548 9512
rect 17588 9472 17589 9512
rect 17547 9463 17589 9472
rect 17931 9512 17973 9521
rect 17931 9472 17932 9512
rect 17972 9472 17973 9512
rect 17931 9463 17973 9472
rect 18315 9512 18357 9521
rect 18315 9472 18316 9512
rect 18356 9472 18357 9512
rect 18315 9463 18357 9472
rect 18699 9512 18741 9521
rect 18699 9472 18700 9512
rect 18740 9472 18741 9512
rect 18699 9463 18741 9472
rect 19083 9512 19125 9521
rect 19083 9472 19084 9512
rect 19124 9472 19125 9512
rect 19083 9463 19125 9472
rect 19467 9512 19509 9521
rect 19467 9472 19468 9512
rect 19508 9472 19509 9512
rect 19467 9463 19509 9472
rect 19851 9512 19893 9521
rect 19851 9472 19852 9512
rect 19892 9472 19893 9512
rect 19851 9463 19893 9472
rect 20235 9512 20277 9521
rect 20235 9472 20236 9512
rect 20276 9472 20277 9512
rect 20235 9463 20277 9472
rect 12123 9344 12165 9353
rect 12123 9304 12124 9344
rect 12164 9304 12165 9344
rect 12123 9295 12165 9304
rect 15291 9344 15333 9353
rect 15291 9304 15292 9344
rect 15332 9304 15333 9344
rect 15291 9295 15333 9304
rect 18075 9344 18117 9353
rect 18075 9304 18076 9344
rect 18116 9304 18117 9344
rect 18075 9295 18117 9304
rect 19995 9344 20037 9353
rect 19995 9304 19996 9344
rect 20036 9304 20037 9344
rect 19995 9295 20037 9304
rect 13083 9260 13125 9269
rect 13083 9220 13084 9260
rect 13124 9220 13125 9260
rect 13083 9211 13125 9220
rect 14811 9260 14853 9269
rect 14811 9220 14812 9260
rect 14852 9220 14853 9260
rect 14811 9211 14853 9220
rect 16059 9260 16101 9269
rect 16059 9220 16060 9260
rect 16100 9220 16101 9260
rect 16059 9211 16101 9220
rect 18843 9260 18885 9269
rect 18843 9220 18844 9260
rect 18884 9220 18885 9260
rect 18843 9211 18885 9220
rect 1152 9092 20452 9116
rect 1152 9052 4928 9092
rect 4968 9052 5010 9092
rect 5050 9052 5092 9092
rect 5132 9052 5174 9092
rect 5214 9052 5256 9092
rect 5296 9052 20048 9092
rect 20088 9052 20130 9092
rect 20170 9052 20212 9092
rect 20252 9052 20294 9092
rect 20334 9052 20376 9092
rect 20416 9052 20452 9092
rect 1152 9028 20452 9052
rect 1467 8924 1509 8933
rect 1467 8884 1468 8924
rect 1508 8884 1509 8924
rect 1467 8875 1509 8884
rect 2715 8924 2757 8933
rect 2715 8884 2716 8924
rect 2756 8884 2757 8924
rect 2715 8875 2757 8884
rect 3195 8924 3237 8933
rect 3195 8884 3196 8924
rect 3236 8884 3237 8924
rect 3195 8875 3237 8884
rect 3579 8924 3621 8933
rect 3579 8884 3580 8924
rect 3620 8884 3621 8924
rect 3579 8875 3621 8884
rect 3963 8924 4005 8933
rect 3963 8884 3964 8924
rect 4004 8884 4005 8924
rect 3963 8875 4005 8884
rect 4347 8924 4389 8933
rect 4347 8884 4348 8924
rect 4388 8884 4389 8924
rect 4347 8875 4389 8884
rect 4731 8924 4773 8933
rect 4731 8884 4732 8924
rect 4772 8884 4773 8924
rect 4731 8875 4773 8884
rect 5115 8924 5157 8933
rect 5115 8884 5116 8924
rect 5156 8884 5157 8924
rect 5115 8875 5157 8884
rect 5883 8924 5925 8933
rect 5883 8884 5884 8924
rect 5924 8884 5925 8924
rect 5883 8875 5925 8884
rect 6267 8924 6309 8933
rect 6267 8884 6268 8924
rect 6308 8884 6309 8924
rect 6267 8875 6309 8884
rect 6651 8924 6693 8933
rect 6651 8884 6652 8924
rect 6692 8884 6693 8924
rect 6651 8875 6693 8884
rect 7035 8924 7077 8933
rect 7035 8884 7036 8924
rect 7076 8884 7077 8924
rect 7035 8875 7077 8884
rect 7419 8924 7461 8933
rect 7419 8884 7420 8924
rect 7460 8884 7461 8924
rect 7419 8875 7461 8884
rect 16059 8924 16101 8933
rect 16059 8884 16060 8924
rect 16100 8884 16101 8924
rect 16059 8875 16101 8884
rect 16923 8924 16965 8933
rect 16923 8884 16924 8924
rect 16964 8884 16965 8924
rect 16923 8875 16965 8884
rect 18459 8924 18501 8933
rect 18459 8884 18460 8924
rect 18500 8884 18501 8924
rect 18459 8875 18501 8884
rect 19611 8924 19653 8933
rect 19611 8884 19612 8924
rect 19652 8884 19653 8924
rect 19611 8875 19653 8884
rect 19995 8924 20037 8933
rect 19995 8884 19996 8924
rect 20036 8884 20037 8924
rect 19995 8875 20037 8884
rect 1947 8840 1989 8849
rect 1947 8800 1948 8840
rect 1988 8800 1989 8840
rect 1947 8791 1989 8800
rect 5499 8840 5541 8849
rect 5499 8800 5500 8840
rect 5540 8800 5541 8840
rect 5499 8791 5541 8800
rect 17307 8840 17349 8849
rect 17307 8800 17308 8840
rect 17348 8800 17349 8840
rect 17307 8791 17349 8800
rect 18843 8840 18885 8849
rect 18843 8800 18844 8840
rect 18884 8800 18885 8840
rect 18843 8791 18885 8800
rect 19515 8840 19557 8849
rect 19515 8800 19516 8840
rect 19556 8800 19557 8840
rect 19515 8791 19557 8800
rect 1227 8672 1269 8681
rect 1227 8632 1228 8672
rect 1268 8632 1269 8672
rect 1227 8623 1269 8632
rect 1611 8672 1653 8681
rect 1611 8632 1612 8672
rect 1652 8632 1653 8672
rect 1611 8623 1653 8632
rect 1851 8672 1893 8681
rect 1851 8632 1852 8672
rect 1892 8632 1893 8672
rect 1851 8623 1893 8632
rect 2187 8672 2229 8681
rect 2187 8632 2188 8672
rect 2228 8632 2229 8672
rect 2187 8623 2229 8632
rect 2571 8672 2613 8681
rect 2571 8632 2572 8672
rect 2612 8632 2613 8672
rect 2571 8623 2613 8632
rect 2955 8672 2997 8681
rect 2955 8632 2956 8672
rect 2996 8632 2997 8672
rect 2955 8623 2997 8632
rect 3435 8672 3477 8681
rect 3435 8632 3436 8672
rect 3476 8632 3477 8672
rect 3435 8623 3477 8632
rect 3819 8672 3861 8681
rect 3819 8632 3820 8672
rect 3860 8632 3861 8672
rect 3819 8623 3861 8632
rect 4203 8672 4245 8681
rect 4203 8632 4204 8672
rect 4244 8632 4245 8672
rect 4203 8623 4245 8632
rect 4587 8672 4629 8681
rect 4587 8632 4588 8672
rect 4628 8632 4629 8672
rect 4587 8623 4629 8632
rect 4971 8672 5013 8681
rect 4971 8632 4972 8672
rect 5012 8632 5013 8672
rect 4971 8623 5013 8632
rect 5355 8672 5397 8681
rect 5355 8632 5356 8672
rect 5396 8632 5397 8672
rect 5355 8623 5397 8632
rect 5739 8672 5781 8681
rect 5739 8632 5740 8672
rect 5780 8632 5781 8672
rect 5739 8623 5781 8632
rect 6123 8672 6165 8681
rect 6123 8632 6124 8672
rect 6164 8632 6165 8672
rect 6123 8623 6165 8632
rect 6507 8672 6549 8681
rect 6507 8632 6508 8672
rect 6548 8632 6549 8672
rect 6507 8623 6549 8632
rect 6891 8672 6933 8681
rect 6891 8632 6892 8672
rect 6932 8632 6933 8672
rect 6891 8623 6933 8632
rect 7275 8672 7317 8681
rect 7275 8632 7276 8672
rect 7316 8632 7317 8672
rect 7275 8623 7317 8632
rect 7659 8672 7701 8681
rect 7659 8632 7660 8672
rect 7700 8632 7701 8672
rect 7659 8623 7701 8632
rect 13323 8672 13365 8681
rect 13323 8632 13324 8672
rect 13364 8632 13365 8672
rect 13323 8623 13365 8632
rect 13563 8672 13605 8681
rect 13563 8632 13564 8672
rect 13604 8632 13605 8672
rect 13563 8623 13605 8632
rect 15819 8672 15861 8681
rect 15819 8632 15820 8672
rect 15860 8632 15861 8672
rect 15819 8623 15861 8632
rect 16203 8672 16245 8681
rect 16203 8632 16204 8672
rect 16244 8632 16245 8672
rect 16203 8623 16245 8632
rect 16587 8672 16629 8681
rect 16587 8632 16588 8672
rect 16628 8632 16629 8672
rect 16587 8623 16629 8632
rect 17163 8672 17205 8681
rect 17163 8632 17164 8672
rect 17204 8632 17205 8672
rect 17163 8623 17205 8632
rect 17547 8672 17589 8681
rect 17547 8632 17548 8672
rect 17588 8632 17589 8672
rect 17547 8623 17589 8632
rect 17691 8672 17733 8681
rect 17691 8632 17692 8672
rect 17732 8632 17733 8672
rect 17691 8623 17733 8632
rect 17931 8672 17973 8681
rect 17931 8632 17932 8672
rect 17972 8632 17973 8672
rect 17931 8623 17973 8632
rect 18075 8672 18117 8681
rect 18075 8632 18076 8672
rect 18116 8632 18117 8672
rect 18075 8623 18117 8632
rect 18315 8672 18357 8681
rect 18315 8632 18316 8672
rect 18356 8632 18357 8672
rect 18315 8623 18357 8632
rect 18699 8672 18741 8681
rect 18699 8632 18700 8672
rect 18740 8632 18741 8672
rect 18699 8623 18741 8632
rect 19083 8672 19125 8681
rect 19083 8632 19084 8672
rect 19124 8632 19125 8672
rect 19083 8623 19125 8632
rect 19275 8672 19317 8681
rect 19275 8632 19276 8672
rect 19316 8632 19317 8672
rect 19275 8623 19317 8632
rect 19851 8672 19893 8681
rect 19851 8632 19852 8672
rect 19892 8632 19893 8672
rect 19851 8623 19893 8632
rect 20235 8672 20277 8681
rect 20235 8632 20236 8672
rect 20276 8632 20277 8672
rect 20235 8623 20277 8632
rect 16827 8588 16869 8597
rect 16827 8548 16828 8588
rect 16868 8548 16869 8588
rect 16827 8539 16869 8548
rect 2331 8504 2373 8513
rect 2331 8464 2332 8504
rect 2372 8464 2373 8504
rect 2331 8455 2373 8464
rect 16443 8504 16485 8513
rect 16443 8464 16444 8504
rect 16484 8464 16485 8504
rect 16443 8455 16485 8464
rect 1152 8336 20448 8360
rect 1152 8296 3688 8336
rect 3728 8296 3770 8336
rect 3810 8296 3852 8336
rect 3892 8296 3934 8336
rect 3974 8296 4016 8336
rect 4056 8296 18808 8336
rect 18848 8296 18890 8336
rect 18930 8296 18972 8336
rect 19012 8296 19054 8336
rect 19094 8296 19136 8336
rect 19176 8296 20448 8336
rect 1152 8272 20448 8296
rect 2043 8168 2085 8177
rect 2043 8128 2044 8168
rect 2084 8128 2085 8168
rect 2043 8119 2085 8128
rect 9915 8168 9957 8177
rect 9915 8128 9916 8168
rect 9956 8128 9957 8168
rect 9915 8119 9957 8128
rect 10299 8168 10341 8177
rect 10299 8128 10300 8168
rect 10340 8128 10341 8168
rect 10299 8119 10341 8128
rect 16923 8168 16965 8177
rect 16923 8128 16924 8168
rect 16964 8128 16965 8168
rect 16923 8119 16965 8128
rect 17307 8168 17349 8177
rect 17307 8128 17308 8168
rect 17348 8128 17349 8168
rect 17307 8119 17349 8128
rect 18075 8168 18117 8177
rect 18075 8128 18076 8168
rect 18116 8128 18117 8168
rect 18075 8119 18117 8128
rect 18555 8168 18597 8177
rect 18555 8128 18556 8168
rect 18596 8128 18597 8168
rect 18555 8119 18597 8128
rect 18939 8084 18981 8093
rect 18939 8044 18940 8084
rect 18980 8044 18981 8084
rect 18939 8035 18981 8044
rect 19611 8084 19653 8093
rect 19611 8044 19612 8084
rect 19652 8044 19653 8084
rect 19611 8035 19653 8044
rect 2283 8000 2325 8009
rect 2283 7960 2284 8000
rect 2324 7960 2325 8000
rect 2283 7951 2325 7960
rect 10155 8000 10197 8009
rect 10155 7960 10156 8000
rect 10196 7960 10197 8000
rect 10155 7951 10197 7960
rect 10539 8000 10581 8009
rect 10539 7960 10540 8000
rect 10580 7960 10581 8000
rect 10539 7951 10581 7960
rect 16299 8000 16341 8009
rect 16299 7960 16300 8000
rect 16340 7960 16341 8000
rect 16299 7951 16341 7960
rect 16683 8000 16725 8009
rect 16683 7960 16684 8000
rect 16724 7960 16725 8000
rect 16683 7951 16725 7960
rect 17067 8000 17109 8009
rect 17067 7960 17068 8000
rect 17108 7960 17109 8000
rect 17067 7951 17109 7960
rect 17451 8000 17493 8009
rect 17451 7960 17452 8000
rect 17492 7960 17493 8000
rect 17451 7951 17493 7960
rect 17835 8000 17877 8009
rect 17835 7960 17836 8000
rect 17876 7960 17877 8000
rect 17835 7951 17877 7960
rect 18411 8000 18453 8009
rect 18411 7960 18412 8000
rect 18452 7960 18453 8000
rect 18411 7951 18453 7960
rect 18795 8000 18837 8009
rect 18795 7960 18796 8000
rect 18836 7960 18837 8000
rect 18795 7951 18837 7960
rect 19179 8000 19221 8009
rect 19179 7960 19180 8000
rect 19220 7960 19221 8000
rect 19179 7951 19221 7960
rect 19371 8000 19413 8009
rect 19371 7960 19372 8000
rect 19412 7960 19413 8000
rect 19371 7951 19413 7960
rect 19755 8000 19797 8009
rect 19755 7960 19756 8000
rect 19796 7960 19797 8000
rect 19755 7951 19797 7960
rect 20139 8000 20181 8009
rect 20139 7960 20140 8000
rect 20180 7960 20181 8000
rect 20139 7951 20181 7960
rect 16539 7748 16581 7757
rect 16539 7708 16540 7748
rect 16580 7708 16581 7748
rect 16539 7699 16581 7708
rect 17691 7748 17733 7757
rect 17691 7708 17692 7748
rect 17732 7708 17733 7748
rect 17691 7699 17733 7708
rect 18171 7748 18213 7757
rect 18171 7708 18172 7748
rect 18212 7708 18213 7748
rect 18171 7699 18213 7708
rect 19995 7748 20037 7757
rect 19995 7708 19996 7748
rect 20036 7708 20037 7748
rect 19995 7699 20037 7708
rect 20379 7748 20421 7757
rect 20379 7708 20380 7748
rect 20420 7708 20421 7748
rect 20379 7699 20421 7708
rect 1152 7580 20452 7604
rect 1152 7540 4928 7580
rect 4968 7540 5010 7580
rect 5050 7540 5092 7580
rect 5132 7540 5174 7580
rect 5214 7540 5256 7580
rect 5296 7540 20048 7580
rect 20088 7540 20130 7580
rect 20170 7540 20212 7580
rect 20252 7540 20294 7580
rect 20334 7540 20376 7580
rect 20416 7540 20452 7580
rect 1152 7516 20452 7540
rect 5883 7412 5925 7421
rect 5883 7372 5884 7412
rect 5924 7372 5925 7412
rect 5883 7363 5925 7372
rect 13947 7412 13989 7421
rect 13947 7372 13948 7412
rect 13988 7372 13989 7412
rect 13947 7363 13989 7372
rect 18555 7412 18597 7421
rect 18555 7372 18556 7412
rect 18596 7372 18597 7412
rect 18555 7363 18597 7372
rect 16059 7328 16101 7337
rect 16059 7288 16060 7328
rect 16100 7288 16101 7328
rect 16059 7279 16101 7288
rect 1947 7160 1989 7169
rect 1947 7120 1948 7160
rect 1988 7120 1989 7160
rect 1947 7111 1989 7120
rect 2187 7160 2229 7169
rect 2187 7120 2188 7160
rect 2228 7120 2229 7160
rect 2187 7111 2229 7120
rect 4347 7160 4389 7169
rect 4347 7120 4348 7160
rect 4388 7120 4389 7160
rect 4347 7111 4389 7120
rect 4587 7160 4629 7169
rect 4587 7120 4588 7160
rect 4628 7120 4629 7160
rect 4587 7111 4629 7120
rect 5211 7160 5253 7169
rect 5211 7120 5212 7160
rect 5252 7120 5253 7160
rect 5211 7111 5253 7120
rect 5451 7160 5493 7169
rect 5451 7120 5452 7160
rect 5492 7120 5493 7160
rect 5451 7111 5493 7120
rect 5643 7160 5685 7169
rect 5643 7120 5644 7160
rect 5684 7120 5685 7160
rect 5643 7111 5685 7120
rect 10155 7160 10197 7169
rect 10155 7120 10156 7160
rect 10196 7120 10197 7160
rect 10155 7111 10197 7120
rect 10299 7160 10341 7169
rect 10299 7120 10300 7160
rect 10340 7120 10341 7160
rect 10299 7111 10341 7120
rect 10539 7160 10581 7169
rect 10539 7120 10540 7160
rect 10580 7120 10581 7160
rect 10539 7111 10581 7120
rect 11835 7160 11877 7169
rect 11835 7120 11836 7160
rect 11876 7120 11877 7160
rect 11835 7111 11877 7120
rect 12075 7160 12117 7169
rect 12075 7120 12076 7160
rect 12116 7120 12117 7160
rect 12075 7111 12117 7120
rect 12459 7160 12501 7169
rect 12459 7120 12460 7160
rect 12500 7120 12501 7160
rect 12459 7111 12501 7120
rect 13563 7160 13605 7169
rect 13563 7120 13564 7160
rect 13604 7120 13605 7160
rect 13563 7111 13605 7120
rect 13803 7160 13845 7169
rect 13803 7120 13804 7160
rect 13844 7120 13845 7160
rect 13803 7111 13845 7120
rect 14187 7160 14229 7169
rect 14187 7120 14188 7160
rect 14228 7120 14229 7160
rect 14187 7111 14229 7120
rect 15387 7160 15429 7169
rect 15387 7120 15388 7160
rect 15428 7120 15429 7160
rect 15387 7111 15429 7120
rect 15627 7160 15669 7169
rect 15627 7120 15628 7160
rect 15668 7120 15669 7160
rect 15627 7111 15669 7120
rect 16299 7160 16341 7169
rect 16299 7120 16300 7160
rect 16340 7120 16341 7160
rect 16299 7111 16341 7120
rect 16875 7160 16917 7169
rect 16875 7120 16876 7160
rect 16916 7120 16917 7160
rect 16875 7111 16917 7120
rect 17259 7160 17301 7169
rect 17259 7120 17260 7160
rect 17300 7120 17301 7160
rect 17259 7111 17301 7120
rect 17547 7160 17589 7169
rect 17547 7120 17548 7160
rect 17588 7120 17589 7160
rect 17547 7111 17589 7120
rect 17787 7160 17829 7169
rect 17787 7120 17788 7160
rect 17828 7120 17829 7160
rect 17787 7111 17829 7120
rect 18123 7160 18165 7169
rect 18123 7120 18124 7160
rect 18164 7120 18165 7160
rect 18123 7111 18165 7120
rect 18315 7160 18357 7169
rect 18315 7120 18316 7160
rect 18356 7120 18357 7160
rect 18315 7111 18357 7120
rect 18699 7160 18741 7169
rect 18699 7120 18700 7160
rect 18740 7120 18741 7160
rect 18699 7111 18741 7120
rect 19083 7160 19125 7169
rect 19083 7120 19084 7160
rect 19124 7120 19125 7160
rect 19083 7111 19125 7120
rect 19659 7160 19701 7169
rect 19659 7120 19660 7160
rect 19700 7120 19701 7160
rect 19659 7111 19701 7120
rect 20139 7160 20181 7169
rect 20139 7120 20140 7160
rect 20180 7120 20181 7160
rect 20139 7111 20181 7120
rect 9915 7076 9957 7085
rect 9915 7036 9916 7076
rect 9956 7036 9957 7076
rect 9915 7027 9957 7036
rect 19323 7076 19365 7085
rect 19323 7036 19324 7076
rect 19364 7036 19365 7076
rect 19323 7027 19365 7036
rect 12219 6992 12261 7001
rect 12219 6952 12220 6992
rect 12260 6952 12261 6992
rect 12219 6943 12261 6952
rect 16635 6992 16677 7001
rect 16635 6952 16636 6992
rect 16676 6952 16677 6992
rect 16635 6943 16677 6952
rect 17019 6992 17061 7001
rect 17019 6952 17020 6992
rect 17060 6952 17061 6992
rect 17019 6943 17061 6952
rect 17883 6992 17925 7001
rect 17883 6952 17884 6992
rect 17924 6952 17925 6992
rect 17883 6943 17925 6952
rect 18939 6992 18981 7001
rect 18939 6952 18940 6992
rect 18980 6952 18981 6992
rect 18939 6943 18981 6952
rect 19419 6992 19461 7001
rect 19419 6952 19420 6992
rect 19460 6952 19461 6992
rect 19419 6943 19461 6952
rect 20379 6992 20421 7001
rect 20379 6952 20380 6992
rect 20420 6952 20421 6992
rect 20379 6943 20421 6952
rect 1152 6824 20448 6848
rect 1152 6784 3688 6824
rect 3728 6784 3770 6824
rect 3810 6784 3852 6824
rect 3892 6784 3934 6824
rect 3974 6784 4016 6824
rect 4056 6784 18808 6824
rect 18848 6784 18890 6824
rect 18930 6784 18972 6824
rect 19012 6784 19054 6824
rect 19094 6784 19136 6824
rect 19176 6784 20448 6824
rect 1152 6760 20448 6784
rect 12699 6656 12741 6665
rect 12699 6616 12700 6656
rect 12740 6616 12741 6656
rect 12699 6607 12741 6616
rect 18651 6656 18693 6665
rect 18651 6616 18652 6656
rect 18692 6616 18693 6656
rect 18651 6607 18693 6616
rect 19035 6656 19077 6665
rect 19035 6616 19036 6656
rect 19076 6616 19077 6656
rect 19035 6607 19077 6616
rect 19419 6656 19461 6665
rect 19419 6616 19420 6656
rect 19460 6616 19461 6656
rect 19419 6607 19461 6616
rect 20379 6656 20421 6665
rect 20379 6616 20380 6656
rect 20420 6616 20421 6656
rect 20379 6607 20421 6616
rect 3339 6488 3381 6497
rect 3339 6448 3340 6488
rect 3380 6448 3381 6488
rect 3339 6439 3381 6448
rect 4395 6488 4437 6497
rect 4395 6448 4396 6488
rect 4436 6448 4437 6488
rect 4395 6439 4437 6448
rect 9147 6488 9189 6497
rect 9147 6448 9148 6488
rect 9188 6448 9189 6488
rect 9147 6439 9189 6448
rect 9387 6488 9429 6497
rect 9387 6448 9388 6488
rect 9428 6448 9429 6488
rect 9387 6439 9429 6448
rect 12939 6488 12981 6497
rect 12939 6448 12940 6488
rect 12980 6448 12981 6488
rect 12939 6439 12981 6448
rect 13323 6488 13365 6497
rect 13323 6448 13324 6488
rect 13364 6448 13365 6488
rect 13323 6439 13365 6448
rect 14667 6488 14709 6497
rect 14667 6448 14668 6488
rect 14708 6448 14709 6488
rect 14667 6439 14709 6448
rect 14907 6488 14949 6497
rect 14907 6448 14908 6488
rect 14948 6448 14949 6488
rect 14907 6439 14949 6448
rect 18411 6488 18453 6497
rect 18411 6448 18412 6488
rect 18452 6448 18453 6488
rect 18411 6439 18453 6448
rect 18795 6488 18837 6497
rect 18795 6448 18796 6488
rect 18836 6448 18837 6488
rect 18795 6439 18837 6448
rect 19179 6488 19221 6497
rect 19179 6448 19180 6488
rect 19220 6448 19221 6488
rect 19179 6439 19221 6448
rect 19755 6488 19797 6497
rect 19755 6448 19756 6488
rect 19796 6448 19797 6488
rect 19755 6439 19797 6448
rect 20139 6488 20181 6497
rect 20139 6448 20140 6488
rect 20180 6448 20181 6488
rect 20139 6439 20181 6448
rect 3579 6320 3621 6329
rect 3579 6280 3580 6320
rect 3620 6280 3621 6320
rect 3579 6271 3621 6280
rect 13083 6320 13125 6329
rect 13083 6280 13084 6320
rect 13124 6280 13125 6320
rect 13083 6271 13125 6280
rect 4635 6236 4677 6245
rect 4635 6196 4636 6236
rect 4676 6196 4677 6236
rect 4635 6187 4677 6196
rect 19515 6236 19557 6245
rect 19515 6196 19516 6236
rect 19556 6196 19557 6236
rect 19515 6187 19557 6196
rect 1152 6068 20452 6092
rect 1152 6028 4928 6068
rect 4968 6028 5010 6068
rect 5050 6028 5092 6068
rect 5132 6028 5174 6068
rect 5214 6028 5256 6068
rect 5296 6028 20048 6068
rect 20088 6028 20130 6068
rect 20170 6028 20212 6068
rect 20252 6028 20294 6068
rect 20334 6028 20376 6068
rect 20416 6028 20452 6068
rect 1152 6004 20452 6028
rect 19131 5900 19173 5909
rect 19131 5860 19132 5900
rect 19172 5860 19173 5900
rect 19131 5851 19173 5860
rect 19995 5900 20037 5909
rect 19995 5860 19996 5900
rect 20036 5860 20037 5900
rect 19995 5851 20037 5860
rect 12315 5816 12357 5825
rect 12315 5776 12316 5816
rect 12356 5776 12357 5816
rect 12315 5767 12357 5776
rect 3195 5648 3237 5657
rect 3195 5608 3196 5648
rect 3236 5608 3237 5648
rect 3195 5599 3237 5608
rect 3435 5648 3477 5657
rect 3435 5608 3436 5648
rect 3476 5608 3477 5648
rect 3435 5599 3477 5608
rect 4779 5648 4821 5657
rect 4779 5608 4780 5648
rect 4820 5608 4821 5648
rect 4779 5599 4821 5608
rect 5835 5648 5877 5657
rect 5835 5608 5836 5648
rect 5876 5608 5877 5648
rect 5835 5599 5877 5608
rect 8283 5648 8325 5657
rect 8283 5608 8284 5648
rect 8324 5608 8325 5648
rect 8283 5599 8325 5608
rect 8523 5648 8565 5657
rect 8523 5608 8524 5648
rect 8564 5608 8565 5648
rect 8523 5599 8565 5608
rect 9291 5648 9333 5657
rect 9291 5608 9292 5648
rect 9332 5608 9333 5648
rect 9291 5599 9333 5608
rect 10635 5648 10677 5657
rect 10635 5608 10636 5648
rect 10676 5608 10677 5648
rect 10635 5599 10677 5608
rect 11019 5648 11061 5657
rect 11019 5608 11020 5648
rect 11060 5608 11061 5648
rect 11019 5599 11061 5608
rect 12075 5648 12117 5657
rect 12075 5608 12076 5648
rect 12116 5608 12117 5648
rect 12075 5599 12117 5608
rect 14955 5648 14997 5657
rect 14955 5608 14956 5648
rect 14996 5608 14997 5648
rect 14955 5599 14997 5608
rect 15195 5648 15237 5657
rect 15195 5608 15196 5648
rect 15236 5608 15237 5648
rect 15195 5599 15237 5608
rect 18219 5648 18261 5657
rect 18219 5608 18220 5648
rect 18260 5608 18261 5648
rect 18219 5599 18261 5608
rect 18795 5648 18837 5657
rect 18795 5608 18796 5648
rect 18836 5608 18837 5648
rect 18795 5599 18837 5608
rect 19371 5648 19413 5657
rect 19371 5608 19372 5648
rect 19412 5608 19413 5648
rect 19371 5599 19413 5608
rect 19755 5648 19797 5657
rect 19755 5608 19756 5648
rect 19796 5608 19797 5648
rect 19755 5599 19797 5608
rect 20139 5648 20181 5657
rect 20139 5608 20140 5648
rect 20180 5608 20181 5648
rect 20139 5599 20181 5608
rect 20379 5648 20421 5657
rect 20379 5608 20380 5648
rect 20420 5608 20421 5648
rect 20379 5599 20421 5608
rect 4539 5564 4581 5573
rect 4539 5524 4540 5564
rect 4580 5524 4581 5564
rect 4539 5515 4581 5524
rect 19035 5564 19077 5573
rect 19035 5524 19036 5564
rect 19076 5524 19077 5564
rect 19035 5515 19077 5524
rect 5595 5480 5637 5489
rect 5595 5440 5596 5480
rect 5636 5440 5637 5480
rect 5595 5431 5637 5440
rect 9531 5480 9573 5489
rect 9531 5440 9532 5480
rect 9572 5440 9573 5480
rect 9531 5431 9573 5440
rect 10875 5480 10917 5489
rect 10875 5440 10876 5480
rect 10916 5440 10917 5480
rect 10875 5431 10917 5440
rect 11259 5480 11301 5489
rect 11259 5440 11260 5480
rect 11300 5440 11301 5480
rect 11259 5431 11301 5440
rect 17979 5480 18021 5489
rect 17979 5440 17980 5480
rect 18020 5440 18021 5480
rect 17979 5431 18021 5440
rect 1152 5312 20448 5336
rect 1152 5272 3688 5312
rect 3728 5272 3770 5312
rect 3810 5272 3852 5312
rect 3892 5272 3934 5312
rect 3974 5272 4016 5312
rect 4056 5272 18808 5312
rect 18848 5272 18890 5312
rect 18930 5272 18972 5312
rect 19012 5272 19054 5312
rect 19094 5272 19136 5312
rect 19176 5272 20448 5312
rect 1152 5248 20448 5272
rect 16251 5144 16293 5153
rect 16251 5104 16252 5144
rect 16292 5104 16293 5144
rect 16251 5095 16293 5104
rect 19995 5144 20037 5153
rect 19995 5104 19996 5144
rect 20036 5104 20037 5144
rect 19995 5095 20037 5104
rect 7035 5060 7077 5069
rect 7035 5020 7036 5060
rect 7076 5020 7077 5060
rect 7035 5011 7077 5020
rect 7611 5060 7653 5069
rect 7611 5020 7612 5060
rect 7652 5020 7653 5060
rect 7611 5011 7653 5020
rect 20379 5060 20421 5069
rect 20379 5020 20380 5060
rect 20420 5020 20421 5060
rect 20379 5011 20421 5020
rect 3723 4976 3765 4985
rect 3723 4936 3724 4976
rect 3764 4936 3765 4976
rect 3723 4927 3765 4936
rect 5163 4976 5205 4985
rect 5163 4936 5164 4976
rect 5204 4936 5205 4976
rect 5163 4927 5205 4936
rect 6651 4976 6693 4985
rect 6651 4936 6652 4976
rect 6692 4936 6693 4976
rect 6651 4927 6693 4936
rect 6891 4976 6933 4985
rect 6891 4936 6892 4976
rect 6932 4936 6933 4976
rect 6891 4927 6933 4936
rect 7275 4976 7317 4985
rect 7275 4936 7276 4976
rect 7316 4936 7317 4976
rect 7275 4927 7317 4936
rect 7851 4976 7893 4985
rect 7851 4936 7852 4976
rect 7892 4936 7893 4976
rect 7851 4927 7893 4936
rect 8091 4976 8133 4985
rect 8091 4936 8092 4976
rect 8132 4936 8133 4976
rect 8091 4927 8133 4936
rect 8331 4976 8373 4985
rect 8331 4936 8332 4976
rect 8372 4936 8373 4976
rect 8331 4927 8373 4936
rect 13803 4976 13845 4985
rect 13803 4936 13804 4976
rect 13844 4936 13845 4976
rect 13803 4927 13845 4936
rect 16011 4976 16053 4985
rect 16011 4936 16012 4976
rect 16052 4936 16053 4976
rect 16011 4927 16053 4936
rect 18699 4976 18741 4985
rect 18699 4936 18700 4976
rect 18740 4936 18741 4976
rect 18699 4927 18741 4936
rect 19035 4976 19077 4985
rect 19035 4936 19036 4976
rect 19076 4936 19077 4976
rect 19035 4927 19077 4936
rect 19275 4976 19317 4985
rect 19275 4936 19276 4976
rect 19316 4936 19317 4976
rect 19275 4927 19317 4936
rect 19755 4976 19797 4985
rect 19755 4936 19756 4976
rect 19796 4936 19797 4976
rect 19755 4927 19797 4936
rect 20139 4976 20181 4985
rect 20139 4936 20140 4976
rect 20180 4936 20181 4976
rect 20139 4927 20181 4936
rect 3963 4808 4005 4817
rect 3963 4768 3964 4808
rect 4004 4768 4005 4808
rect 3963 4759 4005 4768
rect 5403 4724 5445 4733
rect 5403 4684 5404 4724
rect 5444 4684 5445 4724
rect 5403 4675 5445 4684
rect 14043 4724 14085 4733
rect 14043 4684 14044 4724
rect 14084 4684 14085 4724
rect 14043 4675 14085 4684
rect 18939 4724 18981 4733
rect 18939 4684 18940 4724
rect 18980 4684 18981 4724
rect 18939 4675 18981 4684
rect 1152 4556 20452 4580
rect 1152 4516 4928 4556
rect 4968 4516 5010 4556
rect 5050 4516 5092 4556
rect 5132 4516 5174 4556
rect 5214 4516 5256 4556
rect 5296 4516 20048 4556
rect 20088 4516 20130 4556
rect 20170 4516 20212 4556
rect 20252 4516 20294 4556
rect 20334 4516 20376 4556
rect 20416 4516 20452 4556
rect 1152 4492 20452 4516
rect 12123 4304 12165 4313
rect 12123 4264 12124 4304
rect 12164 4264 12165 4304
rect 12123 4255 12165 4264
rect 15387 4304 15429 4313
rect 15387 4264 15388 4304
rect 15428 4264 15429 4304
rect 15387 4255 15429 4264
rect 19131 4304 19173 4313
rect 19131 4264 19132 4304
rect 19172 4264 19173 4304
rect 19131 4255 19173 4264
rect 20379 4304 20421 4313
rect 20379 4264 20380 4304
rect 20420 4264 20421 4304
rect 20379 4255 20421 4264
rect 3867 4136 3909 4145
rect 3867 4096 3868 4136
rect 3908 4096 3909 4136
rect 3867 4087 3909 4096
rect 4107 4136 4149 4145
rect 4107 4096 4108 4136
rect 4148 4096 4149 4136
rect 4107 4087 4149 4096
rect 11883 4136 11925 4145
rect 11883 4096 11884 4136
rect 11924 4096 11925 4136
rect 11883 4087 11925 4096
rect 15147 4136 15189 4145
rect 15147 4096 15148 4136
rect 15188 4096 15189 4136
rect 15147 4087 15189 4096
rect 18795 4136 18837 4145
rect 18795 4096 18796 4136
rect 18836 4096 18837 4136
rect 18795 4087 18837 4096
rect 19371 4136 19413 4145
rect 19371 4096 19372 4136
rect 19412 4096 19413 4136
rect 19371 4087 19413 4096
rect 19594 4136 19652 4137
rect 19594 4096 19603 4136
rect 19643 4096 19652 4136
rect 19594 4095 19652 4096
rect 20139 4136 20181 4145
rect 20139 4096 20140 4136
rect 20180 4096 20181 4136
rect 20139 4087 20181 4096
rect 19035 4052 19077 4061
rect 19035 4012 19036 4052
rect 19076 4012 19077 4052
rect 19035 4003 19077 4012
rect 19803 3968 19845 3977
rect 19803 3928 19804 3968
rect 19844 3928 19845 3968
rect 19803 3919 19845 3928
rect 1152 3800 20448 3824
rect 1152 3760 3688 3800
rect 3728 3760 3770 3800
rect 3810 3760 3852 3800
rect 3892 3760 3934 3800
rect 3974 3760 4016 3800
rect 4056 3760 18808 3800
rect 18848 3760 18890 3800
rect 18930 3760 18972 3800
rect 19012 3760 19054 3800
rect 19094 3760 19136 3800
rect 19176 3760 20448 3800
rect 1152 3736 20448 3760
rect 9147 3632 9189 3641
rect 9147 3592 9148 3632
rect 9188 3592 9189 3632
rect 9147 3583 9189 3592
rect 10971 3632 11013 3641
rect 10971 3592 10972 3632
rect 11012 3592 11013 3632
rect 10971 3583 11013 3592
rect 13659 3632 13701 3641
rect 13659 3592 13660 3632
rect 13700 3592 13701 3632
rect 13659 3583 13701 3592
rect 14043 3632 14085 3641
rect 14043 3592 14044 3632
rect 14084 3592 14085 3632
rect 14043 3583 14085 3592
rect 16827 3632 16869 3641
rect 16827 3592 16828 3632
rect 16868 3592 16869 3632
rect 16827 3583 16869 3592
rect 20379 3632 20421 3641
rect 20379 3592 20380 3632
rect 20420 3592 20421 3632
rect 20379 3583 20421 3592
rect 1899 3464 1941 3473
rect 1899 3424 1900 3464
rect 1940 3424 1941 3464
rect 1899 3415 1941 3424
rect 6315 3464 6357 3473
rect 6315 3424 6316 3464
rect 6356 3424 6357 3464
rect 6315 3415 6357 3424
rect 8523 3464 8565 3473
rect 8523 3424 8524 3464
rect 8564 3424 8565 3464
rect 8523 3415 8565 3424
rect 8907 3464 8949 3473
rect 8907 3424 8908 3464
rect 8948 3424 8949 3464
rect 8907 3415 8949 3424
rect 9963 3464 10005 3473
rect 9963 3424 9964 3464
rect 10004 3424 10005 3464
rect 9963 3415 10005 3424
rect 10731 3464 10773 3473
rect 10731 3424 10732 3464
rect 10772 3424 10773 3464
rect 10731 3415 10773 3424
rect 12075 3464 12117 3473
rect 12075 3424 12076 3464
rect 12116 3424 12117 3464
rect 12075 3415 12117 3424
rect 13419 3464 13461 3473
rect 13419 3424 13420 3464
rect 13460 3424 13461 3464
rect 13419 3415 13461 3424
rect 13803 3464 13845 3473
rect 13803 3424 13804 3464
rect 13844 3424 13845 3464
rect 13803 3415 13845 3424
rect 14955 3464 14997 3473
rect 14955 3424 14956 3464
rect 14996 3424 14997 3464
rect 14955 3415 14997 3424
rect 16587 3464 16629 3473
rect 16587 3424 16588 3464
rect 16628 3424 16629 3464
rect 16587 3415 16629 3424
rect 16971 3464 17013 3473
rect 16971 3424 16972 3464
rect 17012 3424 17013 3464
rect 16971 3415 17013 3424
rect 19371 3464 19413 3473
rect 19371 3424 19372 3464
rect 19412 3424 19413 3464
rect 19371 3415 19413 3424
rect 19786 3464 19844 3465
rect 19786 3424 19795 3464
rect 19835 3424 19844 3464
rect 19786 3423 19844 3424
rect 20139 3464 20181 3473
rect 20139 3424 20140 3464
rect 20180 3424 20181 3464
rect 20139 3415 20181 3424
rect 2139 3296 2181 3305
rect 2139 3256 2140 3296
rect 2180 3256 2181 3296
rect 2139 3247 2181 3256
rect 8763 3296 8805 3305
rect 8763 3256 8764 3296
rect 8804 3256 8805 3296
rect 8763 3247 8805 3256
rect 19611 3296 19653 3305
rect 19611 3256 19612 3296
rect 19652 3256 19653 3296
rect 19611 3247 19653 3256
rect 6555 3212 6597 3221
rect 6555 3172 6556 3212
rect 6596 3172 6597 3212
rect 6555 3163 6597 3172
rect 10203 3212 10245 3221
rect 10203 3172 10204 3212
rect 10244 3172 10245 3212
rect 10203 3163 10245 3172
rect 12315 3212 12357 3221
rect 12315 3172 12316 3212
rect 12356 3172 12357 3212
rect 12315 3163 12357 3172
rect 15195 3212 15237 3221
rect 15195 3172 15196 3212
rect 15236 3172 15237 3212
rect 15195 3163 15237 3172
rect 17211 3212 17253 3221
rect 17211 3172 17212 3212
rect 17252 3172 17253 3212
rect 17211 3163 17253 3172
rect 19995 3212 20037 3221
rect 19995 3172 19996 3212
rect 20036 3172 20037 3212
rect 19995 3163 20037 3172
rect 1152 3044 20452 3068
rect 1152 3004 4928 3044
rect 4968 3004 5010 3044
rect 5050 3004 5092 3044
rect 5132 3004 5174 3044
rect 5214 3004 5256 3044
rect 5296 3004 20048 3044
rect 20088 3004 20130 3044
rect 20170 3004 20212 3044
rect 20252 3004 20294 3044
rect 20334 3004 20376 3044
rect 20416 3004 20452 3044
rect 1152 2980 20452 3004
rect 18843 2876 18885 2885
rect 18843 2836 18844 2876
rect 18884 2836 18885 2876
rect 18843 2827 18885 2836
rect 19995 2876 20037 2885
rect 19995 2836 19996 2876
rect 20036 2836 20037 2876
rect 19995 2827 20037 2836
rect 20379 2876 20421 2885
rect 20379 2836 20380 2876
rect 20420 2836 20421 2876
rect 20379 2827 20421 2836
rect 6603 2624 6645 2633
rect 6603 2584 6604 2624
rect 6644 2584 6645 2624
rect 6603 2575 6645 2584
rect 17163 2624 17205 2633
rect 17163 2584 17164 2624
rect 17204 2584 17205 2624
rect 17163 2575 17205 2584
rect 18123 2624 18165 2633
rect 18123 2584 18124 2624
rect 18164 2584 18165 2624
rect 18123 2575 18165 2584
rect 18603 2624 18645 2633
rect 18603 2584 18604 2624
rect 18644 2584 18645 2624
rect 18603 2575 18645 2584
rect 18987 2624 19029 2633
rect 18987 2584 18988 2624
rect 19028 2584 19029 2624
rect 18987 2575 19029 2584
rect 19371 2624 19413 2633
rect 19371 2584 19372 2624
rect 19412 2584 19413 2624
rect 19371 2575 19413 2584
rect 19755 2624 19797 2633
rect 19755 2584 19756 2624
rect 19796 2584 19797 2624
rect 19755 2575 19797 2584
rect 20139 2624 20181 2633
rect 20139 2584 20140 2624
rect 20180 2584 20181 2624
rect 20139 2575 20181 2584
rect 19227 2540 19269 2549
rect 19227 2500 19228 2540
rect 19268 2500 19269 2540
rect 19227 2491 19269 2500
rect 6843 2456 6885 2465
rect 6843 2416 6844 2456
rect 6884 2416 6885 2456
rect 6843 2407 6885 2416
rect 17403 2456 17445 2465
rect 17403 2416 17404 2456
rect 17444 2416 17445 2456
rect 17403 2407 17445 2416
rect 18363 2456 18405 2465
rect 18363 2416 18364 2456
rect 18404 2416 18405 2456
rect 18363 2407 18405 2416
rect 19611 2456 19653 2465
rect 19611 2416 19612 2456
rect 19652 2416 19653 2456
rect 19611 2407 19653 2416
rect 1152 2288 20448 2312
rect 1152 2248 3688 2288
rect 3728 2248 3770 2288
rect 3810 2248 3852 2288
rect 3892 2248 3934 2288
rect 3974 2248 4016 2288
rect 4056 2248 18808 2288
rect 18848 2248 18890 2288
rect 18930 2248 18972 2288
rect 19012 2248 19054 2288
rect 19094 2248 19136 2288
rect 19176 2248 20448 2288
rect 1152 2224 20448 2248
rect 19995 2120 20037 2129
rect 19995 2080 19996 2120
rect 20036 2080 20037 2120
rect 19995 2071 20037 2080
rect 18555 2036 18597 2045
rect 18555 1996 18556 2036
rect 18596 1996 18597 2036
rect 18555 1987 18597 1996
rect 20379 2036 20421 2045
rect 20379 1996 20380 2036
rect 20420 1996 20421 2036
rect 20379 1987 20421 1996
rect 12939 1952 12981 1961
rect 12939 1912 12940 1952
rect 12980 1912 12981 1952
rect 12939 1903 12981 1912
rect 15339 1952 15381 1961
rect 15339 1912 15340 1952
rect 15380 1912 15381 1952
rect 15339 1903 15381 1912
rect 17931 1952 17973 1961
rect 17931 1912 17932 1952
rect 17972 1912 17973 1952
rect 17931 1903 17973 1912
rect 18315 1952 18357 1961
rect 18315 1912 18316 1952
rect 18356 1912 18357 1952
rect 18315 1903 18357 1912
rect 18987 1952 19029 1961
rect 18987 1912 18988 1952
rect 19028 1912 19029 1952
rect 18987 1903 19029 1912
rect 19371 1952 19413 1961
rect 19371 1912 19372 1952
rect 19412 1912 19413 1952
rect 19371 1903 19413 1912
rect 19755 1952 19797 1961
rect 19755 1912 19756 1952
rect 19796 1912 19797 1952
rect 19755 1903 19797 1912
rect 20139 1952 20181 1961
rect 20139 1912 20140 1952
rect 20180 1912 20181 1952
rect 20139 1903 20181 1912
rect 18171 1784 18213 1793
rect 18171 1744 18172 1784
rect 18212 1744 18213 1784
rect 18171 1735 18213 1744
rect 19227 1784 19269 1793
rect 19227 1744 19228 1784
rect 19268 1744 19269 1784
rect 19227 1735 19269 1744
rect 13179 1700 13221 1709
rect 13179 1660 13180 1700
rect 13220 1660 13221 1700
rect 13179 1651 13221 1660
rect 15579 1700 15621 1709
rect 15579 1660 15580 1700
rect 15620 1660 15621 1700
rect 15579 1651 15621 1660
rect 19611 1700 19653 1709
rect 19611 1660 19612 1700
rect 19652 1660 19653 1700
rect 19611 1651 19653 1660
rect 1152 1532 20452 1556
rect 1152 1492 4928 1532
rect 4968 1492 5010 1532
rect 5050 1492 5092 1532
rect 5132 1492 5174 1532
rect 5214 1492 5256 1532
rect 5296 1492 20048 1532
rect 20088 1492 20130 1532
rect 20170 1492 20212 1532
rect 20252 1492 20294 1532
rect 20334 1492 20376 1532
rect 20416 1492 20452 1532
rect 1152 1468 20452 1492
<< via1 >>
rect 3688 9808 3728 9848
rect 3770 9808 3810 9848
rect 3852 9808 3892 9848
rect 3934 9808 3974 9848
rect 4016 9808 4056 9848
rect 18808 9808 18848 9848
rect 18890 9808 18930 9848
rect 18972 9808 19012 9848
rect 19054 9808 19094 9848
rect 19136 9808 19176 9848
rect 1564 9640 1604 9680
rect 2332 9640 2372 9680
rect 3100 9640 3140 9680
rect 3484 9640 3524 9680
rect 3868 9640 3908 9680
rect 5020 9640 5060 9680
rect 5404 9640 5444 9680
rect 5788 9640 5828 9680
rect 6172 9640 6212 9680
rect 6556 9640 6596 9680
rect 6940 9640 6980 9680
rect 7708 9640 7748 9680
rect 8188 9640 8228 9680
rect 8572 9640 8612 9680
rect 8956 9640 8996 9680
rect 16156 9640 16196 9680
rect 16540 9640 16580 9680
rect 16924 9640 16964 9680
rect 17692 9640 17732 9680
rect 18460 9640 18500 9680
rect 19612 9640 19652 9680
rect 1948 9556 1988 9596
rect 2716 9556 2756 9596
rect 4252 9556 4292 9596
rect 7324 9556 7364 9596
rect 7804 9556 7844 9596
rect 15676 9556 15716 9596
rect 17308 9556 17348 9596
rect 19228 9556 19268 9596
rect 1324 9472 1364 9512
rect 1708 9472 1748 9512
rect 2092 9472 2132 9512
rect 2476 9472 2516 9512
rect 2860 9472 2900 9512
rect 3244 9472 3284 9512
rect 3628 9472 3668 9512
rect 4012 9472 4052 9512
rect 4396 9472 4436 9512
rect 4636 9472 4676 9512
rect 4780 9472 4820 9512
rect 5164 9472 5204 9512
rect 5548 9472 5588 9512
rect 5932 9472 5972 9512
rect 6316 9472 6356 9512
rect 6700 9472 6740 9512
rect 7084 9472 7124 9512
rect 7468 9472 7508 9512
rect 8044 9472 8084 9512
rect 8428 9472 8468 9512
rect 8812 9472 8852 9512
rect 9196 9472 9236 9512
rect 11884 9472 11924 9512
rect 12844 9472 12884 9512
rect 14572 9472 14612 9512
rect 15052 9472 15092 9512
rect 15436 9472 15476 9512
rect 15820 9472 15860 9512
rect 16396 9472 16436 9512
rect 16780 9472 16820 9512
rect 17164 9472 17204 9512
rect 17548 9472 17588 9512
rect 17932 9472 17972 9512
rect 18316 9472 18356 9512
rect 18700 9472 18740 9512
rect 19084 9472 19124 9512
rect 19468 9472 19508 9512
rect 19852 9472 19892 9512
rect 20236 9472 20276 9512
rect 12124 9304 12164 9344
rect 15292 9304 15332 9344
rect 18076 9304 18116 9344
rect 19996 9304 20036 9344
rect 13084 9220 13124 9260
rect 14812 9220 14852 9260
rect 16060 9220 16100 9260
rect 18844 9220 18884 9260
rect 4928 9052 4968 9092
rect 5010 9052 5050 9092
rect 5092 9052 5132 9092
rect 5174 9052 5214 9092
rect 5256 9052 5296 9092
rect 20048 9052 20088 9092
rect 20130 9052 20170 9092
rect 20212 9052 20252 9092
rect 20294 9052 20334 9092
rect 20376 9052 20416 9092
rect 1468 8884 1508 8924
rect 2716 8884 2756 8924
rect 3196 8884 3236 8924
rect 3580 8884 3620 8924
rect 3964 8884 4004 8924
rect 4348 8884 4388 8924
rect 4732 8884 4772 8924
rect 5116 8884 5156 8924
rect 5884 8884 5924 8924
rect 6268 8884 6308 8924
rect 6652 8884 6692 8924
rect 7036 8884 7076 8924
rect 7420 8884 7460 8924
rect 16060 8884 16100 8924
rect 16924 8884 16964 8924
rect 18460 8884 18500 8924
rect 19612 8884 19652 8924
rect 19996 8884 20036 8924
rect 1948 8800 1988 8840
rect 5500 8800 5540 8840
rect 17308 8800 17348 8840
rect 18844 8800 18884 8840
rect 19516 8800 19556 8840
rect 1228 8632 1268 8672
rect 1612 8632 1652 8672
rect 1852 8632 1892 8672
rect 2188 8632 2228 8672
rect 2572 8632 2612 8672
rect 2956 8632 2996 8672
rect 3436 8632 3476 8672
rect 3820 8632 3860 8672
rect 4204 8632 4244 8672
rect 4588 8632 4628 8672
rect 4972 8632 5012 8672
rect 5356 8632 5396 8672
rect 5740 8632 5780 8672
rect 6124 8632 6164 8672
rect 6508 8632 6548 8672
rect 6892 8632 6932 8672
rect 7276 8632 7316 8672
rect 7660 8632 7700 8672
rect 13324 8632 13364 8672
rect 13564 8632 13604 8672
rect 15820 8632 15860 8672
rect 16204 8632 16244 8672
rect 16588 8632 16628 8672
rect 17164 8632 17204 8672
rect 17548 8632 17588 8672
rect 17692 8632 17732 8672
rect 17932 8632 17972 8672
rect 18076 8632 18116 8672
rect 18316 8632 18356 8672
rect 18700 8632 18740 8672
rect 19084 8632 19124 8672
rect 19276 8632 19316 8672
rect 19852 8632 19892 8672
rect 20236 8632 20276 8672
rect 16828 8548 16868 8588
rect 2332 8464 2372 8504
rect 16444 8464 16484 8504
rect 3688 8296 3728 8336
rect 3770 8296 3810 8336
rect 3852 8296 3892 8336
rect 3934 8296 3974 8336
rect 4016 8296 4056 8336
rect 18808 8296 18848 8336
rect 18890 8296 18930 8336
rect 18972 8296 19012 8336
rect 19054 8296 19094 8336
rect 19136 8296 19176 8336
rect 2044 8128 2084 8168
rect 9916 8128 9956 8168
rect 10300 8128 10340 8168
rect 16924 8128 16964 8168
rect 17308 8128 17348 8168
rect 18076 8128 18116 8168
rect 18556 8128 18596 8168
rect 18940 8044 18980 8084
rect 19612 8044 19652 8084
rect 2284 7960 2324 8000
rect 10156 7960 10196 8000
rect 10540 7960 10580 8000
rect 16300 7960 16340 8000
rect 16684 7960 16724 8000
rect 17068 7960 17108 8000
rect 17452 7960 17492 8000
rect 17836 7960 17876 8000
rect 18412 7960 18452 8000
rect 18796 7960 18836 8000
rect 19180 7960 19220 8000
rect 19372 7960 19412 8000
rect 19756 7960 19796 8000
rect 20140 7960 20180 8000
rect 16540 7708 16580 7748
rect 17692 7708 17732 7748
rect 18172 7708 18212 7748
rect 19996 7708 20036 7748
rect 20380 7708 20420 7748
rect 4928 7540 4968 7580
rect 5010 7540 5050 7580
rect 5092 7540 5132 7580
rect 5174 7540 5214 7580
rect 5256 7540 5296 7580
rect 20048 7540 20088 7580
rect 20130 7540 20170 7580
rect 20212 7540 20252 7580
rect 20294 7540 20334 7580
rect 20376 7540 20416 7580
rect 5884 7372 5924 7412
rect 13948 7372 13988 7412
rect 18556 7372 18596 7412
rect 16060 7288 16100 7328
rect 1948 7120 1988 7160
rect 2188 7120 2228 7160
rect 4348 7120 4388 7160
rect 4588 7120 4628 7160
rect 5212 7120 5252 7160
rect 5452 7120 5492 7160
rect 5644 7120 5684 7160
rect 10156 7120 10196 7160
rect 10300 7120 10340 7160
rect 10540 7120 10580 7160
rect 11836 7120 11876 7160
rect 12076 7120 12116 7160
rect 12460 7120 12500 7160
rect 13564 7120 13604 7160
rect 13804 7120 13844 7160
rect 14188 7120 14228 7160
rect 15388 7120 15428 7160
rect 15628 7120 15668 7160
rect 16300 7120 16340 7160
rect 16876 7120 16916 7160
rect 17260 7120 17300 7160
rect 17548 7120 17588 7160
rect 17788 7120 17828 7160
rect 18124 7120 18164 7160
rect 18316 7120 18356 7160
rect 18700 7120 18740 7160
rect 19084 7120 19124 7160
rect 19660 7120 19700 7160
rect 20140 7120 20180 7160
rect 9916 7036 9956 7076
rect 19324 7036 19364 7076
rect 12220 6952 12260 6992
rect 16636 6952 16676 6992
rect 17020 6952 17060 6992
rect 17884 6952 17924 6992
rect 18940 6952 18980 6992
rect 19420 6952 19460 6992
rect 20380 6952 20420 6992
rect 3688 6784 3728 6824
rect 3770 6784 3810 6824
rect 3852 6784 3892 6824
rect 3934 6784 3974 6824
rect 4016 6784 4056 6824
rect 18808 6784 18848 6824
rect 18890 6784 18930 6824
rect 18972 6784 19012 6824
rect 19054 6784 19094 6824
rect 19136 6784 19176 6824
rect 12700 6616 12740 6656
rect 18652 6616 18692 6656
rect 19036 6616 19076 6656
rect 19420 6616 19460 6656
rect 20380 6616 20420 6656
rect 3340 6448 3380 6488
rect 4396 6448 4436 6488
rect 9148 6448 9188 6488
rect 9388 6448 9428 6488
rect 12940 6448 12980 6488
rect 13324 6448 13364 6488
rect 14668 6448 14708 6488
rect 14908 6448 14948 6488
rect 18412 6448 18452 6488
rect 18796 6448 18836 6488
rect 19180 6448 19220 6488
rect 19756 6448 19796 6488
rect 20140 6448 20180 6488
rect 3580 6280 3620 6320
rect 13084 6280 13124 6320
rect 4636 6196 4676 6236
rect 19516 6196 19556 6236
rect 4928 6028 4968 6068
rect 5010 6028 5050 6068
rect 5092 6028 5132 6068
rect 5174 6028 5214 6068
rect 5256 6028 5296 6068
rect 20048 6028 20088 6068
rect 20130 6028 20170 6068
rect 20212 6028 20252 6068
rect 20294 6028 20334 6068
rect 20376 6028 20416 6068
rect 19132 5860 19172 5900
rect 19996 5860 20036 5900
rect 12316 5776 12356 5816
rect 3196 5608 3236 5648
rect 3436 5608 3476 5648
rect 4780 5608 4820 5648
rect 5836 5608 5876 5648
rect 8284 5608 8324 5648
rect 8524 5608 8564 5648
rect 9292 5608 9332 5648
rect 10636 5608 10676 5648
rect 11020 5608 11060 5648
rect 12076 5608 12116 5648
rect 14956 5608 14996 5648
rect 15196 5608 15236 5648
rect 18220 5608 18260 5648
rect 18796 5608 18836 5648
rect 19372 5608 19412 5648
rect 19756 5608 19796 5648
rect 20140 5608 20180 5648
rect 20380 5608 20420 5648
rect 4540 5524 4580 5564
rect 19036 5524 19076 5564
rect 5596 5440 5636 5480
rect 9532 5440 9572 5480
rect 10876 5440 10916 5480
rect 11260 5440 11300 5480
rect 17980 5440 18020 5480
rect 3688 5272 3728 5312
rect 3770 5272 3810 5312
rect 3852 5272 3892 5312
rect 3934 5272 3974 5312
rect 4016 5272 4056 5312
rect 18808 5272 18848 5312
rect 18890 5272 18930 5312
rect 18972 5272 19012 5312
rect 19054 5272 19094 5312
rect 19136 5272 19176 5312
rect 16252 5104 16292 5144
rect 19996 5104 20036 5144
rect 7036 5020 7076 5060
rect 7612 5020 7652 5060
rect 20380 5020 20420 5060
rect 3724 4936 3764 4976
rect 5164 4936 5204 4976
rect 6652 4936 6692 4976
rect 6892 4936 6932 4976
rect 7276 4936 7316 4976
rect 7852 4936 7892 4976
rect 8092 4936 8132 4976
rect 8332 4936 8372 4976
rect 13804 4936 13844 4976
rect 16012 4936 16052 4976
rect 18700 4936 18740 4976
rect 19036 4936 19076 4976
rect 19276 4936 19316 4976
rect 19756 4936 19796 4976
rect 20140 4936 20180 4976
rect 3964 4768 4004 4808
rect 5404 4684 5444 4724
rect 14044 4684 14084 4724
rect 18940 4684 18980 4724
rect 4928 4516 4968 4556
rect 5010 4516 5050 4556
rect 5092 4516 5132 4556
rect 5174 4516 5214 4556
rect 5256 4516 5296 4556
rect 20048 4516 20088 4556
rect 20130 4516 20170 4556
rect 20212 4516 20252 4556
rect 20294 4516 20334 4556
rect 20376 4516 20416 4556
rect 12124 4264 12164 4304
rect 15388 4264 15428 4304
rect 19132 4264 19172 4304
rect 20380 4264 20420 4304
rect 3868 4096 3908 4136
rect 4108 4096 4148 4136
rect 11884 4096 11924 4136
rect 15148 4096 15188 4136
rect 18796 4096 18836 4136
rect 19372 4096 19412 4136
rect 19603 4096 19643 4136
rect 20140 4096 20180 4136
rect 19036 4012 19076 4052
rect 19804 3928 19844 3968
rect 3688 3760 3728 3800
rect 3770 3760 3810 3800
rect 3852 3760 3892 3800
rect 3934 3760 3974 3800
rect 4016 3760 4056 3800
rect 18808 3760 18848 3800
rect 18890 3760 18930 3800
rect 18972 3760 19012 3800
rect 19054 3760 19094 3800
rect 19136 3760 19176 3800
rect 9148 3592 9188 3632
rect 10972 3592 11012 3632
rect 13660 3592 13700 3632
rect 14044 3592 14084 3632
rect 16828 3592 16868 3632
rect 20380 3592 20420 3632
rect 1900 3424 1940 3464
rect 6316 3424 6356 3464
rect 8524 3424 8564 3464
rect 8908 3424 8948 3464
rect 9964 3424 10004 3464
rect 10732 3424 10772 3464
rect 12076 3424 12116 3464
rect 13420 3424 13460 3464
rect 13804 3424 13844 3464
rect 14956 3424 14996 3464
rect 16588 3424 16628 3464
rect 16972 3424 17012 3464
rect 19372 3424 19412 3464
rect 19795 3424 19835 3464
rect 20140 3424 20180 3464
rect 2140 3256 2180 3296
rect 8764 3256 8804 3296
rect 19612 3256 19652 3296
rect 6556 3172 6596 3212
rect 10204 3172 10244 3212
rect 12316 3172 12356 3212
rect 15196 3172 15236 3212
rect 17212 3172 17252 3212
rect 19996 3172 20036 3212
rect 4928 3004 4968 3044
rect 5010 3004 5050 3044
rect 5092 3004 5132 3044
rect 5174 3004 5214 3044
rect 5256 3004 5296 3044
rect 20048 3004 20088 3044
rect 20130 3004 20170 3044
rect 20212 3004 20252 3044
rect 20294 3004 20334 3044
rect 20376 3004 20416 3044
rect 18844 2836 18884 2876
rect 19996 2836 20036 2876
rect 20380 2836 20420 2876
rect 6604 2584 6644 2624
rect 17164 2584 17204 2624
rect 18124 2584 18164 2624
rect 18604 2584 18644 2624
rect 18988 2584 19028 2624
rect 19372 2584 19412 2624
rect 19756 2584 19796 2624
rect 20140 2584 20180 2624
rect 19228 2500 19268 2540
rect 6844 2416 6884 2456
rect 17404 2416 17444 2456
rect 18364 2416 18404 2456
rect 19612 2416 19652 2456
rect 3688 2248 3728 2288
rect 3770 2248 3810 2288
rect 3852 2248 3892 2288
rect 3934 2248 3974 2288
rect 4016 2248 4056 2288
rect 18808 2248 18848 2288
rect 18890 2248 18930 2288
rect 18972 2248 19012 2288
rect 19054 2248 19094 2288
rect 19136 2248 19176 2288
rect 19996 2080 20036 2120
rect 18556 1996 18596 2036
rect 20380 1996 20420 2036
rect 12940 1912 12980 1952
rect 15340 1912 15380 1952
rect 17932 1912 17972 1952
rect 18316 1912 18356 1952
rect 18988 1912 19028 1952
rect 19372 1912 19412 1952
rect 19756 1912 19796 1952
rect 20140 1912 20180 1952
rect 18172 1744 18212 1784
rect 19228 1744 19268 1784
rect 13180 1660 13220 1700
rect 15580 1660 15620 1700
rect 19612 1660 19652 1700
rect 4928 1492 4968 1532
rect 5010 1492 5050 1532
rect 5092 1492 5132 1532
rect 5174 1492 5214 1532
rect 5256 1492 5296 1532
rect 20048 1492 20088 1532
rect 20130 1492 20170 1532
rect 20212 1492 20252 1532
rect 20294 1492 20334 1532
rect 20376 1492 20416 1532
<< metal2 >>
rect 0 11024 90 11044
rect 21510 11024 21600 11044
rect 0 10984 364 11024
rect 404 10984 413 11024
rect 20707 10984 20716 11024
rect 20756 10984 21600 11024
rect 0 10964 90 10984
rect 21510 10964 21600 10984
rect 0 10688 90 10708
rect 21510 10688 21600 10708
rect 0 10648 652 10688
rect 692 10648 701 10688
rect 20515 10648 20524 10688
rect 20564 10648 21600 10688
rect 0 10628 90 10648
rect 21510 10628 21600 10648
rect 0 10352 90 10372
rect 21510 10352 21600 10372
rect 0 10312 268 10352
rect 308 10312 317 10352
rect 20140 10312 21600 10352
rect 0 10292 90 10312
rect 2275 10060 2284 10100
rect 2324 10060 9292 10100
rect 9332 10060 9341 10100
rect 12940 10060 18220 10100
rect 18260 10060 18269 10100
rect 18883 10060 18892 10100
rect 18932 10060 19948 10100
rect 19988 10060 19997 10100
rect 0 10016 90 10036
rect 12940 10016 12980 10060
rect 20140 10016 20180 10312
rect 21510 10292 21600 10312
rect 21510 10016 21600 10036
rect 0 9976 2668 10016
rect 2708 9976 2717 10016
rect 3715 9976 3724 10016
rect 3764 9976 3773 10016
rect 6115 9976 6124 10016
rect 6164 9976 12980 10016
rect 16099 9976 16108 10016
rect 16148 9976 20180 10016
rect 20236 9976 21600 10016
rect 0 9956 90 9976
rect 3724 9932 3764 9976
rect 20236 9932 20276 9976
rect 21510 9956 21600 9976
rect 3532 9892 3764 9932
rect 4780 9892 9868 9932
rect 9908 9892 9917 9932
rect 15235 9892 15244 9932
rect 15284 9892 16820 9932
rect 17827 9892 17836 9932
rect 17876 9892 19268 9932
rect 19363 9892 19372 9932
rect 19412 9892 20276 9932
rect 172 9808 3436 9848
rect 3476 9808 3485 9848
rect 0 9680 90 9700
rect 172 9680 212 9808
rect 1996 9724 2380 9764
rect 2420 9724 2429 9764
rect 2572 9724 2764 9764
rect 2804 9724 2813 9764
rect 1996 9680 2036 9724
rect 2572 9680 2612 9724
rect 3532 9680 3572 9892
rect 3679 9808 3688 9848
rect 3728 9808 3770 9848
rect 3810 9808 3852 9848
rect 3892 9808 3934 9848
rect 3974 9808 4016 9848
rect 4056 9808 4065 9848
rect 0 9640 212 9680
rect 1555 9640 1564 9680
rect 1604 9640 2036 9680
rect 2323 9640 2332 9680
rect 2372 9640 2612 9680
rect 2764 9640 2956 9680
rect 2996 9640 3005 9680
rect 3091 9640 3100 9680
rect 3140 9640 3340 9680
rect 3380 9640 3389 9680
rect 3475 9640 3484 9680
rect 3524 9640 3572 9680
rect 3859 9640 3868 9680
rect 3908 9640 4204 9680
rect 4244 9640 4253 9680
rect 0 9620 90 9640
rect 2764 9596 2804 9640
rect 1939 9556 1948 9596
rect 1988 9556 2572 9596
rect 2612 9556 2621 9596
rect 2707 9556 2716 9596
rect 2756 9556 2804 9596
rect 2860 9556 3244 9596
rect 3284 9556 3293 9596
rect 3340 9556 3724 9596
rect 3764 9556 3773 9596
rect 4243 9556 4252 9596
rect 4292 9556 4492 9596
rect 4532 9556 4541 9596
rect 2860 9512 2900 9556
rect 3340 9512 3380 9556
rect 4780 9512 4820 9892
rect 16780 9848 16820 9892
rect 19228 9848 19268 9892
rect 4876 9808 15724 9848
rect 15764 9808 15773 9848
rect 16003 9808 16012 9848
rect 16052 9808 16724 9848
rect 16780 9808 18412 9848
rect 18452 9808 18461 9848
rect 18799 9808 18808 9848
rect 18848 9808 18890 9848
rect 18930 9808 18972 9848
rect 19012 9808 19054 9848
rect 19094 9808 19136 9848
rect 19176 9808 19185 9848
rect 19228 9808 19796 9848
rect 4876 9512 4916 9808
rect 8428 9724 10732 9764
rect 10772 9724 10781 9764
rect 12259 9724 12268 9764
rect 12308 9724 12980 9764
rect 15811 9724 15820 9764
rect 15860 9724 16340 9764
rect 5011 9640 5020 9680
rect 5060 9640 5260 9680
rect 5300 9640 5309 9680
rect 5395 9640 5404 9680
rect 5444 9640 5644 9680
rect 5684 9640 5693 9680
rect 5779 9640 5788 9680
rect 5828 9640 6028 9680
rect 6068 9640 6077 9680
rect 6163 9640 6172 9680
rect 6212 9640 6412 9680
rect 6452 9640 6461 9680
rect 6547 9640 6556 9680
rect 6596 9640 6796 9680
rect 6836 9640 6845 9680
rect 6931 9640 6940 9680
rect 6980 9640 7180 9680
rect 7220 9640 7229 9680
rect 7625 9640 7708 9680
rect 7748 9640 7756 9680
rect 7796 9640 7805 9680
rect 8131 9640 8140 9680
rect 8180 9640 8188 9680
rect 8228 9640 8311 9680
rect 7315 9556 7324 9596
rect 7364 9556 7564 9596
rect 7604 9556 7613 9596
rect 7795 9556 7804 9596
rect 7844 9556 7948 9596
rect 7988 9556 7997 9596
rect 8428 9512 8468 9724
rect 12940 9680 12980 9724
rect 16300 9680 16340 9724
rect 16684 9680 16724 9808
rect 16771 9724 16780 9764
rect 16820 9724 17300 9764
rect 17347 9724 17356 9764
rect 17396 9724 17972 9764
rect 18307 9724 18316 9764
rect 18356 9724 19028 9764
rect 17260 9680 17300 9724
rect 17932 9680 17972 9724
rect 18988 9680 19028 9724
rect 19756 9680 19796 9808
rect 21510 9680 21600 9700
rect 8515 9640 8524 9680
rect 8564 9640 8572 9680
rect 8612 9640 8695 9680
rect 8899 9640 8908 9680
rect 8948 9640 8956 9680
rect 8996 9640 9079 9680
rect 9187 9640 9196 9680
rect 9236 9640 12884 9680
rect 12940 9640 15572 9680
rect 15619 9640 15628 9680
rect 15668 9640 16156 9680
rect 16196 9640 16205 9680
rect 16300 9640 16540 9680
rect 16580 9640 16589 9680
rect 16684 9640 16924 9680
rect 16964 9640 16973 9680
rect 17260 9640 17692 9680
rect 17732 9640 17741 9680
rect 17932 9640 18460 9680
rect 18500 9640 18509 9680
rect 18988 9640 19612 9680
rect 19652 9640 19661 9680
rect 19756 9640 21600 9680
rect 8812 9556 11500 9596
rect 11540 9556 11549 9596
rect 8812 9512 8852 9556
rect 12844 9512 12884 9640
rect 12940 9556 15476 9596
rect 1315 9472 1324 9512
rect 1364 9472 1556 9512
rect 1699 9472 1708 9512
rect 1748 9472 1757 9512
rect 1891 9472 1900 9512
rect 1940 9472 2092 9512
rect 2132 9472 2141 9512
rect 2467 9472 2476 9512
rect 2516 9472 2525 9512
rect 2851 9472 2860 9512
rect 2900 9472 2909 9512
rect 3235 9472 3244 9512
rect 3284 9472 3380 9512
rect 3497 9472 3628 9512
rect 3668 9472 3677 9512
rect 4003 9472 4012 9512
rect 4052 9472 4061 9512
rect 4265 9472 4396 9512
rect 4436 9472 4445 9512
rect 4627 9472 4636 9512
rect 4676 9472 4724 9512
rect 4771 9472 4780 9512
rect 4820 9472 4829 9512
rect 4876 9472 5164 9512
rect 5204 9472 5213 9512
rect 5417 9472 5548 9512
rect 5588 9472 5597 9512
rect 5923 9472 5932 9512
rect 5972 9472 5981 9512
rect 6185 9472 6316 9512
rect 6356 9472 6365 9512
rect 6569 9472 6700 9512
rect 6740 9472 6749 9512
rect 7075 9472 7084 9512
rect 7124 9472 7255 9512
rect 7459 9472 7468 9512
rect 7508 9472 7639 9512
rect 8035 9472 8044 9512
rect 8084 9472 8093 9512
rect 8419 9472 8428 9512
rect 8468 9472 8477 9512
rect 8803 9472 8812 9512
rect 8852 9472 8861 9512
rect 9187 9472 9196 9512
rect 9236 9472 11308 9512
rect 11348 9472 11357 9512
rect 11875 9472 11884 9512
rect 11924 9472 11933 9512
rect 12835 9472 12844 9512
rect 12884 9472 12893 9512
rect 0 9344 90 9364
rect 0 9304 76 9344
rect 116 9304 125 9344
rect 0 9284 90 9304
rect 1516 9176 1556 9472
rect 1708 9260 1748 9472
rect 2476 9428 2516 9472
rect 4012 9428 4052 9472
rect 2476 9388 3052 9428
rect 3092 9388 3101 9428
rect 3331 9388 3340 9428
rect 3380 9388 4052 9428
rect 4684 9428 4724 9472
rect 5932 9428 5972 9472
rect 8044 9428 8084 9472
rect 4684 9388 4876 9428
rect 4916 9388 4925 9428
rect 5932 9388 6508 9428
rect 6548 9388 6557 9428
rect 8044 9388 11788 9428
rect 11828 9388 11837 9428
rect 11884 9344 11924 9472
rect 12940 9428 12980 9556
rect 15436 9512 15476 9556
rect 14441 9472 14572 9512
rect 14612 9472 14621 9512
rect 15043 9472 15052 9512
rect 15092 9472 15101 9512
rect 15427 9472 15436 9512
rect 15476 9472 15485 9512
rect 2083 9304 2092 9344
rect 2132 9304 11924 9344
rect 11980 9388 12980 9428
rect 15052 9428 15092 9472
rect 15532 9428 15572 9640
rect 21510 9620 21600 9640
rect 15667 9556 15676 9596
rect 15716 9556 16204 9596
rect 16244 9556 16253 9596
rect 16483 9556 16492 9596
rect 16532 9556 17308 9596
rect 17348 9556 17357 9596
rect 17923 9556 17932 9596
rect 17972 9556 19228 9596
rect 19268 9556 19277 9596
rect 15689 9472 15820 9512
rect 15860 9472 15869 9512
rect 16265 9472 16396 9512
rect 16436 9472 16445 9512
rect 16649 9472 16780 9512
rect 16820 9472 16829 9512
rect 17033 9472 17068 9512
rect 17108 9472 17164 9512
rect 17204 9472 17213 9512
rect 17347 9472 17356 9512
rect 17396 9472 17548 9512
rect 17588 9472 17597 9512
rect 17923 9472 17932 9512
rect 17972 9472 17981 9512
rect 18307 9472 18316 9512
rect 18356 9472 18365 9512
rect 18691 9472 18700 9512
rect 18740 9472 18796 9512
rect 18836 9472 18871 9512
rect 18953 9472 19084 9512
rect 19124 9472 19133 9512
rect 19459 9472 19468 9512
rect 19508 9472 19564 9512
rect 19604 9472 19639 9512
rect 19721 9472 19756 9512
rect 19796 9472 19852 9512
rect 19892 9472 19901 9512
rect 20105 9472 20236 9512
rect 20276 9472 20285 9512
rect 17932 9428 17972 9472
rect 18316 9428 18356 9472
rect 15052 9388 15436 9428
rect 15476 9388 15485 9428
rect 15532 9388 17972 9428
rect 18019 9388 18028 9428
rect 18068 9388 18356 9428
rect 18595 9388 18604 9428
rect 18644 9388 20180 9428
rect 11980 9260 12020 9388
rect 20140 9344 20180 9388
rect 21510 9344 21600 9364
rect 12115 9304 12124 9344
rect 12164 9304 14956 9344
rect 14996 9304 15005 9344
rect 15283 9304 15292 9344
rect 15332 9304 17108 9344
rect 17155 9304 17164 9344
rect 17204 9304 18076 9344
rect 18116 9304 18125 9344
rect 18211 9304 18220 9344
rect 18260 9304 19996 9344
rect 20036 9304 20045 9344
rect 20140 9304 21600 9344
rect 17068 9260 17108 9304
rect 21510 9284 21600 9304
rect 1708 9220 2572 9260
rect 2612 9220 2621 9260
rect 4387 9220 4396 9260
rect 4436 9220 10348 9260
rect 10388 9220 10397 9260
rect 11875 9220 11884 9260
rect 11924 9220 12020 9260
rect 13075 9220 13084 9260
rect 13124 9220 14708 9260
rect 14803 9220 14812 9260
rect 14852 9220 15956 9260
rect 16051 9220 16060 9260
rect 16100 9220 17012 9260
rect 17068 9220 17492 9260
rect 17539 9220 17548 9260
rect 17588 9220 18844 9260
rect 18884 9220 18893 9260
rect 18979 9220 18988 9260
rect 19028 9220 20908 9260
rect 20948 9220 20957 9260
rect 14668 9176 14708 9220
rect 15916 9176 15956 9220
rect 16972 9176 17012 9220
rect 17452 9176 17492 9220
rect 1516 9136 4780 9176
rect 4820 9136 4829 9176
rect 6307 9136 6316 9176
rect 6356 9136 14092 9176
rect 14132 9136 14141 9176
rect 14668 9136 14764 9176
rect 14804 9136 14813 9176
rect 15916 9136 16876 9176
rect 16916 9136 16925 9176
rect 16972 9136 17260 9176
rect 17300 9136 17309 9176
rect 17452 9136 20524 9176
rect 20564 9136 20573 9176
rect 1603 9052 1612 9092
rect 1652 9052 4396 9092
rect 4436 9052 4445 9092
rect 4919 9052 4928 9092
rect 4968 9052 5010 9092
rect 5050 9052 5092 9092
rect 5132 9052 5174 9092
rect 5214 9052 5256 9092
rect 5296 9052 5305 9092
rect 6691 9052 6700 9092
rect 6740 9052 10060 9092
rect 10100 9052 10109 9092
rect 15427 9052 15436 9092
rect 15476 9052 17684 9092
rect 18019 9052 18028 9092
rect 18068 9052 19372 9092
rect 19412 9052 19421 9092
rect 20039 9052 20048 9092
rect 20088 9052 20130 9092
rect 20170 9052 20212 9092
rect 20252 9052 20294 9092
rect 20334 9052 20376 9092
rect 20416 9052 20425 9092
rect 0 9008 90 9028
rect 0 8968 4204 9008
rect 4244 8968 4253 9008
rect 5740 8968 10252 9008
rect 10292 8968 10301 9008
rect 12835 8968 12844 9008
rect 12884 8968 17548 9008
rect 17588 8968 17597 9008
rect 0 8948 90 8968
rect 1459 8884 1468 8924
rect 1508 8884 1804 8924
rect 1844 8884 1853 8924
rect 2563 8884 2572 8924
rect 2612 8884 2716 8924
rect 2756 8884 2765 8924
rect 3139 8884 3148 8924
rect 3188 8884 3196 8924
rect 3236 8884 3319 8924
rect 3523 8884 3532 8924
rect 3572 8884 3580 8924
rect 3620 8884 3703 8924
rect 3955 8884 3964 8924
rect 4004 8884 4108 8924
rect 4148 8884 4157 8924
rect 4291 8884 4300 8924
rect 4340 8884 4348 8924
rect 4388 8884 4471 8924
rect 4675 8884 4684 8924
rect 4724 8884 4732 8924
rect 4772 8884 4855 8924
rect 5107 8884 5116 8924
rect 5156 8884 5356 8924
rect 5396 8884 5405 8924
rect 1228 8800 1948 8840
rect 1988 8800 1997 8840
rect 2956 8800 4820 8840
rect 5443 8800 5452 8840
rect 5492 8800 5500 8840
rect 5540 8800 5623 8840
rect 0 8672 90 8692
rect 1228 8672 1268 8800
rect 1996 8716 2188 8756
rect 2228 8716 2237 8756
rect 1996 8672 2036 8716
rect 2956 8672 2996 8800
rect 3139 8716 3148 8756
rect 3188 8716 3724 8756
rect 3764 8716 3773 8756
rect 4780 8672 4820 8800
rect 4972 8716 5644 8756
rect 5684 8716 5693 8756
rect 4972 8672 5012 8716
rect 5740 8672 5780 8968
rect 5827 8884 5836 8924
rect 5876 8884 5884 8924
rect 5924 8884 6007 8924
rect 6211 8884 6220 8924
rect 6260 8884 6268 8924
rect 6308 8884 6391 8924
rect 6595 8884 6604 8924
rect 6644 8884 6652 8924
rect 6692 8884 6775 8924
rect 6979 8884 6988 8924
rect 7028 8884 7036 8924
rect 7076 8884 7159 8924
rect 7363 8884 7372 8924
rect 7412 8884 7420 8924
rect 7460 8884 7543 8924
rect 7651 8884 7660 8924
rect 7700 8884 9100 8924
rect 9140 8884 9149 8924
rect 12556 8884 14188 8924
rect 14228 8884 14237 8924
rect 14755 8884 14764 8924
rect 14804 8884 15340 8924
rect 15380 8884 15389 8924
rect 15977 8884 16060 8924
rect 16100 8884 16108 8924
rect 16148 8884 16157 8924
rect 16579 8884 16588 8924
rect 16628 8884 16924 8924
rect 16964 8884 16973 8924
rect 17251 8884 17260 8924
rect 17300 8884 17452 8924
rect 17492 8884 17501 8924
rect 12556 8840 12596 8884
rect 17644 8840 17684 9052
rect 21510 9008 21600 9028
rect 18307 8968 18316 9008
rect 18356 8968 18644 9008
rect 19555 8968 19564 9008
rect 19604 8968 21600 9008
rect 18604 8924 18644 8968
rect 21510 8948 21600 8968
rect 17731 8884 17740 8924
rect 17780 8884 18460 8924
rect 18500 8884 18509 8924
rect 18604 8884 19612 8924
rect 19652 8884 19661 8924
rect 19939 8884 19948 8924
rect 19988 8884 19996 8924
rect 20036 8884 20119 8924
rect 7276 8800 12596 8840
rect 12940 8800 14380 8840
rect 14420 8800 14429 8840
rect 16963 8800 16972 8840
rect 17012 8800 17308 8840
rect 17348 8800 17357 8840
rect 17644 8800 17780 8840
rect 18115 8800 18124 8840
rect 18164 8800 18844 8840
rect 18884 8800 18893 8840
rect 19507 8800 19516 8840
rect 19556 8800 20620 8840
rect 20660 8800 20669 8840
rect 6508 8716 7180 8756
rect 7220 8716 7229 8756
rect 6508 8672 6548 8716
rect 7276 8672 7316 8800
rect 7372 8716 10828 8756
rect 10868 8716 10877 8756
rect 0 8632 940 8672
rect 980 8632 989 8672
rect 1219 8632 1228 8672
rect 1268 8632 1277 8672
rect 1481 8632 1612 8672
rect 1652 8632 1661 8672
rect 1843 8632 1852 8672
rect 1892 8632 2036 8672
rect 2179 8632 2188 8672
rect 2228 8632 2284 8672
rect 2324 8632 2359 8672
rect 2563 8632 2572 8672
rect 2612 8632 2900 8672
rect 2947 8632 2956 8672
rect 2996 8632 3005 8672
rect 3305 8632 3436 8672
rect 3476 8632 3485 8672
rect 3811 8632 3820 8672
rect 3860 8632 4148 8672
rect 4195 8632 4204 8672
rect 4244 8632 4300 8672
rect 4340 8632 4375 8672
rect 4457 8632 4588 8672
rect 4628 8632 4637 8672
rect 4780 8632 4916 8672
rect 4963 8632 4972 8672
rect 5012 8632 5021 8672
rect 5225 8632 5356 8672
rect 5396 8632 5405 8672
rect 5731 8632 5740 8672
rect 5780 8632 5789 8672
rect 5993 8632 6124 8672
rect 6164 8632 6173 8672
rect 6499 8632 6508 8672
rect 6548 8632 6557 8672
rect 6883 8632 6892 8672
rect 6932 8632 6988 8672
rect 7028 8632 7063 8672
rect 7267 8632 7276 8672
rect 7316 8632 7325 8672
rect 0 8612 90 8632
rect 2860 8504 2900 8632
rect 4108 8588 4148 8632
rect 4876 8588 4916 8632
rect 7372 8588 7412 8716
rect 12940 8672 12980 8800
rect 17740 8756 17780 8800
rect 13324 8716 15436 8756
rect 15476 8716 15485 8756
rect 15820 8716 16588 8756
rect 16628 8716 16637 8756
rect 16867 8716 16876 8756
rect 16916 8716 17684 8756
rect 17740 8716 18068 8756
rect 18403 8716 18412 8756
rect 18452 8716 19412 8756
rect 19843 8716 19852 8756
rect 19892 8716 20276 8756
rect 13324 8672 13364 8716
rect 15820 8672 15860 8716
rect 17644 8672 17684 8716
rect 18028 8672 18068 8716
rect 19372 8672 19412 8716
rect 20236 8672 20276 8716
rect 21510 8672 21600 8692
rect 7651 8632 7660 8672
rect 7700 8632 12980 8672
rect 13315 8632 13324 8672
rect 13364 8632 13373 8672
rect 13555 8632 13564 8672
rect 13604 8632 15628 8672
rect 15668 8632 15677 8672
rect 15811 8632 15820 8672
rect 15860 8632 15869 8672
rect 16073 8632 16204 8672
rect 16244 8632 16253 8672
rect 16457 8632 16492 8672
rect 16532 8632 16588 8672
rect 16628 8632 16637 8672
rect 16963 8632 16972 8672
rect 17012 8632 17164 8672
rect 17204 8632 17213 8672
rect 17417 8632 17548 8672
rect 17588 8632 17597 8672
rect 17644 8632 17692 8672
rect 17732 8632 17741 8672
rect 17801 8632 17932 8672
rect 17972 8632 17981 8672
rect 18028 8632 18076 8672
rect 18116 8632 18125 8672
rect 18185 8632 18316 8672
rect 18356 8632 18365 8672
rect 18691 8632 18700 8672
rect 18740 8632 18749 8672
rect 18883 8632 18892 8672
rect 18932 8632 19084 8672
rect 19124 8632 19133 8672
rect 19180 8632 19276 8672
rect 19316 8632 19325 8672
rect 19372 8632 19852 8672
rect 19892 8632 19901 8672
rect 20227 8632 20236 8672
rect 20276 8632 20285 8672
rect 20515 8632 20524 8672
rect 20564 8632 21600 8672
rect 18700 8588 18740 8632
rect 19180 8588 19220 8632
rect 21510 8612 21600 8632
rect 4108 8548 4204 8588
rect 4244 8548 4253 8588
rect 4876 8548 7412 8588
rect 16675 8548 16684 8588
rect 16724 8548 16828 8588
rect 16868 8548 16877 8588
rect 17251 8548 17260 8588
rect 17300 8548 18028 8588
rect 18068 8548 18077 8588
rect 18403 8548 18412 8588
rect 18452 8548 18740 8588
rect 19171 8548 19180 8588
rect 19220 8548 19229 8588
rect 2201 8464 2284 8504
rect 2324 8464 2332 8504
rect 2372 8464 2381 8504
rect 2860 8464 7660 8504
rect 7700 8464 7709 8504
rect 16435 8464 16444 8504
rect 16484 8464 16820 8504
rect 16780 8420 16820 8464
rect 17164 8464 18220 8504
rect 18260 8464 18269 8504
rect 16780 8380 17068 8420
rect 17108 8380 17117 8420
rect 0 8336 90 8356
rect 17164 8336 17204 8464
rect 0 8296 1132 8336
rect 1172 8296 1181 8336
rect 3679 8296 3688 8336
rect 3728 8296 3770 8336
rect 3810 8296 3852 8336
rect 3892 8296 3934 8336
rect 3974 8296 4016 8336
rect 4056 8296 4065 8336
rect 16291 8296 16300 8336
rect 16340 8296 17204 8336
rect 17932 8380 19564 8420
rect 19604 8380 19613 8420
rect 0 8276 90 8296
rect 15523 8212 15532 8252
rect 15572 8212 17836 8252
rect 17876 8212 17885 8252
rect 17932 8168 17972 8380
rect 21510 8336 21600 8356
rect 18799 8296 18808 8336
rect 18848 8296 18890 8336
rect 18930 8296 18972 8336
rect 19012 8296 19054 8336
rect 19094 8296 19136 8336
rect 19176 8296 19185 8336
rect 19363 8296 19372 8336
rect 19412 8296 21600 8336
rect 21510 8276 21600 8296
rect 18412 8212 19468 8252
rect 19508 8212 19517 8252
rect 18412 8168 18452 8212
rect 1987 8128 1996 8168
rect 2036 8128 2044 8168
rect 2084 8128 2167 8168
rect 9859 8128 9868 8168
rect 9908 8128 9916 8168
rect 9956 8128 10039 8168
rect 10243 8128 10252 8168
rect 10292 8128 10300 8168
rect 10340 8128 10423 8168
rect 16915 8128 16924 8168
rect 16964 8128 17164 8168
rect 17204 8128 17213 8168
rect 17299 8128 17308 8168
rect 17348 8128 17972 8168
rect 18067 8128 18076 8168
rect 18116 8128 18452 8168
rect 18499 8128 18508 8168
rect 18548 8128 18556 8168
rect 18596 8128 18679 8168
rect 10156 8044 11212 8084
rect 11252 8044 11261 8084
rect 15619 8044 15628 8084
rect 15668 8044 18548 8084
rect 18691 8044 18700 8084
rect 18740 8044 18940 8084
rect 18980 8044 18989 8084
rect 19603 8044 19612 8084
rect 19652 8044 20660 8084
rect 0 8000 90 8020
rect 10156 8000 10196 8044
rect 18508 8000 18548 8044
rect 20620 8000 20660 8044
rect 21510 8000 21600 8020
rect 0 7960 268 8000
rect 308 7960 317 8000
rect 2153 7960 2284 8000
rect 2324 7960 2333 8000
rect 10147 7960 10156 8000
rect 10196 7960 10205 8000
rect 10531 7960 10540 8000
rect 10580 7960 11020 8000
rect 11060 7960 11069 8000
rect 16169 7960 16300 8000
rect 16340 7960 16349 8000
rect 16553 7960 16684 8000
rect 16724 7960 16733 8000
rect 16937 7960 17068 8000
rect 17108 7960 17117 8000
rect 17443 7960 17452 8000
rect 17492 7960 17501 8000
rect 17827 7960 17836 8000
rect 17876 7960 17885 8000
rect 18019 7960 18028 8000
rect 18068 7960 18412 8000
rect 18452 7960 18461 8000
rect 18508 7960 18796 8000
rect 18836 7960 18845 8000
rect 19049 7960 19180 8000
rect 19220 7960 19229 8000
rect 19363 7960 19372 8000
rect 19412 7960 19468 8000
rect 19508 7960 19543 8000
rect 19625 7960 19756 8000
rect 19796 7960 19805 8000
rect 20131 7960 20140 8000
rect 20180 7960 20564 8000
rect 20620 7960 21600 8000
rect 0 7940 90 7960
rect 17452 7832 17492 7960
rect 17836 7916 17876 7960
rect 20524 7916 20564 7960
rect 21510 7940 21600 7960
rect 17836 7876 18316 7916
rect 18356 7876 18365 7916
rect 20524 7876 20812 7916
rect 20852 7876 20861 7916
rect 7267 7792 7276 7832
rect 7316 7792 17260 7832
rect 17300 7792 17309 7832
rect 17452 7792 17932 7832
rect 17972 7792 17981 7832
rect 16531 7708 16540 7748
rect 16580 7708 17588 7748
rect 17683 7708 17692 7748
rect 17732 7708 18068 7748
rect 18115 7708 18124 7748
rect 18164 7708 18172 7748
rect 18212 7708 18295 7748
rect 19987 7708 19996 7748
rect 20036 7708 20045 7748
rect 20371 7708 20380 7748
rect 20420 7708 21004 7748
rect 21044 7708 21053 7748
rect 0 7664 90 7684
rect 0 7624 1324 7664
rect 1364 7624 1373 7664
rect 0 7604 90 7624
rect 4919 7540 4928 7580
rect 4968 7540 5010 7580
rect 5050 7540 5092 7580
rect 5132 7540 5174 7580
rect 5214 7540 5256 7580
rect 5296 7540 5305 7580
rect 17548 7496 17588 7708
rect 18028 7664 18068 7708
rect 19996 7664 20036 7708
rect 21510 7664 21600 7684
rect 18028 7624 19660 7664
rect 19700 7624 19709 7664
rect 19996 7624 21600 7664
rect 21510 7604 21600 7624
rect 20039 7540 20048 7580
rect 20088 7540 20130 7580
rect 20170 7540 20212 7580
rect 20252 7540 20294 7580
rect 20334 7540 20376 7580
rect 20416 7540 20425 7580
rect 15715 7456 15724 7496
rect 15764 7456 17492 7496
rect 17548 7456 20716 7496
rect 20756 7456 20765 7496
rect 17452 7412 17492 7456
rect 5875 7372 5884 7412
rect 5924 7372 7948 7412
rect 7988 7372 7997 7412
rect 11491 7372 11500 7412
rect 11540 7372 13948 7412
rect 13988 7372 13997 7412
rect 14467 7372 14476 7412
rect 14516 7372 17012 7412
rect 17452 7372 18124 7412
rect 18164 7372 18173 7412
rect 18547 7372 18556 7412
rect 18596 7372 19372 7412
rect 19412 7372 19421 7412
rect 0 7328 90 7348
rect 0 7288 556 7328
rect 596 7288 605 7328
rect 4588 7288 8812 7328
rect 8852 7288 8861 7328
rect 13891 7288 13900 7328
rect 13940 7288 15764 7328
rect 16003 7288 16012 7328
rect 16052 7288 16060 7328
rect 16100 7288 16183 7328
rect 0 7268 90 7288
rect 4588 7160 4628 7288
rect 5548 7204 5780 7244
rect 5548 7160 5588 7204
rect 5740 7160 5780 7204
rect 12940 7204 13324 7244
rect 13364 7204 13373 7244
rect 13699 7204 13708 7244
rect 13748 7204 14324 7244
rect 12940 7160 12980 7204
rect 1891 7120 1900 7160
rect 1940 7120 1948 7160
rect 1988 7120 2071 7160
rect 2179 7120 2188 7160
rect 2228 7120 2359 7160
rect 4265 7120 4348 7160
rect 4388 7120 4396 7160
rect 4436 7120 4445 7160
rect 4579 7120 4588 7160
rect 4628 7120 4637 7160
rect 4771 7120 4780 7160
rect 4820 7120 5212 7160
rect 5252 7120 5261 7160
rect 5443 7120 5452 7160
rect 5492 7120 5588 7160
rect 5635 7120 5644 7160
rect 5684 7120 5693 7160
rect 5740 7120 8716 7160
rect 8756 7120 8765 7160
rect 10147 7120 10156 7160
rect 10196 7120 10205 7160
rect 10291 7120 10300 7160
rect 10340 7120 10348 7160
rect 10388 7120 10471 7160
rect 10531 7120 10540 7160
rect 10580 7120 11596 7160
rect 11636 7120 11645 7160
rect 11779 7120 11788 7160
rect 11828 7120 11836 7160
rect 11876 7120 11959 7160
rect 12067 7120 12076 7160
rect 12116 7120 12125 7160
rect 12451 7120 12460 7160
rect 12500 7120 12980 7160
rect 13027 7120 13036 7160
rect 13076 7120 13564 7160
rect 13604 7120 13613 7160
rect 13795 7120 13804 7160
rect 13844 7120 13853 7160
rect 14179 7120 14188 7160
rect 14228 7120 14237 7160
rect 5644 7076 5684 7120
rect 10156 7076 10196 7120
rect 12076 7076 12116 7120
rect 13804 7076 13844 7120
rect 1420 7036 2900 7076
rect 0 6992 90 7012
rect 1420 6992 1460 7036
rect 0 6952 1460 6992
rect 2860 6992 2900 7036
rect 4780 7036 5684 7076
rect 5740 7036 9916 7076
rect 9956 7036 9965 7076
rect 10156 7036 11404 7076
rect 11444 7036 11453 7076
rect 12076 7036 12596 7076
rect 12739 7036 12748 7076
rect 12788 7036 13844 7076
rect 2860 6952 4492 6992
rect 4532 6952 4541 6992
rect 0 6932 90 6952
rect 4780 6824 4820 7036
rect 5740 6992 5780 7036
rect 12556 6992 12596 7036
rect 14188 6992 14228 7120
rect 14284 7076 14324 7204
rect 15724 7160 15764 7288
rect 16972 7160 17012 7372
rect 21510 7328 21600 7348
rect 20995 7288 21004 7328
rect 21044 7288 21600 7328
rect 21510 7268 21600 7288
rect 18403 7204 18412 7244
rect 18452 7204 18932 7244
rect 18892 7160 18932 7204
rect 14371 7120 14380 7160
rect 14420 7120 15388 7160
rect 15428 7120 15437 7160
rect 15619 7120 15628 7160
rect 15668 7120 15677 7160
rect 15724 7120 16300 7160
rect 16340 7120 16349 7160
rect 16483 7120 16492 7160
rect 16532 7120 16876 7160
rect 16916 7120 16925 7160
rect 16972 7120 17260 7160
rect 17300 7120 17309 7160
rect 17443 7120 17452 7160
rect 17492 7120 17548 7160
rect 17588 7120 17623 7160
rect 17731 7120 17740 7160
rect 17780 7120 17788 7160
rect 17828 7120 17911 7160
rect 17993 7120 18124 7160
rect 18164 7120 18173 7160
rect 18307 7120 18316 7160
rect 18356 7120 18365 7160
rect 18691 7120 18700 7160
rect 18740 7120 18836 7160
rect 18892 7120 19084 7160
rect 19124 7120 19133 7160
rect 19529 7120 19660 7160
rect 19700 7120 19709 7160
rect 20131 7120 20140 7160
rect 20180 7120 20189 7160
rect 15628 7076 15668 7120
rect 14284 7036 15668 7076
rect 18316 7076 18356 7120
rect 18316 7036 18700 7076
rect 18740 7036 18749 7076
rect 18796 6992 18836 7120
rect 20140 7076 20180 7120
rect 19315 7036 19324 7076
rect 19364 7036 20180 7076
rect 21510 6992 21600 7012
rect 5347 6952 5356 6992
rect 5396 6952 5780 6992
rect 7459 6952 7468 6992
rect 7508 6952 12220 6992
rect 12260 6952 12269 6992
rect 12556 6952 13132 6992
rect 13172 6952 13181 6992
rect 13516 6952 14228 6992
rect 16204 6952 16636 6992
rect 16676 6952 16685 6992
rect 16963 6952 16972 6992
rect 17012 6952 17020 6992
rect 17060 6952 17143 6992
rect 17251 6952 17260 6992
rect 17300 6952 17884 6992
rect 17924 6952 17933 6992
rect 18019 6952 18028 6992
rect 18068 6952 18836 6992
rect 18931 6952 18940 6992
rect 18980 6952 19276 6992
rect 19316 6952 19325 6992
rect 19372 6952 19420 6992
rect 19460 6952 19469 6992
rect 20371 6952 20380 6992
rect 20420 6952 21600 6992
rect 7843 6868 7852 6908
rect 7892 6868 12788 6908
rect 3679 6784 3688 6824
rect 3728 6784 3770 6824
rect 3810 6784 3852 6824
rect 3892 6784 3934 6824
rect 3974 6784 4016 6824
rect 4056 6784 4065 6824
rect 4291 6784 4300 6824
rect 4340 6784 4820 6824
rect 7939 6784 7948 6824
rect 7988 6784 11884 6824
rect 11924 6784 11933 6824
rect 12748 6740 12788 6868
rect 13516 6824 13556 6952
rect 16204 6824 16244 6952
rect 12931 6784 12940 6824
rect 12980 6784 13556 6824
rect 14179 6784 14188 6824
rect 14228 6784 16244 6824
rect 18799 6784 18808 6824
rect 18848 6784 18890 6824
rect 18930 6784 18972 6824
rect 19012 6784 19054 6824
rect 19094 6784 19136 6824
rect 19176 6784 19185 6824
rect 19372 6740 19412 6952
rect 21510 6932 21600 6952
rect 7075 6700 7084 6740
rect 7124 6700 9908 6740
rect 12748 6700 19412 6740
rect 0 6656 90 6676
rect 9868 6656 9908 6700
rect 21510 6656 21600 6676
rect 0 6616 8908 6656
rect 8948 6616 8957 6656
rect 9868 6616 12700 6656
rect 12740 6616 12749 6656
rect 13027 6616 13036 6656
rect 13076 6616 13516 6656
rect 13556 6616 13565 6656
rect 14083 6616 14092 6656
rect 14132 6616 16972 6656
rect 17012 6616 17021 6656
rect 18403 6616 18412 6656
rect 18452 6616 18461 6656
rect 18595 6616 18604 6656
rect 18644 6616 18652 6656
rect 18692 6616 18775 6656
rect 19027 6616 19036 6656
rect 19076 6616 19316 6656
rect 19411 6616 19420 6656
rect 19460 6616 19756 6656
rect 19796 6616 19805 6656
rect 20371 6616 20380 6656
rect 20420 6616 21600 6656
rect 0 6596 90 6616
rect 18412 6572 18452 6616
rect 4483 6532 4492 6572
rect 4532 6532 18452 6572
rect 19276 6488 19316 6616
rect 21510 6596 21600 6616
rect 19660 6532 20524 6572
rect 20564 6532 20573 6572
rect 19660 6488 19700 6532
rect 2947 6448 2956 6488
rect 2996 6448 3340 6488
rect 3380 6448 3389 6488
rect 4387 6448 4396 6488
rect 4436 6448 4780 6488
rect 4820 6448 4829 6488
rect 5635 6448 5644 6488
rect 5684 6448 9148 6488
rect 9188 6448 9197 6488
rect 9379 6448 9388 6488
rect 9428 6448 11692 6488
rect 11732 6448 11741 6488
rect 12876 6448 12940 6488
rect 12980 6448 13036 6488
rect 13076 6448 13111 6488
rect 13193 6448 13228 6488
rect 13268 6448 13324 6488
rect 13364 6448 13373 6488
rect 14659 6448 14668 6488
rect 14708 6448 14717 6488
rect 14899 6448 14908 6488
rect 14948 6448 18220 6488
rect 18260 6448 18269 6488
rect 18403 6448 18412 6488
rect 18452 6448 18583 6488
rect 18787 6448 18796 6488
rect 18836 6448 18845 6488
rect 19171 6448 19180 6488
rect 19220 6448 19229 6488
rect 19276 6448 19700 6488
rect 19747 6448 19756 6488
rect 19796 6448 19927 6488
rect 20131 6448 20140 6488
rect 20180 6448 20908 6488
rect 20948 6448 20957 6488
rect 14668 6404 14708 6448
rect 18796 6404 18836 6448
rect 1507 6364 1516 6404
rect 1556 6364 14708 6404
rect 14755 6364 14764 6404
rect 14804 6364 18124 6404
rect 18164 6364 18173 6404
rect 18499 6364 18508 6404
rect 18548 6364 18836 6404
rect 0 6320 90 6340
rect 19180 6320 19220 6448
rect 21510 6320 21600 6340
rect 0 6280 1420 6320
rect 1460 6280 1469 6320
rect 3571 6280 3580 6320
rect 3620 6280 10676 6320
rect 10723 6280 10732 6320
rect 10772 6280 13084 6320
rect 13124 6280 13133 6320
rect 15148 6280 19220 6320
rect 20515 6280 20524 6320
rect 20564 6280 21600 6320
rect 0 6260 90 6280
rect 10636 6236 10676 6280
rect 4627 6196 4636 6236
rect 4676 6196 8716 6236
rect 8756 6196 8765 6236
rect 10636 6196 13804 6236
rect 13844 6196 13853 6236
rect 15148 6152 15188 6280
rect 21510 6260 21600 6280
rect 18787 6196 18796 6236
rect 18836 6196 19516 6236
rect 19556 6196 19565 6236
rect 1315 6112 1324 6152
rect 1364 6112 15188 6152
rect 4919 6028 4928 6068
rect 4968 6028 5010 6068
rect 5050 6028 5092 6068
rect 5132 6028 5174 6068
rect 5214 6028 5256 6068
rect 5296 6028 5305 6068
rect 7084 6028 8716 6068
rect 8756 6028 8765 6068
rect 8899 6028 8908 6068
rect 8948 6028 14572 6068
rect 14612 6028 14621 6068
rect 14947 6028 14956 6068
rect 14996 6028 18412 6068
rect 18452 6028 18461 6068
rect 20039 6028 20048 6068
rect 20088 6028 20130 6068
rect 20170 6028 20212 6068
rect 20252 6028 20294 6068
rect 20334 6028 20376 6068
rect 20416 6028 20425 6068
rect 0 5984 90 6004
rect 7084 5984 7124 6028
rect 21510 5984 21600 6004
rect 0 5944 212 5984
rect 2179 5944 2188 5984
rect 2228 5944 7124 5984
rect 7171 5944 7180 5984
rect 7220 5944 18796 5984
rect 18836 5944 18845 5984
rect 19996 5944 21600 5984
rect 0 5924 90 5944
rect 172 5816 212 5944
rect 19996 5900 20036 5944
rect 21510 5924 21600 5944
rect 2860 5860 8620 5900
rect 8660 5860 8669 5900
rect 8803 5860 8812 5900
rect 8852 5860 17356 5900
rect 17396 5860 17405 5900
rect 18691 5860 18700 5900
rect 18740 5860 19132 5900
rect 19172 5860 19181 5900
rect 19987 5860 19996 5900
rect 20036 5860 20045 5900
rect 2860 5816 2900 5860
rect 172 5776 2900 5816
rect 9292 5776 11980 5816
rect 12020 5776 12029 5816
rect 12307 5776 12316 5816
rect 12356 5776 13036 5816
rect 13076 5776 13085 5816
rect 15139 5776 15148 5816
rect 15188 5776 19660 5816
rect 19700 5776 19709 5816
rect 9292 5732 9332 5776
rect 3331 5692 3340 5732
rect 3380 5692 6164 5732
rect 0 5648 90 5668
rect 6124 5648 6164 5692
rect 8524 5692 9332 5732
rect 9379 5692 9388 5732
rect 9428 5692 18836 5732
rect 8524 5648 8564 5692
rect 18796 5648 18836 5692
rect 20140 5692 20620 5732
rect 20660 5692 20669 5732
rect 20140 5648 20180 5692
rect 21510 5648 21600 5668
rect 0 5608 1516 5648
rect 1556 5608 1565 5648
rect 3043 5608 3052 5648
rect 3092 5608 3196 5648
rect 3236 5608 3245 5648
rect 3427 5608 3436 5648
rect 3476 5608 4724 5648
rect 4771 5608 4780 5648
rect 4820 5608 5780 5648
rect 5827 5608 5836 5648
rect 5876 5608 5932 5648
rect 5972 5608 6007 5648
rect 6124 5608 8284 5648
rect 8324 5608 8333 5648
rect 8515 5608 8524 5648
rect 8564 5608 8573 5648
rect 9161 5608 9292 5648
rect 9332 5608 9341 5648
rect 9571 5608 9580 5648
rect 9620 5608 10636 5648
rect 10676 5608 10685 5648
rect 11011 5608 11020 5648
rect 11060 5608 11069 5648
rect 12067 5608 12076 5648
rect 12116 5608 14476 5648
rect 14516 5608 14525 5648
rect 14825 5608 14956 5648
rect 14996 5608 15005 5648
rect 15113 5608 15196 5648
rect 15236 5608 15244 5648
rect 15284 5608 15293 5648
rect 16003 5608 16012 5648
rect 16052 5608 18220 5648
rect 18260 5608 18269 5648
rect 18787 5608 18796 5648
rect 18836 5608 18845 5648
rect 19241 5608 19372 5648
rect 19412 5608 19421 5648
rect 19651 5608 19660 5648
rect 19700 5608 19756 5648
rect 19796 5608 19831 5648
rect 20131 5608 20140 5648
rect 20180 5608 20189 5648
rect 20371 5608 20380 5648
rect 20420 5608 20524 5648
rect 20564 5608 20573 5648
rect 20707 5608 20716 5648
rect 20756 5608 21600 5648
rect 0 5588 90 5608
rect 4684 5564 4724 5608
rect 3427 5524 3436 5564
rect 3476 5524 4540 5564
rect 4580 5524 4589 5564
rect 4684 5524 5644 5564
rect 5684 5524 5693 5564
rect 5740 5480 5780 5608
rect 11020 5564 11060 5608
rect 21510 5588 21600 5608
rect 11020 5524 12556 5564
rect 12596 5524 12605 5564
rect 19027 5524 19036 5564
rect 19076 5524 20812 5564
rect 20852 5524 20861 5564
rect 3235 5440 3244 5480
rect 3284 5440 5596 5480
rect 5636 5440 5645 5480
rect 5740 5440 9196 5480
rect 9236 5440 9245 5480
rect 9523 5440 9532 5480
rect 9572 5440 10732 5480
rect 10772 5440 10781 5480
rect 10867 5440 10876 5480
rect 10916 5440 10925 5480
rect 11251 5440 11260 5480
rect 11300 5440 11309 5480
rect 13987 5440 13996 5480
rect 14036 5440 17980 5480
rect 18020 5440 18029 5480
rect 3580 5356 9292 5396
rect 9332 5356 9341 5396
rect 0 5312 90 5332
rect 3580 5312 3620 5356
rect 0 5272 3620 5312
rect 3679 5272 3688 5312
rect 3728 5272 3770 5312
rect 3810 5272 3852 5312
rect 3892 5272 3934 5312
rect 3974 5272 4016 5312
rect 4056 5272 4065 5312
rect 4195 5272 4204 5312
rect 4244 5272 6604 5312
rect 6644 5272 6653 5312
rect 6883 5272 6892 5312
rect 6932 5272 9772 5312
rect 9812 5272 9821 5312
rect 0 5252 90 5272
rect 10876 5228 10916 5440
rect 11260 5396 11300 5440
rect 11260 5356 15916 5396
rect 15956 5356 15965 5396
rect 16108 5356 20812 5396
rect 20852 5356 20861 5396
rect 14851 5272 14860 5312
rect 14900 5272 16012 5312
rect 16052 5272 16061 5312
rect 16108 5228 16148 5356
rect 21510 5312 21600 5332
rect 18799 5272 18808 5312
rect 18848 5272 18890 5312
rect 18930 5272 18972 5312
rect 19012 5272 19054 5312
rect 19094 5272 19136 5312
rect 19176 5272 19185 5312
rect 19996 5272 21600 5312
rect 547 5188 556 5228
rect 596 5188 9388 5228
rect 9428 5188 9437 5228
rect 10876 5188 16148 5228
rect 19996 5144 20036 5272
rect 21510 5252 21600 5272
rect 172 5104 12980 5144
rect 13027 5104 13036 5144
rect 13076 5104 16108 5144
rect 16148 5104 16157 5144
rect 16243 5104 16252 5144
rect 16292 5104 18508 5144
rect 18548 5104 18557 5144
rect 19987 5104 19996 5144
rect 20036 5104 20045 5144
rect 0 4976 90 4996
rect 172 4976 212 5104
rect 4579 5020 4588 5060
rect 4628 5020 7036 5060
rect 7076 5020 7085 5060
rect 7555 5020 7564 5060
rect 7604 5020 7612 5060
rect 7652 5020 7735 5060
rect 7852 5020 9676 5060
rect 9716 5020 9725 5060
rect 7852 4976 7892 5020
rect 12940 4976 12980 5104
rect 15331 5020 15340 5060
rect 15380 5020 19660 5060
rect 19700 5020 19709 5060
rect 20371 5020 20380 5060
rect 20420 5020 20716 5060
rect 20756 5020 20765 5060
rect 21510 4976 21600 4996
rect 0 4936 212 4976
rect 1027 4936 1036 4976
rect 1076 4936 3724 4976
rect 3764 4936 3773 4976
rect 5155 4936 5164 4976
rect 5204 4936 5836 4976
rect 5876 4936 5885 4976
rect 6595 4936 6604 4976
rect 6644 4936 6652 4976
rect 6692 4936 6775 4976
rect 6883 4936 6892 4976
rect 6932 4936 7063 4976
rect 7267 4936 7276 4976
rect 7316 4936 7660 4976
rect 7700 4936 7709 4976
rect 7843 4936 7852 4976
rect 7892 4936 7901 4976
rect 8035 4936 8044 4976
rect 8084 4936 8092 4976
rect 8132 4936 8215 4976
rect 8323 4936 8332 4976
rect 8372 4936 9484 4976
rect 9524 4936 9533 4976
rect 12940 4936 13804 4976
rect 13844 4936 13853 4976
rect 15881 4936 16012 4976
rect 16052 4936 16061 4976
rect 18691 4936 18700 4976
rect 18740 4936 19036 4976
rect 19076 4936 19085 4976
rect 19267 4936 19276 4976
rect 19316 4936 19325 4976
rect 19625 4936 19756 4976
rect 19796 4936 19805 4976
rect 19852 4936 20140 4976
rect 20180 4936 20189 4976
rect 20515 4936 20524 4976
rect 20564 4936 21600 4976
rect 0 4916 90 4936
rect 19276 4892 19316 4936
rect 2860 4852 19316 4892
rect 0 4640 90 4660
rect 2860 4640 2900 4852
rect 19852 4808 19892 4936
rect 21510 4916 21600 4936
rect 3955 4768 3964 4808
rect 4004 4768 16396 4808
rect 16436 4768 16445 4808
rect 18211 4768 18220 4808
rect 18260 4768 19892 4808
rect 5395 4684 5404 4724
rect 5444 4684 6604 4724
rect 6644 4684 6653 4724
rect 6787 4684 6796 4724
rect 6836 4684 7564 4724
rect 7604 4684 7613 4724
rect 14035 4684 14044 4724
rect 14084 4684 18740 4724
rect 18931 4684 18940 4724
rect 18980 4684 19892 4724
rect 0 4600 2900 4640
rect 0 4580 90 4600
rect 4919 4516 4928 4556
rect 4968 4516 5010 4556
rect 5050 4516 5092 4556
rect 5132 4516 5174 4556
rect 5214 4516 5256 4556
rect 5296 4516 5305 4556
rect 7843 4516 7852 4556
rect 7892 4516 12076 4556
rect 12116 4516 12125 4556
rect 2860 4432 16012 4472
rect 16052 4432 16061 4472
rect 2860 4388 2900 4432
rect 18700 4388 18740 4684
rect 19852 4640 19892 4684
rect 21510 4640 21600 4660
rect 19852 4600 21600 4640
rect 21510 4580 21600 4600
rect 20039 4516 20048 4556
rect 20088 4516 20130 4556
rect 20170 4516 20212 4556
rect 20252 4516 20294 4556
rect 20334 4516 20376 4556
rect 20416 4516 20425 4556
rect 931 4348 940 4388
rect 980 4348 2900 4388
rect 3139 4348 3148 4388
rect 3188 4348 6796 4388
rect 6836 4348 6845 4388
rect 6979 4348 6988 4388
rect 7028 4348 13996 4388
rect 14036 4348 14045 4388
rect 18700 4348 20180 4388
rect 0 4304 90 4324
rect 0 4264 10060 4304
rect 10100 4264 10109 4304
rect 12115 4264 12124 4304
rect 12164 4264 12460 4304
rect 12500 4264 12509 4304
rect 15379 4264 15388 4304
rect 15428 4264 17396 4304
rect 17923 4264 17932 4304
rect 17972 4264 19132 4304
rect 19172 4264 19181 4304
rect 19459 4264 19468 4304
rect 19508 4264 19517 4304
rect 0 4244 90 4264
rect 17356 4220 17396 4264
rect 19468 4220 19508 4264
rect 259 4180 268 4220
rect 308 4180 2900 4220
rect 3427 4180 3436 4220
rect 3476 4180 9580 4220
rect 9620 4180 9629 4220
rect 11884 4180 13420 4220
rect 13460 4180 13469 4220
rect 15331 4180 15340 4220
rect 15380 4180 15628 4220
rect 15668 4180 15677 4220
rect 15811 4180 15820 4220
rect 15860 4180 16780 4220
rect 16820 4180 16829 4220
rect 17356 4180 19508 4220
rect 2860 4052 2900 4180
rect 11884 4136 11924 4180
rect 20140 4136 20180 4348
rect 21510 4304 21600 4324
rect 20371 4264 20380 4304
rect 20420 4264 20524 4304
rect 20564 4264 20573 4304
rect 20707 4264 20716 4304
rect 20756 4264 21600 4304
rect 21510 4244 21600 4264
rect 3523 4096 3532 4136
rect 3572 4096 3868 4136
rect 3908 4096 3917 4136
rect 4099 4096 4108 4136
rect 4148 4096 11692 4136
rect 11732 4096 11741 4136
rect 11875 4096 11884 4136
rect 11924 4096 11933 4136
rect 15017 4096 15148 4136
rect 15188 4096 15197 4136
rect 18665 4096 18796 4136
rect 18836 4096 18845 4136
rect 19337 4096 19372 4136
rect 19412 4096 19468 4136
rect 19508 4096 19517 4136
rect 19564 4096 19603 4136
rect 19643 4096 19652 4136
rect 20131 4096 20140 4136
rect 20180 4096 20189 4136
rect 2860 4012 10060 4052
rect 10100 4012 10109 4052
rect 19027 4012 19036 4052
rect 19076 4012 19180 4052
rect 19220 4012 19229 4052
rect 0 3968 90 3988
rect 0 3928 2900 3968
rect 9187 3928 9196 3968
rect 9236 3928 15244 3968
rect 15284 3928 15293 3968
rect 0 3908 90 3928
rect 2860 3884 2900 3928
rect 19564 3884 19604 4096
rect 21510 3968 21600 3988
rect 19795 3928 19804 3968
rect 19844 3928 19892 3968
rect 20035 3928 20044 3968
rect 20084 3928 21600 3968
rect 2860 3844 19604 3884
rect 172 3760 3436 3800
rect 3476 3760 3485 3800
rect 3679 3760 3688 3800
rect 3728 3760 3770 3800
rect 3810 3760 3852 3800
rect 3892 3760 3934 3800
rect 3974 3760 4016 3800
rect 4056 3760 4065 3800
rect 4972 3760 16972 3800
rect 17012 3760 17021 3800
rect 18799 3760 18808 3800
rect 18848 3760 18890 3800
rect 18930 3760 18972 3800
rect 19012 3760 19054 3800
rect 19094 3760 19136 3800
rect 19176 3760 19185 3800
rect 0 3632 90 3652
rect 172 3632 212 3760
rect 4972 3716 5012 3760
rect 1219 3676 1228 3716
rect 1268 3676 5012 3716
rect 9763 3676 9772 3716
rect 9812 3676 12268 3716
rect 12308 3676 12317 3716
rect 12940 3676 15052 3716
rect 15092 3676 15101 3716
rect 16588 3676 19276 3716
rect 19316 3676 19325 3716
rect 12940 3632 12980 3676
rect 16588 3632 16628 3676
rect 0 3592 212 3632
rect 9065 3592 9148 3632
rect 9188 3592 9196 3632
rect 9236 3592 9245 3632
rect 10963 3592 10972 3632
rect 11012 3592 12980 3632
rect 13603 3592 13612 3632
rect 13652 3592 13660 3632
rect 13700 3592 13783 3632
rect 14035 3592 14044 3632
rect 14084 3592 16628 3632
rect 16819 3592 16828 3632
rect 16868 3592 18316 3632
rect 18356 3592 18365 3632
rect 0 3572 90 3592
rect 1315 3508 1324 3548
rect 1364 3508 14996 3548
rect 15043 3508 15052 3548
rect 15092 3508 17644 3548
rect 17684 3508 17693 3548
rect 14956 3464 14996 3508
rect 19852 3464 19892 3928
rect 21510 3908 21600 3928
rect 21510 3632 21600 3652
rect 20371 3592 20380 3632
rect 20420 3592 20716 3632
rect 20756 3592 20765 3632
rect 21091 3592 21100 3632
rect 21140 3592 21600 3632
rect 21510 3572 21600 3592
rect 1891 3424 1900 3464
rect 1940 3424 1996 3464
rect 2036 3424 2071 3464
rect 6307 3424 6316 3464
rect 6356 3424 6796 3464
rect 6836 3424 6845 3464
rect 8393 3424 8524 3464
rect 8564 3424 8573 3464
rect 8707 3424 8716 3464
rect 8756 3424 8908 3464
rect 8948 3424 8957 3464
rect 9833 3424 9964 3464
rect 10004 3424 10013 3464
rect 10723 3424 10732 3464
rect 10772 3424 10781 3464
rect 10828 3424 12076 3464
rect 12116 3424 12125 3464
rect 12940 3424 13420 3464
rect 13460 3424 13469 3464
rect 13795 3424 13804 3464
rect 13844 3424 13853 3464
rect 14947 3424 14956 3464
rect 14996 3424 15005 3464
rect 16579 3424 16588 3464
rect 16628 3424 16637 3464
rect 16841 3424 16972 3464
rect 17012 3424 17021 3464
rect 19241 3424 19372 3464
rect 19412 3424 19421 3464
rect 19786 3424 19795 3464
rect 19835 3424 19892 3464
rect 19939 3424 19948 3464
rect 19988 3424 20140 3464
rect 20180 3424 20189 3464
rect 10732 3380 10772 3424
rect 10828 3380 10868 3424
rect 12940 3380 12980 3424
rect 9667 3340 9676 3380
rect 9716 3340 10772 3380
rect 10819 3340 10828 3380
rect 10868 3340 10877 3380
rect 11587 3340 11596 3380
rect 11636 3340 12980 3380
rect 13804 3380 13844 3424
rect 16588 3380 16628 3424
rect 13804 3340 16396 3380
rect 16436 3340 16445 3380
rect 16588 3340 18796 3380
rect 18836 3340 18845 3380
rect 19555 3340 19564 3380
rect 19604 3340 20716 3380
rect 20756 3340 20765 3380
rect 0 3296 90 3316
rect 21510 3296 21600 3316
rect 0 3256 748 3296
rect 788 3256 797 3296
rect 2131 3256 2140 3296
rect 2180 3256 2900 3296
rect 8755 3256 8764 3296
rect 8804 3256 18508 3296
rect 18548 3256 18557 3296
rect 19603 3256 19612 3296
rect 19652 3256 21600 3296
rect 0 3236 90 3256
rect 2860 3128 2900 3256
rect 21510 3236 21600 3256
rect 6547 3172 6556 3212
rect 6596 3172 9772 3212
rect 9812 3172 9821 3212
rect 10195 3172 10204 3212
rect 10244 3172 10868 3212
rect 12307 3172 12316 3212
rect 12356 3172 15052 3212
rect 15092 3172 15101 3212
rect 15187 3172 15196 3212
rect 15236 3172 16204 3212
rect 16244 3172 16253 3212
rect 17203 3172 17212 3212
rect 17252 3172 19276 3212
rect 19316 3172 19325 3212
rect 19913 3172 19996 3212
rect 20036 3172 20044 3212
rect 20084 3172 20093 3212
rect 10828 3128 10868 3172
rect 2860 3088 8948 3128
rect 10828 3088 18700 3128
rect 18740 3088 18749 3128
rect 4919 3004 4928 3044
rect 4968 3004 5010 3044
rect 5050 3004 5092 3044
rect 5132 3004 5174 3044
rect 5214 3004 5256 3044
rect 5296 3004 5305 3044
rect 8716 3004 8812 3044
rect 8852 3004 8861 3044
rect 0 2960 90 2980
rect 0 2920 8468 2960
rect 0 2900 90 2920
rect 8428 2876 8468 2920
rect 8716 2876 8756 3004
rect 8908 2960 8948 3088
rect 9091 3004 9100 3044
rect 9140 3004 15340 3044
rect 15380 3004 15389 3044
rect 20039 3004 20048 3044
rect 20088 3004 20130 3044
rect 20170 3004 20212 3044
rect 20252 3004 20294 3044
rect 20334 3004 20376 3044
rect 20416 3004 20425 3044
rect 21510 2960 21600 2980
rect 8908 2920 13364 2960
rect 15043 2920 15052 2960
rect 15092 2920 19468 2960
rect 19508 2920 19517 2960
rect 20140 2920 21600 2960
rect 8428 2836 8756 2876
rect 13324 2876 13364 2920
rect 20140 2876 20180 2920
rect 21510 2900 21600 2920
rect 13324 2836 15820 2876
rect 15860 2836 15869 2876
rect 18835 2836 18844 2876
rect 18884 2836 19892 2876
rect 19987 2836 19996 2876
rect 20036 2836 20180 2876
rect 20371 2836 20380 2876
rect 20420 2836 21100 2876
rect 21140 2836 21149 2876
rect 19852 2792 19892 2836
rect 12940 2752 19412 2792
rect 19852 2752 20620 2792
rect 20660 2752 20669 2792
rect 0 2624 90 2644
rect 0 2584 2132 2624
rect 6595 2584 6604 2624
rect 6644 2584 7756 2624
rect 7796 2584 7805 2624
rect 0 2564 90 2584
rect 2092 2540 2132 2584
rect 12940 2540 12980 2752
rect 16195 2668 16204 2708
rect 16244 2668 18644 2708
rect 18691 2668 18700 2708
rect 18740 2668 18749 2708
rect 18604 2624 18644 2668
rect 18700 2624 18740 2668
rect 19372 2624 19412 2752
rect 21510 2624 21600 2644
rect 17033 2584 17164 2624
rect 17204 2584 17213 2624
rect 18115 2584 18124 2624
rect 18164 2584 18173 2624
rect 18595 2584 18604 2624
rect 18644 2584 18653 2624
rect 18700 2584 18988 2624
rect 19028 2584 19037 2624
rect 19363 2584 19372 2624
rect 19412 2584 19421 2624
rect 19555 2584 19564 2624
rect 19604 2584 19756 2624
rect 19796 2584 19805 2624
rect 20131 2584 20140 2624
rect 20180 2584 20812 2624
rect 20852 2584 20861 2624
rect 20995 2584 21004 2624
rect 21044 2584 21600 2624
rect 18124 2540 18164 2584
rect 21510 2564 21600 2584
rect 2092 2500 12980 2540
rect 15532 2500 18164 2540
rect 19219 2500 19228 2540
rect 19268 2500 20428 2540
rect 20468 2500 20477 2540
rect 6835 2416 6844 2456
rect 6884 2416 12844 2456
rect 12884 2416 12893 2456
rect 15532 2372 15572 2500
rect 17395 2416 17404 2456
rect 17444 2416 17684 2456
rect 18355 2416 18364 2456
rect 18404 2416 18740 2456
rect 19603 2416 19612 2456
rect 19652 2416 19661 2456
rect 3532 2332 15572 2372
rect 0 2288 90 2308
rect 3532 2288 3572 2332
rect 0 2248 3572 2288
rect 3679 2248 3688 2288
rect 3728 2248 3770 2288
rect 3810 2248 3852 2288
rect 3892 2248 3934 2288
rect 3974 2248 4016 2288
rect 4056 2248 4065 2288
rect 0 2228 90 2248
rect 739 2164 748 2204
rect 788 2164 17300 2204
rect 1411 2080 1420 2120
rect 1460 2080 17164 2120
rect 17204 2080 17213 2120
rect 0 1952 90 1972
rect 0 1912 9964 1952
rect 10004 1912 10013 1952
rect 12931 1912 12940 1952
rect 12980 1912 12989 1952
rect 15209 1912 15340 1952
rect 15380 1912 15389 1952
rect 0 1892 90 1912
rect 12940 1784 12980 1912
rect 17260 1868 17300 2164
rect 17644 1952 17684 2416
rect 18700 2120 18740 2416
rect 18799 2248 18808 2288
rect 18848 2248 18890 2288
rect 18930 2248 18972 2288
rect 19012 2248 19054 2288
rect 19094 2248 19136 2288
rect 19176 2248 19185 2288
rect 18700 2080 19508 2120
rect 18547 1996 18556 2036
rect 18596 1996 19372 2036
rect 19412 1996 19421 2036
rect 19468 1952 19508 2080
rect 19612 2036 19652 2416
rect 21510 2288 21600 2308
rect 19996 2248 21600 2288
rect 19996 2120 20036 2248
rect 21510 2228 21600 2248
rect 19987 2080 19996 2120
rect 20036 2080 20045 2120
rect 19612 1996 20180 2036
rect 20371 1996 20380 2036
rect 20420 1996 21004 2036
rect 21044 1996 21053 2036
rect 20140 1952 20180 1996
rect 21510 1952 21600 1972
rect 17644 1912 17932 1952
rect 17972 1912 17981 1952
rect 18307 1912 18316 1952
rect 18356 1912 18365 1952
rect 18499 1912 18508 1952
rect 18548 1912 18988 1952
rect 19028 1912 19037 1952
rect 19241 1912 19276 1952
rect 19316 1912 19372 1952
rect 19412 1912 19421 1952
rect 19468 1912 19756 1952
rect 19796 1912 19805 1952
rect 20131 1912 20140 1952
rect 20180 1912 20189 1952
rect 20419 1912 20428 1952
rect 20468 1912 21600 1952
rect 18316 1868 18356 1912
rect 21510 1892 21600 1912
rect 17260 1828 18356 1868
rect 19084 1828 20524 1868
rect 20564 1828 20573 1868
rect 19084 1784 19124 1828
rect 12940 1744 17356 1784
rect 17396 1744 17405 1784
rect 18163 1744 18172 1784
rect 18212 1744 19124 1784
rect 19219 1744 19228 1784
rect 19268 1744 21004 1784
rect 21044 1744 21053 1784
rect 13171 1660 13180 1700
rect 13220 1660 15476 1700
rect 15571 1660 15580 1700
rect 15620 1660 19468 1700
rect 19508 1660 19517 1700
rect 19603 1660 19612 1700
rect 19652 1660 19661 1700
rect 0 1616 90 1636
rect 0 1576 1228 1616
rect 1268 1576 1277 1616
rect 0 1556 90 1576
rect 15436 1532 15476 1660
rect 19612 1616 19652 1660
rect 21510 1616 21600 1636
rect 19612 1576 21600 1616
rect 21510 1556 21600 1576
rect 4919 1492 4928 1532
rect 4968 1492 5010 1532
rect 5050 1492 5092 1532
rect 5132 1492 5174 1532
rect 5214 1492 5256 1532
rect 5296 1492 5305 1532
rect 15436 1492 19756 1532
rect 19796 1492 19805 1532
rect 20039 1492 20048 1532
rect 20088 1492 20130 1532
rect 20170 1492 20212 1532
rect 20252 1492 20294 1532
rect 20334 1492 20376 1532
rect 20416 1492 20425 1532
rect 0 1280 90 1300
rect 21510 1280 21600 1300
rect 0 1240 1324 1280
rect 1364 1240 1373 1280
rect 20611 1240 20620 1280
rect 20660 1240 21600 1280
rect 0 1220 90 1240
rect 21510 1220 21600 1240
rect 0 944 90 964
rect 21510 944 21600 964
rect 0 904 1420 944
rect 1460 904 1469 944
rect 20515 904 20524 944
rect 20564 904 21600 944
rect 0 884 90 904
rect 21510 884 21600 904
rect 0 608 90 628
rect 21510 608 21600 628
rect 0 568 8524 608
rect 8564 568 8573 608
rect 20995 568 21004 608
rect 21044 568 21600 608
rect 0 548 90 568
rect 21510 548 21600 568
<< via2 >>
rect 364 10984 404 11024
rect 20716 10984 20756 11024
rect 652 10648 692 10688
rect 20524 10648 20564 10688
rect 268 10312 308 10352
rect 2284 10060 2324 10100
rect 9292 10060 9332 10100
rect 18220 10060 18260 10100
rect 18892 10060 18932 10100
rect 19948 10060 19988 10100
rect 2668 9976 2708 10016
rect 3724 9976 3764 10016
rect 6124 9976 6164 10016
rect 16108 9976 16148 10016
rect 9868 9892 9908 9932
rect 15244 9892 15284 9932
rect 17836 9892 17876 9932
rect 19372 9892 19412 9932
rect 3436 9808 3476 9848
rect 2380 9724 2420 9764
rect 2764 9724 2804 9764
rect 3688 9808 3728 9848
rect 3770 9808 3810 9848
rect 3852 9808 3892 9848
rect 3934 9808 3974 9848
rect 4016 9808 4056 9848
rect 2956 9640 2996 9680
rect 3340 9640 3380 9680
rect 4204 9640 4244 9680
rect 2572 9556 2612 9596
rect 3244 9556 3284 9596
rect 3724 9556 3764 9596
rect 4492 9556 4532 9596
rect 15724 9808 15764 9848
rect 16012 9808 16052 9848
rect 18412 9808 18452 9848
rect 18808 9808 18848 9848
rect 18890 9808 18930 9848
rect 18972 9808 19012 9848
rect 19054 9808 19094 9848
rect 19136 9808 19176 9848
rect 10732 9724 10772 9764
rect 12268 9724 12308 9764
rect 15820 9724 15860 9764
rect 5260 9640 5300 9680
rect 5644 9640 5684 9680
rect 6028 9640 6068 9680
rect 6412 9640 6452 9680
rect 6796 9640 6836 9680
rect 7180 9640 7220 9680
rect 7756 9640 7796 9680
rect 8140 9640 8180 9680
rect 7564 9556 7604 9596
rect 7948 9556 7988 9596
rect 16780 9724 16820 9764
rect 17356 9724 17396 9764
rect 18316 9724 18356 9764
rect 8524 9640 8564 9680
rect 8908 9640 8948 9680
rect 9196 9640 9236 9680
rect 15628 9640 15668 9680
rect 11500 9556 11540 9596
rect 1900 9472 1940 9512
rect 3628 9472 3668 9512
rect 4396 9472 4436 9512
rect 5548 9472 5588 9512
rect 6316 9472 6356 9512
rect 6700 9472 6740 9512
rect 7084 9472 7124 9512
rect 7468 9472 7508 9512
rect 11308 9472 11348 9512
rect 76 9304 116 9344
rect 3052 9388 3092 9428
rect 3340 9388 3380 9428
rect 4876 9388 4916 9428
rect 6508 9388 6548 9428
rect 11788 9388 11828 9428
rect 14572 9472 14612 9512
rect 2092 9304 2132 9344
rect 16204 9556 16244 9596
rect 16492 9556 16532 9596
rect 17932 9556 17972 9596
rect 15820 9472 15860 9512
rect 16396 9472 16436 9512
rect 16780 9472 16820 9512
rect 17068 9472 17108 9512
rect 17356 9472 17396 9512
rect 18796 9472 18836 9512
rect 19084 9472 19124 9512
rect 19564 9472 19604 9512
rect 19756 9472 19796 9512
rect 20236 9472 20276 9512
rect 15436 9388 15476 9428
rect 18028 9388 18068 9428
rect 18604 9388 18644 9428
rect 14956 9304 14996 9344
rect 17164 9304 17204 9344
rect 18220 9304 18260 9344
rect 2572 9220 2612 9260
rect 4396 9220 4436 9260
rect 10348 9220 10388 9260
rect 11884 9220 11924 9260
rect 17548 9220 17588 9260
rect 18988 9220 19028 9260
rect 20908 9220 20948 9260
rect 4780 9136 4820 9176
rect 6316 9136 6356 9176
rect 14092 9136 14132 9176
rect 14764 9136 14804 9176
rect 16876 9136 16916 9176
rect 17260 9136 17300 9176
rect 20524 9136 20564 9176
rect 1612 9052 1652 9092
rect 4396 9052 4436 9092
rect 4928 9052 4968 9092
rect 5010 9052 5050 9092
rect 5092 9052 5132 9092
rect 5174 9052 5214 9092
rect 5256 9052 5296 9092
rect 6700 9052 6740 9092
rect 10060 9052 10100 9092
rect 15436 9052 15476 9092
rect 18028 9052 18068 9092
rect 19372 9052 19412 9092
rect 20048 9052 20088 9092
rect 20130 9052 20170 9092
rect 20212 9052 20252 9092
rect 20294 9052 20334 9092
rect 20376 9052 20416 9092
rect 4204 8968 4244 9008
rect 10252 8968 10292 9008
rect 12844 8968 12884 9008
rect 17548 8968 17588 9008
rect 1804 8884 1844 8924
rect 2572 8884 2612 8924
rect 3148 8884 3188 8924
rect 3532 8884 3572 8924
rect 4108 8884 4148 8924
rect 4300 8884 4340 8924
rect 4684 8884 4724 8924
rect 5356 8884 5396 8924
rect 5452 8800 5492 8840
rect 2188 8716 2228 8756
rect 3148 8716 3188 8756
rect 3724 8716 3764 8756
rect 5644 8716 5684 8756
rect 5836 8884 5876 8924
rect 6220 8884 6260 8924
rect 6604 8884 6644 8924
rect 6988 8884 7028 8924
rect 7372 8884 7412 8924
rect 7660 8884 7700 8924
rect 9100 8884 9140 8924
rect 14188 8884 14228 8924
rect 14764 8884 14804 8924
rect 15340 8884 15380 8924
rect 16108 8884 16148 8924
rect 16588 8884 16628 8924
rect 17260 8884 17300 8924
rect 17452 8884 17492 8924
rect 18316 8968 18356 9008
rect 19564 8968 19604 9008
rect 17740 8884 17780 8924
rect 19948 8884 19988 8924
rect 14380 8800 14420 8840
rect 16972 8800 17012 8840
rect 18124 8800 18164 8840
rect 20620 8800 20660 8840
rect 7180 8716 7220 8756
rect 10828 8716 10868 8756
rect 940 8632 980 8672
rect 1612 8632 1652 8672
rect 2284 8632 2324 8672
rect 3436 8632 3476 8672
rect 4300 8632 4340 8672
rect 4588 8632 4628 8672
rect 5356 8632 5396 8672
rect 6124 8632 6164 8672
rect 6988 8632 7028 8672
rect 15436 8716 15476 8756
rect 16588 8716 16628 8756
rect 16876 8716 16916 8756
rect 18412 8716 18452 8756
rect 19852 8716 19892 8756
rect 15628 8632 15668 8672
rect 16204 8632 16244 8672
rect 16492 8632 16532 8672
rect 16972 8632 17012 8672
rect 17548 8632 17588 8672
rect 17932 8632 17972 8672
rect 18316 8632 18356 8672
rect 18892 8632 18932 8672
rect 20524 8632 20564 8672
rect 4204 8548 4244 8588
rect 16684 8548 16724 8588
rect 17260 8548 17300 8588
rect 18028 8548 18068 8588
rect 18412 8548 18452 8588
rect 19180 8548 19220 8588
rect 2284 8464 2324 8504
rect 7660 8464 7700 8504
rect 18220 8464 18260 8504
rect 17068 8380 17108 8420
rect 1132 8296 1172 8336
rect 3688 8296 3728 8336
rect 3770 8296 3810 8336
rect 3852 8296 3892 8336
rect 3934 8296 3974 8336
rect 4016 8296 4056 8336
rect 16300 8296 16340 8336
rect 19564 8380 19604 8420
rect 15532 8212 15572 8252
rect 17836 8212 17876 8252
rect 18808 8296 18848 8336
rect 18890 8296 18930 8336
rect 18972 8296 19012 8336
rect 19054 8296 19094 8336
rect 19136 8296 19176 8336
rect 19372 8296 19412 8336
rect 19468 8212 19508 8252
rect 1996 8128 2036 8168
rect 9868 8128 9908 8168
rect 10252 8128 10292 8168
rect 17164 8128 17204 8168
rect 18508 8128 18548 8168
rect 11212 8044 11252 8084
rect 15628 8044 15668 8084
rect 18700 8044 18740 8084
rect 268 7960 308 8000
rect 2284 7960 2324 8000
rect 11020 7960 11060 8000
rect 16300 7960 16340 8000
rect 16684 7960 16724 8000
rect 17068 7960 17108 8000
rect 18028 7960 18068 8000
rect 19180 7960 19220 8000
rect 19468 7960 19508 8000
rect 19756 7960 19796 8000
rect 18316 7876 18356 7916
rect 20812 7876 20852 7916
rect 7276 7792 7316 7832
rect 17260 7792 17300 7832
rect 17932 7792 17972 7832
rect 18124 7708 18164 7748
rect 21004 7708 21044 7748
rect 1324 7624 1364 7664
rect 4928 7540 4968 7580
rect 5010 7540 5050 7580
rect 5092 7540 5132 7580
rect 5174 7540 5214 7580
rect 5256 7540 5296 7580
rect 19660 7624 19700 7664
rect 20048 7540 20088 7580
rect 20130 7540 20170 7580
rect 20212 7540 20252 7580
rect 20294 7540 20334 7580
rect 20376 7540 20416 7580
rect 15724 7456 15764 7496
rect 20716 7456 20756 7496
rect 7948 7372 7988 7412
rect 11500 7372 11540 7412
rect 14476 7372 14516 7412
rect 18124 7372 18164 7412
rect 19372 7372 19412 7412
rect 556 7288 596 7328
rect 8812 7288 8852 7328
rect 13900 7288 13940 7328
rect 16012 7288 16052 7328
rect 13324 7204 13364 7244
rect 13708 7204 13748 7244
rect 1900 7120 1940 7160
rect 2188 7120 2228 7160
rect 4396 7120 4436 7160
rect 4780 7120 4820 7160
rect 8716 7120 8756 7160
rect 10348 7120 10388 7160
rect 11596 7120 11636 7160
rect 11788 7120 11828 7160
rect 13036 7120 13076 7160
rect 11404 7036 11444 7076
rect 12748 7036 12788 7076
rect 4492 6952 4532 6992
rect 21004 7288 21044 7328
rect 18412 7204 18452 7244
rect 14380 7120 14420 7160
rect 16492 7120 16532 7160
rect 17452 7120 17492 7160
rect 17740 7120 17780 7160
rect 18124 7120 18164 7160
rect 19660 7120 19700 7160
rect 18700 7036 18740 7076
rect 5356 6952 5396 6992
rect 7468 6952 7508 6992
rect 13132 6952 13172 6992
rect 16972 6952 17012 6992
rect 17260 6952 17300 6992
rect 18028 6952 18068 6992
rect 19276 6952 19316 6992
rect 7852 6868 7892 6908
rect 3688 6784 3728 6824
rect 3770 6784 3810 6824
rect 3852 6784 3892 6824
rect 3934 6784 3974 6824
rect 4016 6784 4056 6824
rect 4300 6784 4340 6824
rect 7948 6784 7988 6824
rect 11884 6784 11924 6824
rect 12940 6784 12980 6824
rect 14188 6784 14228 6824
rect 18808 6784 18848 6824
rect 18890 6784 18930 6824
rect 18972 6784 19012 6824
rect 19054 6784 19094 6824
rect 19136 6784 19176 6824
rect 7084 6700 7124 6740
rect 8908 6616 8948 6656
rect 13036 6616 13076 6656
rect 13516 6616 13556 6656
rect 14092 6616 14132 6656
rect 16972 6616 17012 6656
rect 18412 6616 18452 6656
rect 18604 6616 18644 6656
rect 19756 6616 19796 6656
rect 4492 6532 4532 6572
rect 20524 6532 20564 6572
rect 2956 6448 2996 6488
rect 4780 6448 4820 6488
rect 5644 6448 5684 6488
rect 11692 6448 11732 6488
rect 13036 6448 13076 6488
rect 13228 6448 13268 6488
rect 18220 6448 18260 6488
rect 18412 6448 18452 6488
rect 19756 6448 19796 6488
rect 20908 6448 20948 6488
rect 1516 6364 1556 6404
rect 14764 6364 14804 6404
rect 18124 6364 18164 6404
rect 18508 6364 18548 6404
rect 1420 6280 1460 6320
rect 10732 6280 10772 6320
rect 20524 6280 20564 6320
rect 8716 6196 8756 6236
rect 13804 6196 13844 6236
rect 18796 6196 18836 6236
rect 1324 6112 1364 6152
rect 4928 6028 4968 6068
rect 5010 6028 5050 6068
rect 5092 6028 5132 6068
rect 5174 6028 5214 6068
rect 5256 6028 5296 6068
rect 8716 6028 8756 6068
rect 8908 6028 8948 6068
rect 14572 6028 14612 6068
rect 14956 6028 14996 6068
rect 18412 6028 18452 6068
rect 20048 6028 20088 6068
rect 20130 6028 20170 6068
rect 20212 6028 20252 6068
rect 20294 6028 20334 6068
rect 20376 6028 20416 6068
rect 2188 5944 2228 5984
rect 7180 5944 7220 5984
rect 18796 5944 18836 5984
rect 8620 5860 8660 5900
rect 8812 5860 8852 5900
rect 17356 5860 17396 5900
rect 18700 5860 18740 5900
rect 11980 5776 12020 5816
rect 13036 5776 13076 5816
rect 15148 5776 15188 5816
rect 19660 5776 19700 5816
rect 3340 5692 3380 5732
rect 9388 5692 9428 5732
rect 20620 5692 20660 5732
rect 1516 5608 1556 5648
rect 3052 5608 3092 5648
rect 5932 5608 5972 5648
rect 9292 5608 9332 5648
rect 9580 5608 9620 5648
rect 14476 5608 14516 5648
rect 14956 5608 14996 5648
rect 15244 5608 15284 5648
rect 16012 5608 16052 5648
rect 19372 5608 19412 5648
rect 19660 5608 19700 5648
rect 20524 5608 20564 5648
rect 20716 5608 20756 5648
rect 3436 5524 3476 5564
rect 5644 5524 5684 5564
rect 12556 5524 12596 5564
rect 20812 5524 20852 5564
rect 3244 5440 3284 5480
rect 9196 5440 9236 5480
rect 10732 5440 10772 5480
rect 13996 5440 14036 5480
rect 9292 5356 9332 5396
rect 3688 5272 3728 5312
rect 3770 5272 3810 5312
rect 3852 5272 3892 5312
rect 3934 5272 3974 5312
rect 4016 5272 4056 5312
rect 4204 5272 4244 5312
rect 6604 5272 6644 5312
rect 6892 5272 6932 5312
rect 9772 5272 9812 5312
rect 15916 5356 15956 5396
rect 20812 5356 20852 5396
rect 14860 5272 14900 5312
rect 16012 5272 16052 5312
rect 18808 5272 18848 5312
rect 18890 5272 18930 5312
rect 18972 5272 19012 5312
rect 19054 5272 19094 5312
rect 19136 5272 19176 5312
rect 556 5188 596 5228
rect 9388 5188 9428 5228
rect 13036 5104 13076 5144
rect 16108 5104 16148 5144
rect 18508 5104 18548 5144
rect 4588 5020 4628 5060
rect 7564 5020 7604 5060
rect 9676 5020 9716 5060
rect 15340 5020 15380 5060
rect 19660 5020 19700 5060
rect 20716 5020 20756 5060
rect 1036 4936 1076 4976
rect 5836 4936 5876 4976
rect 6604 4936 6644 4976
rect 6892 4936 6932 4976
rect 7660 4936 7700 4976
rect 8044 4936 8084 4976
rect 9484 4936 9524 4976
rect 16012 4936 16052 4976
rect 19756 4936 19796 4976
rect 20524 4936 20564 4976
rect 16396 4768 16436 4808
rect 18220 4768 18260 4808
rect 6604 4684 6644 4724
rect 6796 4684 6836 4724
rect 7564 4684 7604 4724
rect 4928 4516 4968 4556
rect 5010 4516 5050 4556
rect 5092 4516 5132 4556
rect 5174 4516 5214 4556
rect 5256 4516 5296 4556
rect 7852 4516 7892 4556
rect 12076 4516 12116 4556
rect 16012 4432 16052 4472
rect 20048 4516 20088 4556
rect 20130 4516 20170 4556
rect 20212 4516 20252 4556
rect 20294 4516 20334 4556
rect 20376 4516 20416 4556
rect 940 4348 980 4388
rect 3148 4348 3188 4388
rect 6796 4348 6836 4388
rect 6988 4348 7028 4388
rect 13996 4348 14036 4388
rect 10060 4264 10100 4304
rect 12460 4264 12500 4304
rect 17932 4264 17972 4304
rect 19468 4264 19508 4304
rect 268 4180 308 4220
rect 3436 4180 3476 4220
rect 9580 4180 9620 4220
rect 13420 4180 13460 4220
rect 15340 4180 15380 4220
rect 15628 4180 15668 4220
rect 15820 4180 15860 4220
rect 16780 4180 16820 4220
rect 20524 4264 20564 4304
rect 20716 4264 20756 4304
rect 3532 4096 3572 4136
rect 11692 4096 11732 4136
rect 15148 4096 15188 4136
rect 18796 4096 18836 4136
rect 19468 4096 19508 4136
rect 10060 4012 10100 4052
rect 19180 4012 19220 4052
rect 9196 3928 9236 3968
rect 15244 3928 15284 3968
rect 20044 3928 20084 3968
rect 3436 3760 3476 3800
rect 3688 3760 3728 3800
rect 3770 3760 3810 3800
rect 3852 3760 3892 3800
rect 3934 3760 3974 3800
rect 4016 3760 4056 3800
rect 16972 3760 17012 3800
rect 18808 3760 18848 3800
rect 18890 3760 18930 3800
rect 18972 3760 19012 3800
rect 19054 3760 19094 3800
rect 19136 3760 19176 3800
rect 1228 3676 1268 3716
rect 9772 3676 9812 3716
rect 12268 3676 12308 3716
rect 15052 3676 15092 3716
rect 19276 3676 19316 3716
rect 9196 3592 9236 3632
rect 13612 3592 13652 3632
rect 18316 3592 18356 3632
rect 1324 3508 1364 3548
rect 15052 3508 15092 3548
rect 17644 3508 17684 3548
rect 20716 3592 20756 3632
rect 21100 3592 21140 3632
rect 1996 3424 2036 3464
rect 6796 3424 6836 3464
rect 8524 3424 8564 3464
rect 8716 3424 8756 3464
rect 9964 3424 10004 3464
rect 16972 3424 17012 3464
rect 19372 3424 19412 3464
rect 19948 3424 19988 3464
rect 9676 3340 9716 3380
rect 10828 3340 10868 3380
rect 11596 3340 11636 3380
rect 16396 3340 16436 3380
rect 18796 3340 18836 3380
rect 19564 3340 19604 3380
rect 20716 3340 20756 3380
rect 748 3256 788 3296
rect 18508 3256 18548 3296
rect 9772 3172 9812 3212
rect 15052 3172 15092 3212
rect 16204 3172 16244 3212
rect 19276 3172 19316 3212
rect 20044 3172 20084 3212
rect 18700 3088 18740 3128
rect 4928 3004 4968 3044
rect 5010 3004 5050 3044
rect 5092 3004 5132 3044
rect 5174 3004 5214 3044
rect 5256 3004 5296 3044
rect 8812 3004 8852 3044
rect 9100 3004 9140 3044
rect 15340 3004 15380 3044
rect 20048 3004 20088 3044
rect 20130 3004 20170 3044
rect 20212 3004 20252 3044
rect 20294 3004 20334 3044
rect 20376 3004 20416 3044
rect 15052 2920 15092 2960
rect 19468 2920 19508 2960
rect 15820 2836 15860 2876
rect 21100 2836 21140 2876
rect 20620 2752 20660 2792
rect 7756 2584 7796 2624
rect 16204 2668 16244 2708
rect 18700 2668 18740 2708
rect 17164 2584 17204 2624
rect 19564 2584 19604 2624
rect 20812 2584 20852 2624
rect 21004 2584 21044 2624
rect 20428 2500 20468 2540
rect 12844 2416 12884 2456
rect 3688 2248 3728 2288
rect 3770 2248 3810 2288
rect 3852 2248 3892 2288
rect 3934 2248 3974 2288
rect 4016 2248 4056 2288
rect 748 2164 788 2204
rect 1420 2080 1460 2120
rect 17164 2080 17204 2120
rect 9964 1912 10004 1952
rect 15340 1912 15380 1952
rect 18808 2248 18848 2288
rect 18890 2248 18930 2288
rect 18972 2248 19012 2288
rect 19054 2248 19094 2288
rect 19136 2248 19176 2288
rect 19372 1996 19412 2036
rect 21004 1996 21044 2036
rect 18508 1912 18548 1952
rect 19276 1912 19316 1952
rect 20428 1912 20468 1952
rect 20524 1828 20564 1868
rect 17356 1744 17396 1784
rect 21004 1744 21044 1784
rect 19468 1660 19508 1700
rect 1228 1576 1268 1616
rect 4928 1492 4968 1532
rect 5010 1492 5050 1532
rect 5092 1492 5132 1532
rect 5174 1492 5214 1532
rect 5256 1492 5296 1532
rect 19756 1492 19796 1532
rect 20048 1492 20088 1532
rect 20130 1492 20170 1532
rect 20212 1492 20252 1532
rect 20294 1492 20334 1532
rect 20376 1492 20416 1532
rect 1324 1240 1364 1280
rect 20620 1240 20660 1280
rect 1420 904 1460 944
rect 20524 904 20564 944
rect 8524 568 8564 608
rect 21004 568 21044 608
<< metal3 >>
rect 1784 11764 1864 11844
rect 1976 11764 2056 11844
rect 2168 11764 2248 11844
rect 2360 11764 2440 11844
rect 2552 11764 2632 11844
rect 2744 11764 2824 11844
rect 2936 11764 3016 11844
rect 3128 11764 3208 11844
rect 3320 11764 3400 11844
rect 3512 11764 3592 11844
rect 3704 11764 3784 11844
rect 3896 11764 3976 11844
rect 4088 11764 4168 11844
rect 4280 11764 4360 11844
rect 4472 11764 4552 11844
rect 4664 11764 4744 11844
rect 4856 11764 4936 11844
rect 5048 11764 5128 11844
rect 5240 11764 5320 11844
rect 5432 11764 5512 11844
rect 5624 11764 5704 11844
rect 5816 11764 5896 11844
rect 6008 11764 6088 11844
rect 6200 11764 6280 11844
rect 6392 11764 6472 11844
rect 6584 11764 6664 11844
rect 6776 11764 6856 11844
rect 6968 11764 7048 11844
rect 7160 11764 7240 11844
rect 7352 11764 7432 11844
rect 7544 11764 7624 11844
rect 7736 11764 7816 11844
rect 7928 11764 8008 11844
rect 8120 11764 8200 11844
rect 8312 11764 8392 11844
rect 8504 11764 8584 11844
rect 8696 11764 8776 11844
rect 8888 11764 8968 11844
rect 9080 11764 9160 11844
rect 9272 11764 9352 11844
rect 9464 11764 9544 11844
rect 9656 11764 9736 11844
rect 9848 11764 9928 11844
rect 10040 11764 10120 11844
rect 10232 11764 10312 11844
rect 10424 11764 10504 11844
rect 10616 11764 10696 11844
rect 10808 11764 10888 11844
rect 11000 11764 11080 11844
rect 11192 11764 11272 11844
rect 11384 11764 11464 11844
rect 11576 11764 11656 11844
rect 11768 11764 11848 11844
rect 11960 11764 12040 11844
rect 12152 11764 12232 11844
rect 12344 11764 12424 11844
rect 12536 11764 12616 11844
rect 12728 11764 12808 11844
rect 12920 11764 13000 11844
rect 13112 11764 13192 11844
rect 13304 11764 13384 11844
rect 13496 11764 13576 11844
rect 13688 11764 13768 11844
rect 13880 11764 13960 11844
rect 14072 11764 14152 11844
rect 14264 11764 14344 11844
rect 14456 11764 14536 11844
rect 14648 11764 14728 11844
rect 14840 11764 14920 11844
rect 15032 11764 15112 11844
rect 15224 11764 15304 11844
rect 15416 11764 15496 11844
rect 15608 11764 15688 11844
rect 15800 11764 15880 11844
rect 15992 11764 16072 11844
rect 16184 11764 16264 11844
rect 16376 11764 16456 11844
rect 16568 11764 16648 11844
rect 16760 11764 16840 11844
rect 16952 11764 17032 11844
rect 17144 11764 17224 11844
rect 17336 11764 17416 11844
rect 17528 11764 17608 11844
rect 17720 11764 17800 11844
rect 17912 11764 17992 11844
rect 18104 11764 18184 11844
rect 18296 11764 18376 11844
rect 18488 11764 18568 11844
rect 18680 11764 18760 11844
rect 18872 11764 18952 11844
rect 19064 11764 19144 11844
rect 19256 11764 19336 11844
rect 19448 11764 19528 11844
rect 364 11024 404 11033
rect 268 10352 308 10361
rect 76 9344 116 9353
rect 76 9209 116 9304
rect 268 8840 308 10312
rect 364 9512 404 10984
rect 364 9463 404 9472
rect 652 10688 692 10697
rect 268 8791 308 8800
rect 652 8672 692 10648
rect 1612 9092 1652 9101
rect 652 8623 692 8632
rect 940 8672 980 8681
rect 268 8000 308 8009
rect 268 4220 308 7960
rect 556 7328 596 7337
rect 556 5228 596 7288
rect 556 5179 596 5188
rect 940 4388 980 8632
rect 1612 8672 1652 9052
rect 1804 8924 1844 11764
rect 1804 8875 1844 8884
rect 1900 9512 1940 9521
rect 1612 8623 1652 8632
rect 1132 8336 1172 8345
rect 1132 5732 1172 8296
rect 1324 7664 1364 7673
rect 1324 6152 1364 7624
rect 1900 7160 1940 9472
rect 1996 8168 2036 11764
rect 2092 9344 2132 9353
rect 2092 9209 2132 9304
rect 2188 8756 2228 11764
rect 2188 8707 2228 8716
rect 2284 10100 2324 10109
rect 2284 8672 2324 10060
rect 2380 9764 2420 11764
rect 2380 9715 2420 9724
rect 2572 9596 2612 11764
rect 2572 9547 2612 9556
rect 2668 10016 2708 10025
rect 2572 9260 2612 9269
rect 2572 8924 2612 9220
rect 2572 8875 2612 8884
rect 2668 8924 2708 9976
rect 2764 9764 2804 11764
rect 2764 9715 2804 9724
rect 2956 9680 2996 11764
rect 2956 9631 2996 9640
rect 2668 8875 2708 8884
rect 3052 9428 3092 9437
rect 2284 8623 2324 8632
rect 1996 8119 2036 8128
rect 2284 8504 2324 8513
rect 2284 8000 2324 8464
rect 2284 7951 2324 7960
rect 1900 7111 1940 7120
rect 2188 7160 2228 7169
rect 1516 6404 1556 6413
rect 1420 6320 1460 6329
rect 1420 6185 1460 6280
rect 1324 6103 1364 6112
rect 1132 5683 1172 5692
rect 1516 5648 1556 6364
rect 2188 5984 2228 7120
rect 2188 5935 2228 5944
rect 2956 6488 2996 6497
rect 1516 5599 1556 5608
rect 940 4339 980 4348
rect 1036 4976 1076 4985
rect 268 4171 308 4180
rect 748 3296 788 3305
rect 748 2204 788 3256
rect 748 2155 788 2164
rect 1036 80 1076 4936
rect 1228 3716 1268 3725
rect 1228 1616 1268 3676
rect 1228 1567 1268 1576
rect 1324 3548 1364 3557
rect 1324 1280 1364 3508
rect 1996 3464 2036 3473
rect 1324 1231 1364 1240
rect 1420 2120 1460 2129
rect 1420 944 1460 2080
rect 1420 895 1460 904
rect 1996 80 2036 3424
rect 2956 80 2996 6448
rect 3052 5648 3092 9388
rect 3148 8924 3188 11764
rect 3340 9680 3380 11764
rect 3340 9631 3380 9640
rect 3436 9848 3476 9857
rect 3148 8875 3188 8884
rect 3244 9596 3284 9605
rect 3052 5599 3092 5608
rect 3148 8756 3188 8765
rect 3148 4388 3188 8716
rect 3244 5480 3284 9556
rect 3340 9428 3380 9437
rect 3340 5732 3380 9388
rect 3436 9428 3476 9808
rect 3436 9379 3476 9388
rect 3532 8924 3572 11764
rect 3724 10016 3764 11764
rect 3916 10184 3956 11764
rect 4108 10268 4148 11764
rect 4108 10228 4244 10268
rect 3916 10144 4148 10184
rect 3724 9967 3764 9976
rect 3688 9848 4056 9857
rect 3728 9808 3770 9848
rect 3810 9808 3852 9848
rect 3892 9808 3934 9848
rect 3974 9808 4016 9848
rect 3688 9799 4056 9808
rect 3724 9596 3764 9605
rect 3532 8875 3572 8884
rect 3628 9512 3668 9521
rect 3340 5683 3380 5692
rect 3436 8672 3476 8681
rect 3436 5564 3476 8632
rect 3628 8504 3668 9472
rect 3724 8756 3764 9556
rect 4108 8924 4148 10144
rect 4204 9680 4244 10228
rect 4204 9631 4244 9640
rect 4108 8875 4148 8884
rect 4204 9008 4244 9017
rect 3724 8707 3764 8716
rect 4204 8756 4244 8968
rect 4300 8924 4340 11764
rect 4492 9596 4532 11764
rect 4492 9547 4532 9556
rect 4396 9512 4436 9521
rect 4396 9260 4436 9472
rect 4396 9211 4436 9220
rect 4300 8875 4340 8884
rect 4396 9092 4436 9101
rect 4204 8707 4244 8716
rect 4300 8672 4340 8681
rect 3436 5515 3476 5524
rect 3532 8464 3668 8504
rect 4204 8588 4244 8597
rect 3244 5431 3284 5440
rect 3148 4339 3188 4348
rect 3436 4220 3476 4229
rect 3436 3800 3476 4180
rect 3532 4136 3572 8464
rect 3688 8336 4056 8345
rect 3728 8296 3770 8336
rect 3810 8296 3852 8336
rect 3892 8296 3934 8336
rect 3974 8296 4016 8336
rect 3688 8287 4056 8296
rect 3688 6824 4056 6833
rect 3728 6784 3770 6824
rect 3810 6784 3852 6824
rect 3892 6784 3934 6824
rect 3974 6784 4016 6824
rect 3688 6775 4056 6784
rect 3688 5312 4056 5321
rect 3728 5272 3770 5312
rect 3810 5272 3852 5312
rect 3892 5272 3934 5312
rect 3974 5272 4016 5312
rect 3688 5263 4056 5272
rect 4204 5312 4244 8548
rect 4300 6992 4340 8632
rect 4396 7160 4436 9052
rect 4684 8924 4724 11764
rect 4876 9428 4916 11764
rect 4876 9379 4916 9388
rect 5068 9260 5108 11764
rect 5260 9680 5300 11764
rect 5260 9631 5300 9640
rect 5068 9220 5396 9260
rect 4684 8875 4724 8884
rect 4780 9176 4820 9185
rect 4396 7111 4436 7120
rect 4588 8672 4628 8681
rect 4300 6943 4340 6952
rect 4492 6992 4532 7001
rect 4204 5263 4244 5272
rect 4300 6824 4340 6833
rect 3532 4087 3572 4096
rect 3436 3751 3476 3760
rect 3688 3800 4056 3809
rect 3728 3760 3770 3800
rect 3810 3760 3852 3800
rect 3892 3760 3934 3800
rect 3974 3760 4016 3800
rect 3688 3751 4056 3760
rect 3688 2288 4056 2297
rect 3728 2248 3770 2288
rect 3810 2248 3852 2288
rect 3892 2248 3934 2288
rect 3974 2248 4016 2288
rect 3688 2239 4056 2248
rect 3916 148 4148 188
rect 3916 80 3956 148
rect 1016 0 1096 80
rect 1976 0 2056 80
rect 2936 0 3016 80
rect 3896 0 3976 80
rect 4108 60 4148 148
rect 4300 60 4340 6784
rect 4492 6572 4532 6952
rect 4492 6523 4532 6532
rect 4588 5060 4628 8632
rect 4780 7160 4820 9136
rect 4928 9092 5296 9101
rect 4968 9052 5010 9092
rect 5050 9052 5092 9092
rect 5132 9052 5174 9092
rect 5214 9052 5256 9092
rect 4928 9043 5296 9052
rect 5356 8924 5396 9220
rect 5356 8875 5396 8884
rect 5452 8840 5492 11764
rect 5644 9680 5684 11764
rect 5644 9631 5684 9640
rect 5452 8791 5492 8800
rect 5548 9512 5588 9521
rect 5356 8672 5396 8681
rect 4928 7580 5296 7589
rect 4968 7540 5010 7580
rect 5050 7540 5092 7580
rect 5132 7540 5174 7580
rect 5214 7540 5256 7580
rect 4928 7531 5296 7540
rect 4780 7111 4820 7120
rect 5356 6992 5396 8632
rect 5356 6943 5396 6952
rect 5548 6908 5588 9472
rect 5836 8924 5876 11764
rect 5836 8875 5876 8884
rect 5932 10016 5972 10025
rect 5548 6859 5588 6868
rect 5644 8756 5684 8765
rect 4588 5011 4628 5020
rect 4780 6488 4820 6497
rect 4780 944 4820 6448
rect 5644 6488 5684 8716
rect 5644 6439 5684 6448
rect 4928 6068 5296 6077
rect 4968 6028 5010 6068
rect 5050 6028 5092 6068
rect 5132 6028 5174 6068
rect 5214 6028 5256 6068
rect 4928 6019 5296 6028
rect 5932 5648 5972 9976
rect 6028 9680 6068 11764
rect 6028 9631 6068 9640
rect 6124 10016 6164 10025
rect 6124 8672 6164 9976
rect 6220 8924 6260 11764
rect 6412 9680 6452 11764
rect 6412 9631 6452 9640
rect 6316 9512 6356 9521
rect 6316 9176 6356 9472
rect 6508 9428 6548 9437
rect 6508 9344 6548 9388
rect 6508 9293 6548 9304
rect 6316 9127 6356 9136
rect 6220 8875 6260 8884
rect 6604 8924 6644 11764
rect 6796 9680 6836 11764
rect 6796 9631 6836 9640
rect 6700 9512 6740 9521
rect 6700 9092 6740 9472
rect 6700 9043 6740 9052
rect 6604 8875 6644 8884
rect 6988 8924 7028 11764
rect 7180 9680 7220 11764
rect 7180 9631 7220 9640
rect 6988 8875 7028 8884
rect 7084 9512 7124 9521
rect 6124 8623 6164 8632
rect 6988 8672 7028 8681
rect 5932 5599 5972 5608
rect 5644 5564 5684 5573
rect 5644 5429 5684 5524
rect 6604 5312 6644 5321
rect 5836 4976 5876 4985
rect 4928 4556 5296 4565
rect 4968 4516 5010 4556
rect 5050 4516 5092 4556
rect 5132 4516 5174 4556
rect 5214 4516 5256 4556
rect 4928 4507 5296 4516
rect 4928 3044 5296 3053
rect 4968 3004 5010 3044
rect 5050 3004 5092 3044
rect 5132 3004 5174 3044
rect 5214 3004 5256 3044
rect 4928 2995 5296 3004
rect 4928 1532 5296 1541
rect 4968 1492 5010 1532
rect 5050 1492 5092 1532
rect 5132 1492 5174 1532
rect 5214 1492 5256 1532
rect 4928 1483 5296 1492
rect 4780 904 4916 944
rect 4876 80 4916 904
rect 5836 80 5876 4936
rect 6604 4976 6644 5272
rect 6604 4927 6644 4936
rect 6892 5312 6932 5321
rect 6892 4976 6932 5272
rect 6892 4927 6932 4936
rect 6604 4724 6644 4733
rect 6604 4640 6644 4684
rect 6604 4589 6644 4600
rect 6796 4724 6836 4733
rect 6796 4388 6836 4684
rect 6796 4339 6836 4348
rect 6988 4388 7028 8632
rect 7084 6740 7124 9472
rect 7276 9344 7316 9353
rect 7084 6691 7124 6700
rect 7180 8756 7220 8765
rect 7180 5984 7220 8716
rect 7276 7832 7316 9304
rect 7372 8924 7412 11764
rect 7564 9596 7604 11764
rect 7756 9680 7796 11764
rect 7756 9631 7796 9640
rect 7564 9547 7604 9556
rect 7948 9596 7988 11764
rect 8140 9680 8180 11764
rect 8140 9631 8180 9640
rect 8332 9680 8372 11764
rect 8332 9631 8372 9640
rect 8524 9680 8564 11764
rect 8524 9631 8564 9640
rect 7948 9547 7988 9556
rect 7372 8875 7412 8884
rect 7468 9512 7508 9521
rect 7276 7783 7316 7792
rect 7468 6992 7508 9472
rect 8620 9512 8660 9521
rect 7660 8924 7700 8933
rect 7660 8504 7700 8884
rect 7660 8455 7700 8464
rect 7468 6943 7508 6952
rect 7948 7412 7988 7421
rect 7852 6908 7892 6917
rect 7852 6773 7892 6868
rect 7948 6824 7988 7372
rect 7948 6775 7988 6784
rect 8044 6992 8084 7001
rect 7180 5935 7220 5944
rect 7564 5060 7604 5069
rect 7564 4724 7604 5020
rect 7564 4675 7604 4684
rect 7660 4976 7700 4985
rect 7660 4556 7700 4936
rect 8044 4976 8084 6952
rect 8620 5900 8660 9472
rect 8716 7160 8756 11764
rect 8908 9848 8948 11764
rect 8812 9808 8948 9848
rect 8812 7328 8852 9808
rect 8908 9680 8948 9689
rect 8908 9545 8948 9640
rect 9100 8924 9140 11764
rect 9292 10100 9332 11764
rect 9292 10051 9332 10060
rect 9196 9680 9236 9689
rect 9196 9512 9236 9640
rect 9196 9463 9236 9472
rect 9100 8875 9140 8884
rect 8812 7279 8852 7288
rect 8716 7111 8756 7120
rect 8908 6656 8948 6665
rect 8716 6236 8756 6245
rect 8756 6196 8852 6236
rect 8716 6187 8756 6196
rect 8716 6068 8756 6077
rect 8716 5933 8756 6028
rect 8620 5851 8660 5860
rect 8812 5900 8852 6196
rect 8908 6068 8948 6616
rect 8908 6019 8948 6028
rect 8812 5851 8852 5860
rect 9388 5732 9428 5741
rect 9292 5648 9332 5657
rect 9196 5480 9236 5489
rect 9196 5345 9236 5440
rect 9292 5396 9332 5608
rect 9292 5347 9332 5356
rect 9388 5228 9428 5692
rect 9388 5179 9428 5188
rect 8044 4927 8084 4936
rect 9484 4976 9524 11764
rect 9484 4927 9524 4936
rect 9580 5648 9620 5657
rect 7852 4556 7892 4565
rect 7660 4516 7852 4556
rect 7852 4507 7892 4516
rect 6988 4339 7028 4348
rect 9580 4220 9620 5608
rect 9676 5060 9716 11764
rect 9868 10100 9908 11764
rect 9772 10060 9908 10100
rect 9772 5312 9812 10060
rect 10060 10016 10100 11764
rect 10060 9967 10100 9976
rect 9868 9932 9908 9941
rect 9868 8168 9908 9892
rect 10252 9176 10292 11764
rect 10156 9136 10292 9176
rect 10348 9260 10388 9269
rect 10060 9092 10100 9101
rect 10060 8957 10100 9052
rect 9868 8119 9908 8128
rect 10156 5480 10196 9136
rect 10252 9008 10292 9017
rect 10252 8168 10292 8968
rect 10252 8119 10292 8128
rect 10348 7160 10388 9220
rect 10348 7111 10388 7120
rect 10444 5564 10484 11764
rect 10636 6068 10676 11764
rect 10732 9764 10772 9773
rect 10732 6320 10772 9724
rect 10828 8756 10868 11764
rect 10828 8707 10868 8716
rect 11020 8000 11060 11764
rect 11212 8084 11252 11764
rect 11212 8035 11252 8044
rect 11308 9512 11348 9521
rect 11020 7951 11060 7960
rect 11308 7160 11348 9472
rect 11308 7111 11348 7120
rect 11404 7076 11444 11764
rect 11500 9596 11540 9605
rect 11500 7412 11540 9556
rect 11500 7363 11540 7372
rect 11596 7160 11636 11764
rect 11788 9596 11828 11764
rect 11596 7111 11636 7120
rect 11692 9556 11828 9596
rect 11404 7027 11444 7036
rect 11692 6488 11732 9556
rect 11788 9428 11828 9437
rect 11788 7160 11828 9388
rect 11788 7111 11828 7120
rect 11884 9260 11924 9269
rect 11884 6824 11924 9220
rect 11884 6775 11924 6784
rect 11692 6439 11732 6448
rect 10732 6271 10772 6280
rect 10636 6019 10676 6028
rect 11980 5816 12020 11764
rect 12172 8420 12212 11764
rect 11980 5767 12020 5776
rect 12076 8380 12212 8420
rect 12268 9764 12308 9773
rect 10444 5515 10484 5524
rect 10156 5431 10196 5440
rect 10732 5480 10772 5489
rect 10732 5345 10772 5440
rect 9772 5263 9812 5272
rect 9676 5011 9716 5020
rect 12076 4556 12116 8380
rect 12076 4507 12116 4516
rect 9580 4171 9620 4180
rect 10060 4304 10100 4313
rect 10060 4169 10100 4264
rect 11692 4136 11732 4145
rect 10060 4052 10100 4061
rect 9196 3968 9236 3977
rect 9196 3632 9236 3928
rect 10060 3917 10100 4012
rect 11692 4001 11732 4096
rect 9196 3583 9236 3592
rect 9772 3716 9812 3725
rect 6796 3464 6836 3473
rect 6796 80 6836 3424
rect 8524 3464 8564 3473
rect 7756 2624 7796 2633
rect 7756 80 7796 2584
rect 8524 608 8564 3424
rect 8524 559 8564 568
rect 8716 3464 8756 3473
rect 8716 80 8756 3424
rect 9676 3380 9716 3389
rect 8812 3044 8852 3053
rect 9100 3044 9140 3053
rect 8852 3004 9100 3044
rect 8812 2995 8852 3004
rect 9100 2995 9140 3004
rect 9676 80 9716 3340
rect 9772 3212 9812 3676
rect 12268 3716 12308 9724
rect 12364 4136 12404 11764
rect 12460 8504 12500 8513
rect 12460 4304 12500 8464
rect 12556 6824 12596 11764
rect 12748 7076 12788 11764
rect 12940 11444 12980 11764
rect 12940 11395 12980 11404
rect 12748 7027 12788 7036
rect 12844 9008 12884 9017
rect 12844 6908 12884 8968
rect 13036 7160 13076 7169
rect 13036 7025 13076 7120
rect 13132 6992 13172 11764
rect 13132 6943 13172 6952
rect 13228 11444 13268 11453
rect 12556 6775 12596 6784
rect 12748 6868 12884 6908
rect 12460 4255 12500 4264
rect 12556 5564 12596 5573
rect 12364 4087 12404 4096
rect 12268 3667 12308 3676
rect 9772 3163 9812 3172
rect 9964 3464 10004 3473
rect 9964 1952 10004 3424
rect 9964 1903 10004 1912
rect 10828 3380 10868 3389
rect 10828 188 10868 3340
rect 10636 148 10868 188
rect 11596 3380 11636 3389
rect 10636 80 10676 148
rect 11596 80 11636 3340
rect 12556 80 12596 5524
rect 12748 2900 12788 6868
rect 12940 6824 12980 6833
rect 12940 6689 12980 6784
rect 13036 6656 13076 6665
rect 13036 6488 13076 6616
rect 13036 6439 13076 6448
rect 13228 6488 13268 11404
rect 13324 7244 13364 11764
rect 13324 7195 13364 7204
rect 13516 6656 13556 11764
rect 13516 6607 13556 6616
rect 13612 8588 13652 8597
rect 13228 6439 13268 6448
rect 13036 5816 13076 5825
rect 13036 5144 13076 5776
rect 13036 5095 13076 5104
rect 13420 4220 13460 4229
rect 13460 4180 13556 4220
rect 13420 4171 13460 4180
rect 12748 2860 12884 2900
rect 12844 2456 12884 2860
rect 12844 2407 12884 2416
rect 13516 80 13556 4180
rect 13612 3632 13652 8548
rect 13708 7244 13748 11764
rect 13708 7195 13748 7204
rect 13804 9512 13844 9521
rect 13804 6236 13844 9472
rect 13900 7328 13940 11764
rect 14092 10100 14132 11764
rect 13900 7279 13940 7288
rect 13996 10060 14132 10100
rect 13996 7160 14036 10060
rect 14284 9512 14324 11764
rect 14284 9472 14420 9512
rect 13996 7111 14036 7120
rect 14092 9176 14132 9185
rect 14092 6656 14132 9136
rect 14380 9008 14420 9472
rect 14476 9176 14516 11764
rect 14476 9127 14516 9136
rect 14572 9512 14612 9521
rect 14380 8968 14516 9008
rect 14188 8924 14228 8933
rect 14188 6824 14228 8884
rect 14380 8840 14420 8849
rect 14380 7160 14420 8800
rect 14476 7412 14516 8968
rect 14476 7363 14516 7372
rect 14380 7111 14420 7120
rect 14188 6775 14228 6784
rect 14092 6607 14132 6616
rect 13804 6187 13844 6196
rect 14572 6068 14612 9472
rect 14668 6404 14708 11764
rect 14860 10100 14900 11764
rect 15052 10436 15092 11764
rect 15052 10396 15188 10436
rect 14860 10060 15092 10100
rect 14956 9344 14996 9353
rect 14764 9176 14804 9185
rect 14764 8924 14804 9136
rect 14764 8875 14804 8884
rect 14860 9176 14900 9185
rect 14764 6404 14804 6413
rect 14668 6364 14764 6404
rect 14764 6355 14804 6364
rect 14572 6019 14612 6028
rect 14476 5648 14516 5657
rect 13996 5480 14036 5489
rect 13996 4388 14036 5440
rect 13996 4339 14036 4348
rect 13612 3583 13652 3592
rect 14476 80 14516 5608
rect 14860 5312 14900 9136
rect 14956 6068 14996 9304
rect 15052 6488 15092 10060
rect 15052 6439 15092 6448
rect 14956 6019 14996 6028
rect 15148 5816 15188 10396
rect 15244 9932 15284 11764
rect 15436 9932 15476 11764
rect 15436 9892 15572 9932
rect 15244 9883 15284 9892
rect 15436 9428 15476 9437
rect 15436 9092 15476 9388
rect 15436 9043 15476 9052
rect 15340 8924 15380 8933
rect 15148 5767 15188 5776
rect 15244 5816 15284 5825
rect 14860 5263 14900 5272
rect 14956 5648 14996 5657
rect 14956 2372 14996 5608
rect 15244 5648 15284 5776
rect 15244 5599 15284 5608
rect 15340 5060 15380 8884
rect 15340 5011 15380 5020
rect 15436 8756 15476 8765
rect 15340 4220 15380 4229
rect 15148 4136 15188 4145
rect 15148 4052 15188 4096
rect 15148 4001 15188 4012
rect 15244 3968 15284 3977
rect 15340 3968 15380 4180
rect 15284 3928 15380 3968
rect 15244 3919 15284 3928
rect 15052 3716 15092 3725
rect 15052 3548 15092 3676
rect 15052 3499 15092 3508
rect 15052 3212 15092 3221
rect 15052 2960 15092 3172
rect 15052 2911 15092 2920
rect 15340 3044 15380 3053
rect 14956 2323 14996 2332
rect 15340 1952 15380 3004
rect 15340 1903 15380 1912
rect 15436 80 15476 8716
rect 15532 8252 15572 9892
rect 15628 9680 15668 11764
rect 15628 9631 15668 9640
rect 15724 9848 15764 9857
rect 15532 8203 15572 8212
rect 15628 8672 15668 8681
rect 15628 8084 15668 8632
rect 15628 8035 15668 8044
rect 15724 7496 15764 9808
rect 15820 9764 15860 11764
rect 16012 9848 16052 11764
rect 16012 9799 16052 9808
rect 16108 10016 16148 10025
rect 15820 9715 15860 9724
rect 15820 9512 15860 9521
rect 15820 9428 15860 9472
rect 15820 9377 15860 9388
rect 15916 9344 15956 9353
rect 15724 7447 15764 7456
rect 15820 9260 15860 9269
rect 15820 7076 15860 9220
rect 15628 7036 15860 7076
rect 15628 4220 15668 7036
rect 15916 5396 15956 9304
rect 16012 9092 16052 9101
rect 16012 7328 16052 9052
rect 16108 8924 16148 9976
rect 16204 9596 16244 11764
rect 16396 10520 16436 11764
rect 16396 10480 16532 10520
rect 16204 9547 16244 9556
rect 16492 9596 16532 10480
rect 16492 9547 16532 9556
rect 16396 9512 16436 9521
rect 16108 8875 16148 8884
rect 16300 9428 16340 9437
rect 16204 8756 16244 8767
rect 16204 8672 16244 8716
rect 16204 8623 16244 8632
rect 16300 8504 16340 9388
rect 16012 7279 16052 7288
rect 16108 8464 16340 8504
rect 15916 5347 15956 5356
rect 16012 5648 16052 5657
rect 16012 5312 16052 5608
rect 16012 5263 16052 5272
rect 16108 5144 16148 8464
rect 16300 8336 16340 8345
rect 16300 8000 16340 8296
rect 16300 7951 16340 7960
rect 16108 5095 16148 5104
rect 16012 4976 16052 4985
rect 16012 4472 16052 4936
rect 16396 4808 16436 9472
rect 16492 8924 16532 8933
rect 16492 8672 16532 8884
rect 16588 8924 16628 11764
rect 16780 9764 16820 11764
rect 16780 9715 16820 9724
rect 16588 8875 16628 8884
rect 16780 9512 16820 9521
rect 16492 8623 16532 8632
rect 16588 8756 16628 8765
rect 16588 8621 16628 8716
rect 16684 8588 16724 8597
rect 16684 8000 16724 8548
rect 16684 7951 16724 7960
rect 16492 7160 16532 7169
rect 16492 7025 16532 7120
rect 16396 4759 16436 4768
rect 16012 4423 16052 4432
rect 15628 4171 15668 4180
rect 15820 4220 15860 4229
rect 15820 2876 15860 4180
rect 16780 4220 16820 9472
rect 16876 9176 16916 9185
rect 16876 9041 16916 9136
rect 16972 8840 17012 11764
rect 17068 9512 17108 9521
rect 17068 9377 17108 9472
rect 17164 9344 17204 11764
rect 17356 9764 17396 11764
rect 17356 9715 17396 9724
rect 17164 9295 17204 9304
rect 17356 9512 17396 9521
rect 17260 9176 17300 9185
rect 17260 8924 17300 9136
rect 17260 8875 17300 8884
rect 16972 8791 17012 8800
rect 16876 8756 16916 8765
rect 16876 8621 16916 8716
rect 16972 8672 17012 8681
rect 16972 7160 17012 8632
rect 17260 8588 17300 8597
rect 17068 8420 17108 8429
rect 17068 8000 17108 8380
rect 17164 8168 17204 8177
rect 17260 8168 17300 8548
rect 17204 8128 17300 8168
rect 17164 8119 17204 8128
rect 17068 7951 17108 7960
rect 16876 7120 17012 7160
rect 17260 7832 17300 7841
rect 16876 4640 16916 7120
rect 16972 6992 17012 7001
rect 16972 6656 17012 6952
rect 17260 6992 17300 7792
rect 17260 6943 17300 6952
rect 16972 6607 17012 6616
rect 17356 5900 17396 9472
rect 17548 9260 17588 11764
rect 17548 9211 17588 9220
rect 17644 9512 17684 9521
rect 17548 9008 17588 9017
rect 17452 8924 17492 8933
rect 17452 7160 17492 8884
rect 17548 8672 17588 8968
rect 17548 8623 17588 8632
rect 17452 7111 17492 7120
rect 17356 5851 17396 5860
rect 16876 4591 16916 4600
rect 16780 4171 16820 4180
rect 16972 3800 17012 3809
rect 16972 3464 17012 3760
rect 17644 3548 17684 9472
rect 17740 8924 17780 11764
rect 17740 8875 17780 8884
rect 17836 9932 17876 9941
rect 17836 8420 17876 9892
rect 17932 9596 17972 11764
rect 17932 9547 17972 9556
rect 18028 9428 18068 9437
rect 18028 9260 18068 9388
rect 18028 9211 18068 9220
rect 18028 9092 18068 9101
rect 17932 8840 17972 8849
rect 17932 8672 17972 8800
rect 17932 8623 17972 8632
rect 18028 8588 18068 9052
rect 18124 8840 18164 11764
rect 18220 10100 18260 10109
rect 18220 9596 18260 10060
rect 18316 9764 18356 11764
rect 18316 9715 18356 9724
rect 18412 9848 18452 9857
rect 18220 9556 18356 9596
rect 18124 8791 18164 8800
rect 18220 9344 18260 9353
rect 18028 8539 18068 8548
rect 18220 8504 18260 9304
rect 18316 9008 18356 9556
rect 18316 8959 18356 8968
rect 18412 8756 18452 9808
rect 18412 8707 18452 8716
rect 18316 8672 18356 8681
rect 18316 8537 18356 8632
rect 18412 8588 18452 8597
rect 18220 8455 18260 8464
rect 18412 8453 18452 8548
rect 17740 8380 17876 8420
rect 17740 7160 17780 8380
rect 17836 8252 17876 8261
rect 17836 8000 17876 8212
rect 18508 8168 18548 11764
rect 18508 8119 18548 8128
rect 18604 9428 18644 9437
rect 18028 8000 18068 8009
rect 17836 7960 18028 8000
rect 18028 7951 18068 7960
rect 18316 7916 18356 7925
rect 17740 7111 17780 7120
rect 17932 7832 17972 7841
rect 17932 4304 17972 7792
rect 18124 7748 18164 7757
rect 18124 7412 18164 7708
rect 18124 7363 18164 7372
rect 18124 7160 18164 7169
rect 18028 6992 18068 7001
rect 18028 5816 18068 6952
rect 18124 6404 18164 7120
rect 18124 6355 18164 6364
rect 18220 6488 18260 6497
rect 18028 5767 18068 5776
rect 18220 4808 18260 6448
rect 18220 4759 18260 4768
rect 17932 4255 17972 4264
rect 18316 3632 18356 7876
rect 18412 7244 18452 7253
rect 18412 6656 18452 7204
rect 18412 6607 18452 6616
rect 18604 6656 18644 9388
rect 18700 8084 18740 11764
rect 18892 10100 18932 11764
rect 18892 10051 18932 10060
rect 19084 10016 19124 11764
rect 19276 10100 19316 11764
rect 19468 10184 19508 11764
rect 20716 11024 20756 11033
rect 20524 10688 20564 10697
rect 19468 10144 19700 10184
rect 19276 10060 19508 10100
rect 19084 9976 19316 10016
rect 18808 9848 19176 9857
rect 18848 9808 18890 9848
rect 18930 9808 18972 9848
rect 19012 9808 19054 9848
rect 19094 9808 19136 9848
rect 18808 9799 19176 9808
rect 18796 9512 18836 9521
rect 18796 9377 18836 9472
rect 19084 9512 19124 9521
rect 18988 9260 19028 9271
rect 18988 9176 19028 9220
rect 18988 9127 19028 9136
rect 18892 8672 18932 8681
rect 18892 8504 18932 8632
rect 18892 8455 18932 8464
rect 19084 8504 19124 9472
rect 19180 8672 19220 8683
rect 19180 8588 19220 8632
rect 19180 8539 19220 8548
rect 19084 8455 19124 8464
rect 18808 8336 19176 8345
rect 18848 8296 18890 8336
rect 18930 8296 18972 8336
rect 19012 8296 19054 8336
rect 19094 8296 19136 8336
rect 18808 8287 19176 8296
rect 18700 8035 18740 8044
rect 19180 8000 19220 8009
rect 18604 6607 18644 6616
rect 18700 7076 18740 7085
rect 18412 6488 18452 6497
rect 18412 6068 18452 6448
rect 18412 6019 18452 6028
rect 18508 6404 18548 6413
rect 18508 5144 18548 6364
rect 18700 5900 18740 7036
rect 19180 6992 19220 7960
rect 19180 6943 19220 6952
rect 19276 6992 19316 9976
rect 19372 9932 19412 9941
rect 19372 9092 19412 9892
rect 19372 9043 19412 9052
rect 19372 8336 19412 8345
rect 19372 7412 19412 8296
rect 19468 8252 19508 10060
rect 19564 9512 19604 9521
rect 19564 9344 19604 9472
rect 19564 9295 19604 9304
rect 19564 9008 19604 9017
rect 19564 8420 19604 8968
rect 19564 8371 19604 8380
rect 19468 8203 19508 8212
rect 19372 7363 19412 7372
rect 19468 8000 19508 8009
rect 19276 6943 19316 6952
rect 18808 6824 19176 6833
rect 18848 6784 18890 6824
rect 18930 6784 18972 6824
rect 19012 6784 19054 6824
rect 19094 6784 19136 6824
rect 18808 6775 19176 6784
rect 19276 6824 19316 6833
rect 18796 6236 18836 6245
rect 18796 5984 18836 6196
rect 18796 5935 18836 5944
rect 18700 5851 18740 5860
rect 18808 5312 19176 5321
rect 18848 5272 18890 5312
rect 18930 5272 18972 5312
rect 19012 5272 19054 5312
rect 19094 5272 19136 5312
rect 18808 5263 19176 5272
rect 18508 5095 18548 5104
rect 18796 4304 18836 4313
rect 18796 4136 18836 4264
rect 18796 4087 18836 4096
rect 19180 4052 19220 4147
rect 19180 4003 19220 4012
rect 18808 3800 19176 3809
rect 18848 3760 18890 3800
rect 18930 3760 18972 3800
rect 19012 3760 19054 3800
rect 19094 3760 19136 3800
rect 18808 3751 19176 3760
rect 19276 3716 19316 6784
rect 19372 5648 19412 5657
rect 19372 5513 19412 5608
rect 19276 3667 19316 3676
rect 19372 5396 19412 5405
rect 19372 3632 19412 5356
rect 19468 4304 19508 7960
rect 19660 7664 19700 10144
rect 19948 10100 19988 10109
rect 19756 9512 19796 9521
rect 19756 9428 19796 9472
rect 19756 9377 19796 9388
rect 19948 8924 19988 10060
rect 20236 9596 20276 9607
rect 20236 9512 20276 9556
rect 20236 9463 20276 9472
rect 20524 9176 20564 10648
rect 20524 9127 20564 9136
rect 20048 9092 20416 9101
rect 20088 9052 20130 9092
rect 20170 9052 20212 9092
rect 20252 9052 20294 9092
rect 20334 9052 20376 9092
rect 20048 9043 20416 9052
rect 19948 8875 19988 8884
rect 20620 8840 20660 8849
rect 19852 8756 19892 8765
rect 19660 7615 19700 7624
rect 19756 8000 19796 8009
rect 19660 7160 19700 7169
rect 19660 5816 19700 7120
rect 19756 6656 19796 7960
rect 19756 6607 19796 6616
rect 19756 6488 19796 6497
rect 19756 6353 19796 6448
rect 19660 5767 19700 5776
rect 19660 5648 19700 5657
rect 19660 5060 19700 5608
rect 19660 5011 19700 5020
rect 19756 5480 19796 5489
rect 19756 4976 19796 5440
rect 19756 4927 19796 4936
rect 19468 4255 19508 4264
rect 19468 4136 19508 4145
rect 19468 3716 19508 4096
rect 19468 3676 19604 3716
rect 19372 3592 19508 3632
rect 18316 3583 18356 3592
rect 17644 3499 17684 3508
rect 16972 3415 17012 3424
rect 19372 3464 19412 3473
rect 16396 3380 16436 3389
rect 15820 2827 15860 2836
rect 16204 3212 16244 3221
rect 16204 2708 16244 3172
rect 16204 2659 16244 2668
rect 16396 80 16436 3340
rect 18796 3380 18836 3389
rect 18508 3296 18548 3305
rect 17164 2624 17204 2633
rect 17164 2120 17204 2584
rect 17164 2071 17204 2080
rect 18316 2372 18356 2381
rect 17356 1784 17396 1793
rect 17356 80 17396 1744
rect 18316 80 18356 2332
rect 18508 1952 18548 3256
rect 18700 3128 18740 3137
rect 18700 2708 18740 3088
rect 18700 2659 18740 2668
rect 18796 2456 18836 3340
rect 18508 1903 18548 1912
rect 18700 2416 18836 2456
rect 19276 3212 19316 3221
rect 18700 104 18740 2416
rect 18808 2288 19176 2297
rect 18848 2248 18890 2288
rect 18930 2248 18972 2288
rect 19012 2248 19054 2288
rect 19094 2248 19136 2288
rect 18808 2239 19176 2248
rect 19276 1952 19316 3172
rect 19372 2036 19412 3424
rect 19468 2960 19508 3592
rect 19564 3380 19604 3676
rect 19564 3331 19604 3340
rect 19468 2911 19508 2920
rect 19852 2900 19892 8716
rect 20524 8672 20564 8681
rect 20048 7580 20416 7589
rect 20088 7540 20130 7580
rect 20170 7540 20212 7580
rect 20252 7540 20294 7580
rect 20334 7540 20376 7580
rect 20048 7531 20416 7540
rect 20524 6572 20564 8632
rect 20524 6523 20564 6532
rect 20524 6320 20564 6329
rect 20048 6068 20416 6077
rect 20088 6028 20130 6068
rect 20170 6028 20212 6068
rect 20252 6028 20294 6068
rect 20334 6028 20376 6068
rect 20048 6019 20416 6028
rect 20524 5648 20564 6280
rect 20620 5732 20660 8800
rect 20716 7496 20756 10984
rect 20908 9260 20948 9269
rect 20716 7447 20756 7456
rect 20812 7916 20852 7925
rect 20620 5683 20660 5692
rect 20524 5599 20564 5608
rect 20716 5648 20756 5657
rect 20716 5060 20756 5608
rect 20812 5564 20852 7876
rect 20908 6488 20948 9220
rect 21004 7748 21044 7757
rect 21004 7328 21044 7708
rect 21004 7279 21044 7288
rect 20908 6439 20948 6448
rect 20812 5515 20852 5524
rect 20716 5011 20756 5020
rect 20812 5396 20852 5405
rect 20524 4976 20564 4985
rect 20048 4556 20416 4565
rect 20088 4516 20130 4556
rect 20170 4516 20212 4556
rect 20252 4516 20294 4556
rect 20334 4516 20376 4556
rect 20048 4507 20416 4516
rect 20524 4304 20564 4936
rect 20524 4255 20564 4264
rect 20716 4304 20756 4313
rect 19948 4052 19988 4061
rect 19948 3464 19988 4012
rect 19948 3415 19988 3424
rect 20044 3968 20084 3977
rect 20044 3212 20084 3928
rect 20716 3632 20756 4264
rect 20716 3583 20756 3592
rect 20044 3163 20084 3172
rect 20716 3380 20756 3389
rect 20048 3044 20416 3053
rect 20088 3004 20130 3044
rect 20170 3004 20212 3044
rect 20252 3004 20294 3044
rect 20334 3004 20376 3044
rect 20048 2995 20416 3004
rect 19756 2860 19892 2900
rect 19372 1987 19412 1996
rect 19564 2624 19604 2633
rect 19276 1903 19316 1912
rect 19468 1700 19508 1709
rect 19564 1700 19604 2584
rect 19508 1660 19604 1700
rect 19468 1651 19508 1660
rect 19756 1532 19796 2860
rect 20620 2792 20660 2801
rect 20428 2540 20468 2549
rect 20428 1952 20468 2500
rect 20428 1903 20468 1912
rect 20524 1868 20564 1877
rect 19756 1483 19796 1492
rect 20048 1532 20416 1541
rect 20088 1492 20130 1532
rect 20170 1492 20212 1532
rect 20252 1492 20294 1532
rect 20334 1492 20376 1532
rect 20048 1483 20416 1492
rect 20524 944 20564 1828
rect 20620 1280 20660 2752
rect 20620 1231 20660 1240
rect 20524 895 20564 904
rect 20236 148 20468 188
rect 4108 20 4340 60
rect 4856 0 4936 80
rect 5816 0 5896 80
rect 6776 0 6856 80
rect 7736 0 7816 80
rect 8696 0 8776 80
rect 9656 0 9736 80
rect 10616 0 10696 80
rect 11576 0 11656 80
rect 12536 0 12616 80
rect 13496 0 13576 80
rect 14456 0 14536 80
rect 15416 0 15496 80
rect 16376 0 16456 80
rect 17336 0 17416 80
rect 18296 0 18376 80
rect 19276 104 19316 113
rect 18700 55 18740 64
rect 19256 64 19276 80
rect 20236 80 20276 148
rect 19316 64 19336 80
rect 19256 0 19336 64
rect 20216 0 20296 80
rect 20428 60 20468 148
rect 20716 60 20756 3340
rect 20812 2624 20852 5356
rect 21100 3632 21140 3641
rect 21100 2876 21140 3592
rect 21100 2827 21140 2836
rect 20812 2575 20852 2584
rect 21004 2624 21044 2633
rect 21004 2036 21044 2584
rect 21004 1987 21044 1996
rect 21004 1784 21044 1793
rect 21004 608 21044 1744
rect 21004 559 21044 568
rect 20428 20 20756 60
<< via3 >>
rect 76 9304 116 9344
rect 364 9472 404 9512
rect 268 8800 308 8840
rect 652 8632 692 8672
rect 2092 9304 2132 9344
rect 2668 8884 2708 8924
rect 1420 6280 1460 6320
rect 1132 5692 1172 5732
rect 3436 9388 3476 9428
rect 3688 9808 3728 9848
rect 3770 9808 3810 9848
rect 3852 9808 3892 9848
rect 3934 9808 3974 9848
rect 4016 9808 4056 9848
rect 4204 8716 4244 8756
rect 3688 8296 3728 8336
rect 3770 8296 3810 8336
rect 3852 8296 3892 8336
rect 3934 8296 3974 8336
rect 4016 8296 4056 8336
rect 3688 6784 3728 6824
rect 3770 6784 3810 6824
rect 3852 6784 3892 6824
rect 3934 6784 3974 6824
rect 4016 6784 4056 6824
rect 3688 5272 3728 5312
rect 3770 5272 3810 5312
rect 3852 5272 3892 5312
rect 3934 5272 3974 5312
rect 4016 5272 4056 5312
rect 4300 6952 4340 6992
rect 3688 3760 3728 3800
rect 3770 3760 3810 3800
rect 3852 3760 3892 3800
rect 3934 3760 3974 3800
rect 4016 3760 4056 3800
rect 3688 2248 3728 2288
rect 3770 2248 3810 2288
rect 3852 2248 3892 2288
rect 3934 2248 3974 2288
rect 4016 2248 4056 2288
rect 4928 9052 4968 9092
rect 5010 9052 5050 9092
rect 5092 9052 5132 9092
rect 5174 9052 5214 9092
rect 5256 9052 5296 9092
rect 4928 7540 4968 7580
rect 5010 7540 5050 7580
rect 5092 7540 5132 7580
rect 5174 7540 5214 7580
rect 5256 7540 5296 7580
rect 5932 9976 5972 10016
rect 5548 6868 5588 6908
rect 4928 6028 4968 6068
rect 5010 6028 5050 6068
rect 5092 6028 5132 6068
rect 5174 6028 5214 6068
rect 5256 6028 5296 6068
rect 6508 9304 6548 9344
rect 5644 5524 5684 5564
rect 4928 4516 4968 4556
rect 5010 4516 5050 4556
rect 5092 4516 5132 4556
rect 5174 4516 5214 4556
rect 5256 4516 5296 4556
rect 4928 3004 4968 3044
rect 5010 3004 5050 3044
rect 5092 3004 5132 3044
rect 5174 3004 5214 3044
rect 5256 3004 5296 3044
rect 4928 1492 4968 1532
rect 5010 1492 5050 1532
rect 5092 1492 5132 1532
rect 5174 1492 5214 1532
rect 5256 1492 5296 1532
rect 6604 4600 6644 4640
rect 7276 9304 7316 9344
rect 8332 9640 8372 9680
rect 8620 9472 8660 9512
rect 7852 6868 7892 6908
rect 8044 6952 8084 6992
rect 8908 9640 8948 9680
rect 9196 9472 9236 9512
rect 8716 6028 8756 6068
rect 9196 5440 9236 5480
rect 10060 9976 10100 10016
rect 10060 9052 10100 9092
rect 11308 7120 11348 7160
rect 10636 6028 10676 6068
rect 10444 5524 10484 5564
rect 10156 5440 10196 5480
rect 10732 5440 10772 5480
rect 10060 4264 10100 4304
rect 11692 4096 11732 4136
rect 10060 4012 10100 4052
rect 12460 8464 12500 8504
rect 12940 11404 12980 11444
rect 13036 7120 13076 7160
rect 13228 11404 13268 11444
rect 12556 6784 12596 6824
rect 12364 4096 12404 4136
rect 12940 6784 12980 6824
rect 13612 8548 13652 8588
rect 13804 9472 13844 9512
rect 13996 7120 14036 7160
rect 14476 9136 14516 9176
rect 14860 9136 14900 9176
rect 15052 6448 15092 6488
rect 15244 5776 15284 5816
rect 15148 4012 15188 4052
rect 14956 2332 14996 2372
rect 15820 9388 15860 9428
rect 15916 9304 15956 9344
rect 15820 9220 15860 9260
rect 16012 9052 16052 9092
rect 16300 9388 16340 9428
rect 16204 8716 16244 8756
rect 16492 8884 16532 8924
rect 16588 8716 16628 8756
rect 16492 7120 16532 7160
rect 16876 9136 16916 9176
rect 17068 9472 17108 9512
rect 16876 8716 16916 8756
rect 17644 9472 17684 9512
rect 16876 4600 16916 4640
rect 18028 9220 18068 9260
rect 17932 8800 17972 8840
rect 18316 8632 18356 8672
rect 18412 8548 18452 8588
rect 18028 5776 18068 5816
rect 18808 9808 18848 9848
rect 18890 9808 18930 9848
rect 18972 9808 19012 9848
rect 19054 9808 19094 9848
rect 19136 9808 19176 9848
rect 18796 9472 18836 9512
rect 18988 9136 19028 9176
rect 18892 8464 18932 8504
rect 19180 8632 19220 8672
rect 19084 8464 19124 8504
rect 18808 8296 18848 8336
rect 18890 8296 18930 8336
rect 18972 8296 19012 8336
rect 19054 8296 19094 8336
rect 19136 8296 19176 8336
rect 19180 6952 19220 6992
rect 19564 9304 19604 9344
rect 18808 6784 18848 6824
rect 18890 6784 18930 6824
rect 18972 6784 19012 6824
rect 19054 6784 19094 6824
rect 19136 6784 19176 6824
rect 19276 6784 19316 6824
rect 18808 5272 18848 5312
rect 18890 5272 18930 5312
rect 18972 5272 19012 5312
rect 19054 5272 19094 5312
rect 19136 5272 19176 5312
rect 18796 4264 18836 4304
rect 19180 4012 19220 4052
rect 18808 3760 18848 3800
rect 18890 3760 18930 3800
rect 18972 3760 19012 3800
rect 19054 3760 19094 3800
rect 19136 3760 19176 3800
rect 19372 5608 19412 5648
rect 19372 5356 19412 5396
rect 19756 9388 19796 9428
rect 20236 9556 20276 9596
rect 20048 9052 20088 9092
rect 20130 9052 20170 9092
rect 20212 9052 20252 9092
rect 20294 9052 20334 9092
rect 20376 9052 20416 9092
rect 19756 6448 19796 6488
rect 19756 5440 19796 5480
rect 18316 2332 18356 2372
rect 18808 2248 18848 2288
rect 18890 2248 18930 2288
rect 18972 2248 19012 2288
rect 19054 2248 19094 2288
rect 19136 2248 19176 2288
rect 20048 7540 20088 7580
rect 20130 7540 20170 7580
rect 20212 7540 20252 7580
rect 20294 7540 20334 7580
rect 20376 7540 20416 7580
rect 20048 6028 20088 6068
rect 20130 6028 20170 6068
rect 20212 6028 20252 6068
rect 20294 6028 20334 6068
rect 20376 6028 20416 6068
rect 20048 4516 20088 4556
rect 20130 4516 20170 4556
rect 20212 4516 20252 4556
rect 20294 4516 20334 4556
rect 20376 4516 20416 4556
rect 19948 4012 19988 4052
rect 20048 3004 20088 3044
rect 20130 3004 20170 3044
rect 20212 3004 20252 3044
rect 20294 3004 20334 3044
rect 20376 3004 20416 3044
rect 20048 1492 20088 1532
rect 20130 1492 20170 1532
rect 20212 1492 20252 1532
rect 20294 1492 20334 1532
rect 20376 1492 20416 1532
rect 18700 64 18740 104
rect 19276 64 19316 104
<< metal4 >>
rect 12931 11404 12940 11444
rect 12980 11404 13228 11444
rect 13268 11404 13277 11444
rect 5923 9976 5932 10016
rect 5972 9976 10060 10016
rect 10100 9976 10109 10016
rect 3679 9808 3688 9848
rect 3728 9808 3770 9848
rect 3810 9808 3852 9848
rect 3892 9808 3934 9848
rect 3974 9808 4016 9848
rect 4056 9808 4065 9848
rect 18799 9808 18808 9848
rect 18848 9808 18890 9848
rect 18930 9808 18972 9848
rect 19012 9808 19054 9848
rect 19094 9808 19136 9848
rect 19176 9808 19185 9848
rect 8323 9640 8332 9680
rect 8372 9640 8908 9680
rect 8948 9640 8957 9680
rect 2860 9556 20236 9596
rect 20276 9556 20285 9596
rect 2860 9512 2900 9556
rect 355 9472 364 9512
rect 404 9472 2900 9512
rect 8611 9472 8620 9512
rect 8660 9472 9196 9512
rect 9236 9472 9245 9512
rect 13795 9472 13804 9512
rect 13844 9472 17068 9512
rect 17108 9472 17117 9512
rect 17635 9472 17644 9512
rect 17684 9472 18796 9512
rect 18836 9472 18845 9512
rect 3427 9388 3436 9428
rect 3476 9388 15820 9428
rect 15860 9388 15869 9428
rect 16291 9388 16300 9428
rect 16340 9388 19756 9428
rect 19796 9388 19805 9428
rect 67 9304 76 9344
rect 116 9304 2092 9344
rect 2132 9304 2141 9344
rect 6499 9304 6508 9344
rect 6548 9304 7276 9344
rect 7316 9304 7325 9344
rect 15907 9304 15916 9344
rect 15956 9304 19564 9344
rect 19604 9304 19613 9344
rect 15811 9220 15820 9260
rect 15860 9220 18028 9260
rect 18068 9220 18077 9260
rect 14467 9136 14476 9176
rect 14516 9136 14860 9176
rect 14900 9136 14909 9176
rect 16867 9136 16876 9176
rect 16916 9136 18988 9176
rect 19028 9136 19037 9176
rect 4919 9052 4928 9092
rect 4968 9052 5010 9092
rect 5050 9052 5092 9092
rect 5132 9052 5174 9092
rect 5214 9052 5256 9092
rect 5296 9052 5305 9092
rect 10051 9052 10060 9092
rect 10100 9052 16012 9092
rect 16052 9052 16061 9092
rect 20039 9052 20048 9092
rect 20088 9052 20130 9092
rect 20170 9052 20212 9092
rect 20252 9052 20294 9092
rect 20334 9052 20376 9092
rect 20416 9052 20425 9092
rect 2659 8884 2668 8924
rect 2708 8884 16492 8924
rect 16532 8884 16541 8924
rect 259 8800 268 8840
rect 308 8800 17932 8840
rect 17972 8800 17981 8840
rect 4195 8716 4204 8756
rect 4244 8716 16204 8756
rect 16244 8716 16253 8756
rect 16579 8716 16588 8756
rect 16628 8716 16876 8756
rect 16916 8716 16925 8756
rect 643 8632 652 8672
rect 692 8632 18316 8672
rect 18356 8632 18365 8672
rect 19171 8632 19180 8672
rect 19220 8632 19276 8672
rect 19316 8632 19325 8672
rect 13603 8548 13612 8588
rect 13652 8548 18412 8588
rect 18452 8548 18461 8588
rect 12451 8464 12460 8504
rect 12500 8464 18892 8504
rect 18932 8464 18941 8504
rect 19075 8464 19084 8504
rect 19124 8464 19372 8504
rect 19412 8464 19421 8504
rect 3679 8296 3688 8336
rect 3728 8296 3770 8336
rect 3810 8296 3852 8336
rect 3892 8296 3934 8336
rect 3974 8296 4016 8336
rect 4056 8296 4065 8336
rect 18799 8296 18808 8336
rect 18848 8296 18890 8336
rect 18930 8296 18972 8336
rect 19012 8296 19054 8336
rect 19094 8296 19136 8336
rect 19176 8296 19185 8336
rect 4919 7540 4928 7580
rect 4968 7540 5010 7580
rect 5050 7540 5092 7580
rect 5132 7540 5174 7580
rect 5214 7540 5256 7580
rect 5296 7540 5305 7580
rect 20039 7540 20048 7580
rect 20088 7540 20130 7580
rect 20170 7540 20212 7580
rect 20252 7540 20294 7580
rect 20334 7540 20376 7580
rect 20416 7540 20425 7580
rect 11299 7120 11308 7160
rect 11348 7120 13036 7160
rect 13076 7120 13085 7160
rect 13987 7120 13996 7160
rect 14036 7120 16492 7160
rect 16532 7120 16541 7160
rect 4291 6952 4300 6992
rect 4340 6952 8044 6992
rect 8084 6952 8093 6992
rect 19171 6952 19180 6992
rect 19220 6952 19229 6992
rect 19180 6908 19220 6952
rect 5539 6868 5548 6908
rect 5588 6868 7852 6908
rect 7892 6868 7901 6908
rect 19180 6868 19316 6908
rect 19276 6824 19316 6868
rect 3679 6784 3688 6824
rect 3728 6784 3770 6824
rect 3810 6784 3852 6824
rect 3892 6784 3934 6824
rect 3974 6784 4016 6824
rect 4056 6784 4065 6824
rect 12547 6784 12556 6824
rect 12596 6784 12940 6824
rect 12980 6784 12989 6824
rect 18799 6784 18808 6824
rect 18848 6784 18890 6824
rect 18930 6784 18972 6824
rect 19012 6784 19054 6824
rect 19094 6784 19136 6824
rect 19176 6784 19185 6824
rect 19267 6784 19276 6824
rect 19316 6784 19325 6824
rect 15043 6448 15052 6488
rect 15092 6448 19756 6488
rect 19796 6448 19805 6488
rect 1411 6280 1420 6320
rect 1460 6280 19276 6320
rect 19316 6280 19325 6320
rect 4919 6028 4928 6068
rect 4968 6028 5010 6068
rect 5050 6028 5092 6068
rect 5132 6028 5174 6068
rect 5214 6028 5256 6068
rect 5296 6028 5305 6068
rect 8707 6028 8716 6068
rect 8756 6028 10636 6068
rect 10676 6028 10685 6068
rect 20039 6028 20048 6068
rect 20088 6028 20130 6068
rect 20170 6028 20212 6068
rect 20252 6028 20294 6068
rect 20334 6028 20376 6068
rect 20416 6028 20425 6068
rect 15235 5776 15244 5816
rect 15284 5776 18028 5816
rect 18068 5776 18077 5816
rect 1123 5692 1132 5732
rect 1172 5692 2900 5732
rect 2860 5648 2900 5692
rect 2860 5608 19372 5648
rect 19412 5608 19421 5648
rect 5635 5524 5644 5564
rect 5684 5524 10444 5564
rect 10484 5524 10493 5564
rect 9187 5440 9196 5480
rect 9236 5440 10156 5480
rect 10196 5440 10205 5480
rect 10723 5440 10732 5480
rect 10772 5440 19756 5480
rect 19796 5440 19805 5480
rect 19277 5356 19372 5396
rect 19412 5356 19421 5396
rect 3679 5272 3688 5312
rect 3728 5272 3770 5312
rect 3810 5272 3852 5312
rect 3892 5272 3934 5312
rect 3974 5272 4016 5312
rect 4056 5272 4065 5312
rect 18799 5272 18808 5312
rect 18848 5272 18890 5312
rect 18930 5272 18972 5312
rect 19012 5272 19054 5312
rect 19094 5272 19136 5312
rect 19176 5272 19185 5312
rect 6595 4600 6604 4640
rect 6644 4600 16876 4640
rect 16916 4600 16925 4640
rect 4919 4516 4928 4556
rect 4968 4516 5010 4556
rect 5050 4516 5092 4556
rect 5132 4516 5174 4556
rect 5214 4516 5256 4556
rect 5296 4516 5305 4556
rect 20039 4516 20048 4556
rect 20088 4516 20130 4556
rect 20170 4516 20212 4556
rect 20252 4516 20294 4556
rect 20334 4516 20376 4556
rect 20416 4516 20425 4556
rect 10051 4264 10060 4304
rect 10100 4264 18796 4304
rect 18836 4264 18845 4304
rect 11683 4096 11692 4136
rect 11732 4096 12364 4136
rect 12404 4096 12413 4136
rect 10051 4012 10060 4052
rect 10100 4012 15148 4052
rect 15188 4012 15197 4052
rect 19171 4012 19180 4052
rect 19220 4012 19948 4052
rect 19988 4012 19997 4052
rect 3679 3760 3688 3800
rect 3728 3760 3770 3800
rect 3810 3760 3852 3800
rect 3892 3760 3934 3800
rect 3974 3760 4016 3800
rect 4056 3760 4065 3800
rect 18799 3760 18808 3800
rect 18848 3760 18890 3800
rect 18930 3760 18972 3800
rect 19012 3760 19054 3800
rect 19094 3760 19136 3800
rect 19176 3760 19185 3800
rect 4919 3004 4928 3044
rect 4968 3004 5010 3044
rect 5050 3004 5092 3044
rect 5132 3004 5174 3044
rect 5214 3004 5256 3044
rect 5296 3004 5305 3044
rect 20039 3004 20048 3044
rect 20088 3004 20130 3044
rect 20170 3004 20212 3044
rect 20252 3004 20294 3044
rect 20334 3004 20376 3044
rect 20416 3004 20425 3044
rect 14947 2332 14956 2372
rect 14996 2332 18316 2372
rect 18356 2332 18365 2372
rect 3679 2248 3688 2288
rect 3728 2248 3770 2288
rect 3810 2248 3852 2288
rect 3892 2248 3934 2288
rect 3974 2248 4016 2288
rect 4056 2248 4065 2288
rect 18799 2248 18808 2288
rect 18848 2248 18890 2288
rect 18930 2248 18972 2288
rect 19012 2248 19054 2288
rect 19094 2248 19136 2288
rect 19176 2248 19185 2288
rect 4919 1492 4928 1532
rect 4968 1492 5010 1532
rect 5050 1492 5092 1532
rect 5132 1492 5174 1532
rect 5214 1492 5256 1532
rect 5296 1492 5305 1532
rect 20039 1492 20048 1532
rect 20088 1492 20130 1532
rect 20170 1492 20212 1532
rect 20252 1492 20294 1532
rect 20334 1492 20376 1532
rect 20416 1492 20425 1532
rect 18691 64 18700 104
rect 18740 64 19276 104
rect 19316 64 19325 104
<< via4 >>
rect 3688 9808 3728 9848
rect 3770 9808 3810 9848
rect 3852 9808 3892 9848
rect 3934 9808 3974 9848
rect 4016 9808 4056 9848
rect 18808 9808 18848 9848
rect 18890 9808 18930 9848
rect 18972 9808 19012 9848
rect 19054 9808 19094 9848
rect 19136 9808 19176 9848
rect 4928 9052 4968 9092
rect 5010 9052 5050 9092
rect 5092 9052 5132 9092
rect 5174 9052 5214 9092
rect 5256 9052 5296 9092
rect 20048 9052 20088 9092
rect 20130 9052 20170 9092
rect 20212 9052 20252 9092
rect 20294 9052 20334 9092
rect 20376 9052 20416 9092
rect 19276 8632 19316 8672
rect 19372 8464 19412 8504
rect 3688 8296 3728 8336
rect 3770 8296 3810 8336
rect 3852 8296 3892 8336
rect 3934 8296 3974 8336
rect 4016 8296 4056 8336
rect 18808 8296 18848 8336
rect 18890 8296 18930 8336
rect 18972 8296 19012 8336
rect 19054 8296 19094 8336
rect 19136 8296 19176 8336
rect 4928 7540 4968 7580
rect 5010 7540 5050 7580
rect 5092 7540 5132 7580
rect 5174 7540 5214 7580
rect 5256 7540 5296 7580
rect 20048 7540 20088 7580
rect 20130 7540 20170 7580
rect 20212 7540 20252 7580
rect 20294 7540 20334 7580
rect 20376 7540 20416 7580
rect 3688 6784 3728 6824
rect 3770 6784 3810 6824
rect 3852 6784 3892 6824
rect 3934 6784 3974 6824
rect 4016 6784 4056 6824
rect 18808 6784 18848 6824
rect 18890 6784 18930 6824
rect 18972 6784 19012 6824
rect 19054 6784 19094 6824
rect 19136 6784 19176 6824
rect 19276 6280 19316 6320
rect 4928 6028 4968 6068
rect 5010 6028 5050 6068
rect 5092 6028 5132 6068
rect 5174 6028 5214 6068
rect 5256 6028 5296 6068
rect 20048 6028 20088 6068
rect 20130 6028 20170 6068
rect 20212 6028 20252 6068
rect 20294 6028 20334 6068
rect 20376 6028 20416 6068
rect 19372 5356 19412 5396
rect 3688 5272 3728 5312
rect 3770 5272 3810 5312
rect 3852 5272 3892 5312
rect 3934 5272 3974 5312
rect 4016 5272 4056 5312
rect 18808 5272 18848 5312
rect 18890 5272 18930 5312
rect 18972 5272 19012 5312
rect 19054 5272 19094 5312
rect 19136 5272 19176 5312
rect 4928 4516 4968 4556
rect 5010 4516 5050 4556
rect 5092 4516 5132 4556
rect 5174 4516 5214 4556
rect 5256 4516 5296 4556
rect 20048 4516 20088 4556
rect 20130 4516 20170 4556
rect 20212 4516 20252 4556
rect 20294 4516 20334 4556
rect 20376 4516 20416 4556
rect 3688 3760 3728 3800
rect 3770 3760 3810 3800
rect 3852 3760 3892 3800
rect 3934 3760 3974 3800
rect 4016 3760 4056 3800
rect 18808 3760 18848 3800
rect 18890 3760 18930 3800
rect 18972 3760 19012 3800
rect 19054 3760 19094 3800
rect 19136 3760 19176 3800
rect 4928 3004 4968 3044
rect 5010 3004 5050 3044
rect 5092 3004 5132 3044
rect 5174 3004 5214 3044
rect 5256 3004 5296 3044
rect 20048 3004 20088 3044
rect 20130 3004 20170 3044
rect 20212 3004 20252 3044
rect 20294 3004 20334 3044
rect 20376 3004 20416 3044
rect 3688 2248 3728 2288
rect 3770 2248 3810 2288
rect 3852 2248 3892 2288
rect 3934 2248 3974 2288
rect 4016 2248 4056 2288
rect 18808 2248 18848 2288
rect 18890 2248 18930 2288
rect 18972 2248 19012 2288
rect 19054 2248 19094 2288
rect 19136 2248 19176 2288
rect 4928 1492 4968 1532
rect 5010 1492 5050 1532
rect 5092 1492 5132 1532
rect 5174 1492 5214 1532
rect 5256 1492 5296 1532
rect 20048 1492 20088 1532
rect 20130 1492 20170 1532
rect 20212 1492 20252 1532
rect 20294 1492 20334 1532
rect 20376 1492 20416 1532
<< metal5 >>
rect 3652 9848 4092 11844
rect 3652 9808 3688 9848
rect 3728 9808 3770 9848
rect 3810 9808 3852 9848
rect 3892 9808 3934 9848
rect 3974 9808 4016 9848
rect 4056 9808 4092 9848
rect 3652 8336 4092 9808
rect 3652 8296 3688 8336
rect 3728 8296 3770 8336
rect 3810 8296 3852 8336
rect 3892 8296 3934 8336
rect 3974 8296 4016 8336
rect 4056 8296 4092 8336
rect 3652 6824 4092 8296
rect 3652 6784 3688 6824
rect 3728 6784 3770 6824
rect 3810 6784 3852 6824
rect 3892 6784 3934 6824
rect 3974 6784 4016 6824
rect 4056 6784 4092 6824
rect 3652 5312 4092 6784
rect 3652 5272 3688 5312
rect 3728 5272 3770 5312
rect 3810 5272 3852 5312
rect 3892 5272 3934 5312
rect 3974 5272 4016 5312
rect 4056 5272 4092 5312
rect 3652 3800 4092 5272
rect 3652 3760 3688 3800
rect 3728 3760 3770 3800
rect 3810 3760 3852 3800
rect 3892 3760 3934 3800
rect 3974 3760 4016 3800
rect 4056 3760 4092 3800
rect 3652 2288 4092 3760
rect 3652 2248 3688 2288
rect 3728 2248 3770 2288
rect 3810 2248 3852 2288
rect 3892 2248 3934 2288
rect 3974 2248 4016 2288
rect 4056 2248 4092 2288
rect 3652 0 4092 2248
rect 4892 9092 5332 11844
rect 4892 9052 4928 9092
rect 4968 9052 5010 9092
rect 5050 9052 5092 9092
rect 5132 9052 5174 9092
rect 5214 9052 5256 9092
rect 5296 9052 5332 9092
rect 4892 7580 5332 9052
rect 4892 7540 4928 7580
rect 4968 7540 5010 7580
rect 5050 7540 5092 7580
rect 5132 7540 5174 7580
rect 5214 7540 5256 7580
rect 5296 7540 5332 7580
rect 4892 6068 5332 7540
rect 4892 6028 4928 6068
rect 4968 6028 5010 6068
rect 5050 6028 5092 6068
rect 5132 6028 5174 6068
rect 5214 6028 5256 6068
rect 5296 6028 5332 6068
rect 4892 4556 5332 6028
rect 4892 4516 4928 4556
rect 4968 4516 5010 4556
rect 5050 4516 5092 4556
rect 5132 4516 5174 4556
rect 5214 4516 5256 4556
rect 5296 4516 5332 4556
rect 4892 3044 5332 4516
rect 4892 3004 4928 3044
rect 4968 3004 5010 3044
rect 5050 3004 5092 3044
rect 5132 3004 5174 3044
rect 5214 3004 5256 3044
rect 5296 3004 5332 3044
rect 4892 1532 5332 3004
rect 4892 1492 4928 1532
rect 4968 1492 5010 1532
rect 5050 1492 5092 1532
rect 5132 1492 5174 1532
rect 5214 1492 5256 1532
rect 5296 1492 5332 1532
rect 4892 0 5332 1492
rect 18772 9848 19212 11844
rect 18772 9808 18808 9848
rect 18848 9808 18890 9848
rect 18930 9808 18972 9848
rect 19012 9808 19054 9848
rect 19094 9808 19136 9848
rect 19176 9808 19212 9848
rect 18772 8336 19212 9808
rect 20012 9092 20452 11844
rect 20012 9052 20048 9092
rect 20088 9052 20130 9092
rect 20170 9052 20212 9092
rect 20252 9052 20294 9092
rect 20334 9052 20376 9092
rect 20416 9052 20452 9092
rect 18772 8296 18808 8336
rect 18848 8296 18890 8336
rect 18930 8296 18972 8336
rect 19012 8296 19054 8336
rect 19094 8296 19136 8336
rect 19176 8296 19212 8336
rect 18772 6824 19212 8296
rect 18772 6784 18808 6824
rect 18848 6784 18890 6824
rect 18930 6784 18972 6824
rect 19012 6784 19054 6824
rect 19094 6784 19136 6824
rect 19176 6784 19212 6824
rect 18772 5312 19212 6784
rect 19276 8672 19316 8681
rect 19276 6320 19316 8632
rect 19276 6271 19316 6280
rect 19372 8504 19412 8513
rect 19372 5396 19412 8464
rect 19372 5347 19412 5356
rect 20012 7580 20452 9052
rect 20012 7540 20048 7580
rect 20088 7540 20130 7580
rect 20170 7540 20212 7580
rect 20252 7540 20294 7580
rect 20334 7540 20376 7580
rect 20416 7540 20452 7580
rect 20012 6068 20452 7540
rect 20012 6028 20048 6068
rect 20088 6028 20130 6068
rect 20170 6028 20212 6068
rect 20252 6028 20294 6068
rect 20334 6028 20376 6068
rect 20416 6028 20452 6068
rect 18772 5272 18808 5312
rect 18848 5272 18890 5312
rect 18930 5272 18972 5312
rect 19012 5272 19054 5312
rect 19094 5272 19136 5312
rect 19176 5272 19212 5312
rect 18772 3800 19212 5272
rect 18772 3760 18808 3800
rect 18848 3760 18890 3800
rect 18930 3760 18972 3800
rect 19012 3760 19054 3800
rect 19094 3760 19136 3800
rect 19176 3760 19212 3800
rect 18772 2288 19212 3760
rect 18772 2248 18808 2288
rect 18848 2248 18890 2288
rect 18930 2248 18972 2288
rect 19012 2248 19054 2288
rect 19094 2248 19136 2288
rect 19176 2248 19212 2288
rect 18772 0 19212 2248
rect 20012 4556 20452 6028
rect 20012 4516 20048 4556
rect 20088 4516 20130 4556
rect 20170 4516 20212 4556
rect 20252 4516 20294 4556
rect 20334 4516 20376 4556
rect 20416 4516 20452 4556
rect 20012 3044 20452 4516
rect 20012 3004 20048 3044
rect 20088 3004 20130 3044
rect 20170 3004 20212 3044
rect 20252 3004 20294 3044
rect 20334 3004 20376 3044
rect 20416 3004 20452 3044
rect 20012 1532 20452 3004
rect 20012 1492 20048 1532
rect 20088 1492 20130 1532
rect 20170 1492 20212 1532
rect 20252 1492 20294 1532
rect 20334 1492 20376 1532
rect 20416 1492 20452 1532
rect 20012 0 20452 1492
use sg13g2_buf_1  _00_
timestamp 1676381911
transform 1 0 8448 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  _01_
timestamp 1676381911
transform 1 0 17088 0 -1 3024
box -48 -56 432 834
use sg13g2_buf_1  _02_
timestamp 1676381911
transform 1 0 14880 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  _03_
timestamp 1676381911
transform 1 0 16896 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  _04_
timestamp 1676381911
transform 1 0 9888 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  _05_
timestamp 1676381911
transform 1 0 18048 0 -1 3024
box -48 -56 432 834
use sg13g2_buf_1  _06_
timestamp 1676381911
transform 1 0 19296 0 -1 3024
box -48 -56 432 834
use sg13g2_buf_1  _07_
timestamp 1676381911
transform 1 0 15264 0 1 1512
box -48 -56 432 834
use sg13g2_buf_1  _08_
timestamp 1676381911
transform 1 0 18240 0 1 1512
box -48 -56 432 834
use sg13g2_buf_1  _09_
timestamp 1676381911
transform 1 0 10560 0 -1 6048
box -48 -56 432 834
use sg13g2_buf_1  _10_
timestamp 1676381911
transform 1 0 19488 0 -1 4536
box -48 -56 432 834
use sg13g2_buf_1  _11_
timestamp 1676381911
transform 1 0 18720 0 -1 4536
box -48 -56 432 834
use sg13g2_buf_1  _12_
timestamp 1676381911
transform -1 0 19392 0 1 4536
box -48 -56 432 834
use sg13g2_buf_1  _13_
timestamp 1676381911
transform 1 0 13728 0 1 4536
box -48 -56 432 834
use sg13g2_buf_1  _14_
timestamp 1676381911
transform 1 0 9216 0 -1 6048
box -48 -56 432 834
use sg13g2_buf_1  _15_
timestamp 1676381911
transform 1 0 14592 0 1 6048
box -48 -56 432 834
use sg13g2_buf_1  _16_
timestamp 1676381911
transform 1 0 12768 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  _17_
timestamp 1676381911
transform 1 0 19200 0 -1 9072
box -48 -56 432 834
use sg13g2_buf_1  _18_
timestamp 1676381911
transform 1 0 14496 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  _19_
timestamp 1676381911
transform 1 0 19008 0 -1 7560
box -48 -56 432 834
use sg13g2_buf_1  _20_
timestamp 1676381911
transform 1 0 18720 0 -1 6048
box -48 -56 432 834
use sg13g2_buf_1  _21_
timestamp 1676381911
transform 1 0 19104 0 1 6048
box -48 -56 432 834
use sg13g2_buf_1  _22_
timestamp 1676381911
transform 1 0 15072 0 -1 4536
box -48 -56 432 834
use sg13g2_buf_1  _23_
timestamp 1676381911
transform -1 0 19488 0 -1 6048
box -48 -56 432 834
use sg13g2_buf_1  _24_
timestamp 1676381911
transform 1 0 15936 0 1 4536
box -48 -56 432 834
use sg13g2_buf_1  _25_
timestamp 1676381911
transform 1 0 16128 0 -1 9072
box -48 -56 432 834
use sg13g2_buf_1  _26_
timestamp 1676381911
transform 1 0 11808 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  _27_
timestamp 1676381911
transform 1 0 15744 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  _28_
timestamp 1676381911
transform 1 0 16512 0 -1 9072
box -48 -56 432 834
use sg13g2_buf_1  _29_
timestamp 1676381911
transform -1 0 18048 0 -1 9072
box -48 -56 432 834
use sg13g2_buf_1  _30_
timestamp 1676381911
transform -1 0 18432 0 -1 9072
box -48 -56 432 834
use sg13g2_buf_1  _31_
timestamp 1676381911
transform -1 0 20352 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  _32_
timestamp 1676381911
transform 1 0 1824 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  _33_
timestamp 1676381911
transform 1 0 3264 0 1 6048
box -48 -56 432 834
use sg13g2_buf_1  _34_
timestamp 1676381911
transform 1 0 5568 0 -1 7560
box -48 -56 432 834
use sg13g2_buf_1  _35_
timestamp 1676381911
transform 1 0 4320 0 1 6048
box -48 -56 432 834
use sg13g2_buf_1  _36_
timestamp 1676381911
transform 1 0 5088 0 1 4536
box -48 -56 432 834
use sg13g2_buf_1  _37_
timestamp 1676381911
transform 1 0 6240 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  _38_
timestamp 1676381911
transform 1 0 6528 0 -1 3024
box -48 -56 432 834
use sg13g2_buf_1  _39_
timestamp 1676381911
transform 1 0 8832 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  _40_
timestamp 1676381911
transform 1 0 10656 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  _41_
timestamp 1676381911
transform 1 0 12000 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  _42_
timestamp 1676381911
transform 1 0 13344 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  _43_
timestamp 1676381911
transform 1 0 10944 0 -1 6048
box -48 -56 432 834
use sg13g2_buf_1  _44_
timestamp 1676381911
transform 1 0 11808 0 -1 4536
box -48 -56 432 834
use sg13g2_buf_1  _45_
timestamp 1676381911
transform 1 0 12000 0 -1 6048
box -48 -56 432 834
use sg13g2_buf_1  _46_
timestamp 1676381911
transform 1 0 13248 0 -1 9072
box -48 -56 432 834
use sg13g2_buf_1  _47_
timestamp 1676381911
transform 1 0 13728 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  _48_
timestamp 1676381911
transform 1 0 12864 0 1 1512
box -48 -56 432 834
use sg13g2_buf_1  _49_
timestamp 1676381911
transform 1 0 14880 0 -1 6048
box -48 -56 432 834
use sg13g2_buf_1  _50_
timestamp 1676381911
transform 1 0 16512 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  _51_
timestamp 1676381911
transform -1 0 19488 0 -1 4536
box -48 -56 432 834
use sg13g2_buf_1  _52_
timestamp 1676381911
transform -1 0 2304 0 -1 9072
box -48 -56 432 834
use sg13g2_buf_1  _53_
timestamp 1676381911
transform -1 0 2688 0 -1 9072
box -48 -56 432 834
use sg13g2_buf_1  _54_
timestamp 1676381911
transform -1 0 4704 0 -1 7560
box -48 -56 432 834
use sg13g2_buf_1  _55_
timestamp 1676381911
transform -1 0 5568 0 -1 7560
box -48 -56 432 834
use sg13g2_buf_1  _56_
timestamp 1676381911
transform -1 0 3072 0 -1 9072
box -48 -56 432 834
use sg13g2_buf_1  _57_
timestamp 1676381911
transform -1 0 2304 0 -1 7560
box -48 -56 432 834
use sg13g2_buf_1  _58_
timestamp 1676381911
transform -1 0 3552 0 -1 6048
box -48 -56 432 834
use sg13g2_buf_1  _59_
timestamp 1676381911
transform -1 0 4896 0 -1 6048
box -48 -56 432 834
use sg13g2_buf_1  _60_
timestamp 1676381911
transform -1 0 5952 0 -1 6048
box -48 -56 432 834
use sg13g2_buf_1  _61_
timestamp 1676381911
transform -1 0 7008 0 1 4536
box -48 -56 432 834
use sg13g2_buf_1  _62_
timestamp 1676381911
transform -1 0 7968 0 1 4536
box -48 -56 432 834
use sg13g2_buf_1  _63_
timestamp 1676381911
transform -1 0 8448 0 1 4536
box -48 -56 432 834
use sg13g2_buf_1  _64_
timestamp 1676381911
transform -1 0 4224 0 -1 4536
box -48 -56 432 834
use sg13g2_buf_1  _65_
timestamp 1676381911
transform -1 0 7392 0 1 4536
box -48 -56 432 834
use sg13g2_buf_1  _66_
timestamp 1676381911
transform -1 0 8640 0 -1 6048
box -48 -56 432 834
use sg13g2_buf_1  _67_
timestamp 1676381911
transform -1 0 9504 0 1 6048
box -48 -56 432 834
use sg13g2_buf_1  _68_
timestamp 1676381911
transform -1 0 10656 0 -1 7560
box -48 -56 432 834
use sg13g2_buf_1  _69_
timestamp 1676381911
transform -1 0 10272 0 -1 7560
box -48 -56 432 834
use sg13g2_buf_1  _70_
timestamp 1676381911
transform -1 0 10272 0 1 7560
box -48 -56 432 834
use sg13g2_buf_1  _71_
timestamp 1676381911
transform -1 0 10656 0 1 7560
box -48 -56 432 834
use sg13g2_buf_1  _72_
timestamp 1676381911
transform -1 0 18528 0 1 7560
box -48 -56 432 834
use sg13g2_buf_1  _73_
timestamp 1676381911
transform -1 0 19968 0 -1 9072
box -48 -56 432 834
use sg13g2_buf_1  _74_
timestamp 1676381911
transform -1 0 19776 0 -1 7560
box -48 -56 432 834
use sg13g2_buf_1  _75_
timestamp 1676381911
transform -1 0 19872 0 1 6048
box -48 -56 432 834
use sg13g2_buf_1  _76_
timestamp 1676381911
transform -1 0 18240 0 -1 7560
box -48 -56 432 834
use sg13g2_buf_1  _77_
timestamp 1676381911
transform -1 0 18336 0 -1 6048
box -48 -56 432 834
use sg13g2_buf_1  _78_
timestamp 1676381911
transform -1 0 17376 0 -1 7560
box -48 -56 432 834
use sg13g2_buf_1  _79_
timestamp 1676381911
transform -1 0 16992 0 -1 7560
box -48 -56 432 834
use sg13g2_buf_1  _80_
timestamp 1676381911
transform -1 0 16416 0 -1 7560
box -48 -56 432 834
use sg13g2_buf_1  _81_
timestamp 1676381911
transform -1 0 15744 0 -1 7560
box -48 -56 432 834
use sg13g2_buf_1  _82_
timestamp 1676381911
transform -1 0 13056 0 1 6048
box -48 -56 432 834
use sg13g2_buf_1  _83_
timestamp 1676381911
transform -1 0 12576 0 -1 7560
box -48 -56 432 834
use sg13g2_buf_1  _84_
timestamp 1676381911
transform -1 0 12192 0 -1 7560
box -48 -56 432 834
use sg13g2_buf_1  _85_
timestamp 1676381911
transform -1 0 13440 0 1 6048
box -48 -56 432 834
use sg13g2_buf_1  _86_
timestamp 1676381911
transform -1 0 13920 0 -1 7560
box -48 -56 432 834
use sg13g2_buf_1  _87_
timestamp 1676381911
transform -1 0 14304 0 -1 7560
box -48 -56 432 834
use sg13g2_buf_1  _88_
timestamp 1676381911
transform 1 0 3648 0 1 4536
box -48 -56 432 834
use sg13g2_decap_8  FILLER_0_0
timestamp 1679581782
transform 1 0 1152 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_7
timestamp 1679581782
transform 1 0 1824 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_14
timestamp 1679581782
transform 1 0 2496 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_21
timestamp 1679581782
transform 1 0 3168 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_28
timestamp 1679581782
transform 1 0 3840 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_35
timestamp 1679581782
transform 1 0 4512 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_42
timestamp 1679581782
transform 1 0 5184 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_49
timestamp 1679581782
transform 1 0 5856 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_56
timestamp 1679581782
transform 1 0 6528 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_63
timestamp 1679581782
transform 1 0 7200 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_70
timestamp 1679581782
transform 1 0 7872 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_77
timestamp 1679581782
transform 1 0 8544 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_84
timestamp 1679581782
transform 1 0 9216 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_91
timestamp 1679581782
transform 1 0 9888 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_98
timestamp 1679581782
transform 1 0 10560 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_105
timestamp 1679581782
transform 1 0 11232 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_112
timestamp 1679581782
transform 1 0 11904 0 1 1512
box -48 -56 720 834
use sg13g2_fill_2  FILLER_0_119
timestamp 1677580104
transform 1 0 12576 0 1 1512
box -48 -56 240 834
use sg13g2_fill_1  FILLER_0_121
timestamp 1677579658
transform 1 0 12768 0 1 1512
box -48 -56 144 834
use sg13g2_decap_8  FILLER_0_126
timestamp 1679581782
transform 1 0 13248 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_133
timestamp 1679581782
transform 1 0 13920 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_140
timestamp 1679581782
transform 1 0 14592 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_151
timestamp 1679581782
transform 1 0 15648 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_158
timestamp 1679581782
transform 1 0 16320 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_165
timestamp 1679581782
transform 1 0 16992 0 1 1512
box -48 -56 720 834
use sg13g2_fill_2  FILLER_0_172
timestamp 1677580104
transform 1 0 17664 0 1 1512
box -48 -56 240 834
use sg13g2_fill_2  FILLER_0_182
timestamp 1677580104
transform 1 0 18624 0 1 1512
box -48 -56 240 834
use sg13g2_fill_1  FILLER_0_184
timestamp 1677579658
transform 1 0 18816 0 1 1512
box -48 -56 144 834
use sg13g2_decap_8  FILLER_1_0
timestamp 1679581782
transform 1 0 1152 0 -1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_7
timestamp 1679581782
transform 1 0 1824 0 -1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_14
timestamp 1679581782
transform 1 0 2496 0 -1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_21
timestamp 1679581782
transform 1 0 3168 0 -1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_28
timestamp 1679581782
transform 1 0 3840 0 -1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_35
timestamp 1679581782
transform 1 0 4512 0 -1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_42
timestamp 1679581782
transform 1 0 5184 0 -1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_49
timestamp 1679581782
transform 1 0 5856 0 -1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_60
timestamp 1679581782
transform 1 0 6912 0 -1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_67
timestamp 1679581782
transform 1 0 7584 0 -1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_74
timestamp 1679581782
transform 1 0 8256 0 -1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_81
timestamp 1679581782
transform 1 0 8928 0 -1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_88
timestamp 1679581782
transform 1 0 9600 0 -1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_95
timestamp 1679581782
transform 1 0 10272 0 -1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_102
timestamp 1679581782
transform 1 0 10944 0 -1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_109
timestamp 1679581782
transform 1 0 11616 0 -1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_116
timestamp 1679581782
transform 1 0 12288 0 -1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_123
timestamp 1679581782
transform 1 0 12960 0 -1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_130
timestamp 1679581782
transform 1 0 13632 0 -1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_137
timestamp 1679581782
transform 1 0 14304 0 -1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_144
timestamp 1679581782
transform 1 0 14976 0 -1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_151
timestamp 1679581782
transform 1 0 15648 0 -1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_158
timestamp 1679581782
transform 1 0 16320 0 -1 3024
box -48 -56 720 834
use sg13g2_fill_1  FILLER_1_165
timestamp 1677579658
transform 1 0 16992 0 -1 3024
box -48 -56 144 834
use sg13g2_decap_4  FILLER_1_170
timestamp 1679577901
transform 1 0 17472 0 -1 3024
box -48 -56 432 834
use sg13g2_fill_2  FILLER_1_174
timestamp 1677580104
transform 1 0 17856 0 -1 3024
box -48 -56 240 834
use sg13g2_fill_1  FILLER_1_180
timestamp 1677579658
transform 1 0 18432 0 -1 3024
box -48 -56 144 834
use sg13g2_decap_8  FILLER_2_0
timestamp 1679581782
transform 1 0 1152 0 1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_11
timestamp 1679581782
transform 1 0 2208 0 1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_18
timestamp 1679581782
transform 1 0 2880 0 1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_25
timestamp 1679581782
transform 1 0 3552 0 1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_32
timestamp 1679581782
transform 1 0 4224 0 1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_39
timestamp 1679581782
transform 1 0 4896 0 1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_46
timestamp 1679581782
transform 1 0 5568 0 1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_57
timestamp 1679581782
transform 1 0 6624 0 1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_64
timestamp 1679581782
transform 1 0 7296 0 1 3024
box -48 -56 720 834
use sg13g2_decap_4  FILLER_2_71
timestamp 1679577901
transform 1 0 7968 0 1 3024
box -48 -56 432 834
use sg13g2_fill_1  FILLER_2_75
timestamp 1677579658
transform 1 0 8352 0 1 3024
box -48 -56 144 834
use sg13g2_decap_8  FILLER_2_84
timestamp 1679581782
transform 1 0 9216 0 1 3024
box -48 -56 720 834
use sg13g2_decap_4  FILLER_2_95
timestamp 1679577901
transform 1 0 10272 0 1 3024
box -48 -56 432 834
use sg13g2_decap_8  FILLER_2_103
timestamp 1679581782
transform 1 0 11040 0 1 3024
box -48 -56 720 834
use sg13g2_fill_2  FILLER_2_110
timestamp 1677580104
transform 1 0 11712 0 1 3024
box -48 -56 240 834
use sg13g2_fill_1  FILLER_2_112
timestamp 1677579658
transform 1 0 11904 0 1 3024
box -48 -56 144 834
use sg13g2_decap_8  FILLER_2_117
timestamp 1679581782
transform 1 0 12384 0 1 3024
box -48 -56 720 834
use sg13g2_fill_2  FILLER_2_124
timestamp 1677580104
transform 1 0 13056 0 1 3024
box -48 -56 240 834
use sg13g2_fill_1  FILLER_2_126
timestamp 1677579658
transform 1 0 13248 0 1 3024
box -48 -56 144 834
use sg13g2_decap_8  FILLER_2_135
timestamp 1679581782
transform 1 0 14112 0 1 3024
box -48 -56 720 834
use sg13g2_fill_1  FILLER_2_142
timestamp 1677579658
transform 1 0 14784 0 1 3024
box -48 -56 144 834
use sg13g2_decap_8  FILLER_2_147
timestamp 1679581782
transform 1 0 15264 0 1 3024
box -48 -56 720 834
use sg13g2_decap_4  FILLER_2_154
timestamp 1679577901
transform 1 0 15936 0 1 3024
box -48 -56 432 834
use sg13g2_fill_2  FILLER_2_158
timestamp 1677580104
transform 1 0 16320 0 1 3024
box -48 -56 240 834
use sg13g2_decap_8  FILLER_2_168
timestamp 1679581782
transform 1 0 17280 0 1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_175
timestamp 1679581782
transform 1 0 17952 0 1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_182
timestamp 1679581782
transform 1 0 18624 0 1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_0
timestamp 1679581782
transform 1 0 1152 0 -1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_7
timestamp 1679581782
transform 1 0 1824 0 -1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_14
timestamp 1679581782
transform 1 0 2496 0 -1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_21
timestamp 1679581782
transform 1 0 3168 0 -1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_32
timestamp 1679581782
transform 1 0 4224 0 -1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_39
timestamp 1679581782
transform 1 0 4896 0 -1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_46
timestamp 1679581782
transform 1 0 5568 0 -1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_53
timestamp 1679581782
transform 1 0 6240 0 -1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_60
timestamp 1679581782
transform 1 0 6912 0 -1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_67
timestamp 1679581782
transform 1 0 7584 0 -1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_74
timestamp 1679581782
transform 1 0 8256 0 -1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_81
timestamp 1679581782
transform 1 0 8928 0 -1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_88
timestamp 1679581782
transform 1 0 9600 0 -1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_95
timestamp 1679581782
transform 1 0 10272 0 -1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_102
timestamp 1679581782
transform 1 0 10944 0 -1 4536
box -48 -56 720 834
use sg13g2_fill_2  FILLER_3_109
timestamp 1677580104
transform 1 0 11616 0 -1 4536
box -48 -56 240 834
use sg13g2_decap_8  FILLER_3_115
timestamp 1679581782
transform 1 0 12192 0 -1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_122
timestamp 1679581782
transform 1 0 12864 0 -1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_129
timestamp 1679581782
transform 1 0 13536 0 -1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_136
timestamp 1679581782
transform 1 0 14208 0 -1 4536
box -48 -56 720 834
use sg13g2_fill_2  FILLER_3_143
timestamp 1677580104
transform 1 0 14880 0 -1 4536
box -48 -56 240 834
use sg13g2_decap_8  FILLER_3_149
timestamp 1679581782
transform 1 0 15456 0 -1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_156
timestamp 1679581782
transform 1 0 16128 0 -1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_163
timestamp 1679581782
transform 1 0 16800 0 -1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_170
timestamp 1679581782
transform 1 0 17472 0 -1 4536
box -48 -56 720 834
use sg13g2_decap_4  FILLER_3_177
timestamp 1679577901
transform 1 0 18144 0 -1 4536
box -48 -56 432 834
use sg13g2_fill_2  FILLER_3_181
timestamp 1677580104
transform 1 0 18528 0 -1 4536
box -48 -56 240 834
use sg13g2_fill_2  FILLER_3_195
timestamp 1677580104
transform 1 0 19872 0 -1 4536
box -48 -56 240 834
use sg13g2_decap_8  FILLER_4_0
timestamp 1679581782
transform 1 0 1152 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_7
timestamp 1679581782
transform 1 0 1824 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_14
timestamp 1679581782
transform 1 0 2496 0 1 4536
box -48 -56 720 834
use sg13g2_decap_4  FILLER_4_21
timestamp 1679577901
transform 1 0 3168 0 1 4536
box -48 -56 432 834
use sg13g2_fill_1  FILLER_4_25
timestamp 1677579658
transform 1 0 3552 0 1 4536
box -48 -56 144 834
use sg13g2_decap_8  FILLER_4_30
timestamp 1679581782
transform 1 0 4032 0 1 4536
box -48 -56 720 834
use sg13g2_decap_4  FILLER_4_37
timestamp 1679577901
transform 1 0 4704 0 1 4536
box -48 -56 432 834
use sg13g2_decap_8  FILLER_4_45
timestamp 1679581782
transform 1 0 5472 0 1 4536
box -48 -56 720 834
use sg13g2_decap_4  FILLER_4_52
timestamp 1679577901
transform 1 0 6144 0 1 4536
box -48 -56 432 834
use sg13g2_fill_1  FILLER_4_56
timestamp 1677579658
transform 1 0 6528 0 1 4536
box -48 -56 144 834
use sg13g2_fill_2  FILLER_4_65
timestamp 1677580104
transform 1 0 7392 0 1 4536
box -48 -56 240 834
use sg13g2_fill_1  FILLER_4_71
timestamp 1677579658
transform 1 0 7968 0 1 4536
box -48 -56 144 834
use sg13g2_decap_8  FILLER_4_76
timestamp 1679581782
transform 1 0 8448 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_83
timestamp 1679581782
transform 1 0 9120 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_90
timestamp 1679581782
transform 1 0 9792 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_97
timestamp 1679581782
transform 1 0 10464 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_104
timestamp 1679581782
transform 1 0 11136 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_111
timestamp 1679581782
transform 1 0 11808 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_118
timestamp 1679581782
transform 1 0 12480 0 1 4536
box -48 -56 720 834
use sg13g2_decap_4  FILLER_4_125
timestamp 1679577901
transform 1 0 13152 0 1 4536
box -48 -56 432 834
use sg13g2_fill_2  FILLER_4_129
timestamp 1677580104
transform 1 0 13536 0 1 4536
box -48 -56 240 834
use sg13g2_decap_8  FILLER_4_135
timestamp 1679581782
transform 1 0 14112 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_142
timestamp 1679581782
transform 1 0 14784 0 1 4536
box -48 -56 720 834
use sg13g2_decap_4  FILLER_4_149
timestamp 1679577901
transform 1 0 15456 0 1 4536
box -48 -56 432 834
use sg13g2_fill_1  FILLER_4_153
timestamp 1677579658
transform 1 0 15840 0 1 4536
box -48 -56 144 834
use sg13g2_decap_8  FILLER_4_158
timestamp 1679581782
transform 1 0 16320 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_165
timestamp 1679581782
transform 1 0 16992 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_172
timestamp 1679581782
transform 1 0 17664 0 1 4536
box -48 -56 720 834
use sg13g2_fill_2  FILLER_4_179
timestamp 1677580104
transform 1 0 18336 0 1 4536
box -48 -56 240 834
use sg13g2_fill_1  FILLER_4_181
timestamp 1677579658
transform 1 0 18528 0 1 4536
box -48 -56 144 834
use sg13g2_fill_2  FILLER_4_190
timestamp 1677580104
transform 1 0 19392 0 1 4536
box -48 -56 240 834
use sg13g2_fill_1  FILLER_4_192
timestamp 1677579658
transform 1 0 19584 0 1 4536
box -48 -56 144 834
use sg13g2_decap_8  FILLER_5_0
timestamp 1679581782
transform 1 0 1152 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_7
timestamp 1679581782
transform 1 0 1824 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_14
timestamp 1679581782
transform 1 0 2496 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_25
timestamp 1679581782
transform 1 0 3552 0 -1 6048
box -48 -56 720 834
use sg13g2_fill_2  FILLER_5_32
timestamp 1677580104
transform 1 0 4224 0 -1 6048
box -48 -56 240 834
use sg13g2_fill_1  FILLER_5_34
timestamp 1677579658
transform 1 0 4416 0 -1 6048
box -48 -56 144 834
use sg13g2_decap_8  FILLER_5_39
timestamp 1679581782
transform 1 0 4896 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_50
timestamp 1679581782
transform 1 0 5952 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_57
timestamp 1679581782
transform 1 0 6624 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_64
timestamp 1679581782
transform 1 0 7296 0 -1 6048
box -48 -56 720 834
use sg13g2_fill_2  FILLER_5_71
timestamp 1677580104
transform 1 0 7968 0 -1 6048
box -48 -56 240 834
use sg13g2_fill_1  FILLER_5_73
timestamp 1677579658
transform 1 0 8160 0 -1 6048
box -48 -56 144 834
use sg13g2_decap_4  FILLER_5_78
timestamp 1679577901
transform 1 0 8640 0 -1 6048
box -48 -56 432 834
use sg13g2_fill_2  FILLER_5_82
timestamp 1677580104
transform 1 0 9024 0 -1 6048
box -48 -56 240 834
use sg13g2_decap_8  FILLER_5_88
timestamp 1679581782
transform 1 0 9600 0 -1 6048
box -48 -56 720 834
use sg13g2_fill_2  FILLER_5_95
timestamp 1677580104
transform 1 0 10272 0 -1 6048
box -48 -56 240 834
use sg13g2_fill_1  FILLER_5_97
timestamp 1677579658
transform 1 0 10464 0 -1 6048
box -48 -56 144 834
use sg13g2_decap_8  FILLER_5_106
timestamp 1679581782
transform 1 0 11328 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_117
timestamp 1679581782
transform 1 0 12384 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_124
timestamp 1679581782
transform 1 0 13056 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_131
timestamp 1679581782
transform 1 0 13728 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_4  FILLER_5_138
timestamp 1679577901
transform 1 0 14400 0 -1 6048
box -48 -56 432 834
use sg13g2_fill_1  FILLER_5_142
timestamp 1677579658
transform 1 0 14784 0 -1 6048
box -48 -56 144 834
use sg13g2_decap_8  FILLER_5_147
timestamp 1679581782
transform 1 0 15264 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_154
timestamp 1679581782
transform 1 0 15936 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_161
timestamp 1679581782
transform 1 0 16608 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_168
timestamp 1679581782
transform 1 0 17280 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_4  FILLER_5_179
timestamp 1679577901
transform 1 0 18336 0 -1 6048
box -48 -56 432 834
use sg13g2_fill_2  FILLER_5_191
timestamp 1677580104
transform 1 0 19488 0 -1 6048
box -48 -56 240 834
use sg13g2_decap_8  FILLER_6_0
timestamp 1679581782
transform 1 0 1152 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_7
timestamp 1679581782
transform 1 0 1824 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_14
timestamp 1679581782
transform 1 0 2496 0 1 6048
box -48 -56 720 834
use sg13g2_fill_1  FILLER_6_21
timestamp 1677579658
transform 1 0 3168 0 1 6048
box -48 -56 144 834
use sg13g2_decap_8  FILLER_6_26
timestamp 1679581782
transform 1 0 3648 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_37
timestamp 1679581782
transform 1 0 4704 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_44
timestamp 1679581782
transform 1 0 5376 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_51
timestamp 1679581782
transform 1 0 6048 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_58
timestamp 1679581782
transform 1 0 6720 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_65
timestamp 1679581782
transform 1 0 7392 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_72
timestamp 1679581782
transform 1 0 8064 0 1 6048
box -48 -56 720 834
use sg13g2_decap_4  FILLER_6_79
timestamp 1679577901
transform 1 0 8736 0 1 6048
box -48 -56 432 834
use sg13g2_decap_8  FILLER_6_87
timestamp 1679581782
transform 1 0 9504 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_94
timestamp 1679581782
transform 1 0 10176 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_101
timestamp 1679581782
transform 1 0 10848 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_108
timestamp 1679581782
transform 1 0 11520 0 1 6048
box -48 -56 720 834
use sg13g2_decap_4  FILLER_6_115
timestamp 1679577901
transform 1 0 12192 0 1 6048
box -48 -56 432 834
use sg13g2_fill_1  FILLER_6_119
timestamp 1677579658
transform 1 0 12576 0 1 6048
box -48 -56 144 834
use sg13g2_decap_8  FILLER_6_128
timestamp 1679581782
transform 1 0 13440 0 1 6048
box -48 -56 720 834
use sg13g2_decap_4  FILLER_6_135
timestamp 1679577901
transform 1 0 14112 0 1 6048
box -48 -56 432 834
use sg13g2_fill_1  FILLER_6_139
timestamp 1677579658
transform 1 0 14496 0 1 6048
box -48 -56 144 834
use sg13g2_decap_8  FILLER_6_144
timestamp 1679581782
transform 1 0 14976 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_151
timestamp 1679581782
transform 1 0 15648 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_158
timestamp 1679581782
transform 1 0 16320 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_165
timestamp 1679581782
transform 1 0 16992 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_172
timestamp 1679581782
transform 1 0 17664 0 1 6048
box -48 -56 720 834
use sg13g2_fill_2  FILLER_6_195
timestamp 1677580104
transform 1 0 19872 0 1 6048
box -48 -56 240 834
use sg13g2_decap_8  FILLER_7_0
timestamp 1679581782
transform 1 0 1152 0 -1 7560
box -48 -56 720 834
use sg13g2_fill_1  FILLER_7_7
timestamp 1677579658
transform 1 0 1824 0 -1 7560
box -48 -56 144 834
use sg13g2_decap_8  FILLER_7_12
timestamp 1679581782
transform 1 0 2304 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_19
timestamp 1679581782
transform 1 0 2976 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_26
timestamp 1679581782
transform 1 0 3648 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_4  FILLER_7_37
timestamp 1679577901
transform 1 0 4704 0 -1 7560
box -48 -56 432 834
use sg13g2_fill_1  FILLER_7_41
timestamp 1677579658
transform 1 0 5088 0 -1 7560
box -48 -56 144 834
use sg13g2_decap_8  FILLER_7_50
timestamp 1679581782
transform 1 0 5952 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_57
timestamp 1679581782
transform 1 0 6624 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_64
timestamp 1679581782
transform 1 0 7296 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_71
timestamp 1679581782
transform 1 0 7968 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_78
timestamp 1679581782
transform 1 0 8640 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_4  FILLER_7_85
timestamp 1679577901
transform 1 0 9312 0 -1 7560
box -48 -56 432 834
use sg13g2_fill_2  FILLER_7_89
timestamp 1677580104
transform 1 0 9696 0 -1 7560
box -48 -56 240 834
use sg13g2_decap_8  FILLER_7_99
timestamp 1679581782
transform 1 0 10656 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_4  FILLER_7_106
timestamp 1679577901
transform 1 0 11328 0 -1 7560
box -48 -56 432 834
use sg13g2_fill_1  FILLER_7_110
timestamp 1677579658
transform 1 0 11712 0 -1 7560
box -48 -56 144 834
use sg13g2_decap_8  FILLER_7_119
timestamp 1679581782
transform 1 0 12576 0 -1 7560
box -48 -56 720 834
use sg13g2_fill_2  FILLER_7_126
timestamp 1677580104
transform 1 0 13248 0 -1 7560
box -48 -56 240 834
use sg13g2_fill_1  FILLER_7_128
timestamp 1677579658
transform 1 0 13440 0 -1 7560
box -48 -56 144 834
use sg13g2_decap_8  FILLER_7_137
timestamp 1679581782
transform 1 0 14304 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_4  FILLER_7_144
timestamp 1679577901
transform 1 0 14976 0 -1 7560
box -48 -56 432 834
use sg13g2_fill_2  FILLER_7_152
timestamp 1677580104
transform 1 0 15744 0 -1 7560
box -48 -56 240 834
use sg13g2_fill_1  FILLER_7_154
timestamp 1677579658
transform 1 0 15936 0 -1 7560
box -48 -56 144 834
use sg13g2_fill_2  FILLER_7_159
timestamp 1677580104
transform 1 0 16416 0 -1 7560
box -48 -56 240 834
use sg13g2_fill_1  FILLER_7_169
timestamp 1677579658
transform 1 0 17376 0 -1 7560
box -48 -56 144 834
use sg13g2_fill_2  FILLER_7_194
timestamp 1677580104
transform 1 0 19776 0 -1 7560
box -48 -56 240 834
use sg13g2_fill_1  FILLER_7_196
timestamp 1677579658
transform 1 0 19968 0 -1 7560
box -48 -56 144 834
use sg13g2_decap_8  FILLER_8_0
timestamp 1679581782
transform 1 0 1152 0 1 7560
box -48 -56 720 834
use sg13g2_fill_2  FILLER_8_7
timestamp 1677580104
transform 1 0 1824 0 1 7560
box -48 -56 240 834
use sg13g2_decap_8  FILLER_8_13
timestamp 1679581782
transform 1 0 2400 0 1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_20
timestamp 1679581782
transform 1 0 3072 0 1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_27
timestamp 1679581782
transform 1 0 3744 0 1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_34
timestamp 1679581782
transform 1 0 4416 0 1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_41
timestamp 1679581782
transform 1 0 5088 0 1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_48
timestamp 1679581782
transform 1 0 5760 0 1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_55
timestamp 1679581782
transform 1 0 6432 0 1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_62
timestamp 1679581782
transform 1 0 7104 0 1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_69
timestamp 1679581782
transform 1 0 7776 0 1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_76
timestamp 1679581782
transform 1 0 8448 0 1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_83
timestamp 1679581782
transform 1 0 9120 0 1 7560
box -48 -56 720 834
use sg13g2_fill_1  FILLER_8_90
timestamp 1677579658
transform 1 0 9792 0 1 7560
box -48 -56 144 834
use sg13g2_decap_8  FILLER_8_99
timestamp 1679581782
transform 1 0 10656 0 1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_106
timestamp 1679581782
transform 1 0 11328 0 1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_113
timestamp 1679581782
transform 1 0 12000 0 1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_120
timestamp 1679581782
transform 1 0 12672 0 1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_127
timestamp 1679581782
transform 1 0 13344 0 1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_134
timestamp 1679581782
transform 1 0 14016 0 1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_141
timestamp 1679581782
transform 1 0 14688 0 1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_148
timestamp 1679581782
transform 1 0 15360 0 1 7560
box -48 -56 720 834
use sg13g2_fill_2  FILLER_8_155
timestamp 1677580104
transform 1 0 16032 0 1 7560
box -48 -56 240 834
use sg13g2_fill_1  FILLER_9_20
timestamp 1677579658
transform 1 0 3072 0 -1 9072
box -48 -56 144 834
use sg13g2_decap_8  FILLER_9_69
timestamp 1679581782
transform 1 0 7776 0 -1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_76
timestamp 1679581782
transform 1 0 8448 0 -1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_83
timestamp 1679581782
transform 1 0 9120 0 -1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_90
timestamp 1679581782
transform 1 0 9792 0 -1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_97
timestamp 1679581782
transform 1 0 10464 0 -1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_104
timestamp 1679581782
transform 1 0 11136 0 -1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_111
timestamp 1679581782
transform 1 0 11808 0 -1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_118
timestamp 1679581782
transform 1 0 12480 0 -1 9072
box -48 -56 720 834
use sg13g2_fill_1  FILLER_9_125
timestamp 1677579658
transform 1 0 13152 0 -1 9072
box -48 -56 144 834
use sg13g2_decap_8  FILLER_9_130
timestamp 1679581782
transform 1 0 13632 0 -1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_137
timestamp 1679581782
transform 1 0 14304 0 -1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_144
timestamp 1679581782
transform 1 0 14976 0 -1 9072
box -48 -56 720 834
use sg13g2_fill_1  FILLER_9_151
timestamp 1677579658
transform 1 0 15648 0 -1 9072
box -48 -56 144 834
use sg13g2_fill_1  FILLER_9_200
timestamp 1677579658
transform 1 0 20352 0 -1 9072
box -48 -56 144 834
use sg13g2_fill_1  FILLER_10_0
timestamp 1677579658
transform 1 0 1152 0 1 9072
box -48 -56 144 834
use sg13g2_decap_8  FILLER_10_85
timestamp 1679581782
transform 1 0 9312 0 1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_92
timestamp 1679581782
transform 1 0 9984 0 1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_99
timestamp 1679581782
transform 1 0 10656 0 1 9072
box -48 -56 720 834
use sg13g2_decap_4  FILLER_10_106
timestamp 1679577901
transform 1 0 11328 0 1 9072
box -48 -56 432 834
use sg13g2_fill_1  FILLER_10_110
timestamp 1677579658
transform 1 0 11712 0 1 9072
box -48 -56 144 834
use sg13g2_decap_4  FILLER_10_115
timestamp 1679577901
transform 1 0 12192 0 1 9072
box -48 -56 432 834
use sg13g2_fill_2  FILLER_10_119
timestamp 1677580104
transform 1 0 12576 0 1 9072
box -48 -56 240 834
use sg13g2_decap_8  FILLER_10_125
timestamp 1679581782
transform 1 0 13152 0 1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_132
timestamp 1679581782
transform 1 0 13824 0 1 9072
box -48 -56 720 834
use sg13g2_fill_1  FILLER_10_143
timestamp 1677579658
transform 1 0 14880 0 1 9072
box -48 -56 144 834
use sg13g2_fill_1  FILLER_10_200
timestamp 1677579658
transform 1 0 20352 0 1 9072
box -48 -56 144 834
use sg13g2_buf_1  output1
timestamp 1676381911
transform 1 0 18912 0 1 1512
box -48 -56 432 834
use sg13g2_buf_1  output2
timestamp 1676381911
transform 1 0 19680 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  output3
timestamp 1676381911
transform 1 0 20064 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  output4
timestamp 1676381911
transform 1 0 18624 0 1 4536
box -48 -56 432 834
use sg13g2_buf_1  output5
timestamp 1676381911
transform 1 0 20064 0 -1 4536
box -48 -56 432 834
use sg13g2_buf_1  output6
timestamp 1676381911
transform 1 0 19680 0 1 4536
box -48 -56 432 834
use sg13g2_buf_1  output7
timestamp 1676381911
transform 1 0 20064 0 1 4536
box -48 -56 432 834
use sg13g2_buf_1  output8
timestamp 1676381911
transform 1 0 19680 0 -1 6048
box -48 -56 432 834
use sg13g2_buf_1  output9
timestamp 1676381911
transform 1 0 20064 0 -1 6048
box -48 -56 432 834
use sg13g2_buf_1  output10
timestamp 1676381911
transform 1 0 20064 0 1 6048
box -48 -56 432 834
use sg13g2_buf_1  output11
timestamp 1676381911
transform 1 0 20064 0 -1 7560
box -48 -56 432 834
use sg13g2_buf_1  output12
timestamp 1676381911
transform 1 0 17856 0 1 1512
box -48 -56 432 834
use sg13g2_buf_1  output13
timestamp 1676381911
transform 1 0 20064 0 1 7560
box -48 -56 432 834
use sg13g2_buf_1  output14
timestamp 1676381911
transform 1 0 19680 0 1 7560
box -48 -56 432 834
use sg13g2_buf_1  output15
timestamp 1676381911
transform 1 0 19296 0 1 7560
box -48 -56 432 834
use sg13g2_buf_1  output16
timestamp 1676381911
transform 1 0 18240 0 -1 7560
box -48 -56 432 834
use sg13g2_buf_1  output17
timestamp 1676381911
transform 1 0 18720 0 1 6048
box -48 -56 432 834
use sg13g2_buf_1  output18
timestamp 1676381911
transform 1 0 16992 0 1 7560
box -48 -56 432 834
use sg13g2_buf_1  output19
timestamp 1676381911
transform 1 0 18336 0 1 6048
box -48 -56 432 834
use sg13g2_buf_1  output20
timestamp 1676381911
transform 1 0 17472 0 -1 7560
box -48 -56 432 834
use sg13g2_buf_1  output21
timestamp 1676381911
transform 1 0 16608 0 1 7560
box -48 -56 432 834
use sg13g2_buf_1  output22
timestamp 1676381911
transform 1 0 15744 0 -1 9072
box -48 -56 432 834
use sg13g2_buf_1  output23
timestamp 1676381911
transform 1 0 18528 0 -1 3024
box -48 -56 432 834
use sg13g2_buf_1  output24
timestamp 1676381911
transform 1 0 14976 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  output25
timestamp 1676381911
transform 1 0 16224 0 1 7560
box -48 -56 432 834
use sg13g2_buf_1  output26
timestamp 1676381911
transform 1 0 19296 0 1 1512
box -48 -56 432 834
use sg13g2_buf_1  output27
timestamp 1676381911
transform 1 0 18912 0 -1 3024
box -48 -56 432 834
use sg13g2_buf_1  output28
timestamp 1676381911
transform 1 0 19680 0 1 1512
box -48 -56 432 834
use sg13g2_buf_1  output29
timestamp 1676381911
transform 1 0 20064 0 1 1512
box -48 -56 432 834
use sg13g2_buf_1  output30
timestamp 1676381911
transform 1 0 19680 0 -1 3024
box -48 -56 432 834
use sg13g2_buf_1  output31
timestamp 1676381911
transform 1 0 19296 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  output32
timestamp 1676381911
transform 1 0 20064 0 -1 3024
box -48 -56 432 834
use sg13g2_buf_1  output33
timestamp 1676381911
transform -1 0 16896 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  output34
timestamp 1676381911
transform -1 0 18816 0 -1 9072
box -48 -56 432 834
use sg13g2_buf_1  output35
timestamp 1676381911
transform -1 0 19584 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  output36
timestamp 1676381911
transform -1 0 19200 0 -1 9072
box -48 -56 432 834
use sg13g2_buf_1  output37
timestamp 1676381911
transform -1 0 19968 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  output38
timestamp 1676381911
transform -1 0 18912 0 1 7560
box -48 -56 432 834
use sg13g2_buf_1  output39
timestamp 1676381911
transform -1 0 19296 0 1 7560
box -48 -56 432 834
use sg13g2_buf_1  output40
timestamp 1676381911
transform -1 0 20352 0 -1 9072
box -48 -56 432 834
use sg13g2_buf_1  output41
timestamp 1676381911
transform 1 0 18624 0 -1 7560
box -48 -56 432 834
use sg13g2_buf_1  output42
timestamp 1676381911
transform 1 0 17760 0 1 7560
box -48 -56 432 834
use sg13g2_buf_1  output43
timestamp 1676381911
transform 1 0 17376 0 1 7560
box -48 -56 432 834
use sg13g2_buf_1  output44
timestamp 1676381911
transform -1 0 17280 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  output45
timestamp 1676381911
transform 1 0 15360 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  output46
timestamp 1676381911
transform -1 0 17664 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  output47
timestamp 1676381911
transform -1 0 17280 0 -1 9072
box -48 -56 432 834
use sg13g2_buf_1  output48
timestamp 1676381911
transform -1 0 18048 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  output49
timestamp 1676381911
transform -1 0 17664 0 -1 9072
box -48 -56 432 834
use sg13g2_buf_1  output50
timestamp 1676381911
transform -1 0 18432 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  output51
timestamp 1676381911
transform -1 0 18816 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  output52
timestamp 1676381911
transform -1 0 19200 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  output53
timestamp 1676381911
transform 1 0 1152 0 -1 9072
box -48 -56 432 834
use sg13g2_buf_1  output54
timestamp 1676381911
transform -1 0 2400 0 1 7560
box -48 -56 432 834
use sg13g2_buf_1  output55
timestamp 1676381911
transform 1 0 1536 0 -1 9072
box -48 -56 432 834
use sg13g2_buf_1  output56
timestamp 1676381911
transform 1 0 1248 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  output57
timestamp 1676381911
transform 1 0 1632 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  output58
timestamp 1676381911
transform 1 0 2016 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  output59
timestamp 1676381911
transform 1 0 2400 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  output60
timestamp 1676381911
transform -1 0 3552 0 -1 9072
box -48 -56 432 834
use sg13g2_buf_1  output61
timestamp 1676381911
transform 1 0 2784 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  output62
timestamp 1676381911
transform -1 0 3936 0 -1 9072
box -48 -56 432 834
use sg13g2_buf_1  output63
timestamp 1676381911
transform 1 0 3168 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  output64
timestamp 1676381911
transform -1 0 4320 0 -1 9072
box -48 -56 432 834
use sg13g2_buf_1  output65
timestamp 1676381911
transform 1 0 3552 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  output66
timestamp 1676381911
transform -1 0 4704 0 -1 9072
box -48 -56 432 834
use sg13g2_buf_1  output67
timestamp 1676381911
transform 1 0 3936 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  output68
timestamp 1676381911
transform -1 0 5088 0 -1 9072
box -48 -56 432 834
use sg13g2_buf_1  output69
timestamp 1676381911
transform 1 0 4320 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  output70
timestamp 1676381911
transform -1 0 5472 0 -1 9072
box -48 -56 432 834
use sg13g2_buf_1  output71
timestamp 1676381911
transform 1 0 4704 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  output72
timestamp 1676381911
transform -1 0 5856 0 -1 9072
box -48 -56 432 834
use sg13g2_buf_1  output73
timestamp 1676381911
transform 1 0 5088 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  output74
timestamp 1676381911
transform 1 0 7008 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  output75
timestamp 1676381911
transform 1 0 7392 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  output76
timestamp 1676381911
transform -1 0 8160 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  output77
timestamp 1676381911
transform -1 0 8544 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  output78
timestamp 1676381911
transform -1 0 9312 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  output79
timestamp 1676381911
transform -1 0 8928 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  output80
timestamp 1676381911
transform -1 0 6240 0 -1 9072
box -48 -56 432 834
use sg13g2_buf_1  output81
timestamp 1676381911
transform 1 0 5472 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  output82
timestamp 1676381911
transform -1 0 6624 0 -1 9072
box -48 -56 432 834
use sg13g2_buf_1  output83
timestamp 1676381911
transform 1 0 5856 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  output84
timestamp 1676381911
transform -1 0 7008 0 -1 9072
box -48 -56 432 834
use sg13g2_buf_1  output85
timestamp 1676381911
transform 1 0 6240 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  output86
timestamp 1676381911
transform -1 0 7392 0 -1 9072
box -48 -56 432 834
use sg13g2_buf_1  output87
timestamp 1676381911
transform 1 0 6624 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  output88
timestamp 1676381911
transform -1 0 7776 0 -1 9072
box -48 -56 432 834
use sg13g2_buf_1  output89
timestamp 1676381911
transform -1 0 16512 0 1 9072
box -48 -56 432 834
<< labels >>
flabel metal2 s 0 548 90 628 0 FreeSans 320 0 0 0 FrameData[0]
port 0 nsew signal input
flabel metal2 s 0 3908 90 3988 0 FreeSans 320 0 0 0 FrameData[10]
port 1 nsew signal input
flabel metal2 s 0 4244 90 4324 0 FreeSans 320 0 0 0 FrameData[11]
port 2 nsew signal input
flabel metal2 s 0 4580 90 4660 0 FreeSans 320 0 0 0 FrameData[12]
port 3 nsew signal input
flabel metal2 s 0 4916 90 4996 0 FreeSans 320 0 0 0 FrameData[13]
port 4 nsew signal input
flabel metal2 s 0 5252 90 5332 0 FreeSans 320 0 0 0 FrameData[14]
port 5 nsew signal input
flabel metal2 s 0 5588 90 5668 0 FreeSans 320 0 0 0 FrameData[15]
port 6 nsew signal input
flabel metal2 s 0 5924 90 6004 0 FreeSans 320 0 0 0 FrameData[16]
port 7 nsew signal input
flabel metal2 s 0 6260 90 6340 0 FreeSans 320 0 0 0 FrameData[17]
port 8 nsew signal input
flabel metal2 s 0 6596 90 6676 0 FreeSans 320 0 0 0 FrameData[18]
port 9 nsew signal input
flabel metal2 s 0 6932 90 7012 0 FreeSans 320 0 0 0 FrameData[19]
port 10 nsew signal input
flabel metal2 s 0 884 90 964 0 FreeSans 320 0 0 0 FrameData[1]
port 11 nsew signal input
flabel metal2 s 0 7268 90 7348 0 FreeSans 320 0 0 0 FrameData[20]
port 12 nsew signal input
flabel metal2 s 0 7604 90 7684 0 FreeSans 320 0 0 0 FrameData[21]
port 13 nsew signal input
flabel metal2 s 0 7940 90 8020 0 FreeSans 320 0 0 0 FrameData[22]
port 14 nsew signal input
flabel metal2 s 0 8276 90 8356 0 FreeSans 320 0 0 0 FrameData[23]
port 15 nsew signal input
flabel metal2 s 0 8612 90 8692 0 FreeSans 320 0 0 0 FrameData[24]
port 16 nsew signal input
flabel metal2 s 0 8948 90 9028 0 FreeSans 320 0 0 0 FrameData[25]
port 17 nsew signal input
flabel metal2 s 0 9284 90 9364 0 FreeSans 320 0 0 0 FrameData[26]
port 18 nsew signal input
flabel metal2 s 0 9620 90 9700 0 FreeSans 320 0 0 0 FrameData[27]
port 19 nsew signal input
flabel metal2 s 0 9956 90 10036 0 FreeSans 320 0 0 0 FrameData[28]
port 20 nsew signal input
flabel metal2 s 0 10292 90 10372 0 FreeSans 320 0 0 0 FrameData[29]
port 21 nsew signal input
flabel metal2 s 0 1220 90 1300 0 FreeSans 320 0 0 0 FrameData[2]
port 22 nsew signal input
flabel metal2 s 0 10628 90 10708 0 FreeSans 320 0 0 0 FrameData[30]
port 23 nsew signal input
flabel metal2 s 0 10964 90 11044 0 FreeSans 320 0 0 0 FrameData[31]
port 24 nsew signal input
flabel metal2 s 0 1556 90 1636 0 FreeSans 320 0 0 0 FrameData[3]
port 25 nsew signal input
flabel metal2 s 0 1892 90 1972 0 FreeSans 320 0 0 0 FrameData[4]
port 26 nsew signal input
flabel metal2 s 0 2228 90 2308 0 FreeSans 320 0 0 0 FrameData[5]
port 27 nsew signal input
flabel metal2 s 0 2564 90 2644 0 FreeSans 320 0 0 0 FrameData[6]
port 28 nsew signal input
flabel metal2 s 0 2900 90 2980 0 FreeSans 320 0 0 0 FrameData[7]
port 29 nsew signal input
flabel metal2 s 0 3236 90 3316 0 FreeSans 320 0 0 0 FrameData[8]
port 30 nsew signal input
flabel metal2 s 0 3572 90 3652 0 FreeSans 320 0 0 0 FrameData[9]
port 31 nsew signal input
flabel metal2 s 21510 548 21600 628 0 FreeSans 320 0 0 0 FrameData_O[0]
port 32 nsew signal output
flabel metal2 s 21510 3908 21600 3988 0 FreeSans 320 0 0 0 FrameData_O[10]
port 33 nsew signal output
flabel metal2 s 21510 4244 21600 4324 0 FreeSans 320 0 0 0 FrameData_O[11]
port 34 nsew signal output
flabel metal2 s 21510 4580 21600 4660 0 FreeSans 320 0 0 0 FrameData_O[12]
port 35 nsew signal output
flabel metal2 s 21510 4916 21600 4996 0 FreeSans 320 0 0 0 FrameData_O[13]
port 36 nsew signal output
flabel metal2 s 21510 5252 21600 5332 0 FreeSans 320 0 0 0 FrameData_O[14]
port 37 nsew signal output
flabel metal2 s 21510 5588 21600 5668 0 FreeSans 320 0 0 0 FrameData_O[15]
port 38 nsew signal output
flabel metal2 s 21510 5924 21600 6004 0 FreeSans 320 0 0 0 FrameData_O[16]
port 39 nsew signal output
flabel metal2 s 21510 6260 21600 6340 0 FreeSans 320 0 0 0 FrameData_O[17]
port 40 nsew signal output
flabel metal2 s 21510 6596 21600 6676 0 FreeSans 320 0 0 0 FrameData_O[18]
port 41 nsew signal output
flabel metal2 s 21510 6932 21600 7012 0 FreeSans 320 0 0 0 FrameData_O[19]
port 42 nsew signal output
flabel metal2 s 21510 884 21600 964 0 FreeSans 320 0 0 0 FrameData_O[1]
port 43 nsew signal output
flabel metal2 s 21510 7268 21600 7348 0 FreeSans 320 0 0 0 FrameData_O[20]
port 44 nsew signal output
flabel metal2 s 21510 7604 21600 7684 0 FreeSans 320 0 0 0 FrameData_O[21]
port 45 nsew signal output
flabel metal2 s 21510 7940 21600 8020 0 FreeSans 320 0 0 0 FrameData_O[22]
port 46 nsew signal output
flabel metal2 s 21510 8276 21600 8356 0 FreeSans 320 0 0 0 FrameData_O[23]
port 47 nsew signal output
flabel metal2 s 21510 8612 21600 8692 0 FreeSans 320 0 0 0 FrameData_O[24]
port 48 nsew signal output
flabel metal2 s 21510 8948 21600 9028 0 FreeSans 320 0 0 0 FrameData_O[25]
port 49 nsew signal output
flabel metal2 s 21510 9284 21600 9364 0 FreeSans 320 0 0 0 FrameData_O[26]
port 50 nsew signal output
flabel metal2 s 21510 9620 21600 9700 0 FreeSans 320 0 0 0 FrameData_O[27]
port 51 nsew signal output
flabel metal2 s 21510 9956 21600 10036 0 FreeSans 320 0 0 0 FrameData_O[28]
port 52 nsew signal output
flabel metal2 s 21510 10292 21600 10372 0 FreeSans 320 0 0 0 FrameData_O[29]
port 53 nsew signal output
flabel metal2 s 21510 1220 21600 1300 0 FreeSans 320 0 0 0 FrameData_O[2]
port 54 nsew signal output
flabel metal2 s 21510 10628 21600 10708 0 FreeSans 320 0 0 0 FrameData_O[30]
port 55 nsew signal output
flabel metal2 s 21510 10964 21600 11044 0 FreeSans 320 0 0 0 FrameData_O[31]
port 56 nsew signal output
flabel metal2 s 21510 1556 21600 1636 0 FreeSans 320 0 0 0 FrameData_O[3]
port 57 nsew signal output
flabel metal2 s 21510 1892 21600 1972 0 FreeSans 320 0 0 0 FrameData_O[4]
port 58 nsew signal output
flabel metal2 s 21510 2228 21600 2308 0 FreeSans 320 0 0 0 FrameData_O[5]
port 59 nsew signal output
flabel metal2 s 21510 2564 21600 2644 0 FreeSans 320 0 0 0 FrameData_O[6]
port 60 nsew signal output
flabel metal2 s 21510 2900 21600 2980 0 FreeSans 320 0 0 0 FrameData_O[7]
port 61 nsew signal output
flabel metal2 s 21510 3236 21600 3316 0 FreeSans 320 0 0 0 FrameData_O[8]
port 62 nsew signal output
flabel metal2 s 21510 3572 21600 3652 0 FreeSans 320 0 0 0 FrameData_O[9]
port 63 nsew signal output
flabel metal3 s 1976 0 2056 80 0 FreeSans 320 0 0 0 FrameStrobe[0]
port 64 nsew signal input
flabel metal3 s 11576 0 11656 80 0 FreeSans 320 0 0 0 FrameStrobe[10]
port 65 nsew signal input
flabel metal3 s 12536 0 12616 80 0 FreeSans 320 0 0 0 FrameStrobe[11]
port 66 nsew signal input
flabel metal3 s 13496 0 13576 80 0 FreeSans 320 0 0 0 FrameStrobe[12]
port 67 nsew signal input
flabel metal3 s 14456 0 14536 80 0 FreeSans 320 0 0 0 FrameStrobe[13]
port 68 nsew signal input
flabel metal3 s 15416 0 15496 80 0 FreeSans 320 0 0 0 FrameStrobe[14]
port 69 nsew signal input
flabel metal3 s 16376 0 16456 80 0 FreeSans 320 0 0 0 FrameStrobe[15]
port 70 nsew signal input
flabel metal3 s 17336 0 17416 80 0 FreeSans 320 0 0 0 FrameStrobe[16]
port 71 nsew signal input
flabel metal3 s 18296 0 18376 80 0 FreeSans 320 0 0 0 FrameStrobe[17]
port 72 nsew signal input
flabel metal3 s 19256 0 19336 80 0 FreeSans 320 0 0 0 FrameStrobe[18]
port 73 nsew signal input
flabel metal3 s 20216 0 20296 80 0 FreeSans 320 0 0 0 FrameStrobe[19]
port 74 nsew signal input
flabel metal3 s 2936 0 3016 80 0 FreeSans 320 0 0 0 FrameStrobe[1]
port 75 nsew signal input
flabel metal3 s 3896 0 3976 80 0 FreeSans 320 0 0 0 FrameStrobe[2]
port 76 nsew signal input
flabel metal3 s 4856 0 4936 80 0 FreeSans 320 0 0 0 FrameStrobe[3]
port 77 nsew signal input
flabel metal3 s 5816 0 5896 80 0 FreeSans 320 0 0 0 FrameStrobe[4]
port 78 nsew signal input
flabel metal3 s 6776 0 6856 80 0 FreeSans 320 0 0 0 FrameStrobe[5]
port 79 nsew signal input
flabel metal3 s 7736 0 7816 80 0 FreeSans 320 0 0 0 FrameStrobe[6]
port 80 nsew signal input
flabel metal3 s 8696 0 8776 80 0 FreeSans 320 0 0 0 FrameStrobe[7]
port 81 nsew signal input
flabel metal3 s 9656 0 9736 80 0 FreeSans 320 0 0 0 FrameStrobe[8]
port 82 nsew signal input
flabel metal3 s 10616 0 10696 80 0 FreeSans 320 0 0 0 FrameStrobe[9]
port 83 nsew signal input
flabel metal3 s 15800 11764 15880 11844 0 FreeSans 320 0 0 0 FrameStrobe_O[0]
port 84 nsew signal output
flabel metal3 s 17720 11764 17800 11844 0 FreeSans 320 0 0 0 FrameStrobe_O[10]
port 85 nsew signal output
flabel metal3 s 17912 11764 17992 11844 0 FreeSans 320 0 0 0 FrameStrobe_O[11]
port 86 nsew signal output
flabel metal3 s 18104 11764 18184 11844 0 FreeSans 320 0 0 0 FrameStrobe_O[12]
port 87 nsew signal output
flabel metal3 s 18296 11764 18376 11844 0 FreeSans 320 0 0 0 FrameStrobe_O[13]
port 88 nsew signal output
flabel metal3 s 18488 11764 18568 11844 0 FreeSans 320 0 0 0 FrameStrobe_O[14]
port 89 nsew signal output
flabel metal3 s 18680 11764 18760 11844 0 FreeSans 320 0 0 0 FrameStrobe_O[15]
port 90 nsew signal output
flabel metal3 s 18872 11764 18952 11844 0 FreeSans 320 0 0 0 FrameStrobe_O[16]
port 91 nsew signal output
flabel metal3 s 19064 11764 19144 11844 0 FreeSans 320 0 0 0 FrameStrobe_O[17]
port 92 nsew signal output
flabel metal3 s 19256 11764 19336 11844 0 FreeSans 320 0 0 0 FrameStrobe_O[18]
port 93 nsew signal output
flabel metal3 s 19448 11764 19528 11844 0 FreeSans 320 0 0 0 FrameStrobe_O[19]
port 94 nsew signal output
flabel metal3 s 15992 11764 16072 11844 0 FreeSans 320 0 0 0 FrameStrobe_O[1]
port 95 nsew signal output
flabel metal3 s 16184 11764 16264 11844 0 FreeSans 320 0 0 0 FrameStrobe_O[2]
port 96 nsew signal output
flabel metal3 s 16376 11764 16456 11844 0 FreeSans 320 0 0 0 FrameStrobe_O[3]
port 97 nsew signal output
flabel metal3 s 16568 11764 16648 11844 0 FreeSans 320 0 0 0 FrameStrobe_O[4]
port 98 nsew signal output
flabel metal3 s 16760 11764 16840 11844 0 FreeSans 320 0 0 0 FrameStrobe_O[5]
port 99 nsew signal output
flabel metal3 s 16952 11764 17032 11844 0 FreeSans 320 0 0 0 FrameStrobe_O[6]
port 100 nsew signal output
flabel metal3 s 17144 11764 17224 11844 0 FreeSans 320 0 0 0 FrameStrobe_O[7]
port 101 nsew signal output
flabel metal3 s 17336 11764 17416 11844 0 FreeSans 320 0 0 0 FrameStrobe_O[8]
port 102 nsew signal output
flabel metal3 s 17528 11764 17608 11844 0 FreeSans 320 0 0 0 FrameStrobe_O[9]
port 103 nsew signal output
flabel metal3 s 1784 11764 1864 11844 0 FreeSans 320 0 0 0 N1BEG[0]
port 104 nsew signal output
flabel metal3 s 1976 11764 2056 11844 0 FreeSans 320 0 0 0 N1BEG[1]
port 105 nsew signal output
flabel metal3 s 2168 11764 2248 11844 0 FreeSans 320 0 0 0 N1BEG[2]
port 106 nsew signal output
flabel metal3 s 2360 11764 2440 11844 0 FreeSans 320 0 0 0 N1BEG[3]
port 107 nsew signal output
flabel metal3 s 2552 11764 2632 11844 0 FreeSans 320 0 0 0 N2BEG[0]
port 108 nsew signal output
flabel metal3 s 2744 11764 2824 11844 0 FreeSans 320 0 0 0 N2BEG[1]
port 109 nsew signal output
flabel metal3 s 2936 11764 3016 11844 0 FreeSans 320 0 0 0 N2BEG[2]
port 110 nsew signal output
flabel metal3 s 3128 11764 3208 11844 0 FreeSans 320 0 0 0 N2BEG[3]
port 111 nsew signal output
flabel metal3 s 3320 11764 3400 11844 0 FreeSans 320 0 0 0 N2BEG[4]
port 112 nsew signal output
flabel metal3 s 3512 11764 3592 11844 0 FreeSans 320 0 0 0 N2BEG[5]
port 113 nsew signal output
flabel metal3 s 3704 11764 3784 11844 0 FreeSans 320 0 0 0 N2BEG[6]
port 114 nsew signal output
flabel metal3 s 3896 11764 3976 11844 0 FreeSans 320 0 0 0 N2BEG[7]
port 115 nsew signal output
flabel metal3 s 4088 11764 4168 11844 0 FreeSans 320 0 0 0 N2BEGb[0]
port 116 nsew signal output
flabel metal3 s 4280 11764 4360 11844 0 FreeSans 320 0 0 0 N2BEGb[1]
port 117 nsew signal output
flabel metal3 s 4472 11764 4552 11844 0 FreeSans 320 0 0 0 N2BEGb[2]
port 118 nsew signal output
flabel metal3 s 4664 11764 4744 11844 0 FreeSans 320 0 0 0 N2BEGb[3]
port 119 nsew signal output
flabel metal3 s 4856 11764 4936 11844 0 FreeSans 320 0 0 0 N2BEGb[4]
port 120 nsew signal output
flabel metal3 s 5048 11764 5128 11844 0 FreeSans 320 0 0 0 N2BEGb[5]
port 121 nsew signal output
flabel metal3 s 5240 11764 5320 11844 0 FreeSans 320 0 0 0 N2BEGb[6]
port 122 nsew signal output
flabel metal3 s 5432 11764 5512 11844 0 FreeSans 320 0 0 0 N2BEGb[7]
port 123 nsew signal output
flabel metal3 s 5624 11764 5704 11844 0 FreeSans 320 0 0 0 N4BEG[0]
port 124 nsew signal output
flabel metal3 s 7544 11764 7624 11844 0 FreeSans 320 0 0 0 N4BEG[10]
port 125 nsew signal output
flabel metal3 s 7736 11764 7816 11844 0 FreeSans 320 0 0 0 N4BEG[11]
port 126 nsew signal output
flabel metal3 s 7928 11764 8008 11844 0 FreeSans 320 0 0 0 N4BEG[12]
port 127 nsew signal output
flabel metal3 s 8120 11764 8200 11844 0 FreeSans 320 0 0 0 N4BEG[13]
port 128 nsew signal output
flabel metal3 s 8312 11764 8392 11844 0 FreeSans 320 0 0 0 N4BEG[14]
port 129 nsew signal output
flabel metal3 s 8504 11764 8584 11844 0 FreeSans 320 0 0 0 N4BEG[15]
port 130 nsew signal output
flabel metal3 s 5816 11764 5896 11844 0 FreeSans 320 0 0 0 N4BEG[1]
port 131 nsew signal output
flabel metal3 s 6008 11764 6088 11844 0 FreeSans 320 0 0 0 N4BEG[2]
port 132 nsew signal output
flabel metal3 s 6200 11764 6280 11844 0 FreeSans 320 0 0 0 N4BEG[3]
port 133 nsew signal output
flabel metal3 s 6392 11764 6472 11844 0 FreeSans 320 0 0 0 N4BEG[4]
port 134 nsew signal output
flabel metal3 s 6584 11764 6664 11844 0 FreeSans 320 0 0 0 N4BEG[5]
port 135 nsew signal output
flabel metal3 s 6776 11764 6856 11844 0 FreeSans 320 0 0 0 N4BEG[6]
port 136 nsew signal output
flabel metal3 s 6968 11764 7048 11844 0 FreeSans 320 0 0 0 N4BEG[7]
port 137 nsew signal output
flabel metal3 s 7160 11764 7240 11844 0 FreeSans 320 0 0 0 N4BEG[8]
port 138 nsew signal output
flabel metal3 s 7352 11764 7432 11844 0 FreeSans 320 0 0 0 N4BEG[9]
port 139 nsew signal output
flabel metal3 s 8696 11764 8776 11844 0 FreeSans 320 0 0 0 S1END[0]
port 140 nsew signal input
flabel metal3 s 8888 11764 8968 11844 0 FreeSans 320 0 0 0 S1END[1]
port 141 nsew signal input
flabel metal3 s 9080 11764 9160 11844 0 FreeSans 320 0 0 0 S1END[2]
port 142 nsew signal input
flabel metal3 s 9272 11764 9352 11844 0 FreeSans 320 0 0 0 S1END[3]
port 143 nsew signal input
flabel metal3 s 11000 11764 11080 11844 0 FreeSans 320 0 0 0 S2END[0]
port 144 nsew signal input
flabel metal3 s 11192 11764 11272 11844 0 FreeSans 320 0 0 0 S2END[1]
port 145 nsew signal input
flabel metal3 s 11384 11764 11464 11844 0 FreeSans 320 0 0 0 S2END[2]
port 146 nsew signal input
flabel metal3 s 11576 11764 11656 11844 0 FreeSans 320 0 0 0 S2END[3]
port 147 nsew signal input
flabel metal3 s 11768 11764 11848 11844 0 FreeSans 320 0 0 0 S2END[4]
port 148 nsew signal input
flabel metal3 s 11960 11764 12040 11844 0 FreeSans 320 0 0 0 S2END[5]
port 149 nsew signal input
flabel metal3 s 12152 11764 12232 11844 0 FreeSans 320 0 0 0 S2END[6]
port 150 nsew signal input
flabel metal3 s 12344 11764 12424 11844 0 FreeSans 320 0 0 0 S2END[7]
port 151 nsew signal input
flabel metal3 s 9464 11764 9544 11844 0 FreeSans 320 0 0 0 S2MID[0]
port 152 nsew signal input
flabel metal3 s 9656 11764 9736 11844 0 FreeSans 320 0 0 0 S2MID[1]
port 153 nsew signal input
flabel metal3 s 9848 11764 9928 11844 0 FreeSans 320 0 0 0 S2MID[2]
port 154 nsew signal input
flabel metal3 s 10040 11764 10120 11844 0 FreeSans 320 0 0 0 S2MID[3]
port 155 nsew signal input
flabel metal3 s 10232 11764 10312 11844 0 FreeSans 320 0 0 0 S2MID[4]
port 156 nsew signal input
flabel metal3 s 10424 11764 10504 11844 0 FreeSans 320 0 0 0 S2MID[5]
port 157 nsew signal input
flabel metal3 s 10616 11764 10696 11844 0 FreeSans 320 0 0 0 S2MID[6]
port 158 nsew signal input
flabel metal3 s 10808 11764 10888 11844 0 FreeSans 320 0 0 0 S2MID[7]
port 159 nsew signal input
flabel metal3 s 12536 11764 12616 11844 0 FreeSans 320 0 0 0 S4END[0]
port 160 nsew signal input
flabel metal3 s 14456 11764 14536 11844 0 FreeSans 320 0 0 0 S4END[10]
port 161 nsew signal input
flabel metal3 s 14648 11764 14728 11844 0 FreeSans 320 0 0 0 S4END[11]
port 162 nsew signal input
flabel metal3 s 14840 11764 14920 11844 0 FreeSans 320 0 0 0 S4END[12]
port 163 nsew signal input
flabel metal3 s 15032 11764 15112 11844 0 FreeSans 320 0 0 0 S4END[13]
port 164 nsew signal input
flabel metal3 s 15224 11764 15304 11844 0 FreeSans 320 0 0 0 S4END[14]
port 165 nsew signal input
flabel metal3 s 15416 11764 15496 11844 0 FreeSans 320 0 0 0 S4END[15]
port 166 nsew signal input
flabel metal3 s 12728 11764 12808 11844 0 FreeSans 320 0 0 0 S4END[1]
port 167 nsew signal input
flabel metal3 s 12920 11764 13000 11844 0 FreeSans 320 0 0 0 S4END[2]
port 168 nsew signal input
flabel metal3 s 13112 11764 13192 11844 0 FreeSans 320 0 0 0 S4END[3]
port 169 nsew signal input
flabel metal3 s 13304 11764 13384 11844 0 FreeSans 320 0 0 0 S4END[4]
port 170 nsew signal input
flabel metal3 s 13496 11764 13576 11844 0 FreeSans 320 0 0 0 S4END[5]
port 171 nsew signal input
flabel metal3 s 13688 11764 13768 11844 0 FreeSans 320 0 0 0 S4END[6]
port 172 nsew signal input
flabel metal3 s 13880 11764 13960 11844 0 FreeSans 320 0 0 0 S4END[7]
port 173 nsew signal input
flabel metal3 s 14072 11764 14152 11844 0 FreeSans 320 0 0 0 S4END[8]
port 174 nsew signal input
flabel metal3 s 14264 11764 14344 11844 0 FreeSans 320 0 0 0 S4END[9]
port 175 nsew signal input
flabel metal3 s 1016 0 1096 80 0 FreeSans 320 0 0 0 UserCLK
port 176 nsew signal input
flabel metal3 s 15608 11764 15688 11844 0 FreeSans 320 0 0 0 UserCLKo
port 177 nsew signal output
flabel metal5 s 4892 0 5332 11844 0 FreeSans 2560 90 0 0 VGND
port 178 nsew ground bidirectional
flabel metal5 s 4892 0 5332 40 0 FreeSans 320 0 0 0 VGND
port 178 nsew ground bidirectional
flabel metal5 s 4892 11804 5332 11844 0 FreeSans 320 0 0 0 VGND
port 178 nsew ground bidirectional
flabel metal5 s 20012 0 20452 11844 0 FreeSans 2560 90 0 0 VGND
port 178 nsew ground bidirectional
flabel metal5 s 20012 0 20452 40 0 FreeSans 320 0 0 0 VGND
port 178 nsew ground bidirectional
flabel metal5 s 20012 11804 20452 11844 0 FreeSans 320 0 0 0 VGND
port 178 nsew ground bidirectional
flabel metal5 s 3652 0 4092 11844 0 FreeSans 2560 90 0 0 VPWR
port 179 nsew power bidirectional
flabel metal5 s 3652 0 4092 40 0 FreeSans 320 0 0 0 VPWR
port 179 nsew power bidirectional
flabel metal5 s 3652 11804 4092 11844 0 FreeSans 320 0 0 0 VPWR
port 179 nsew power bidirectional
flabel metal5 s 18772 0 19212 11844 0 FreeSans 2560 90 0 0 VPWR
port 179 nsew power bidirectional
flabel metal5 s 18772 0 19212 40 0 FreeSans 320 0 0 0 VPWR
port 179 nsew power bidirectional
flabel metal5 s 18772 11804 19212 11844 0 FreeSans 320 0 0 0 VPWR
port 179 nsew power bidirectional
rlabel metal1 10802 9072 10802 9072 0 VGND
rlabel metal1 10800 9828 10800 9828 0 VPWR
rlabel metal2 4304 588 4304 588 0 FrameData[0]
rlabel metal2 1472 3948 1472 3948 0 FrameData[10]
rlabel metal2 5072 4284 5072 4284 0 FrameData[11]
rlabel metal2 19296 4914 19296 4914 0 FrameData[12]
rlabel metal2 128 4956 128 4956 0 FrameData[13]
rlabel metal2 1832 5292 1832 5292 0 FrameData[14]
rlabel metal2 800 5628 800 5628 0 FrameData[15]
rlabel metal2 128 5964 128 5964 0 FrameData[16]
rlabel metal2 752 6300 752 6300 0 FrameData[17]
rlabel metal3 14592 7770 14592 7770 0 FrameData[18]
rlabel metal2 752 6972 752 6972 0 FrameData[19]
rlabel metal2 752 924 752 924 0 FrameData[1]
rlabel metal2 320 7308 320 7308 0 FrameData[20]
rlabel metal2 704 7644 704 7644 0 FrameData[21]
rlabel metal2 176 7980 176 7980 0 FrameData[22]
rlabel metal2 608 8316 608 8316 0 FrameData[23]
rlabel metal2 512 8652 512 8652 0 FrameData[24]
rlabel metal3 16224 8694 16224 8694 0 FrameData[25]
rlabel metal2 11904 9408 11904 9408 0 FrameData[26]
rlabel metal2 128 9660 128 9660 0 FrameData[27]
rlabel metal2 1376 9996 1376 9996 0 FrameData[28]
rlabel metal2 176 10332 176 10332 0 FrameData[29]
rlabel metal2 704 1260 704 1260 0 FrameData[2]
rlabel metal2 368 10668 368 10668 0 FrameData[30]
rlabel metal2 224 11004 224 11004 0 FrameData[31]
rlabel metal2 656 1596 656 1596 0 FrameData[3]
rlabel metal2 5024 1932 5024 1932 0 FrameData[4]
rlabel metal2 1808 2268 1808 2268 0 FrameData[5]
rlabel metal2 1088 2604 1088 2604 0 FrameData[6]
rlabel metal2 8592 2856 8592 2856 0 FrameData[7]
rlabel metal2 17280 2016 17280 2016 0 FrameData[8]
rlabel metal2 128 3612 128 3612 0 FrameData[9]
rlabel metal2 21279 588 21279 588 0 FrameData_O[0]
rlabel metal2 20040 3192 20040 3192 0 FrameData_O[10]
rlabel metal2 20568 3612 20568 3612 0 FrameData_O[11]
rlabel metal2 20703 4620 20703 4620 0 FrameData_O[12]
rlabel metal2 20472 4284 20472 4284 0 FrameData_O[13]
rlabel metal2 20016 5208 20016 5208 0 FrameData_O[14]
rlabel metal2 20568 5040 20568 5040 0 FrameData_O[15]
rlabel metal2 20016 5922 20016 5922 0 FrameData_O[16]
rlabel metal2 20472 5628 20472 5628 0 FrameData_O[17]
rlabel metal2 20967 6636 20967 6636 0 FrameData_O[18]
rlabel metal2 20967 6972 20967 6972 0 FrameData_O[19]
rlabel metal2 21039 924 21039 924 0 FrameData_O[1]
rlabel metal2 21279 7308 21279 7308 0 FrameData_O[20]
rlabel metal2 20775 7644 20775 7644 0 FrameData_O[21]
rlabel metal2 21087 7980 21087 7980 0 FrameData_O[22]
rlabel metal2 18984 7392 18984 7392 0 FrameData_O[23]
rlabel metal2 19176 6636 19176 6636 0 FrameData_O[24]
rlabel metal2 17640 8148 17640 8148 0 FrameData_O[25]
rlabel metal2 18648 6636 18648 6636 0 FrameData_O[26]
rlabel metal2 17784 7140 17784 7140 0 FrameData_O[27]
rlabel metal2 17064 8148 17064 8148 0 FrameData_O[28]
rlabel metal2 16104 8904 16104 8904 0 FrameData_O[29]
rlabel metal2 21087 1260 21087 1260 0 FrameData_O[2]
rlabel metal2 16200 9324 16200 9324 0 FrameData_O[30]
rlabel metal2 17064 7728 17064 7728 0 FrameData_O[31]
rlabel metal2 20583 1596 20583 1596 0 FrameData_O[3]
rlabel metal2 20991 1932 20991 1932 0 FrameData_O[4]
rlabel metal2 20016 2184 20016 2184 0 FrameData_O[5]
rlabel metal2 20712 2016 20712 2016 0 FrameData_O[6]
rlabel metal2 20088 2856 20088 2856 0 FrameData_O[7]
rlabel metal2 20583 3276 20583 3276 0 FrameData_O[8]
rlabel metal2 20760 2856 20760 2856 0 FrameData_O[9]
rlabel metal2 1968 3444 1968 3444 0 FrameStrobe[0]
rlabel metal2 13200 3444 13200 3444 0 FrameStrobe[10]
rlabel metal2 11808 5544 11808 5544 0 FrameStrobe[11]
rlabel metal3 13488 4200 13488 4200 0 FrameStrobe[12]
rlabel metal3 14496 2844 14496 2844 0 FrameStrobe[13]
rlabel metal2 14400 8736 14400 8736 0 FrameStrobe[14]
rlabel metal2 15120 3360 15120 3360 0 FrameStrobe[15]
rlabel metal2 12960 1848 12960 1848 0 FrameStrobe[16]
rlabel metal3 18336 1206 18336 1206 0 FrameStrobe[17]
rlabel via3 19296 72 19296 72 0 FrameStrobe[18]
rlabel metal3 20256 114 20256 114 0 FrameStrobe[19]
rlabel metal2 3168 6468 3168 6468 0 FrameStrobe[1]
rlabel metal3 3936 114 3936 114 0 FrameStrobe[2]
rlabel metal3 4896 492 4896 492 0 FrameStrobe[3]
rlabel metal2 5520 4956 5520 4956 0 FrameStrobe[4]
rlabel metal2 6576 3444 6576 3444 0 FrameStrobe[5]
rlabel metal3 7776 1332 7776 1332 0 FrameStrobe[6]
rlabel metal2 8832 3444 8832 3444 0 FrameStrobe[7]
rlabel metal2 10224 3360 10224 3360 0 FrameStrobe[8]
rlabel metal3 10656 114 10656 114 0 FrameStrobe[9]
rlabel metal2 16440 9660 16440 9660 0 FrameStrobe_O[0]
rlabel metal2 18120 8904 18120 8904 0 FrameStrobe_O[10]
rlabel metal2 18600 9576 18600 9576 0 FrameStrobe_O[11]
rlabel metal2 18504 8820 18504 8820 0 FrameStrobe_O[12]
rlabel metal2 19320 9660 19320 9660 0 FrameStrobe_O[13]
rlabel metal2 18552 8148 18552 8148 0 FrameStrobe_O[14]
rlabel metal2 18840 8064 18840 8064 0 FrameStrobe_O[15]
rlabel metal2 19992 8904 19992 8904 0 FrameStrobe_O[16]
rlabel metal2 19128 6972 19128 6972 0 FrameStrobe_O[17]
rlabel metal2 18264 8148 18264 8148 0 FrameStrobe_O[18]
rlabel metal2 17880 7728 17880 7728 0 FrameStrobe_O[19]
rlabel metal2 16824 9660 16824 9660 0 FrameStrobe_O[1]
rlabel metal2 15960 9576 15960 9576 0 FrameStrobe_O[2]
rlabel metal2 16920 9576 16920 9576 0 FrameStrobe_O[3]
rlabel metal2 16776 8904 16776 8904 0 FrameStrobe_O[4]
rlabel metal2 17496 9660 17496 9660 0 FrameStrobe_O[5]
rlabel metal2 17160 8820 17160 8820 0 FrameStrobe_O[6]
rlabel metal2 17640 9324 17640 9324 0 FrameStrobe_O[7]
rlabel metal2 18216 9660 18216 9660 0 FrameStrobe_O[8]
rlabel metal2 18216 9240 18216 9240 0 FrameStrobe_O[9]
rlabel metal2 1656 8904 1656 8904 0 N1BEG[0]
rlabel metal2 2040 8148 2040 8148 0 N1BEG[1]
rlabel metal2 1944 8652 1944 8652 0 N1BEG[2]
rlabel metal2 1800 9660 1800 9660 0 N1BEG[3]
rlabel metal2 2280 9576 2280 9576 0 N2BEG[0]
rlabel metal2 2472 9660 2472 9660 0 N2BEG[1]
rlabel metal2 2760 9576 2760 9576 0 N2BEG[2]
rlabel metal2 3192 8904 3192 8904 0 N2BEG[3]
rlabel metal2 3240 9660 3240 9660 0 N2BEG[4]
rlabel metal2 3576 8904 3576 8904 0 N2BEG[5]
rlabel metal2 3528 9660 3528 9660 0 N2BEG[6]
rlabel metal2 4056 8904 4056 8904 0 N2BEG[7]
rlabel metal2 4056 9660 4056 9660 0 N2BEGb[0]
rlabel metal2 4344 8904 4344 8904 0 N2BEGb[1]
rlabel metal2 4392 9576 4392 9576 0 N2BEGb[2]
rlabel metal2 4728 8904 4728 8904 0 N2BEGb[3]
rlabel metal2 4680 9492 4680 9492 0 N2BEGb[4]
rlabel metal2 5256 8904 5256 8904 0 N2BEGb[5]
rlabel metal2 5160 9660 5160 9660 0 N2BEGb[6]
rlabel metal2 5496 8820 5496 8820 0 N2BEGb[7]
rlabel metal2 5544 9660 5544 9660 0 N4BEG[0]
rlabel metal2 7464 9576 7464 9576 0 N4BEG[10]
rlabel metal2 7752 9660 7752 9660 0 N4BEG[11]
rlabel metal2 7896 9576 7896 9576 0 N4BEG[12]
rlabel metal2 8184 9660 8184 9660 0 N4BEG[13]
rlabel metal2 8952 9660 8952 9660 0 N4BEG[14]
rlabel metal2 8568 9660 8568 9660 0 N4BEG[15]
rlabel metal2 5880 8904 5880 8904 0 N4BEG[1]
rlabel metal2 5928 9660 5928 9660 0 N4BEG[2]
rlabel metal2 6264 8904 6264 8904 0 N4BEG[3]
rlabel metal2 6312 9660 6312 9660 0 N4BEG[4]
rlabel metal2 6648 8904 6648 8904 0 N4BEG[5]
rlabel metal2 6696 9660 6696 9660 0 N4BEG[6]
rlabel metal2 7032 8904 7032 8904 0 N4BEG[7]
rlabel metal2 7080 9660 7080 9660 0 N4BEG[8]
rlabel metal2 7416 8904 7416 8904 0 N4BEG[9]
rlabel metal3 8736 9462 8736 9462 0 S1END[0]
rlabel metal3 8928 10806 8928 10806 0 S1END[1]
rlabel metal2 2736 8652 2736 8652 0 S1END[2]
rlabel metal3 2304 9366 2304 9366 0 S1END[3]
rlabel metal3 11040 9882 11040 9882 0 S2END[0]
rlabel metal3 11232 9924 11232 9924 0 S2END[1]
rlabel metal3 11424 9420 11424 9420 0 S2END[2]
rlabel metal3 11616 9462 11616 9462 0 S2END[3]
rlabel metal3 11808 10680 11808 10680 0 S2END[4]
rlabel metal3 12000 8790 12000 8790 0 S2END[5]
rlabel metal3 12192 10092 12192 10092 0 S2END[6]
rlabel metal3 12384 7950 12384 7950 0 S2END[7]
rlabel metal3 9504 8370 9504 8370 0 S2MID[0]
rlabel metal3 9696 8412 9696 8412 0 S2MID[1]
rlabel metal3 9888 10932 9888 10932 0 S2MID[2]
rlabel metal4 8016 9996 8016 9996 0 S2MID[3]
rlabel metal3 10272 10470 10272 10470 0 S2MID[4]
rlabel metal3 10464 8664 10464 8664 0 S2MID[5]
rlabel metal3 2208 6552 2208 6552 0 S2MID[6]
rlabel metal3 10848 10260 10848 10260 0 S2MID[7]
rlabel metal2 13536 6888 13536 6888 0 S4END[0]
rlabel metal3 14496 10470 14496 10470 0 S4END[10]
rlabel metal3 14688 9084 14688 9084 0 S4END[11]
rlabel metal3 14880 10932 14880 10932 0 S4END[12]
rlabel metal3 15072 11100 15072 11100 0 S4END[13]
rlabel metal3 15264 10848 15264 10848 0 S4END[14]
rlabel metal3 15456 10848 15456 10848 0 S4END[15]
rlabel metal2 13824 7098 13824 7098 0 S4END[1]
rlabel metal3 13248 8946 13248 8946 0 S4END[2]
rlabel metal3 13152 9378 13152 9378 0 S4END[3]
rlabel metal3 13344 9504 13344 9504 0 S4END[4]
rlabel metal3 13056 6552 13056 6552 0 S4END[5]
rlabel metal3 13728 9504 13728 9504 0 S4END[6]
rlabel metal3 13920 9546 13920 9546 0 S4END[7]
rlabel metal3 14112 10932 14112 10932 0 S4END[8]
rlabel metal3 14304 10638 14304 10638 0 S4END[9]
rlabel metal3 1056 2508 1056 2508 0 UserCLK
rlabel metal2 15912 9660 15912 9660 0 UserCLKo
rlabel metal2 18768 1932 18768 1932 0 net1
rlabel metal2 20544 6468 20544 6468 0 net10
rlabel metal2 20160 7098 20160 7098 0 net11
rlabel metal2 17808 1932 17808 1932 0 net12
rlabel metal2 19944 5544 19944 5544 0 net13
rlabel metal2 19608 6636 19608 6636 0 net14
rlabel metal2 16392 4284 16392 4284 0 net15
rlabel metal2 18936 5880 18936 5880 0 net16
rlabel metal2 17400 5124 17400 5124 0 net17
rlabel metal3 17088 8190 17088 8190 0 net18
rlabel metal3 14976 7686 14976 7686 0 net19
rlabel metal2 19848 3444 19848 3444 0 net2
rlabel metal2 17520 7140 17520 7140 0 net20
rlabel metal3 16704 8274 16704 8274 0 net21
rlabel metal2 15840 8694 15840 8694 0 net22
rlabel metal2 17424 2688 17424 2688 0 net23
rlabel metal2 18072 8652 18072 8652 0 net24
rlabel metal3 16320 8148 16320 8148 0 net25
rlabel metal2 19344 1932 19344 1932 0 net26
rlabel metal2 18720 2646 18720 2646 0 net27
rlabel metal2 19632 1932 19632 1932 0 net28
rlabel metal2 20160 1974 20160 1974 0 net29
rlabel metal2 20064 3444 20064 3444 0 net3
rlabel metal2 17544 1680 17544 1680 0 net30
rlabel metal2 18984 2016 18984 2016 0 net31
rlabel metal3 20832 3990 20832 3990 0 net32
rlabel metal2 14592 2856 14592 2856 0 net33
rlabel metal2 13656 3612 13656 3612 0 net34
rlabel metal2 11280 5418 11280 5418 0 net35
rlabel metal2 12312 4284 12312 4284 0 net36
rlabel metal3 13056 5460 13056 5460 0 net37
rlabel metal2 18672 7980 18672 7980 0 net38
rlabel metal2 15336 3612 15336 3612 0 net39
rlabel metal2 18888 4956 18888 4956 0 net4
rlabel metal2 14328 1680 14328 1680 0 net40
rlabel metal2 15240 5628 15240 5628 0 net41
rlabel metal2 17592 3612 17592 3612 0 net42
rlabel metal2 18552 4284 18552 4284 0 net43
rlabel metal3 13824 7854 13824 7854 0 net44
rlabel metal2 15456 9534 15456 9534 0 net45
rlabel metal3 17376 7686 17376 7686 0 net46
rlabel metal3 6624 4662 6624 4662 0 net47
rlabel metal2 15552 9534 15552 9534 0 net48
rlabel metal2 9864 2436 9864 2436 0 net49
rlabel metal2 20160 4242 20160 4242 0 net5
rlabel metal3 15312 3948 15312 3948 0 net50
rlabel metal3 15072 3612 15072 3612 0 net51
rlabel metal3 15072 3066 15072 3066 0 net52
rlabel metal2 1248 8736 1248 8736 0 net53
rlabel metal3 2304 8232 2304 8232 0 net54
rlabel metal3 1632 8862 1632 8862 0 net55
rlabel metal2 1536 9324 1536 9324 0 net56
rlabel metal2 2664 8904 2664 8904 0 net57
rlabel metal2 1944 7140 1944 7140 0 net58
rlabel metal2 2496 9450 2496 9450 0 net59
rlabel metal4 15264 5460 15264 5460 0 net6
rlabel metal2 4008 5544 4008 5544 0 net60
rlabel metal2 4440 5460 4440 5460 0 net61
rlabel metal2 6648 4956 6648 4956 0 net62
rlabel metal2 7608 5040 7608 5040 0 net63
rlabel metal2 8088 4956 8088 4956 0 net64
rlabel metal2 3720 4116 3720 4116 0 net65
rlabel metal2 5832 5040 5832 5040 0 net66
rlabel metal2 7224 5628 7224 5628 0 net67
rlabel metal2 7416 6468 7416 6468 0 net68
rlabel metal2 10344 7140 10344 7140 0 net69
rlabel metal2 20016 4956 20016 4956 0 net7
rlabel metal2 7848 7056 7848 7056 0 net70
rlabel metal2 9912 8148 9912 8148 0 net71
rlabel metal2 10296 8148 10296 8148 0 net72
rlabel metal2 18168 7728 18168 7728 0 net73
rlabel metal2 11304 6636 11304 6636 0 net74
rlabel metal2 9864 6972 9864 6972 0 net75
rlabel metal2 11832 7140 11832 7140 0 net76
rlabel metal3 10752 8022 10752 8022 0 net77
rlabel metal2 13320 7140 13320 7140 0 net78
rlabel metal3 11520 8484 11520 8484 0 net79
rlabel metal2 19728 5628 19728 5628 0 net8
rlabel metal2 19128 8904 19128 8904 0 net80
rlabel metal2 19392 6846 19392 6846 0 net81
rlabel metal3 7200 7350 7200 7350 0 net82
rlabel metal2 17592 6972 17592 6972 0 net83
rlabel metal3 7008 6510 7008 6510 0 net84
rlabel metal2 17016 6972 17016 6972 0 net85
rlabel metal2 16440 6972 16440 6972 0 net86
rlabel metal3 6720 9282 6720 9282 0 net87
rlabel metal2 14904 7140 14904 7140 0 net88
rlabel metal3 16416 7140 16416 7140 0 net89
rlabel metal2 20160 5670 20160 5670 0 net9
<< properties >>
string FIXED_BBOX 0 0 21600 11844
<< end >>
