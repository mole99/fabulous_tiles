magic
tech ihp-sg13g2
magscale 1 2
timestamp 1743708260
<< metal1 >>
rect 1152 10604 52128 10628
rect 1152 10564 4928 10604
rect 4968 10564 5010 10604
rect 5050 10564 5092 10604
rect 5132 10564 5174 10604
rect 5214 10564 5256 10604
rect 5296 10564 20048 10604
rect 20088 10564 20130 10604
rect 20170 10564 20212 10604
rect 20252 10564 20294 10604
rect 20334 10564 20376 10604
rect 20416 10564 35168 10604
rect 35208 10564 35250 10604
rect 35290 10564 35332 10604
rect 35372 10564 35414 10604
rect 35454 10564 35496 10604
rect 35536 10564 50288 10604
rect 50328 10564 50370 10604
rect 50410 10564 50452 10604
rect 50492 10564 50534 10604
rect 50574 10564 50616 10604
rect 50656 10564 52128 10604
rect 1152 10540 52128 10564
rect 1659 10436 1701 10445
rect 1659 10396 1660 10436
rect 1700 10396 1701 10436
rect 1659 10387 1701 10396
rect 4155 10436 4197 10445
rect 4155 10396 4156 10436
rect 4196 10396 4197 10436
rect 4155 10387 4197 10396
rect 6651 10436 6693 10445
rect 6651 10396 6652 10436
rect 6692 10396 6693 10436
rect 6651 10387 6693 10396
rect 9147 10436 9189 10445
rect 9147 10396 9148 10436
rect 9188 10396 9189 10436
rect 9147 10387 9189 10396
rect 11643 10436 11685 10445
rect 11643 10396 11644 10436
rect 11684 10396 11685 10436
rect 11643 10387 11685 10396
rect 14139 10436 14181 10445
rect 14139 10396 14140 10436
rect 14180 10396 14181 10436
rect 14139 10387 14181 10396
rect 16635 10436 16677 10445
rect 16635 10396 16636 10436
rect 16676 10396 16677 10436
rect 16635 10387 16677 10396
rect 19131 10436 19173 10445
rect 19131 10396 19132 10436
rect 19172 10396 19173 10436
rect 19131 10387 19173 10396
rect 21627 10436 21669 10445
rect 21627 10396 21628 10436
rect 21668 10396 21669 10436
rect 21627 10387 21669 10396
rect 24123 10436 24165 10445
rect 24123 10396 24124 10436
rect 24164 10396 24165 10436
rect 24123 10387 24165 10396
rect 26619 10436 26661 10445
rect 26619 10396 26620 10436
rect 26660 10396 26661 10436
rect 26619 10387 26661 10396
rect 29115 10436 29157 10445
rect 29115 10396 29116 10436
rect 29156 10396 29157 10436
rect 29115 10387 29157 10396
rect 31611 10436 31653 10445
rect 31611 10396 31612 10436
rect 31652 10396 31653 10436
rect 31611 10387 31653 10396
rect 34107 10436 34149 10445
rect 34107 10396 34108 10436
rect 34148 10396 34149 10436
rect 34107 10387 34149 10396
rect 39099 10436 39141 10445
rect 39099 10396 39100 10436
rect 39140 10396 39141 10436
rect 39099 10387 39141 10396
rect 41595 10436 41637 10445
rect 41595 10396 41596 10436
rect 41636 10396 41637 10436
rect 41595 10387 41637 10396
rect 44091 10436 44133 10445
rect 44091 10396 44092 10436
rect 44132 10396 44133 10436
rect 44091 10387 44133 10396
rect 46587 10436 46629 10445
rect 46587 10396 46588 10436
rect 46628 10396 46629 10436
rect 46587 10387 46629 10396
rect 49083 10436 49125 10445
rect 49083 10396 49084 10436
rect 49124 10396 49125 10436
rect 49083 10387 49125 10396
rect 50523 10436 50565 10445
rect 50523 10396 50524 10436
rect 50564 10396 50565 10436
rect 50523 10387 50565 10396
rect 50907 10436 50949 10445
rect 50907 10396 50908 10436
rect 50948 10396 50949 10436
rect 50907 10387 50949 10396
rect 51771 10436 51813 10445
rect 51771 10396 51772 10436
rect 51812 10396 51813 10436
rect 51771 10387 51813 10396
rect 51291 10352 51333 10361
rect 51291 10312 51292 10352
rect 51332 10312 51333 10352
rect 51291 10303 51333 10312
rect 1899 10184 1941 10193
rect 1899 10144 1900 10184
rect 1940 10144 1941 10184
rect 1899 10135 1941 10144
rect 4395 10184 4437 10193
rect 4395 10144 4396 10184
rect 4436 10144 4437 10184
rect 4395 10135 4437 10144
rect 6891 10184 6933 10193
rect 6891 10144 6892 10184
rect 6932 10144 6933 10184
rect 6891 10135 6933 10144
rect 9387 10184 9429 10193
rect 9387 10144 9388 10184
rect 9428 10144 9429 10184
rect 9387 10135 9429 10144
rect 11883 10184 11925 10193
rect 11883 10144 11884 10184
rect 11924 10144 11925 10184
rect 11883 10135 11925 10144
rect 14379 10184 14421 10193
rect 14379 10144 14380 10184
rect 14420 10144 14421 10184
rect 14379 10135 14421 10144
rect 16875 10184 16917 10193
rect 16875 10144 16876 10184
rect 16916 10144 16917 10184
rect 16875 10135 16917 10144
rect 19371 10184 19413 10193
rect 19371 10144 19372 10184
rect 19412 10144 19413 10184
rect 19371 10135 19413 10144
rect 21867 10184 21909 10193
rect 21867 10144 21868 10184
rect 21908 10144 21909 10184
rect 21867 10135 21909 10144
rect 24363 10184 24405 10193
rect 24363 10144 24364 10184
rect 24404 10144 24405 10184
rect 24363 10135 24405 10144
rect 26859 10184 26901 10193
rect 26859 10144 26860 10184
rect 26900 10144 26901 10184
rect 26859 10135 26901 10144
rect 29355 10184 29397 10193
rect 29355 10144 29356 10184
rect 29396 10144 29397 10184
rect 29355 10135 29397 10144
rect 31851 10184 31893 10193
rect 31851 10144 31852 10184
rect 31892 10144 31893 10184
rect 31851 10135 31893 10144
rect 34347 10184 34389 10193
rect 34347 10144 34348 10184
rect 34388 10144 34389 10184
rect 34347 10135 34389 10144
rect 36603 10184 36645 10193
rect 36603 10144 36604 10184
rect 36644 10144 36645 10184
rect 36603 10135 36645 10144
rect 36843 10184 36885 10193
rect 36843 10144 36844 10184
rect 36884 10144 36885 10184
rect 36843 10135 36885 10144
rect 39339 10184 39381 10193
rect 39339 10144 39340 10184
rect 39380 10144 39381 10184
rect 39339 10135 39381 10144
rect 41835 10184 41877 10193
rect 41835 10144 41836 10184
rect 41876 10144 41877 10184
rect 41835 10135 41877 10144
rect 44331 10184 44373 10193
rect 44331 10144 44332 10184
rect 44372 10144 44373 10184
rect 44331 10135 44373 10144
rect 46827 10184 46869 10193
rect 46827 10144 46828 10184
rect 46868 10144 46869 10184
rect 46827 10135 46869 10144
rect 49323 10184 49365 10193
rect 49323 10144 49324 10184
rect 49364 10144 49365 10184
rect 49323 10135 49365 10144
rect 49611 10184 49653 10193
rect 49611 10144 49612 10184
rect 49652 10144 49653 10184
rect 49611 10135 49653 10144
rect 50091 10184 50133 10193
rect 50091 10144 50092 10184
rect 50132 10144 50133 10184
rect 50091 10135 50133 10144
rect 50283 10184 50325 10193
rect 50283 10144 50284 10184
rect 50324 10144 50325 10184
rect 50283 10135 50325 10144
rect 50667 10184 50709 10193
rect 50667 10144 50668 10184
rect 50708 10144 50709 10184
rect 50667 10135 50709 10144
rect 51051 10184 51093 10193
rect 51051 10144 51052 10184
rect 51092 10144 51093 10184
rect 51051 10135 51093 10144
rect 51435 10184 51477 10193
rect 51435 10144 51436 10184
rect 51476 10144 51477 10184
rect 51435 10135 51477 10144
rect 52011 10184 52053 10193
rect 52011 10144 52012 10184
rect 52052 10144 52053 10184
rect 52011 10135 52053 10144
rect 49851 10100 49893 10109
rect 49851 10060 49852 10100
rect 49892 10060 49893 10100
rect 49851 10051 49893 10060
rect 51675 10016 51717 10025
rect 51675 9976 51676 10016
rect 51716 9976 51717 10016
rect 51675 9967 51717 9976
rect 1152 9848 52128 9872
rect 1152 9808 3688 9848
rect 3728 9808 3770 9848
rect 3810 9808 3852 9848
rect 3892 9808 3934 9848
rect 3974 9808 4016 9848
rect 4056 9808 18808 9848
rect 18848 9808 18890 9848
rect 18930 9808 18972 9848
rect 19012 9808 19054 9848
rect 19094 9808 19136 9848
rect 19176 9808 33928 9848
rect 33968 9808 34010 9848
rect 34050 9808 34092 9848
rect 34132 9808 34174 9848
rect 34214 9808 34256 9848
rect 34296 9808 49048 9848
rect 49088 9808 49130 9848
rect 49170 9808 49212 9848
rect 49252 9808 49294 9848
rect 49334 9808 49376 9848
rect 49416 9808 52128 9848
rect 1152 9784 52128 9808
rect 13851 9680 13893 9689
rect 13851 9640 13852 9680
rect 13892 9640 13893 9680
rect 13851 9631 13893 9640
rect 15771 9680 15813 9689
rect 15771 9640 15772 9680
rect 15812 9640 15813 9680
rect 15771 9631 15813 9640
rect 18459 9680 18501 9689
rect 18459 9640 18460 9680
rect 18500 9640 18501 9680
rect 18459 9631 18501 9640
rect 20859 9680 20901 9689
rect 20859 9640 20860 9680
rect 20900 9640 20901 9680
rect 20859 9631 20901 9640
rect 23163 9680 23205 9689
rect 23163 9640 23164 9680
rect 23204 9640 23205 9680
rect 23163 9631 23205 9640
rect 24027 9680 24069 9689
rect 24027 9640 24028 9680
rect 24068 9640 24069 9680
rect 24027 9631 24069 9640
rect 25371 9680 25413 9689
rect 25371 9640 25372 9680
rect 25412 9640 25413 9680
rect 25371 9631 25413 9640
rect 26907 9680 26949 9689
rect 26907 9640 26908 9680
rect 26948 9640 26949 9680
rect 26907 9631 26949 9640
rect 27867 9680 27909 9689
rect 27867 9640 27868 9680
rect 27908 9640 27909 9680
rect 27867 9631 27909 9640
rect 29115 9680 29157 9689
rect 29115 9640 29116 9680
rect 29156 9640 29157 9680
rect 29115 9631 29157 9640
rect 29691 9680 29733 9689
rect 29691 9640 29692 9680
rect 29732 9640 29733 9680
rect 29691 9631 29733 9640
rect 41595 9680 41637 9689
rect 41595 9640 41596 9680
rect 41636 9640 41637 9680
rect 41595 9631 41637 9640
rect 43419 9680 43461 9689
rect 43419 9640 43420 9680
rect 43460 9640 43461 9680
rect 43419 9631 43461 9640
rect 43995 9680 44037 9689
rect 43995 9640 43996 9680
rect 44036 9640 44037 9680
rect 43995 9631 44037 9640
rect 44955 9680 44997 9689
rect 44955 9640 44956 9680
rect 44996 9640 44997 9680
rect 44955 9631 44997 9640
rect 46203 9680 46245 9689
rect 46203 9640 46204 9680
rect 46244 9640 46245 9680
rect 46203 9631 46245 9640
rect 46683 9680 46725 9689
rect 46683 9640 46684 9680
rect 46724 9640 46725 9680
rect 46683 9631 46725 9640
rect 48219 9680 48261 9689
rect 48219 9640 48220 9680
rect 48260 9640 48261 9680
rect 48219 9631 48261 9640
rect 48891 9680 48933 9689
rect 48891 9640 48892 9680
rect 48932 9640 48933 9680
rect 48891 9631 48933 9640
rect 50811 9680 50853 9689
rect 50811 9640 50812 9680
rect 50852 9640 50853 9680
rect 50811 9631 50853 9640
rect 51195 9680 51237 9689
rect 51195 9640 51196 9680
rect 51236 9640 51237 9680
rect 51195 9631 51237 9640
rect 40635 9596 40677 9605
rect 40635 9556 40636 9596
rect 40676 9556 40677 9596
rect 40635 9547 40677 9556
rect 13707 9512 13749 9521
rect 13707 9472 13708 9512
rect 13748 9472 13749 9512
rect 13707 9463 13749 9472
rect 14091 9512 14133 9521
rect 14091 9472 14092 9512
rect 14132 9472 14133 9512
rect 14091 9463 14133 9472
rect 14283 9512 14325 9521
rect 14283 9472 14284 9512
rect 14324 9472 14325 9512
rect 14283 9463 14325 9472
rect 14523 9512 14565 9521
rect 14523 9472 14524 9512
rect 14564 9472 14565 9512
rect 14523 9463 14565 9472
rect 15627 9512 15669 9521
rect 15627 9472 15628 9512
rect 15668 9472 15669 9512
rect 15627 9463 15669 9472
rect 16011 9512 16053 9521
rect 16011 9472 16012 9512
rect 16052 9472 16053 9512
rect 16011 9463 16053 9472
rect 18699 9512 18741 9521
rect 18699 9472 18700 9512
rect 18740 9472 18741 9512
rect 18699 9463 18741 9472
rect 21099 9512 21141 9521
rect 21099 9472 21100 9512
rect 21140 9472 21141 9512
rect 21099 9463 21141 9472
rect 23403 9512 23445 9521
rect 23403 9472 23404 9512
rect 23444 9472 23445 9512
rect 23403 9463 23445 9472
rect 23787 9512 23829 9521
rect 23787 9472 23788 9512
rect 23828 9472 23829 9512
rect 23787 9463 23829 9472
rect 25611 9512 25653 9521
rect 25611 9472 25612 9512
rect 25652 9472 25653 9512
rect 25611 9463 25653 9472
rect 26187 9512 26229 9521
rect 26187 9472 26188 9512
rect 26228 9472 26229 9512
rect 26187 9463 26229 9472
rect 26667 9512 26709 9521
rect 26667 9472 26668 9512
rect 26708 9472 26709 9512
rect 26667 9463 26709 9472
rect 28107 9512 28149 9521
rect 28107 9472 28108 9512
rect 28148 9472 28149 9512
rect 28107 9463 28149 9472
rect 28875 9512 28917 9521
rect 28875 9472 28876 9512
rect 28916 9472 28917 9512
rect 28875 9463 28917 9472
rect 29931 9512 29973 9521
rect 29931 9472 29932 9512
rect 29972 9472 29973 9512
rect 29931 9463 29973 9472
rect 30219 9512 30261 9521
rect 30219 9472 30220 9512
rect 30260 9472 30261 9512
rect 30219 9463 30261 9472
rect 30459 9512 30501 9521
rect 30459 9472 30460 9512
rect 30500 9472 30501 9512
rect 30459 9463 30501 9472
rect 40299 9512 40341 9521
rect 40299 9472 40300 9512
rect 40340 9472 40341 9512
rect 40299 9463 40341 9472
rect 40875 9512 40917 9521
rect 40875 9472 40876 9512
rect 40916 9472 40917 9512
rect 40875 9463 40917 9472
rect 41835 9512 41877 9521
rect 41835 9472 41836 9512
rect 41876 9472 41877 9512
rect 41835 9463 41877 9472
rect 42795 9512 42837 9521
rect 42795 9472 42796 9512
rect 42836 9472 42837 9512
rect 42795 9463 42837 9472
rect 43659 9512 43701 9521
rect 43659 9472 43660 9512
rect 43700 9472 43701 9512
rect 43659 9463 43701 9472
rect 44235 9512 44277 9521
rect 44235 9472 44236 9512
rect 44276 9472 44277 9512
rect 44235 9463 44277 9472
rect 45195 9512 45237 9521
rect 45195 9472 45196 9512
rect 45236 9472 45237 9512
rect 45195 9463 45237 9472
rect 46491 9512 46533 9521
rect 46491 9472 46492 9512
rect 46532 9472 46533 9512
rect 46491 9463 46533 9472
rect 46923 9512 46965 9521
rect 46923 9472 46924 9512
rect 46964 9472 46965 9512
rect 46923 9463 46965 9472
rect 47307 9512 47349 9521
rect 47307 9472 47308 9512
rect 47348 9472 47349 9512
rect 47307 9463 47349 9472
rect 48459 9512 48501 9521
rect 48459 9472 48460 9512
rect 48500 9472 48501 9512
rect 48459 9463 48501 9472
rect 48651 9512 48693 9521
rect 48651 9472 48652 9512
rect 48692 9472 48693 9512
rect 48651 9463 48693 9472
rect 50571 9512 50613 9521
rect 50571 9472 50572 9512
rect 50612 9472 50613 9512
rect 50571 9463 50613 9472
rect 50955 9512 50997 9521
rect 50955 9472 50956 9512
rect 50996 9472 50997 9512
rect 50955 9463 50997 9472
rect 51435 9512 51477 9521
rect 51435 9472 51436 9512
rect 51476 9472 51477 9512
rect 51435 9463 51477 9472
rect 51819 9512 51861 9521
rect 51819 9472 51820 9512
rect 51860 9472 51861 9512
rect 51819 9463 51861 9472
rect 40059 9344 40101 9353
rect 40059 9304 40060 9344
rect 40100 9304 40101 9344
rect 40059 9295 40101 9304
rect 15610 9260 15668 9261
rect 15610 9220 15619 9260
rect 15659 9220 15668 9260
rect 15610 9219 15668 9220
rect 26427 9260 26469 9269
rect 26427 9220 26428 9260
rect 26468 9220 26469 9260
rect 26427 9211 26469 9220
rect 42555 9260 42597 9269
rect 42555 9220 42556 9260
rect 42596 9220 42597 9260
rect 42555 9211 42597 9220
rect 47067 9260 47109 9269
rect 47067 9220 47068 9260
rect 47108 9220 47109 9260
rect 47067 9211 47109 9220
rect 50266 9260 50324 9261
rect 50266 9220 50275 9260
rect 50315 9220 50324 9260
rect 50266 9219 50324 9220
rect 51675 9260 51717 9269
rect 51675 9220 51676 9260
rect 51716 9220 51717 9260
rect 51675 9211 51717 9220
rect 52059 9260 52101 9269
rect 52059 9220 52060 9260
rect 52100 9220 52101 9260
rect 52059 9211 52101 9220
rect 1152 9092 52128 9116
rect 1152 9052 4928 9092
rect 4968 9052 5010 9092
rect 5050 9052 5092 9092
rect 5132 9052 5174 9092
rect 5214 9052 5256 9092
rect 5296 9052 20048 9092
rect 20088 9052 20130 9092
rect 20170 9052 20212 9092
rect 20252 9052 20294 9092
rect 20334 9052 20376 9092
rect 20416 9052 35168 9092
rect 35208 9052 35250 9092
rect 35290 9052 35332 9092
rect 35372 9052 35414 9092
rect 35454 9052 35496 9092
rect 35536 9052 50288 9092
rect 50328 9052 50370 9092
rect 50410 9052 50452 9092
rect 50492 9052 50534 9092
rect 50574 9052 50616 9092
rect 50656 9052 52128 9092
rect 1152 9028 52128 9052
rect 33723 8924 33765 8933
rect 33723 8884 33724 8924
rect 33764 8884 33765 8924
rect 33723 8875 33765 8884
rect 25851 8840 25893 8849
rect 25851 8800 25852 8840
rect 25892 8800 25893 8840
rect 25851 8791 25893 8800
rect 28347 8840 28389 8849
rect 28347 8800 28348 8840
rect 28388 8800 28389 8840
rect 28347 8791 28389 8800
rect 25611 8672 25653 8681
rect 25611 8632 25612 8672
rect 25652 8632 25653 8672
rect 25611 8623 25653 8632
rect 27723 8672 27765 8681
rect 27723 8632 27724 8672
rect 27764 8632 27765 8672
rect 27723 8623 27765 8632
rect 27963 8672 28005 8681
rect 27963 8632 27964 8672
rect 28004 8632 28005 8672
rect 27963 8623 28005 8632
rect 28107 8672 28149 8681
rect 28107 8632 28108 8672
rect 28148 8632 28149 8672
rect 28107 8623 28149 8632
rect 33291 8672 33333 8681
rect 33291 8632 33292 8672
rect 33332 8632 33333 8672
rect 33291 8623 33333 8632
rect 33483 8672 33525 8681
rect 33483 8632 33484 8672
rect 33524 8632 33525 8672
rect 33483 8623 33525 8632
rect 33963 8672 34005 8681
rect 33963 8632 33964 8672
rect 34004 8632 34005 8672
rect 33963 8623 34005 8632
rect 34251 8672 34293 8681
rect 34251 8632 34252 8672
rect 34292 8632 34293 8672
rect 34251 8623 34293 8632
rect 34539 8672 34581 8681
rect 34539 8632 34540 8672
rect 34580 8632 34581 8672
rect 34539 8623 34581 8632
rect 34827 8672 34869 8681
rect 34827 8632 34828 8672
rect 34868 8632 34869 8672
rect 34827 8623 34869 8632
rect 35115 8672 35157 8681
rect 35115 8632 35116 8672
rect 35156 8632 35157 8672
rect 35115 8623 35157 8632
rect 35403 8672 35445 8681
rect 35403 8632 35404 8672
rect 35444 8632 35445 8672
rect 35403 8623 35445 8632
rect 35691 8672 35733 8681
rect 35691 8632 35692 8672
rect 35732 8632 35733 8672
rect 35691 8623 35733 8632
rect 35883 8672 35925 8681
rect 35883 8632 35884 8672
rect 35924 8632 35925 8672
rect 35883 8623 35925 8632
rect 51435 8672 51477 8681
rect 51435 8632 51436 8672
rect 51476 8632 51477 8672
rect 51435 8623 51477 8632
rect 51675 8672 51717 8681
rect 51675 8632 51676 8672
rect 51716 8632 51717 8672
rect 51675 8623 51717 8632
rect 51819 8672 51861 8681
rect 51819 8632 51820 8672
rect 51860 8632 51861 8672
rect 51819 8623 51861 8632
rect 52059 8672 52101 8681
rect 52059 8632 52060 8672
rect 52100 8632 52101 8672
rect 52059 8623 52101 8632
rect 1152 8336 52128 8360
rect 1152 8296 3688 8336
rect 3728 8296 3770 8336
rect 3810 8296 3852 8336
rect 3892 8296 3934 8336
rect 3974 8296 4016 8336
rect 4056 8296 18808 8336
rect 18848 8296 18890 8336
rect 18930 8296 18972 8336
rect 19012 8296 19054 8336
rect 19094 8296 19136 8336
rect 19176 8296 33928 8336
rect 33968 8296 34010 8336
rect 34050 8296 34092 8336
rect 34132 8296 34174 8336
rect 34214 8296 34256 8336
rect 34296 8296 49048 8336
rect 49088 8296 49130 8336
rect 49170 8296 49212 8336
rect 49252 8296 49294 8336
rect 49334 8296 49376 8336
rect 49416 8296 52128 8336
rect 1152 8272 52128 8296
rect 23547 8168 23589 8177
rect 23547 8128 23548 8168
rect 23588 8128 23589 8168
rect 23547 8119 23589 8128
rect 28251 8168 28293 8177
rect 28251 8128 28252 8168
rect 28292 8128 28293 8168
rect 28251 8119 28293 8128
rect 31707 8084 31749 8093
rect 31707 8044 31708 8084
rect 31748 8044 31749 8084
rect 31707 8035 31749 8044
rect 23307 8000 23349 8009
rect 23307 7960 23308 8000
rect 23348 7960 23349 8000
rect 23307 7951 23349 7960
rect 28011 8000 28053 8009
rect 28011 7960 28012 8000
rect 28052 7960 28053 8000
rect 28011 7951 28053 7960
rect 31467 8000 31509 8009
rect 31467 7960 31468 8000
rect 31508 7960 31509 8000
rect 31467 7951 31509 7960
rect 35211 8000 35253 8009
rect 35211 7960 35212 8000
rect 35252 7960 35253 8000
rect 35211 7951 35253 7960
rect 51435 8000 51477 8009
rect 51435 7960 51436 8000
rect 51476 7960 51477 8000
rect 51435 7951 51477 7960
rect 51819 8000 51861 8009
rect 51819 7960 51820 8000
rect 51860 7960 51861 8000
rect 51819 7951 51861 7960
rect 51675 7832 51717 7841
rect 51675 7792 51676 7832
rect 51716 7792 51717 7832
rect 51675 7783 51717 7792
rect 33466 7748 33524 7749
rect 33466 7708 33475 7748
rect 33515 7708 33524 7748
rect 33466 7707 33524 7708
rect 35451 7748 35493 7757
rect 35451 7708 35452 7748
rect 35492 7708 35493 7748
rect 35451 7699 35493 7708
rect 52059 7748 52101 7757
rect 52059 7708 52060 7748
rect 52100 7708 52101 7748
rect 52059 7699 52101 7708
rect 1152 7580 52128 7604
rect 1152 7540 4928 7580
rect 4968 7540 5010 7580
rect 5050 7540 5092 7580
rect 5132 7540 5174 7580
rect 5214 7540 5256 7580
rect 5296 7540 20048 7580
rect 20088 7540 20130 7580
rect 20170 7540 20212 7580
rect 20252 7540 20294 7580
rect 20334 7540 20376 7580
rect 20416 7540 35168 7580
rect 35208 7540 35250 7580
rect 35290 7540 35332 7580
rect 35372 7540 35414 7580
rect 35454 7540 35496 7580
rect 35536 7540 50288 7580
rect 50328 7540 50370 7580
rect 50410 7540 50452 7580
rect 50492 7540 50534 7580
rect 50574 7540 50616 7580
rect 50656 7540 52128 7580
rect 1152 7516 52128 7540
rect 35211 7328 35253 7337
rect 35211 7288 35212 7328
rect 35252 7288 35253 7328
rect 35211 7279 35253 7288
rect 35499 7328 35541 7337
rect 35499 7288 35500 7328
rect 35540 7288 35541 7328
rect 35499 7279 35541 7288
rect 18891 7160 18933 7169
rect 18891 7120 18892 7160
rect 18932 7120 18933 7160
rect 18891 7111 18933 7120
rect 23595 7160 23637 7169
rect 23595 7120 23596 7160
rect 23636 7120 23637 7160
rect 23595 7111 23637 7120
rect 23835 7160 23877 7169
rect 23835 7120 23836 7160
rect 23876 7120 23877 7160
rect 23835 7111 23877 7120
rect 29739 7160 29781 7169
rect 29739 7120 29740 7160
rect 29780 7120 29781 7160
rect 29739 7111 29781 7120
rect 30219 7160 30261 7169
rect 30219 7120 30220 7160
rect 30260 7120 30261 7160
rect 30219 7111 30261 7120
rect 51435 7160 51477 7169
rect 51435 7120 51436 7160
rect 51476 7120 51477 7160
rect 51435 7111 51477 7120
rect 51819 7160 51861 7169
rect 51819 7120 51820 7160
rect 51860 7120 51861 7160
rect 51819 7111 51861 7120
rect 52059 7160 52101 7169
rect 52059 7120 52060 7160
rect 52100 7120 52101 7160
rect 52059 7111 52101 7120
rect 30459 7076 30501 7085
rect 30459 7036 30460 7076
rect 30500 7036 30501 7076
rect 30459 7027 30501 7036
rect 19131 6992 19173 7001
rect 19131 6952 19132 6992
rect 19172 6952 19173 6992
rect 19131 6943 19173 6952
rect 29979 6992 30021 7001
rect 29979 6952 29980 6992
rect 30020 6952 30021 6992
rect 29979 6943 30021 6952
rect 51675 6992 51717 7001
rect 51675 6952 51676 6992
rect 51716 6952 51717 6992
rect 51675 6943 51717 6952
rect 1152 6824 52128 6848
rect 1152 6784 3688 6824
rect 3728 6784 3770 6824
rect 3810 6784 3852 6824
rect 3892 6784 3934 6824
rect 3974 6784 4016 6824
rect 4056 6784 18808 6824
rect 18848 6784 18890 6824
rect 18930 6784 18972 6824
rect 19012 6784 19054 6824
rect 19094 6784 19136 6824
rect 19176 6784 33928 6824
rect 33968 6784 34010 6824
rect 34050 6784 34092 6824
rect 34132 6784 34174 6824
rect 34214 6784 34256 6824
rect 34296 6784 49048 6824
rect 49088 6784 49130 6824
rect 49170 6784 49212 6824
rect 49252 6784 49294 6824
rect 49334 6784 49376 6824
rect 49416 6784 52128 6824
rect 1152 6760 52128 6784
rect 25659 6572 25701 6581
rect 25659 6532 25660 6572
rect 25700 6532 25701 6572
rect 25659 6523 25701 6532
rect 22731 6488 22773 6497
rect 22731 6448 22732 6488
rect 22772 6448 22773 6488
rect 22731 6439 22773 6448
rect 25419 6488 25461 6497
rect 25419 6448 25420 6488
rect 25460 6448 25461 6488
rect 25419 6439 25461 6448
rect 25803 6488 25845 6497
rect 25803 6448 25804 6488
rect 25844 6448 25845 6488
rect 25803 6439 25845 6448
rect 35499 6488 35541 6497
rect 35499 6448 35500 6488
rect 35540 6448 35541 6488
rect 35499 6439 35541 6448
rect 35787 6488 35829 6497
rect 35787 6448 35788 6488
rect 35828 6448 35829 6488
rect 35787 6439 35829 6448
rect 36171 6488 36213 6497
rect 36171 6448 36172 6488
rect 36212 6448 36213 6488
rect 36171 6439 36213 6448
rect 36459 6488 36501 6497
rect 36459 6448 36460 6488
rect 36500 6448 36501 6488
rect 36459 6439 36501 6448
rect 36747 6488 36789 6497
rect 36747 6448 36748 6488
rect 36788 6448 36789 6488
rect 36747 6439 36789 6448
rect 37035 6488 37077 6497
rect 37035 6448 37036 6488
rect 37076 6448 37077 6488
rect 37035 6439 37077 6448
rect 37323 6488 37365 6497
rect 37323 6448 37324 6488
rect 37364 6448 37365 6488
rect 37323 6439 37365 6448
rect 37611 6488 37653 6497
rect 37611 6448 37612 6488
rect 37652 6448 37653 6488
rect 37611 6439 37653 6448
rect 37899 6488 37941 6497
rect 37899 6448 37900 6488
rect 37940 6448 37941 6488
rect 37899 6439 37941 6448
rect 38283 6488 38325 6497
rect 38283 6448 38284 6488
rect 38324 6448 38325 6488
rect 38283 6439 38325 6448
rect 51435 6488 51477 6497
rect 51435 6448 51436 6488
rect 51476 6448 51477 6488
rect 51435 6439 51477 6448
rect 51819 6488 51861 6497
rect 51819 6448 51820 6488
rect 51860 6448 51861 6488
rect 51819 6439 51861 6448
rect 52059 6488 52101 6497
rect 52059 6448 52060 6488
rect 52100 6448 52101 6488
rect 52059 6439 52101 6448
rect 26043 6320 26085 6329
rect 26043 6280 26044 6320
rect 26084 6280 26085 6320
rect 26043 6271 26085 6280
rect 22971 6236 23013 6245
rect 22971 6196 22972 6236
rect 23012 6196 23013 6236
rect 22971 6187 23013 6196
rect 36027 6236 36069 6245
rect 36027 6196 36028 6236
rect 36068 6196 36069 6236
rect 36027 6187 36069 6196
rect 38523 6236 38565 6245
rect 38523 6196 38524 6236
rect 38564 6196 38565 6236
rect 38523 6187 38565 6196
rect 51675 6236 51717 6245
rect 51675 6196 51676 6236
rect 51716 6196 51717 6236
rect 51675 6187 51717 6196
rect 1152 6068 52128 6092
rect 1152 6028 4928 6068
rect 4968 6028 5010 6068
rect 5050 6028 5092 6068
rect 5132 6028 5174 6068
rect 5214 6028 5256 6068
rect 5296 6028 20048 6068
rect 20088 6028 20130 6068
rect 20170 6028 20212 6068
rect 20252 6028 20294 6068
rect 20334 6028 20376 6068
rect 20416 6028 35168 6068
rect 35208 6028 35250 6068
rect 35290 6028 35332 6068
rect 35372 6028 35414 6068
rect 35454 6028 35496 6068
rect 35536 6028 50288 6068
rect 50328 6028 50370 6068
rect 50410 6028 50452 6068
rect 50492 6028 50534 6068
rect 50574 6028 50616 6068
rect 50656 6028 52128 6068
rect 1152 6004 52128 6028
rect 35787 5816 35829 5825
rect 35787 5776 35788 5816
rect 35828 5776 35829 5816
rect 35787 5767 35829 5776
rect 36075 5816 36117 5825
rect 36075 5776 36076 5816
rect 36116 5776 36117 5816
rect 36075 5767 36117 5776
rect 52059 5816 52101 5825
rect 52059 5776 52060 5816
rect 52100 5776 52101 5816
rect 52059 5767 52101 5776
rect 23883 5648 23925 5657
rect 23883 5608 23884 5648
rect 23924 5608 23925 5648
rect 23883 5599 23925 5608
rect 24123 5648 24165 5657
rect 24123 5608 24124 5648
rect 24164 5608 24165 5648
rect 24123 5599 24165 5608
rect 27819 5648 27861 5657
rect 27819 5608 27820 5648
rect 27860 5608 27861 5648
rect 27819 5599 27861 5608
rect 51435 5648 51477 5657
rect 51435 5608 51436 5648
rect 51476 5608 51477 5648
rect 51435 5599 51477 5608
rect 51819 5648 51861 5657
rect 51819 5608 51820 5648
rect 51860 5608 51861 5648
rect 51819 5599 51861 5608
rect 51675 5564 51717 5573
rect 51675 5524 51676 5564
rect 51716 5524 51717 5564
rect 51675 5515 51717 5524
rect 28059 5480 28101 5489
rect 28059 5440 28060 5480
rect 28100 5440 28101 5480
rect 28059 5431 28101 5440
rect 1152 5312 52128 5336
rect 1152 5272 3688 5312
rect 3728 5272 3770 5312
rect 3810 5272 3852 5312
rect 3892 5272 3934 5312
rect 3974 5272 4016 5312
rect 4056 5272 18808 5312
rect 18848 5272 18890 5312
rect 18930 5272 18972 5312
rect 19012 5272 19054 5312
rect 19094 5272 19136 5312
rect 19176 5272 33928 5312
rect 33968 5272 34010 5312
rect 34050 5272 34092 5312
rect 34132 5272 34174 5312
rect 34214 5272 34256 5312
rect 34296 5272 49048 5312
rect 49088 5272 49130 5312
rect 49170 5272 49212 5312
rect 49252 5272 49294 5312
rect 49334 5272 49376 5312
rect 49416 5272 52128 5312
rect 1152 5248 52128 5272
rect 52059 5144 52101 5153
rect 52059 5104 52060 5144
rect 52100 5104 52101 5144
rect 52059 5095 52101 5104
rect 14667 4976 14709 4985
rect 14667 4936 14668 4976
rect 14708 4936 14709 4976
rect 14667 4927 14709 4936
rect 15243 4976 15285 4985
rect 15243 4936 15244 4976
rect 15284 4936 15285 4976
rect 15243 4927 15285 4936
rect 24171 4976 24213 4985
rect 24171 4936 24172 4976
rect 24212 4936 24213 4976
rect 24171 4927 24213 4936
rect 24843 4976 24885 4985
rect 24843 4936 24844 4976
rect 24884 4936 24885 4976
rect 24843 4927 24885 4936
rect 25227 4976 25269 4985
rect 25227 4936 25228 4976
rect 25268 4936 25269 4976
rect 25227 4927 25269 4936
rect 30027 4976 30069 4985
rect 30027 4936 30028 4976
rect 30068 4936 30069 4976
rect 30027 4927 30069 4936
rect 51435 4976 51477 4985
rect 51435 4936 51436 4976
rect 51476 4936 51477 4976
rect 51435 4927 51477 4936
rect 51819 4976 51861 4985
rect 51819 4936 51820 4976
rect 51860 4936 51861 4976
rect 51819 4927 51861 4936
rect 30267 4808 30309 4817
rect 30267 4768 30268 4808
rect 30308 4768 30309 4808
rect 30267 4759 30309 4768
rect 51675 4808 51717 4817
rect 51675 4768 51676 4808
rect 51716 4768 51717 4808
rect 51675 4759 51717 4768
rect 14907 4724 14949 4733
rect 14907 4684 14908 4724
rect 14948 4684 14949 4724
rect 14907 4675 14949 4684
rect 15483 4724 15525 4733
rect 15483 4684 15484 4724
rect 15524 4684 15525 4724
rect 15483 4675 15525 4684
rect 24411 4724 24453 4733
rect 24411 4684 24412 4724
rect 24452 4684 24453 4724
rect 24411 4675 24453 4684
rect 25083 4724 25125 4733
rect 25083 4684 25084 4724
rect 25124 4684 25125 4724
rect 25083 4675 25125 4684
rect 25467 4724 25509 4733
rect 25467 4684 25468 4724
rect 25508 4684 25509 4724
rect 25467 4675 25509 4684
rect 1152 4556 52128 4580
rect 1152 4516 4928 4556
rect 4968 4516 5010 4556
rect 5050 4516 5092 4556
rect 5132 4516 5174 4556
rect 5214 4516 5256 4556
rect 5296 4516 20048 4556
rect 20088 4516 20130 4556
rect 20170 4516 20212 4556
rect 20252 4516 20294 4556
rect 20334 4516 20376 4556
rect 20416 4516 35168 4556
rect 35208 4516 35250 4556
rect 35290 4516 35332 4556
rect 35372 4516 35414 4556
rect 35454 4516 35496 4556
rect 35536 4516 50288 4556
rect 50328 4516 50370 4556
rect 50410 4516 50452 4556
rect 50492 4516 50534 4556
rect 50574 4516 50616 4556
rect 50656 4516 52128 4556
rect 1152 4492 52128 4516
rect 52059 4304 52101 4313
rect 52059 4264 52060 4304
rect 52100 4264 52101 4304
rect 52059 4255 52101 4264
rect 13419 4136 13461 4145
rect 13419 4096 13420 4136
rect 13460 4096 13461 4136
rect 13419 4087 13461 4096
rect 16395 4136 16437 4145
rect 16395 4096 16396 4136
rect 16436 4096 16437 4136
rect 16395 4087 16437 4096
rect 16875 4136 16917 4145
rect 16875 4096 16876 4136
rect 16916 4096 16917 4136
rect 16875 4087 16917 4096
rect 19179 4136 19221 4145
rect 19179 4096 19180 4136
rect 19220 4096 19221 4136
rect 19179 4087 19221 4096
rect 23019 4136 23061 4145
rect 23019 4096 23020 4136
rect 23060 4096 23061 4136
rect 23019 4087 23061 4096
rect 28011 4136 28053 4145
rect 28011 4096 28012 4136
rect 28052 4096 28053 4136
rect 28011 4087 28053 4096
rect 38859 4136 38901 4145
rect 38859 4096 38860 4136
rect 38900 4096 38901 4136
rect 38859 4087 38901 4096
rect 50859 4136 50901 4145
rect 50859 4096 50860 4136
rect 50900 4096 50901 4136
rect 50859 4087 50901 4096
rect 51051 4136 51093 4145
rect 51051 4096 51052 4136
rect 51092 4096 51093 4136
rect 51051 4087 51093 4096
rect 51435 4136 51477 4145
rect 51435 4096 51436 4136
rect 51476 4096 51477 4136
rect 51435 4087 51477 4096
rect 51819 4136 51861 4145
rect 51819 4096 51820 4136
rect 51860 4096 51861 4136
rect 51819 4087 51861 4096
rect 28251 4052 28293 4061
rect 28251 4012 28252 4052
rect 28292 4012 28293 4052
rect 28251 4003 28293 4012
rect 51675 4052 51717 4061
rect 51675 4012 51676 4052
rect 51716 4012 51717 4052
rect 51675 4003 51717 4012
rect 13659 3968 13701 3977
rect 13659 3928 13660 3968
rect 13700 3928 13701 3968
rect 13659 3919 13701 3928
rect 16635 3968 16677 3977
rect 16635 3928 16636 3968
rect 16676 3928 16677 3968
rect 16635 3919 16677 3928
rect 17115 3968 17157 3977
rect 17115 3928 17116 3968
rect 17156 3928 17157 3968
rect 17115 3919 17157 3928
rect 19419 3968 19461 3977
rect 19419 3928 19420 3968
rect 19460 3928 19461 3968
rect 19419 3919 19461 3928
rect 23259 3968 23301 3977
rect 23259 3928 23260 3968
rect 23300 3928 23301 3968
rect 23259 3919 23301 3928
rect 38619 3968 38661 3977
rect 38619 3928 38620 3968
rect 38660 3928 38661 3968
rect 38619 3919 38661 3928
rect 51291 3968 51333 3977
rect 51291 3928 51292 3968
rect 51332 3928 51333 3968
rect 51291 3919 51333 3928
rect 1152 3800 52128 3824
rect 1152 3760 3688 3800
rect 3728 3760 3770 3800
rect 3810 3760 3852 3800
rect 3892 3760 3934 3800
rect 3974 3760 4016 3800
rect 4056 3760 18808 3800
rect 18848 3760 18890 3800
rect 18930 3760 18972 3800
rect 19012 3760 19054 3800
rect 19094 3760 19136 3800
rect 19176 3760 33928 3800
rect 33968 3760 34010 3800
rect 34050 3760 34092 3800
rect 34132 3760 34174 3800
rect 34214 3760 34256 3800
rect 34296 3760 49048 3800
rect 49088 3760 49130 3800
rect 49170 3760 49212 3800
rect 49252 3760 49294 3800
rect 49334 3760 49376 3800
rect 49416 3760 52128 3800
rect 1152 3736 52128 3760
rect 22779 3632 22821 3641
rect 22779 3592 22780 3632
rect 22820 3592 22821 3632
rect 22779 3583 22821 3592
rect 52059 3632 52101 3641
rect 52059 3592 52060 3632
rect 52100 3592 52101 3632
rect 52059 3583 52101 3592
rect 19803 3548 19845 3557
rect 19803 3508 19804 3548
rect 19844 3508 19845 3548
rect 19803 3499 19845 3508
rect 14187 3464 14229 3473
rect 14187 3424 14188 3464
rect 14228 3424 14229 3464
rect 14187 3415 14229 3424
rect 14667 3464 14709 3473
rect 14667 3424 14668 3464
rect 14708 3424 14709 3464
rect 14667 3415 14709 3424
rect 17115 3464 17157 3473
rect 17115 3424 17116 3464
rect 17156 3424 17157 3464
rect 17115 3415 17157 3424
rect 19563 3464 19605 3473
rect 19563 3424 19564 3464
rect 19604 3424 19605 3464
rect 19563 3415 19605 3424
rect 21291 3464 21333 3473
rect 21291 3424 21292 3464
rect 21332 3424 21333 3464
rect 21291 3415 21333 3424
rect 21531 3464 21573 3473
rect 21531 3424 21532 3464
rect 21572 3424 21573 3464
rect 21531 3415 21573 3424
rect 21706 3464 21764 3465
rect 21706 3424 21715 3464
rect 21755 3424 21764 3464
rect 21706 3423 21764 3424
rect 22539 3464 22581 3473
rect 22539 3424 22540 3464
rect 22580 3424 22581 3464
rect 22539 3415 22581 3424
rect 28203 3464 28245 3473
rect 28203 3424 28204 3464
rect 28244 3424 28245 3464
rect 28203 3415 28245 3424
rect 29643 3464 29685 3473
rect 29643 3424 29644 3464
rect 29684 3424 29685 3464
rect 29643 3415 29685 3424
rect 30411 3464 30453 3473
rect 30411 3424 30412 3464
rect 30452 3424 30453 3464
rect 30411 3415 30453 3424
rect 30795 3464 30837 3473
rect 30795 3424 30796 3464
rect 30836 3424 30837 3464
rect 30795 3415 30837 3424
rect 31210 3464 31268 3465
rect 31210 3424 31219 3464
rect 31259 3424 31268 3464
rect 31210 3423 31268 3424
rect 31659 3464 31701 3473
rect 31659 3424 31660 3464
rect 31700 3424 31701 3464
rect 31659 3415 31701 3424
rect 32427 3464 32469 3473
rect 32427 3424 32428 3464
rect 32468 3424 32469 3464
rect 32427 3415 32469 3424
rect 32907 3464 32949 3473
rect 32907 3424 32908 3464
rect 32948 3424 32949 3464
rect 32907 3415 32949 3424
rect 33771 3464 33813 3473
rect 33771 3424 33772 3464
rect 33812 3424 33813 3464
rect 33771 3415 33813 3424
rect 35019 3464 35061 3473
rect 35019 3424 35020 3464
rect 35060 3424 35061 3464
rect 35019 3415 35061 3424
rect 35722 3464 35780 3465
rect 35722 3424 35731 3464
rect 35771 3424 35780 3464
rect 35722 3423 35780 3424
rect 36267 3464 36309 3473
rect 36267 3424 36268 3464
rect 36308 3424 36309 3464
rect 36267 3415 36309 3424
rect 36939 3464 36981 3473
rect 36939 3424 36940 3464
rect 36980 3424 36981 3464
rect 36939 3415 36981 3424
rect 37707 3464 37749 3473
rect 37707 3424 37708 3464
rect 37748 3424 37749 3464
rect 37707 3415 37749 3424
rect 41739 3464 41781 3473
rect 41739 3424 41740 3464
rect 41780 3424 41781 3464
rect 41739 3415 41781 3424
rect 42027 3464 42069 3473
rect 42027 3424 42028 3464
rect 42068 3424 42069 3464
rect 42027 3415 42069 3424
rect 42411 3464 42453 3473
rect 42411 3424 42412 3464
rect 42452 3424 42453 3464
rect 42411 3415 42453 3424
rect 42699 3464 42741 3473
rect 42699 3424 42700 3464
rect 42740 3424 42741 3464
rect 42699 3415 42741 3424
rect 42987 3464 43029 3473
rect 42987 3424 42988 3464
rect 43028 3424 43029 3464
rect 42987 3415 43029 3424
rect 43275 3464 43317 3473
rect 43275 3424 43276 3464
rect 43316 3424 43317 3464
rect 43275 3415 43317 3424
rect 43563 3464 43605 3473
rect 43563 3424 43564 3464
rect 43604 3424 43605 3464
rect 43563 3415 43605 3424
rect 43851 3464 43893 3473
rect 43851 3424 43852 3464
rect 43892 3424 43893 3464
rect 43851 3415 43893 3424
rect 44139 3464 44181 3473
rect 44139 3424 44140 3464
rect 44180 3424 44181 3464
rect 44139 3415 44181 3424
rect 44427 3464 44469 3473
rect 44427 3424 44428 3464
rect 44468 3424 44469 3464
rect 44427 3415 44469 3424
rect 44715 3464 44757 3473
rect 44715 3424 44716 3464
rect 44756 3424 44757 3464
rect 44715 3415 44757 3424
rect 51435 3464 51477 3473
rect 51435 3424 51436 3464
rect 51476 3424 51477 3464
rect 51435 3415 51477 3424
rect 51819 3464 51861 3473
rect 51819 3424 51820 3464
rect 51860 3424 51861 3464
rect 51819 3415 51861 3424
rect 31035 3296 31077 3305
rect 31035 3256 31036 3296
rect 31076 3256 31077 3296
rect 31035 3247 31077 3256
rect 31419 3296 31461 3305
rect 31419 3256 31420 3296
rect 31460 3256 31461 3296
rect 31419 3247 31461 3256
rect 42267 3296 42309 3305
rect 42267 3256 42268 3296
rect 42308 3256 42309 3296
rect 42267 3247 42309 3256
rect 49995 3296 50037 3305
rect 49995 3256 49996 3296
rect 50036 3256 50037 3296
rect 49995 3247 50037 3256
rect 50283 3296 50325 3305
rect 50283 3256 50284 3296
rect 50324 3256 50325 3296
rect 50283 3247 50325 3256
rect 50859 3296 50901 3305
rect 50859 3256 50860 3296
rect 50900 3256 50901 3296
rect 50859 3247 50901 3256
rect 14427 3212 14469 3221
rect 14427 3172 14428 3212
rect 14468 3172 14469 3212
rect 14427 3163 14469 3172
rect 14907 3212 14949 3221
rect 14907 3172 14908 3212
rect 14948 3172 14949 3212
rect 14907 3163 14949 3172
rect 17403 3212 17445 3221
rect 17403 3172 17404 3212
rect 17444 3172 17445 3212
rect 17403 3163 17445 3172
rect 21915 3212 21957 3221
rect 21915 3172 21916 3212
rect 21956 3172 21957 3212
rect 21915 3163 21957 3172
rect 28443 3212 28485 3221
rect 28443 3172 28444 3212
rect 28484 3172 28485 3212
rect 28443 3163 28485 3172
rect 29883 3212 29925 3221
rect 29883 3172 29884 3212
rect 29924 3172 29925 3212
rect 29883 3163 29925 3172
rect 30651 3212 30693 3221
rect 30651 3172 30652 3212
rect 30692 3172 30693 3212
rect 30651 3163 30693 3172
rect 31899 3212 31941 3221
rect 31899 3172 31900 3212
rect 31940 3172 31941 3212
rect 31899 3163 31941 3172
rect 32667 3212 32709 3221
rect 32667 3172 32668 3212
rect 32708 3172 32709 3212
rect 32667 3163 32709 3172
rect 33147 3212 33189 3221
rect 33147 3172 33148 3212
rect 33188 3172 33189 3212
rect 33147 3163 33189 3172
rect 34011 3212 34053 3221
rect 34011 3172 34012 3212
rect 34052 3172 34053 3212
rect 34011 3163 34053 3172
rect 35259 3212 35301 3221
rect 35259 3172 35260 3212
rect 35300 3172 35301 3212
rect 35259 3163 35301 3172
rect 35547 3212 35589 3221
rect 35547 3172 35548 3212
rect 35588 3172 35589 3212
rect 35547 3163 35589 3172
rect 36027 3212 36069 3221
rect 36027 3172 36028 3212
rect 36068 3172 36069 3212
rect 36027 3163 36069 3172
rect 36699 3212 36741 3221
rect 36699 3172 36700 3212
rect 36740 3172 36741 3212
rect 36699 3163 36741 3172
rect 37467 3212 37509 3221
rect 37467 3172 37468 3212
rect 37508 3172 37509 3212
rect 37467 3163 37509 3172
rect 41722 3212 41780 3213
rect 41722 3172 41731 3212
rect 41771 3172 41780 3212
rect 41722 3171 41780 3172
rect 50554 3212 50612 3213
rect 50554 3172 50563 3212
rect 50603 3172 50612 3212
rect 50554 3171 50612 3172
rect 51226 3212 51284 3213
rect 51226 3172 51235 3212
rect 51275 3172 51284 3212
rect 51226 3171 51284 3172
rect 51675 3212 51717 3221
rect 51675 3172 51676 3212
rect 51716 3172 51717 3212
rect 51675 3163 51717 3172
rect 1152 3044 52128 3068
rect 1152 3004 4928 3044
rect 4968 3004 5010 3044
rect 5050 3004 5092 3044
rect 5132 3004 5174 3044
rect 5214 3004 5256 3044
rect 5296 3004 20048 3044
rect 20088 3004 20130 3044
rect 20170 3004 20212 3044
rect 20252 3004 20294 3044
rect 20334 3004 20376 3044
rect 20416 3004 35168 3044
rect 35208 3004 35250 3044
rect 35290 3004 35332 3044
rect 35372 3004 35414 3044
rect 35454 3004 35496 3044
rect 35536 3004 50288 3044
rect 50328 3004 50370 3044
rect 50410 3004 50452 3044
rect 50492 3004 50534 3044
rect 50574 3004 50616 3044
rect 50656 3004 52128 3044
rect 1152 2980 52128 3004
rect 14331 2876 14373 2885
rect 14331 2836 14332 2876
rect 14372 2836 14373 2876
rect 14331 2827 14373 2836
rect 23259 2876 23301 2885
rect 23259 2836 23260 2876
rect 23300 2836 23301 2876
rect 23259 2827 23301 2836
rect 49978 2876 50036 2877
rect 49978 2836 49987 2876
rect 50027 2836 50036 2876
rect 49978 2835 50036 2836
rect 18459 2792 18501 2801
rect 18459 2752 18460 2792
rect 18500 2752 18501 2792
rect 18459 2743 18501 2752
rect 20763 2792 20805 2801
rect 20763 2752 20764 2792
rect 20804 2752 20805 2792
rect 20763 2743 20805 2752
rect 23739 2792 23781 2801
rect 23739 2752 23740 2792
rect 23780 2752 23781 2792
rect 23739 2743 23781 2752
rect 52059 2792 52101 2801
rect 52059 2752 52060 2792
rect 52100 2752 52101 2792
rect 52059 2743 52101 2752
rect 2187 2624 2229 2633
rect 2187 2584 2188 2624
rect 2228 2584 2229 2624
rect 2187 2575 2229 2584
rect 7275 2624 7317 2633
rect 7275 2584 7276 2624
rect 7316 2584 7317 2624
rect 7275 2575 7317 2584
rect 11787 2624 11829 2633
rect 11787 2584 11788 2624
rect 11828 2584 11829 2624
rect 11787 2575 11829 2584
rect 13131 2624 13173 2633
rect 13131 2584 13132 2624
rect 13172 2584 13173 2624
rect 13131 2575 13173 2584
rect 14091 2624 14133 2633
rect 14091 2584 14092 2624
rect 14132 2584 14133 2624
rect 14091 2575 14133 2584
rect 14667 2624 14709 2633
rect 14667 2584 14668 2624
rect 14708 2584 14709 2624
rect 14667 2575 14709 2584
rect 18219 2624 18261 2633
rect 18219 2584 18220 2624
rect 18260 2584 18261 2624
rect 18219 2575 18261 2584
rect 18603 2624 18645 2633
rect 18603 2584 18604 2624
rect 18644 2584 18645 2624
rect 18603 2575 18645 2584
rect 20523 2624 20565 2633
rect 20523 2584 20524 2624
rect 20564 2584 20565 2624
rect 20523 2575 20565 2584
rect 20907 2624 20949 2633
rect 20907 2584 20908 2624
rect 20948 2584 20949 2624
rect 20907 2575 20949 2584
rect 23019 2624 23061 2633
rect 23019 2584 23020 2624
rect 23060 2584 23061 2624
rect 23019 2575 23061 2584
rect 23499 2624 23541 2633
rect 23499 2584 23500 2624
rect 23540 2584 23541 2624
rect 23499 2575 23541 2584
rect 24075 2624 24117 2633
rect 24075 2584 24076 2624
rect 24116 2584 24117 2624
rect 24075 2575 24117 2584
rect 24555 2624 24597 2633
rect 24555 2584 24556 2624
rect 24596 2584 24597 2624
rect 24555 2575 24597 2584
rect 24795 2624 24837 2633
rect 24795 2584 24796 2624
rect 24836 2584 24837 2624
rect 24795 2575 24837 2584
rect 24939 2624 24981 2633
rect 24939 2584 24940 2624
rect 24980 2584 24981 2624
rect 24939 2575 24981 2584
rect 25611 2624 25653 2633
rect 25611 2584 25612 2624
rect 25652 2584 25653 2624
rect 25611 2575 25653 2584
rect 27051 2624 27093 2633
rect 27051 2584 27052 2624
rect 27092 2584 27093 2624
rect 27051 2575 27093 2584
rect 28395 2624 28437 2633
rect 28395 2584 28396 2624
rect 28436 2584 28437 2624
rect 28395 2575 28437 2584
rect 28779 2624 28821 2633
rect 28779 2584 28780 2624
rect 28820 2584 28821 2624
rect 28779 2575 28821 2584
rect 33387 2624 33429 2633
rect 33387 2584 33388 2624
rect 33428 2584 33429 2624
rect 33387 2575 33429 2584
rect 34251 2624 34293 2633
rect 34251 2584 34252 2624
rect 34292 2584 34293 2624
rect 34251 2575 34293 2584
rect 34635 2624 34677 2633
rect 34635 2584 34636 2624
rect 34676 2584 34677 2624
rect 34635 2575 34677 2584
rect 39531 2624 39573 2633
rect 39531 2584 39532 2624
rect 39572 2584 39573 2624
rect 39531 2575 39573 2584
rect 40011 2624 40053 2633
rect 40011 2584 40012 2624
rect 40052 2584 40053 2624
rect 40011 2575 40053 2584
rect 49035 2624 49077 2633
rect 49035 2584 49036 2624
rect 49076 2584 49077 2624
rect 49035 2575 49077 2584
rect 49323 2624 49365 2633
rect 49323 2584 49324 2624
rect 49364 2584 49365 2624
rect 49323 2575 49365 2584
rect 49611 2624 49653 2633
rect 49611 2584 49612 2624
rect 49652 2584 49653 2624
rect 49611 2575 49653 2584
rect 49899 2624 49941 2633
rect 49899 2584 49900 2624
rect 49940 2584 49941 2624
rect 49899 2575 49941 2584
rect 50187 2624 50229 2633
rect 50187 2584 50188 2624
rect 50228 2584 50229 2624
rect 50187 2575 50229 2584
rect 50475 2624 50517 2633
rect 50475 2584 50476 2624
rect 50516 2584 50517 2624
rect 50475 2575 50517 2584
rect 50763 2624 50805 2633
rect 50763 2584 50764 2624
rect 50804 2584 50805 2624
rect 50763 2575 50805 2584
rect 51051 2624 51093 2633
rect 51051 2584 51052 2624
rect 51092 2584 51093 2624
rect 51051 2575 51093 2584
rect 51435 2624 51477 2633
rect 51435 2584 51436 2624
rect 51476 2584 51477 2624
rect 51435 2575 51477 2584
rect 51819 2624 51861 2633
rect 51819 2584 51820 2624
rect 51860 2584 51861 2624
rect 51819 2575 51861 2584
rect 7515 2540 7557 2549
rect 7515 2500 7516 2540
rect 7556 2500 7557 2540
rect 7515 2491 7557 2500
rect 51675 2540 51717 2549
rect 51675 2500 51676 2540
rect 51716 2500 51717 2540
rect 51675 2491 51717 2500
rect 2427 2456 2469 2465
rect 2427 2416 2428 2456
rect 2468 2416 2469 2456
rect 2427 2407 2469 2416
rect 12027 2456 12069 2465
rect 12027 2416 12028 2456
rect 12068 2416 12069 2456
rect 12027 2407 12069 2416
rect 13371 2456 13413 2465
rect 13371 2416 13372 2456
rect 13412 2416 13413 2456
rect 13371 2407 13413 2416
rect 14907 2456 14949 2465
rect 14907 2416 14908 2456
rect 14948 2416 14949 2456
rect 14907 2407 14949 2416
rect 18843 2456 18885 2465
rect 18843 2416 18844 2456
rect 18884 2416 18885 2456
rect 18843 2407 18885 2416
rect 21147 2456 21189 2465
rect 21147 2416 21148 2456
rect 21188 2416 21189 2456
rect 21147 2407 21189 2416
rect 24315 2456 24357 2465
rect 24315 2416 24316 2456
rect 24356 2416 24357 2456
rect 24315 2407 24357 2416
rect 25179 2456 25221 2465
rect 25179 2416 25180 2456
rect 25220 2416 25221 2456
rect 25179 2407 25221 2416
rect 25851 2456 25893 2465
rect 25851 2416 25852 2456
rect 25892 2416 25893 2456
rect 25851 2407 25893 2416
rect 27291 2456 27333 2465
rect 27291 2416 27292 2456
rect 27332 2416 27333 2456
rect 27291 2407 27333 2416
rect 28635 2456 28677 2465
rect 28635 2416 28636 2456
rect 28676 2416 28677 2456
rect 28635 2407 28677 2416
rect 29019 2456 29061 2465
rect 29019 2416 29020 2456
rect 29060 2416 29061 2456
rect 29019 2407 29061 2416
rect 33627 2456 33669 2465
rect 33627 2416 33628 2456
rect 33668 2416 33669 2456
rect 33627 2407 33669 2416
rect 34491 2456 34533 2465
rect 34491 2416 34492 2456
rect 34532 2416 34533 2456
rect 34491 2407 34533 2416
rect 34875 2456 34917 2465
rect 34875 2416 34876 2456
rect 34916 2416 34917 2456
rect 34875 2407 34917 2416
rect 39291 2456 39333 2465
rect 39291 2416 39292 2456
rect 39332 2416 39333 2456
rect 39291 2407 39333 2416
rect 39771 2456 39813 2465
rect 39771 2416 39772 2456
rect 39812 2416 39813 2456
rect 39771 2407 39813 2416
rect 51291 2456 51333 2465
rect 51291 2416 51292 2456
rect 51332 2416 51333 2456
rect 51291 2407 51333 2416
rect 1152 2288 52128 2312
rect 1152 2248 3688 2288
rect 3728 2248 3770 2288
rect 3810 2248 3852 2288
rect 3892 2248 3934 2288
rect 3974 2248 4016 2288
rect 4056 2248 18808 2288
rect 18848 2248 18890 2288
rect 18930 2248 18972 2288
rect 19012 2248 19054 2288
rect 19094 2248 19136 2288
rect 19176 2248 33928 2288
rect 33968 2248 34010 2288
rect 34050 2248 34092 2288
rect 34132 2248 34174 2288
rect 34214 2248 34256 2288
rect 34296 2248 49048 2288
rect 49088 2248 49130 2288
rect 49170 2248 49212 2288
rect 49252 2248 49294 2288
rect 49334 2248 49376 2288
rect 49416 2248 52128 2288
rect 1152 2224 52128 2248
rect 52059 2120 52101 2129
rect 52059 2080 52060 2120
rect 52100 2080 52101 2120
rect 52059 2071 52101 2080
rect 23019 1952 23061 1961
rect 23019 1912 23020 1952
rect 23060 1912 23061 1952
rect 23019 1903 23061 1912
rect 23403 1952 23445 1961
rect 23403 1912 23404 1952
rect 23444 1912 23445 1952
rect 23403 1903 23445 1912
rect 23787 1952 23829 1961
rect 23787 1912 23788 1952
rect 23828 1912 23829 1952
rect 23787 1903 23829 1912
rect 24171 1952 24213 1961
rect 24171 1912 24172 1952
rect 24212 1912 24213 1952
rect 24171 1903 24213 1912
rect 24555 1952 24597 1961
rect 24555 1912 24556 1952
rect 24596 1912 24597 1952
rect 24555 1903 24597 1912
rect 24939 1952 24981 1961
rect 24939 1912 24940 1952
rect 24980 1912 24981 1952
rect 24939 1903 24981 1912
rect 25323 1952 25365 1961
rect 25323 1912 25324 1952
rect 25364 1912 25365 1952
rect 25323 1903 25365 1912
rect 25707 1952 25749 1961
rect 25707 1912 25708 1952
rect 25748 1912 25749 1952
rect 25707 1903 25749 1912
rect 26091 1952 26133 1961
rect 26091 1912 26092 1952
rect 26132 1912 26133 1952
rect 26091 1903 26133 1912
rect 26475 1952 26517 1961
rect 26475 1912 26476 1952
rect 26516 1912 26517 1952
rect 26475 1903 26517 1912
rect 26859 1952 26901 1961
rect 26859 1912 26860 1952
rect 26900 1912 26901 1952
rect 26859 1903 26901 1912
rect 27243 1952 27285 1961
rect 27243 1912 27244 1952
rect 27284 1912 27285 1952
rect 27243 1903 27285 1912
rect 27627 1952 27669 1961
rect 27627 1912 27628 1952
rect 27668 1912 27669 1952
rect 27627 1903 27669 1912
rect 28011 1952 28053 1961
rect 28011 1912 28012 1952
rect 28052 1912 28053 1952
rect 28011 1903 28053 1912
rect 28395 1952 28437 1961
rect 28395 1912 28396 1952
rect 28436 1912 28437 1952
rect 28395 1903 28437 1912
rect 28827 1952 28869 1961
rect 28827 1912 28828 1952
rect 28868 1912 28869 1952
rect 28827 1903 28869 1912
rect 29163 1952 29205 1961
rect 29163 1912 29164 1952
rect 29204 1912 29205 1952
rect 29163 1903 29205 1912
rect 29547 1952 29589 1961
rect 29547 1912 29548 1952
rect 29588 1912 29589 1952
rect 29547 1903 29589 1912
rect 29931 1952 29973 1961
rect 29931 1912 29932 1952
rect 29972 1912 29973 1952
rect 29931 1903 29973 1912
rect 30315 1952 30357 1961
rect 30315 1912 30316 1952
rect 30356 1912 30357 1952
rect 30315 1903 30357 1912
rect 30699 1952 30741 1961
rect 30699 1912 30700 1952
rect 30740 1912 30741 1952
rect 30699 1903 30741 1912
rect 31083 1952 31125 1961
rect 31083 1912 31084 1952
rect 31124 1912 31125 1952
rect 31083 1903 31125 1912
rect 31467 1952 31509 1961
rect 31467 1912 31468 1952
rect 31508 1912 31509 1952
rect 31467 1903 31509 1912
rect 31851 1952 31893 1961
rect 31851 1912 31852 1952
rect 31892 1912 31893 1952
rect 31851 1903 31893 1912
rect 32235 1952 32277 1961
rect 32235 1912 32236 1952
rect 32276 1912 32277 1952
rect 32235 1903 32277 1912
rect 32619 1952 32661 1961
rect 32619 1912 32620 1952
rect 32660 1912 32661 1952
rect 32619 1903 32661 1912
rect 33003 1952 33045 1961
rect 33003 1912 33004 1952
rect 33044 1912 33045 1952
rect 33003 1903 33045 1912
rect 33387 1952 33429 1961
rect 33387 1912 33388 1952
rect 33428 1912 33429 1952
rect 33387 1903 33429 1912
rect 33771 1952 33813 1961
rect 33771 1912 33772 1952
rect 33812 1912 33813 1952
rect 33771 1903 33813 1912
rect 34155 1952 34197 1961
rect 34155 1912 34156 1952
rect 34196 1912 34197 1952
rect 34155 1903 34197 1912
rect 34474 1952 34532 1953
rect 34474 1912 34483 1952
rect 34523 1912 34532 1952
rect 34474 1911 34532 1912
rect 34858 1952 34916 1953
rect 34858 1912 34867 1952
rect 34907 1912 34916 1952
rect 34858 1911 34916 1912
rect 35307 1952 35349 1961
rect 35307 1912 35308 1952
rect 35348 1912 35349 1952
rect 35307 1903 35349 1912
rect 35691 1952 35733 1961
rect 35691 1912 35692 1952
rect 35732 1912 35733 1952
rect 35691 1903 35733 1912
rect 36075 1952 36117 1961
rect 36075 1912 36076 1952
rect 36116 1912 36117 1952
rect 36075 1903 36117 1912
rect 36459 1952 36501 1961
rect 36459 1912 36460 1952
rect 36500 1912 36501 1952
rect 36459 1903 36501 1912
rect 36843 1952 36885 1961
rect 36843 1912 36844 1952
rect 36884 1912 36885 1952
rect 36843 1903 36885 1912
rect 37227 1952 37269 1961
rect 37227 1912 37228 1952
rect 37268 1912 37269 1952
rect 37227 1903 37269 1912
rect 37611 1952 37653 1961
rect 37611 1912 37612 1952
rect 37652 1912 37653 1952
rect 37611 1903 37653 1912
rect 37995 1952 38037 1961
rect 37995 1912 37996 1952
rect 38036 1912 38037 1952
rect 37995 1903 38037 1912
rect 38379 1952 38421 1961
rect 38379 1912 38380 1952
rect 38420 1912 38421 1952
rect 38379 1903 38421 1912
rect 38763 1952 38805 1961
rect 38763 1912 38764 1952
rect 38804 1912 38805 1952
rect 38763 1903 38805 1912
rect 39147 1952 39189 1961
rect 39147 1912 39148 1952
rect 39188 1912 39189 1952
rect 39147 1903 39189 1912
rect 39531 1952 39573 1961
rect 39531 1912 39532 1952
rect 39572 1912 39573 1952
rect 39531 1903 39573 1912
rect 39915 1952 39957 1961
rect 39915 1912 39916 1952
rect 39956 1912 39957 1952
rect 39915 1903 39957 1912
rect 40299 1952 40341 1961
rect 40299 1912 40300 1952
rect 40340 1912 40341 1952
rect 40299 1903 40341 1912
rect 40683 1952 40725 1961
rect 40683 1912 40684 1952
rect 40724 1912 40725 1952
rect 40683 1903 40725 1912
rect 41067 1952 41109 1961
rect 41067 1912 41068 1952
rect 41108 1912 41109 1952
rect 41067 1903 41109 1912
rect 41451 1952 41493 1961
rect 41451 1912 41452 1952
rect 41492 1912 41493 1952
rect 41451 1903 41493 1912
rect 41835 1952 41877 1961
rect 41835 1912 41836 1952
rect 41876 1912 41877 1952
rect 41835 1903 41877 1912
rect 42219 1952 42261 1961
rect 42219 1912 42220 1952
rect 42260 1912 42261 1952
rect 42219 1903 42261 1912
rect 42603 1952 42645 1961
rect 42603 1912 42604 1952
rect 42644 1912 42645 1952
rect 42603 1903 42645 1912
rect 49995 1952 50037 1961
rect 49995 1912 49996 1952
rect 50036 1912 50037 1952
rect 49995 1903 50037 1912
rect 50379 1952 50421 1961
rect 50379 1912 50380 1952
rect 50420 1912 50421 1952
rect 50379 1903 50421 1912
rect 51051 1952 51093 1961
rect 51051 1912 51052 1952
rect 51092 1912 51093 1952
rect 51051 1903 51093 1912
rect 51627 1952 51669 1961
rect 51627 1912 51628 1952
rect 51668 1912 51669 1952
rect 51627 1903 51669 1912
rect 51819 1952 51861 1961
rect 51819 1912 51820 1952
rect 51860 1912 51861 1952
rect 51819 1903 51861 1912
rect 50859 1868 50901 1877
rect 50859 1828 50860 1868
rect 50900 1828 50901 1868
rect 50859 1819 50901 1828
rect 48651 1784 48693 1793
rect 48651 1744 48652 1784
rect 48692 1744 48693 1784
rect 48651 1735 48693 1744
rect 48939 1784 48981 1793
rect 48939 1744 48940 1784
rect 48980 1744 48981 1784
rect 48939 1735 48981 1744
rect 49227 1784 49269 1793
rect 49227 1744 49228 1784
rect 49268 1744 49269 1784
rect 49227 1735 49269 1744
rect 49515 1784 49557 1793
rect 49515 1744 49516 1784
rect 49556 1744 49557 1784
rect 49515 1735 49557 1744
rect 49803 1784 49845 1793
rect 49803 1744 49804 1784
rect 49844 1744 49845 1784
rect 49803 1735 49845 1744
rect 50235 1784 50277 1793
rect 50235 1744 50236 1784
rect 50276 1744 50277 1784
rect 50235 1735 50277 1744
rect 51291 1784 51333 1793
rect 51291 1744 51292 1784
rect 51332 1744 51333 1784
rect 51291 1735 51333 1744
rect 22779 1700 22821 1709
rect 22779 1660 22780 1700
rect 22820 1660 22821 1700
rect 22779 1651 22821 1660
rect 23163 1700 23205 1709
rect 23163 1660 23164 1700
rect 23204 1660 23205 1700
rect 23163 1651 23205 1660
rect 23547 1700 23589 1709
rect 23547 1660 23548 1700
rect 23588 1660 23589 1700
rect 23547 1651 23589 1660
rect 23931 1700 23973 1709
rect 23931 1660 23932 1700
rect 23972 1660 23973 1700
rect 23931 1651 23973 1660
rect 24315 1700 24357 1709
rect 24315 1660 24316 1700
rect 24356 1660 24357 1700
rect 24315 1651 24357 1660
rect 24699 1700 24741 1709
rect 24699 1660 24700 1700
rect 24740 1660 24741 1700
rect 24699 1651 24741 1660
rect 25083 1700 25125 1709
rect 25083 1660 25084 1700
rect 25124 1660 25125 1700
rect 25083 1651 25125 1660
rect 25467 1700 25509 1709
rect 25467 1660 25468 1700
rect 25508 1660 25509 1700
rect 25467 1651 25509 1660
rect 25851 1700 25893 1709
rect 25851 1660 25852 1700
rect 25892 1660 25893 1700
rect 25851 1651 25893 1660
rect 26235 1700 26277 1709
rect 26235 1660 26236 1700
rect 26276 1660 26277 1700
rect 26235 1651 26277 1660
rect 26619 1700 26661 1709
rect 26619 1660 26620 1700
rect 26660 1660 26661 1700
rect 26619 1651 26661 1660
rect 27003 1700 27045 1709
rect 27003 1660 27004 1700
rect 27044 1660 27045 1700
rect 27003 1651 27045 1660
rect 27387 1700 27429 1709
rect 27387 1660 27388 1700
rect 27428 1660 27429 1700
rect 27387 1651 27429 1660
rect 27771 1700 27813 1709
rect 27771 1660 27772 1700
rect 27812 1660 27813 1700
rect 27771 1651 27813 1660
rect 28155 1700 28197 1709
rect 28155 1660 28156 1700
rect 28196 1660 28197 1700
rect 28155 1651 28197 1660
rect 28539 1700 28581 1709
rect 28539 1660 28540 1700
rect 28580 1660 28581 1700
rect 28539 1651 28581 1660
rect 28923 1700 28965 1709
rect 28923 1660 28924 1700
rect 28964 1660 28965 1700
rect 28923 1651 28965 1660
rect 29307 1700 29349 1709
rect 29307 1660 29308 1700
rect 29348 1660 29349 1700
rect 29307 1651 29349 1660
rect 29691 1700 29733 1709
rect 29691 1660 29692 1700
rect 29732 1660 29733 1700
rect 29691 1651 29733 1660
rect 30075 1700 30117 1709
rect 30075 1660 30076 1700
rect 30116 1660 30117 1700
rect 30075 1651 30117 1660
rect 30459 1700 30501 1709
rect 30459 1660 30460 1700
rect 30500 1660 30501 1700
rect 30459 1651 30501 1660
rect 30843 1700 30885 1709
rect 30843 1660 30844 1700
rect 30884 1660 30885 1700
rect 30843 1651 30885 1660
rect 31227 1700 31269 1709
rect 31227 1660 31228 1700
rect 31268 1660 31269 1700
rect 31227 1651 31269 1660
rect 31611 1700 31653 1709
rect 31611 1660 31612 1700
rect 31652 1660 31653 1700
rect 31611 1651 31653 1660
rect 31995 1700 32037 1709
rect 31995 1660 31996 1700
rect 32036 1660 32037 1700
rect 31995 1651 32037 1660
rect 32379 1700 32421 1709
rect 32379 1660 32380 1700
rect 32420 1660 32421 1700
rect 32379 1651 32421 1660
rect 32763 1700 32805 1709
rect 32763 1660 32764 1700
rect 32804 1660 32805 1700
rect 32763 1651 32805 1660
rect 33147 1700 33189 1709
rect 33147 1660 33148 1700
rect 33188 1660 33189 1700
rect 33147 1651 33189 1660
rect 33531 1700 33573 1709
rect 33531 1660 33532 1700
rect 33572 1660 33573 1700
rect 33531 1651 33573 1660
rect 33915 1700 33957 1709
rect 33915 1660 33916 1700
rect 33956 1660 33957 1700
rect 33915 1651 33957 1660
rect 34299 1700 34341 1709
rect 34299 1660 34300 1700
rect 34340 1660 34341 1700
rect 34299 1651 34341 1660
rect 34683 1700 34725 1709
rect 34683 1660 34684 1700
rect 34724 1660 34725 1700
rect 34683 1651 34725 1660
rect 35067 1700 35109 1709
rect 35067 1660 35068 1700
rect 35108 1660 35109 1700
rect 35067 1651 35109 1660
rect 35451 1700 35493 1709
rect 35451 1660 35452 1700
rect 35492 1660 35493 1700
rect 35451 1651 35493 1660
rect 35835 1700 35877 1709
rect 35835 1660 35836 1700
rect 35876 1660 35877 1700
rect 35835 1651 35877 1660
rect 36219 1700 36261 1709
rect 36219 1660 36220 1700
rect 36260 1660 36261 1700
rect 36219 1651 36261 1660
rect 36603 1700 36645 1709
rect 36603 1660 36604 1700
rect 36644 1660 36645 1700
rect 36603 1651 36645 1660
rect 36987 1700 37029 1709
rect 36987 1660 36988 1700
rect 37028 1660 37029 1700
rect 36987 1651 37029 1660
rect 37371 1700 37413 1709
rect 37371 1660 37372 1700
rect 37412 1660 37413 1700
rect 37371 1651 37413 1660
rect 37755 1700 37797 1709
rect 37755 1660 37756 1700
rect 37796 1660 37797 1700
rect 37755 1651 37797 1660
rect 38139 1700 38181 1709
rect 38139 1660 38140 1700
rect 38180 1660 38181 1700
rect 38139 1651 38181 1660
rect 38523 1700 38565 1709
rect 38523 1660 38524 1700
rect 38564 1660 38565 1700
rect 38523 1651 38565 1660
rect 38907 1700 38949 1709
rect 38907 1660 38908 1700
rect 38948 1660 38949 1700
rect 38907 1651 38949 1660
rect 39291 1700 39333 1709
rect 39291 1660 39292 1700
rect 39332 1660 39333 1700
rect 39291 1651 39333 1660
rect 39675 1700 39717 1709
rect 39675 1660 39676 1700
rect 39716 1660 39717 1700
rect 39675 1651 39717 1660
rect 40059 1700 40101 1709
rect 40059 1660 40060 1700
rect 40100 1660 40101 1700
rect 40059 1651 40101 1660
rect 40443 1700 40485 1709
rect 40443 1660 40444 1700
rect 40484 1660 40485 1700
rect 40443 1651 40485 1660
rect 40827 1700 40869 1709
rect 40827 1660 40828 1700
rect 40868 1660 40869 1700
rect 40827 1651 40869 1660
rect 41211 1700 41253 1709
rect 41211 1660 41212 1700
rect 41252 1660 41253 1700
rect 41211 1651 41253 1660
rect 41595 1700 41637 1709
rect 41595 1660 41596 1700
rect 41636 1660 41637 1700
rect 41595 1651 41637 1660
rect 41979 1700 42021 1709
rect 41979 1660 41980 1700
rect 42020 1660 42021 1700
rect 41979 1651 42021 1660
rect 42363 1700 42405 1709
rect 42363 1660 42364 1700
rect 42404 1660 42405 1700
rect 42363 1651 42405 1660
rect 50619 1700 50661 1709
rect 50619 1660 50620 1700
rect 50660 1660 50661 1700
rect 50619 1651 50661 1660
rect 1152 1532 52128 1556
rect 1152 1492 4928 1532
rect 4968 1492 5010 1532
rect 5050 1492 5092 1532
rect 5132 1492 5174 1532
rect 5214 1492 5256 1532
rect 5296 1492 20048 1532
rect 20088 1492 20130 1532
rect 20170 1492 20212 1532
rect 20252 1492 20294 1532
rect 20334 1492 20376 1532
rect 20416 1492 35168 1532
rect 35208 1492 35250 1532
rect 35290 1492 35332 1532
rect 35372 1492 35414 1532
rect 35454 1492 35496 1532
rect 35536 1492 50288 1532
rect 50328 1492 50370 1532
rect 50410 1492 50452 1532
rect 50492 1492 50534 1532
rect 50574 1492 50616 1532
rect 50656 1492 52128 1532
rect 1152 1468 52128 1492
<< via1 >>
rect 4928 10564 4968 10604
rect 5010 10564 5050 10604
rect 5092 10564 5132 10604
rect 5174 10564 5214 10604
rect 5256 10564 5296 10604
rect 20048 10564 20088 10604
rect 20130 10564 20170 10604
rect 20212 10564 20252 10604
rect 20294 10564 20334 10604
rect 20376 10564 20416 10604
rect 35168 10564 35208 10604
rect 35250 10564 35290 10604
rect 35332 10564 35372 10604
rect 35414 10564 35454 10604
rect 35496 10564 35536 10604
rect 50288 10564 50328 10604
rect 50370 10564 50410 10604
rect 50452 10564 50492 10604
rect 50534 10564 50574 10604
rect 50616 10564 50656 10604
rect 1660 10396 1700 10436
rect 4156 10396 4196 10436
rect 6652 10396 6692 10436
rect 9148 10396 9188 10436
rect 11644 10396 11684 10436
rect 14140 10396 14180 10436
rect 16636 10396 16676 10436
rect 19132 10396 19172 10436
rect 21628 10396 21668 10436
rect 24124 10396 24164 10436
rect 26620 10396 26660 10436
rect 29116 10396 29156 10436
rect 31612 10396 31652 10436
rect 34108 10396 34148 10436
rect 39100 10396 39140 10436
rect 41596 10396 41636 10436
rect 44092 10396 44132 10436
rect 46588 10396 46628 10436
rect 49084 10396 49124 10436
rect 50524 10396 50564 10436
rect 50908 10396 50948 10436
rect 51772 10396 51812 10436
rect 51292 10312 51332 10352
rect 1900 10144 1940 10184
rect 4396 10144 4436 10184
rect 6892 10144 6932 10184
rect 9388 10144 9428 10184
rect 11884 10144 11924 10184
rect 14380 10144 14420 10184
rect 16876 10144 16916 10184
rect 19372 10144 19412 10184
rect 21868 10144 21908 10184
rect 24364 10144 24404 10184
rect 26860 10144 26900 10184
rect 29356 10144 29396 10184
rect 31852 10144 31892 10184
rect 34348 10144 34388 10184
rect 36604 10144 36644 10184
rect 36844 10144 36884 10184
rect 39340 10144 39380 10184
rect 41836 10144 41876 10184
rect 44332 10144 44372 10184
rect 46828 10144 46868 10184
rect 49324 10144 49364 10184
rect 49612 10144 49652 10184
rect 50092 10144 50132 10184
rect 50284 10144 50324 10184
rect 50668 10144 50708 10184
rect 51052 10144 51092 10184
rect 51436 10144 51476 10184
rect 52012 10144 52052 10184
rect 49852 10060 49892 10100
rect 51676 9976 51716 10016
rect 3688 9808 3728 9848
rect 3770 9808 3810 9848
rect 3852 9808 3892 9848
rect 3934 9808 3974 9848
rect 4016 9808 4056 9848
rect 18808 9808 18848 9848
rect 18890 9808 18930 9848
rect 18972 9808 19012 9848
rect 19054 9808 19094 9848
rect 19136 9808 19176 9848
rect 33928 9808 33968 9848
rect 34010 9808 34050 9848
rect 34092 9808 34132 9848
rect 34174 9808 34214 9848
rect 34256 9808 34296 9848
rect 49048 9808 49088 9848
rect 49130 9808 49170 9848
rect 49212 9808 49252 9848
rect 49294 9808 49334 9848
rect 49376 9808 49416 9848
rect 13852 9640 13892 9680
rect 15772 9640 15812 9680
rect 18460 9640 18500 9680
rect 20860 9640 20900 9680
rect 23164 9640 23204 9680
rect 24028 9640 24068 9680
rect 25372 9640 25412 9680
rect 26908 9640 26948 9680
rect 27868 9640 27908 9680
rect 29116 9640 29156 9680
rect 29692 9640 29732 9680
rect 41596 9640 41636 9680
rect 43420 9640 43460 9680
rect 43996 9640 44036 9680
rect 44956 9640 44996 9680
rect 46204 9640 46244 9680
rect 46684 9640 46724 9680
rect 48220 9640 48260 9680
rect 48892 9640 48932 9680
rect 50812 9640 50852 9680
rect 51196 9640 51236 9680
rect 40636 9556 40676 9596
rect 13708 9472 13748 9512
rect 14092 9472 14132 9512
rect 14284 9472 14324 9512
rect 14524 9472 14564 9512
rect 15628 9472 15668 9512
rect 16012 9472 16052 9512
rect 18700 9472 18740 9512
rect 21100 9472 21140 9512
rect 23404 9472 23444 9512
rect 23788 9472 23828 9512
rect 25612 9472 25652 9512
rect 26188 9472 26228 9512
rect 26668 9472 26708 9512
rect 28108 9472 28148 9512
rect 28876 9472 28916 9512
rect 29932 9472 29972 9512
rect 30220 9472 30260 9512
rect 30460 9472 30500 9512
rect 40300 9472 40340 9512
rect 40876 9472 40916 9512
rect 41836 9472 41876 9512
rect 42796 9472 42836 9512
rect 43660 9472 43700 9512
rect 44236 9472 44276 9512
rect 45196 9472 45236 9512
rect 46492 9472 46532 9512
rect 46924 9472 46964 9512
rect 47308 9472 47348 9512
rect 48460 9472 48500 9512
rect 48652 9472 48692 9512
rect 50572 9472 50612 9512
rect 50956 9472 50996 9512
rect 51436 9472 51476 9512
rect 51820 9472 51860 9512
rect 40060 9304 40100 9344
rect 15619 9220 15659 9260
rect 26428 9220 26468 9260
rect 42556 9220 42596 9260
rect 47068 9220 47108 9260
rect 50275 9220 50315 9260
rect 51676 9220 51716 9260
rect 52060 9220 52100 9260
rect 4928 9052 4968 9092
rect 5010 9052 5050 9092
rect 5092 9052 5132 9092
rect 5174 9052 5214 9092
rect 5256 9052 5296 9092
rect 20048 9052 20088 9092
rect 20130 9052 20170 9092
rect 20212 9052 20252 9092
rect 20294 9052 20334 9092
rect 20376 9052 20416 9092
rect 35168 9052 35208 9092
rect 35250 9052 35290 9092
rect 35332 9052 35372 9092
rect 35414 9052 35454 9092
rect 35496 9052 35536 9092
rect 50288 9052 50328 9092
rect 50370 9052 50410 9092
rect 50452 9052 50492 9092
rect 50534 9052 50574 9092
rect 50616 9052 50656 9092
rect 33724 8884 33764 8924
rect 25852 8800 25892 8840
rect 28348 8800 28388 8840
rect 25612 8632 25652 8672
rect 27724 8632 27764 8672
rect 27964 8632 28004 8672
rect 28108 8632 28148 8672
rect 33292 8632 33332 8672
rect 33484 8632 33524 8672
rect 33964 8632 34004 8672
rect 34252 8632 34292 8672
rect 34540 8632 34580 8672
rect 34828 8632 34868 8672
rect 35116 8632 35156 8672
rect 35404 8632 35444 8672
rect 35692 8632 35732 8672
rect 35884 8632 35924 8672
rect 51436 8632 51476 8672
rect 51676 8632 51716 8672
rect 51820 8632 51860 8672
rect 52060 8632 52100 8672
rect 3688 8296 3728 8336
rect 3770 8296 3810 8336
rect 3852 8296 3892 8336
rect 3934 8296 3974 8336
rect 4016 8296 4056 8336
rect 18808 8296 18848 8336
rect 18890 8296 18930 8336
rect 18972 8296 19012 8336
rect 19054 8296 19094 8336
rect 19136 8296 19176 8336
rect 33928 8296 33968 8336
rect 34010 8296 34050 8336
rect 34092 8296 34132 8336
rect 34174 8296 34214 8336
rect 34256 8296 34296 8336
rect 49048 8296 49088 8336
rect 49130 8296 49170 8336
rect 49212 8296 49252 8336
rect 49294 8296 49334 8336
rect 49376 8296 49416 8336
rect 23548 8128 23588 8168
rect 28252 8128 28292 8168
rect 31708 8044 31748 8084
rect 23308 7960 23348 8000
rect 28012 7960 28052 8000
rect 31468 7960 31508 8000
rect 35212 7960 35252 8000
rect 51436 7960 51476 8000
rect 51820 7960 51860 8000
rect 51676 7792 51716 7832
rect 33475 7708 33515 7748
rect 35452 7708 35492 7748
rect 52060 7708 52100 7748
rect 4928 7540 4968 7580
rect 5010 7540 5050 7580
rect 5092 7540 5132 7580
rect 5174 7540 5214 7580
rect 5256 7540 5296 7580
rect 20048 7540 20088 7580
rect 20130 7540 20170 7580
rect 20212 7540 20252 7580
rect 20294 7540 20334 7580
rect 20376 7540 20416 7580
rect 35168 7540 35208 7580
rect 35250 7540 35290 7580
rect 35332 7540 35372 7580
rect 35414 7540 35454 7580
rect 35496 7540 35536 7580
rect 50288 7540 50328 7580
rect 50370 7540 50410 7580
rect 50452 7540 50492 7580
rect 50534 7540 50574 7580
rect 50616 7540 50656 7580
rect 35212 7288 35252 7328
rect 35500 7288 35540 7328
rect 18892 7120 18932 7160
rect 23596 7120 23636 7160
rect 23836 7120 23876 7160
rect 29740 7120 29780 7160
rect 30220 7120 30260 7160
rect 51436 7120 51476 7160
rect 51820 7120 51860 7160
rect 52060 7120 52100 7160
rect 30460 7036 30500 7076
rect 19132 6952 19172 6992
rect 29980 6952 30020 6992
rect 51676 6952 51716 6992
rect 3688 6784 3728 6824
rect 3770 6784 3810 6824
rect 3852 6784 3892 6824
rect 3934 6784 3974 6824
rect 4016 6784 4056 6824
rect 18808 6784 18848 6824
rect 18890 6784 18930 6824
rect 18972 6784 19012 6824
rect 19054 6784 19094 6824
rect 19136 6784 19176 6824
rect 33928 6784 33968 6824
rect 34010 6784 34050 6824
rect 34092 6784 34132 6824
rect 34174 6784 34214 6824
rect 34256 6784 34296 6824
rect 49048 6784 49088 6824
rect 49130 6784 49170 6824
rect 49212 6784 49252 6824
rect 49294 6784 49334 6824
rect 49376 6784 49416 6824
rect 25660 6532 25700 6572
rect 22732 6448 22772 6488
rect 25420 6448 25460 6488
rect 25804 6448 25844 6488
rect 35500 6448 35540 6488
rect 35788 6448 35828 6488
rect 36172 6448 36212 6488
rect 36460 6448 36500 6488
rect 36748 6448 36788 6488
rect 37036 6448 37076 6488
rect 37324 6448 37364 6488
rect 37612 6448 37652 6488
rect 37900 6448 37940 6488
rect 38284 6448 38324 6488
rect 51436 6448 51476 6488
rect 51820 6448 51860 6488
rect 52060 6448 52100 6488
rect 26044 6280 26084 6320
rect 22972 6196 23012 6236
rect 36028 6196 36068 6236
rect 38524 6196 38564 6236
rect 51676 6196 51716 6236
rect 4928 6028 4968 6068
rect 5010 6028 5050 6068
rect 5092 6028 5132 6068
rect 5174 6028 5214 6068
rect 5256 6028 5296 6068
rect 20048 6028 20088 6068
rect 20130 6028 20170 6068
rect 20212 6028 20252 6068
rect 20294 6028 20334 6068
rect 20376 6028 20416 6068
rect 35168 6028 35208 6068
rect 35250 6028 35290 6068
rect 35332 6028 35372 6068
rect 35414 6028 35454 6068
rect 35496 6028 35536 6068
rect 50288 6028 50328 6068
rect 50370 6028 50410 6068
rect 50452 6028 50492 6068
rect 50534 6028 50574 6068
rect 50616 6028 50656 6068
rect 35788 5776 35828 5816
rect 36076 5776 36116 5816
rect 52060 5776 52100 5816
rect 23884 5608 23924 5648
rect 24124 5608 24164 5648
rect 27820 5608 27860 5648
rect 51436 5608 51476 5648
rect 51820 5608 51860 5648
rect 51676 5524 51716 5564
rect 28060 5440 28100 5480
rect 3688 5272 3728 5312
rect 3770 5272 3810 5312
rect 3852 5272 3892 5312
rect 3934 5272 3974 5312
rect 4016 5272 4056 5312
rect 18808 5272 18848 5312
rect 18890 5272 18930 5312
rect 18972 5272 19012 5312
rect 19054 5272 19094 5312
rect 19136 5272 19176 5312
rect 33928 5272 33968 5312
rect 34010 5272 34050 5312
rect 34092 5272 34132 5312
rect 34174 5272 34214 5312
rect 34256 5272 34296 5312
rect 49048 5272 49088 5312
rect 49130 5272 49170 5312
rect 49212 5272 49252 5312
rect 49294 5272 49334 5312
rect 49376 5272 49416 5312
rect 52060 5104 52100 5144
rect 14668 4936 14708 4976
rect 15244 4936 15284 4976
rect 24172 4936 24212 4976
rect 24844 4936 24884 4976
rect 25228 4936 25268 4976
rect 30028 4936 30068 4976
rect 51436 4936 51476 4976
rect 51820 4936 51860 4976
rect 30268 4768 30308 4808
rect 51676 4768 51716 4808
rect 14908 4684 14948 4724
rect 15484 4684 15524 4724
rect 24412 4684 24452 4724
rect 25084 4684 25124 4724
rect 25468 4684 25508 4724
rect 4928 4516 4968 4556
rect 5010 4516 5050 4556
rect 5092 4516 5132 4556
rect 5174 4516 5214 4556
rect 5256 4516 5296 4556
rect 20048 4516 20088 4556
rect 20130 4516 20170 4556
rect 20212 4516 20252 4556
rect 20294 4516 20334 4556
rect 20376 4516 20416 4556
rect 35168 4516 35208 4556
rect 35250 4516 35290 4556
rect 35332 4516 35372 4556
rect 35414 4516 35454 4556
rect 35496 4516 35536 4556
rect 50288 4516 50328 4556
rect 50370 4516 50410 4556
rect 50452 4516 50492 4556
rect 50534 4516 50574 4556
rect 50616 4516 50656 4556
rect 52060 4264 52100 4304
rect 13420 4096 13460 4136
rect 16396 4096 16436 4136
rect 16876 4096 16916 4136
rect 19180 4096 19220 4136
rect 23020 4096 23060 4136
rect 28012 4096 28052 4136
rect 38860 4096 38900 4136
rect 50860 4096 50900 4136
rect 51052 4096 51092 4136
rect 51436 4096 51476 4136
rect 51820 4096 51860 4136
rect 28252 4012 28292 4052
rect 51676 4012 51716 4052
rect 13660 3928 13700 3968
rect 16636 3928 16676 3968
rect 17116 3928 17156 3968
rect 19420 3928 19460 3968
rect 23260 3928 23300 3968
rect 38620 3928 38660 3968
rect 51292 3928 51332 3968
rect 3688 3760 3728 3800
rect 3770 3760 3810 3800
rect 3852 3760 3892 3800
rect 3934 3760 3974 3800
rect 4016 3760 4056 3800
rect 18808 3760 18848 3800
rect 18890 3760 18930 3800
rect 18972 3760 19012 3800
rect 19054 3760 19094 3800
rect 19136 3760 19176 3800
rect 33928 3760 33968 3800
rect 34010 3760 34050 3800
rect 34092 3760 34132 3800
rect 34174 3760 34214 3800
rect 34256 3760 34296 3800
rect 49048 3760 49088 3800
rect 49130 3760 49170 3800
rect 49212 3760 49252 3800
rect 49294 3760 49334 3800
rect 49376 3760 49416 3800
rect 22780 3592 22820 3632
rect 52060 3592 52100 3632
rect 19804 3508 19844 3548
rect 14188 3424 14228 3464
rect 14668 3424 14708 3464
rect 17116 3424 17156 3464
rect 19564 3424 19604 3464
rect 21292 3424 21332 3464
rect 21532 3424 21572 3464
rect 21715 3424 21755 3464
rect 22540 3424 22580 3464
rect 28204 3424 28244 3464
rect 29644 3424 29684 3464
rect 30412 3424 30452 3464
rect 30796 3424 30836 3464
rect 31219 3424 31259 3464
rect 31660 3424 31700 3464
rect 32428 3424 32468 3464
rect 32908 3424 32948 3464
rect 33772 3424 33812 3464
rect 35020 3424 35060 3464
rect 35731 3424 35771 3464
rect 36268 3424 36308 3464
rect 36940 3424 36980 3464
rect 37708 3424 37748 3464
rect 41740 3424 41780 3464
rect 42028 3424 42068 3464
rect 42412 3424 42452 3464
rect 42700 3424 42740 3464
rect 42988 3424 43028 3464
rect 43276 3424 43316 3464
rect 43564 3424 43604 3464
rect 43852 3424 43892 3464
rect 44140 3424 44180 3464
rect 44428 3424 44468 3464
rect 44716 3424 44756 3464
rect 51436 3424 51476 3464
rect 51820 3424 51860 3464
rect 31036 3256 31076 3296
rect 31420 3256 31460 3296
rect 42268 3256 42308 3296
rect 49996 3256 50036 3296
rect 50284 3256 50324 3296
rect 50860 3256 50900 3296
rect 14428 3172 14468 3212
rect 14908 3172 14948 3212
rect 17404 3172 17444 3212
rect 21916 3172 21956 3212
rect 28444 3172 28484 3212
rect 29884 3172 29924 3212
rect 30652 3172 30692 3212
rect 31900 3172 31940 3212
rect 32668 3172 32708 3212
rect 33148 3172 33188 3212
rect 34012 3172 34052 3212
rect 35260 3172 35300 3212
rect 35548 3172 35588 3212
rect 36028 3172 36068 3212
rect 36700 3172 36740 3212
rect 37468 3172 37508 3212
rect 41731 3172 41771 3212
rect 50563 3172 50603 3212
rect 51235 3172 51275 3212
rect 51676 3172 51716 3212
rect 4928 3004 4968 3044
rect 5010 3004 5050 3044
rect 5092 3004 5132 3044
rect 5174 3004 5214 3044
rect 5256 3004 5296 3044
rect 20048 3004 20088 3044
rect 20130 3004 20170 3044
rect 20212 3004 20252 3044
rect 20294 3004 20334 3044
rect 20376 3004 20416 3044
rect 35168 3004 35208 3044
rect 35250 3004 35290 3044
rect 35332 3004 35372 3044
rect 35414 3004 35454 3044
rect 35496 3004 35536 3044
rect 50288 3004 50328 3044
rect 50370 3004 50410 3044
rect 50452 3004 50492 3044
rect 50534 3004 50574 3044
rect 50616 3004 50656 3044
rect 14332 2836 14372 2876
rect 23260 2836 23300 2876
rect 49987 2836 50027 2876
rect 18460 2752 18500 2792
rect 20764 2752 20804 2792
rect 23740 2752 23780 2792
rect 52060 2752 52100 2792
rect 2188 2584 2228 2624
rect 7276 2584 7316 2624
rect 11788 2584 11828 2624
rect 13132 2584 13172 2624
rect 14092 2584 14132 2624
rect 14668 2584 14708 2624
rect 18220 2584 18260 2624
rect 18604 2584 18644 2624
rect 20524 2584 20564 2624
rect 20908 2584 20948 2624
rect 23020 2584 23060 2624
rect 23500 2584 23540 2624
rect 24076 2584 24116 2624
rect 24556 2584 24596 2624
rect 24796 2584 24836 2624
rect 24940 2584 24980 2624
rect 25612 2584 25652 2624
rect 27052 2584 27092 2624
rect 28396 2584 28436 2624
rect 28780 2584 28820 2624
rect 33388 2584 33428 2624
rect 34252 2584 34292 2624
rect 34636 2584 34676 2624
rect 39532 2584 39572 2624
rect 40012 2584 40052 2624
rect 49036 2584 49076 2624
rect 49324 2584 49364 2624
rect 49612 2584 49652 2624
rect 49900 2584 49940 2624
rect 50188 2584 50228 2624
rect 50476 2584 50516 2624
rect 50764 2584 50804 2624
rect 51052 2584 51092 2624
rect 51436 2584 51476 2624
rect 51820 2584 51860 2624
rect 7516 2500 7556 2540
rect 51676 2500 51716 2540
rect 2428 2416 2468 2456
rect 12028 2416 12068 2456
rect 13372 2416 13412 2456
rect 14908 2416 14948 2456
rect 18844 2416 18884 2456
rect 21148 2416 21188 2456
rect 24316 2416 24356 2456
rect 25180 2416 25220 2456
rect 25852 2416 25892 2456
rect 27292 2416 27332 2456
rect 28636 2416 28676 2456
rect 29020 2416 29060 2456
rect 33628 2416 33668 2456
rect 34492 2416 34532 2456
rect 34876 2416 34916 2456
rect 39292 2416 39332 2456
rect 39772 2416 39812 2456
rect 51292 2416 51332 2456
rect 3688 2248 3728 2288
rect 3770 2248 3810 2288
rect 3852 2248 3892 2288
rect 3934 2248 3974 2288
rect 4016 2248 4056 2288
rect 18808 2248 18848 2288
rect 18890 2248 18930 2288
rect 18972 2248 19012 2288
rect 19054 2248 19094 2288
rect 19136 2248 19176 2288
rect 33928 2248 33968 2288
rect 34010 2248 34050 2288
rect 34092 2248 34132 2288
rect 34174 2248 34214 2288
rect 34256 2248 34296 2288
rect 49048 2248 49088 2288
rect 49130 2248 49170 2288
rect 49212 2248 49252 2288
rect 49294 2248 49334 2288
rect 49376 2248 49416 2288
rect 52060 2080 52100 2120
rect 23020 1912 23060 1952
rect 23404 1912 23444 1952
rect 23788 1912 23828 1952
rect 24172 1912 24212 1952
rect 24556 1912 24596 1952
rect 24940 1912 24980 1952
rect 25324 1912 25364 1952
rect 25708 1912 25748 1952
rect 26092 1912 26132 1952
rect 26476 1912 26516 1952
rect 26860 1912 26900 1952
rect 27244 1912 27284 1952
rect 27628 1912 27668 1952
rect 28012 1912 28052 1952
rect 28396 1912 28436 1952
rect 28828 1912 28868 1952
rect 29164 1912 29204 1952
rect 29548 1912 29588 1952
rect 29932 1912 29972 1952
rect 30316 1912 30356 1952
rect 30700 1912 30740 1952
rect 31084 1912 31124 1952
rect 31468 1912 31508 1952
rect 31852 1912 31892 1952
rect 32236 1912 32276 1952
rect 32620 1912 32660 1952
rect 33004 1912 33044 1952
rect 33388 1912 33428 1952
rect 33772 1912 33812 1952
rect 34156 1912 34196 1952
rect 34483 1912 34523 1952
rect 34867 1912 34907 1952
rect 35308 1912 35348 1952
rect 35692 1912 35732 1952
rect 36076 1912 36116 1952
rect 36460 1912 36500 1952
rect 36844 1912 36884 1952
rect 37228 1912 37268 1952
rect 37612 1912 37652 1952
rect 37996 1912 38036 1952
rect 38380 1912 38420 1952
rect 38764 1912 38804 1952
rect 39148 1912 39188 1952
rect 39532 1912 39572 1952
rect 39916 1912 39956 1952
rect 40300 1912 40340 1952
rect 40684 1912 40724 1952
rect 41068 1912 41108 1952
rect 41452 1912 41492 1952
rect 41836 1912 41876 1952
rect 42220 1912 42260 1952
rect 42604 1912 42644 1952
rect 49996 1912 50036 1952
rect 50380 1912 50420 1952
rect 51052 1912 51092 1952
rect 51628 1912 51668 1952
rect 51820 1912 51860 1952
rect 50860 1828 50900 1868
rect 48652 1744 48692 1784
rect 48940 1744 48980 1784
rect 49228 1744 49268 1784
rect 49516 1744 49556 1784
rect 49804 1744 49844 1784
rect 50236 1744 50276 1784
rect 51292 1744 51332 1784
rect 22780 1660 22820 1700
rect 23164 1660 23204 1700
rect 23548 1660 23588 1700
rect 23932 1660 23972 1700
rect 24316 1660 24356 1700
rect 24700 1660 24740 1700
rect 25084 1660 25124 1700
rect 25468 1660 25508 1700
rect 25852 1660 25892 1700
rect 26236 1660 26276 1700
rect 26620 1660 26660 1700
rect 27004 1660 27044 1700
rect 27388 1660 27428 1700
rect 27772 1660 27812 1700
rect 28156 1660 28196 1700
rect 28540 1660 28580 1700
rect 28924 1660 28964 1700
rect 29308 1660 29348 1700
rect 29692 1660 29732 1700
rect 30076 1660 30116 1700
rect 30460 1660 30500 1700
rect 30844 1660 30884 1700
rect 31228 1660 31268 1700
rect 31612 1660 31652 1700
rect 31996 1660 32036 1700
rect 32380 1660 32420 1700
rect 32764 1660 32804 1700
rect 33148 1660 33188 1700
rect 33532 1660 33572 1700
rect 33916 1660 33956 1700
rect 34300 1660 34340 1700
rect 34684 1660 34724 1700
rect 35068 1660 35108 1700
rect 35452 1660 35492 1700
rect 35836 1660 35876 1700
rect 36220 1660 36260 1700
rect 36604 1660 36644 1700
rect 36988 1660 37028 1700
rect 37372 1660 37412 1700
rect 37756 1660 37796 1700
rect 38140 1660 38180 1700
rect 38524 1660 38564 1700
rect 38908 1660 38948 1700
rect 39292 1660 39332 1700
rect 39676 1660 39716 1700
rect 40060 1660 40100 1700
rect 40444 1660 40484 1700
rect 40828 1660 40868 1700
rect 41212 1660 41252 1700
rect 41596 1660 41636 1700
rect 41980 1660 42020 1700
rect 42364 1660 42404 1700
rect 50620 1660 50660 1700
rect 4928 1492 4968 1532
rect 5010 1492 5050 1532
rect 5092 1492 5132 1532
rect 5174 1492 5214 1532
rect 5256 1492 5296 1532
rect 20048 1492 20088 1532
rect 20130 1492 20170 1532
rect 20212 1492 20252 1532
rect 20294 1492 20334 1532
rect 20376 1492 20416 1532
rect 35168 1492 35208 1532
rect 35250 1492 35290 1532
rect 35332 1492 35372 1532
rect 35414 1492 35454 1532
rect 35496 1492 35536 1532
rect 50288 1492 50328 1532
rect 50370 1492 50410 1532
rect 50452 1492 50492 1532
rect 50534 1492 50574 1532
rect 50616 1492 50656 1532
<< metal2 >>
rect 0 11192 90 11212
rect 53190 11192 53280 11212
rect 0 11152 844 11192
rect 884 11152 893 11192
rect 50947 11152 50956 11192
rect 50996 11152 53280 11192
rect 0 11132 90 11152
rect 53190 11132 53280 11152
rect 0 10856 90 10876
rect 53190 10856 53280 10876
rect 0 10816 23596 10856
rect 23636 10816 23645 10856
rect 51043 10816 51052 10856
rect 51092 10816 53280 10856
rect 0 10796 90 10816
rect 53190 10796 53280 10816
rect 4919 10564 4928 10604
rect 4968 10564 5010 10604
rect 5050 10564 5092 10604
rect 5132 10564 5174 10604
rect 5214 10564 5256 10604
rect 5296 10564 5305 10604
rect 20039 10564 20048 10604
rect 20088 10564 20130 10604
rect 20170 10564 20212 10604
rect 20252 10564 20294 10604
rect 20334 10564 20376 10604
rect 20416 10564 20425 10604
rect 35159 10564 35168 10604
rect 35208 10564 35250 10604
rect 35290 10564 35332 10604
rect 35372 10564 35414 10604
rect 35454 10564 35496 10604
rect 35536 10564 35545 10604
rect 39139 10564 39148 10604
rect 39188 10564 46156 10604
rect 46196 10564 46205 10604
rect 50279 10564 50288 10604
rect 50328 10564 50370 10604
rect 50410 10564 50452 10604
rect 50492 10564 50534 10604
rect 50574 10564 50616 10604
rect 50656 10564 50665 10604
rect 0 10520 90 10540
rect 53190 10520 53280 10540
rect 0 10480 14284 10520
rect 14324 10480 14333 10520
rect 36931 10480 36940 10520
rect 36980 10480 44908 10520
rect 44948 10480 44957 10520
rect 50524 10480 51244 10520
rect 51284 10480 51293 10520
rect 51427 10480 51436 10520
rect 51476 10480 53280 10520
rect 0 10460 90 10480
rect 50524 10436 50564 10480
rect 53190 10460 53280 10480
rect 1603 10396 1612 10436
rect 1652 10396 1660 10436
rect 1700 10396 1783 10436
rect 4099 10396 4108 10436
rect 4148 10396 4156 10436
rect 4196 10396 4279 10436
rect 6595 10396 6604 10436
rect 6644 10396 6652 10436
rect 6692 10396 6775 10436
rect 9091 10396 9100 10436
rect 9140 10396 9148 10436
rect 9188 10396 9271 10436
rect 11587 10396 11596 10436
rect 11636 10396 11644 10436
rect 11684 10396 11767 10436
rect 14083 10396 14092 10436
rect 14132 10396 14140 10436
rect 14180 10396 14263 10436
rect 16579 10396 16588 10436
rect 16628 10396 16636 10436
rect 16676 10396 16759 10436
rect 19075 10396 19084 10436
rect 19124 10396 19132 10436
rect 19172 10396 19255 10436
rect 21571 10396 21580 10436
rect 21620 10396 21628 10436
rect 21668 10396 21751 10436
rect 24067 10396 24076 10436
rect 24116 10396 24124 10436
rect 24164 10396 24247 10436
rect 26563 10396 26572 10436
rect 26612 10396 26620 10436
rect 26660 10396 26743 10436
rect 29059 10396 29068 10436
rect 29108 10396 29116 10436
rect 29156 10396 29239 10436
rect 31555 10396 31564 10436
rect 31604 10396 31612 10436
rect 31652 10396 31735 10436
rect 34051 10396 34060 10436
rect 34100 10396 34108 10436
rect 34148 10396 34231 10436
rect 36748 10396 36980 10436
rect 39043 10396 39052 10436
rect 39092 10396 39100 10436
rect 39140 10396 39223 10436
rect 41539 10396 41548 10436
rect 41588 10396 41596 10436
rect 41636 10396 41719 10436
rect 44035 10396 44044 10436
rect 44084 10396 44092 10436
rect 44132 10396 44215 10436
rect 46531 10396 46540 10436
rect 46580 10396 46588 10436
rect 46628 10396 46711 10436
rect 49027 10396 49036 10436
rect 49076 10396 49084 10436
rect 49124 10396 49207 10436
rect 50515 10396 50524 10436
rect 50564 10396 50573 10436
rect 50899 10396 50908 10436
rect 50948 10396 51052 10436
rect 51092 10396 51101 10436
rect 51523 10396 51532 10436
rect 51572 10396 51772 10436
rect 51812 10396 51821 10436
rect 36748 10352 36788 10396
rect 24163 10312 24172 10352
rect 24212 10312 36788 10352
rect 36940 10352 36980 10396
rect 36940 10312 50708 10352
rect 51283 10312 51292 10352
rect 51332 10312 53108 10352
rect 1612 10228 26668 10268
rect 26708 10228 26717 10268
rect 34348 10228 36748 10268
rect 36788 10228 36797 10268
rect 39340 10228 44620 10268
rect 44660 10228 44669 10268
rect 0 10184 90 10204
rect 1612 10184 1652 10228
rect 34348 10184 34388 10228
rect 39340 10184 39380 10228
rect 50668 10184 50708 10312
rect 53068 10184 53108 10312
rect 53190 10184 53280 10204
rect 0 10144 1652 10184
rect 1769 10144 1900 10184
rect 1940 10144 1949 10184
rect 4265 10144 4396 10184
rect 4436 10144 4445 10184
rect 6761 10144 6892 10184
rect 6932 10144 6941 10184
rect 9257 10144 9388 10184
rect 9428 10144 9437 10184
rect 11875 10144 11884 10184
rect 11924 10144 13612 10184
rect 13652 10144 13661 10184
rect 14249 10144 14380 10184
rect 14420 10144 14429 10184
rect 16867 10144 16876 10184
rect 16916 10144 18412 10184
rect 18452 10144 18461 10184
rect 19363 10144 19372 10184
rect 19412 10144 20812 10184
rect 20852 10144 20861 10184
rect 21859 10144 21868 10184
rect 21908 10144 23116 10184
rect 23156 10144 23165 10184
rect 24355 10144 24364 10184
rect 24404 10144 25228 10184
rect 25268 10144 25277 10184
rect 26851 10144 26860 10184
rect 26900 10144 27820 10184
rect 27860 10144 27869 10184
rect 29225 10144 29356 10184
rect 29396 10144 29405 10184
rect 31843 10144 31852 10184
rect 31892 10144 33140 10184
rect 34339 10144 34348 10184
rect 34388 10144 34397 10184
rect 36547 10144 36556 10184
rect 36596 10144 36604 10184
rect 36644 10144 36727 10184
rect 36835 10144 36844 10184
rect 36884 10144 39148 10184
rect 39188 10144 39197 10184
rect 39331 10144 39340 10184
rect 39380 10144 39389 10184
rect 41827 10144 41836 10184
rect 41876 10144 43372 10184
rect 43412 10144 43421 10184
rect 44323 10144 44332 10184
rect 44372 10144 46636 10184
rect 46676 10144 46685 10184
rect 46819 10144 46828 10184
rect 46868 10144 48172 10184
rect 48212 10144 48221 10184
rect 48931 10144 48940 10184
rect 48980 10144 49324 10184
rect 49364 10144 49373 10184
rect 49603 10144 49612 10184
rect 49652 10144 49661 10184
rect 49961 10144 50092 10184
rect 50132 10144 50284 10184
rect 50324 10144 50333 10184
rect 50659 10144 50668 10184
rect 50708 10144 50717 10184
rect 50921 10144 51052 10184
rect 51092 10144 51101 10184
rect 51305 10144 51436 10184
rect 51476 10144 51485 10184
rect 51619 10144 51628 10184
rect 51668 10144 52012 10184
rect 52052 10144 52061 10184
rect 53068 10144 53280 10184
rect 0 10124 90 10144
rect 33100 10100 33140 10144
rect 49612 10100 49652 10144
rect 53190 10124 53280 10144
rect 15427 10060 15436 10100
rect 15476 10060 26572 10100
rect 26612 10060 26621 10100
rect 27715 10060 27724 10100
rect 27764 10060 30700 10100
rect 30740 10060 30749 10100
rect 33100 10060 43948 10100
rect 43988 10060 43997 10100
rect 47491 10060 47500 10100
rect 47540 10060 49652 10100
rect 49843 10060 49852 10100
rect 49892 10060 51532 10100
rect 51572 10060 51581 10100
rect 172 9976 24268 10016
rect 24308 9976 24317 10016
rect 26947 9976 26956 10016
rect 26996 9976 29012 10016
rect 29155 9976 29164 10016
rect 29204 9976 37996 10016
rect 38036 9976 38045 10016
rect 38092 9976 51052 10016
rect 51092 9976 51101 10016
rect 51667 9976 51676 10016
rect 51716 9976 53108 10016
rect 0 9848 90 9868
rect 172 9848 212 9976
rect 28972 9932 29012 9976
rect 38092 9932 38132 9976
rect 7180 9892 28876 9932
rect 28916 9892 28925 9932
rect 28972 9892 38132 9932
rect 38188 9892 46348 9932
rect 46388 9892 46397 9932
rect 50371 9892 50380 9932
rect 50420 9892 51436 9932
rect 51476 9892 51485 9932
rect 0 9808 212 9848
rect 3679 9808 3688 9848
rect 3728 9808 3770 9848
rect 3810 9808 3852 9848
rect 3892 9808 3934 9848
rect 3974 9808 4016 9848
rect 4056 9808 4065 9848
rect 0 9788 90 9808
rect 7180 9764 7220 9892
rect 38188 9848 38228 9892
rect 53068 9848 53108 9976
rect 53190 9848 53280 9868
rect 18799 9808 18808 9848
rect 18848 9808 18890 9848
rect 18930 9808 18972 9848
rect 19012 9808 19054 9848
rect 19094 9808 19136 9848
rect 19176 9808 19185 9848
rect 19363 9808 19372 9848
rect 19412 9808 27724 9848
rect 27764 9808 27773 9848
rect 27907 9808 27916 9848
rect 27956 9808 30028 9848
rect 30068 9808 30077 9848
rect 33919 9808 33928 9848
rect 33968 9808 34010 9848
rect 34050 9808 34092 9848
rect 34132 9808 34174 9848
rect 34214 9808 34256 9848
rect 34296 9808 34305 9848
rect 35011 9808 35020 9848
rect 35060 9808 38228 9848
rect 38275 9808 38284 9848
rect 38324 9808 47500 9848
rect 47540 9808 47549 9848
rect 49039 9808 49048 9848
rect 49088 9808 49130 9848
rect 49170 9808 49212 9848
rect 49252 9808 49294 9848
rect 49334 9808 49376 9848
rect 49416 9808 49425 9848
rect 53068 9808 53280 9848
rect 53190 9788 53280 9808
rect 835 9724 844 9764
rect 884 9724 7220 9764
rect 9379 9724 9388 9764
rect 9428 9724 37900 9764
rect 37940 9724 37949 9764
rect 38083 9724 38092 9764
rect 38132 9724 50612 9764
rect 13603 9640 13612 9680
rect 13652 9640 13852 9680
rect 13892 9640 13901 9680
rect 14371 9640 14380 9680
rect 14420 9640 15772 9680
rect 15812 9640 15821 9680
rect 18403 9640 18412 9680
rect 18452 9640 18460 9680
rect 18500 9640 18583 9680
rect 20803 9640 20812 9680
rect 20852 9640 20860 9680
rect 20900 9640 20983 9680
rect 23107 9640 23116 9680
rect 23156 9640 23164 9680
rect 23204 9640 23287 9680
rect 24019 9640 24028 9680
rect 24068 9640 24172 9680
rect 24212 9640 24221 9680
rect 25219 9640 25228 9680
rect 25268 9640 25372 9680
rect 25412 9640 25421 9680
rect 26825 9640 26908 9680
rect 26948 9640 26956 9680
rect 26996 9640 27005 9680
rect 27811 9640 27820 9680
rect 27860 9640 27868 9680
rect 27908 9640 27991 9680
rect 29033 9640 29116 9680
rect 29156 9640 29164 9680
rect 29204 9640 29213 9680
rect 29347 9640 29356 9680
rect 29396 9640 29692 9680
rect 29732 9640 29741 9680
rect 29836 9640 41596 9680
rect 41636 9640 41645 9680
rect 41740 9640 43084 9680
rect 43124 9640 43133 9680
rect 43363 9640 43372 9680
rect 43412 9640 43420 9680
rect 43460 9640 43543 9680
rect 43939 9640 43948 9680
rect 43988 9640 43996 9680
rect 44036 9640 44119 9680
rect 44899 9640 44908 9680
rect 44948 9640 44956 9680
rect 44996 9640 45079 9680
rect 46147 9640 46156 9680
rect 46196 9640 46204 9680
rect 46244 9640 46327 9680
rect 46627 9640 46636 9680
rect 46676 9640 46684 9680
rect 46724 9640 46807 9680
rect 48163 9640 48172 9680
rect 48212 9640 48220 9680
rect 48260 9640 48343 9680
rect 48809 9640 48892 9680
rect 48932 9640 48940 9680
rect 48980 9640 48989 9680
rect 29836 9596 29876 9640
rect 6883 9556 6892 9596
rect 6932 9556 29876 9596
rect 30019 9556 30028 9596
rect 30068 9556 40636 9596
rect 40676 9556 40685 9596
rect 0 9512 90 9532
rect 41740 9512 41780 9640
rect 41836 9556 43468 9596
rect 43508 9556 43517 9596
rect 43564 9556 43852 9596
rect 43892 9556 43901 9596
rect 45196 9556 47692 9596
rect 47732 9556 47741 9596
rect 41836 9512 41876 9556
rect 43564 9512 43604 9556
rect 45196 9512 45236 9556
rect 50572 9512 50612 9724
rect 50803 9640 50812 9680
rect 50852 9640 50956 9680
rect 50996 9640 51005 9680
rect 51187 9640 51196 9680
rect 51236 9640 51628 9680
rect 51668 9640 51677 9680
rect 51523 9556 51532 9596
rect 51572 9556 51956 9596
rect 51916 9512 51956 9556
rect 53190 9512 53280 9532
rect 0 9472 7220 9512
rect 13699 9472 13708 9512
rect 13748 9472 14092 9512
rect 14132 9472 14141 9512
rect 14275 9472 14284 9512
rect 14324 9472 14455 9512
rect 14515 9472 14524 9512
rect 14564 9472 15572 9512
rect 15619 9472 15628 9512
rect 15668 9472 16012 9512
rect 16052 9472 16061 9512
rect 18569 9472 18700 9512
rect 18740 9472 18749 9512
rect 21091 9472 21100 9512
rect 21140 9472 21292 9512
rect 21332 9472 21341 9512
rect 23395 9472 23404 9512
rect 23444 9472 23453 9512
rect 23587 9472 23596 9512
rect 23636 9472 23788 9512
rect 23828 9472 23837 9512
rect 25481 9472 25612 9512
rect 25652 9472 25661 9512
rect 26057 9472 26188 9512
rect 26228 9472 26237 9512
rect 26537 9472 26668 9512
rect 26708 9472 26717 9512
rect 28099 9472 28108 9512
rect 28148 9472 28588 9512
rect 28628 9472 28637 9512
rect 28745 9472 28876 9512
rect 28916 9472 28925 9512
rect 29801 9472 29932 9512
rect 29972 9472 29981 9512
rect 30089 9472 30220 9512
rect 30260 9472 30269 9512
rect 30451 9472 30460 9512
rect 30500 9472 38284 9512
rect 38324 9472 38333 9512
rect 40291 9472 40300 9512
rect 40340 9472 40349 9512
rect 40867 9472 40876 9512
rect 40916 9472 41780 9512
rect 41827 9472 41836 9512
rect 41876 9472 41885 9512
rect 42787 9472 42796 9512
rect 42836 9472 43604 9512
rect 43651 9472 43660 9512
rect 43700 9472 44180 9512
rect 44227 9472 44236 9512
rect 44276 9472 44285 9512
rect 45187 9472 45196 9512
rect 45236 9472 45245 9512
rect 46483 9472 46492 9512
rect 46532 9472 46868 9512
rect 46915 9472 46924 9512
rect 46964 9472 47252 9512
rect 47299 9472 47308 9512
rect 47348 9472 47357 9512
rect 48451 9472 48460 9512
rect 48500 9472 48596 9512
rect 48643 9472 48652 9512
rect 48692 9472 49996 9512
rect 50036 9472 50045 9512
rect 50563 9472 50572 9512
rect 50612 9472 50621 9512
rect 50825 9472 50956 9512
rect 50996 9472 51005 9512
rect 51427 9472 51436 9512
rect 51476 9472 51485 9512
rect 51619 9472 51628 9512
rect 51668 9472 51820 9512
rect 51860 9472 51869 9512
rect 51916 9472 53280 9512
rect 0 9452 90 9472
rect 7180 9428 7220 9472
rect 15532 9428 15572 9472
rect 23404 9428 23444 9472
rect 40300 9428 40340 9472
rect 44140 9428 44180 9472
rect 44236 9428 44276 9472
rect 7180 9388 15436 9428
rect 15476 9388 15485 9428
rect 15532 9388 19372 9428
rect 19412 9388 19421 9428
rect 23404 9388 23788 9428
rect 23828 9388 23837 9428
rect 23971 9388 23980 9428
rect 24020 9388 28396 9428
rect 28436 9388 28445 9428
rect 30691 9388 30700 9428
rect 30740 9388 40244 9428
rect 40300 9388 42700 9428
rect 42740 9388 42749 9428
rect 44131 9388 44140 9428
rect 44180 9388 44189 9428
rect 44236 9388 46156 9428
rect 46196 9388 46205 9428
rect 40204 9344 40244 9388
rect 46828 9344 46868 9472
rect 47212 9428 47252 9472
rect 47308 9428 47348 9472
rect 48556 9428 48596 9472
rect 47203 9388 47212 9428
rect 47252 9388 47261 9428
rect 47308 9388 48460 9428
rect 48500 9388 48509 9428
rect 48556 9388 49612 9428
rect 49652 9388 49661 9428
rect 4387 9304 4396 9344
rect 4436 9304 27916 9344
rect 27956 9304 27965 9344
rect 28204 9304 40060 9344
rect 40100 9304 40109 9344
rect 40204 9304 43564 9344
rect 43604 9304 43613 9344
rect 46828 9304 48076 9344
rect 48116 9304 48125 9344
rect 1891 9220 1900 9260
rect 1940 9220 7220 9260
rect 15610 9220 15619 9260
rect 15659 9220 20140 9260
rect 20180 9220 20189 9260
rect 26297 9220 26380 9260
rect 26420 9220 26428 9260
rect 26468 9220 26477 9260
rect 0 9176 90 9196
rect 7180 9176 7220 9220
rect 28204 9176 28244 9304
rect 28579 9220 28588 9260
rect 28628 9220 38228 9260
rect 38275 9220 38284 9260
rect 38324 9220 42556 9260
rect 42596 9220 42605 9260
rect 44611 9220 44620 9260
rect 44660 9220 47068 9260
rect 47108 9220 47117 9260
rect 47203 9220 47212 9260
rect 47252 9220 48940 9260
rect 48980 9220 48989 9260
rect 49036 9220 50092 9260
rect 50132 9220 50275 9260
rect 50315 9220 50324 9260
rect 0 9136 212 9176
rect 7180 9136 20524 9176
rect 20564 9136 20573 9176
rect 20803 9136 20812 9176
rect 20852 9136 28244 9176
rect 28291 9136 28300 9176
rect 28340 9136 38132 9176
rect 0 9116 90 9136
rect 172 9008 212 9136
rect 4919 9052 4928 9092
rect 4968 9052 5010 9092
rect 5050 9052 5092 9092
rect 5132 9052 5174 9092
rect 5214 9052 5256 9092
rect 5296 9052 5305 9092
rect 20039 9052 20048 9092
rect 20088 9052 20130 9092
rect 20170 9052 20212 9092
rect 20252 9052 20294 9092
rect 20334 9052 20376 9092
rect 20416 9052 20425 9092
rect 28387 9052 28396 9092
rect 28436 9052 35020 9092
rect 35060 9052 35069 9092
rect 35159 9052 35168 9092
rect 35208 9052 35250 9092
rect 35290 9052 35332 9092
rect 35372 9052 35414 9092
rect 35454 9052 35496 9092
rect 35536 9052 35545 9092
rect 38092 9008 38132 9136
rect 38188 9092 38228 9220
rect 43180 9136 45964 9176
rect 46004 9136 46013 9176
rect 46147 9136 46156 9176
rect 46196 9136 47308 9176
rect 47348 9136 47357 9176
rect 43180 9092 43220 9136
rect 38188 9052 43220 9092
rect 44131 9052 44140 9092
rect 44180 9052 48844 9092
rect 48884 9052 48893 9092
rect 49036 9008 49076 9220
rect 50279 9052 50288 9092
rect 50328 9052 50370 9092
rect 50410 9052 50452 9092
rect 50492 9052 50534 9092
rect 50574 9052 50616 9092
rect 50656 9052 50665 9092
rect 172 8968 28108 9008
rect 28148 8968 28157 9008
rect 29923 8968 29932 9008
rect 29972 8968 37996 9008
rect 38036 8968 38045 9008
rect 38092 8968 44620 9008
rect 44660 8968 44669 9008
rect 46147 8968 46156 9008
rect 46196 8968 49076 9008
rect 739 8884 748 8924
rect 788 8884 7220 8924
rect 0 8840 90 8860
rect 7180 8840 7220 8884
rect 23020 8884 26188 8924
rect 26228 8884 26237 8924
rect 26563 8884 26572 8924
rect 26612 8884 30220 8924
rect 30260 8884 30269 8924
rect 33715 8884 33724 8924
rect 33764 8884 47212 8924
rect 47252 8884 47261 8924
rect 23020 8840 23060 8884
rect 51436 8840 51476 9472
rect 53190 9452 53280 9472
rect 51667 9220 51676 9260
rect 51716 9220 51725 9260
rect 52051 9220 52060 9260
rect 52100 9220 52684 9260
rect 52724 9220 52733 9260
rect 51676 9176 51716 9220
rect 53190 9176 53280 9196
rect 51676 9136 53280 9176
rect 53190 9116 53280 9136
rect 53190 8840 53280 8860
rect 0 8800 1228 8840
rect 1268 8800 1277 8840
rect 7180 8800 23060 8840
rect 25843 8800 25852 8840
rect 25892 8800 28244 8840
rect 28339 8800 28348 8840
rect 28388 8800 51476 8840
rect 52675 8800 52684 8840
rect 52724 8800 53280 8840
rect 0 8780 90 8800
rect 28204 8756 28244 8800
rect 53190 8780 53280 8800
rect 7180 8716 27764 8756
rect 28204 8716 43276 8756
rect 43316 8716 43325 8756
rect 43555 8716 43564 8756
rect 43604 8716 46156 8756
rect 46196 8716 46205 8756
rect 46339 8716 46348 8756
rect 46388 8716 51476 8756
rect 7180 8672 7220 8716
rect 27724 8672 27764 8716
rect 51436 8672 51476 8716
rect 1123 8632 1132 8672
rect 1172 8632 7220 8672
rect 24259 8632 24268 8672
rect 24308 8632 25612 8672
rect 25652 8632 25661 8672
rect 26371 8632 26380 8672
rect 26420 8632 27340 8672
rect 27380 8632 27389 8672
rect 27715 8632 27724 8672
rect 27764 8632 27773 8672
rect 27833 8632 27916 8672
rect 27956 8632 27964 8672
rect 28004 8632 28013 8672
rect 28099 8632 28108 8672
rect 28148 8632 28279 8672
rect 33187 8632 33196 8672
rect 33236 8632 33292 8672
rect 33332 8632 33484 8672
rect 33524 8632 33964 8672
rect 34004 8632 34252 8672
rect 34292 8632 34540 8672
rect 34580 8632 34828 8672
rect 34868 8632 35116 8672
rect 35156 8632 35404 8672
rect 35444 8632 35692 8672
rect 35732 8632 35884 8672
rect 35924 8632 35933 8672
rect 37987 8632 37996 8672
rect 38036 8632 46924 8672
rect 46964 8632 46973 8672
rect 51427 8632 51436 8672
rect 51476 8632 51485 8672
rect 51667 8632 51676 8672
rect 51716 8632 51764 8672
rect 51811 8632 51820 8672
rect 51860 8632 51991 8672
rect 52051 8632 52060 8672
rect 52100 8632 53164 8672
rect 53204 8632 53213 8672
rect 51724 8588 51764 8632
rect 51724 8548 52532 8588
rect 0 8504 90 8524
rect 52492 8504 52532 8548
rect 53190 8504 53280 8524
rect 0 8464 23348 8504
rect 52492 8464 53280 8504
rect 0 8444 90 8464
rect 3679 8296 3688 8336
rect 3728 8296 3770 8336
rect 3810 8296 3852 8336
rect 3892 8296 3934 8336
rect 3974 8296 4016 8336
rect 4056 8296 4065 8336
rect 18799 8296 18808 8336
rect 18848 8296 18890 8336
rect 18930 8296 18972 8336
rect 19012 8296 19054 8336
rect 19094 8296 19136 8336
rect 19176 8296 19185 8336
rect 0 8168 90 8188
rect 0 8128 1324 8168
rect 1364 8128 1373 8168
rect 0 8108 90 8128
rect 1219 8044 1228 8084
rect 1268 8044 23252 8084
rect 355 7960 364 8000
rect 404 7960 7220 8000
rect 7180 7916 7220 7960
rect 23212 7916 23252 8044
rect 23308 8000 23348 8464
rect 53190 8444 53280 8464
rect 33919 8296 33928 8336
rect 33968 8296 34010 8336
rect 34050 8296 34092 8336
rect 34132 8296 34174 8336
rect 34214 8296 34256 8336
rect 34296 8296 34305 8336
rect 49039 8296 49048 8336
rect 49088 8296 49130 8336
rect 49170 8296 49212 8336
rect 49252 8296 49294 8336
rect 49334 8296 49376 8336
rect 49416 8296 49425 8336
rect 53190 8168 53280 8188
rect 23539 8128 23548 8168
rect 23588 8128 23980 8168
rect 24020 8128 24029 8168
rect 28243 8128 28252 8168
rect 28292 8128 51628 8168
rect 51668 8128 51677 8168
rect 53155 8128 53164 8168
rect 53204 8128 53280 8168
rect 53190 8108 53280 8128
rect 23875 8044 23884 8084
rect 23924 8044 31604 8084
rect 31699 8044 31708 8084
rect 31748 8044 38092 8084
rect 38132 8044 38141 8084
rect 23299 7960 23308 8000
rect 23348 7960 23357 8000
rect 28003 7960 28012 8000
rect 28052 7960 28061 8000
rect 31459 7960 31468 8000
rect 31508 7960 31517 8000
rect 28012 7916 28052 7960
rect 7180 7876 23060 7916
rect 23212 7876 28052 7916
rect 0 7832 90 7852
rect 23020 7832 23060 7876
rect 31468 7832 31508 7960
rect 31564 7916 31604 8044
rect 34819 7960 34828 8000
rect 34868 7960 35212 8000
rect 35252 7960 35261 8000
rect 43180 7960 51436 8000
rect 51476 7960 51485 8000
rect 51811 7960 51820 8000
rect 51860 7960 51869 8000
rect 43180 7916 43220 7960
rect 51820 7916 51860 7960
rect 31564 7876 34924 7916
rect 34964 7876 34973 7916
rect 35020 7876 35252 7916
rect 35299 7876 35308 7916
rect 35348 7876 43220 7916
rect 46060 7876 51860 7916
rect 35020 7832 35060 7876
rect 0 7792 21580 7832
rect 21620 7792 21629 7832
rect 23020 7792 31508 7832
rect 33100 7792 35060 7832
rect 35212 7832 35252 7876
rect 46060 7832 46100 7876
rect 53190 7832 53280 7852
rect 35212 7792 46100 7832
rect 51667 7792 51676 7832
rect 51716 7792 53280 7832
rect 0 7772 90 7792
rect 33100 7748 33140 7792
rect 53190 7772 53280 7792
rect 25699 7708 25708 7748
rect 25748 7708 33140 7748
rect 33187 7708 33196 7748
rect 33236 7708 33475 7748
rect 33515 7708 33524 7748
rect 35443 7708 35452 7748
rect 35492 7708 44236 7748
rect 44276 7708 44285 7748
rect 52051 7708 52060 7748
rect 52100 7708 52109 7748
rect 52060 7664 52100 7708
rect 38083 7624 38092 7664
rect 38132 7624 50804 7664
rect 52060 7624 53164 7664
rect 53204 7624 53213 7664
rect 50764 7580 50804 7624
rect 4919 7540 4928 7580
rect 4968 7540 5010 7580
rect 5050 7540 5092 7580
rect 5132 7540 5174 7580
rect 5214 7540 5256 7580
rect 5296 7540 5305 7580
rect 20039 7540 20048 7580
rect 20088 7540 20130 7580
rect 20170 7540 20212 7580
rect 20252 7540 20294 7580
rect 20334 7540 20376 7580
rect 20416 7540 20425 7580
rect 35159 7540 35168 7580
rect 35208 7540 35250 7580
rect 35290 7540 35332 7580
rect 35372 7540 35414 7580
rect 35454 7540 35496 7580
rect 35536 7540 35545 7580
rect 50279 7540 50288 7580
rect 50328 7540 50370 7580
rect 50410 7540 50452 7580
rect 50492 7540 50534 7580
rect 50574 7540 50616 7580
rect 50656 7540 50665 7580
rect 50764 7540 52012 7580
rect 52052 7540 52061 7580
rect 0 7496 90 7516
rect 53190 7496 53280 7516
rect 0 7456 22924 7496
rect 22964 7456 22973 7496
rect 53155 7456 53164 7496
rect 53204 7456 53280 7496
rect 0 7436 90 7456
rect 53190 7436 53280 7456
rect 23020 7288 34828 7328
rect 34868 7288 35212 7328
rect 35252 7288 35500 7328
rect 35540 7288 35549 7328
rect 23020 7244 23060 7288
rect 451 7204 460 7244
rect 500 7204 23060 7244
rect 29644 7204 30356 7244
rect 0 7160 90 7180
rect 29644 7160 29684 7204
rect 30316 7160 30356 7204
rect 35116 7204 35636 7244
rect 35116 7160 35156 7204
rect 0 7120 1228 7160
rect 1268 7120 1277 7160
rect 10723 7120 10732 7160
rect 10772 7120 18892 7160
rect 18932 7120 18941 7160
rect 21571 7120 21580 7160
rect 21620 7120 23596 7160
rect 23636 7120 23645 7160
rect 23753 7120 23836 7160
rect 23876 7120 23884 7160
rect 23924 7120 23933 7160
rect 24163 7120 24172 7160
rect 24212 7120 29684 7160
rect 29731 7120 29740 7160
rect 29780 7120 29789 7160
rect 29836 7120 30220 7160
rect 30260 7120 30269 7160
rect 30316 7120 35156 7160
rect 35596 7160 35636 7204
rect 53190 7160 53280 7180
rect 35596 7120 51436 7160
rect 51476 7120 51485 7160
rect 51811 7120 51820 7160
rect 51860 7120 51916 7160
rect 51956 7120 51991 7160
rect 52051 7120 52060 7160
rect 52100 7120 53280 7160
rect 0 7100 90 7120
rect 29740 7076 29780 7120
rect 1027 7036 1036 7076
rect 1076 7036 29780 7076
rect 19123 6952 19132 6992
rect 19172 6952 19948 6992
rect 19988 6952 19997 6992
rect 0 6824 90 6844
rect 0 6784 3572 6824
rect 3679 6784 3688 6824
rect 3728 6784 3770 6824
rect 3810 6784 3852 6824
rect 3892 6784 3934 6824
rect 3974 6784 4016 6824
rect 4056 6784 4065 6824
rect 18799 6784 18808 6824
rect 18848 6784 18890 6824
rect 18930 6784 18972 6824
rect 19012 6784 19054 6824
rect 19094 6784 19136 6824
rect 19176 6784 19185 6824
rect 0 6764 90 6784
rect 3532 6740 3572 6784
rect 3532 6700 21580 6740
rect 21620 6700 21629 6740
rect 29836 6656 29876 7120
rect 53190 7100 53280 7120
rect 30451 7036 30460 7076
rect 30500 7036 51820 7076
rect 51860 7036 51869 7076
rect 29971 6952 29980 6992
rect 30020 6952 33140 6992
rect 51667 6952 51676 6992
rect 51716 6952 53108 6992
rect 33100 6908 33140 6952
rect 33100 6868 51436 6908
rect 51476 6868 51485 6908
rect 53068 6824 53108 6952
rect 53190 6824 53280 6844
rect 33919 6784 33928 6824
rect 33968 6784 34010 6824
rect 34050 6784 34092 6824
rect 34132 6784 34174 6824
rect 34214 6784 34256 6824
rect 34296 6784 34305 6824
rect 49039 6784 49048 6824
rect 49088 6784 49130 6824
rect 49170 6784 49212 6824
rect 49252 6784 49294 6824
rect 49334 6784 49376 6824
rect 49416 6784 49425 6824
rect 53068 6784 53280 6824
rect 53190 6764 53280 6784
rect 1315 6616 1324 6656
rect 1364 6616 29876 6656
rect 25577 6532 25660 6572
rect 25700 6532 25708 6572
rect 25748 6532 25757 6572
rect 0 6488 90 6508
rect 53190 6488 53280 6508
rect 0 6448 1420 6488
rect 1460 6448 1469 6488
rect 22601 6448 22732 6488
rect 22772 6448 22781 6488
rect 22915 6448 22924 6488
rect 22964 6448 25420 6488
rect 25460 6448 25469 6488
rect 25673 6448 25804 6488
rect 25844 6448 25853 6488
rect 35491 6448 35500 6488
rect 35540 6448 35788 6488
rect 35828 6448 36172 6488
rect 36212 6448 36460 6488
rect 36500 6448 36748 6488
rect 36788 6448 37036 6488
rect 37076 6448 37324 6488
rect 37364 6448 37612 6488
rect 37652 6448 37900 6488
rect 37940 6448 37949 6488
rect 38275 6448 38284 6488
rect 38324 6448 38333 6488
rect 43180 6448 51436 6488
rect 51476 6448 51485 6488
rect 51689 6448 51820 6488
rect 51860 6448 51869 6488
rect 52051 6448 52060 6488
rect 52100 6448 53280 6488
rect 0 6428 90 6448
rect 38284 6404 38324 6448
rect 259 6364 268 6404
rect 308 6364 7220 6404
rect 7180 6320 7220 6364
rect 20140 6364 38324 6404
rect 20140 6320 20180 6364
rect 43180 6320 43220 6448
rect 53190 6428 53280 6448
rect 7180 6280 20180 6320
rect 26035 6280 26044 6320
rect 26084 6280 43220 6320
rect 22841 6196 22924 6236
rect 22964 6196 22972 6236
rect 23012 6196 23021 6236
rect 35980 6196 36028 6236
rect 36068 6196 36077 6236
rect 38515 6196 38524 6236
rect 38564 6196 47500 6236
rect 47540 6196 47549 6236
rect 51667 6196 51676 6236
rect 51716 6196 51725 6236
rect 0 6152 90 6172
rect 35980 6152 36020 6196
rect 51676 6152 51716 6196
rect 53190 6152 53280 6172
rect 0 6112 25804 6152
rect 25844 6112 25853 6152
rect 35980 6112 50804 6152
rect 51676 6112 53280 6152
rect 0 6092 90 6112
rect 50764 6068 50804 6112
rect 53190 6092 53280 6112
rect 4919 6028 4928 6068
rect 4968 6028 5010 6068
rect 5050 6028 5092 6068
rect 5132 6028 5174 6068
rect 5214 6028 5256 6068
rect 5296 6028 5305 6068
rect 20039 6028 20048 6068
rect 20088 6028 20130 6068
rect 20170 6028 20212 6068
rect 20252 6028 20294 6068
rect 20334 6028 20376 6068
rect 20416 6028 20425 6068
rect 35159 6028 35168 6068
rect 35208 6028 35250 6068
rect 35290 6028 35332 6068
rect 35372 6028 35414 6068
rect 35454 6028 35496 6068
rect 35536 6028 35545 6068
rect 50279 6028 50288 6068
rect 50328 6028 50370 6068
rect 50410 6028 50452 6068
rect 50492 6028 50534 6068
rect 50574 6028 50616 6068
rect 50656 6028 50665 6068
rect 50764 6028 52108 6068
rect 52148 6028 52157 6068
rect 0 5816 90 5836
rect 53190 5816 53280 5836
rect 0 5776 22732 5816
rect 22772 5776 22781 5816
rect 35657 5776 35788 5816
rect 35828 5776 36076 5816
rect 36116 5776 36125 5816
rect 52051 5776 52060 5816
rect 52100 5776 53280 5816
rect 0 5756 90 5776
rect 53190 5756 53280 5776
rect 22915 5692 22924 5732
rect 22964 5692 51860 5732
rect 51820 5648 51860 5692
rect 21571 5608 21580 5648
rect 21620 5608 23884 5648
rect 23924 5608 23933 5648
rect 24041 5608 24124 5648
rect 24164 5608 24172 5648
rect 24212 5608 24221 5648
rect 27689 5608 27820 5648
rect 27860 5608 27869 5648
rect 43180 5608 51436 5648
rect 51476 5608 51485 5648
rect 51811 5608 51820 5648
rect 51860 5608 51869 5648
rect 43180 5564 43220 5608
rect 19939 5524 19948 5564
rect 19988 5524 23060 5564
rect 0 5480 90 5500
rect 0 5440 10732 5480
rect 10772 5440 10781 5480
rect 0 5420 90 5440
rect 23020 5396 23060 5524
rect 27916 5524 43220 5564
rect 51667 5524 51676 5564
rect 51716 5524 52532 5564
rect 27916 5396 27956 5524
rect 52492 5480 52532 5524
rect 53190 5480 53280 5500
rect 28051 5440 28060 5480
rect 28100 5440 33140 5480
rect 52492 5440 53280 5480
rect 23020 5356 27956 5396
rect 33100 5396 33140 5440
rect 53190 5420 53280 5440
rect 33100 5356 51916 5396
rect 51956 5356 51965 5396
rect 3679 5272 3688 5312
rect 3728 5272 3770 5312
rect 3810 5272 3852 5312
rect 3892 5272 3934 5312
rect 3974 5272 4016 5312
rect 4056 5272 4065 5312
rect 18799 5272 18808 5312
rect 18848 5272 18890 5312
rect 18930 5272 18972 5312
rect 19012 5272 19054 5312
rect 19094 5272 19136 5312
rect 19176 5272 19185 5312
rect 33919 5272 33928 5312
rect 33968 5272 34010 5312
rect 34050 5272 34092 5312
rect 34132 5272 34174 5312
rect 34214 5272 34256 5312
rect 34296 5272 34305 5312
rect 49039 5272 49048 5312
rect 49088 5272 49130 5312
rect 49170 5272 49212 5312
rect 49252 5272 49294 5312
rect 49334 5272 49376 5312
rect 49416 5272 49425 5312
rect 1219 5188 1228 5228
rect 1268 5188 27820 5228
rect 27860 5188 27869 5228
rect 0 5144 90 5164
rect 53190 5144 53280 5164
rect 0 5104 1132 5144
rect 1172 5104 1181 5144
rect 7180 5104 15092 5144
rect 27907 5104 27916 5144
rect 27956 5104 33140 5144
rect 52051 5104 52060 5144
rect 52100 5104 53280 5144
rect 0 5084 90 5104
rect 7180 5060 7220 5104
rect 1411 5020 1420 5060
rect 1460 5020 7220 5060
rect 15052 5060 15092 5104
rect 15052 5020 30068 5060
rect 30028 4976 30068 5020
rect 33100 4976 33140 5104
rect 53190 5084 53280 5104
rect 43180 5020 51860 5060
rect 43180 4976 43220 5020
rect 51820 4976 51860 5020
rect 14537 4936 14668 4976
rect 14708 4936 14717 4976
rect 15235 4936 15244 4976
rect 15284 4936 18124 4976
rect 18164 4936 18173 4976
rect 24041 4936 24172 4976
rect 24212 4936 24221 4976
rect 24835 4936 24844 4976
rect 24884 4936 24893 4976
rect 25219 4936 25228 4976
rect 25268 4936 25277 4976
rect 30019 4936 30028 4976
rect 30068 4936 30077 4976
rect 33100 4936 43220 4976
rect 51305 4936 51436 4976
rect 51476 4936 51485 4976
rect 51811 4936 51820 4976
rect 51860 4936 51869 4976
rect 24844 4892 24884 4936
rect 5443 4852 5452 4892
rect 5492 4852 24884 4892
rect 0 4808 90 4828
rect 25228 4808 25268 4936
rect 43180 4852 51820 4892
rect 51860 4852 51869 4892
rect 43180 4808 43220 4852
rect 53190 4808 53280 4828
rect 0 4768 1036 4808
rect 1076 4768 1085 4808
rect 5827 4768 5836 4808
rect 5876 4768 25268 4808
rect 30259 4768 30268 4808
rect 30308 4768 43220 4808
rect 51667 4768 51676 4808
rect 51716 4768 53280 4808
rect 0 4748 90 4768
rect 53190 4748 53280 4768
rect 14899 4684 14908 4724
rect 14948 4684 15340 4724
rect 15380 4684 15389 4724
rect 15475 4684 15484 4724
rect 15524 4684 15628 4724
rect 15668 4684 15677 4724
rect 24403 4684 24412 4724
rect 24452 4684 24844 4724
rect 24884 4684 24893 4724
rect 25075 4684 25084 4724
rect 25124 4684 25364 4724
rect 25459 4684 25468 4724
rect 25508 4684 25516 4724
rect 25556 4684 25639 4724
rect 25324 4640 25364 4684
rect 14659 4600 14668 4640
rect 14708 4600 17740 4640
rect 17780 4600 17789 4640
rect 25324 4600 26092 4640
rect 26132 4600 26141 4640
rect 4919 4516 4928 4556
rect 4968 4516 5010 4556
rect 5050 4516 5092 4556
rect 5132 4516 5174 4556
rect 5214 4516 5256 4556
rect 5296 4516 5305 4556
rect 20039 4516 20048 4556
rect 20088 4516 20130 4556
rect 20170 4516 20212 4556
rect 20252 4516 20294 4556
rect 20334 4516 20376 4556
rect 20416 4516 20425 4556
rect 35159 4516 35168 4556
rect 35208 4516 35250 4556
rect 35290 4516 35332 4556
rect 35372 4516 35414 4556
rect 35454 4516 35496 4556
rect 35536 4516 35545 4556
rect 50279 4516 50288 4556
rect 50328 4516 50370 4556
rect 50410 4516 50452 4556
rect 50492 4516 50534 4556
rect 50574 4516 50616 4556
rect 50656 4516 50665 4556
rect 0 4472 90 4492
rect 53190 4472 53280 4492
rect 0 4432 364 4472
rect 404 4432 413 4472
rect 6211 4432 6220 4472
rect 6260 4432 24172 4472
rect 24212 4432 24221 4472
rect 52060 4432 53280 4472
rect 0 4412 90 4432
rect 22819 4348 22828 4388
rect 22868 4348 23156 4388
rect 27331 4348 27340 4388
rect 27380 4348 33044 4388
rect 6595 4264 6604 4304
rect 6644 4264 23060 4304
rect 11587 4180 11596 4220
rect 11636 4180 12980 4220
rect 13699 4180 13708 4220
rect 13748 4180 16300 4220
rect 16340 4180 16349 4220
rect 16396 4180 18508 4220
rect 18548 4180 18557 4220
rect 18691 4180 18700 4220
rect 18740 4180 22924 4220
rect 22964 4180 22973 4220
rect 0 4136 90 4156
rect 0 4096 460 4136
rect 500 4096 509 4136
rect 0 4076 90 4096
rect 12940 4052 12980 4180
rect 16396 4136 16436 4180
rect 23020 4136 23060 4264
rect 23116 4220 23156 4348
rect 33004 4304 33044 4348
rect 52060 4304 52100 4432
rect 53190 4412 53280 4432
rect 23299 4264 23308 4304
rect 23348 4264 32908 4304
rect 32948 4264 32957 4304
rect 33004 4264 43220 4304
rect 44227 4264 44236 4304
rect 44276 4264 51476 4304
rect 52051 4264 52060 4304
rect 52100 4264 52109 4304
rect 23116 4180 38900 4220
rect 38860 4136 38900 4180
rect 13411 4096 13420 4136
rect 13460 4096 16204 4136
rect 16244 4096 16253 4136
rect 16387 4096 16396 4136
rect 16436 4096 16445 4136
rect 16867 4096 16876 4136
rect 16916 4096 18316 4136
rect 18356 4096 18365 4136
rect 18700 4096 18932 4136
rect 19171 4096 19180 4136
rect 19220 4096 19660 4136
rect 19700 4096 19709 4136
rect 19843 4096 19852 4136
rect 19892 4096 22964 4136
rect 23011 4096 23020 4136
rect 23060 4096 23069 4136
rect 27881 4096 28012 4136
rect 28052 4096 28061 4136
rect 28195 4096 28204 4136
rect 28244 4096 35020 4136
rect 35060 4096 35069 4136
rect 38851 4096 38860 4136
rect 38900 4096 38909 4136
rect 18700 4052 18740 4096
rect 12940 4012 18740 4052
rect 18892 4052 18932 4096
rect 18892 4012 22636 4052
rect 22676 4012 22685 4052
rect 13651 3928 13660 3968
rect 13700 3928 14380 3968
rect 14420 3928 14429 3968
rect 16627 3928 16636 3968
rect 16676 3928 16876 3968
rect 16916 3928 16925 3968
rect 17107 3928 17116 3968
rect 17156 3928 18412 3968
rect 18452 3928 18461 3968
rect 19411 3928 19420 3968
rect 19460 3928 20716 3968
rect 20756 3928 20765 3968
rect 12739 3844 12748 3884
rect 12788 3844 18604 3884
rect 18644 3844 18653 3884
rect 18700 3844 22732 3884
rect 22772 3844 22781 3884
rect 0 3800 90 3820
rect 18700 3800 18740 3844
rect 22924 3800 22964 4096
rect 28243 4012 28252 4052
rect 28292 4012 28340 4052
rect 28387 4012 28396 4052
rect 28436 4012 36940 4052
rect 36980 4012 36989 4052
rect 28300 3968 28340 4012
rect 23251 3928 23260 3968
rect 23300 3928 24076 3968
rect 24116 3928 24125 3968
rect 28300 3928 29164 3968
rect 29204 3928 29213 3968
rect 37795 3928 37804 3968
rect 37844 3928 38620 3968
rect 38660 3928 38669 3968
rect 43180 3884 43220 4264
rect 47491 4180 47500 4220
rect 47540 4180 51092 4220
rect 51052 4136 51092 4180
rect 51436 4136 51476 4264
rect 53190 4136 53280 4156
rect 50729 4096 50860 4136
rect 50900 4096 50909 4136
rect 51043 4096 51052 4136
rect 51092 4096 51101 4136
rect 51427 4096 51436 4136
rect 51476 4096 51485 4136
rect 51811 4096 51820 4136
rect 51860 4096 52012 4136
rect 52052 4096 52061 4136
rect 52492 4096 53280 4136
rect 52492 4052 52532 4096
rect 53190 4076 53280 4096
rect 51667 4012 51676 4052
rect 51716 4012 52532 4052
rect 51283 3928 51292 3968
rect 51332 3928 51956 3968
rect 23107 3844 23116 3884
rect 23156 3844 28012 3884
rect 28052 3844 28061 3884
rect 28291 3844 28300 3884
rect 28340 3844 31372 3884
rect 31412 3844 31421 3884
rect 43180 3844 51860 3884
rect 0 3760 748 3800
rect 788 3760 797 3800
rect 3679 3760 3688 3800
rect 3728 3760 3770 3800
rect 3810 3760 3852 3800
rect 3892 3760 3934 3800
rect 3974 3760 4016 3800
rect 4056 3760 4065 3800
rect 14275 3760 14284 3800
rect 14324 3760 18740 3800
rect 18799 3760 18808 3800
rect 18848 3760 18890 3800
rect 18930 3760 18972 3800
rect 19012 3760 19054 3800
rect 19094 3760 19136 3800
rect 19176 3760 19185 3800
rect 21955 3760 21964 3800
rect 22004 3760 22828 3800
rect 22868 3760 22877 3800
rect 22924 3760 30988 3800
rect 31028 3760 31037 3800
rect 33919 3760 33928 3800
rect 33968 3760 34010 3800
rect 34050 3760 34092 3800
rect 34132 3760 34174 3800
rect 34214 3760 34256 3800
rect 34296 3760 34305 3800
rect 49039 3760 49048 3800
rect 49088 3760 49130 3800
rect 49170 3760 49212 3800
rect 49252 3760 49294 3800
rect 49334 3760 49376 3800
rect 49416 3760 49425 3800
rect 0 3740 90 3760
rect 13027 3676 13036 3716
rect 13076 3676 20140 3716
rect 20180 3676 20189 3716
rect 23203 3676 23212 3716
rect 23252 3676 30220 3716
rect 30260 3676 30269 3716
rect 4099 3592 4108 3632
rect 4148 3592 17108 3632
rect 18307 3592 18316 3632
rect 18356 3592 18796 3632
rect 18836 3592 18845 3632
rect 18892 3592 20620 3632
rect 20660 3592 20669 3632
rect 20803 3592 20812 3632
rect 20852 3592 22580 3632
rect 22771 3592 22780 3632
rect 22820 3592 22924 3632
rect 22964 3592 22973 3632
rect 23107 3592 23116 3632
rect 23156 3592 32428 3632
rect 32468 3592 32477 3632
rect 10435 3508 10444 3548
rect 10484 3508 12940 3548
rect 12980 3508 12989 3548
rect 14188 3508 16972 3548
rect 17012 3508 17021 3548
rect 0 3464 90 3484
rect 14188 3464 14228 3508
rect 17068 3464 17108 3592
rect 18892 3548 18932 3592
rect 17251 3508 17260 3548
rect 17300 3508 18932 3548
rect 19795 3508 19804 3548
rect 19844 3508 22060 3548
rect 22100 3508 22109 3548
rect 22540 3464 22580 3592
rect 23203 3508 23212 3548
rect 23252 3508 31700 3548
rect 31660 3464 31700 3508
rect 36076 3508 36404 3548
rect 0 3424 268 3464
rect 308 3424 317 3464
rect 14179 3424 14188 3464
rect 14228 3424 14237 3464
rect 14659 3424 14668 3464
rect 14708 3424 16780 3464
rect 16820 3424 16829 3464
rect 17068 3424 17116 3464
rect 17156 3424 17165 3464
rect 18403 3424 18412 3464
rect 18452 3424 18700 3464
rect 18740 3424 18749 3464
rect 19433 3424 19564 3464
rect 19604 3424 19613 3464
rect 20515 3424 20524 3464
rect 20564 3424 21292 3464
rect 21332 3424 21341 3464
rect 21449 3424 21532 3464
rect 21572 3424 21580 3464
rect 21620 3424 21629 3464
rect 21706 3424 21715 3464
rect 21755 3424 21772 3464
rect 21812 3424 21895 3464
rect 22531 3424 22540 3464
rect 22580 3424 22589 3464
rect 25891 3424 25900 3464
rect 25940 3424 28204 3464
rect 28244 3424 28253 3464
rect 28963 3424 28972 3464
rect 29012 3424 29644 3464
rect 29684 3424 29693 3464
rect 30211 3424 30220 3464
rect 30260 3424 30412 3464
rect 30452 3424 30461 3464
rect 30595 3424 30604 3464
rect 30644 3424 30796 3464
rect 30836 3424 30845 3464
rect 30979 3424 30988 3464
rect 31028 3424 31219 3464
rect 31259 3424 31268 3464
rect 31651 3424 31660 3464
rect 31700 3424 31709 3464
rect 32297 3424 32428 3464
rect 32468 3424 32477 3464
rect 32777 3424 32908 3464
rect 32948 3424 32957 3464
rect 33641 3424 33772 3464
rect 33812 3424 33821 3464
rect 34889 3424 35020 3464
rect 35060 3424 35069 3464
rect 35203 3424 35212 3464
rect 35252 3424 35731 3464
rect 35771 3424 35780 3464
rect 0 3404 90 3424
rect 36076 3380 36116 3508
rect 10819 3340 10828 3380
rect 10868 3340 28012 3380
rect 28052 3340 28061 3380
rect 28108 3340 31180 3380
rect 31220 3340 31229 3380
rect 31276 3340 36116 3380
rect 36172 3424 36268 3464
rect 36308 3424 36317 3464
rect 28108 3296 28148 3340
rect 31276 3296 31316 3340
rect 36172 3296 36212 3424
rect 36364 3380 36404 3508
rect 51820 3464 51860 3844
rect 51916 3464 51956 3928
rect 53190 3800 53280 3820
rect 52060 3760 53280 3800
rect 52060 3632 52100 3760
rect 53190 3740 53280 3760
rect 52051 3592 52060 3632
rect 52100 3592 52109 3632
rect 53190 3464 53280 3484
rect 36809 3424 36940 3464
rect 36980 3424 36989 3464
rect 37577 3424 37708 3464
rect 37748 3424 37757 3464
rect 41731 3424 41740 3464
rect 41780 3424 42028 3464
rect 42068 3424 42412 3464
rect 42452 3424 42700 3464
rect 42740 3424 42988 3464
rect 43028 3424 43276 3464
rect 43316 3424 43564 3464
rect 43604 3424 43852 3464
rect 43892 3424 44140 3464
rect 44180 3424 44428 3464
rect 44468 3424 44716 3464
rect 44756 3424 44765 3464
rect 47203 3424 47212 3464
rect 47252 3424 51436 3464
rect 51476 3424 51485 3464
rect 51811 3424 51820 3464
rect 51860 3424 51869 3464
rect 51916 3424 53280 3464
rect 53190 3404 53280 3424
rect 36364 3340 44716 3380
rect 44756 3340 44765 3380
rect 11203 3256 11212 3296
rect 11252 3256 28148 3296
rect 31027 3256 31036 3296
rect 31076 3256 31316 3296
rect 31411 3256 31420 3296
rect 31460 3256 32236 3296
rect 32276 3256 32285 3296
rect 36172 3256 36308 3296
rect 42259 3256 42268 3296
rect 42308 3256 49420 3296
rect 49460 3256 49469 3296
rect 49987 3256 49996 3296
rect 50036 3256 50188 3296
rect 50228 3256 50284 3296
rect 50324 3256 50860 3296
rect 50900 3256 50909 3296
rect 14419 3172 14428 3212
rect 14468 3172 14668 3212
rect 14708 3172 14717 3212
rect 14899 3172 14908 3212
rect 14948 3172 15724 3212
rect 15764 3172 15773 3212
rect 16771 3172 16780 3212
rect 16820 3172 17260 3212
rect 17300 3172 17309 3212
rect 17395 3172 17404 3212
rect 17444 3172 21484 3212
rect 21524 3172 21533 3212
rect 21907 3172 21916 3212
rect 21956 3172 22444 3212
rect 22484 3172 22493 3212
rect 28435 3172 28444 3212
rect 28484 3172 28684 3212
rect 28724 3172 28733 3212
rect 29875 3172 29884 3212
rect 29924 3172 30316 3212
rect 30356 3172 30365 3212
rect 30643 3172 30652 3212
rect 30692 3172 31660 3212
rect 31700 3172 31709 3212
rect 31891 3172 31900 3212
rect 31940 3172 32524 3212
rect 32564 3172 32573 3212
rect 32659 3172 32668 3212
rect 32708 3172 33004 3212
rect 33044 3172 33053 3212
rect 33139 3172 33148 3212
rect 33188 3172 33388 3212
rect 33428 3172 33437 3212
rect 34003 3172 34012 3212
rect 34052 3172 34348 3212
rect 34388 3172 34397 3212
rect 35011 3172 35020 3212
rect 35060 3172 35260 3212
rect 35300 3172 35309 3212
rect 35539 3172 35548 3212
rect 35588 3172 35692 3212
rect 35732 3172 35741 3212
rect 36019 3172 36028 3212
rect 36068 3172 36076 3212
rect 36116 3172 36199 3212
rect 0 3128 90 3148
rect 36268 3128 36308 3256
rect 36451 3172 36460 3212
rect 36500 3172 36700 3212
rect 36740 3172 36749 3212
rect 37459 3172 37468 3212
rect 37508 3172 37516 3212
rect 37556 3172 37639 3212
rect 41609 3172 41731 3212
rect 41780 3172 41789 3212
rect 50554 3172 50563 3212
rect 50603 3172 50860 3212
rect 50900 3172 51235 3212
rect 51275 3172 51436 3212
rect 51476 3172 51485 3212
rect 51667 3172 51676 3212
rect 51716 3172 51725 3212
rect 50572 3128 50612 3172
rect 0 3088 27956 3128
rect 28003 3088 28012 3128
rect 28052 3088 36308 3128
rect 50188 3088 50612 3128
rect 51676 3128 51716 3172
rect 53190 3128 53280 3148
rect 51676 3088 53280 3128
rect 0 3068 90 3088
rect 27916 3044 27956 3088
rect 4919 3004 4928 3044
rect 4968 3004 5010 3044
rect 5050 3004 5092 3044
rect 5132 3004 5174 3044
rect 5214 3004 5256 3044
rect 5296 3004 5305 3044
rect 14563 3004 14572 3044
rect 14612 3004 19852 3044
rect 19892 3004 19901 3044
rect 20039 3004 20048 3044
rect 20088 3004 20130 3044
rect 20170 3004 20212 3044
rect 20252 3004 20294 3044
rect 20334 3004 20376 3044
rect 20416 3004 20425 3044
rect 22723 3004 22732 3044
rect 22772 3004 27860 3044
rect 27916 3004 33100 3044
rect 33140 3004 33149 3044
rect 35159 3004 35168 3044
rect 35208 3004 35250 3044
rect 35290 3004 35332 3044
rect 35372 3004 35414 3044
rect 35454 3004 35496 3044
rect 35536 3004 35545 3044
rect 27820 2960 27860 3004
rect 6979 2920 6988 2960
rect 7028 2920 21772 2960
rect 21812 2920 21821 2960
rect 22435 2920 22444 2960
rect 22484 2920 24556 2960
rect 24596 2920 24605 2960
rect 27820 2920 30260 2960
rect 31651 2920 31660 2960
rect 31700 2920 49516 2960
rect 49556 2920 49565 2960
rect 30220 2876 30260 2920
rect 50188 2876 50228 3088
rect 53190 3068 53280 3088
rect 50279 3004 50288 3044
rect 50328 3004 50370 3044
rect 50410 3004 50452 3044
rect 50492 3004 50534 3044
rect 50574 3004 50616 3044
rect 50656 3004 50665 3044
rect 11788 2836 14188 2876
rect 14228 2836 14237 2876
rect 14323 2836 14332 2876
rect 14372 2836 21332 2876
rect 0 2792 90 2812
rect 0 2752 1420 2792
rect 1460 2752 1469 2792
rect 0 2732 90 2752
rect 11788 2624 11828 2836
rect 13132 2752 15436 2792
rect 15476 2752 15485 2792
rect 18451 2752 18460 2792
rect 18500 2752 20620 2792
rect 20660 2752 20669 2792
rect 20755 2752 20764 2792
rect 20804 2752 20948 2792
rect 13132 2624 13172 2752
rect 20908 2708 20948 2752
rect 21292 2708 21332 2836
rect 21484 2836 23116 2876
rect 23156 2836 23165 2876
rect 23251 2836 23260 2876
rect 23300 2836 26860 2876
rect 26900 2836 26909 2876
rect 30220 2836 37708 2876
rect 37748 2836 37757 2876
rect 49978 2836 49987 2876
rect 50027 2836 50228 2876
rect 21484 2792 21524 2836
rect 53190 2792 53280 2812
rect 21379 2752 21388 2792
rect 21428 2752 21524 2792
rect 23731 2752 23740 2792
rect 23780 2752 26476 2792
rect 26516 2752 26525 2792
rect 26659 2752 26668 2792
rect 26708 2752 30260 2792
rect 30307 2752 30316 2792
rect 30356 2752 42412 2792
rect 42452 2752 42461 2792
rect 44707 2752 44716 2792
rect 44756 2752 51092 2792
rect 52051 2752 52060 2792
rect 52100 2752 53280 2792
rect 30220 2708 30260 2752
rect 14092 2668 16204 2708
rect 16244 2668 16253 2708
rect 19939 2668 19948 2708
rect 19988 2668 20660 2708
rect 20908 2668 21236 2708
rect 21292 2668 24460 2708
rect 24500 2668 24509 2708
rect 24844 2668 28012 2708
rect 28052 2668 28061 2708
rect 30220 2668 31468 2708
rect 31508 2668 31517 2708
rect 31564 2668 39148 2708
rect 39188 2668 39197 2708
rect 14092 2624 14132 2668
rect 20620 2624 20660 2668
rect 21196 2624 21236 2668
rect 24844 2624 24884 2668
rect 31564 2624 31604 2668
rect 51052 2624 51092 2752
rect 53190 2732 53280 2752
rect 739 2584 748 2624
rect 788 2584 2188 2624
rect 2228 2584 2237 2624
rect 7180 2584 7276 2624
rect 7316 2584 7325 2624
rect 11779 2584 11788 2624
rect 11828 2584 11837 2624
rect 13123 2584 13132 2624
rect 13172 2584 13181 2624
rect 14083 2584 14092 2624
rect 14132 2584 14141 2624
rect 14659 2584 14668 2624
rect 14708 2584 15820 2624
rect 15860 2584 15869 2624
rect 18089 2584 18220 2624
rect 18260 2584 18269 2624
rect 18595 2584 18604 2624
rect 18644 2584 19276 2624
rect 19316 2584 19325 2624
rect 19459 2584 19468 2624
rect 19508 2584 20524 2624
rect 20564 2584 20573 2624
rect 20620 2584 20908 2624
rect 20948 2584 20957 2624
rect 21196 2584 21868 2624
rect 21908 2584 21917 2624
rect 23011 2584 23020 2624
rect 23060 2584 23191 2624
rect 23299 2584 23308 2624
rect 23348 2584 23500 2624
rect 23540 2584 23549 2624
rect 23683 2584 23692 2624
rect 23732 2584 24076 2624
rect 24116 2584 24125 2624
rect 24547 2584 24556 2624
rect 24596 2584 24652 2624
rect 24692 2584 24727 2624
rect 24787 2584 24796 2624
rect 24836 2584 24884 2624
rect 24931 2584 24940 2624
rect 24980 2584 25111 2624
rect 25219 2584 25228 2624
rect 25268 2584 25612 2624
rect 25652 2584 25661 2624
rect 25891 2584 25900 2624
rect 25940 2584 27052 2624
rect 27092 2584 27101 2624
rect 27235 2584 27244 2624
rect 27284 2584 28396 2624
rect 28436 2584 28445 2624
rect 28649 2584 28780 2624
rect 28820 2584 28829 2624
rect 29059 2584 29068 2624
rect 29108 2584 31604 2624
rect 31651 2584 31660 2624
rect 31700 2584 33388 2624
rect 33428 2584 33437 2624
rect 34121 2584 34252 2624
rect 34292 2584 34301 2624
rect 34505 2584 34540 2624
rect 34580 2584 34636 2624
rect 34676 2584 34685 2624
rect 36259 2584 36268 2624
rect 36308 2584 39532 2624
rect 39572 2584 39581 2624
rect 39715 2584 39724 2624
rect 39764 2584 40012 2624
rect 40052 2584 40061 2624
rect 49027 2584 49036 2624
rect 49076 2584 49324 2624
rect 49364 2584 49612 2624
rect 49652 2584 49708 2624
rect 49748 2584 49900 2624
rect 49940 2584 49949 2624
rect 50057 2584 50188 2624
rect 50228 2584 50476 2624
rect 50516 2584 50764 2624
rect 50804 2584 50813 2624
rect 51043 2584 51052 2624
rect 51092 2584 51101 2624
rect 51427 2584 51436 2624
rect 51476 2584 51485 2624
rect 51811 2584 51820 2624
rect 51860 2584 52108 2624
rect 52148 2584 52157 2624
rect 0 2456 90 2476
rect 0 2416 1420 2456
rect 1460 2416 1469 2456
rect 2419 2416 2428 2456
rect 2468 2416 4780 2456
rect 4820 2416 4829 2456
rect 0 2396 90 2416
rect 7180 2372 7220 2584
rect 49036 2540 49076 2584
rect 51436 2540 51476 2584
rect 7507 2500 7516 2540
rect 7556 2500 49076 2540
rect 49411 2500 49420 2540
rect 49460 2500 51476 2540
rect 51667 2500 51676 2540
rect 51716 2500 52724 2540
rect 52684 2456 52724 2500
rect 53190 2456 53280 2476
rect 12019 2416 12028 2456
rect 12068 2416 13268 2456
rect 13363 2416 13372 2456
rect 13412 2416 14804 2456
rect 14899 2416 14908 2456
rect 14948 2416 14957 2456
rect 18835 2416 18844 2456
rect 18884 2416 20852 2456
rect 21139 2416 21148 2456
rect 21188 2416 22924 2456
rect 22964 2416 22973 2456
rect 23107 2416 23116 2456
rect 23156 2416 24172 2456
rect 24212 2416 24221 2456
rect 24307 2416 24316 2456
rect 24356 2416 25036 2456
rect 25076 2416 25085 2456
rect 25171 2416 25180 2456
rect 25220 2416 25420 2456
rect 25460 2416 25469 2456
rect 25843 2416 25852 2456
rect 25892 2416 27188 2456
rect 27283 2416 27292 2456
rect 27332 2416 28532 2456
rect 28627 2416 28636 2456
rect 28676 2416 28916 2456
rect 29011 2416 29020 2456
rect 29060 2416 30316 2456
rect 30356 2416 30365 2456
rect 33619 2416 33628 2456
rect 33668 2416 33716 2456
rect 2668 2332 7220 2372
rect 0 2120 90 2140
rect 2668 2120 2708 2332
rect 3679 2248 3688 2288
rect 3728 2248 3770 2288
rect 3810 2248 3852 2288
rect 3892 2248 3934 2288
rect 3974 2248 4016 2288
rect 4056 2248 4065 2288
rect 13228 2204 13268 2416
rect 14764 2288 14804 2416
rect 14908 2372 14948 2416
rect 14908 2332 20428 2372
rect 20468 2332 20477 2372
rect 20812 2288 20852 2416
rect 27148 2372 27188 2416
rect 28492 2372 28532 2416
rect 28876 2372 28916 2416
rect 21091 2332 21100 2372
rect 21140 2332 25652 2372
rect 25699 2332 25708 2372
rect 25748 2332 27052 2372
rect 27092 2332 27101 2372
rect 27148 2332 28396 2372
rect 28436 2332 28445 2372
rect 28492 2332 28780 2372
rect 28820 2332 28829 2372
rect 28876 2332 29836 2372
rect 29876 2332 29885 2372
rect 25612 2288 25652 2332
rect 14764 2248 18412 2288
rect 18452 2248 18461 2288
rect 18799 2248 18808 2288
rect 18848 2248 18890 2288
rect 18930 2248 18972 2288
rect 19012 2248 19054 2288
rect 19094 2248 19136 2288
rect 19176 2248 19185 2288
rect 20812 2248 23020 2288
rect 23060 2248 23069 2288
rect 23203 2248 23212 2288
rect 23252 2248 25364 2288
rect 25612 2248 31892 2288
rect 25324 2204 25364 2248
rect 2755 2164 2764 2204
rect 2804 2164 12980 2204
rect 13228 2164 20908 2204
rect 20948 2164 20957 2204
rect 21004 2164 24308 2204
rect 0 2080 2708 2120
rect 12940 2120 12980 2164
rect 12940 2080 19468 2120
rect 19508 2080 19517 2120
rect 0 2060 90 2080
rect 8899 1996 8908 2036
rect 8948 1996 20620 2036
rect 20660 1996 20669 2036
rect 21004 1952 21044 2164
rect 24268 2120 24308 2164
rect 24748 2164 25228 2204
rect 25268 2164 25277 2204
rect 25324 2164 31124 2204
rect 24748 2120 24788 2164
rect 21859 2080 21868 2120
rect 21908 2080 24212 2120
rect 24268 2080 24788 2120
rect 25027 2080 25036 2120
rect 25076 2080 26996 2120
rect 21187 1996 21196 2036
rect 21236 1996 23444 2036
rect 23404 1952 23444 1996
rect 24172 1952 24212 2080
rect 24835 1996 24844 2036
rect 24884 1996 25364 2036
rect 25324 1952 25364 1996
rect 26956 1952 26996 2080
rect 29347 1996 29356 2036
rect 29396 1996 30740 2036
rect 30700 1952 30740 1996
rect 31084 1952 31124 2164
rect 31852 1952 31892 2248
rect 33676 1952 33716 2416
rect 34444 2416 34492 2456
rect 34532 2416 34541 2456
rect 34828 2416 34876 2456
rect 34916 2416 34925 2456
rect 37603 2416 37612 2456
rect 37652 2416 39292 2456
rect 39332 2416 39341 2456
rect 39427 2416 39436 2456
rect 39476 2416 39772 2456
rect 39812 2416 39821 2456
rect 51283 2416 51292 2456
rect 51332 2416 52588 2456
rect 52628 2416 52637 2456
rect 52684 2416 53280 2456
rect 33919 2248 33928 2288
rect 33968 2248 34010 2288
rect 34050 2248 34092 2288
rect 34132 2248 34174 2288
rect 34214 2248 34256 2288
rect 34296 2248 34305 2288
rect 34444 1952 34484 2416
rect 34828 1952 34868 2416
rect 53190 2396 53280 2416
rect 49039 2248 49048 2288
rect 49088 2248 49130 2288
rect 49170 2248 49212 2288
rect 49252 2248 49294 2288
rect 49334 2248 49376 2288
rect 49416 2248 49425 2288
rect 53190 2120 53280 2140
rect 34915 2080 34924 2120
rect 34964 2080 39572 2120
rect 42403 2080 42412 2120
rect 42452 2080 50420 2120
rect 52051 2080 52060 2120
rect 52100 2080 53280 2120
rect 39532 2036 39572 2080
rect 36844 1996 37516 2036
rect 37556 1996 37565 2036
rect 37996 1996 39436 2036
rect 39476 1996 39485 2036
rect 39532 1996 39956 2036
rect 40003 1996 40012 2036
rect 40052 1996 40724 2036
rect 36844 1952 36884 1996
rect 37996 1952 38036 1996
rect 39916 1952 39956 1996
rect 40684 1952 40724 1996
rect 50380 1952 50420 2080
rect 53190 2060 53280 2080
rect 9283 1912 9292 1952
rect 9332 1912 21044 1952
rect 21475 1912 21484 1952
rect 21524 1912 23020 1952
rect 23060 1912 23069 1952
rect 23395 1912 23404 1952
rect 23444 1912 23453 1952
rect 23779 1912 23788 1952
rect 23828 1912 23837 1952
rect 24163 1912 24172 1952
rect 24212 1912 24221 1952
rect 24425 1912 24556 1952
rect 24596 1912 24605 1952
rect 24931 1912 24940 1952
rect 24980 1912 24989 1952
rect 25315 1912 25324 1952
rect 25364 1912 25373 1952
rect 25507 1912 25516 1952
rect 25556 1912 25708 1952
rect 25748 1912 25757 1952
rect 25961 1912 26092 1952
rect 26132 1912 26141 1952
rect 26345 1912 26476 1952
rect 26516 1912 26525 1952
rect 26729 1912 26860 1952
rect 26900 1912 26909 1952
rect 26956 1912 27244 1952
rect 27284 1912 27293 1952
rect 27619 1912 27628 1952
rect 27668 1912 27677 1952
rect 27881 1912 28012 1952
rect 28052 1912 28061 1952
rect 28265 1912 28396 1952
rect 28436 1912 28445 1952
rect 28771 1912 28780 1952
rect 28820 1912 28828 1952
rect 28868 1912 28951 1952
rect 29155 1912 29164 1952
rect 29204 1912 29335 1952
rect 29539 1912 29548 1952
rect 29588 1912 29597 1952
rect 29827 1912 29836 1952
rect 29876 1912 29932 1952
rect 29972 1912 30007 1952
rect 30185 1912 30316 1952
rect 30356 1912 30365 1952
rect 30691 1912 30700 1952
rect 30740 1912 30749 1952
rect 31075 1912 31084 1952
rect 31124 1912 31133 1952
rect 31337 1912 31468 1952
rect 31508 1912 31517 1952
rect 31843 1912 31852 1952
rect 31892 1912 31901 1952
rect 32105 1912 32236 1952
rect 32276 1912 32285 1952
rect 32489 1912 32524 1952
rect 32564 1912 32620 1952
rect 32660 1912 32669 1952
rect 32873 1912 33004 1952
rect 33044 1912 33053 1952
rect 33257 1912 33388 1952
rect 33428 1912 33437 1952
rect 33676 1912 33772 1952
rect 33812 1912 33821 1952
rect 34147 1912 34156 1952
rect 34196 1912 34348 1952
rect 34388 1912 34397 1952
rect 34444 1912 34483 1952
rect 34523 1912 34532 1952
rect 34828 1912 34867 1952
rect 34907 1912 34916 1952
rect 35011 1912 35020 1952
rect 35060 1912 35308 1952
rect 35348 1912 35357 1952
rect 35561 1912 35692 1952
rect 35732 1912 35741 1952
rect 35945 1912 36076 1952
rect 36116 1912 36125 1952
rect 36329 1912 36460 1952
rect 36500 1912 36509 1952
rect 36835 1912 36844 1952
rect 36884 1912 36893 1952
rect 37219 1912 37228 1952
rect 37268 1912 37460 1952
rect 37603 1912 37612 1952
rect 37652 1912 37783 1952
rect 37987 1912 37996 1952
rect 38036 1912 38045 1952
rect 38249 1912 38380 1952
rect 38420 1912 38429 1952
rect 38755 1912 38764 1952
rect 38804 1912 38813 1952
rect 39017 1912 39148 1952
rect 39188 1912 39197 1952
rect 39401 1912 39532 1952
rect 39572 1912 39581 1952
rect 39907 1912 39916 1952
rect 39956 1912 39965 1952
rect 40169 1912 40300 1952
rect 40340 1912 40349 1952
rect 40675 1912 40684 1952
rect 40724 1912 40733 1952
rect 40937 1912 41068 1952
rect 41108 1912 41117 1952
rect 41321 1912 41452 1952
rect 41492 1912 41501 1952
rect 41705 1912 41836 1952
rect 41876 1912 41885 1952
rect 42089 1912 42220 1952
rect 42260 1912 42269 1952
rect 42473 1912 42604 1952
rect 42644 1912 42653 1952
rect 49507 1912 49516 1952
rect 49556 1912 49996 1952
rect 50036 1912 50045 1952
rect 50371 1912 50380 1952
rect 50420 1912 50429 1952
rect 50860 1912 51052 1952
rect 51092 1912 51101 1952
rect 51427 1912 51436 1952
rect 51476 1912 51628 1952
rect 51668 1912 51820 1952
rect 51860 1912 51869 1952
rect 23788 1868 23828 1912
rect 24940 1868 24980 1912
rect 27628 1868 27668 1912
rect 29548 1868 29588 1912
rect 3523 1828 3532 1868
rect 3572 1828 18220 1868
rect 18260 1828 18269 1868
rect 18403 1828 18412 1868
rect 18452 1828 21772 1868
rect 21812 1828 21821 1868
rect 22051 1828 22060 1868
rect 22100 1828 23828 1868
rect 24067 1828 24076 1868
rect 24116 1828 24980 1868
rect 25411 1828 25420 1868
rect 25460 1828 27668 1868
rect 28675 1828 28684 1868
rect 28724 1828 29588 1868
rect 37420 1868 37460 1912
rect 38764 1868 38804 1912
rect 50860 1868 50900 1912
rect 37420 1828 37804 1868
rect 37844 1828 37853 1868
rect 37987 1828 37996 1868
rect 38036 1828 38804 1868
rect 49228 1828 50188 1868
rect 50228 1828 50860 1868
rect 50900 1828 50909 1868
rect 51148 1828 52436 1868
rect 0 1784 90 1804
rect 49228 1784 49268 1828
rect 51148 1784 51188 1828
rect 52396 1784 52436 1828
rect 53190 1784 53280 1804
rect 0 1744 1420 1784
rect 1460 1744 1469 1784
rect 4771 1744 4780 1784
rect 4820 1744 48652 1784
rect 48692 1744 48940 1784
rect 48980 1744 49228 1784
rect 49268 1744 49277 1784
rect 49507 1744 49516 1784
rect 49556 1744 49708 1784
rect 49748 1744 49804 1784
rect 49844 1744 49908 1784
rect 50227 1744 50236 1784
rect 50276 1744 51188 1784
rect 51283 1744 51292 1784
rect 51332 1744 52300 1784
rect 52340 1744 52349 1784
rect 52396 1744 53280 1784
rect 0 1724 90 1744
rect 53190 1724 53280 1744
rect 7180 1660 10100 1700
rect 18403 1660 18412 1700
rect 18452 1660 22540 1700
rect 22580 1660 22589 1700
rect 22649 1660 22732 1700
rect 22772 1660 22780 1700
rect 22820 1660 22829 1700
rect 23107 1660 23116 1700
rect 23156 1660 23164 1700
rect 23204 1660 23287 1700
rect 23417 1660 23500 1700
rect 23540 1660 23548 1700
rect 23588 1660 23597 1700
rect 23801 1660 23884 1700
rect 23924 1660 23932 1700
rect 23972 1660 23981 1700
rect 24185 1660 24268 1700
rect 24308 1660 24316 1700
rect 24356 1660 24365 1700
rect 24569 1660 24652 1700
rect 24692 1660 24700 1700
rect 24740 1660 24749 1700
rect 24953 1660 25036 1700
rect 25076 1660 25084 1700
rect 25124 1660 25133 1700
rect 25337 1660 25420 1700
rect 25460 1660 25468 1700
rect 25508 1660 25517 1700
rect 25721 1660 25804 1700
rect 25844 1660 25852 1700
rect 25892 1660 25901 1700
rect 26105 1660 26188 1700
rect 26228 1660 26236 1700
rect 26276 1660 26285 1700
rect 26489 1660 26572 1700
rect 26612 1660 26620 1700
rect 26660 1660 26669 1700
rect 26873 1660 26956 1700
rect 26996 1660 27004 1700
rect 27044 1660 27053 1700
rect 27257 1660 27340 1700
rect 27380 1660 27388 1700
rect 27428 1660 27437 1700
rect 27641 1660 27724 1700
rect 27764 1660 27772 1700
rect 27812 1660 27821 1700
rect 28025 1660 28108 1700
rect 28148 1660 28156 1700
rect 28196 1660 28205 1700
rect 28409 1660 28492 1700
rect 28532 1660 28540 1700
rect 28580 1660 28589 1700
rect 28793 1660 28876 1700
rect 28916 1660 28924 1700
rect 28964 1660 28973 1700
rect 29177 1660 29260 1700
rect 29300 1660 29308 1700
rect 29348 1660 29357 1700
rect 29561 1660 29644 1700
rect 29684 1660 29692 1700
rect 29732 1660 29741 1700
rect 29945 1660 30028 1700
rect 30068 1660 30076 1700
rect 30116 1660 30125 1700
rect 30329 1660 30412 1700
rect 30452 1660 30460 1700
rect 30500 1660 30509 1700
rect 30713 1660 30796 1700
rect 30836 1660 30844 1700
rect 30884 1660 30893 1700
rect 31097 1660 31180 1700
rect 31220 1660 31228 1700
rect 31268 1660 31277 1700
rect 31481 1660 31564 1700
rect 31604 1660 31612 1700
rect 31652 1660 31661 1700
rect 31865 1660 31948 1700
rect 31988 1660 31996 1700
rect 32036 1660 32045 1700
rect 32249 1660 32332 1700
rect 32372 1660 32380 1700
rect 32420 1660 32429 1700
rect 32633 1660 32716 1700
rect 32756 1660 32764 1700
rect 32804 1660 32813 1700
rect 32988 1660 33100 1700
rect 33140 1660 33148 1700
rect 33188 1660 33197 1700
rect 33401 1660 33484 1700
rect 33524 1660 33532 1700
rect 33572 1660 33581 1700
rect 33785 1660 33868 1700
rect 33908 1660 33916 1700
rect 33956 1660 33965 1700
rect 34169 1660 34252 1700
rect 34292 1660 34300 1700
rect 34340 1660 34349 1700
rect 34553 1660 34636 1700
rect 34676 1660 34684 1700
rect 34724 1660 34733 1700
rect 34937 1660 35020 1700
rect 35060 1660 35068 1700
rect 35108 1660 35117 1700
rect 35443 1660 35452 1700
rect 35492 1660 35596 1700
rect 35636 1660 35645 1700
rect 35779 1660 35788 1700
rect 35828 1660 35836 1700
rect 35876 1660 35959 1700
rect 36089 1660 36172 1700
rect 36212 1660 36220 1700
rect 36260 1660 36269 1700
rect 36473 1660 36556 1700
rect 36596 1660 36604 1700
rect 36644 1660 36653 1700
rect 36857 1660 36940 1700
rect 36980 1660 36988 1700
rect 37028 1660 37037 1700
rect 37241 1660 37324 1700
rect 37364 1660 37372 1700
rect 37412 1660 37421 1700
rect 37625 1660 37708 1700
rect 37748 1660 37756 1700
rect 37796 1660 37805 1700
rect 38009 1660 38092 1700
rect 38132 1660 38140 1700
rect 38180 1660 38189 1700
rect 38393 1660 38476 1700
rect 38516 1660 38524 1700
rect 38564 1660 38573 1700
rect 38777 1660 38860 1700
rect 38900 1660 38908 1700
rect 38948 1660 38957 1700
rect 39161 1660 39244 1700
rect 39284 1660 39292 1700
rect 39332 1660 39341 1700
rect 39545 1660 39628 1700
rect 39668 1660 39676 1700
rect 39716 1660 39725 1700
rect 39929 1660 40012 1700
rect 40052 1660 40060 1700
rect 40100 1660 40109 1700
rect 40313 1660 40396 1700
rect 40436 1660 40444 1700
rect 40484 1660 40493 1700
rect 40697 1660 40780 1700
rect 40820 1660 40828 1700
rect 40868 1660 40877 1700
rect 41081 1660 41164 1700
rect 41204 1660 41212 1700
rect 41252 1660 41261 1700
rect 41465 1660 41548 1700
rect 41588 1660 41596 1700
rect 41636 1660 41645 1700
rect 41849 1660 41932 1700
rect 41972 1660 41980 1700
rect 42020 1660 42029 1700
rect 42233 1660 42316 1700
rect 42356 1660 42364 1700
rect 42404 1660 42413 1700
rect 50611 1660 50620 1700
rect 50660 1660 50708 1700
rect 7180 1616 7220 1660
rect 4291 1576 4300 1616
rect 4340 1576 7220 1616
rect 4919 1492 4928 1532
rect 4968 1492 5010 1532
rect 5050 1492 5092 1532
rect 5132 1492 5174 1532
rect 5214 1492 5256 1532
rect 5296 1492 5305 1532
rect 0 1448 90 1468
rect 10060 1448 10100 1660
rect 50668 1616 50708 1660
rect 18412 1576 23692 1616
rect 23732 1576 23741 1616
rect 24163 1576 24172 1616
rect 24212 1576 29492 1616
rect 29539 1576 29548 1616
rect 29588 1576 35636 1616
rect 35971 1576 35980 1616
rect 36020 1576 39532 1616
rect 39572 1576 39581 1616
rect 50668 1576 51916 1616
rect 51956 1576 51965 1616
rect 18412 1448 18452 1576
rect 29452 1532 29492 1576
rect 35596 1532 35636 1576
rect 20039 1492 20048 1532
rect 20088 1492 20130 1532
rect 20170 1492 20212 1532
rect 20252 1492 20294 1532
rect 20334 1492 20376 1532
rect 20416 1492 20425 1532
rect 20611 1492 20620 1532
rect 20660 1492 24308 1532
rect 24451 1492 24460 1532
rect 24500 1492 29356 1532
rect 29396 1492 29405 1532
rect 29452 1492 34924 1532
rect 34964 1492 34973 1532
rect 35159 1492 35168 1532
rect 35208 1492 35250 1532
rect 35290 1492 35332 1532
rect 35372 1492 35414 1532
rect 35454 1492 35496 1532
rect 35536 1492 35545 1532
rect 35596 1492 37900 1532
rect 37940 1492 37949 1532
rect 50279 1492 50288 1532
rect 50328 1492 50370 1532
rect 50410 1492 50452 1532
rect 50492 1492 50534 1532
rect 50574 1492 50616 1532
rect 50656 1492 50665 1532
rect 24268 1448 24308 1492
rect 53190 1448 53280 1468
rect 0 1408 1420 1448
rect 1460 1408 1469 1448
rect 10060 1408 18452 1448
rect 22915 1408 22924 1448
rect 22964 1408 23060 1448
rect 24268 1408 25900 1448
rect 25940 1408 25949 1448
rect 52579 1408 52588 1448
rect 52628 1408 53280 1448
rect 0 1388 90 1408
rect 23020 1280 23060 1408
rect 53190 1388 53280 1408
rect 23020 1240 29068 1280
rect 29108 1240 29117 1280
rect 0 1112 90 1132
rect 53190 1112 53280 1132
rect 0 1072 1420 1112
rect 1460 1072 1469 1112
rect 51907 1072 51916 1112
rect 51956 1072 53280 1112
rect 0 1052 90 1072
rect 53190 1052 53280 1072
rect 0 776 90 796
rect 53190 776 53280 796
rect 0 736 748 776
rect 788 736 797 776
rect 52291 736 52300 776
rect 52340 736 53280 776
rect 0 716 90 736
rect 53190 716 53280 736
rect 21571 316 21580 356
rect 21620 316 36268 356
rect 36308 316 36317 356
rect 9667 232 9676 272
rect 9716 232 24748 272
rect 24788 232 24797 272
rect 25603 232 25612 272
rect 25652 232 46156 272
rect 46196 232 46205 272
rect 21283 148 21292 188
rect 21332 148 23060 188
rect 23779 148 23788 188
rect 23828 148 45772 188
rect 45812 148 45821 188
rect 23020 104 23060 148
rect 23020 64 45388 104
rect 45428 64 45437 104
<< via2 >>
rect 844 11152 884 11192
rect 50956 11152 50996 11192
rect 23596 10816 23636 10856
rect 51052 10816 51092 10856
rect 4928 10564 4968 10604
rect 5010 10564 5050 10604
rect 5092 10564 5132 10604
rect 5174 10564 5214 10604
rect 5256 10564 5296 10604
rect 20048 10564 20088 10604
rect 20130 10564 20170 10604
rect 20212 10564 20252 10604
rect 20294 10564 20334 10604
rect 20376 10564 20416 10604
rect 35168 10564 35208 10604
rect 35250 10564 35290 10604
rect 35332 10564 35372 10604
rect 35414 10564 35454 10604
rect 35496 10564 35536 10604
rect 39148 10564 39188 10604
rect 46156 10564 46196 10604
rect 50288 10564 50328 10604
rect 50370 10564 50410 10604
rect 50452 10564 50492 10604
rect 50534 10564 50574 10604
rect 50616 10564 50656 10604
rect 14284 10480 14324 10520
rect 36940 10480 36980 10520
rect 44908 10480 44948 10520
rect 51244 10480 51284 10520
rect 51436 10480 51476 10520
rect 1612 10396 1652 10436
rect 4108 10396 4148 10436
rect 6604 10396 6644 10436
rect 9100 10396 9140 10436
rect 11596 10396 11636 10436
rect 14092 10396 14132 10436
rect 16588 10396 16628 10436
rect 19084 10396 19124 10436
rect 21580 10396 21620 10436
rect 24076 10396 24116 10436
rect 26572 10396 26612 10436
rect 29068 10396 29108 10436
rect 31564 10396 31604 10436
rect 34060 10396 34100 10436
rect 39052 10396 39092 10436
rect 41548 10396 41588 10436
rect 44044 10396 44084 10436
rect 46540 10396 46580 10436
rect 49036 10396 49076 10436
rect 51052 10396 51092 10436
rect 51532 10396 51572 10436
rect 24172 10312 24212 10352
rect 26668 10228 26708 10268
rect 36748 10228 36788 10268
rect 44620 10228 44660 10268
rect 1900 10144 1940 10184
rect 4396 10144 4436 10184
rect 6892 10144 6932 10184
rect 9388 10144 9428 10184
rect 13612 10144 13652 10184
rect 14380 10144 14420 10184
rect 18412 10144 18452 10184
rect 20812 10144 20852 10184
rect 23116 10144 23156 10184
rect 25228 10144 25268 10184
rect 27820 10144 27860 10184
rect 29356 10144 29396 10184
rect 36556 10144 36596 10184
rect 39148 10144 39188 10184
rect 43372 10144 43412 10184
rect 46636 10144 46676 10184
rect 48172 10144 48212 10184
rect 48940 10144 48980 10184
rect 50092 10144 50132 10184
rect 51052 10144 51092 10184
rect 51436 10144 51476 10184
rect 51628 10144 51668 10184
rect 15436 10060 15476 10100
rect 26572 10060 26612 10100
rect 27724 10060 27764 10100
rect 30700 10060 30740 10100
rect 43948 10060 43988 10100
rect 47500 10060 47540 10100
rect 51532 10060 51572 10100
rect 24268 9976 24308 10016
rect 26956 9976 26996 10016
rect 29164 9976 29204 10016
rect 37996 9976 38036 10016
rect 51052 9976 51092 10016
rect 28876 9892 28916 9932
rect 46348 9892 46388 9932
rect 50380 9892 50420 9932
rect 51436 9892 51476 9932
rect 3688 9808 3728 9848
rect 3770 9808 3810 9848
rect 3852 9808 3892 9848
rect 3934 9808 3974 9848
rect 4016 9808 4056 9848
rect 18808 9808 18848 9848
rect 18890 9808 18930 9848
rect 18972 9808 19012 9848
rect 19054 9808 19094 9848
rect 19136 9808 19176 9848
rect 19372 9808 19412 9848
rect 27724 9808 27764 9848
rect 27916 9808 27956 9848
rect 30028 9808 30068 9848
rect 33928 9808 33968 9848
rect 34010 9808 34050 9848
rect 34092 9808 34132 9848
rect 34174 9808 34214 9848
rect 34256 9808 34296 9848
rect 35020 9808 35060 9848
rect 38284 9808 38324 9848
rect 47500 9808 47540 9848
rect 49048 9808 49088 9848
rect 49130 9808 49170 9848
rect 49212 9808 49252 9848
rect 49294 9808 49334 9848
rect 49376 9808 49416 9848
rect 844 9724 884 9764
rect 9388 9724 9428 9764
rect 37900 9724 37940 9764
rect 38092 9724 38132 9764
rect 13612 9640 13652 9680
rect 14380 9640 14420 9680
rect 18412 9640 18452 9680
rect 20812 9640 20852 9680
rect 23116 9640 23156 9680
rect 24172 9640 24212 9680
rect 25228 9640 25268 9680
rect 26956 9640 26996 9680
rect 27820 9640 27860 9680
rect 29164 9640 29204 9680
rect 29356 9640 29396 9680
rect 43084 9640 43124 9680
rect 43372 9640 43412 9680
rect 43948 9640 43988 9680
rect 44908 9640 44948 9680
rect 46156 9640 46196 9680
rect 46636 9640 46676 9680
rect 48172 9640 48212 9680
rect 48940 9640 48980 9680
rect 6892 9556 6932 9596
rect 30028 9556 30068 9596
rect 43468 9556 43508 9596
rect 43852 9556 43892 9596
rect 47692 9556 47732 9596
rect 50956 9640 50996 9680
rect 51628 9640 51668 9680
rect 51532 9556 51572 9596
rect 14092 9472 14132 9512
rect 14284 9472 14324 9512
rect 18700 9472 18740 9512
rect 21292 9472 21332 9512
rect 23596 9472 23636 9512
rect 25612 9472 25652 9512
rect 26188 9472 26228 9512
rect 26668 9472 26708 9512
rect 28588 9472 28628 9512
rect 28876 9472 28916 9512
rect 29932 9472 29972 9512
rect 30220 9472 30260 9512
rect 38284 9472 38324 9512
rect 49996 9472 50036 9512
rect 50956 9472 50996 9512
rect 51628 9472 51668 9512
rect 15436 9388 15476 9428
rect 19372 9388 19412 9428
rect 23788 9388 23828 9428
rect 23980 9388 24020 9428
rect 28396 9388 28436 9428
rect 30700 9388 30740 9428
rect 42700 9388 42740 9428
rect 44140 9388 44180 9428
rect 46156 9388 46196 9428
rect 47212 9388 47252 9428
rect 48460 9388 48500 9428
rect 49612 9388 49652 9428
rect 4396 9304 4436 9344
rect 27916 9304 27956 9344
rect 43564 9304 43604 9344
rect 48076 9304 48116 9344
rect 1900 9220 1940 9260
rect 20140 9220 20180 9260
rect 26380 9220 26420 9260
rect 28588 9220 28628 9260
rect 38284 9220 38324 9260
rect 44620 9220 44660 9260
rect 47212 9220 47252 9260
rect 48940 9220 48980 9260
rect 50092 9220 50132 9260
rect 20524 9136 20564 9176
rect 20812 9136 20852 9176
rect 28300 9136 28340 9176
rect 4928 9052 4968 9092
rect 5010 9052 5050 9092
rect 5092 9052 5132 9092
rect 5174 9052 5214 9092
rect 5256 9052 5296 9092
rect 20048 9052 20088 9092
rect 20130 9052 20170 9092
rect 20212 9052 20252 9092
rect 20294 9052 20334 9092
rect 20376 9052 20416 9092
rect 28396 9052 28436 9092
rect 35020 9052 35060 9092
rect 35168 9052 35208 9092
rect 35250 9052 35290 9092
rect 35332 9052 35372 9092
rect 35414 9052 35454 9092
rect 35496 9052 35536 9092
rect 45964 9136 46004 9176
rect 46156 9136 46196 9176
rect 47308 9136 47348 9176
rect 44140 9052 44180 9092
rect 48844 9052 48884 9092
rect 50288 9052 50328 9092
rect 50370 9052 50410 9092
rect 50452 9052 50492 9092
rect 50534 9052 50574 9092
rect 50616 9052 50656 9092
rect 28108 8968 28148 9008
rect 29932 8968 29972 9008
rect 37996 8968 38036 9008
rect 44620 8968 44660 9008
rect 46156 8968 46196 9008
rect 748 8884 788 8924
rect 26188 8884 26228 8924
rect 26572 8884 26612 8924
rect 30220 8884 30260 8924
rect 47212 8884 47252 8924
rect 52684 9220 52724 9260
rect 1228 8800 1268 8840
rect 52684 8800 52724 8840
rect 43276 8716 43316 8756
rect 43564 8716 43604 8756
rect 46156 8716 46196 8756
rect 46348 8716 46388 8756
rect 1132 8632 1172 8672
rect 24268 8632 24308 8672
rect 26380 8632 26420 8672
rect 27340 8632 27380 8672
rect 27916 8632 27956 8672
rect 28108 8632 28148 8672
rect 33196 8632 33236 8672
rect 37996 8632 38036 8672
rect 46924 8632 46964 8672
rect 51820 8632 51860 8672
rect 53164 8632 53204 8672
rect 3688 8296 3728 8336
rect 3770 8296 3810 8336
rect 3852 8296 3892 8336
rect 3934 8296 3974 8336
rect 4016 8296 4056 8336
rect 18808 8296 18848 8336
rect 18890 8296 18930 8336
rect 18972 8296 19012 8336
rect 19054 8296 19094 8336
rect 19136 8296 19176 8336
rect 1324 8128 1364 8168
rect 1228 8044 1268 8084
rect 364 7960 404 8000
rect 33928 8296 33968 8336
rect 34010 8296 34050 8336
rect 34092 8296 34132 8336
rect 34174 8296 34214 8336
rect 34256 8296 34296 8336
rect 49048 8296 49088 8336
rect 49130 8296 49170 8336
rect 49212 8296 49252 8336
rect 49294 8296 49334 8336
rect 49376 8296 49416 8336
rect 23980 8128 24020 8168
rect 51628 8128 51668 8168
rect 53164 8128 53204 8168
rect 23884 8044 23924 8084
rect 38092 8044 38132 8084
rect 34828 7960 34868 8000
rect 34924 7876 34964 7916
rect 35308 7876 35348 7916
rect 21580 7792 21620 7832
rect 25708 7708 25748 7748
rect 33196 7708 33236 7748
rect 44236 7708 44276 7748
rect 38092 7624 38132 7664
rect 53164 7624 53204 7664
rect 4928 7540 4968 7580
rect 5010 7540 5050 7580
rect 5092 7540 5132 7580
rect 5174 7540 5214 7580
rect 5256 7540 5296 7580
rect 20048 7540 20088 7580
rect 20130 7540 20170 7580
rect 20212 7540 20252 7580
rect 20294 7540 20334 7580
rect 20376 7540 20416 7580
rect 35168 7540 35208 7580
rect 35250 7540 35290 7580
rect 35332 7540 35372 7580
rect 35414 7540 35454 7580
rect 35496 7540 35536 7580
rect 50288 7540 50328 7580
rect 50370 7540 50410 7580
rect 50452 7540 50492 7580
rect 50534 7540 50574 7580
rect 50616 7540 50656 7580
rect 52012 7540 52052 7580
rect 22924 7456 22964 7496
rect 53164 7456 53204 7496
rect 34828 7288 34868 7328
rect 460 7204 500 7244
rect 1228 7120 1268 7160
rect 10732 7120 10772 7160
rect 21580 7120 21620 7160
rect 23884 7120 23924 7160
rect 24172 7120 24212 7160
rect 51916 7120 51956 7160
rect 1036 7036 1076 7076
rect 19948 6952 19988 6992
rect 3688 6784 3728 6824
rect 3770 6784 3810 6824
rect 3852 6784 3892 6824
rect 3934 6784 3974 6824
rect 4016 6784 4056 6824
rect 18808 6784 18848 6824
rect 18890 6784 18930 6824
rect 18972 6784 19012 6824
rect 19054 6784 19094 6824
rect 19136 6784 19176 6824
rect 21580 6700 21620 6740
rect 51820 7036 51860 7076
rect 51436 6868 51476 6908
rect 33928 6784 33968 6824
rect 34010 6784 34050 6824
rect 34092 6784 34132 6824
rect 34174 6784 34214 6824
rect 34256 6784 34296 6824
rect 49048 6784 49088 6824
rect 49130 6784 49170 6824
rect 49212 6784 49252 6824
rect 49294 6784 49334 6824
rect 49376 6784 49416 6824
rect 1324 6616 1364 6656
rect 25708 6532 25748 6572
rect 1420 6448 1460 6488
rect 22732 6448 22772 6488
rect 22924 6448 22964 6488
rect 25804 6448 25844 6488
rect 35788 6448 35828 6488
rect 51820 6448 51860 6488
rect 268 6364 308 6404
rect 22924 6196 22964 6236
rect 47500 6196 47540 6236
rect 25804 6112 25844 6152
rect 4928 6028 4968 6068
rect 5010 6028 5050 6068
rect 5092 6028 5132 6068
rect 5174 6028 5214 6068
rect 5256 6028 5296 6068
rect 20048 6028 20088 6068
rect 20130 6028 20170 6068
rect 20212 6028 20252 6068
rect 20294 6028 20334 6068
rect 20376 6028 20416 6068
rect 35168 6028 35208 6068
rect 35250 6028 35290 6068
rect 35332 6028 35372 6068
rect 35414 6028 35454 6068
rect 35496 6028 35536 6068
rect 50288 6028 50328 6068
rect 50370 6028 50410 6068
rect 50452 6028 50492 6068
rect 50534 6028 50574 6068
rect 50616 6028 50656 6068
rect 52108 6028 52148 6068
rect 22732 5776 22772 5816
rect 35788 5776 35828 5816
rect 22924 5692 22964 5732
rect 21580 5608 21620 5648
rect 24172 5608 24212 5648
rect 27820 5608 27860 5648
rect 19948 5524 19988 5564
rect 10732 5440 10772 5480
rect 51916 5356 51956 5396
rect 3688 5272 3728 5312
rect 3770 5272 3810 5312
rect 3852 5272 3892 5312
rect 3934 5272 3974 5312
rect 4016 5272 4056 5312
rect 18808 5272 18848 5312
rect 18890 5272 18930 5312
rect 18972 5272 19012 5312
rect 19054 5272 19094 5312
rect 19136 5272 19176 5312
rect 33928 5272 33968 5312
rect 34010 5272 34050 5312
rect 34092 5272 34132 5312
rect 34174 5272 34214 5312
rect 34256 5272 34296 5312
rect 49048 5272 49088 5312
rect 49130 5272 49170 5312
rect 49212 5272 49252 5312
rect 49294 5272 49334 5312
rect 49376 5272 49416 5312
rect 1228 5188 1268 5228
rect 27820 5188 27860 5228
rect 1132 5104 1172 5144
rect 27916 5104 27956 5144
rect 1420 5020 1460 5060
rect 14668 4936 14708 4976
rect 18124 4936 18164 4976
rect 24172 4936 24212 4976
rect 51436 4936 51476 4976
rect 5452 4852 5492 4892
rect 51820 4852 51860 4892
rect 1036 4768 1076 4808
rect 5836 4768 5876 4808
rect 15340 4684 15380 4724
rect 15628 4684 15668 4724
rect 24844 4684 24884 4724
rect 25516 4684 25556 4724
rect 14668 4600 14708 4640
rect 17740 4600 17780 4640
rect 26092 4600 26132 4640
rect 4928 4516 4968 4556
rect 5010 4516 5050 4556
rect 5092 4516 5132 4556
rect 5174 4516 5214 4556
rect 5256 4516 5296 4556
rect 20048 4516 20088 4556
rect 20130 4516 20170 4556
rect 20212 4516 20252 4556
rect 20294 4516 20334 4556
rect 20376 4516 20416 4556
rect 35168 4516 35208 4556
rect 35250 4516 35290 4556
rect 35332 4516 35372 4556
rect 35414 4516 35454 4556
rect 35496 4516 35536 4556
rect 50288 4516 50328 4556
rect 50370 4516 50410 4556
rect 50452 4516 50492 4556
rect 50534 4516 50574 4556
rect 50616 4516 50656 4556
rect 364 4432 404 4472
rect 6220 4432 6260 4472
rect 24172 4432 24212 4472
rect 22828 4348 22868 4388
rect 27340 4348 27380 4388
rect 6604 4264 6644 4304
rect 11596 4180 11636 4220
rect 13708 4180 13748 4220
rect 16300 4180 16340 4220
rect 18508 4180 18548 4220
rect 18700 4180 18740 4220
rect 22924 4180 22964 4220
rect 460 4096 500 4136
rect 23308 4264 23348 4304
rect 32908 4264 32948 4304
rect 44236 4264 44276 4304
rect 16204 4096 16244 4136
rect 18316 4096 18356 4136
rect 19660 4096 19700 4136
rect 19852 4096 19892 4136
rect 28012 4096 28052 4136
rect 28204 4096 28244 4136
rect 35020 4096 35060 4136
rect 22636 4012 22676 4052
rect 14380 3928 14420 3968
rect 16876 3928 16916 3968
rect 18412 3928 18452 3968
rect 20716 3928 20756 3968
rect 12748 3844 12788 3884
rect 18604 3844 18644 3884
rect 22732 3844 22772 3884
rect 28396 4012 28436 4052
rect 36940 4012 36980 4052
rect 24076 3928 24116 3968
rect 29164 3928 29204 3968
rect 37804 3928 37844 3968
rect 47500 4180 47540 4220
rect 50860 4096 50900 4136
rect 52012 4096 52052 4136
rect 23116 3844 23156 3884
rect 28012 3844 28052 3884
rect 28300 3844 28340 3884
rect 31372 3844 31412 3884
rect 748 3760 788 3800
rect 3688 3760 3728 3800
rect 3770 3760 3810 3800
rect 3852 3760 3892 3800
rect 3934 3760 3974 3800
rect 4016 3760 4056 3800
rect 14284 3760 14324 3800
rect 18808 3760 18848 3800
rect 18890 3760 18930 3800
rect 18972 3760 19012 3800
rect 19054 3760 19094 3800
rect 19136 3760 19176 3800
rect 21964 3760 22004 3800
rect 22828 3760 22868 3800
rect 30988 3760 31028 3800
rect 33928 3760 33968 3800
rect 34010 3760 34050 3800
rect 34092 3760 34132 3800
rect 34174 3760 34214 3800
rect 34256 3760 34296 3800
rect 49048 3760 49088 3800
rect 49130 3760 49170 3800
rect 49212 3760 49252 3800
rect 49294 3760 49334 3800
rect 49376 3760 49416 3800
rect 13036 3676 13076 3716
rect 20140 3676 20180 3716
rect 23212 3676 23252 3716
rect 30220 3676 30260 3716
rect 4108 3592 4148 3632
rect 18316 3592 18356 3632
rect 18796 3592 18836 3632
rect 20620 3592 20660 3632
rect 20812 3592 20852 3632
rect 22924 3592 22964 3632
rect 23116 3592 23156 3632
rect 32428 3592 32468 3632
rect 10444 3508 10484 3548
rect 12940 3508 12980 3548
rect 16972 3508 17012 3548
rect 17260 3508 17300 3548
rect 22060 3508 22100 3548
rect 23212 3508 23252 3548
rect 268 3424 308 3464
rect 16780 3424 16820 3464
rect 18412 3424 18452 3464
rect 18700 3424 18740 3464
rect 19564 3424 19604 3464
rect 20524 3424 20564 3464
rect 21580 3424 21620 3464
rect 21772 3424 21812 3464
rect 25900 3424 25940 3464
rect 28972 3424 29012 3464
rect 30220 3424 30260 3464
rect 30604 3424 30644 3464
rect 30988 3424 31028 3464
rect 32428 3424 32468 3464
rect 32908 3424 32948 3464
rect 33772 3424 33812 3464
rect 35020 3424 35060 3464
rect 35212 3424 35252 3464
rect 10828 3340 10868 3380
rect 28012 3340 28052 3380
rect 31180 3340 31220 3380
rect 36940 3424 36980 3464
rect 37708 3424 37748 3464
rect 47212 3424 47252 3464
rect 44716 3340 44756 3380
rect 11212 3256 11252 3296
rect 32236 3256 32276 3296
rect 49420 3256 49460 3296
rect 50188 3256 50228 3296
rect 14668 3172 14708 3212
rect 15724 3172 15764 3212
rect 16780 3172 16820 3212
rect 17260 3172 17300 3212
rect 21484 3172 21524 3212
rect 22444 3172 22484 3212
rect 28684 3172 28724 3212
rect 30316 3172 30356 3212
rect 31660 3172 31700 3212
rect 32524 3172 32564 3212
rect 33004 3172 33044 3212
rect 33388 3172 33428 3212
rect 34348 3172 34388 3212
rect 35020 3172 35060 3212
rect 35692 3172 35732 3212
rect 36076 3172 36116 3212
rect 36460 3172 36500 3212
rect 37516 3172 37556 3212
rect 41740 3172 41771 3212
rect 41771 3172 41780 3212
rect 50860 3172 50900 3212
rect 51436 3172 51476 3212
rect 28012 3088 28052 3128
rect 4928 3004 4968 3044
rect 5010 3004 5050 3044
rect 5092 3004 5132 3044
rect 5174 3004 5214 3044
rect 5256 3004 5296 3044
rect 14572 3004 14612 3044
rect 19852 3004 19892 3044
rect 20048 3004 20088 3044
rect 20130 3004 20170 3044
rect 20212 3004 20252 3044
rect 20294 3004 20334 3044
rect 20376 3004 20416 3044
rect 22732 3004 22772 3044
rect 33100 3004 33140 3044
rect 35168 3004 35208 3044
rect 35250 3004 35290 3044
rect 35332 3004 35372 3044
rect 35414 3004 35454 3044
rect 35496 3004 35536 3044
rect 6988 2920 7028 2960
rect 21772 2920 21812 2960
rect 22444 2920 22484 2960
rect 24556 2920 24596 2960
rect 31660 2920 31700 2960
rect 49516 2920 49556 2960
rect 50288 3004 50328 3044
rect 50370 3004 50410 3044
rect 50452 3004 50492 3044
rect 50534 3004 50574 3044
rect 50616 3004 50656 3044
rect 14188 2836 14228 2876
rect 1420 2752 1460 2792
rect 15436 2752 15476 2792
rect 20620 2752 20660 2792
rect 23116 2836 23156 2876
rect 26860 2836 26900 2876
rect 37708 2836 37748 2876
rect 21388 2752 21428 2792
rect 26476 2752 26516 2792
rect 26668 2752 26708 2792
rect 30316 2752 30356 2792
rect 42412 2752 42452 2792
rect 44716 2752 44756 2792
rect 16204 2668 16244 2708
rect 19948 2668 19988 2708
rect 24460 2668 24500 2708
rect 28012 2668 28052 2708
rect 31468 2668 31508 2708
rect 39148 2668 39188 2708
rect 748 2584 788 2624
rect 15820 2584 15860 2624
rect 18220 2584 18260 2624
rect 19276 2584 19316 2624
rect 19468 2584 19508 2624
rect 21868 2584 21908 2624
rect 23020 2584 23060 2624
rect 23308 2584 23348 2624
rect 23692 2584 23732 2624
rect 24652 2584 24692 2624
rect 24940 2584 24980 2624
rect 25228 2584 25268 2624
rect 25900 2584 25940 2624
rect 27244 2584 27284 2624
rect 28780 2584 28820 2624
rect 29068 2584 29108 2624
rect 31660 2584 31700 2624
rect 34252 2584 34292 2624
rect 34540 2584 34580 2624
rect 36268 2584 36308 2624
rect 39724 2584 39764 2624
rect 49708 2584 49748 2624
rect 50188 2584 50228 2624
rect 52108 2584 52148 2624
rect 1420 2416 1460 2456
rect 4780 2416 4820 2456
rect 49420 2500 49460 2540
rect 22924 2416 22964 2456
rect 23116 2416 23156 2456
rect 24172 2416 24212 2456
rect 25036 2416 25076 2456
rect 25420 2416 25460 2456
rect 30316 2416 30356 2456
rect 3688 2248 3728 2288
rect 3770 2248 3810 2288
rect 3852 2248 3892 2288
rect 3934 2248 3974 2288
rect 4016 2248 4056 2288
rect 20428 2332 20468 2372
rect 21100 2332 21140 2372
rect 25708 2332 25748 2372
rect 27052 2332 27092 2372
rect 28396 2332 28436 2372
rect 28780 2332 28820 2372
rect 29836 2332 29876 2372
rect 18412 2248 18452 2288
rect 18808 2248 18848 2288
rect 18890 2248 18930 2288
rect 18972 2248 19012 2288
rect 19054 2248 19094 2288
rect 19136 2248 19176 2288
rect 23020 2248 23060 2288
rect 23212 2248 23252 2288
rect 2764 2164 2804 2204
rect 20908 2164 20948 2204
rect 19468 2080 19508 2120
rect 8908 1996 8948 2036
rect 20620 1996 20660 2036
rect 25228 2164 25268 2204
rect 21868 2080 21908 2120
rect 25036 2080 25076 2120
rect 21196 1996 21236 2036
rect 24844 1996 24884 2036
rect 29356 1996 29396 2036
rect 37612 2416 37652 2456
rect 39436 2416 39476 2456
rect 52588 2416 52628 2456
rect 33928 2248 33968 2288
rect 34010 2248 34050 2288
rect 34092 2248 34132 2288
rect 34174 2248 34214 2288
rect 34256 2248 34296 2288
rect 49048 2248 49088 2288
rect 49130 2248 49170 2288
rect 49212 2248 49252 2288
rect 49294 2248 49334 2288
rect 49376 2248 49416 2288
rect 34924 2080 34964 2120
rect 42412 2080 42452 2120
rect 37516 1996 37556 2036
rect 39436 1996 39476 2036
rect 40012 1996 40052 2036
rect 9292 1912 9332 1952
rect 21484 1912 21524 1952
rect 24556 1912 24596 1952
rect 25516 1912 25556 1952
rect 26092 1912 26132 1952
rect 26476 1912 26516 1952
rect 26860 1912 26900 1952
rect 28012 1912 28052 1952
rect 28396 1912 28436 1952
rect 28780 1912 28820 1952
rect 29164 1912 29204 1952
rect 29836 1912 29876 1952
rect 30316 1912 30356 1952
rect 31468 1912 31508 1952
rect 32236 1912 32276 1952
rect 32524 1912 32564 1952
rect 33004 1912 33044 1952
rect 33388 1912 33428 1952
rect 34348 1912 34388 1952
rect 35020 1912 35060 1952
rect 35692 1912 35732 1952
rect 36076 1912 36116 1952
rect 36460 1912 36500 1952
rect 37612 1912 37652 1952
rect 38380 1912 38420 1952
rect 39148 1912 39188 1952
rect 39532 1912 39572 1952
rect 40300 1912 40340 1952
rect 41068 1912 41108 1952
rect 41452 1912 41492 1952
rect 41836 1912 41876 1952
rect 42220 1912 42260 1952
rect 42604 1912 42644 1952
rect 49516 1912 49556 1952
rect 51436 1912 51476 1952
rect 3532 1828 3572 1868
rect 18220 1828 18260 1868
rect 18412 1828 18452 1868
rect 21772 1828 21812 1868
rect 22060 1828 22100 1868
rect 24076 1828 24116 1868
rect 25420 1828 25460 1868
rect 28684 1828 28724 1868
rect 37804 1828 37844 1868
rect 37996 1828 38036 1868
rect 50188 1828 50228 1868
rect 1420 1744 1460 1784
rect 4780 1744 4820 1784
rect 49708 1744 49748 1784
rect 52300 1744 52340 1784
rect 18412 1660 18452 1700
rect 22540 1660 22580 1700
rect 22732 1660 22772 1700
rect 23116 1660 23156 1700
rect 23500 1660 23540 1700
rect 23884 1660 23924 1700
rect 24268 1660 24308 1700
rect 24652 1660 24692 1700
rect 25036 1660 25076 1700
rect 25420 1660 25460 1700
rect 25804 1660 25844 1700
rect 26188 1660 26228 1700
rect 26572 1660 26612 1700
rect 26956 1660 26996 1700
rect 27340 1660 27380 1700
rect 27724 1660 27764 1700
rect 28108 1660 28148 1700
rect 28492 1660 28532 1700
rect 28876 1660 28916 1700
rect 29260 1660 29300 1700
rect 29644 1660 29684 1700
rect 30028 1660 30068 1700
rect 30412 1660 30452 1700
rect 30796 1660 30836 1700
rect 31180 1660 31220 1700
rect 31564 1660 31604 1700
rect 31948 1660 31988 1700
rect 32332 1660 32372 1700
rect 32716 1660 32756 1700
rect 33100 1660 33140 1700
rect 33484 1660 33524 1700
rect 33868 1660 33908 1700
rect 34252 1660 34292 1700
rect 34636 1660 34676 1700
rect 35020 1660 35060 1700
rect 35596 1660 35636 1700
rect 35788 1660 35828 1700
rect 36172 1660 36212 1700
rect 36556 1660 36596 1700
rect 36940 1660 36980 1700
rect 37324 1660 37364 1700
rect 37708 1660 37748 1700
rect 38092 1660 38132 1700
rect 38476 1660 38516 1700
rect 38860 1660 38900 1700
rect 39244 1660 39284 1700
rect 39628 1660 39668 1700
rect 40012 1660 40052 1700
rect 40396 1660 40436 1700
rect 40780 1660 40820 1700
rect 41164 1660 41204 1700
rect 41548 1660 41588 1700
rect 41932 1660 41972 1700
rect 42316 1660 42356 1700
rect 4300 1576 4340 1616
rect 4928 1492 4968 1532
rect 5010 1492 5050 1532
rect 5092 1492 5132 1532
rect 5174 1492 5214 1532
rect 5256 1492 5296 1532
rect 23692 1576 23732 1616
rect 24172 1576 24212 1616
rect 29548 1576 29588 1616
rect 35980 1576 36020 1616
rect 39532 1576 39572 1616
rect 51916 1576 51956 1616
rect 20048 1492 20088 1532
rect 20130 1492 20170 1532
rect 20212 1492 20252 1532
rect 20294 1492 20334 1532
rect 20376 1492 20416 1532
rect 20620 1492 20660 1532
rect 24460 1492 24500 1532
rect 29356 1492 29396 1532
rect 34924 1492 34964 1532
rect 35168 1492 35208 1532
rect 35250 1492 35290 1532
rect 35332 1492 35372 1532
rect 35414 1492 35454 1532
rect 35496 1492 35536 1532
rect 37900 1492 37940 1532
rect 50288 1492 50328 1532
rect 50370 1492 50410 1532
rect 50452 1492 50492 1532
rect 50534 1492 50574 1532
rect 50616 1492 50656 1532
rect 1420 1408 1460 1448
rect 22924 1408 22964 1448
rect 25900 1408 25940 1448
rect 52588 1408 52628 1448
rect 29068 1240 29108 1280
rect 1420 1072 1460 1112
rect 51916 1072 51956 1112
rect 748 736 788 776
rect 52300 736 52340 776
rect 21580 316 21620 356
rect 36268 316 36308 356
rect 9676 232 9716 272
rect 24748 232 24788 272
rect 25612 232 25652 272
rect 46156 232 46196 272
rect 21292 148 21332 188
rect 23788 148 23828 188
rect 45772 148 45812 188
rect 45388 64 45428 104
<< metal3 >>
rect 1592 12100 1672 12180
rect 4088 12100 4168 12180
rect 6584 12100 6664 12180
rect 9080 12100 9160 12180
rect 11576 12100 11656 12180
rect 14072 12100 14152 12180
rect 16568 12100 16648 12180
rect 19064 12100 19144 12180
rect 21560 12100 21640 12180
rect 24056 12100 24136 12180
rect 26552 12100 26632 12180
rect 29048 12100 29128 12180
rect 31544 12100 31624 12180
rect 34040 12100 34120 12180
rect 36536 12100 36616 12180
rect 39032 12100 39112 12180
rect 41528 12100 41608 12180
rect 44024 12100 44104 12180
rect 46520 12100 46600 12180
rect 49016 12100 49096 12180
rect 51512 12100 51592 12180
rect 844 11192 884 11201
rect 844 9764 884 11152
rect 1612 10436 1652 12100
rect 1612 10387 1652 10396
rect 4108 10436 4148 12100
rect 4928 10604 5296 10613
rect 4968 10564 5010 10604
rect 5050 10564 5092 10604
rect 5132 10564 5174 10604
rect 5214 10564 5256 10604
rect 4928 10555 5296 10564
rect 4108 10387 4148 10396
rect 6604 10436 6644 12100
rect 6604 10387 6644 10396
rect 9100 10436 9140 12100
rect 9100 10387 9140 10396
rect 11596 10436 11636 12100
rect 11596 10387 11636 10396
rect 14092 10436 14132 12100
rect 14092 10387 14132 10396
rect 14284 10520 14324 10529
rect 844 9715 884 9724
rect 1900 10184 1940 10193
rect 1900 9260 1940 10144
rect 4396 10184 4436 10193
rect 3688 9848 4056 9857
rect 3728 9808 3770 9848
rect 3810 9808 3852 9848
rect 3892 9808 3934 9848
rect 3974 9808 4016 9848
rect 3688 9799 4056 9808
rect 4396 9344 4436 10144
rect 6892 10184 6932 10193
rect 6892 9596 6932 10144
rect 9388 10184 9428 10193
rect 9388 9764 9428 10144
rect 9388 9715 9428 9724
rect 13612 10184 13652 10193
rect 13612 9680 13652 10144
rect 13612 9631 13652 9640
rect 6892 9547 6932 9556
rect 4396 9295 4436 9304
rect 14092 9512 14132 9521
rect 1900 9211 1940 9220
rect 4928 9092 5296 9101
rect 4968 9052 5010 9092
rect 5050 9052 5092 9092
rect 5132 9052 5174 9092
rect 5214 9052 5256 9092
rect 4928 9043 5296 9052
rect 748 8924 788 8933
rect 364 8000 404 8009
rect 268 6404 308 6413
rect 268 3464 308 6364
rect 364 4472 404 7960
rect 364 4423 404 4432
rect 460 7244 500 7253
rect 460 4136 500 7204
rect 460 4087 500 4096
rect 748 3800 788 8884
rect 1228 8840 1268 8849
rect 1132 8672 1172 8681
rect 1036 7076 1076 7085
rect 1036 4808 1076 7036
rect 1132 5144 1172 8632
rect 1228 8084 1268 8800
rect 3688 8336 4056 8345
rect 3728 8296 3770 8336
rect 3810 8296 3852 8336
rect 3892 8296 3934 8336
rect 3974 8296 4016 8336
rect 3688 8287 4056 8296
rect 1228 8035 1268 8044
rect 1324 8168 1364 8177
rect 1228 7160 1268 7169
rect 1228 5228 1268 7120
rect 1324 6656 1364 8128
rect 4928 7580 5296 7589
rect 4968 7540 5010 7580
rect 5050 7540 5092 7580
rect 5132 7540 5174 7580
rect 5214 7540 5256 7580
rect 4928 7531 5296 7540
rect 10732 7160 10772 7169
rect 3688 6824 4056 6833
rect 3728 6784 3770 6824
rect 3810 6784 3852 6824
rect 3892 6784 3934 6824
rect 3974 6784 4016 6824
rect 3688 6775 4056 6784
rect 1324 6607 1364 6616
rect 1228 5179 1268 5188
rect 1420 6488 1460 6497
rect 1132 5095 1172 5104
rect 1420 5060 1460 6448
rect 4928 6068 5296 6077
rect 4968 6028 5010 6068
rect 5050 6028 5092 6068
rect 5132 6028 5174 6068
rect 5214 6028 5256 6068
rect 4928 6019 5296 6028
rect 10732 5480 10772 7120
rect 10732 5431 10772 5440
rect 3688 5312 4056 5321
rect 3728 5272 3770 5312
rect 3810 5272 3852 5312
rect 3892 5272 3934 5312
rect 3974 5272 4016 5312
rect 3688 5263 4056 5272
rect 1420 5011 1460 5020
rect 1036 4759 1076 4768
rect 5452 4892 5492 4901
rect 4928 4556 5296 4565
rect 4968 4516 5010 4556
rect 5050 4516 5092 4556
rect 5132 4516 5174 4556
rect 5214 4516 5256 4556
rect 4928 4507 5296 4516
rect 748 3751 788 3760
rect 3688 3800 4056 3809
rect 3728 3760 3770 3800
rect 3810 3760 3852 3800
rect 3892 3760 3934 3800
rect 3974 3760 4016 3800
rect 3688 3751 4056 3760
rect 268 3415 308 3424
rect 4108 3632 4148 3641
rect 1420 2792 1460 2801
rect 1420 2657 1460 2752
rect 748 2624 788 2633
rect 748 776 788 2584
rect 1420 2456 1460 2465
rect 1420 2321 1460 2416
rect 3688 2288 4056 2297
rect 3728 2248 3770 2288
rect 3810 2248 3852 2288
rect 3892 2248 3934 2288
rect 3974 2248 4016 2288
rect 3688 2239 4056 2248
rect 2764 2204 2804 2213
rect 1420 1784 1460 1793
rect 1420 1649 1460 1744
rect 1420 1448 1460 1457
rect 1420 1313 1460 1408
rect 1420 1112 1460 1121
rect 1420 977 1460 1072
rect 748 727 788 736
rect 2764 80 2804 2164
rect 3148 1868 3188 1877
rect 3148 80 3188 1828
rect 3532 1868 3572 1877
rect 3532 80 3572 1828
rect 4108 188 4148 3592
rect 4928 3044 5296 3053
rect 4968 3004 5010 3044
rect 5050 3004 5092 3044
rect 5132 3004 5174 3044
rect 5214 3004 5256 3044
rect 4928 2995 5296 3004
rect 4780 2456 4820 2465
rect 4780 1784 4820 2416
rect 4780 1735 4820 1744
rect 3916 148 4148 188
rect 4300 1616 4340 1625
rect 3916 80 3956 148
rect 4300 80 4340 1576
rect 4928 1532 5296 1541
rect 4968 1492 5010 1532
rect 5050 1492 5092 1532
rect 5132 1492 5174 1532
rect 5214 1492 5256 1532
rect 4928 1483 5296 1492
rect 4684 524 4724 533
rect 4684 80 4724 484
rect 5068 440 5108 449
rect 5068 80 5108 400
rect 5452 80 5492 4852
rect 5836 4808 5876 4817
rect 5836 80 5876 4768
rect 6220 4472 6260 4481
rect 6220 80 6260 4432
rect 6604 4304 6644 4313
rect 6604 80 6644 4264
rect 11596 4220 11636 4229
rect 8524 4136 8564 4145
rect 6988 2960 7028 2969
rect 6988 80 7028 2920
rect 8140 2960 8180 2969
rect 7372 2624 7412 2633
rect 7372 80 7412 2584
rect 7756 1616 7796 1625
rect 7756 80 7796 1576
rect 8140 80 8180 2920
rect 8524 80 8564 4096
rect 10444 3548 10484 3557
rect 8908 2036 8948 2045
rect 8908 80 8948 1996
rect 9292 1952 9332 1961
rect 9292 80 9332 1912
rect 10060 356 10100 365
rect 9676 272 9716 281
rect 9676 80 9716 232
rect 10060 80 10100 316
rect 10444 80 10484 3508
rect 10828 3380 10868 3389
rect 10828 80 10868 3340
rect 11212 3296 11252 3305
rect 11212 80 11252 3256
rect 11596 80 11636 4180
rect 13708 4220 13748 4229
rect 12748 3884 12788 3893
rect 12364 2540 12404 2549
rect 11980 272 12020 281
rect 11980 80 12020 232
rect 12364 80 12404 2500
rect 12748 80 12788 3844
rect 13036 3716 13076 3725
rect 12940 3548 12980 3557
rect 13036 3548 13076 3676
rect 12980 3508 13076 3548
rect 12940 3499 12980 3508
rect 13132 1700 13172 1709
rect 13132 80 13172 1660
rect 13708 188 13748 4180
rect 13516 148 13748 188
rect 13900 3548 13940 3557
rect 13516 80 13556 148
rect 13900 80 13940 3508
rect 14092 104 14132 9472
rect 14284 9512 14324 10480
rect 16588 10436 16628 12100
rect 16588 10387 16628 10396
rect 19084 10436 19124 12100
rect 20048 10604 20416 10613
rect 20088 10564 20130 10604
rect 20170 10564 20212 10604
rect 20252 10564 20294 10604
rect 20334 10564 20376 10604
rect 20048 10555 20416 10564
rect 19084 10387 19124 10396
rect 21580 10436 21620 12100
rect 21580 10387 21620 10396
rect 23596 10856 23636 10865
rect 14380 10184 14420 10193
rect 14380 9680 14420 10144
rect 18412 10184 18452 10193
rect 14380 9631 14420 9640
rect 15436 10100 15476 10109
rect 14284 9463 14324 9472
rect 15436 9428 15476 10060
rect 18412 9680 18452 10144
rect 20812 10184 20852 10193
rect 18808 9848 19176 9857
rect 18848 9808 18890 9848
rect 18930 9808 18972 9848
rect 19012 9808 19054 9848
rect 19094 9808 19136 9848
rect 18808 9799 19176 9808
rect 19372 9848 19412 9857
rect 18412 9631 18452 9640
rect 15436 9379 15476 9388
rect 18700 9512 18740 9521
rect 18700 9377 18740 9472
rect 19372 9428 19412 9808
rect 20812 9680 20852 10144
rect 20812 9631 20852 9640
rect 23116 10184 23156 10193
rect 23116 9680 23156 10144
rect 23116 9631 23156 9640
rect 19372 9379 19412 9388
rect 21292 9512 21332 9521
rect 20140 9260 20180 9355
rect 20140 9211 20180 9220
rect 20524 9176 20564 9185
rect 20812 9176 20852 9185
rect 20564 9136 20812 9176
rect 20524 9127 20564 9136
rect 20812 9127 20852 9136
rect 20048 9092 20416 9101
rect 20088 9052 20130 9092
rect 20170 9052 20212 9092
rect 20252 9052 20294 9092
rect 20334 9052 20376 9092
rect 20048 9043 20416 9052
rect 18808 8336 19176 8345
rect 18848 8296 18890 8336
rect 18930 8296 18972 8336
rect 19012 8296 19054 8336
rect 19094 8296 19136 8336
rect 18808 8287 19176 8296
rect 20048 7580 20416 7589
rect 20088 7540 20130 7580
rect 20170 7540 20212 7580
rect 20252 7540 20294 7580
rect 20334 7540 20376 7580
rect 20048 7531 20416 7540
rect 19948 6992 19988 7001
rect 18808 6824 19176 6833
rect 18848 6784 18890 6824
rect 18930 6784 18972 6824
rect 19012 6784 19054 6824
rect 19094 6784 19136 6824
rect 18808 6775 19176 6784
rect 19948 5564 19988 6952
rect 20048 6068 20416 6077
rect 20088 6028 20130 6068
rect 20170 6028 20212 6068
rect 20252 6028 20294 6068
rect 20334 6028 20376 6068
rect 20048 6019 20416 6028
rect 19948 5515 19988 5524
rect 18808 5312 19176 5321
rect 18848 5272 18890 5312
rect 18930 5272 18972 5312
rect 19012 5272 19054 5312
rect 19094 5272 19136 5312
rect 18808 5263 19176 5272
rect 14668 4976 14708 4985
rect 14668 4640 14708 4936
rect 18124 4976 18164 4985
rect 14668 4591 14708 4600
rect 15340 4724 15380 4733
rect 14380 3968 14420 3977
rect 14284 3800 14324 3809
rect 14188 2876 14228 2885
rect 14188 2741 14228 2836
rect 2744 0 2824 80
rect 3128 0 3208 80
rect 3512 0 3592 80
rect 3896 0 3976 80
rect 4280 0 4360 80
rect 4664 0 4744 80
rect 5048 0 5128 80
rect 5432 0 5512 80
rect 5816 0 5896 80
rect 6200 0 6280 80
rect 6584 0 6664 80
rect 6968 0 7048 80
rect 7352 0 7432 80
rect 7736 0 7816 80
rect 8120 0 8200 80
rect 8504 0 8584 80
rect 8888 0 8968 80
rect 9272 0 9352 80
rect 9656 0 9736 80
rect 10040 0 10120 80
rect 10424 0 10504 80
rect 10808 0 10888 80
rect 11192 0 11272 80
rect 11576 0 11656 80
rect 11960 0 12040 80
rect 12344 0 12424 80
rect 12728 0 12808 80
rect 13112 0 13192 80
rect 13496 0 13576 80
rect 13880 0 13960 80
rect 14284 80 14324 3760
rect 14380 1532 14420 3928
rect 14668 3212 14708 3221
rect 14380 1483 14420 1492
rect 14572 3044 14612 3053
rect 14572 608 14612 3004
rect 14668 2036 14708 3172
rect 14668 1987 14708 1996
rect 15052 2876 15092 2885
rect 14572 568 14708 608
rect 14668 80 14708 568
rect 15052 80 15092 2836
rect 15340 2204 15380 4684
rect 15628 4724 15668 4733
rect 15340 2155 15380 2164
rect 15436 2792 15476 2801
rect 15436 80 15476 2752
rect 15628 2372 15668 4684
rect 17740 4640 17780 4649
rect 16300 4220 16340 4229
rect 16204 4136 16244 4145
rect 15628 2323 15668 2332
rect 15724 3212 15764 3221
rect 15724 2120 15764 3172
rect 16204 2900 16244 4096
rect 16300 3884 16340 4180
rect 16300 3835 16340 3844
rect 16876 3968 16916 3977
rect 16780 3464 16820 3473
rect 16780 3212 16820 3424
rect 16780 3163 16820 3172
rect 16204 2860 16628 2900
rect 16204 2708 16244 2717
rect 15724 2071 15764 2080
rect 15820 2624 15860 2633
rect 15820 80 15860 2584
rect 16204 80 16244 2668
rect 16588 80 16628 2860
rect 16876 2876 16916 3928
rect 16876 2827 16916 2836
rect 16972 3548 17012 3557
rect 16972 80 17012 3508
rect 17260 3548 17300 3557
rect 17260 3413 17300 3508
rect 17260 3212 17300 3221
rect 17260 2900 17300 3172
rect 17260 2860 17396 2900
rect 17356 80 17396 2860
rect 17740 80 17780 4600
rect 18124 80 18164 4936
rect 20048 4556 20416 4565
rect 20088 4516 20130 4556
rect 20170 4516 20212 4556
rect 20252 4516 20294 4556
rect 20334 4516 20376 4556
rect 20048 4507 20416 4516
rect 18508 4220 18548 4229
rect 18316 4136 18356 4145
rect 18316 3632 18356 4096
rect 18316 3583 18356 3592
rect 18412 3968 18452 3977
rect 18412 3464 18452 3928
rect 18412 3415 18452 3424
rect 18220 2624 18260 2633
rect 18220 1868 18260 2584
rect 18220 1819 18260 1828
rect 18412 2288 18452 2297
rect 18412 1868 18452 2248
rect 18412 1819 18452 1828
rect 18412 1700 18452 1709
rect 18412 356 18452 1660
rect 18412 307 18452 316
rect 18508 80 18548 4180
rect 18700 4220 18740 4229
rect 18604 3884 18644 3893
rect 18700 3884 18740 4180
rect 18644 3844 18740 3884
rect 19660 4136 19700 4145
rect 18604 3835 18644 3844
rect 18808 3800 19176 3809
rect 18848 3760 18890 3800
rect 18930 3760 18972 3800
rect 19012 3760 19054 3800
rect 19094 3760 19136 3800
rect 18808 3751 19176 3760
rect 18796 3632 18836 3641
rect 18700 3464 18740 3473
rect 18700 2708 18740 3424
rect 18700 2659 18740 2668
rect 18796 2456 18836 3592
rect 19564 3464 19604 3473
rect 19372 2708 19412 2717
rect 18700 2416 18836 2456
rect 19276 2624 19316 2633
rect 18700 188 18740 2416
rect 18808 2288 19176 2297
rect 18848 2248 18890 2288
rect 18930 2248 18972 2288
rect 19012 2248 19054 2288
rect 19094 2248 19136 2288
rect 18808 2239 19176 2248
rect 18700 148 18932 188
rect 18892 80 18932 148
rect 19276 80 19316 2584
rect 19372 1868 19412 2668
rect 19468 2624 19508 2633
rect 19468 2120 19508 2584
rect 19468 2071 19508 2080
rect 19564 1952 19604 3424
rect 19660 2876 19700 4096
rect 19852 4136 19892 4145
rect 19852 3044 19892 4096
rect 20716 3968 20756 3977
rect 20140 3716 20180 3725
rect 20140 3581 20180 3676
rect 20620 3632 20660 3641
rect 20620 3497 20660 3592
rect 20524 3464 20564 3473
rect 19852 2995 19892 3004
rect 20048 3044 20416 3053
rect 20088 3004 20130 3044
rect 20170 3004 20212 3044
rect 20252 3004 20294 3044
rect 20334 3004 20376 3044
rect 20048 2995 20416 3004
rect 19660 2836 19892 2876
rect 19852 2120 19892 2836
rect 19564 1903 19604 1912
rect 19660 2080 19892 2120
rect 19948 2708 19988 2717
rect 19372 1819 19412 1828
rect 19660 80 19700 2080
rect 19852 1952 19892 1961
rect 19852 1532 19892 1912
rect 19852 1483 19892 1492
rect 19948 1364 19988 2668
rect 20428 2372 20468 2381
rect 20428 2237 20468 2332
rect 20048 1532 20416 1541
rect 20088 1492 20130 1532
rect 20170 1492 20212 1532
rect 20252 1492 20294 1532
rect 20334 1492 20376 1532
rect 20048 1483 20416 1492
rect 19948 1324 20084 1364
rect 20044 80 20084 1324
rect 20524 1112 20564 3424
rect 20620 2792 20660 2801
rect 20620 2708 20660 2752
rect 20620 2657 20660 2668
rect 20620 2036 20660 2045
rect 20620 1532 20660 1996
rect 20716 1616 20756 3928
rect 20716 1567 20756 1576
rect 20812 3632 20852 3641
rect 20620 1483 20660 1492
rect 20428 1072 20564 1112
rect 20428 80 20468 1072
rect 20812 80 20852 3592
rect 21196 2708 21236 2717
rect 21100 2372 21140 2381
rect 20908 2332 21100 2372
rect 20908 2204 20948 2332
rect 21100 2323 21140 2332
rect 20908 2155 20948 2164
rect 21196 2036 21236 2668
rect 21196 1987 21236 1996
rect 21196 356 21236 365
rect 21196 80 21236 316
rect 21292 188 21332 9472
rect 23596 9512 23636 10816
rect 24076 10436 24116 12100
rect 24076 10387 24116 10396
rect 26572 10436 26612 12100
rect 26572 10387 26612 10396
rect 29068 10436 29108 12100
rect 29068 10387 29108 10396
rect 31564 10436 31604 12100
rect 31564 10387 31604 10396
rect 34060 10436 34100 12100
rect 35168 10604 35536 10613
rect 35208 10564 35250 10604
rect 35290 10564 35332 10604
rect 35372 10564 35414 10604
rect 35454 10564 35496 10604
rect 35168 10555 35536 10564
rect 34060 10387 34100 10396
rect 24172 10352 24212 10361
rect 24172 9680 24212 10312
rect 26668 10268 26708 10277
rect 25228 10184 25268 10193
rect 24172 9631 24212 9640
rect 24268 10016 24308 10025
rect 23596 9463 23636 9472
rect 23788 9428 23828 9437
rect 21580 7832 21620 7841
rect 21580 7160 21620 7792
rect 21580 7111 21620 7120
rect 22924 7496 22964 7505
rect 21580 6740 21620 6749
rect 21580 5648 21620 6700
rect 22732 6488 22772 6497
rect 22732 5816 22772 6448
rect 22924 6488 22964 7456
rect 22924 6439 22964 6448
rect 22732 5767 22772 5776
rect 22924 6236 22964 6245
rect 22924 5732 22964 6196
rect 22924 5683 22964 5692
rect 21580 5599 21620 5608
rect 22828 4388 22868 4397
rect 22636 4052 22676 4147
rect 22636 4003 22676 4012
rect 22732 3884 22772 3893
rect 21964 3800 22004 3809
rect 21580 3464 21620 3473
rect 21580 3329 21620 3424
rect 21772 3464 21812 3473
rect 21484 3212 21524 3221
rect 21388 2792 21428 2801
rect 21388 2372 21428 2752
rect 21388 2323 21428 2332
rect 21484 1952 21524 3172
rect 21772 2960 21812 3424
rect 21772 2911 21812 2920
rect 21484 1903 21524 1912
rect 21772 2708 21812 2717
rect 21772 1868 21812 2668
rect 21868 2624 21908 2633
rect 21868 2120 21908 2584
rect 21868 2071 21908 2080
rect 21772 1819 21812 1828
rect 21292 139 21332 148
rect 21580 356 21620 365
rect 21580 80 21620 316
rect 21964 80 22004 3760
rect 22060 3548 22100 3557
rect 22060 1868 22100 3508
rect 22732 3548 22772 3844
rect 22828 3800 22868 4348
rect 23308 4304 23348 4313
rect 22924 4220 22964 4229
rect 22924 4085 22964 4180
rect 23212 4220 23252 4229
rect 23116 4052 23156 4061
rect 23116 3884 23156 4012
rect 23116 3835 23156 3844
rect 22828 3751 22868 3760
rect 22924 3800 22964 3809
rect 22924 3632 22964 3760
rect 23212 3716 23252 4180
rect 23308 3884 23348 4264
rect 23308 3835 23348 3844
rect 23212 3667 23252 3676
rect 22924 3583 22964 3592
rect 23116 3632 23156 3641
rect 22732 3499 22772 3508
rect 23116 3497 23156 3592
rect 23212 3548 23252 3557
rect 23212 3413 23252 3508
rect 22444 3212 22484 3221
rect 22444 2960 22484 3172
rect 22444 2911 22484 2920
rect 22732 3044 22772 3053
rect 22732 2456 22772 3004
rect 23116 2876 23156 2885
rect 23156 2836 23252 2876
rect 23116 2827 23156 2836
rect 23020 2624 23060 2633
rect 22060 1819 22100 1828
rect 22348 2416 22772 2456
rect 22828 2584 23020 2624
rect 22348 80 22388 2416
rect 22540 2288 22580 2297
rect 22540 1700 22580 2248
rect 22540 1651 22580 1660
rect 22732 1700 22772 1709
rect 22732 80 22772 1660
rect 22828 524 22868 2584
rect 23020 2575 23060 2584
rect 22924 2456 22964 2465
rect 22924 1448 22964 2416
rect 23116 2456 23156 2465
rect 23020 2288 23060 2297
rect 23116 2288 23156 2416
rect 23060 2248 23156 2288
rect 23212 2288 23252 2836
rect 23020 2239 23060 2248
rect 23212 2239 23252 2248
rect 23308 2624 23348 2633
rect 22924 1399 22964 1408
rect 23116 1700 23156 1709
rect 22828 475 22868 484
rect 23116 80 23156 1660
rect 23308 440 23348 2584
rect 23692 2624 23732 2633
rect 23308 391 23348 400
rect 23500 1700 23540 1709
rect 23500 80 23540 1660
rect 23692 1616 23732 2584
rect 23692 1567 23732 1576
rect 23788 188 23828 9388
rect 23980 9428 24020 9437
rect 23980 8168 24020 9388
rect 24268 8672 24308 9976
rect 25228 9680 25268 10144
rect 25228 9631 25268 9640
rect 26572 10100 26612 10109
rect 24268 8623 24308 8632
rect 25612 9512 25652 9521
rect 23980 8119 24020 8128
rect 23884 8084 23924 8093
rect 23884 7160 23924 8044
rect 23884 7111 23924 7120
rect 24172 7160 24212 7169
rect 24172 5648 24212 7120
rect 24172 5599 24212 5608
rect 24172 4976 24212 4985
rect 24172 4472 24212 4936
rect 24172 4423 24212 4432
rect 24844 4724 24884 4733
rect 24076 3968 24116 3977
rect 24076 1868 24116 3928
rect 24556 2960 24596 2969
rect 24460 2708 24500 2717
rect 24076 1819 24116 1828
rect 24172 2456 24212 2465
rect 23788 139 23828 148
rect 23884 1700 23924 1709
rect 23884 80 23924 1660
rect 24172 1616 24212 2416
rect 24172 1567 24212 1576
rect 24268 1700 24308 1709
rect 24268 80 24308 1660
rect 24460 1532 24500 2668
rect 24556 1952 24596 2920
rect 24652 2624 24692 2633
rect 24692 2584 24788 2624
rect 24652 2575 24692 2584
rect 24556 1903 24596 1912
rect 24460 1483 24500 1492
rect 24652 1700 24692 1709
rect 24652 80 24692 1660
rect 24748 272 24788 2584
rect 24844 2036 24884 4684
rect 25516 4724 25556 4733
rect 24940 2624 24980 2633
rect 24940 2288 24980 2584
rect 25228 2624 25268 2633
rect 24940 2239 24980 2248
rect 25036 2456 25076 2465
rect 25036 2120 25076 2416
rect 25228 2204 25268 2584
rect 25228 2155 25268 2164
rect 25420 2456 25460 2465
rect 25036 2071 25076 2080
rect 24844 1987 24884 1996
rect 25420 1868 25460 2416
rect 25516 1952 25556 4684
rect 25516 1903 25556 1912
rect 25420 1819 25460 1828
rect 24748 223 24788 232
rect 25036 1700 25076 1709
rect 25036 80 25076 1660
rect 25420 1700 25460 1709
rect 25420 80 25460 1660
rect 25612 272 25652 9472
rect 26188 9512 26228 9521
rect 26188 8924 26228 9472
rect 26188 8875 26228 8884
rect 26380 9260 26420 9269
rect 26380 8672 26420 9220
rect 26572 8924 26612 10060
rect 26668 9512 26708 10228
rect 27820 10184 27860 10193
rect 27724 10100 27764 10109
rect 26956 10016 26996 10025
rect 26956 9680 26996 9976
rect 27724 9848 27764 10060
rect 27724 9799 27764 9808
rect 26956 9631 26996 9640
rect 27820 9680 27860 10144
rect 29356 10184 29396 10193
rect 29164 10016 29204 10025
rect 28876 9932 28916 9941
rect 27820 9631 27860 9640
rect 27916 9848 27956 9857
rect 26668 9463 26708 9472
rect 27916 9344 27956 9808
rect 28588 9512 28628 9521
rect 27916 9295 27956 9304
rect 28396 9428 28436 9437
rect 28300 9260 28340 9271
rect 28300 9176 28340 9220
rect 28300 9127 28340 9136
rect 28396 9092 28436 9388
rect 28588 9260 28628 9472
rect 28876 9512 28916 9892
rect 29164 9680 29204 9976
rect 29164 9631 29204 9640
rect 29356 9680 29396 10144
rect 36556 10184 36596 12100
rect 36940 10520 36980 10529
rect 36748 10480 36940 10520
rect 36748 10268 36788 10480
rect 36940 10471 36980 10480
rect 39052 10436 39092 12100
rect 39052 10387 39092 10396
rect 39148 10604 39188 10613
rect 36748 10219 36788 10228
rect 36556 10135 36596 10144
rect 39148 10184 39188 10564
rect 41548 10436 41588 12100
rect 41548 10387 41588 10396
rect 44044 10436 44084 12100
rect 46156 10604 46196 10613
rect 44044 10387 44084 10396
rect 44908 10520 44948 10529
rect 44620 10268 44660 10277
rect 39148 10135 39188 10144
rect 43372 10184 43412 10193
rect 30700 10100 30740 10109
rect 29356 9631 29396 9640
rect 30028 9848 30068 9857
rect 30028 9596 30068 9808
rect 30028 9547 30068 9556
rect 28876 9463 28916 9472
rect 29932 9512 29972 9521
rect 28588 9211 28628 9220
rect 28396 9043 28436 9052
rect 26572 8875 26612 8884
rect 28108 9008 28148 9017
rect 26380 8623 26420 8632
rect 27340 8672 27380 8681
rect 25708 7748 25748 7757
rect 25708 6572 25748 7708
rect 25708 6523 25748 6532
rect 25804 6488 25844 6497
rect 25804 6152 25844 6448
rect 25804 6103 25844 6112
rect 26092 4640 26132 4649
rect 25900 3464 25940 3473
rect 25900 2960 25940 3424
rect 25900 2911 25940 2920
rect 25900 2624 25940 2633
rect 25708 2372 25748 2381
rect 25708 1532 25748 2332
rect 25708 1483 25748 1492
rect 25804 1700 25844 1709
rect 25612 223 25652 232
rect 25804 80 25844 1660
rect 25900 1448 25940 2584
rect 26092 1952 26132 4600
rect 27340 4388 27380 8632
rect 27916 8672 27956 8681
rect 27820 5648 27860 5657
rect 27820 5228 27860 5608
rect 27820 5179 27860 5188
rect 27916 5144 27956 8632
rect 28108 8672 28148 8968
rect 29932 9008 29972 9472
rect 29932 8959 29972 8968
rect 30220 9512 30260 9521
rect 30220 8924 30260 9472
rect 30700 9428 30740 10060
rect 37996 10016 38036 10025
rect 38036 9976 38132 10016
rect 37996 9967 38036 9976
rect 33928 9848 34296 9857
rect 33968 9808 34010 9848
rect 34050 9808 34092 9848
rect 34132 9808 34174 9848
rect 34214 9808 34256 9848
rect 33928 9799 34296 9808
rect 35020 9848 35060 9857
rect 30700 9379 30740 9388
rect 35020 9092 35060 9808
rect 37900 9764 37940 9773
rect 38092 9764 38132 9976
rect 43276 9932 43316 9941
rect 37940 9724 38036 9764
rect 37900 9715 37940 9724
rect 37996 9344 38036 9724
rect 38092 9715 38132 9724
rect 38284 9848 38324 9857
rect 38284 9512 38324 9808
rect 38284 9463 38324 9472
rect 43084 9680 43124 9689
rect 42700 9428 42740 9437
rect 37996 9304 38324 9344
rect 38284 9260 38324 9304
rect 38284 9211 38324 9220
rect 35020 9043 35060 9052
rect 35168 9092 35536 9101
rect 35208 9052 35250 9092
rect 35290 9052 35332 9092
rect 35372 9052 35414 9092
rect 35454 9052 35496 9092
rect 35168 9043 35536 9052
rect 30220 8875 30260 8884
rect 37996 9008 38036 9017
rect 28108 8623 28148 8632
rect 33196 8672 33236 8681
rect 27916 5095 27956 5104
rect 33196 7748 33236 8632
rect 37996 8672 38036 8968
rect 37996 8623 38036 8632
rect 33928 8336 34296 8345
rect 33968 8296 34010 8336
rect 34050 8296 34092 8336
rect 34132 8296 34174 8336
rect 34214 8296 34256 8336
rect 33928 8287 34296 8296
rect 38092 8084 38132 8093
rect 27340 4339 27380 4348
rect 32908 4304 32948 4313
rect 28012 4136 28052 4145
rect 28012 4001 28052 4096
rect 28204 4136 28244 4145
rect 28012 3884 28052 3893
rect 28204 3884 28244 4096
rect 28396 4052 28436 4061
rect 28052 3844 28244 3884
rect 28300 3884 28340 3893
rect 28012 3835 28052 3844
rect 28300 3800 28340 3844
rect 28300 3749 28340 3760
rect 28396 3716 28436 4012
rect 28396 3667 28436 3676
rect 29164 3968 29204 3977
rect 28972 3464 29012 3473
rect 28012 3380 28052 3389
rect 28012 3128 28052 3340
rect 28012 3079 28052 3088
rect 28684 3212 28724 3221
rect 26860 2876 26900 2885
rect 26092 1903 26132 1912
rect 26476 2792 26516 2801
rect 26476 1952 26516 2752
rect 26668 2792 26708 2801
rect 26668 2708 26708 2752
rect 26668 2657 26708 2668
rect 26476 1903 26516 1912
rect 26860 1952 26900 2836
rect 28012 2708 28052 2717
rect 27244 2624 27284 2633
rect 27052 2584 27244 2624
rect 27052 2372 27092 2584
rect 27244 2575 27284 2584
rect 27052 2323 27092 2332
rect 26860 1903 26900 1912
rect 28012 1952 28052 2668
rect 28012 1903 28052 1912
rect 28108 2708 28148 2717
rect 28108 1868 28148 2668
rect 28396 2372 28436 2381
rect 28396 1952 28436 2332
rect 28396 1903 28436 1912
rect 28108 1819 28148 1828
rect 28684 1868 28724 3172
rect 28780 2624 28820 2633
rect 28780 2489 28820 2584
rect 28780 2372 28820 2381
rect 28780 1952 28820 2332
rect 28780 1903 28820 1912
rect 28684 1819 28724 1828
rect 25900 1399 25940 1408
rect 26188 1700 26228 1709
rect 26188 80 26228 1660
rect 26572 1700 26612 1709
rect 26572 80 26612 1660
rect 26956 1700 26996 1709
rect 26956 80 26996 1660
rect 27340 1700 27380 1709
rect 27340 80 27380 1660
rect 27724 1700 27764 1709
rect 27724 80 27764 1660
rect 28108 1700 28148 1709
rect 28108 80 28148 1660
rect 28492 1700 28532 1709
rect 28492 80 28532 1660
rect 28876 1700 28916 1709
rect 28876 80 28916 1660
rect 28972 1112 29012 3424
rect 29068 2624 29108 2633
rect 29068 1280 29108 2584
rect 29164 1952 29204 3928
rect 31372 3884 31412 3893
rect 30220 3716 30260 3811
rect 30220 3667 30260 3676
rect 30988 3800 31028 3809
rect 29548 3464 29588 3473
rect 29164 1903 29204 1912
rect 29356 2036 29396 2045
rect 29068 1231 29108 1240
rect 29260 1700 29300 1709
rect 28972 1063 29012 1072
rect 29260 80 29300 1660
rect 29356 1532 29396 1996
rect 29548 1616 29588 3424
rect 30220 3464 30260 3473
rect 29836 2372 29876 2381
rect 29836 1952 29876 2332
rect 29836 1903 29876 1912
rect 30220 1784 30260 3424
rect 30604 3464 30644 3473
rect 30316 3212 30356 3221
rect 30316 2792 30356 3172
rect 30316 2743 30356 2752
rect 30316 2456 30356 2465
rect 30316 1952 30356 2416
rect 30316 1903 30356 1912
rect 30220 1735 30260 1744
rect 29548 1567 29588 1576
rect 29644 1700 29684 1709
rect 29356 1483 29396 1492
rect 29644 80 29684 1660
rect 30028 1700 30068 1709
rect 30028 80 30068 1660
rect 30412 1700 30452 1709
rect 30412 80 30452 1660
rect 30604 1448 30644 3424
rect 30988 3464 31028 3760
rect 31372 3749 31412 3844
rect 30988 3415 31028 3424
rect 32428 3632 32468 3641
rect 32428 3464 32468 3592
rect 32428 3415 32468 3424
rect 32908 3464 32948 4264
rect 32908 3415 32948 3424
rect 31180 3380 31220 3389
rect 31180 3245 31220 3340
rect 32236 3296 32276 3305
rect 31660 3212 31700 3221
rect 31660 2960 31700 3172
rect 31660 2911 31700 2920
rect 31468 2708 31508 2717
rect 31468 1952 31508 2668
rect 31468 1903 31508 1912
rect 31660 2624 31700 2633
rect 30604 1399 30644 1408
rect 30796 1700 30836 1709
rect 30796 80 30836 1660
rect 31180 1700 31220 1709
rect 31180 80 31220 1660
rect 31564 1700 31604 1709
rect 31564 80 31604 1660
rect 31660 1700 31700 2584
rect 32236 1952 32276 3256
rect 32236 1903 32276 1912
rect 32524 3212 32564 3221
rect 32524 1952 32564 3172
rect 32524 1903 32564 1912
rect 33004 3212 33044 3221
rect 33004 1952 33044 3172
rect 33100 3128 33140 3137
rect 33100 3044 33140 3088
rect 33196 3128 33236 7708
rect 34828 8000 34868 8009
rect 34828 7328 34868 7960
rect 34924 7916 34964 7925
rect 35308 7916 35348 7925
rect 34964 7876 35308 7916
rect 34924 7867 34964 7876
rect 35308 7867 35348 7876
rect 38092 7664 38132 8044
rect 38092 7615 38132 7624
rect 35168 7580 35536 7589
rect 35208 7540 35250 7580
rect 35290 7540 35332 7580
rect 35372 7540 35414 7580
rect 35454 7540 35496 7580
rect 35168 7531 35536 7540
rect 34828 7279 34868 7288
rect 33928 6824 34296 6833
rect 33968 6784 34010 6824
rect 34050 6784 34092 6824
rect 34132 6784 34174 6824
rect 34214 6784 34256 6824
rect 33928 6775 34296 6784
rect 35788 6488 35828 6497
rect 35168 6068 35536 6077
rect 35208 6028 35250 6068
rect 35290 6028 35332 6068
rect 35372 6028 35414 6068
rect 35454 6028 35496 6068
rect 35168 6019 35536 6028
rect 35788 5816 35828 6448
rect 33928 5312 34296 5321
rect 33968 5272 34010 5312
rect 34050 5272 34092 5312
rect 34132 5272 34174 5312
rect 34214 5272 34256 5312
rect 33928 5263 34296 5272
rect 35168 4556 35536 4565
rect 35208 4516 35250 4556
rect 35290 4516 35332 4556
rect 35372 4516 35414 4556
rect 35454 4516 35496 4556
rect 35168 4507 35536 4516
rect 35020 4136 35060 4145
rect 33928 3800 34296 3809
rect 33968 3760 34010 3800
rect 34050 3760 34092 3800
rect 34132 3760 34174 3800
rect 34214 3760 34256 3800
rect 33928 3751 34296 3760
rect 33772 3716 33812 3725
rect 33772 3464 33812 3676
rect 33772 3415 33812 3424
rect 35020 3464 35060 4096
rect 35020 3415 35060 3424
rect 35212 3464 35252 3473
rect 35212 3380 35252 3424
rect 35212 3329 35252 3340
rect 33196 3079 33236 3088
rect 33388 3212 33428 3221
rect 33100 2993 33140 3004
rect 33004 1903 33044 1912
rect 33388 1952 33428 3172
rect 34348 3212 34388 3221
rect 34252 2624 34292 2633
rect 34252 2540 34292 2584
rect 34252 2489 34292 2500
rect 33928 2288 34296 2297
rect 33968 2248 34010 2288
rect 34050 2248 34092 2288
rect 34132 2248 34174 2288
rect 34214 2248 34256 2288
rect 33928 2239 34296 2248
rect 33388 1903 33428 1912
rect 34348 1952 34388 3172
rect 35020 3212 35060 3221
rect 34348 1903 34388 1912
rect 34540 2624 34580 2633
rect 31660 1651 31700 1660
rect 31948 1700 31988 1709
rect 31948 80 31988 1660
rect 32332 1700 32372 1709
rect 32332 80 32372 1660
rect 32716 1700 32756 1709
rect 33100 1700 33140 1709
rect 32716 80 32756 1660
rect 33004 1660 33100 1700
rect 33004 440 33044 1660
rect 33100 1651 33140 1660
rect 33484 1700 33524 1709
rect 33004 400 33140 440
rect 33100 80 33140 400
rect 33484 80 33524 1660
rect 33868 1700 33908 1709
rect 33868 80 33908 1660
rect 34252 1700 34292 1709
rect 34252 80 34292 1660
rect 34540 272 34580 2584
rect 34924 2120 34964 2129
rect 34540 223 34580 232
rect 34636 1700 34676 1709
rect 34636 80 34676 1660
rect 34924 1532 34964 2080
rect 35020 1952 35060 3172
rect 35692 3212 35732 3221
rect 35168 3044 35536 3053
rect 35208 3004 35250 3044
rect 35290 3004 35332 3044
rect 35372 3004 35414 3044
rect 35454 3004 35496 3044
rect 35168 2995 35536 3004
rect 35020 1903 35060 1912
rect 35692 1952 35732 3172
rect 35788 2792 35828 5776
rect 36940 4052 36980 4061
rect 36940 3464 36980 4012
rect 37804 3968 37844 3977
rect 36940 3415 36980 3424
rect 37708 3464 37748 3473
rect 35788 2743 35828 2752
rect 36076 3212 36116 3221
rect 35692 1903 35732 1912
rect 36076 1952 36116 3172
rect 36460 3212 36500 3221
rect 36076 1903 36116 1912
rect 36268 2624 36308 2633
rect 35980 1868 36020 1877
rect 34924 1483 34964 1492
rect 35020 1700 35060 1709
rect 35020 80 35060 1660
rect 35596 1700 35636 1709
rect 35168 1532 35536 1541
rect 35208 1492 35250 1532
rect 35290 1492 35332 1532
rect 35372 1492 35414 1532
rect 35454 1492 35496 1532
rect 35168 1483 35536 1492
rect 35596 188 35636 1660
rect 35404 148 35636 188
rect 35788 1700 35828 1709
rect 35404 80 35444 148
rect 35788 80 35828 1660
rect 35980 1616 36020 1828
rect 35980 1567 36020 1576
rect 36172 1700 36212 1709
rect 36172 80 36212 1660
rect 36268 356 36308 2584
rect 36460 1952 36500 3172
rect 37516 3212 37556 3221
rect 37516 2036 37556 3172
rect 37708 2876 37748 3424
rect 37708 2827 37748 2836
rect 37516 1987 37556 1996
rect 37612 2456 37652 2465
rect 36460 1903 36500 1912
rect 37612 1952 37652 2416
rect 37612 1903 37652 1912
rect 37804 1868 37844 3928
rect 38380 3884 38420 3893
rect 38380 1952 38420 3844
rect 41740 3212 41780 3221
rect 40012 2876 40052 2885
rect 38380 1903 38420 1912
rect 39148 2708 39188 2717
rect 39148 1952 39188 2668
rect 39724 2624 39764 2633
rect 39436 2456 39476 2465
rect 39436 2036 39476 2416
rect 39436 1987 39476 1996
rect 39148 1903 39188 1912
rect 39532 1952 39572 1961
rect 37804 1819 37844 1828
rect 37996 1868 38036 1877
rect 36268 307 36308 316
rect 36556 1700 36596 1709
rect 36556 80 36596 1660
rect 36940 1700 36980 1709
rect 36940 80 36980 1660
rect 37324 1700 37364 1709
rect 37324 80 37364 1660
rect 37708 1700 37748 1709
rect 37708 80 37748 1660
rect 37900 1532 37940 1541
rect 37996 1532 38036 1828
rect 37940 1492 38036 1532
rect 38092 1700 38132 1709
rect 37900 1483 37940 1492
rect 38092 80 38132 1660
rect 38476 1700 38516 1709
rect 38476 80 38516 1660
rect 38860 1700 38900 1709
rect 38860 80 38900 1660
rect 39244 1700 39284 1709
rect 39244 80 39284 1660
rect 39532 1616 39572 1912
rect 39532 1567 39572 1576
rect 39628 1700 39668 1709
rect 39628 80 39668 1660
rect 39724 356 39764 2584
rect 40012 2036 40052 2836
rect 40012 1987 40052 1996
rect 40300 2708 40340 2717
rect 40300 1952 40340 2668
rect 41740 2456 41780 3172
rect 41740 2407 41780 2416
rect 42412 2792 42452 2801
rect 40300 1903 40340 1912
rect 41068 2372 41108 2381
rect 41068 1952 41108 2332
rect 41068 1903 41108 1912
rect 41452 2204 41492 2213
rect 41452 1952 41492 2164
rect 41452 1903 41492 1912
rect 41836 2120 41876 2129
rect 41836 1952 41876 2080
rect 42412 2120 42452 2752
rect 42412 2071 42452 2080
rect 41836 1903 41876 1912
rect 42220 2036 42260 2047
rect 42220 1952 42260 1996
rect 42220 1903 42260 1912
rect 42604 1952 42644 1961
rect 42604 1817 42644 1912
rect 39724 307 39764 316
rect 40012 1700 40052 1709
rect 40012 80 40052 1660
rect 40396 1700 40436 1709
rect 40396 80 40436 1660
rect 40780 1700 40820 1709
rect 40780 80 40820 1660
rect 41164 1700 41204 1709
rect 41164 80 41204 1660
rect 41548 1700 41588 1709
rect 41548 80 41588 1660
rect 41932 1700 41972 1709
rect 41932 80 41972 1660
rect 42316 1700 42356 1709
rect 42316 80 42356 1660
rect 42700 80 42740 9388
rect 43084 80 43124 9640
rect 43276 8756 43316 9892
rect 43372 9680 43412 10144
rect 43372 9631 43412 9640
rect 43948 10100 43988 10109
rect 43948 9680 43988 10060
rect 43948 9631 43988 9640
rect 43276 8707 43316 8716
rect 43468 9596 43508 9605
rect 43468 80 43508 9556
rect 43852 9596 43892 9605
rect 43564 9344 43604 9353
rect 43564 8756 43604 9304
rect 43564 8707 43604 8716
rect 43852 80 43892 9556
rect 44140 9428 44180 9437
rect 44140 9092 44180 9388
rect 44620 9260 44660 10228
rect 44908 9680 44948 10480
rect 44908 9631 44948 9640
rect 46156 9680 46196 10564
rect 46540 10436 46580 12100
rect 46540 10387 46580 10396
rect 49036 10436 49076 12100
rect 50956 11192 50996 11201
rect 50288 10604 50656 10613
rect 50328 10564 50370 10604
rect 50410 10564 50452 10604
rect 50492 10564 50534 10604
rect 50574 10564 50616 10604
rect 50288 10555 50656 10564
rect 49036 10387 49076 10396
rect 46636 10184 46676 10193
rect 46156 9631 46196 9640
rect 46348 9932 46388 9941
rect 44620 9211 44660 9220
rect 46156 9428 46196 9437
rect 45964 9176 46004 9185
rect 46156 9176 46196 9388
rect 46004 9136 46100 9176
rect 45964 9127 46004 9136
rect 44140 9043 44180 9052
rect 44620 9008 44660 9017
rect 44236 7748 44276 7757
rect 44236 4304 44276 7708
rect 44236 4255 44276 4264
rect 44236 104 44276 113
rect 14092 55 14132 64
rect 14264 0 14344 80
rect 14648 0 14728 80
rect 15032 0 15112 80
rect 15416 0 15496 80
rect 15800 0 15880 80
rect 16184 0 16264 80
rect 16568 0 16648 80
rect 16952 0 17032 80
rect 17336 0 17416 80
rect 17720 0 17800 80
rect 18104 0 18184 80
rect 18488 0 18568 80
rect 18872 0 18952 80
rect 19256 0 19336 80
rect 19640 0 19720 80
rect 20024 0 20104 80
rect 20408 0 20488 80
rect 20792 0 20872 80
rect 21176 0 21256 80
rect 21560 0 21640 80
rect 21944 0 22024 80
rect 22328 0 22408 80
rect 22712 0 22792 80
rect 23096 0 23176 80
rect 23480 0 23560 80
rect 23864 0 23944 80
rect 24248 0 24328 80
rect 24632 0 24712 80
rect 25016 0 25096 80
rect 25400 0 25480 80
rect 25784 0 25864 80
rect 26168 0 26248 80
rect 26552 0 26632 80
rect 26936 0 27016 80
rect 27320 0 27400 80
rect 27704 0 27784 80
rect 28088 0 28168 80
rect 28472 0 28552 80
rect 28856 0 28936 80
rect 29240 0 29320 80
rect 29624 0 29704 80
rect 30008 0 30088 80
rect 30392 0 30472 80
rect 30776 0 30856 80
rect 31160 0 31240 80
rect 31544 0 31624 80
rect 31928 0 32008 80
rect 32312 0 32392 80
rect 32696 0 32776 80
rect 33080 0 33160 80
rect 33464 0 33544 80
rect 33848 0 33928 80
rect 34232 0 34312 80
rect 34616 0 34696 80
rect 35000 0 35080 80
rect 35384 0 35464 80
rect 35768 0 35848 80
rect 36152 0 36232 80
rect 36536 0 36616 80
rect 36920 0 37000 80
rect 37304 0 37384 80
rect 37688 0 37768 80
rect 38072 0 38152 80
rect 38456 0 38536 80
rect 38840 0 38920 80
rect 39224 0 39304 80
rect 39608 0 39688 80
rect 39992 0 40072 80
rect 40376 0 40456 80
rect 40760 0 40840 80
rect 41144 0 41224 80
rect 41528 0 41608 80
rect 41912 0 41992 80
rect 42296 0 42376 80
rect 42680 0 42760 80
rect 43064 0 43144 80
rect 43448 0 43528 80
rect 43832 0 43912 80
rect 44216 64 44236 80
rect 44620 80 44660 8968
rect 44716 3380 44756 3389
rect 44716 2792 44756 3340
rect 46060 2900 46100 9136
rect 46156 9127 46196 9136
rect 46156 9008 46196 9017
rect 46156 8756 46196 8968
rect 46156 8707 46196 8716
rect 46348 8756 46388 9892
rect 46636 9680 46676 10144
rect 48172 10184 48212 10193
rect 47500 10100 47540 10109
rect 47500 9848 47540 10060
rect 47500 9799 47540 9808
rect 46636 9631 46676 9640
rect 48172 9680 48212 10144
rect 48172 9631 48212 9640
rect 48940 10184 48980 10193
rect 48940 9680 48980 10144
rect 50092 10184 50132 10193
rect 49048 9848 49416 9857
rect 49088 9808 49130 9848
rect 49170 9808 49212 9848
rect 49252 9808 49294 9848
rect 49334 9808 49376 9848
rect 49048 9799 49416 9808
rect 48940 9631 48980 9640
rect 47692 9596 47732 9605
rect 47212 9428 47252 9437
rect 47212 9260 47252 9388
rect 47212 9211 47252 9220
rect 47308 9176 47348 9185
rect 46348 8707 46388 8716
rect 47212 8924 47252 8933
rect 46924 8672 46964 8681
rect 46060 2860 46580 2900
rect 44716 2743 44756 2752
rect 46156 272 46196 281
rect 45004 188 45044 197
rect 45004 80 45044 148
rect 45772 188 45812 197
rect 45388 104 45428 113
rect 44276 64 44296 80
rect 44216 0 44296 64
rect 44600 0 44680 80
rect 44984 0 45064 80
rect 45368 64 45388 80
rect 45772 80 45812 148
rect 46156 80 46196 232
rect 46540 80 46580 2860
rect 46924 80 46964 8632
rect 47212 3464 47252 8884
rect 47212 3415 47252 3424
rect 47308 80 47348 9136
rect 47500 6236 47540 6245
rect 47500 4220 47540 6196
rect 47500 4171 47540 4180
rect 47692 80 47732 9556
rect 49996 9512 50036 9521
rect 48460 9428 48500 9437
rect 48076 9344 48116 9353
rect 48076 80 48116 9304
rect 48460 80 48500 9388
rect 49612 9428 49652 9437
rect 48940 9260 48980 9269
rect 48844 9092 48884 9101
rect 48844 80 48884 9052
rect 48940 2120 48980 9220
rect 49048 8336 49416 8345
rect 49088 8296 49130 8336
rect 49170 8296 49212 8336
rect 49252 8296 49294 8336
rect 49334 8296 49376 8336
rect 49048 8287 49416 8296
rect 49048 6824 49416 6833
rect 49088 6784 49130 6824
rect 49170 6784 49212 6824
rect 49252 6784 49294 6824
rect 49334 6784 49376 6824
rect 49048 6775 49416 6784
rect 49048 5312 49416 5321
rect 49088 5272 49130 5312
rect 49170 5272 49212 5312
rect 49252 5272 49294 5312
rect 49334 5272 49376 5312
rect 49048 5263 49416 5272
rect 49048 3800 49416 3809
rect 49088 3760 49130 3800
rect 49170 3760 49212 3800
rect 49252 3760 49294 3800
rect 49334 3760 49376 3800
rect 49048 3751 49416 3760
rect 49420 3296 49460 3305
rect 49420 2540 49460 3256
rect 49420 2491 49460 2500
rect 49516 2960 49556 2969
rect 49048 2288 49416 2297
rect 49088 2248 49130 2288
rect 49170 2248 49212 2288
rect 49252 2248 49294 2288
rect 49334 2248 49376 2288
rect 49048 2239 49416 2248
rect 48940 2080 49268 2120
rect 49228 80 49268 2080
rect 49516 1952 49556 2920
rect 49516 1903 49556 1912
rect 49612 80 49652 9388
rect 49708 2624 49748 2633
rect 49708 1784 49748 2584
rect 49708 1735 49748 1744
rect 49996 80 50036 9472
rect 50092 9260 50132 10144
rect 50380 9932 50420 9941
rect 50380 9797 50420 9892
rect 50956 9680 50996 11152
rect 51052 10856 51092 10865
rect 51052 10436 51092 10816
rect 51244 10520 51284 10529
rect 51436 10520 51476 10529
rect 51284 10480 51436 10520
rect 51244 10471 51284 10480
rect 51436 10471 51476 10480
rect 51052 10387 51092 10396
rect 51532 10436 51572 12100
rect 51532 10387 51572 10396
rect 51052 10184 51092 10193
rect 51052 10016 51092 10144
rect 51052 9967 51092 9976
rect 51436 10184 51476 10193
rect 51436 9932 51476 10144
rect 51628 10184 51668 10193
rect 51436 9883 51476 9892
rect 51532 10100 51572 10109
rect 50956 9631 50996 9640
rect 51532 9596 51572 10060
rect 51628 9680 51668 10144
rect 51628 9631 51668 9640
rect 51532 9547 51572 9556
rect 50092 9211 50132 9220
rect 50956 9512 50996 9521
rect 50288 9092 50656 9101
rect 50328 9052 50370 9092
rect 50410 9052 50452 9092
rect 50492 9052 50534 9092
rect 50574 9052 50616 9092
rect 50288 9043 50656 9052
rect 50288 7580 50656 7589
rect 50328 7540 50370 7580
rect 50410 7540 50452 7580
rect 50492 7540 50534 7580
rect 50574 7540 50616 7580
rect 50288 7531 50656 7540
rect 50288 6068 50656 6077
rect 50328 6028 50370 6068
rect 50410 6028 50452 6068
rect 50492 6028 50534 6068
rect 50574 6028 50616 6068
rect 50288 6019 50656 6028
rect 50288 4556 50656 4565
rect 50328 4516 50370 4556
rect 50410 4516 50452 4556
rect 50492 4516 50534 4556
rect 50574 4516 50616 4556
rect 50288 4507 50656 4516
rect 50860 4136 50900 4145
rect 50188 3296 50228 3305
rect 50188 2624 50228 3256
rect 50860 3212 50900 4096
rect 50860 3163 50900 3172
rect 50288 3044 50656 3053
rect 50328 3004 50370 3044
rect 50410 3004 50452 3044
rect 50492 3004 50534 3044
rect 50574 3004 50616 3044
rect 50288 2995 50656 3004
rect 50188 1868 50228 2584
rect 50188 1819 50228 1828
rect 50288 1532 50656 1541
rect 50328 1492 50370 1532
rect 50410 1492 50452 1532
rect 50492 1492 50534 1532
rect 50574 1492 50616 1532
rect 50288 1483 50656 1492
rect 50380 104 50420 113
rect 45428 64 45448 80
rect 45368 0 45448 64
rect 45752 0 45832 80
rect 46136 0 46216 80
rect 46520 0 46600 80
rect 46904 0 46984 80
rect 47288 0 47368 80
rect 47672 0 47752 80
rect 48056 0 48136 80
rect 48440 0 48520 80
rect 48824 0 48904 80
rect 49208 0 49288 80
rect 49592 0 49672 80
rect 49976 0 50056 80
rect 50360 64 50380 80
rect 50956 104 50996 9472
rect 51628 9512 51668 9521
rect 51628 8168 51668 9472
rect 52684 9260 52724 9269
rect 52684 8840 52724 9220
rect 52684 8791 52724 8800
rect 51628 8119 51668 8128
rect 51820 8672 51860 8681
rect 51820 7076 51860 8632
rect 53164 8672 53204 8681
rect 53164 8168 53204 8632
rect 53164 8119 53204 8128
rect 53164 7664 53204 7673
rect 52012 7580 52052 7589
rect 51820 7027 51860 7036
rect 51916 7160 51956 7169
rect 51436 6908 51476 6917
rect 51436 4976 51476 6868
rect 51436 4927 51476 4936
rect 51820 6488 51860 6497
rect 51820 4892 51860 6448
rect 51916 5396 51956 7120
rect 51916 5347 51956 5356
rect 51820 4843 51860 4852
rect 52012 4136 52052 7540
rect 53164 7496 53204 7624
rect 53164 7447 53204 7456
rect 52012 4087 52052 4096
rect 52108 6068 52148 6077
rect 51436 3212 51476 3221
rect 51436 1952 51476 3172
rect 52108 2624 52148 6028
rect 52108 2575 52148 2584
rect 51436 1903 51476 1912
rect 52588 2456 52628 2465
rect 52300 1784 52340 1793
rect 51916 1616 51956 1625
rect 51916 1112 51956 1576
rect 51916 1063 51956 1072
rect 52300 776 52340 1744
rect 52588 1448 52628 2416
rect 52588 1399 52628 1408
rect 52300 727 52340 736
rect 50420 64 50440 80
rect 50360 0 50440 64
rect 50956 55 50996 64
<< via3 >>
rect 4928 10564 4968 10604
rect 5010 10564 5050 10604
rect 5092 10564 5132 10604
rect 5174 10564 5214 10604
rect 5256 10564 5296 10604
rect 3688 9808 3728 9848
rect 3770 9808 3810 9848
rect 3852 9808 3892 9848
rect 3934 9808 3974 9848
rect 4016 9808 4056 9848
rect 4928 9052 4968 9092
rect 5010 9052 5050 9092
rect 5092 9052 5132 9092
rect 5174 9052 5214 9092
rect 5256 9052 5296 9092
rect 3688 8296 3728 8336
rect 3770 8296 3810 8336
rect 3852 8296 3892 8336
rect 3934 8296 3974 8336
rect 4016 8296 4056 8336
rect 4928 7540 4968 7580
rect 5010 7540 5050 7580
rect 5092 7540 5132 7580
rect 5174 7540 5214 7580
rect 5256 7540 5296 7580
rect 3688 6784 3728 6824
rect 3770 6784 3810 6824
rect 3852 6784 3892 6824
rect 3934 6784 3974 6824
rect 4016 6784 4056 6824
rect 4928 6028 4968 6068
rect 5010 6028 5050 6068
rect 5092 6028 5132 6068
rect 5174 6028 5214 6068
rect 5256 6028 5296 6068
rect 3688 5272 3728 5312
rect 3770 5272 3810 5312
rect 3852 5272 3892 5312
rect 3934 5272 3974 5312
rect 4016 5272 4056 5312
rect 4928 4516 4968 4556
rect 5010 4516 5050 4556
rect 5092 4516 5132 4556
rect 5174 4516 5214 4556
rect 5256 4516 5296 4556
rect 3688 3760 3728 3800
rect 3770 3760 3810 3800
rect 3852 3760 3892 3800
rect 3934 3760 3974 3800
rect 4016 3760 4056 3800
rect 1420 2752 1460 2792
rect 1420 2416 1460 2456
rect 3688 2248 3728 2288
rect 3770 2248 3810 2288
rect 3852 2248 3892 2288
rect 3934 2248 3974 2288
rect 4016 2248 4056 2288
rect 1420 1744 1460 1784
rect 1420 1408 1460 1448
rect 1420 1072 1460 1112
rect 3148 1828 3188 1868
rect 4928 3004 4968 3044
rect 5010 3004 5050 3044
rect 5092 3004 5132 3044
rect 5174 3004 5214 3044
rect 5256 3004 5296 3044
rect 4928 1492 4968 1532
rect 5010 1492 5050 1532
rect 5092 1492 5132 1532
rect 5174 1492 5214 1532
rect 5256 1492 5296 1532
rect 4684 484 4724 524
rect 5068 400 5108 440
rect 8524 4096 8564 4136
rect 8140 2920 8180 2960
rect 7372 2584 7412 2624
rect 7756 1576 7796 1616
rect 10060 316 10100 356
rect 12364 2500 12404 2540
rect 11980 232 12020 272
rect 13132 1660 13172 1700
rect 13900 3508 13940 3548
rect 20048 10564 20088 10604
rect 20130 10564 20170 10604
rect 20212 10564 20252 10604
rect 20294 10564 20334 10604
rect 20376 10564 20416 10604
rect 18808 9808 18848 9848
rect 18890 9808 18930 9848
rect 18972 9808 19012 9848
rect 19054 9808 19094 9848
rect 19136 9808 19176 9848
rect 18700 9472 18740 9512
rect 20140 9220 20180 9260
rect 20048 9052 20088 9092
rect 20130 9052 20170 9092
rect 20212 9052 20252 9092
rect 20294 9052 20334 9092
rect 20376 9052 20416 9092
rect 18808 8296 18848 8336
rect 18890 8296 18930 8336
rect 18972 8296 19012 8336
rect 19054 8296 19094 8336
rect 19136 8296 19176 8336
rect 20048 7540 20088 7580
rect 20130 7540 20170 7580
rect 20212 7540 20252 7580
rect 20294 7540 20334 7580
rect 20376 7540 20416 7580
rect 18808 6784 18848 6824
rect 18890 6784 18930 6824
rect 18972 6784 19012 6824
rect 19054 6784 19094 6824
rect 19136 6784 19176 6824
rect 20048 6028 20088 6068
rect 20130 6028 20170 6068
rect 20212 6028 20252 6068
rect 20294 6028 20334 6068
rect 20376 6028 20416 6068
rect 18808 5272 18848 5312
rect 18890 5272 18930 5312
rect 18972 5272 19012 5312
rect 19054 5272 19094 5312
rect 19136 5272 19176 5312
rect 14188 2836 14228 2876
rect 14092 64 14132 104
rect 14380 1492 14420 1532
rect 14668 1996 14708 2036
rect 15052 2836 15092 2876
rect 15340 2164 15380 2204
rect 15628 2332 15668 2372
rect 16300 3844 16340 3884
rect 15724 2080 15764 2120
rect 16876 2836 16916 2876
rect 17260 3508 17300 3548
rect 20048 4516 20088 4556
rect 20130 4516 20170 4556
rect 20212 4516 20252 4556
rect 20294 4516 20334 4556
rect 20376 4516 20416 4556
rect 18412 316 18452 356
rect 18808 3760 18848 3800
rect 18890 3760 18930 3800
rect 18972 3760 19012 3800
rect 19054 3760 19094 3800
rect 19136 3760 19176 3800
rect 18700 2668 18740 2708
rect 19372 2668 19412 2708
rect 18808 2248 18848 2288
rect 18890 2248 18930 2288
rect 18972 2248 19012 2288
rect 19054 2248 19094 2288
rect 19136 2248 19176 2288
rect 20140 3676 20180 3716
rect 20620 3592 20660 3632
rect 20048 3004 20088 3044
rect 20130 3004 20170 3044
rect 20212 3004 20252 3044
rect 20294 3004 20334 3044
rect 20376 3004 20416 3044
rect 19564 1912 19604 1952
rect 19372 1828 19412 1868
rect 19852 1912 19892 1952
rect 19852 1492 19892 1532
rect 20428 2332 20468 2372
rect 20048 1492 20088 1532
rect 20130 1492 20170 1532
rect 20212 1492 20252 1532
rect 20294 1492 20334 1532
rect 20376 1492 20416 1532
rect 20620 2668 20660 2708
rect 20716 1576 20756 1616
rect 21196 2668 21236 2708
rect 21196 316 21236 356
rect 35168 10564 35208 10604
rect 35250 10564 35290 10604
rect 35332 10564 35372 10604
rect 35414 10564 35454 10604
rect 35496 10564 35536 10604
rect 22636 4012 22676 4052
rect 21580 3424 21620 3464
rect 21388 2332 21428 2372
rect 21772 2668 21812 2708
rect 22924 4180 22964 4220
rect 23212 4180 23252 4220
rect 23116 4012 23156 4052
rect 22924 3760 22964 3800
rect 23308 3844 23348 3884
rect 23116 3592 23156 3632
rect 22732 3508 22772 3548
rect 23212 3508 23252 3548
rect 22540 2248 22580 2288
rect 22828 484 22868 524
rect 23308 400 23348 440
rect 24940 2248 24980 2288
rect 28300 9220 28340 9260
rect 25900 2920 25940 2960
rect 25708 1492 25748 1532
rect 33928 9808 33968 9848
rect 34010 9808 34050 9848
rect 34092 9808 34132 9848
rect 34174 9808 34214 9848
rect 34256 9808 34296 9848
rect 43276 9892 43316 9932
rect 35168 9052 35208 9092
rect 35250 9052 35290 9092
rect 35332 9052 35372 9092
rect 35414 9052 35454 9092
rect 35496 9052 35536 9092
rect 33928 8296 33968 8336
rect 34010 8296 34050 8336
rect 34092 8296 34132 8336
rect 34174 8296 34214 8336
rect 34256 8296 34296 8336
rect 28012 4096 28052 4136
rect 28300 3760 28340 3800
rect 28396 3676 28436 3716
rect 26668 2668 26708 2708
rect 28108 2668 28148 2708
rect 28108 1828 28148 1868
rect 28780 2584 28820 2624
rect 31372 3844 31412 3884
rect 30220 3676 30260 3716
rect 29548 3424 29588 3464
rect 28972 1072 29012 1112
rect 30220 1744 30260 1784
rect 31180 3340 31220 3380
rect 30604 1408 30644 1448
rect 33100 3088 33140 3128
rect 35168 7540 35208 7580
rect 35250 7540 35290 7580
rect 35332 7540 35372 7580
rect 35414 7540 35454 7580
rect 35496 7540 35536 7580
rect 33928 6784 33968 6824
rect 34010 6784 34050 6824
rect 34092 6784 34132 6824
rect 34174 6784 34214 6824
rect 34256 6784 34296 6824
rect 35168 6028 35208 6068
rect 35250 6028 35290 6068
rect 35332 6028 35372 6068
rect 35414 6028 35454 6068
rect 35496 6028 35536 6068
rect 33928 5272 33968 5312
rect 34010 5272 34050 5312
rect 34092 5272 34132 5312
rect 34174 5272 34214 5312
rect 34256 5272 34296 5312
rect 35168 4516 35208 4556
rect 35250 4516 35290 4556
rect 35332 4516 35372 4556
rect 35414 4516 35454 4556
rect 35496 4516 35536 4556
rect 33928 3760 33968 3800
rect 34010 3760 34050 3800
rect 34092 3760 34132 3800
rect 34174 3760 34214 3800
rect 34256 3760 34296 3800
rect 33772 3676 33812 3716
rect 35212 3340 35252 3380
rect 33196 3088 33236 3128
rect 34252 2500 34292 2540
rect 33928 2248 33968 2288
rect 34010 2248 34050 2288
rect 34092 2248 34132 2288
rect 34174 2248 34214 2288
rect 34256 2248 34296 2288
rect 31660 1660 31700 1700
rect 34540 232 34580 272
rect 35168 3004 35208 3044
rect 35250 3004 35290 3044
rect 35332 3004 35372 3044
rect 35414 3004 35454 3044
rect 35496 3004 35536 3044
rect 35788 2752 35828 2792
rect 35980 1828 36020 1868
rect 35168 1492 35208 1532
rect 35250 1492 35290 1532
rect 35332 1492 35372 1532
rect 35414 1492 35454 1532
rect 35496 1492 35536 1532
rect 38380 3844 38420 3884
rect 40012 2836 40052 2876
rect 40300 2668 40340 2708
rect 41740 2416 41780 2456
rect 41068 2332 41108 2372
rect 41452 2164 41492 2204
rect 41836 2080 41876 2120
rect 42220 1996 42260 2036
rect 42604 1912 42644 1952
rect 39724 316 39764 356
rect 50288 10564 50328 10604
rect 50370 10564 50410 10604
rect 50452 10564 50492 10604
rect 50534 10564 50574 10604
rect 50616 10564 50656 10604
rect 44236 64 44276 104
rect 49048 9808 49088 9848
rect 49130 9808 49170 9848
rect 49212 9808 49252 9848
rect 49294 9808 49334 9848
rect 49376 9808 49416 9848
rect 45004 148 45044 188
rect 49048 8296 49088 8336
rect 49130 8296 49170 8336
rect 49212 8296 49252 8336
rect 49294 8296 49334 8336
rect 49376 8296 49416 8336
rect 49048 6784 49088 6824
rect 49130 6784 49170 6824
rect 49212 6784 49252 6824
rect 49294 6784 49334 6824
rect 49376 6784 49416 6824
rect 49048 5272 49088 5312
rect 49130 5272 49170 5312
rect 49212 5272 49252 5312
rect 49294 5272 49334 5312
rect 49376 5272 49416 5312
rect 49048 3760 49088 3800
rect 49130 3760 49170 3800
rect 49212 3760 49252 3800
rect 49294 3760 49334 3800
rect 49376 3760 49416 3800
rect 49048 2248 49088 2288
rect 49130 2248 49170 2288
rect 49212 2248 49252 2288
rect 49294 2248 49334 2288
rect 49376 2248 49416 2288
rect 50380 9892 50420 9932
rect 50288 9052 50328 9092
rect 50370 9052 50410 9092
rect 50452 9052 50492 9092
rect 50534 9052 50574 9092
rect 50616 9052 50656 9092
rect 50288 7540 50328 7580
rect 50370 7540 50410 7580
rect 50452 7540 50492 7580
rect 50534 7540 50574 7580
rect 50616 7540 50656 7580
rect 50288 6028 50328 6068
rect 50370 6028 50410 6068
rect 50452 6028 50492 6068
rect 50534 6028 50574 6068
rect 50616 6028 50656 6068
rect 50288 4516 50328 4556
rect 50370 4516 50410 4556
rect 50452 4516 50492 4556
rect 50534 4516 50574 4556
rect 50616 4516 50656 4556
rect 50288 3004 50328 3044
rect 50370 3004 50410 3044
rect 50452 3004 50492 3044
rect 50534 3004 50574 3044
rect 50616 3004 50656 3044
rect 50288 1492 50328 1532
rect 50370 1492 50410 1532
rect 50452 1492 50492 1532
rect 50534 1492 50574 1532
rect 50616 1492 50656 1532
rect 50380 64 50420 104
rect 50956 64 50996 104
<< metal4 >>
rect 4919 10564 4928 10604
rect 4968 10564 5010 10604
rect 5050 10564 5092 10604
rect 5132 10564 5174 10604
rect 5214 10564 5256 10604
rect 5296 10564 5305 10604
rect 20039 10564 20048 10604
rect 20088 10564 20130 10604
rect 20170 10564 20212 10604
rect 20252 10564 20294 10604
rect 20334 10564 20376 10604
rect 20416 10564 20425 10604
rect 35159 10564 35168 10604
rect 35208 10564 35250 10604
rect 35290 10564 35332 10604
rect 35372 10564 35414 10604
rect 35454 10564 35496 10604
rect 35536 10564 35545 10604
rect 50279 10564 50288 10604
rect 50328 10564 50370 10604
rect 50410 10564 50452 10604
rect 50492 10564 50534 10604
rect 50574 10564 50616 10604
rect 50656 10564 50665 10604
rect 43267 9892 43276 9932
rect 43316 9892 50380 9932
rect 50420 9892 50429 9932
rect 3679 9808 3688 9848
rect 3728 9808 3770 9848
rect 3810 9808 3852 9848
rect 3892 9808 3934 9848
rect 3974 9808 4016 9848
rect 4056 9808 4065 9848
rect 18799 9808 18808 9848
rect 18848 9808 18890 9848
rect 18930 9808 18972 9848
rect 19012 9808 19054 9848
rect 19094 9808 19136 9848
rect 19176 9808 19185 9848
rect 33919 9808 33928 9848
rect 33968 9808 34010 9848
rect 34050 9808 34092 9848
rect 34132 9808 34174 9848
rect 34214 9808 34256 9848
rect 34296 9808 34305 9848
rect 49039 9808 49048 9848
rect 49088 9808 49130 9848
rect 49170 9808 49212 9848
rect 49252 9808 49294 9848
rect 49334 9808 49376 9848
rect 49416 9808 49425 9848
rect 18691 9472 18700 9512
rect 18740 9472 19468 9512
rect 19508 9472 19517 9512
rect 20131 9220 20140 9260
rect 20180 9220 28300 9260
rect 28340 9220 28349 9260
rect 4919 9052 4928 9092
rect 4968 9052 5010 9092
rect 5050 9052 5092 9092
rect 5132 9052 5174 9092
rect 5214 9052 5256 9092
rect 5296 9052 5305 9092
rect 20039 9052 20048 9092
rect 20088 9052 20130 9092
rect 20170 9052 20212 9092
rect 20252 9052 20294 9092
rect 20334 9052 20376 9092
rect 20416 9052 20425 9092
rect 35159 9052 35168 9092
rect 35208 9052 35250 9092
rect 35290 9052 35332 9092
rect 35372 9052 35414 9092
rect 35454 9052 35496 9092
rect 35536 9052 35545 9092
rect 50279 9052 50288 9092
rect 50328 9052 50370 9092
rect 50410 9052 50452 9092
rect 50492 9052 50534 9092
rect 50574 9052 50616 9092
rect 50656 9052 50665 9092
rect 3679 8296 3688 8336
rect 3728 8296 3770 8336
rect 3810 8296 3852 8336
rect 3892 8296 3934 8336
rect 3974 8296 4016 8336
rect 4056 8296 4065 8336
rect 18799 8296 18808 8336
rect 18848 8296 18890 8336
rect 18930 8296 18972 8336
rect 19012 8296 19054 8336
rect 19094 8296 19136 8336
rect 19176 8296 19185 8336
rect 33919 8296 33928 8336
rect 33968 8296 34010 8336
rect 34050 8296 34092 8336
rect 34132 8296 34174 8336
rect 34214 8296 34256 8336
rect 34296 8296 34305 8336
rect 49039 8296 49048 8336
rect 49088 8296 49130 8336
rect 49170 8296 49212 8336
rect 49252 8296 49294 8336
rect 49334 8296 49376 8336
rect 49416 8296 49425 8336
rect 4919 7540 4928 7580
rect 4968 7540 5010 7580
rect 5050 7540 5092 7580
rect 5132 7540 5174 7580
rect 5214 7540 5256 7580
rect 5296 7540 5305 7580
rect 20039 7540 20048 7580
rect 20088 7540 20130 7580
rect 20170 7540 20212 7580
rect 20252 7540 20294 7580
rect 20334 7540 20376 7580
rect 20416 7540 20425 7580
rect 35159 7540 35168 7580
rect 35208 7540 35250 7580
rect 35290 7540 35332 7580
rect 35372 7540 35414 7580
rect 35454 7540 35496 7580
rect 35536 7540 35545 7580
rect 50279 7540 50288 7580
rect 50328 7540 50370 7580
rect 50410 7540 50452 7580
rect 50492 7540 50534 7580
rect 50574 7540 50616 7580
rect 50656 7540 50665 7580
rect 3679 6784 3688 6824
rect 3728 6784 3770 6824
rect 3810 6784 3852 6824
rect 3892 6784 3934 6824
rect 3974 6784 4016 6824
rect 4056 6784 4065 6824
rect 18799 6784 18808 6824
rect 18848 6784 18890 6824
rect 18930 6784 18972 6824
rect 19012 6784 19054 6824
rect 19094 6784 19136 6824
rect 19176 6784 19185 6824
rect 33919 6784 33928 6824
rect 33968 6784 34010 6824
rect 34050 6784 34092 6824
rect 34132 6784 34174 6824
rect 34214 6784 34256 6824
rect 34296 6784 34305 6824
rect 49039 6784 49048 6824
rect 49088 6784 49130 6824
rect 49170 6784 49212 6824
rect 49252 6784 49294 6824
rect 49334 6784 49376 6824
rect 49416 6784 49425 6824
rect 4919 6028 4928 6068
rect 4968 6028 5010 6068
rect 5050 6028 5092 6068
rect 5132 6028 5174 6068
rect 5214 6028 5256 6068
rect 5296 6028 5305 6068
rect 20039 6028 20048 6068
rect 20088 6028 20130 6068
rect 20170 6028 20212 6068
rect 20252 6028 20294 6068
rect 20334 6028 20376 6068
rect 20416 6028 20425 6068
rect 35159 6028 35168 6068
rect 35208 6028 35250 6068
rect 35290 6028 35332 6068
rect 35372 6028 35414 6068
rect 35454 6028 35496 6068
rect 35536 6028 35545 6068
rect 50279 6028 50288 6068
rect 50328 6028 50370 6068
rect 50410 6028 50452 6068
rect 50492 6028 50534 6068
rect 50574 6028 50616 6068
rect 50656 6028 50665 6068
rect 3679 5272 3688 5312
rect 3728 5272 3770 5312
rect 3810 5272 3852 5312
rect 3892 5272 3934 5312
rect 3974 5272 4016 5312
rect 4056 5272 4065 5312
rect 18799 5272 18808 5312
rect 18848 5272 18890 5312
rect 18930 5272 18972 5312
rect 19012 5272 19054 5312
rect 19094 5272 19136 5312
rect 19176 5272 19185 5312
rect 33919 5272 33928 5312
rect 33968 5272 34010 5312
rect 34050 5272 34092 5312
rect 34132 5272 34174 5312
rect 34214 5272 34256 5312
rect 34296 5272 34305 5312
rect 49039 5272 49048 5312
rect 49088 5272 49130 5312
rect 49170 5272 49212 5312
rect 49252 5272 49294 5312
rect 49334 5272 49376 5312
rect 49416 5272 49425 5312
rect 4919 4516 4928 4556
rect 4968 4516 5010 4556
rect 5050 4516 5092 4556
rect 5132 4516 5174 4556
rect 5214 4516 5256 4556
rect 5296 4516 5305 4556
rect 20039 4516 20048 4556
rect 20088 4516 20130 4556
rect 20170 4516 20212 4556
rect 20252 4516 20294 4556
rect 20334 4516 20376 4556
rect 20416 4516 20425 4556
rect 35159 4516 35168 4556
rect 35208 4516 35250 4556
rect 35290 4516 35332 4556
rect 35372 4516 35414 4556
rect 35454 4516 35496 4556
rect 35536 4516 35545 4556
rect 50279 4516 50288 4556
rect 50328 4516 50370 4556
rect 50410 4516 50452 4556
rect 50492 4516 50534 4556
rect 50574 4516 50616 4556
rect 50656 4516 50665 4556
rect 22915 4180 22924 4220
rect 22964 4180 23212 4220
rect 23252 4180 23261 4220
rect 8515 4096 8524 4136
rect 8564 4096 28012 4136
rect 28052 4096 28061 4136
rect 22627 4012 22636 4052
rect 22676 4012 23116 4052
rect 23156 4012 23165 4052
rect 16291 3844 16300 3884
rect 16340 3844 23308 3884
rect 23348 3844 23357 3884
rect 31363 3844 31372 3884
rect 31412 3844 38380 3884
rect 38420 3844 38429 3884
rect 3679 3760 3688 3800
rect 3728 3760 3770 3800
rect 3810 3760 3852 3800
rect 3892 3760 3934 3800
rect 3974 3760 4016 3800
rect 4056 3760 4065 3800
rect 18799 3760 18808 3800
rect 18848 3760 18890 3800
rect 18930 3760 18972 3800
rect 19012 3760 19054 3800
rect 19094 3760 19136 3800
rect 19176 3760 19185 3800
rect 22915 3760 22924 3800
rect 22964 3760 28300 3800
rect 28340 3760 28349 3800
rect 33919 3760 33928 3800
rect 33968 3760 34010 3800
rect 34050 3760 34092 3800
rect 34132 3760 34174 3800
rect 34214 3760 34256 3800
rect 34296 3760 34305 3800
rect 49039 3760 49048 3800
rect 49088 3760 49130 3800
rect 49170 3760 49212 3800
rect 49252 3760 49294 3800
rect 49334 3760 49376 3800
rect 49416 3760 49425 3800
rect 20131 3676 20140 3716
rect 20180 3676 28396 3716
rect 28436 3676 28445 3716
rect 30211 3676 30220 3716
rect 30260 3676 33772 3716
rect 33812 3676 33821 3716
rect 20611 3592 20620 3632
rect 20660 3592 23116 3632
rect 23156 3592 23165 3632
rect 13891 3508 13900 3548
rect 13940 3508 17260 3548
rect 17300 3508 17309 3548
rect 22723 3508 22732 3548
rect 22772 3508 23212 3548
rect 23252 3508 23261 3548
rect 21571 3424 21580 3464
rect 21620 3424 29548 3464
rect 29588 3424 29597 3464
rect 31171 3340 31180 3380
rect 31220 3340 35212 3380
rect 35252 3340 35261 3380
rect 33072 3088 33100 3128
rect 33140 3088 33196 3128
rect 33236 3088 33245 3128
rect 4919 3004 4928 3044
rect 4968 3004 5010 3044
rect 5050 3004 5092 3044
rect 5132 3004 5174 3044
rect 5214 3004 5256 3044
rect 5296 3004 5305 3044
rect 20039 3004 20048 3044
rect 20088 3004 20130 3044
rect 20170 3004 20212 3044
rect 20252 3004 20294 3044
rect 20334 3004 20376 3044
rect 20416 3004 20425 3044
rect 35159 3004 35168 3044
rect 35208 3004 35250 3044
rect 35290 3004 35332 3044
rect 35372 3004 35414 3044
rect 35454 3004 35496 3044
rect 35536 3004 35545 3044
rect 50279 3004 50288 3044
rect 50328 3004 50370 3044
rect 50410 3004 50452 3044
rect 50492 3004 50534 3044
rect 50574 3004 50616 3044
rect 50656 3004 50665 3044
rect 8131 2920 8140 2960
rect 8180 2920 25900 2960
rect 25940 2920 25949 2960
rect 14179 2836 14188 2876
rect 14228 2836 15052 2876
rect 15092 2836 15101 2876
rect 16867 2836 16876 2876
rect 16916 2836 40012 2876
rect 40052 2836 40061 2876
rect 1411 2752 1420 2792
rect 1460 2752 35788 2792
rect 35828 2752 35837 2792
rect 18691 2668 18700 2708
rect 18740 2668 19372 2708
rect 19412 2668 19421 2708
rect 20611 2668 20620 2708
rect 20660 2668 21196 2708
rect 21236 2668 21245 2708
rect 21763 2668 21772 2708
rect 21812 2668 26668 2708
rect 26708 2668 26717 2708
rect 28099 2668 28108 2708
rect 28148 2668 40300 2708
rect 40340 2668 40349 2708
rect 7363 2584 7372 2624
rect 7412 2584 28780 2624
rect 28820 2584 28829 2624
rect 12355 2500 12364 2540
rect 12404 2500 34252 2540
rect 34292 2500 34301 2540
rect 1411 2416 1420 2456
rect 1460 2416 41740 2456
rect 41780 2416 41789 2456
rect 15619 2332 15628 2372
rect 15668 2332 19316 2372
rect 20419 2332 20428 2372
rect 20468 2332 21388 2372
rect 21428 2332 21437 2372
rect 21484 2332 41068 2372
rect 41108 2332 41117 2372
rect 19276 2288 19316 2332
rect 21484 2288 21524 2332
rect 3679 2248 3688 2288
rect 3728 2248 3770 2288
rect 3810 2248 3852 2288
rect 3892 2248 3934 2288
rect 3974 2248 4016 2288
rect 4056 2248 4065 2288
rect 18799 2248 18808 2288
rect 18848 2248 18890 2288
rect 18930 2248 18972 2288
rect 19012 2248 19054 2288
rect 19094 2248 19136 2288
rect 19176 2248 19185 2288
rect 19276 2248 21524 2288
rect 22531 2248 22540 2288
rect 22580 2248 24940 2288
rect 24980 2248 24989 2288
rect 33919 2248 33928 2288
rect 33968 2248 34010 2288
rect 34050 2248 34092 2288
rect 34132 2248 34174 2288
rect 34214 2248 34256 2288
rect 34296 2248 34305 2288
rect 49039 2248 49048 2288
rect 49088 2248 49130 2288
rect 49170 2248 49212 2288
rect 49252 2248 49294 2288
rect 49334 2248 49376 2288
rect 49416 2248 49425 2288
rect 15331 2164 15340 2204
rect 15380 2164 41452 2204
rect 41492 2164 41501 2204
rect 15715 2080 15724 2120
rect 15764 2080 41836 2120
rect 41876 2080 41885 2120
rect 14659 1996 14668 2036
rect 14708 1996 42220 2036
rect 42260 1996 42269 2036
rect 12940 1912 19564 1952
rect 19604 1912 19613 1952
rect 19843 1912 19852 1952
rect 19892 1912 42604 1952
rect 42644 1912 42653 1952
rect 12940 1868 12980 1912
rect 3139 1828 3148 1868
rect 3188 1828 12980 1868
rect 19363 1828 19372 1868
rect 19412 1828 28108 1868
rect 28148 1828 28157 1868
rect 33100 1828 35980 1868
rect 36020 1828 36029 1868
rect 1411 1744 1420 1784
rect 1460 1744 30220 1784
rect 30260 1744 30269 1784
rect 13123 1660 13132 1700
rect 13172 1660 31660 1700
rect 31700 1660 31709 1700
rect 33100 1616 33140 1828
rect 7747 1576 7756 1616
rect 7796 1576 20564 1616
rect 20707 1576 20716 1616
rect 20756 1576 33140 1616
rect 20524 1532 20564 1576
rect 4919 1492 4928 1532
rect 4968 1492 5010 1532
rect 5050 1492 5092 1532
rect 5132 1492 5174 1532
rect 5214 1492 5256 1532
rect 5296 1492 5305 1532
rect 14371 1492 14380 1532
rect 14420 1492 19852 1532
rect 19892 1492 19901 1532
rect 20039 1492 20048 1532
rect 20088 1492 20130 1532
rect 20170 1492 20212 1532
rect 20252 1492 20294 1532
rect 20334 1492 20376 1532
rect 20416 1492 20425 1532
rect 20524 1492 25708 1532
rect 25748 1492 25757 1532
rect 35159 1492 35168 1532
rect 35208 1492 35250 1532
rect 35290 1492 35332 1532
rect 35372 1492 35414 1532
rect 35454 1492 35496 1532
rect 35536 1492 35545 1532
rect 50279 1492 50288 1532
rect 50328 1492 50370 1532
rect 50410 1492 50452 1532
rect 50492 1492 50534 1532
rect 50574 1492 50616 1532
rect 50656 1492 50665 1532
rect 1411 1408 1420 1448
rect 1460 1408 30604 1448
rect 30644 1408 30653 1448
rect 1411 1072 1420 1112
rect 1460 1072 28972 1112
rect 29012 1072 29021 1112
rect 4675 484 4684 524
rect 4724 484 22828 524
rect 22868 484 22877 524
rect 5059 400 5068 440
rect 5108 400 23308 440
rect 23348 400 23357 440
rect 10051 316 10060 356
rect 10100 316 18412 356
rect 18452 316 18461 356
rect 21187 316 21196 356
rect 21236 316 39724 356
rect 39764 316 39773 356
rect 11971 232 11980 272
rect 12020 232 34540 272
rect 34580 232 34589 272
rect 19459 148 19468 188
rect 19508 148 45004 188
rect 45044 148 45053 188
rect 14083 64 14092 104
rect 14132 64 44236 104
rect 44276 64 44285 104
rect 50371 64 50380 104
rect 50420 64 50956 104
rect 50996 64 51005 104
<< via4 >>
rect 4928 10564 4968 10604
rect 5010 10564 5050 10604
rect 5092 10564 5132 10604
rect 5174 10564 5214 10604
rect 5256 10564 5296 10604
rect 20048 10564 20088 10604
rect 20130 10564 20170 10604
rect 20212 10564 20252 10604
rect 20294 10564 20334 10604
rect 20376 10564 20416 10604
rect 35168 10564 35208 10604
rect 35250 10564 35290 10604
rect 35332 10564 35372 10604
rect 35414 10564 35454 10604
rect 35496 10564 35536 10604
rect 50288 10564 50328 10604
rect 50370 10564 50410 10604
rect 50452 10564 50492 10604
rect 50534 10564 50574 10604
rect 50616 10564 50656 10604
rect 3688 9808 3728 9848
rect 3770 9808 3810 9848
rect 3852 9808 3892 9848
rect 3934 9808 3974 9848
rect 4016 9808 4056 9848
rect 18808 9808 18848 9848
rect 18890 9808 18930 9848
rect 18972 9808 19012 9848
rect 19054 9808 19094 9848
rect 19136 9808 19176 9848
rect 33928 9808 33968 9848
rect 34010 9808 34050 9848
rect 34092 9808 34132 9848
rect 34174 9808 34214 9848
rect 34256 9808 34296 9848
rect 49048 9808 49088 9848
rect 49130 9808 49170 9848
rect 49212 9808 49252 9848
rect 49294 9808 49334 9848
rect 49376 9808 49416 9848
rect 19468 9472 19508 9512
rect 4928 9052 4968 9092
rect 5010 9052 5050 9092
rect 5092 9052 5132 9092
rect 5174 9052 5214 9092
rect 5256 9052 5296 9092
rect 20048 9052 20088 9092
rect 20130 9052 20170 9092
rect 20212 9052 20252 9092
rect 20294 9052 20334 9092
rect 20376 9052 20416 9092
rect 35168 9052 35208 9092
rect 35250 9052 35290 9092
rect 35332 9052 35372 9092
rect 35414 9052 35454 9092
rect 35496 9052 35536 9092
rect 50288 9052 50328 9092
rect 50370 9052 50410 9092
rect 50452 9052 50492 9092
rect 50534 9052 50574 9092
rect 50616 9052 50656 9092
rect 3688 8296 3728 8336
rect 3770 8296 3810 8336
rect 3852 8296 3892 8336
rect 3934 8296 3974 8336
rect 4016 8296 4056 8336
rect 18808 8296 18848 8336
rect 18890 8296 18930 8336
rect 18972 8296 19012 8336
rect 19054 8296 19094 8336
rect 19136 8296 19176 8336
rect 33928 8296 33968 8336
rect 34010 8296 34050 8336
rect 34092 8296 34132 8336
rect 34174 8296 34214 8336
rect 34256 8296 34296 8336
rect 49048 8296 49088 8336
rect 49130 8296 49170 8336
rect 49212 8296 49252 8336
rect 49294 8296 49334 8336
rect 49376 8296 49416 8336
rect 4928 7540 4968 7580
rect 5010 7540 5050 7580
rect 5092 7540 5132 7580
rect 5174 7540 5214 7580
rect 5256 7540 5296 7580
rect 20048 7540 20088 7580
rect 20130 7540 20170 7580
rect 20212 7540 20252 7580
rect 20294 7540 20334 7580
rect 20376 7540 20416 7580
rect 35168 7540 35208 7580
rect 35250 7540 35290 7580
rect 35332 7540 35372 7580
rect 35414 7540 35454 7580
rect 35496 7540 35536 7580
rect 50288 7540 50328 7580
rect 50370 7540 50410 7580
rect 50452 7540 50492 7580
rect 50534 7540 50574 7580
rect 50616 7540 50656 7580
rect 3688 6784 3728 6824
rect 3770 6784 3810 6824
rect 3852 6784 3892 6824
rect 3934 6784 3974 6824
rect 4016 6784 4056 6824
rect 18808 6784 18848 6824
rect 18890 6784 18930 6824
rect 18972 6784 19012 6824
rect 19054 6784 19094 6824
rect 19136 6784 19176 6824
rect 33928 6784 33968 6824
rect 34010 6784 34050 6824
rect 34092 6784 34132 6824
rect 34174 6784 34214 6824
rect 34256 6784 34296 6824
rect 49048 6784 49088 6824
rect 49130 6784 49170 6824
rect 49212 6784 49252 6824
rect 49294 6784 49334 6824
rect 49376 6784 49416 6824
rect 4928 6028 4968 6068
rect 5010 6028 5050 6068
rect 5092 6028 5132 6068
rect 5174 6028 5214 6068
rect 5256 6028 5296 6068
rect 20048 6028 20088 6068
rect 20130 6028 20170 6068
rect 20212 6028 20252 6068
rect 20294 6028 20334 6068
rect 20376 6028 20416 6068
rect 35168 6028 35208 6068
rect 35250 6028 35290 6068
rect 35332 6028 35372 6068
rect 35414 6028 35454 6068
rect 35496 6028 35536 6068
rect 50288 6028 50328 6068
rect 50370 6028 50410 6068
rect 50452 6028 50492 6068
rect 50534 6028 50574 6068
rect 50616 6028 50656 6068
rect 3688 5272 3728 5312
rect 3770 5272 3810 5312
rect 3852 5272 3892 5312
rect 3934 5272 3974 5312
rect 4016 5272 4056 5312
rect 18808 5272 18848 5312
rect 18890 5272 18930 5312
rect 18972 5272 19012 5312
rect 19054 5272 19094 5312
rect 19136 5272 19176 5312
rect 33928 5272 33968 5312
rect 34010 5272 34050 5312
rect 34092 5272 34132 5312
rect 34174 5272 34214 5312
rect 34256 5272 34296 5312
rect 49048 5272 49088 5312
rect 49130 5272 49170 5312
rect 49212 5272 49252 5312
rect 49294 5272 49334 5312
rect 49376 5272 49416 5312
rect 4928 4516 4968 4556
rect 5010 4516 5050 4556
rect 5092 4516 5132 4556
rect 5174 4516 5214 4556
rect 5256 4516 5296 4556
rect 20048 4516 20088 4556
rect 20130 4516 20170 4556
rect 20212 4516 20252 4556
rect 20294 4516 20334 4556
rect 20376 4516 20416 4556
rect 35168 4516 35208 4556
rect 35250 4516 35290 4556
rect 35332 4516 35372 4556
rect 35414 4516 35454 4556
rect 35496 4516 35536 4556
rect 50288 4516 50328 4556
rect 50370 4516 50410 4556
rect 50452 4516 50492 4556
rect 50534 4516 50574 4556
rect 50616 4516 50656 4556
rect 3688 3760 3728 3800
rect 3770 3760 3810 3800
rect 3852 3760 3892 3800
rect 3934 3760 3974 3800
rect 4016 3760 4056 3800
rect 18808 3760 18848 3800
rect 18890 3760 18930 3800
rect 18972 3760 19012 3800
rect 19054 3760 19094 3800
rect 19136 3760 19176 3800
rect 33928 3760 33968 3800
rect 34010 3760 34050 3800
rect 34092 3760 34132 3800
rect 34174 3760 34214 3800
rect 34256 3760 34296 3800
rect 49048 3760 49088 3800
rect 49130 3760 49170 3800
rect 49212 3760 49252 3800
rect 49294 3760 49334 3800
rect 49376 3760 49416 3800
rect 4928 3004 4968 3044
rect 5010 3004 5050 3044
rect 5092 3004 5132 3044
rect 5174 3004 5214 3044
rect 5256 3004 5296 3044
rect 20048 3004 20088 3044
rect 20130 3004 20170 3044
rect 20212 3004 20252 3044
rect 20294 3004 20334 3044
rect 20376 3004 20416 3044
rect 35168 3004 35208 3044
rect 35250 3004 35290 3044
rect 35332 3004 35372 3044
rect 35414 3004 35454 3044
rect 35496 3004 35536 3044
rect 50288 3004 50328 3044
rect 50370 3004 50410 3044
rect 50452 3004 50492 3044
rect 50534 3004 50574 3044
rect 50616 3004 50656 3044
rect 3688 2248 3728 2288
rect 3770 2248 3810 2288
rect 3852 2248 3892 2288
rect 3934 2248 3974 2288
rect 4016 2248 4056 2288
rect 18808 2248 18848 2288
rect 18890 2248 18930 2288
rect 18972 2248 19012 2288
rect 19054 2248 19094 2288
rect 19136 2248 19176 2288
rect 33928 2248 33968 2288
rect 34010 2248 34050 2288
rect 34092 2248 34132 2288
rect 34174 2248 34214 2288
rect 34256 2248 34296 2288
rect 49048 2248 49088 2288
rect 49130 2248 49170 2288
rect 49212 2248 49252 2288
rect 49294 2248 49334 2288
rect 49376 2248 49416 2288
rect 4928 1492 4968 1532
rect 5010 1492 5050 1532
rect 5092 1492 5132 1532
rect 5174 1492 5214 1532
rect 5256 1492 5296 1532
rect 20048 1492 20088 1532
rect 20130 1492 20170 1532
rect 20212 1492 20252 1532
rect 20294 1492 20334 1532
rect 20376 1492 20416 1532
rect 35168 1492 35208 1532
rect 35250 1492 35290 1532
rect 35332 1492 35372 1532
rect 35414 1492 35454 1532
rect 35496 1492 35536 1532
rect 50288 1492 50328 1532
rect 50370 1492 50410 1532
rect 50452 1492 50492 1532
rect 50534 1492 50574 1532
rect 50616 1492 50656 1532
rect 19468 148 19508 188
<< metal5 >>
rect 3652 9848 4092 12180
rect 3652 9808 3688 9848
rect 3728 9808 3770 9848
rect 3810 9808 3852 9848
rect 3892 9808 3934 9848
rect 3974 9808 4016 9848
rect 4056 9808 4092 9848
rect 3652 8336 4092 9808
rect 3652 8296 3688 8336
rect 3728 8296 3770 8336
rect 3810 8296 3852 8336
rect 3892 8296 3934 8336
rect 3974 8296 4016 8336
rect 4056 8296 4092 8336
rect 3652 6824 4092 8296
rect 3652 6784 3688 6824
rect 3728 6784 3770 6824
rect 3810 6784 3852 6824
rect 3892 6784 3934 6824
rect 3974 6784 4016 6824
rect 4056 6784 4092 6824
rect 3652 5312 4092 6784
rect 3652 5272 3688 5312
rect 3728 5272 3770 5312
rect 3810 5272 3852 5312
rect 3892 5272 3934 5312
rect 3974 5272 4016 5312
rect 4056 5272 4092 5312
rect 3652 3800 4092 5272
rect 3652 3760 3688 3800
rect 3728 3760 3770 3800
rect 3810 3760 3852 3800
rect 3892 3760 3934 3800
rect 3974 3760 4016 3800
rect 4056 3760 4092 3800
rect 3652 2288 4092 3760
rect 3652 2248 3688 2288
rect 3728 2248 3770 2288
rect 3810 2248 3852 2288
rect 3892 2248 3934 2288
rect 3974 2248 4016 2288
rect 4056 2248 4092 2288
rect 3652 0 4092 2248
rect 4892 10604 5332 12180
rect 4892 10564 4928 10604
rect 4968 10564 5010 10604
rect 5050 10564 5092 10604
rect 5132 10564 5174 10604
rect 5214 10564 5256 10604
rect 5296 10564 5332 10604
rect 4892 9092 5332 10564
rect 4892 9052 4928 9092
rect 4968 9052 5010 9092
rect 5050 9052 5092 9092
rect 5132 9052 5174 9092
rect 5214 9052 5256 9092
rect 5296 9052 5332 9092
rect 4892 7580 5332 9052
rect 4892 7540 4928 7580
rect 4968 7540 5010 7580
rect 5050 7540 5092 7580
rect 5132 7540 5174 7580
rect 5214 7540 5256 7580
rect 5296 7540 5332 7580
rect 4892 6068 5332 7540
rect 4892 6028 4928 6068
rect 4968 6028 5010 6068
rect 5050 6028 5092 6068
rect 5132 6028 5174 6068
rect 5214 6028 5256 6068
rect 5296 6028 5332 6068
rect 4892 4556 5332 6028
rect 4892 4516 4928 4556
rect 4968 4516 5010 4556
rect 5050 4516 5092 4556
rect 5132 4516 5174 4556
rect 5214 4516 5256 4556
rect 5296 4516 5332 4556
rect 4892 3044 5332 4516
rect 4892 3004 4928 3044
rect 4968 3004 5010 3044
rect 5050 3004 5092 3044
rect 5132 3004 5174 3044
rect 5214 3004 5256 3044
rect 5296 3004 5332 3044
rect 4892 1532 5332 3004
rect 4892 1492 4928 1532
rect 4968 1492 5010 1532
rect 5050 1492 5092 1532
rect 5132 1492 5174 1532
rect 5214 1492 5256 1532
rect 5296 1492 5332 1532
rect 4892 0 5332 1492
rect 18772 9848 19212 12180
rect 18772 9808 18808 9848
rect 18848 9808 18890 9848
rect 18930 9808 18972 9848
rect 19012 9808 19054 9848
rect 19094 9808 19136 9848
rect 19176 9808 19212 9848
rect 18772 8336 19212 9808
rect 20012 10604 20452 12180
rect 20012 10564 20048 10604
rect 20088 10564 20130 10604
rect 20170 10564 20212 10604
rect 20252 10564 20294 10604
rect 20334 10564 20376 10604
rect 20416 10564 20452 10604
rect 18772 8296 18808 8336
rect 18848 8296 18890 8336
rect 18930 8296 18972 8336
rect 19012 8296 19054 8336
rect 19094 8296 19136 8336
rect 19176 8296 19212 8336
rect 18772 6824 19212 8296
rect 18772 6784 18808 6824
rect 18848 6784 18890 6824
rect 18930 6784 18972 6824
rect 19012 6784 19054 6824
rect 19094 6784 19136 6824
rect 19176 6784 19212 6824
rect 18772 5312 19212 6784
rect 18772 5272 18808 5312
rect 18848 5272 18890 5312
rect 18930 5272 18972 5312
rect 19012 5272 19054 5312
rect 19094 5272 19136 5312
rect 19176 5272 19212 5312
rect 18772 3800 19212 5272
rect 18772 3760 18808 3800
rect 18848 3760 18890 3800
rect 18930 3760 18972 3800
rect 19012 3760 19054 3800
rect 19094 3760 19136 3800
rect 19176 3760 19212 3800
rect 18772 2288 19212 3760
rect 18772 2248 18808 2288
rect 18848 2248 18890 2288
rect 18930 2248 18972 2288
rect 19012 2248 19054 2288
rect 19094 2248 19136 2288
rect 19176 2248 19212 2288
rect 18772 0 19212 2248
rect 19468 9512 19508 9521
rect 19468 188 19508 9472
rect 19468 139 19508 148
rect 20012 9092 20452 10564
rect 20012 9052 20048 9092
rect 20088 9052 20130 9092
rect 20170 9052 20212 9092
rect 20252 9052 20294 9092
rect 20334 9052 20376 9092
rect 20416 9052 20452 9092
rect 20012 7580 20452 9052
rect 20012 7540 20048 7580
rect 20088 7540 20130 7580
rect 20170 7540 20212 7580
rect 20252 7540 20294 7580
rect 20334 7540 20376 7580
rect 20416 7540 20452 7580
rect 20012 6068 20452 7540
rect 20012 6028 20048 6068
rect 20088 6028 20130 6068
rect 20170 6028 20212 6068
rect 20252 6028 20294 6068
rect 20334 6028 20376 6068
rect 20416 6028 20452 6068
rect 20012 4556 20452 6028
rect 20012 4516 20048 4556
rect 20088 4516 20130 4556
rect 20170 4516 20212 4556
rect 20252 4516 20294 4556
rect 20334 4516 20376 4556
rect 20416 4516 20452 4556
rect 20012 3044 20452 4516
rect 20012 3004 20048 3044
rect 20088 3004 20130 3044
rect 20170 3004 20212 3044
rect 20252 3004 20294 3044
rect 20334 3004 20376 3044
rect 20416 3004 20452 3044
rect 20012 1532 20452 3004
rect 20012 1492 20048 1532
rect 20088 1492 20130 1532
rect 20170 1492 20212 1532
rect 20252 1492 20294 1532
rect 20334 1492 20376 1532
rect 20416 1492 20452 1532
rect 20012 0 20452 1492
rect 33892 9848 34332 12180
rect 33892 9808 33928 9848
rect 33968 9808 34010 9848
rect 34050 9808 34092 9848
rect 34132 9808 34174 9848
rect 34214 9808 34256 9848
rect 34296 9808 34332 9848
rect 33892 8336 34332 9808
rect 33892 8296 33928 8336
rect 33968 8296 34010 8336
rect 34050 8296 34092 8336
rect 34132 8296 34174 8336
rect 34214 8296 34256 8336
rect 34296 8296 34332 8336
rect 33892 6824 34332 8296
rect 33892 6784 33928 6824
rect 33968 6784 34010 6824
rect 34050 6784 34092 6824
rect 34132 6784 34174 6824
rect 34214 6784 34256 6824
rect 34296 6784 34332 6824
rect 33892 5312 34332 6784
rect 33892 5272 33928 5312
rect 33968 5272 34010 5312
rect 34050 5272 34092 5312
rect 34132 5272 34174 5312
rect 34214 5272 34256 5312
rect 34296 5272 34332 5312
rect 33892 3800 34332 5272
rect 33892 3760 33928 3800
rect 33968 3760 34010 3800
rect 34050 3760 34092 3800
rect 34132 3760 34174 3800
rect 34214 3760 34256 3800
rect 34296 3760 34332 3800
rect 33892 2288 34332 3760
rect 33892 2248 33928 2288
rect 33968 2248 34010 2288
rect 34050 2248 34092 2288
rect 34132 2248 34174 2288
rect 34214 2248 34256 2288
rect 34296 2248 34332 2288
rect 33892 0 34332 2248
rect 35132 10604 35572 12180
rect 35132 10564 35168 10604
rect 35208 10564 35250 10604
rect 35290 10564 35332 10604
rect 35372 10564 35414 10604
rect 35454 10564 35496 10604
rect 35536 10564 35572 10604
rect 35132 9092 35572 10564
rect 35132 9052 35168 9092
rect 35208 9052 35250 9092
rect 35290 9052 35332 9092
rect 35372 9052 35414 9092
rect 35454 9052 35496 9092
rect 35536 9052 35572 9092
rect 35132 7580 35572 9052
rect 35132 7540 35168 7580
rect 35208 7540 35250 7580
rect 35290 7540 35332 7580
rect 35372 7540 35414 7580
rect 35454 7540 35496 7580
rect 35536 7540 35572 7580
rect 35132 6068 35572 7540
rect 35132 6028 35168 6068
rect 35208 6028 35250 6068
rect 35290 6028 35332 6068
rect 35372 6028 35414 6068
rect 35454 6028 35496 6068
rect 35536 6028 35572 6068
rect 35132 4556 35572 6028
rect 35132 4516 35168 4556
rect 35208 4516 35250 4556
rect 35290 4516 35332 4556
rect 35372 4516 35414 4556
rect 35454 4516 35496 4556
rect 35536 4516 35572 4556
rect 35132 3044 35572 4516
rect 35132 3004 35168 3044
rect 35208 3004 35250 3044
rect 35290 3004 35332 3044
rect 35372 3004 35414 3044
rect 35454 3004 35496 3044
rect 35536 3004 35572 3044
rect 35132 1532 35572 3004
rect 35132 1492 35168 1532
rect 35208 1492 35250 1532
rect 35290 1492 35332 1532
rect 35372 1492 35414 1532
rect 35454 1492 35496 1532
rect 35536 1492 35572 1532
rect 35132 0 35572 1492
rect 49012 9848 49452 12180
rect 49012 9808 49048 9848
rect 49088 9808 49130 9848
rect 49170 9808 49212 9848
rect 49252 9808 49294 9848
rect 49334 9808 49376 9848
rect 49416 9808 49452 9848
rect 49012 8336 49452 9808
rect 49012 8296 49048 8336
rect 49088 8296 49130 8336
rect 49170 8296 49212 8336
rect 49252 8296 49294 8336
rect 49334 8296 49376 8336
rect 49416 8296 49452 8336
rect 49012 6824 49452 8296
rect 49012 6784 49048 6824
rect 49088 6784 49130 6824
rect 49170 6784 49212 6824
rect 49252 6784 49294 6824
rect 49334 6784 49376 6824
rect 49416 6784 49452 6824
rect 49012 5312 49452 6784
rect 49012 5272 49048 5312
rect 49088 5272 49130 5312
rect 49170 5272 49212 5312
rect 49252 5272 49294 5312
rect 49334 5272 49376 5312
rect 49416 5272 49452 5312
rect 49012 3800 49452 5272
rect 49012 3760 49048 3800
rect 49088 3760 49130 3800
rect 49170 3760 49212 3800
rect 49252 3760 49294 3800
rect 49334 3760 49376 3800
rect 49416 3760 49452 3800
rect 49012 2288 49452 3760
rect 49012 2248 49048 2288
rect 49088 2248 49130 2288
rect 49170 2248 49212 2288
rect 49252 2248 49294 2288
rect 49334 2248 49376 2288
rect 49416 2248 49452 2288
rect 49012 0 49452 2248
rect 50252 10604 50692 12180
rect 50252 10564 50288 10604
rect 50328 10564 50370 10604
rect 50410 10564 50452 10604
rect 50492 10564 50534 10604
rect 50574 10564 50616 10604
rect 50656 10564 50692 10604
rect 50252 9092 50692 10564
rect 50252 9052 50288 9092
rect 50328 9052 50370 9092
rect 50410 9052 50452 9092
rect 50492 9052 50534 9092
rect 50574 9052 50616 9092
rect 50656 9052 50692 9092
rect 50252 7580 50692 9052
rect 50252 7540 50288 7580
rect 50328 7540 50370 7580
rect 50410 7540 50452 7580
rect 50492 7540 50534 7580
rect 50574 7540 50616 7580
rect 50656 7540 50692 7580
rect 50252 6068 50692 7540
rect 50252 6028 50288 6068
rect 50328 6028 50370 6068
rect 50410 6028 50452 6068
rect 50492 6028 50534 6068
rect 50574 6028 50616 6068
rect 50656 6028 50692 6068
rect 50252 4556 50692 6028
rect 50252 4516 50288 4556
rect 50328 4516 50370 4556
rect 50410 4516 50452 4556
rect 50492 4516 50534 4556
rect 50574 4516 50616 4556
rect 50656 4516 50692 4556
rect 50252 3044 50692 4516
rect 50252 3004 50288 3044
rect 50328 3004 50370 3044
rect 50410 3004 50452 3044
rect 50492 3004 50534 3044
rect 50574 3004 50616 3044
rect 50656 3004 50692 3044
rect 50252 1532 50692 3004
rect 50252 1492 50288 1532
rect 50328 1492 50370 1532
rect 50410 1492 50452 1532
rect 50492 1492 50534 1532
rect 50574 1492 50616 1532
rect 50656 1492 50692 1532
rect 50252 0 50692 1492
use sg13g2_buf_1  _000_
timestamp 1676381911
transform 1 0 2112 0 -1 3024
box -48 -56 432 834
use sg13g2_buf_1  _001_
timestamp 1676381911
transform 1 0 29568 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  _002_
timestamp 1676381911
transform 1 0 30720 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  _003_
timestamp 1676381911
transform 1 0 30336 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  _004_
timestamp 1676381911
transform 1 0 7200 0 -1 3024
box -48 -56 432 834
use sg13g2_buf_1  _005_
timestamp 1676381911
transform 1 0 41952 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  _006_
timestamp 1676381911
transform 1 0 35712 0 1 6048
box -48 -56 432 834
use sg13g2_buf_1  _007_
timestamp 1676381911
transform 1 0 33408 0 -1 9072
box -48 -56 432 834
use sg13g2_buf_1  _008_
timestamp 1676381911
transform 1 0 38208 0 1 6048
box -48 -56 432 834
use sg13g2_buf_1  _009_
timestamp 1676381911
transform 1 0 26112 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  _010_
timestamp 1676381911
transform 1 0 35136 0 1 7560
box -48 -56 432 834
use sg13g2_buf_1  _011_
timestamp 1676381911
transform 1 0 31392 0 1 7560
box -48 -56 432 834
use sg13g2_buf_1  _012_
timestamp 1676381911
transform 1 0 29664 0 -1 7560
box -48 -56 432 834
use sg13g2_buf_1  _013_
timestamp 1676381911
transform 1 0 27648 0 -1 9072
box -48 -56 432 834
use sg13g2_buf_1  _014_
timestamp 1676381911
transform 1 0 18816 0 -1 7560
box -48 -56 432 834
use sg13g2_buf_1  _015_
timestamp 1676381911
transform 1 0 22656 0 1 6048
box -48 -56 432 834
use sg13g2_buf_1  _016_
timestamp 1676381911
transform 1 0 25728 0 1 6048
box -48 -56 432 834
use sg13g2_buf_1  _017_
timestamp 1676381911
transform 1 0 29952 0 1 4536
box -48 -56 432 834
use sg13g2_buf_1  _018_
timestamp 1676381911
transform 1 0 23808 0 -1 6048
box -48 -56 432 834
use sg13g2_buf_1  _019_
timestamp 1676381911
transform 1 0 27744 0 -1 6048
box -48 -56 432 834
use sg13g2_buf_1  _020_
timestamp 1676381911
transform 1 0 25344 0 1 6048
box -48 -56 432 834
use sg13g2_buf_1  _021_
timestamp 1676381911
transform 1 0 23520 0 -1 7560
box -48 -56 432 834
use sg13g2_buf_1  _022_
timestamp 1676381911
transform 1 0 30144 0 -1 7560
box -48 -56 432 834
use sg13g2_buf_1  _023_
timestamp 1676381911
transform 1 0 23232 0 1 7560
box -48 -56 432 834
use sg13g2_buf_1  _024_
timestamp 1676381911
transform 1 0 27936 0 1 7560
box -48 -56 432 834
use sg13g2_buf_1  _025_
timestamp 1676381911
transform 1 0 28032 0 -1 9072
box -48 -56 432 834
use sg13g2_buf_1  _026_
timestamp 1676381911
transform 1 0 30144 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  _027_
timestamp 1676381911
transform 1 0 25536 0 -1 9072
box -48 -56 432 834
use sg13g2_buf_1  _028_
timestamp 1676381911
transform 1 0 26592 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  _029_
timestamp 1676381911
transform 1 0 14208 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  _030_
timestamp 1676381911
transform 1 0 23712 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  _031_
timestamp 1676381911
transform 1 0 28800 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  _032_
timestamp 1676381911
transform -1 0 40992 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  _033_
timestamp 1676381911
transform -1 0 41952 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  _034_
timestamp 1676381911
transform -1 0 42912 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  _035_
timestamp 1676381911
transform -1 0 14208 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  _036_
timestamp 1676381911
transform -1 0 16128 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  _037_
timestamp 1676381911
transform -1 0 18816 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  _038_
timestamp 1676381911
transform -1 0 21216 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  _039_
timestamp 1676381911
transform -1 0 23520 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  _040_
timestamp 1676381911
transform -1 0 25728 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  _041_
timestamp 1676381911
transform -1 0 28224 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  _042_
timestamp 1676381911
transform -1 0 30048 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  _043_
timestamp 1676381911
transform -1 0 44352 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  _044_
timestamp 1676381911
transform -1 0 45312 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  _045_
timestamp 1676381911
transform -1 0 46560 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  _046_
timestamp 1676381911
transform -1 0 47424 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  _047_
timestamp 1676381911
transform -1 0 43776 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  _048_
timestamp 1676381911
transform -1 0 47040 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  _049_
timestamp 1676381911
transform -1 0 48576 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  _050_
timestamp 1676381911
transform 1 0 48576 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  _051_
timestamp 1676381911
transform 1 0 50880 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  _052_
timestamp 1676381911
transform 1 0 17088 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  _053_
timestamp 1676381911
transform 1 0 18144 0 -1 3024
box -48 -56 432 834
use sg13g2_buf_1  _054_
timestamp 1676381911
transform 1 0 19488 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  _055_
timestamp 1676381911
transform 1 0 20448 0 -1 3024
box -48 -56 432 834
use sg13g2_buf_1  _056_
timestamp 1676381911
transform 1 0 21600 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  _057_
timestamp 1676381911
transform 1 0 22944 0 -1 4536
box -48 -56 432 834
use sg13g2_buf_1  _058_
timestamp 1676381911
transform 1 0 24096 0 1 4536
box -48 -56 432 834
use sg13g2_buf_1  _059_
timestamp 1676381911
transform 1 0 25152 0 1 4536
box -48 -56 432 834
use sg13g2_buf_1  _060_
timestamp 1676381911
transform 1 0 24768 0 1 4536
box -48 -56 432 834
use sg13g2_buf_1  _061_
timestamp 1676381911
transform 1 0 23424 0 -1 3024
box -48 -56 432 834
use sg13g2_buf_1  _062_
timestamp 1676381911
transform 1 0 22944 0 -1 3024
box -48 -56 432 834
use sg13g2_buf_1  _063_
timestamp 1676381911
transform 1 0 24000 0 -1 3024
box -48 -56 432 834
use sg13g2_buf_1  _064_
timestamp 1676381911
transform 1 0 24864 0 -1 3024
box -48 -56 432 834
use sg13g2_buf_1  _065_
timestamp 1676381911
transform 1 0 24480 0 -1 3024
box -48 -56 432 834
use sg13g2_buf_1  _066_
timestamp 1676381911
transform 1 0 25536 0 -1 3024
box -48 -56 432 834
use sg13g2_buf_1  _067_
timestamp 1676381911
transform 1 0 26976 0 -1 3024
box -48 -56 432 834
use sg13g2_buf_1  _068_
timestamp 1676381911
transform 1 0 27936 0 -1 4536
box -48 -56 432 834
use sg13g2_buf_1  _069_
timestamp 1676381911
transform 1 0 28128 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  _070_
timestamp 1676381911
transform 1 0 28320 0 -1 3024
box -48 -56 432 834
use sg13g2_buf_1  _071_
timestamp 1676381911
transform 1 0 28704 0 -1 3024
box -48 -56 432 834
use sg13g2_buf_1  _072_
timestamp 1676381911
transform 1 0 14016 0 -1 3024
box -48 -56 432 834
use sg13g2_buf_1  _073_
timestamp 1676381911
transform 1 0 14592 0 -1 3024
box -48 -56 432 834
use sg13g2_buf_1  _074_
timestamp 1676381911
transform 1 0 13056 0 -1 3024
box -48 -56 432 834
use sg13g2_buf_1  _075_
timestamp 1676381911
transform 1 0 11712 0 -1 3024
box -48 -56 432 834
use sg13g2_buf_1  _076_
timestamp 1676381911
transform 1 0 31104 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  _077_
timestamp 1676381911
transform 1 0 31584 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  _078_
timestamp 1676381911
transform 1 0 32352 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  _079_
timestamp 1676381911
transform 1 0 32832 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  _080_
timestamp 1676381911
transform 1 0 33312 0 -1 3024
box -48 -56 432 834
use sg13g2_buf_1  _081_
timestamp 1676381911
transform 1 0 33696 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  _082_
timestamp 1676381911
transform 1 0 34176 0 -1 3024
box -48 -56 432 834
use sg13g2_buf_1  _083_
timestamp 1676381911
transform 1 0 34560 0 -1 3024
box -48 -56 432 834
use sg13g2_buf_1  _084_
timestamp 1676381911
transform 1 0 34944 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  _085_
timestamp 1676381911
transform -1 0 35904 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  _086_
timestamp 1676381911
transform -1 0 36384 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  _087_
timestamp 1676381911
transform -1 0 37056 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  _088_
timestamp 1676381911
transform -1 0 37824 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  _089_
timestamp 1676381911
transform -1 0 38976 0 -1 4536
box -48 -56 432 834
use sg13g2_buf_1  _090_
timestamp 1676381911
transform -1 0 39648 0 -1 3024
box -48 -56 432 834
use sg13g2_buf_1  _091_
timestamp 1676381911
transform -1 0 40128 0 -1 3024
box -48 -56 432 834
use sg13g2_buf_1  _092_
timestamp 1676381911
transform 1 0 22464 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  _093_
timestamp 1676381911
transform 1 0 21216 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  _094_
timestamp 1676381911
transform 1 0 20832 0 -1 3024
box -48 -56 432 834
use sg13g2_buf_1  _095_
timestamp 1676381911
transform 1 0 19104 0 -1 4536
box -48 -56 432 834
use sg13g2_buf_1  _096_
timestamp 1676381911
transform 1 0 18528 0 -1 3024
box -48 -56 432 834
use sg13g2_buf_1  _097_
timestamp 1676381911
transform 1 0 16800 0 -1 4536
box -48 -56 432 834
use sg13g2_buf_1  _098_
timestamp 1676381911
transform 1 0 16320 0 -1 4536
box -48 -56 432 834
use sg13g2_buf_1  _099_
timestamp 1676381911
transform 1 0 15168 0 1 4536
box -48 -56 432 834
use sg13g2_buf_1  _100_
timestamp 1676381911
transform 1 0 14592 0 1 4536
box -48 -56 432 834
use sg13g2_buf_1  _101_
timestamp 1676381911
transform 1 0 14592 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  _102_
timestamp 1676381911
transform 1 0 14112 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  _103_
timestamp 1676381911
transform 1 0 13344 0 -1 4536
box -48 -56 432 834
use sg13g2_buf_1  _104_
timestamp 1676381911
transform -1 0 40416 0 1 9072
box -48 -56 432 834
use sg13g2_antennanp  ANTENNA_1
timestamp 1679999689
transform 1 0 35424 0 -1 7560
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_2
timestamp 1679999689
transform 1 0 44640 0 1 3024
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_3
timestamp 1679999689
transform 1 0 36000 0 -1 6048
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_4
timestamp 1679999689
transform 1 0 33408 0 1 7560
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_5
timestamp 1679999689
transform 1 0 50688 0 -1 3024
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_6
timestamp 1679999689
transform -1 0 49920 0 1 1512
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_7
timestamp 1679999689
transform -1 0 13824 0 1 9072
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_8
timestamp 1679999689
transform -1 0 15744 0 1 9072
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_9
timestamp 1679999689
transform 1 0 35136 0 -1 7560
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_10
timestamp 1679999689
transform 1 0 44352 0 1 3024
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_11
timestamp 1679999689
transform 1 0 35712 0 -1 6048
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_12
timestamp 1679999689
transform 1 0 35808 0 -1 9072
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_13
timestamp 1679999689
transform 1 0 50400 0 -1 3024
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_14
timestamp 1679999689
transform 1 0 50208 0 1 9072
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_15
timestamp 1679999689
transform 1 0 51072 0 1 3024
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_16
timestamp 1679999689
transform 1 0 44064 0 1 3024
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_17
timestamp 1679999689
transform 1 0 37824 0 1 6048
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_18
timestamp 1679999689
transform -1 0 35808 0 -1 9072
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_19
timestamp 1679999689
transform 1 0 50112 0 -1 3024
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_20
timestamp 1679999689
transform -1 0 50208 0 -1 10584
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_21
timestamp 1679999689
transform -1 0 49632 0 1 1512
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_22
timestamp 1679999689
transform 1 0 43776 0 1 3024
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_23
timestamp 1679999689
transform 1 0 37536 0 1 6048
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_24
timestamp 1679999689
transform -1 0 35520 0 -1 9072
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_25
timestamp 1679999689
transform -1 0 50976 0 1 3024
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_26
timestamp 1679999689
transform 1 0 49824 0 -1 3024
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_27
timestamp 1679999689
transform 1 0 43488 0 1 3024
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_28
timestamp 1679999689
transform 1 0 37248 0 1 6048
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_29
timestamp 1679999689
transform -1 0 35232 0 -1 9072
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_30
timestamp 1679999689
transform -1 0 49344 0 1 1512
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_31
timestamp 1679999689
transform 1 0 49536 0 -1 3024
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_32
timestamp 1679999689
transform 1 0 43200 0 1 3024
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_33
timestamp 1679999689
transform 1 0 36960 0 1 6048
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_34
timestamp 1679999689
transform -1 0 34944 0 -1 9072
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_35
timestamp 1679999689
transform -1 0 49056 0 1 1512
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_36
timestamp 1679999689
transform 1 0 50400 0 1 3024
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_37
timestamp 1679999689
transform 1 0 42912 0 1 3024
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_38
timestamp 1679999689
transform 1 0 36672 0 1 6048
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_39
timestamp 1679999689
transform -1 0 34656 0 -1 9072
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_40
timestamp 1679999689
transform -1 0 50400 0 1 3024
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_41
timestamp 1679999689
transform 1 0 49248 0 -1 3024
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_42
timestamp 1679999689
transform 1 0 42624 0 1 3024
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_43
timestamp 1679999689
transform 1 0 36384 0 1 6048
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_44
timestamp 1679999689
transform -1 0 34368 0 -1 9072
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_45
timestamp 1679999689
transform -1 0 48768 0 1 1512
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_46
timestamp 1679999689
transform -1 0 50976 0 -1 4536
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_47
timestamp 1679999689
transform 1 0 42336 0 1 3024
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_48
timestamp 1679999689
transform 1 0 36096 0 1 6048
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_49
timestamp 1679999689
transform -1 0 34080 0 -1 9072
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_50
timestamp 1679999689
transform -1 0 50112 0 1 3024
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_51
timestamp 1679999689
transform 1 0 48960 0 -1 3024
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_52
timestamp 1679999689
transform 1 0 41664 0 1 3024
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_53
timestamp 1679999689
transform 1 0 35424 0 1 6048
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_54
timestamp 1679999689
transform -1 0 33408 0 -1 9072
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_55
timestamp 1679999689
transform -1 0 50976 0 1 1512
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_56
timestamp 1679999689
transform -1 0 51744 0 1 1512
box -48 -56 336 834
use sg13g2_decap_8  FILLER_0_0
timestamp 1679581782
transform 1 0 1152 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_7
timestamp 1679581782
transform 1 0 1824 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_14
timestamp 1679581782
transform 1 0 2496 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_21
timestamp 1679581782
transform 1 0 3168 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_28
timestamp 1679581782
transform 1 0 3840 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_35
timestamp 1679581782
transform 1 0 4512 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_42
timestamp 1679581782
transform 1 0 5184 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_49
timestamp 1679581782
transform 1 0 5856 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_56
timestamp 1679581782
transform 1 0 6528 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_63
timestamp 1679581782
transform 1 0 7200 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_70
timestamp 1679581782
transform 1 0 7872 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_77
timestamp 1679581782
transform 1 0 8544 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_84
timestamp 1679581782
transform 1 0 9216 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_91
timestamp 1679581782
transform 1 0 9888 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_98
timestamp 1679581782
transform 1 0 10560 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_105
timestamp 1679581782
transform 1 0 11232 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_112
timestamp 1679581782
transform 1 0 11904 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_119
timestamp 1679581782
transform 1 0 12576 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_126
timestamp 1679581782
transform 1 0 13248 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_133
timestamp 1679581782
transform 1 0 13920 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_140
timestamp 1679581782
transform 1 0 14592 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_147
timestamp 1679581782
transform 1 0 15264 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_154
timestamp 1679581782
transform 1 0 15936 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_161
timestamp 1679581782
transform 1 0 16608 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_168
timestamp 1679581782
transform 1 0 17280 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_175
timestamp 1679581782
transform 1 0 17952 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_182
timestamp 1679581782
transform 1 0 18624 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_189
timestamp 1679581782
transform 1 0 19296 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_196
timestamp 1679581782
transform 1 0 19968 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_203
timestamp 1679581782
transform 1 0 20640 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_210
timestamp 1679581782
transform 1 0 21312 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_217
timestamp 1679581782
transform 1 0 21984 0 1 1512
box -48 -56 720 834
use sg13g2_fill_1  FILLER_0_224
timestamp 1677579658
transform 1 0 22656 0 1 1512
box -48 -56 144 834
use sg13g2_decap_8  FILLER_0_433
timestamp 1679581782
transform 1 0 42720 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_440
timestamp 1679581782
transform 1 0 43392 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_447
timestamp 1679581782
transform 1 0 44064 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_454
timestamp 1679581782
transform 1 0 44736 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_461
timestamp 1679581782
transform 1 0 45408 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_468
timestamp 1679581782
transform 1 0 46080 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_475
timestamp 1679581782
transform 1 0 46752 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_482
timestamp 1679581782
transform 1 0 47424 0 1 1512
box -48 -56 720 834
use sg13g2_decap_4  FILLER_0_489
timestamp 1679577901
transform 1 0 48096 0 1 1512
box -48 -56 432 834
use sg13g2_fill_1  FILLER_0_523
timestamp 1677579658
transform 1 0 51360 0 1 1512
box -48 -56 144 834
use sg13g2_decap_8  FILLER_1_0
timestamp 1679581782
transform 1 0 1152 0 -1 3024
box -48 -56 720 834
use sg13g2_fill_2  FILLER_1_7
timestamp 1677580104
transform 1 0 1824 0 -1 3024
box -48 -56 240 834
use sg13g2_fill_1  FILLER_1_9
timestamp 1677579658
transform 1 0 2016 0 -1 3024
box -48 -56 144 834
use sg13g2_decap_8  FILLER_1_14
timestamp 1679581782
transform 1 0 2496 0 -1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_21
timestamp 1679581782
transform 1 0 3168 0 -1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_28
timestamp 1679581782
transform 1 0 3840 0 -1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_35
timestamp 1679581782
transform 1 0 4512 0 -1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_42
timestamp 1679581782
transform 1 0 5184 0 -1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_49
timestamp 1679581782
transform 1 0 5856 0 -1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_56
timestamp 1679581782
transform 1 0 6528 0 -1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_67
timestamp 1679581782
transform 1 0 7584 0 -1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_74
timestamp 1679581782
transform 1 0 8256 0 -1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_81
timestamp 1679581782
transform 1 0 8928 0 -1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_88
timestamp 1679581782
transform 1 0 9600 0 -1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_95
timestamp 1679581782
transform 1 0 10272 0 -1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_102
timestamp 1679581782
transform 1 0 10944 0 -1 3024
box -48 -56 720 834
use sg13g2_fill_1  FILLER_1_109
timestamp 1677579658
transform 1 0 11616 0 -1 3024
box -48 -56 144 834
use sg13g2_decap_8  FILLER_1_114
timestamp 1679581782
transform 1 0 12096 0 -1 3024
box -48 -56 720 834
use sg13g2_fill_2  FILLER_1_121
timestamp 1677580104
transform 1 0 12768 0 -1 3024
box -48 -56 240 834
use sg13g2_fill_1  FILLER_1_123
timestamp 1677579658
transform 1 0 12960 0 -1 3024
box -48 -56 144 834
use sg13g2_decap_4  FILLER_1_128
timestamp 1679577901
transform 1 0 13440 0 -1 3024
box -48 -56 432 834
use sg13g2_fill_2  FILLER_1_132
timestamp 1677580104
transform 1 0 13824 0 -1 3024
box -48 -56 240 834
use sg13g2_fill_2  FILLER_1_138
timestamp 1677580104
transform 1 0 14400 0 -1 3024
box -48 -56 240 834
use sg13g2_decap_8  FILLER_1_144
timestamp 1679581782
transform 1 0 14976 0 -1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_151
timestamp 1679581782
transform 1 0 15648 0 -1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_158
timestamp 1679581782
transform 1 0 16320 0 -1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_165
timestamp 1679581782
transform 1 0 16992 0 -1 3024
box -48 -56 720 834
use sg13g2_decap_4  FILLER_1_172
timestamp 1679577901
transform 1 0 17664 0 -1 3024
box -48 -56 432 834
use sg13g2_fill_1  FILLER_1_176
timestamp 1677579658
transform 1 0 18048 0 -1 3024
box -48 -56 144 834
use sg13g2_decap_8  FILLER_1_185
timestamp 1679581782
transform 1 0 18912 0 -1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_192
timestamp 1679581782
transform 1 0 19584 0 -1 3024
box -48 -56 720 834
use sg13g2_fill_2  FILLER_1_199
timestamp 1677580104
transform 1 0 20256 0 -1 3024
box -48 -56 240 834
use sg13g2_decap_8  FILLER_1_209
timestamp 1679581782
transform 1 0 21216 0 -1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_216
timestamp 1679581782
transform 1 0 21888 0 -1 3024
box -48 -56 720 834
use sg13g2_decap_4  FILLER_1_223
timestamp 1679577901
transform 1 0 22560 0 -1 3024
box -48 -56 432 834
use sg13g2_fill_1  FILLER_1_231
timestamp 1677579658
transform 1 0 23328 0 -1 3024
box -48 -56 144 834
use sg13g2_fill_2  FILLER_1_236
timestamp 1677580104
transform 1 0 23808 0 -1 3024
box -48 -56 240 834
use sg13g2_fill_1  FILLER_1_242
timestamp 1677579658
transform 1 0 24384 0 -1 3024
box -48 -56 144 834
use sg13g2_fill_2  FILLER_1_251
timestamp 1677580104
transform 1 0 25248 0 -1 3024
box -48 -56 240 834
use sg13g2_fill_1  FILLER_1_253
timestamp 1677579658
transform 1 0 25440 0 -1 3024
box -48 -56 144 834
use sg13g2_decap_8  FILLER_1_258
timestamp 1679581782
transform 1 0 25920 0 -1 3024
box -48 -56 720 834
use sg13g2_decap_4  FILLER_1_265
timestamp 1679577901
transform 1 0 26592 0 -1 3024
box -48 -56 432 834
use sg13g2_decap_8  FILLER_1_273
timestamp 1679581782
transform 1 0 27360 0 -1 3024
box -48 -56 720 834
use sg13g2_fill_2  FILLER_1_280
timestamp 1677580104
transform 1 0 28032 0 -1 3024
box -48 -56 240 834
use sg13g2_fill_1  FILLER_1_282
timestamp 1677579658
transform 1 0 28224 0 -1 3024
box -48 -56 144 834
use sg13g2_decap_8  FILLER_1_291
timestamp 1679581782
transform 1 0 29088 0 -1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_298
timestamp 1679581782
transform 1 0 29760 0 -1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_305
timestamp 1679581782
transform 1 0 30432 0 -1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_312
timestamp 1679581782
transform 1 0 31104 0 -1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_319
timestamp 1679581782
transform 1 0 31776 0 -1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_326
timestamp 1679581782
transform 1 0 32448 0 -1 3024
box -48 -56 720 834
use sg13g2_fill_2  FILLER_1_333
timestamp 1677580104
transform 1 0 33120 0 -1 3024
box -48 -56 240 834
use sg13g2_decap_4  FILLER_1_339
timestamp 1679577901
transform 1 0 33696 0 -1 3024
box -48 -56 432 834
use sg13g2_fill_1  FILLER_1_343
timestamp 1677579658
transform 1 0 34080 0 -1 3024
box -48 -56 144 834
use sg13g2_decap_8  FILLER_1_352
timestamp 1679581782
transform 1 0 34944 0 -1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_359
timestamp 1679581782
transform 1 0 35616 0 -1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_366
timestamp 1679581782
transform 1 0 36288 0 -1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_373
timestamp 1679581782
transform 1 0 36960 0 -1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_380
timestamp 1679581782
transform 1 0 37632 0 -1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_387
timestamp 1679581782
transform 1 0 38304 0 -1 3024
box -48 -56 720 834
use sg13g2_fill_2  FILLER_1_394
timestamp 1677580104
transform 1 0 38976 0 -1 3024
box -48 -56 240 834
use sg13g2_fill_1  FILLER_1_396
timestamp 1677579658
transform 1 0 39168 0 -1 3024
box -48 -56 144 834
use sg13g2_fill_1  FILLER_1_401
timestamp 1677579658
transform 1 0 39648 0 -1 3024
box -48 -56 144 834
use sg13g2_decap_8  FILLER_1_406
timestamp 1679581782
transform 1 0 40128 0 -1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_413
timestamp 1679581782
transform 1 0 40800 0 -1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_420
timestamp 1679581782
transform 1 0 41472 0 -1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_427
timestamp 1679581782
transform 1 0 42144 0 -1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_434
timestamp 1679581782
transform 1 0 42816 0 -1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_441
timestamp 1679581782
transform 1 0 43488 0 -1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_448
timestamp 1679581782
transform 1 0 44160 0 -1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_455
timestamp 1679581782
transform 1 0 44832 0 -1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_462
timestamp 1679581782
transform 1 0 45504 0 -1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_469
timestamp 1679581782
transform 1 0 46176 0 -1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_476
timestamp 1679581782
transform 1 0 46848 0 -1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_483
timestamp 1679581782
transform 1 0 47520 0 -1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_490
timestamp 1679581782
transform 1 0 48192 0 -1 3024
box -48 -56 720 834
use sg13g2_fill_1  FILLER_1_497
timestamp 1677579658
transform 1 0 48864 0 -1 3024
box -48 -56 144 834
use sg13g2_decap_8  FILLER_2_0
timestamp 1679581782
transform 1 0 1152 0 1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_7
timestamp 1679581782
transform 1 0 1824 0 1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_14
timestamp 1679581782
transform 1 0 2496 0 1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_21
timestamp 1679581782
transform 1 0 3168 0 1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_28
timestamp 1679581782
transform 1 0 3840 0 1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_35
timestamp 1679581782
transform 1 0 4512 0 1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_42
timestamp 1679581782
transform 1 0 5184 0 1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_49
timestamp 1679581782
transform 1 0 5856 0 1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_56
timestamp 1679581782
transform 1 0 6528 0 1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_63
timestamp 1679581782
transform 1 0 7200 0 1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_70
timestamp 1679581782
transform 1 0 7872 0 1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_77
timestamp 1679581782
transform 1 0 8544 0 1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_84
timestamp 1679581782
transform 1 0 9216 0 1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_91
timestamp 1679581782
transform 1 0 9888 0 1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_98
timestamp 1679581782
transform 1 0 10560 0 1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_105
timestamp 1679581782
transform 1 0 11232 0 1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_112
timestamp 1679581782
transform 1 0 11904 0 1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_119
timestamp 1679581782
transform 1 0 12576 0 1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_126
timestamp 1679581782
transform 1 0 13248 0 1 3024
box -48 -56 720 834
use sg13g2_fill_2  FILLER_2_133
timestamp 1677580104
transform 1 0 13920 0 1 3024
box -48 -56 240 834
use sg13g2_fill_1  FILLER_2_139
timestamp 1677579658
transform 1 0 14496 0 1 3024
box -48 -56 144 834
use sg13g2_decap_8  FILLER_2_144
timestamp 1679581782
transform 1 0 14976 0 1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_151
timestamp 1679581782
transform 1 0 15648 0 1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_158
timestamp 1679581782
transform 1 0 16320 0 1 3024
box -48 -56 720 834
use sg13g2_fill_1  FILLER_2_165
timestamp 1677579658
transform 1 0 16992 0 1 3024
box -48 -56 144 834
use sg13g2_decap_8  FILLER_2_170
timestamp 1679581782
transform 1 0 17472 0 1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_177
timestamp 1679581782
transform 1 0 18144 0 1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_184
timestamp 1679581782
transform 1 0 18816 0 1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_195
timestamp 1679581782
transform 1 0 19872 0 1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_202
timestamp 1679581782
transform 1 0 20544 0 1 3024
box -48 -56 720 834
use sg13g2_decap_4  FILLER_2_217
timestamp 1679577901
transform 1 0 21984 0 1 3024
box -48 -56 432 834
use sg13g2_fill_1  FILLER_2_221
timestamp 1677579658
transform 1 0 22368 0 1 3024
box -48 -56 144 834
use sg13g2_decap_8  FILLER_2_226
timestamp 1679581782
transform 1 0 22848 0 1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_233
timestamp 1679581782
transform 1 0 23520 0 1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_240
timestamp 1679581782
transform 1 0 24192 0 1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_247
timestamp 1679581782
transform 1 0 24864 0 1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_254
timestamp 1679581782
transform 1 0 25536 0 1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_261
timestamp 1679581782
transform 1 0 26208 0 1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_268
timestamp 1679581782
transform 1 0 26880 0 1 3024
box -48 -56 720 834
use sg13g2_decap_4  FILLER_2_275
timestamp 1679577901
transform 1 0 27552 0 1 3024
box -48 -56 432 834
use sg13g2_fill_2  FILLER_2_279
timestamp 1677580104
transform 1 0 27936 0 1 3024
box -48 -56 240 834
use sg13g2_decap_8  FILLER_2_285
timestamp 1679581782
transform 1 0 28512 0 1 3024
box -48 -56 720 834
use sg13g2_decap_4  FILLER_2_292
timestamp 1679577901
transform 1 0 29184 0 1 3024
box -48 -56 432 834
use sg13g2_decap_4  FILLER_2_300
timestamp 1679577901
transform 1 0 29952 0 1 3024
box -48 -56 432 834
use sg13g2_fill_1  FILLER_2_316
timestamp 1677579658
transform 1 0 31488 0 1 3024
box -48 -56 144 834
use sg13g2_decap_4  FILLER_2_321
timestamp 1679577901
transform 1 0 31968 0 1 3024
box -48 -56 432 834
use sg13g2_fill_1  FILLER_2_329
timestamp 1677579658
transform 1 0 32736 0 1 3024
box -48 -56 144 834
use sg13g2_decap_4  FILLER_2_334
timestamp 1679577901
transform 1 0 33216 0 1 3024
box -48 -56 432 834
use sg13g2_fill_1  FILLER_2_338
timestamp 1677579658
transform 1 0 33600 0 1 3024
box -48 -56 144 834
use sg13g2_decap_8  FILLER_2_343
timestamp 1679581782
transform 1 0 34080 0 1 3024
box -48 -56 720 834
use sg13g2_fill_2  FILLER_2_350
timestamp 1677580104
transform 1 0 34752 0 1 3024
box -48 -56 240 834
use sg13g2_fill_2  FILLER_2_356
timestamp 1677580104
transform 1 0 35328 0 1 3024
box -48 -56 240 834
use sg13g2_fill_1  FILLER_2_362
timestamp 1677579658
transform 1 0 35904 0 1 3024
box -48 -56 144 834
use sg13g2_fill_2  FILLER_2_367
timestamp 1677580104
transform 1 0 36384 0 1 3024
box -48 -56 240 834
use sg13g2_fill_1  FILLER_2_369
timestamp 1677579658
transform 1 0 36576 0 1 3024
box -48 -56 144 834
use sg13g2_decap_4  FILLER_2_374
timestamp 1679577901
transform 1 0 37056 0 1 3024
box -48 -56 432 834
use sg13g2_decap_8  FILLER_2_382
timestamp 1679581782
transform 1 0 37824 0 1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_389
timestamp 1679581782
transform 1 0 38496 0 1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_396
timestamp 1679581782
transform 1 0 39168 0 1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_403
timestamp 1679581782
transform 1 0 39840 0 1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_410
timestamp 1679581782
transform 1 0 40512 0 1 3024
box -48 -56 720 834
use sg13g2_decap_4  FILLER_2_417
timestamp 1679577901
transform 1 0 41184 0 1 3024
box -48 -56 432 834
use sg13g2_fill_1  FILLER_2_421
timestamp 1677579658
transform 1 0 41568 0 1 3024
box -48 -56 144 834
use sg13g2_decap_8  FILLER_2_456
timestamp 1679581782
transform 1 0 44928 0 1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_463
timestamp 1679581782
transform 1 0 45600 0 1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_470
timestamp 1679581782
transform 1 0 46272 0 1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_477
timestamp 1679581782
transform 1 0 46944 0 1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_484
timestamp 1679581782
transform 1 0 47616 0 1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_491
timestamp 1679581782
transform 1 0 48288 0 1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_498
timestamp 1679581782
transform 1 0 48960 0 1 3024
box -48 -56 720 834
use sg13g2_fill_2  FILLER_2_505
timestamp 1677580104
transform 1 0 49632 0 1 3024
box -48 -56 240 834
use sg13g2_fill_1  FILLER_2_519
timestamp 1677579658
transform 1 0 50976 0 1 3024
box -48 -56 144 834
use sg13g2_decap_8  FILLER_3_0
timestamp 1679581782
transform 1 0 1152 0 -1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_7
timestamp 1679581782
transform 1 0 1824 0 -1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_14
timestamp 1679581782
transform 1 0 2496 0 -1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_21
timestamp 1679581782
transform 1 0 3168 0 -1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_28
timestamp 1679581782
transform 1 0 3840 0 -1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_35
timestamp 1679581782
transform 1 0 4512 0 -1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_42
timestamp 1679581782
transform 1 0 5184 0 -1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_49
timestamp 1679581782
transform 1 0 5856 0 -1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_56
timestamp 1679581782
transform 1 0 6528 0 -1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_63
timestamp 1679581782
transform 1 0 7200 0 -1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_70
timestamp 1679581782
transform 1 0 7872 0 -1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_77
timestamp 1679581782
transform 1 0 8544 0 -1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_84
timestamp 1679581782
transform 1 0 9216 0 -1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_91
timestamp 1679581782
transform 1 0 9888 0 -1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_98
timestamp 1679581782
transform 1 0 10560 0 -1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_105
timestamp 1679581782
transform 1 0 11232 0 -1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_112
timestamp 1679581782
transform 1 0 11904 0 -1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_119
timestamp 1679581782
transform 1 0 12576 0 -1 4536
box -48 -56 720 834
use sg13g2_fill_1  FILLER_3_126
timestamp 1677579658
transform 1 0 13248 0 -1 4536
box -48 -56 144 834
use sg13g2_decap_8  FILLER_3_131
timestamp 1679581782
transform 1 0 13728 0 -1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_138
timestamp 1679581782
transform 1 0 14400 0 -1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_145
timestamp 1679581782
transform 1 0 15072 0 -1 4536
box -48 -56 720 834
use sg13g2_decap_4  FILLER_3_152
timestamp 1679577901
transform 1 0 15744 0 -1 4536
box -48 -56 432 834
use sg13g2_fill_2  FILLER_3_156
timestamp 1677580104
transform 1 0 16128 0 -1 4536
box -48 -56 240 834
use sg13g2_fill_1  FILLER_3_162
timestamp 1677579658
transform 1 0 16704 0 -1 4536
box -48 -56 144 834
use sg13g2_decap_8  FILLER_3_167
timestamp 1679581782
transform 1 0 17184 0 -1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_174
timestamp 1679581782
transform 1 0 17856 0 -1 4536
box -48 -56 720 834
use sg13g2_decap_4  FILLER_3_181
timestamp 1679577901
transform 1 0 18528 0 -1 4536
box -48 -56 432 834
use sg13g2_fill_2  FILLER_3_185
timestamp 1677580104
transform 1 0 18912 0 -1 4536
box -48 -56 240 834
use sg13g2_decap_8  FILLER_3_191
timestamp 1679581782
transform 1 0 19488 0 -1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_198
timestamp 1679581782
transform 1 0 20160 0 -1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_205
timestamp 1679581782
transform 1 0 20832 0 -1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_212
timestamp 1679581782
transform 1 0 21504 0 -1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_219
timestamp 1679581782
transform 1 0 22176 0 -1 4536
box -48 -56 720 834
use sg13g2_fill_1  FILLER_3_226
timestamp 1677579658
transform 1 0 22848 0 -1 4536
box -48 -56 144 834
use sg13g2_decap_8  FILLER_3_231
timestamp 1679581782
transform 1 0 23328 0 -1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_238
timestamp 1679581782
transform 1 0 24000 0 -1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_245
timestamp 1679581782
transform 1 0 24672 0 -1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_252
timestamp 1679581782
transform 1 0 25344 0 -1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_259
timestamp 1679581782
transform 1 0 26016 0 -1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_266
timestamp 1679581782
transform 1 0 26688 0 -1 4536
box -48 -56 720 834
use sg13g2_decap_4  FILLER_3_273
timestamp 1679577901
transform 1 0 27360 0 -1 4536
box -48 -56 432 834
use sg13g2_fill_2  FILLER_3_277
timestamp 1677580104
transform 1 0 27744 0 -1 4536
box -48 -56 240 834
use sg13g2_decap_8  FILLER_3_283
timestamp 1679581782
transform 1 0 28320 0 -1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_290
timestamp 1679581782
transform 1 0 28992 0 -1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_297
timestamp 1679581782
transform 1 0 29664 0 -1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_304
timestamp 1679581782
transform 1 0 30336 0 -1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_311
timestamp 1679581782
transform 1 0 31008 0 -1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_318
timestamp 1679581782
transform 1 0 31680 0 -1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_325
timestamp 1679581782
transform 1 0 32352 0 -1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_332
timestamp 1679581782
transform 1 0 33024 0 -1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_339
timestamp 1679581782
transform 1 0 33696 0 -1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_346
timestamp 1679581782
transform 1 0 34368 0 -1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_353
timestamp 1679581782
transform 1 0 35040 0 -1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_360
timestamp 1679581782
transform 1 0 35712 0 -1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_367
timestamp 1679581782
transform 1 0 36384 0 -1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_374
timestamp 1679581782
transform 1 0 37056 0 -1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_381
timestamp 1679581782
transform 1 0 37728 0 -1 4536
box -48 -56 720 834
use sg13g2_fill_2  FILLER_3_388
timestamp 1677580104
transform 1 0 38400 0 -1 4536
box -48 -56 240 834
use sg13g2_decap_8  FILLER_3_394
timestamp 1679581782
transform 1 0 38976 0 -1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_401
timestamp 1679581782
transform 1 0 39648 0 -1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_408
timestamp 1679581782
transform 1 0 40320 0 -1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_415
timestamp 1679581782
transform 1 0 40992 0 -1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_422
timestamp 1679581782
transform 1 0 41664 0 -1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_429
timestamp 1679581782
transform 1 0 42336 0 -1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_436
timestamp 1679581782
transform 1 0 43008 0 -1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_443
timestamp 1679581782
transform 1 0 43680 0 -1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_450
timestamp 1679581782
transform 1 0 44352 0 -1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_457
timestamp 1679581782
transform 1 0 45024 0 -1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_464
timestamp 1679581782
transform 1 0 45696 0 -1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_471
timestamp 1679581782
transform 1 0 46368 0 -1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_478
timestamp 1679581782
transform 1 0 47040 0 -1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_485
timestamp 1679581782
transform 1 0 47712 0 -1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_492
timestamp 1679581782
transform 1 0 48384 0 -1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_499
timestamp 1679581782
transform 1 0 49056 0 -1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_506
timestamp 1679581782
transform 1 0 49728 0 -1 4536
box -48 -56 720 834
use sg13g2_fill_2  FILLER_3_513
timestamp 1677580104
transform 1 0 50400 0 -1 4536
box -48 -56 240 834
use sg13g2_fill_1  FILLER_3_515
timestamp 1677579658
transform 1 0 50592 0 -1 4536
box -48 -56 144 834
use sg13g2_decap_8  FILLER_4_0
timestamp 1679581782
transform 1 0 1152 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_7
timestamp 1679581782
transform 1 0 1824 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_14
timestamp 1679581782
transform 1 0 2496 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_21
timestamp 1679581782
transform 1 0 3168 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_28
timestamp 1679581782
transform 1 0 3840 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_35
timestamp 1679581782
transform 1 0 4512 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_42
timestamp 1679581782
transform 1 0 5184 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_49
timestamp 1679581782
transform 1 0 5856 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_56
timestamp 1679581782
transform 1 0 6528 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_63
timestamp 1679581782
transform 1 0 7200 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_70
timestamp 1679581782
transform 1 0 7872 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_77
timestamp 1679581782
transform 1 0 8544 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_84
timestamp 1679581782
transform 1 0 9216 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_91
timestamp 1679581782
transform 1 0 9888 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_98
timestamp 1679581782
transform 1 0 10560 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_105
timestamp 1679581782
transform 1 0 11232 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_112
timestamp 1679581782
transform 1 0 11904 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_119
timestamp 1679581782
transform 1 0 12576 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_126
timestamp 1679581782
transform 1 0 13248 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_133
timestamp 1679581782
transform 1 0 13920 0 1 4536
box -48 -56 720 834
use sg13g2_fill_2  FILLER_4_144
timestamp 1677580104
transform 1 0 14976 0 1 4536
box -48 -56 240 834
use sg13g2_decap_8  FILLER_4_150
timestamp 1679581782
transform 1 0 15552 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_157
timestamp 1679581782
transform 1 0 16224 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_164
timestamp 1679581782
transform 1 0 16896 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_171
timestamp 1679581782
transform 1 0 17568 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_178
timestamp 1679581782
transform 1 0 18240 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_185
timestamp 1679581782
transform 1 0 18912 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_192
timestamp 1679581782
transform 1 0 19584 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_199
timestamp 1679581782
transform 1 0 20256 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_206
timestamp 1679581782
transform 1 0 20928 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_213
timestamp 1679581782
transform 1 0 21600 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_220
timestamp 1679581782
transform 1 0 22272 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_227
timestamp 1679581782
transform 1 0 22944 0 1 4536
box -48 -56 720 834
use sg13g2_decap_4  FILLER_4_234
timestamp 1679577901
transform 1 0 23616 0 1 4536
box -48 -56 432 834
use sg13g2_fill_1  FILLER_4_238
timestamp 1677579658
transform 1 0 24000 0 1 4536
box -48 -56 144 834
use sg13g2_fill_2  FILLER_4_243
timestamp 1677580104
transform 1 0 24480 0 1 4536
box -48 -56 240 834
use sg13g2_fill_1  FILLER_4_245
timestamp 1677579658
transform 1 0 24672 0 1 4536
box -48 -56 144 834
use sg13g2_decap_8  FILLER_4_254
timestamp 1679581782
transform 1 0 25536 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_261
timestamp 1679581782
transform 1 0 26208 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_268
timestamp 1679581782
transform 1 0 26880 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_275
timestamp 1679581782
transform 1 0 27552 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_282
timestamp 1679581782
transform 1 0 28224 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_289
timestamp 1679581782
transform 1 0 28896 0 1 4536
box -48 -56 720 834
use sg13g2_decap_4  FILLER_4_296
timestamp 1679577901
transform 1 0 29568 0 1 4536
box -48 -56 432 834
use sg13g2_decap_8  FILLER_4_304
timestamp 1679581782
transform 1 0 30336 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_311
timestamp 1679581782
transform 1 0 31008 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_318
timestamp 1679581782
transform 1 0 31680 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_325
timestamp 1679581782
transform 1 0 32352 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_332
timestamp 1679581782
transform 1 0 33024 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_339
timestamp 1679581782
transform 1 0 33696 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_346
timestamp 1679581782
transform 1 0 34368 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_353
timestamp 1679581782
transform 1 0 35040 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_360
timestamp 1679581782
transform 1 0 35712 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_367
timestamp 1679581782
transform 1 0 36384 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_374
timestamp 1679581782
transform 1 0 37056 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_381
timestamp 1679581782
transform 1 0 37728 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_388
timestamp 1679581782
transform 1 0 38400 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_395
timestamp 1679581782
transform 1 0 39072 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_402
timestamp 1679581782
transform 1 0 39744 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_409
timestamp 1679581782
transform 1 0 40416 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_416
timestamp 1679581782
transform 1 0 41088 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_423
timestamp 1679581782
transform 1 0 41760 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_430
timestamp 1679581782
transform 1 0 42432 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_437
timestamp 1679581782
transform 1 0 43104 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_444
timestamp 1679581782
transform 1 0 43776 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_451
timestamp 1679581782
transform 1 0 44448 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_458
timestamp 1679581782
transform 1 0 45120 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_465
timestamp 1679581782
transform 1 0 45792 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_472
timestamp 1679581782
transform 1 0 46464 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_479
timestamp 1679581782
transform 1 0 47136 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_486
timestamp 1679581782
transform 1 0 47808 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_493
timestamp 1679581782
transform 1 0 48480 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_500
timestamp 1679581782
transform 1 0 49152 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_507
timestamp 1679581782
transform 1 0 49824 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_514
timestamp 1679581782
transform 1 0 50496 0 1 4536
box -48 -56 720 834
use sg13g2_fill_2  FILLER_4_521
timestamp 1677580104
transform 1 0 51168 0 1 4536
box -48 -56 240 834
use sg13g2_decap_8  FILLER_5_0
timestamp 1679581782
transform 1 0 1152 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_7
timestamp 1679581782
transform 1 0 1824 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_14
timestamp 1679581782
transform 1 0 2496 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_21
timestamp 1679581782
transform 1 0 3168 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_28
timestamp 1679581782
transform 1 0 3840 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_35
timestamp 1679581782
transform 1 0 4512 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_42
timestamp 1679581782
transform 1 0 5184 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_49
timestamp 1679581782
transform 1 0 5856 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_56
timestamp 1679581782
transform 1 0 6528 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_63
timestamp 1679581782
transform 1 0 7200 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_70
timestamp 1679581782
transform 1 0 7872 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_77
timestamp 1679581782
transform 1 0 8544 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_84
timestamp 1679581782
transform 1 0 9216 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_91
timestamp 1679581782
transform 1 0 9888 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_98
timestamp 1679581782
transform 1 0 10560 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_105
timestamp 1679581782
transform 1 0 11232 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_112
timestamp 1679581782
transform 1 0 11904 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_119
timestamp 1679581782
transform 1 0 12576 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_126
timestamp 1679581782
transform 1 0 13248 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_133
timestamp 1679581782
transform 1 0 13920 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_140
timestamp 1679581782
transform 1 0 14592 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_147
timestamp 1679581782
transform 1 0 15264 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_154
timestamp 1679581782
transform 1 0 15936 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_161
timestamp 1679581782
transform 1 0 16608 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_168
timestamp 1679581782
transform 1 0 17280 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_175
timestamp 1679581782
transform 1 0 17952 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_182
timestamp 1679581782
transform 1 0 18624 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_189
timestamp 1679581782
transform 1 0 19296 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_196
timestamp 1679581782
transform 1 0 19968 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_203
timestamp 1679581782
transform 1 0 20640 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_210
timestamp 1679581782
transform 1 0 21312 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_217
timestamp 1679581782
transform 1 0 21984 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_224
timestamp 1679581782
transform 1 0 22656 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_4  FILLER_5_231
timestamp 1679577901
transform 1 0 23328 0 -1 6048
box -48 -56 432 834
use sg13g2_fill_1  FILLER_5_235
timestamp 1677579658
transform 1 0 23712 0 -1 6048
box -48 -56 144 834
use sg13g2_decap_8  FILLER_5_240
timestamp 1679581782
transform 1 0 24192 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_247
timestamp 1679581782
transform 1 0 24864 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_254
timestamp 1679581782
transform 1 0 25536 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_261
timestamp 1679581782
transform 1 0 26208 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_268
timestamp 1679581782
transform 1 0 26880 0 -1 6048
box -48 -56 720 834
use sg13g2_fill_2  FILLER_5_275
timestamp 1677580104
transform 1 0 27552 0 -1 6048
box -48 -56 240 834
use sg13g2_decap_8  FILLER_5_281
timestamp 1679581782
transform 1 0 28128 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_288
timestamp 1679581782
transform 1 0 28800 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_295
timestamp 1679581782
transform 1 0 29472 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_302
timestamp 1679581782
transform 1 0 30144 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_309
timestamp 1679581782
transform 1 0 30816 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_316
timestamp 1679581782
transform 1 0 31488 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_323
timestamp 1679581782
transform 1 0 32160 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_330
timestamp 1679581782
transform 1 0 32832 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_337
timestamp 1679581782
transform 1 0 33504 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_344
timestamp 1679581782
transform 1 0 34176 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_351
timestamp 1679581782
transform 1 0 34848 0 -1 6048
box -48 -56 720 834
use sg13g2_fill_2  FILLER_5_358
timestamp 1677580104
transform 1 0 35520 0 -1 6048
box -48 -56 240 834
use sg13g2_decap_8  FILLER_5_366
timestamp 1679581782
transform 1 0 36288 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_373
timestamp 1679581782
transform 1 0 36960 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_380
timestamp 1679581782
transform 1 0 37632 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_387
timestamp 1679581782
transform 1 0 38304 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_394
timestamp 1679581782
transform 1 0 38976 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_401
timestamp 1679581782
transform 1 0 39648 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_408
timestamp 1679581782
transform 1 0 40320 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_415
timestamp 1679581782
transform 1 0 40992 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_422
timestamp 1679581782
transform 1 0 41664 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_429
timestamp 1679581782
transform 1 0 42336 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_436
timestamp 1679581782
transform 1 0 43008 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_443
timestamp 1679581782
transform 1 0 43680 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_450
timestamp 1679581782
transform 1 0 44352 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_457
timestamp 1679581782
transform 1 0 45024 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_464
timestamp 1679581782
transform 1 0 45696 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_471
timestamp 1679581782
transform 1 0 46368 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_478
timestamp 1679581782
transform 1 0 47040 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_485
timestamp 1679581782
transform 1 0 47712 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_492
timestamp 1679581782
transform 1 0 48384 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_499
timestamp 1679581782
transform 1 0 49056 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_506
timestamp 1679581782
transform 1 0 49728 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_513
timestamp 1679581782
transform 1 0 50400 0 -1 6048
box -48 -56 720 834
use sg13g2_fill_2  FILLER_5_520
timestamp 1677580104
transform 1 0 51072 0 -1 6048
box -48 -56 240 834
use sg13g2_fill_1  FILLER_5_522
timestamp 1677579658
transform 1 0 51264 0 -1 6048
box -48 -56 144 834
use sg13g2_decap_8  FILLER_6_0
timestamp 1679581782
transform 1 0 1152 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_7
timestamp 1679581782
transform 1 0 1824 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_14
timestamp 1679581782
transform 1 0 2496 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_21
timestamp 1679581782
transform 1 0 3168 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_28
timestamp 1679581782
transform 1 0 3840 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_35
timestamp 1679581782
transform 1 0 4512 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_42
timestamp 1679581782
transform 1 0 5184 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_49
timestamp 1679581782
transform 1 0 5856 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_56
timestamp 1679581782
transform 1 0 6528 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_63
timestamp 1679581782
transform 1 0 7200 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_70
timestamp 1679581782
transform 1 0 7872 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_77
timestamp 1679581782
transform 1 0 8544 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_84
timestamp 1679581782
transform 1 0 9216 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_91
timestamp 1679581782
transform 1 0 9888 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_98
timestamp 1679581782
transform 1 0 10560 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_105
timestamp 1679581782
transform 1 0 11232 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_112
timestamp 1679581782
transform 1 0 11904 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_119
timestamp 1679581782
transform 1 0 12576 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_126
timestamp 1679581782
transform 1 0 13248 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_133
timestamp 1679581782
transform 1 0 13920 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_140
timestamp 1679581782
transform 1 0 14592 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_147
timestamp 1679581782
transform 1 0 15264 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_154
timestamp 1679581782
transform 1 0 15936 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_161
timestamp 1679581782
transform 1 0 16608 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_168
timestamp 1679581782
transform 1 0 17280 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_175
timestamp 1679581782
transform 1 0 17952 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_182
timestamp 1679581782
transform 1 0 18624 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_189
timestamp 1679581782
transform 1 0 19296 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_196
timestamp 1679581782
transform 1 0 19968 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_203
timestamp 1679581782
transform 1 0 20640 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_210
timestamp 1679581782
transform 1 0 21312 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_217
timestamp 1679581782
transform 1 0 21984 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_228
timestamp 1679581782
transform 1 0 23040 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_235
timestamp 1679581782
transform 1 0 23712 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_242
timestamp 1679581782
transform 1 0 24384 0 1 6048
box -48 -56 720 834
use sg13g2_fill_2  FILLER_6_249
timestamp 1677580104
transform 1 0 25056 0 1 6048
box -48 -56 240 834
use sg13g2_fill_1  FILLER_6_251
timestamp 1677579658
transform 1 0 25248 0 1 6048
box -48 -56 144 834
use sg13g2_decap_8  FILLER_6_260
timestamp 1679581782
transform 1 0 26112 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_267
timestamp 1679581782
transform 1 0 26784 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_274
timestamp 1679581782
transform 1 0 27456 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_281
timestamp 1679581782
transform 1 0 28128 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_288
timestamp 1679581782
transform 1 0 28800 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_295
timestamp 1679581782
transform 1 0 29472 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_302
timestamp 1679581782
transform 1 0 30144 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_309
timestamp 1679581782
transform 1 0 30816 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_316
timestamp 1679581782
transform 1 0 31488 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_323
timestamp 1679581782
transform 1 0 32160 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_330
timestamp 1679581782
transform 1 0 32832 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_337
timestamp 1679581782
transform 1 0 33504 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_344
timestamp 1679581782
transform 1 0 34176 0 1 6048
box -48 -56 720 834
use sg13g2_decap_4  FILLER_6_351
timestamp 1679577901
transform 1 0 34848 0 1 6048
box -48 -56 432 834
use sg13g2_fill_2  FILLER_6_355
timestamp 1677580104
transform 1 0 35232 0 1 6048
box -48 -56 240 834
use sg13g2_fill_1  FILLER_6_385
timestamp 1677579658
transform 1 0 38112 0 1 6048
box -48 -56 144 834
use sg13g2_decap_8  FILLER_6_390
timestamp 1679581782
transform 1 0 38592 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_397
timestamp 1679581782
transform 1 0 39264 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_404
timestamp 1679581782
transform 1 0 39936 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_411
timestamp 1679581782
transform 1 0 40608 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_418
timestamp 1679581782
transform 1 0 41280 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_425
timestamp 1679581782
transform 1 0 41952 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_432
timestamp 1679581782
transform 1 0 42624 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_439
timestamp 1679581782
transform 1 0 43296 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_446
timestamp 1679581782
transform 1 0 43968 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_453
timestamp 1679581782
transform 1 0 44640 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_460
timestamp 1679581782
transform 1 0 45312 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_467
timestamp 1679581782
transform 1 0 45984 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_474
timestamp 1679581782
transform 1 0 46656 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_481
timestamp 1679581782
transform 1 0 47328 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_488
timestamp 1679581782
transform 1 0 48000 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_495
timestamp 1679581782
transform 1 0 48672 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_502
timestamp 1679581782
transform 1 0 49344 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_509
timestamp 1679581782
transform 1 0 50016 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_516
timestamp 1679581782
transform 1 0 50688 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_0
timestamp 1679581782
transform 1 0 1152 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_7
timestamp 1679581782
transform 1 0 1824 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_14
timestamp 1679581782
transform 1 0 2496 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_21
timestamp 1679581782
transform 1 0 3168 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_28
timestamp 1679581782
transform 1 0 3840 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_35
timestamp 1679581782
transform 1 0 4512 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_42
timestamp 1679581782
transform 1 0 5184 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_49
timestamp 1679581782
transform 1 0 5856 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_56
timestamp 1679581782
transform 1 0 6528 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_63
timestamp 1679581782
transform 1 0 7200 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_70
timestamp 1679581782
transform 1 0 7872 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_77
timestamp 1679581782
transform 1 0 8544 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_84
timestamp 1679581782
transform 1 0 9216 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_91
timestamp 1679581782
transform 1 0 9888 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_98
timestamp 1679581782
transform 1 0 10560 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_105
timestamp 1679581782
transform 1 0 11232 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_112
timestamp 1679581782
transform 1 0 11904 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_119
timestamp 1679581782
transform 1 0 12576 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_126
timestamp 1679581782
transform 1 0 13248 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_133
timestamp 1679581782
transform 1 0 13920 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_140
timestamp 1679581782
transform 1 0 14592 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_147
timestamp 1679581782
transform 1 0 15264 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_154
timestamp 1679581782
transform 1 0 15936 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_161
timestamp 1679581782
transform 1 0 16608 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_168
timestamp 1679581782
transform 1 0 17280 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_175
timestamp 1679581782
transform 1 0 17952 0 -1 7560
box -48 -56 720 834
use sg13g2_fill_2  FILLER_7_182
timestamp 1677580104
transform 1 0 18624 0 -1 7560
box -48 -56 240 834
use sg13g2_decap_8  FILLER_7_188
timestamp 1679581782
transform 1 0 19200 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_195
timestamp 1679581782
transform 1 0 19872 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_202
timestamp 1679581782
transform 1 0 20544 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_209
timestamp 1679581782
transform 1 0 21216 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_216
timestamp 1679581782
transform 1 0 21888 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_223
timestamp 1679581782
transform 1 0 22560 0 -1 7560
box -48 -56 720 834
use sg13g2_fill_2  FILLER_7_230
timestamp 1677580104
transform 1 0 23232 0 -1 7560
box -48 -56 240 834
use sg13g2_fill_1  FILLER_7_232
timestamp 1677579658
transform 1 0 23424 0 -1 7560
box -48 -56 144 834
use sg13g2_decap_8  FILLER_7_237
timestamp 1679581782
transform 1 0 23904 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_244
timestamp 1679581782
transform 1 0 24576 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_251
timestamp 1679581782
transform 1 0 25248 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_258
timestamp 1679581782
transform 1 0 25920 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_265
timestamp 1679581782
transform 1 0 26592 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_272
timestamp 1679581782
transform 1 0 27264 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_279
timestamp 1679581782
transform 1 0 27936 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_286
timestamp 1679581782
transform 1 0 28608 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_4  FILLER_7_293
timestamp 1679577901
transform 1 0 29280 0 -1 7560
box -48 -56 432 834
use sg13g2_fill_1  FILLER_7_301
timestamp 1677579658
transform 1 0 30048 0 -1 7560
box -48 -56 144 834
use sg13g2_decap_8  FILLER_7_306
timestamp 1679581782
transform 1 0 30528 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_313
timestamp 1679581782
transform 1 0 31200 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_320
timestamp 1679581782
transform 1 0 31872 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_327
timestamp 1679581782
transform 1 0 32544 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_334
timestamp 1679581782
transform 1 0 33216 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_341
timestamp 1679581782
transform 1 0 33888 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_4  FILLER_7_348
timestamp 1679577901
transform 1 0 34560 0 -1 7560
box -48 -56 432 834
use sg13g2_fill_2  FILLER_7_352
timestamp 1677580104
transform 1 0 34944 0 -1 7560
box -48 -56 240 834
use sg13g2_decap_8  FILLER_7_360
timestamp 1679581782
transform 1 0 35712 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_367
timestamp 1679581782
transform 1 0 36384 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_374
timestamp 1679581782
transform 1 0 37056 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_381
timestamp 1679581782
transform 1 0 37728 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_388
timestamp 1679581782
transform 1 0 38400 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_395
timestamp 1679581782
transform 1 0 39072 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_402
timestamp 1679581782
transform 1 0 39744 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_409
timestamp 1679581782
transform 1 0 40416 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_416
timestamp 1679581782
transform 1 0 41088 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_423
timestamp 1679581782
transform 1 0 41760 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_430
timestamp 1679581782
transform 1 0 42432 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_437
timestamp 1679581782
transform 1 0 43104 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_444
timestamp 1679581782
transform 1 0 43776 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_451
timestamp 1679581782
transform 1 0 44448 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_458
timestamp 1679581782
transform 1 0 45120 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_465
timestamp 1679581782
transform 1 0 45792 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_472
timestamp 1679581782
transform 1 0 46464 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_479
timestamp 1679581782
transform 1 0 47136 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_486
timestamp 1679581782
transform 1 0 47808 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_493
timestamp 1679581782
transform 1 0 48480 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_500
timestamp 1679581782
transform 1 0 49152 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_507
timestamp 1679581782
transform 1 0 49824 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_514
timestamp 1679581782
transform 1 0 50496 0 -1 7560
box -48 -56 720 834
use sg13g2_fill_2  FILLER_7_521
timestamp 1677580104
transform 1 0 51168 0 -1 7560
box -48 -56 240 834
use sg13g2_decap_8  FILLER_8_0
timestamp 1679581782
transform 1 0 1152 0 1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_7
timestamp 1679581782
transform 1 0 1824 0 1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_14
timestamp 1679581782
transform 1 0 2496 0 1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_21
timestamp 1679581782
transform 1 0 3168 0 1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_28
timestamp 1679581782
transform 1 0 3840 0 1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_35
timestamp 1679581782
transform 1 0 4512 0 1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_42
timestamp 1679581782
transform 1 0 5184 0 1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_49
timestamp 1679581782
transform 1 0 5856 0 1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_56
timestamp 1679581782
transform 1 0 6528 0 1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_63
timestamp 1679581782
transform 1 0 7200 0 1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_70
timestamp 1679581782
transform 1 0 7872 0 1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_77
timestamp 1679581782
transform 1 0 8544 0 1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_84
timestamp 1679581782
transform 1 0 9216 0 1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_91
timestamp 1679581782
transform 1 0 9888 0 1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_98
timestamp 1679581782
transform 1 0 10560 0 1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_105
timestamp 1679581782
transform 1 0 11232 0 1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_112
timestamp 1679581782
transform 1 0 11904 0 1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_119
timestamp 1679581782
transform 1 0 12576 0 1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_126
timestamp 1679581782
transform 1 0 13248 0 1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_133
timestamp 1679581782
transform 1 0 13920 0 1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_140
timestamp 1679581782
transform 1 0 14592 0 1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_147
timestamp 1679581782
transform 1 0 15264 0 1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_154
timestamp 1679581782
transform 1 0 15936 0 1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_161
timestamp 1679581782
transform 1 0 16608 0 1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_168
timestamp 1679581782
transform 1 0 17280 0 1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_175
timestamp 1679581782
transform 1 0 17952 0 1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_182
timestamp 1679581782
transform 1 0 18624 0 1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_189
timestamp 1679581782
transform 1 0 19296 0 1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_196
timestamp 1679581782
transform 1 0 19968 0 1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_203
timestamp 1679581782
transform 1 0 20640 0 1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_210
timestamp 1679581782
transform 1 0 21312 0 1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_217
timestamp 1679581782
transform 1 0 21984 0 1 7560
box -48 -56 720 834
use sg13g2_decap_4  FILLER_8_224
timestamp 1679577901
transform 1 0 22656 0 1 7560
box -48 -56 432 834
use sg13g2_fill_2  FILLER_8_228
timestamp 1677580104
transform 1 0 23040 0 1 7560
box -48 -56 240 834
use sg13g2_decap_8  FILLER_8_234
timestamp 1679581782
transform 1 0 23616 0 1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_241
timestamp 1679581782
transform 1 0 24288 0 1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_248
timestamp 1679581782
transform 1 0 24960 0 1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_255
timestamp 1679581782
transform 1 0 25632 0 1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_262
timestamp 1679581782
transform 1 0 26304 0 1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_269
timestamp 1679581782
transform 1 0 26976 0 1 7560
box -48 -56 720 834
use sg13g2_fill_2  FILLER_8_276
timestamp 1677580104
transform 1 0 27648 0 1 7560
box -48 -56 240 834
use sg13g2_fill_1  FILLER_8_278
timestamp 1677579658
transform 1 0 27840 0 1 7560
box -48 -56 144 834
use sg13g2_decap_8  FILLER_8_283
timestamp 1679581782
transform 1 0 28320 0 1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_290
timestamp 1679581782
transform 1 0 28992 0 1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_297
timestamp 1679581782
transform 1 0 29664 0 1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_304
timestamp 1679581782
transform 1 0 30336 0 1 7560
box -48 -56 720 834
use sg13g2_decap_4  FILLER_8_311
timestamp 1679577901
transform 1 0 31008 0 1 7560
box -48 -56 432 834
use sg13g2_decap_8  FILLER_8_319
timestamp 1679581782
transform 1 0 31776 0 1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_326
timestamp 1679581782
transform 1 0 32448 0 1 7560
box -48 -56 720 834
use sg13g2_fill_2  FILLER_8_333
timestamp 1677580104
transform 1 0 33120 0 1 7560
box -48 -56 240 834
use sg13g2_fill_1  FILLER_8_335
timestamp 1677579658
transform 1 0 33312 0 1 7560
box -48 -56 144 834
use sg13g2_decap_8  FILLER_8_339
timestamp 1679581782
transform 1 0 33696 0 1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_346
timestamp 1679581782
transform 1 0 34368 0 1 7560
box -48 -56 720 834
use sg13g2_fill_1  FILLER_8_353
timestamp 1677579658
transform 1 0 35040 0 1 7560
box -48 -56 144 834
use sg13g2_decap_8  FILLER_8_358
timestamp 1679581782
transform 1 0 35520 0 1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_365
timestamp 1679581782
transform 1 0 36192 0 1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_372
timestamp 1679581782
transform 1 0 36864 0 1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_379
timestamp 1679581782
transform 1 0 37536 0 1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_386
timestamp 1679581782
transform 1 0 38208 0 1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_393
timestamp 1679581782
transform 1 0 38880 0 1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_400
timestamp 1679581782
transform 1 0 39552 0 1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_407
timestamp 1679581782
transform 1 0 40224 0 1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_414
timestamp 1679581782
transform 1 0 40896 0 1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_421
timestamp 1679581782
transform 1 0 41568 0 1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_428
timestamp 1679581782
transform 1 0 42240 0 1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_435
timestamp 1679581782
transform 1 0 42912 0 1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_442
timestamp 1679581782
transform 1 0 43584 0 1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_449
timestamp 1679581782
transform 1 0 44256 0 1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_456
timestamp 1679581782
transform 1 0 44928 0 1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_463
timestamp 1679581782
transform 1 0 45600 0 1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_470
timestamp 1679581782
transform 1 0 46272 0 1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_477
timestamp 1679581782
transform 1 0 46944 0 1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_484
timestamp 1679581782
transform 1 0 47616 0 1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_491
timestamp 1679581782
transform 1 0 48288 0 1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_498
timestamp 1679581782
transform 1 0 48960 0 1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_505
timestamp 1679581782
transform 1 0 49632 0 1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_512
timestamp 1679581782
transform 1 0 50304 0 1 7560
box -48 -56 720 834
use sg13g2_decap_4  FILLER_8_519
timestamp 1679577901
transform 1 0 50976 0 1 7560
box -48 -56 432 834
use sg13g2_decap_8  FILLER_9_0
timestamp 1679581782
transform 1 0 1152 0 -1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_7
timestamp 1679581782
transform 1 0 1824 0 -1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_14
timestamp 1679581782
transform 1 0 2496 0 -1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_21
timestamp 1679581782
transform 1 0 3168 0 -1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_28
timestamp 1679581782
transform 1 0 3840 0 -1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_35
timestamp 1679581782
transform 1 0 4512 0 -1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_42
timestamp 1679581782
transform 1 0 5184 0 -1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_49
timestamp 1679581782
transform 1 0 5856 0 -1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_56
timestamp 1679581782
transform 1 0 6528 0 -1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_63
timestamp 1679581782
transform 1 0 7200 0 -1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_70
timestamp 1679581782
transform 1 0 7872 0 -1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_77
timestamp 1679581782
transform 1 0 8544 0 -1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_84
timestamp 1679581782
transform 1 0 9216 0 -1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_91
timestamp 1679581782
transform 1 0 9888 0 -1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_98
timestamp 1679581782
transform 1 0 10560 0 -1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_105
timestamp 1679581782
transform 1 0 11232 0 -1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_112
timestamp 1679581782
transform 1 0 11904 0 -1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_119
timestamp 1679581782
transform 1 0 12576 0 -1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_126
timestamp 1679581782
transform 1 0 13248 0 -1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_133
timestamp 1679581782
transform 1 0 13920 0 -1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_140
timestamp 1679581782
transform 1 0 14592 0 -1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_147
timestamp 1679581782
transform 1 0 15264 0 -1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_154
timestamp 1679581782
transform 1 0 15936 0 -1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_161
timestamp 1679581782
transform 1 0 16608 0 -1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_168
timestamp 1679581782
transform 1 0 17280 0 -1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_175
timestamp 1679581782
transform 1 0 17952 0 -1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_182
timestamp 1679581782
transform 1 0 18624 0 -1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_189
timestamp 1679581782
transform 1 0 19296 0 -1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_196
timestamp 1679581782
transform 1 0 19968 0 -1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_203
timestamp 1679581782
transform 1 0 20640 0 -1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_210
timestamp 1679581782
transform 1 0 21312 0 -1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_217
timestamp 1679581782
transform 1 0 21984 0 -1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_224
timestamp 1679581782
transform 1 0 22656 0 -1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_231
timestamp 1679581782
transform 1 0 23328 0 -1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_238
timestamp 1679581782
transform 1 0 24000 0 -1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_245
timestamp 1679581782
transform 1 0 24672 0 -1 9072
box -48 -56 720 834
use sg13g2_fill_2  FILLER_9_252
timestamp 1677580104
transform 1 0 25344 0 -1 9072
box -48 -56 240 834
use sg13g2_decap_8  FILLER_9_258
timestamp 1679581782
transform 1 0 25920 0 -1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_265
timestamp 1679581782
transform 1 0 26592 0 -1 9072
box -48 -56 720 834
use sg13g2_decap_4  FILLER_9_272
timestamp 1679577901
transform 1 0 27264 0 -1 9072
box -48 -56 432 834
use sg13g2_decap_8  FILLER_9_284
timestamp 1679581782
transform 1 0 28416 0 -1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_291
timestamp 1679581782
transform 1 0 29088 0 -1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_298
timestamp 1679581782
transform 1 0 29760 0 -1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_305
timestamp 1679581782
transform 1 0 30432 0 -1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_312
timestamp 1679581782
transform 1 0 31104 0 -1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_319
timestamp 1679581782
transform 1 0 31776 0 -1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_326
timestamp 1679581782
transform 1 0 32448 0 -1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_364
timestamp 1679581782
transform 1 0 36096 0 -1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_371
timestamp 1679581782
transform 1 0 36768 0 -1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_378
timestamp 1679581782
transform 1 0 37440 0 -1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_385
timestamp 1679581782
transform 1 0 38112 0 -1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_392
timestamp 1679581782
transform 1 0 38784 0 -1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_399
timestamp 1679581782
transform 1 0 39456 0 -1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_406
timestamp 1679581782
transform 1 0 40128 0 -1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_413
timestamp 1679581782
transform 1 0 40800 0 -1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_420
timestamp 1679581782
transform 1 0 41472 0 -1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_427
timestamp 1679581782
transform 1 0 42144 0 -1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_434
timestamp 1679581782
transform 1 0 42816 0 -1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_441
timestamp 1679581782
transform 1 0 43488 0 -1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_448
timestamp 1679581782
transform 1 0 44160 0 -1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_455
timestamp 1679581782
transform 1 0 44832 0 -1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_462
timestamp 1679581782
transform 1 0 45504 0 -1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_469
timestamp 1679581782
transform 1 0 46176 0 -1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_476
timestamp 1679581782
transform 1 0 46848 0 -1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_483
timestamp 1679581782
transform 1 0 47520 0 -1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_490
timestamp 1679581782
transform 1 0 48192 0 -1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_497
timestamp 1679581782
transform 1 0 48864 0 -1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_504
timestamp 1679581782
transform 1 0 49536 0 -1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_511
timestamp 1679581782
transform 1 0 50208 0 -1 9072
box -48 -56 720 834
use sg13g2_decap_4  FILLER_9_518
timestamp 1679577901
transform 1 0 50880 0 -1 9072
box -48 -56 432 834
use sg13g2_fill_1  FILLER_9_522
timestamp 1677579658
transform 1 0 51264 0 -1 9072
box -48 -56 144 834
use sg13g2_decap_8  FILLER_10_0
timestamp 1679581782
transform 1 0 1152 0 1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_7
timestamp 1679581782
transform 1 0 1824 0 1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_14
timestamp 1679581782
transform 1 0 2496 0 1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_21
timestamp 1679581782
transform 1 0 3168 0 1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_28
timestamp 1679581782
transform 1 0 3840 0 1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_35
timestamp 1679581782
transform 1 0 4512 0 1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_42
timestamp 1679581782
transform 1 0 5184 0 1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_49
timestamp 1679581782
transform 1 0 5856 0 1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_56
timestamp 1679581782
transform 1 0 6528 0 1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_63
timestamp 1679581782
transform 1 0 7200 0 1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_70
timestamp 1679581782
transform 1 0 7872 0 1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_77
timestamp 1679581782
transform 1 0 8544 0 1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_84
timestamp 1679581782
transform 1 0 9216 0 1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_91
timestamp 1679581782
transform 1 0 9888 0 1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_98
timestamp 1679581782
transform 1 0 10560 0 1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_105
timestamp 1679581782
transform 1 0 11232 0 1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_112
timestamp 1679581782
transform 1 0 11904 0 1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_119
timestamp 1679581782
transform 1 0 12576 0 1 9072
box -48 -56 720 834
use sg13g2_fill_2  FILLER_10_126
timestamp 1677580104
transform 1 0 13248 0 1 9072
box -48 -56 240 834
use sg13g2_fill_1  FILLER_10_128
timestamp 1677579658
transform 1 0 13440 0 1 9072
box -48 -56 144 834
use sg13g2_decap_8  FILLER_10_140
timestamp 1679581782
transform 1 0 14592 0 1 9072
box -48 -56 720 834
use sg13g2_fill_2  FILLER_10_147
timestamp 1677580104
transform 1 0 15264 0 1 9072
box -48 -56 240 834
use sg13g2_decap_8  FILLER_10_156
timestamp 1679581782
transform 1 0 16128 0 1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_163
timestamp 1679581782
transform 1 0 16800 0 1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_170
timestamp 1679581782
transform 1 0 17472 0 1 9072
box -48 -56 720 834
use sg13g2_fill_2  FILLER_10_177
timestamp 1677580104
transform 1 0 18144 0 1 9072
box -48 -56 240 834
use sg13g2_fill_1  FILLER_10_179
timestamp 1677579658
transform 1 0 18336 0 1 9072
box -48 -56 144 834
use sg13g2_decap_8  FILLER_10_184
timestamp 1679581782
transform 1 0 18816 0 1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_191
timestamp 1679581782
transform 1 0 19488 0 1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_198
timestamp 1679581782
transform 1 0 20160 0 1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_209
timestamp 1679581782
transform 1 0 21216 0 1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_216
timestamp 1679581782
transform 1 0 21888 0 1 9072
box -48 -56 720 834
use sg13g2_decap_4  FILLER_10_223
timestamp 1679577901
transform 1 0 22560 0 1 9072
box -48 -56 432 834
use sg13g2_fill_2  FILLER_10_227
timestamp 1677580104
transform 1 0 22944 0 1 9072
box -48 -56 240 834
use sg13g2_fill_2  FILLER_10_233
timestamp 1677580104
transform 1 0 23520 0 1 9072
box -48 -56 240 834
use sg13g2_decap_8  FILLER_10_239
timestamp 1679581782
transform 1 0 24096 0 1 9072
box -48 -56 720 834
use sg13g2_decap_4  FILLER_10_246
timestamp 1679577901
transform 1 0 24768 0 1 9072
box -48 -56 432 834
use sg13g2_fill_2  FILLER_10_250
timestamp 1677580104
transform 1 0 25152 0 1 9072
box -48 -56 240 834
use sg13g2_decap_4  FILLER_10_256
timestamp 1679577901
transform 1 0 25728 0 1 9072
box -48 -56 432 834
use sg13g2_fill_1  FILLER_10_264
timestamp 1677579658
transform 1 0 26496 0 1 9072
box -48 -56 144 834
use sg13g2_decap_8  FILLER_10_269
timestamp 1679581782
transform 1 0 26976 0 1 9072
box -48 -56 720 834
use sg13g2_fill_2  FILLER_10_276
timestamp 1677580104
transform 1 0 27648 0 1 9072
box -48 -56 240 834
use sg13g2_decap_4  FILLER_10_282
timestamp 1679577901
transform 1 0 28224 0 1 9072
box -48 -56 432 834
use sg13g2_fill_2  FILLER_10_286
timestamp 1677580104
transform 1 0 28608 0 1 9072
box -48 -56 240 834
use sg13g2_decap_4  FILLER_10_292
timestamp 1679577901
transform 1 0 29184 0 1 9072
box -48 -56 432 834
use sg13g2_fill_1  FILLER_10_296
timestamp 1677579658
transform 1 0 29568 0 1 9072
box -48 -56 144 834
use sg13g2_fill_1  FILLER_10_301
timestamp 1677579658
transform 1 0 30048 0 1 9072
box -48 -56 144 834
use sg13g2_decap_8  FILLER_10_306
timestamp 1679581782
transform 1 0 30528 0 1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_313
timestamp 1679581782
transform 1 0 31200 0 1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_320
timestamp 1679581782
transform 1 0 31872 0 1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_327
timestamp 1679581782
transform 1 0 32544 0 1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_334
timestamp 1679581782
transform 1 0 33216 0 1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_341
timestamp 1679581782
transform 1 0 33888 0 1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_348
timestamp 1679581782
transform 1 0 34560 0 1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_355
timestamp 1679581782
transform 1 0 35232 0 1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_362
timestamp 1679581782
transform 1 0 35904 0 1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_369
timestamp 1679581782
transform 1 0 36576 0 1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_376
timestamp 1679581782
transform 1 0 37248 0 1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_383
timestamp 1679581782
transform 1 0 37920 0 1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_390
timestamp 1679581782
transform 1 0 38592 0 1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_397
timestamp 1679581782
transform 1 0 39264 0 1 9072
box -48 -56 720 834
use sg13g2_fill_1  FILLER_10_404
timestamp 1677579658
transform 1 0 39936 0 1 9072
box -48 -56 144 834
use sg13g2_fill_2  FILLER_10_409
timestamp 1677580104
transform 1 0 40416 0 1 9072
box -48 -56 240 834
use sg13g2_decap_4  FILLER_10_415
timestamp 1679577901
transform 1 0 40992 0 1 9072
box -48 -56 432 834
use sg13g2_fill_2  FILLER_10_419
timestamp 1677580104
transform 1 0 41376 0 1 9072
box -48 -56 240 834
use sg13g2_decap_4  FILLER_10_425
timestamp 1679577901
transform 1 0 41952 0 1 9072
box -48 -56 432 834
use sg13g2_fill_2  FILLER_10_429
timestamp 1677580104
transform 1 0 42336 0 1 9072
box -48 -56 240 834
use sg13g2_decap_4  FILLER_10_435
timestamp 1679577901
transform 1 0 42912 0 1 9072
box -48 -56 432 834
use sg13g2_fill_1  FILLER_10_439
timestamp 1677579658
transform 1 0 43296 0 1 9072
box -48 -56 144 834
use sg13g2_fill_2  FILLER_10_444
timestamp 1677580104
transform 1 0 43776 0 1 9072
box -48 -56 240 834
use sg13g2_decap_4  FILLER_10_450
timestamp 1679577901
transform 1 0 44352 0 1 9072
box -48 -56 432 834
use sg13g2_fill_2  FILLER_10_454
timestamp 1677580104
transform 1 0 44736 0 1 9072
box -48 -56 240 834
use sg13g2_decap_8  FILLER_10_460
timestamp 1679581782
transform 1 0 45312 0 1 9072
box -48 -56 720 834
use sg13g2_fill_2  FILLER_10_467
timestamp 1677580104
transform 1 0 45984 0 1 9072
box -48 -56 240 834
use sg13g2_fill_1  FILLER_10_473
timestamp 1677579658
transform 1 0 46560 0 1 9072
box -48 -56 144 834
use sg13g2_decap_8  FILLER_10_482
timestamp 1679581782
transform 1 0 47424 0 1 9072
box -48 -56 720 834
use sg13g2_fill_1  FILLER_10_489
timestamp 1677579658
transform 1 0 48096 0 1 9072
box -48 -56 144 834
use sg13g2_decap_8  FILLER_10_498
timestamp 1679581782
transform 1 0 48960 0 1 9072
box -48 -56 720 834
use sg13g2_decap_4  FILLER_10_505
timestamp 1679577901
transform 1 0 49632 0 1 9072
box -48 -56 432 834
use sg13g2_fill_2  FILLER_10_509
timestamp 1677580104
transform 1 0 50016 0 1 9072
box -48 -56 240 834
use sg13g2_fill_1  FILLER_10_522
timestamp 1677579658
transform 1 0 51264 0 1 9072
box -48 -56 144 834
use sg13g2_decap_4  FILLER_11_0
timestamp 1679577901
transform 1 0 1152 0 -1 10584
box -48 -56 432 834
use sg13g2_fill_1  FILLER_11_4
timestamp 1677579658
transform 1 0 1536 0 -1 10584
box -48 -56 144 834
use sg13g2_decap_8  FILLER_11_9
timestamp 1679581782
transform 1 0 2016 0 -1 10584
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_16
timestamp 1679581782
transform 1 0 2688 0 -1 10584
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_23
timestamp 1679581782
transform 1 0 3360 0 -1 10584
box -48 -56 720 834
use sg13g2_fill_1  FILLER_11_30
timestamp 1677579658
transform 1 0 4032 0 -1 10584
box -48 -56 144 834
use sg13g2_decap_8  FILLER_11_35
timestamp 1679581782
transform 1 0 4512 0 -1 10584
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_42
timestamp 1679581782
transform 1 0 5184 0 -1 10584
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_49
timestamp 1679581782
transform 1 0 5856 0 -1 10584
box -48 -56 720 834
use sg13g2_fill_1  FILLER_11_56
timestamp 1677579658
transform 1 0 6528 0 -1 10584
box -48 -56 144 834
use sg13g2_decap_8  FILLER_11_61
timestamp 1679581782
transform 1 0 7008 0 -1 10584
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_68
timestamp 1679581782
transform 1 0 7680 0 -1 10584
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_75
timestamp 1679581782
transform 1 0 8352 0 -1 10584
box -48 -56 720 834
use sg13g2_fill_1  FILLER_11_82
timestamp 1677579658
transform 1 0 9024 0 -1 10584
box -48 -56 144 834
use sg13g2_decap_8  FILLER_11_87
timestamp 1679581782
transform 1 0 9504 0 -1 10584
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_94
timestamp 1679581782
transform 1 0 10176 0 -1 10584
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_101
timestamp 1679581782
transform 1 0 10848 0 -1 10584
box -48 -56 720 834
use sg13g2_fill_1  FILLER_11_108
timestamp 1677579658
transform 1 0 11520 0 -1 10584
box -48 -56 144 834
use sg13g2_decap_8  FILLER_11_113
timestamp 1679581782
transform 1 0 12000 0 -1 10584
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_120
timestamp 1679581782
transform 1 0 12672 0 -1 10584
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_127
timestamp 1679581782
transform 1 0 13344 0 -1 10584
box -48 -56 720 834
use sg13g2_fill_1  FILLER_11_134
timestamp 1677579658
transform 1 0 14016 0 -1 10584
box -48 -56 144 834
use sg13g2_decap_8  FILLER_11_139
timestamp 1679581782
transform 1 0 14496 0 -1 10584
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_146
timestamp 1679581782
transform 1 0 15168 0 -1 10584
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_153
timestamp 1679581782
transform 1 0 15840 0 -1 10584
box -48 -56 720 834
use sg13g2_fill_1  FILLER_11_160
timestamp 1677579658
transform 1 0 16512 0 -1 10584
box -48 -56 144 834
use sg13g2_decap_8  FILLER_11_165
timestamp 1679581782
transform 1 0 16992 0 -1 10584
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_172
timestamp 1679581782
transform 1 0 17664 0 -1 10584
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_179
timestamp 1679581782
transform 1 0 18336 0 -1 10584
box -48 -56 720 834
use sg13g2_fill_1  FILLER_11_186
timestamp 1677579658
transform 1 0 19008 0 -1 10584
box -48 -56 144 834
use sg13g2_decap_8  FILLER_11_191
timestamp 1679581782
transform 1 0 19488 0 -1 10584
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_198
timestamp 1679581782
transform 1 0 20160 0 -1 10584
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_205
timestamp 1679581782
transform 1 0 20832 0 -1 10584
box -48 -56 720 834
use sg13g2_fill_1  FILLER_11_212
timestamp 1677579658
transform 1 0 21504 0 -1 10584
box -48 -56 144 834
use sg13g2_decap_8  FILLER_11_217
timestamp 1679581782
transform 1 0 21984 0 -1 10584
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_224
timestamp 1679581782
transform 1 0 22656 0 -1 10584
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_231
timestamp 1679581782
transform 1 0 23328 0 -1 10584
box -48 -56 720 834
use sg13g2_fill_1  FILLER_11_238
timestamp 1677579658
transform 1 0 24000 0 -1 10584
box -48 -56 144 834
use sg13g2_decap_8  FILLER_11_243
timestamp 1679581782
transform 1 0 24480 0 -1 10584
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_250
timestamp 1679581782
transform 1 0 25152 0 -1 10584
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_257
timestamp 1679581782
transform 1 0 25824 0 -1 10584
box -48 -56 720 834
use sg13g2_fill_1  FILLER_11_264
timestamp 1677579658
transform 1 0 26496 0 -1 10584
box -48 -56 144 834
use sg13g2_decap_8  FILLER_11_269
timestamp 1679581782
transform 1 0 26976 0 -1 10584
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_276
timestamp 1679581782
transform 1 0 27648 0 -1 10584
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_283
timestamp 1679581782
transform 1 0 28320 0 -1 10584
box -48 -56 720 834
use sg13g2_fill_1  FILLER_11_290
timestamp 1677579658
transform 1 0 28992 0 -1 10584
box -48 -56 144 834
use sg13g2_decap_8  FILLER_11_295
timestamp 1679581782
transform 1 0 29472 0 -1 10584
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_302
timestamp 1679581782
transform 1 0 30144 0 -1 10584
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_309
timestamp 1679581782
transform 1 0 30816 0 -1 10584
box -48 -56 720 834
use sg13g2_fill_1  FILLER_11_316
timestamp 1677579658
transform 1 0 31488 0 -1 10584
box -48 -56 144 834
use sg13g2_decap_8  FILLER_11_321
timestamp 1679581782
transform 1 0 31968 0 -1 10584
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_328
timestamp 1679581782
transform 1 0 32640 0 -1 10584
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_335
timestamp 1679581782
transform 1 0 33312 0 -1 10584
box -48 -56 720 834
use sg13g2_fill_1  FILLER_11_342
timestamp 1677579658
transform 1 0 33984 0 -1 10584
box -48 -56 144 834
use sg13g2_decap_8  FILLER_11_347
timestamp 1679581782
transform 1 0 34464 0 -1 10584
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_354
timestamp 1679581782
transform 1 0 35136 0 -1 10584
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_361
timestamp 1679581782
transform 1 0 35808 0 -1 10584
box -48 -56 720 834
use sg13g2_fill_1  FILLER_11_368
timestamp 1677579658
transform 1 0 36480 0 -1 10584
box -48 -56 144 834
use sg13g2_decap_8  FILLER_11_373
timestamp 1679581782
transform 1 0 36960 0 -1 10584
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_380
timestamp 1679581782
transform 1 0 37632 0 -1 10584
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_387
timestamp 1679581782
transform 1 0 38304 0 -1 10584
box -48 -56 720 834
use sg13g2_fill_1  FILLER_11_394
timestamp 1677579658
transform 1 0 38976 0 -1 10584
box -48 -56 144 834
use sg13g2_decap_8  FILLER_11_399
timestamp 1679581782
transform 1 0 39456 0 -1 10584
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_406
timestamp 1679581782
transform 1 0 40128 0 -1 10584
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_413
timestamp 1679581782
transform 1 0 40800 0 -1 10584
box -48 -56 720 834
use sg13g2_fill_1  FILLER_11_420
timestamp 1677579658
transform 1 0 41472 0 -1 10584
box -48 -56 144 834
use sg13g2_decap_8  FILLER_11_425
timestamp 1679581782
transform 1 0 41952 0 -1 10584
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_432
timestamp 1679581782
transform 1 0 42624 0 -1 10584
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_439
timestamp 1679581782
transform 1 0 43296 0 -1 10584
box -48 -56 720 834
use sg13g2_fill_1  FILLER_11_446
timestamp 1677579658
transform 1 0 43968 0 -1 10584
box -48 -56 144 834
use sg13g2_decap_8  FILLER_11_451
timestamp 1679581782
transform 1 0 44448 0 -1 10584
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_458
timestamp 1679581782
transform 1 0 45120 0 -1 10584
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_465
timestamp 1679581782
transform 1 0 45792 0 -1 10584
box -48 -56 720 834
use sg13g2_fill_1  FILLER_11_472
timestamp 1677579658
transform 1 0 46464 0 -1 10584
box -48 -56 144 834
use sg13g2_decap_8  FILLER_11_477
timestamp 1679581782
transform 1 0 46944 0 -1 10584
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_484
timestamp 1679581782
transform 1 0 47616 0 -1 10584
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_491
timestamp 1679581782
transform 1 0 48288 0 -1 10584
box -48 -56 720 834
use sg13g2_fill_1  FILLER_11_498
timestamp 1677579658
transform 1 0 48960 0 -1 10584
box -48 -56 144 834
use sg13g2_fill_1  FILLER_11_503
timestamp 1677579658
transform 1 0 49440 0 -1 10584
box -48 -56 144 834
use sg13g2_buf_1  output1
timestamp 1676381911
transform 1 0 50976 0 1 1512
box -48 -56 432 834
use sg13g2_buf_1  output2
timestamp 1676381911
transform 1 0 51360 0 -1 4536
box -48 -56 432 834
use sg13g2_buf_1  output3
timestamp 1676381911
transform 1 0 51744 0 -1 4536
box -48 -56 432 834
use sg13g2_buf_1  output4
timestamp 1676381911
transform 1 0 51360 0 1 4536
box -48 -56 432 834
use sg13g2_buf_1  output5
timestamp 1676381911
transform 1 0 51744 0 1 4536
box -48 -56 432 834
use sg13g2_buf_1  output6
timestamp 1676381911
transform 1 0 51360 0 -1 6048
box -48 -56 432 834
use sg13g2_buf_1  output7
timestamp 1676381911
transform 1 0 51744 0 -1 6048
box -48 -56 432 834
use sg13g2_buf_1  output8
timestamp 1676381911
transform 1 0 51360 0 1 6048
box -48 -56 432 834
use sg13g2_buf_1  output9
timestamp 1676381911
transform 1 0 51744 0 1 6048
box -48 -56 432 834
use sg13g2_buf_1  output10
timestamp 1676381911
transform 1 0 51360 0 -1 7560
box -48 -56 432 834
use sg13g2_buf_1  output11
timestamp 1676381911
transform 1 0 51744 0 -1 7560
box -48 -56 432 834
use sg13g2_buf_1  output12
timestamp 1676381911
transform 1 0 50304 0 1 1512
box -48 -56 432 834
use sg13g2_buf_1  output13
timestamp 1676381911
transform 1 0 51744 0 1 7560
box -48 -56 432 834
use sg13g2_buf_1  output14
timestamp 1676381911
transform 1 0 51360 0 1 7560
box -48 -56 432 834
use sg13g2_buf_1  output15
timestamp 1676381911
transform 1 0 51744 0 -1 9072
box -48 -56 432 834
use sg13g2_buf_1  output16
timestamp 1676381911
transform 1 0 51360 0 -1 9072
box -48 -56 432 834
use sg13g2_buf_1  output17
timestamp 1676381911
transform 1 0 51744 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  output18
timestamp 1676381911
transform 1 0 51360 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  output19
timestamp 1676381911
transform 1 0 49536 0 -1 10584
box -48 -56 432 834
use sg13g2_buf_1  output20
timestamp 1676381911
transform 1 0 51360 0 -1 10584
box -48 -56 432 834
use sg13g2_buf_1  output21
timestamp 1676381911
transform 1 0 50976 0 -1 10584
box -48 -56 432 834
use sg13g2_buf_1  output22
timestamp 1676381911
transform 1 0 50208 0 -1 10584
box -48 -56 432 834
use sg13g2_buf_1  output23
timestamp 1676381911
transform 1 0 50976 0 -1 3024
box -48 -56 432 834
use sg13g2_buf_1  output24
timestamp 1676381911
transform 1 0 50592 0 -1 10584
box -48 -56 432 834
use sg13g2_buf_1  output25
timestamp 1676381911
transform 1 0 50496 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  output26
timestamp 1676381911
transform 1 0 49920 0 1 1512
box -48 -56 432 834
use sg13g2_buf_1  output27
timestamp 1676381911
transform 1 0 51744 0 1 1512
box -48 -56 432 834
use sg13g2_buf_1  output28
timestamp 1676381911
transform 1 0 51360 0 -1 3024
box -48 -56 432 834
use sg13g2_buf_1  output29
timestamp 1676381911
transform 1 0 51744 0 -1 3024
box -48 -56 432 834
use sg13g2_buf_1  output30
timestamp 1676381911
transform 1 0 51360 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  output31
timestamp 1676381911
transform 1 0 50976 0 -1 4536
box -48 -56 432 834
use sg13g2_buf_1  output32
timestamp 1676381911
transform 1 0 51744 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  output33
timestamp 1676381911
transform -1 0 4512 0 -1 10584
box -48 -56 432 834
use sg13g2_buf_1  output34
timestamp 1676381911
transform -1 0 29472 0 -1 10584
box -48 -56 432 834
use sg13g2_buf_1  output35
timestamp 1676381911
transform -1 0 31968 0 -1 10584
box -48 -56 432 834
use sg13g2_buf_1  output36
timestamp 1676381911
transform -1 0 34464 0 -1 10584
box -48 -56 432 834
use sg13g2_buf_1  output37
timestamp 1676381911
transform -1 0 36960 0 -1 10584
box -48 -56 432 834
use sg13g2_buf_1  output38
timestamp 1676381911
transform -1 0 39456 0 -1 10584
box -48 -56 432 834
use sg13g2_buf_1  output39
timestamp 1676381911
transform -1 0 41952 0 -1 10584
box -48 -56 432 834
use sg13g2_buf_1  output40
timestamp 1676381911
transform -1 0 44448 0 -1 10584
box -48 -56 432 834
use sg13g2_buf_1  output41
timestamp 1676381911
transform -1 0 46944 0 -1 10584
box -48 -56 432 834
use sg13g2_buf_1  output42
timestamp 1676381911
transform -1 0 49440 0 -1 10584
box -48 -56 432 834
use sg13g2_buf_1  output43
timestamp 1676381911
transform -1 0 52128 0 -1 10584
box -48 -56 432 834
use sg13g2_buf_1  output44
timestamp 1676381911
transform -1 0 7008 0 -1 10584
box -48 -56 432 834
use sg13g2_buf_1  output45
timestamp 1676381911
transform -1 0 9504 0 -1 10584
box -48 -56 432 834
use sg13g2_buf_1  output46
timestamp 1676381911
transform -1 0 12000 0 -1 10584
box -48 -56 432 834
use sg13g2_buf_1  output47
timestamp 1676381911
transform -1 0 14496 0 -1 10584
box -48 -56 432 834
use sg13g2_buf_1  output48
timestamp 1676381911
transform -1 0 16992 0 -1 10584
box -48 -56 432 834
use sg13g2_buf_1  output49
timestamp 1676381911
transform -1 0 19488 0 -1 10584
box -48 -56 432 834
use sg13g2_buf_1  output50
timestamp 1676381911
transform -1 0 21984 0 -1 10584
box -48 -56 432 834
use sg13g2_buf_1  output51
timestamp 1676381911
transform -1 0 24480 0 -1 10584
box -48 -56 432 834
use sg13g2_buf_1  output52
timestamp 1676381911
transform -1 0 26976 0 -1 10584
box -48 -56 432 834
use sg13g2_buf_1  output53
timestamp 1676381911
transform -1 0 23136 0 1 1512
box -48 -56 432 834
use sg13g2_buf_1  output54
timestamp 1676381911
transform -1 0 23520 0 1 1512
box -48 -56 432 834
use sg13g2_buf_1  output55
timestamp 1676381911
transform -1 0 23904 0 1 1512
box -48 -56 432 834
use sg13g2_buf_1  output56
timestamp 1676381911
transform -1 0 24288 0 1 1512
box -48 -56 432 834
use sg13g2_buf_1  output57
timestamp 1676381911
transform -1 0 24672 0 1 1512
box -48 -56 432 834
use sg13g2_buf_1  output58
timestamp 1676381911
transform -1 0 25056 0 1 1512
box -48 -56 432 834
use sg13g2_buf_1  output59
timestamp 1676381911
transform -1 0 25440 0 1 1512
box -48 -56 432 834
use sg13g2_buf_1  output60
timestamp 1676381911
transform -1 0 25824 0 1 1512
box -48 -56 432 834
use sg13g2_buf_1  output61
timestamp 1676381911
transform -1 0 26208 0 1 1512
box -48 -56 432 834
use sg13g2_buf_1  output62
timestamp 1676381911
transform -1 0 26592 0 1 1512
box -48 -56 432 834
use sg13g2_buf_1  output63
timestamp 1676381911
transform -1 0 26976 0 1 1512
box -48 -56 432 834
use sg13g2_buf_1  output64
timestamp 1676381911
transform -1 0 27360 0 1 1512
box -48 -56 432 834
use sg13g2_buf_1  output65
timestamp 1676381911
transform -1 0 27744 0 1 1512
box -48 -56 432 834
use sg13g2_buf_1  output66
timestamp 1676381911
transform -1 0 28128 0 1 1512
box -48 -56 432 834
use sg13g2_buf_1  output67
timestamp 1676381911
transform -1 0 28512 0 1 1512
box -48 -56 432 834
use sg13g2_buf_1  output68
timestamp 1676381911
transform -1 0 28896 0 1 1512
box -48 -56 432 834
use sg13g2_buf_1  output69
timestamp 1676381911
transform -1 0 29280 0 1 1512
box -48 -56 432 834
use sg13g2_buf_1  output70
timestamp 1676381911
transform -1 0 29664 0 1 1512
box -48 -56 432 834
use sg13g2_buf_1  output71
timestamp 1676381911
transform -1 0 30048 0 1 1512
box -48 -56 432 834
use sg13g2_buf_1  output72
timestamp 1676381911
transform -1 0 30432 0 1 1512
box -48 -56 432 834
use sg13g2_buf_1  output73
timestamp 1676381911
transform -1 0 30816 0 1 1512
box -48 -56 432 834
use sg13g2_buf_1  output74
timestamp 1676381911
transform -1 0 34656 0 1 1512
box -48 -56 432 834
use sg13g2_buf_1  output75
timestamp 1676381911
transform -1 0 35040 0 1 1512
box -48 -56 432 834
use sg13g2_buf_1  output76
timestamp 1676381911
transform -1 0 35424 0 1 1512
box -48 -56 432 834
use sg13g2_buf_1  output77
timestamp 1676381911
transform -1 0 35808 0 1 1512
box -48 -56 432 834
use sg13g2_buf_1  output78
timestamp 1676381911
transform -1 0 36192 0 1 1512
box -48 -56 432 834
use sg13g2_buf_1  output79
timestamp 1676381911
transform -1 0 36576 0 1 1512
box -48 -56 432 834
use sg13g2_buf_1  output80
timestamp 1676381911
transform -1 0 31200 0 1 1512
box -48 -56 432 834
use sg13g2_buf_1  output81
timestamp 1676381911
transform -1 0 31584 0 1 1512
box -48 -56 432 834
use sg13g2_buf_1  output82
timestamp 1676381911
transform -1 0 31968 0 1 1512
box -48 -56 432 834
use sg13g2_buf_1  output83
timestamp 1676381911
transform -1 0 32352 0 1 1512
box -48 -56 432 834
use sg13g2_buf_1  output84
timestamp 1676381911
transform -1 0 32736 0 1 1512
box -48 -56 432 834
use sg13g2_buf_1  output85
timestamp 1676381911
transform -1 0 33120 0 1 1512
box -48 -56 432 834
use sg13g2_buf_1  output86
timestamp 1676381911
transform -1 0 33504 0 1 1512
box -48 -56 432 834
use sg13g2_buf_1  output87
timestamp 1676381911
transform -1 0 33888 0 1 1512
box -48 -56 432 834
use sg13g2_buf_1  output88
timestamp 1676381911
transform -1 0 34272 0 1 1512
box -48 -56 432 834
use sg13g2_buf_1  output89
timestamp 1676381911
transform -1 0 36960 0 1 1512
box -48 -56 432 834
use sg13g2_buf_1  output90
timestamp 1676381911
transform -1 0 40800 0 1 1512
box -48 -56 432 834
use sg13g2_buf_1  output91
timestamp 1676381911
transform -1 0 41184 0 1 1512
box -48 -56 432 834
use sg13g2_buf_1  output92
timestamp 1676381911
transform -1 0 41568 0 1 1512
box -48 -56 432 834
use sg13g2_buf_1  output93
timestamp 1676381911
transform -1 0 41952 0 1 1512
box -48 -56 432 834
use sg13g2_buf_1  output94
timestamp 1676381911
transform -1 0 42336 0 1 1512
box -48 -56 432 834
use sg13g2_buf_1  output95
timestamp 1676381911
transform -1 0 42720 0 1 1512
box -48 -56 432 834
use sg13g2_buf_1  output96
timestamp 1676381911
transform -1 0 37344 0 1 1512
box -48 -56 432 834
use sg13g2_buf_1  output97
timestamp 1676381911
transform -1 0 37728 0 1 1512
box -48 -56 432 834
use sg13g2_buf_1  output98
timestamp 1676381911
transform -1 0 38112 0 1 1512
box -48 -56 432 834
use sg13g2_buf_1  output99
timestamp 1676381911
transform -1 0 38496 0 1 1512
box -48 -56 432 834
use sg13g2_buf_1  output100
timestamp 1676381911
transform -1 0 38880 0 1 1512
box -48 -56 432 834
use sg13g2_buf_1  output101
timestamp 1676381911
transform -1 0 39264 0 1 1512
box -48 -56 432 834
use sg13g2_buf_1  output102
timestamp 1676381911
transform -1 0 39648 0 1 1512
box -48 -56 432 834
use sg13g2_buf_1  output103
timestamp 1676381911
transform -1 0 40032 0 1 1512
box -48 -56 432 834
use sg13g2_buf_1  output104
timestamp 1676381911
transform -1 0 40416 0 1 1512
box -48 -56 432 834
use sg13g2_buf_1  output105
timestamp 1676381911
transform -1 0 2016 0 -1 10584
box -48 -56 432 834
<< labels >>
flabel metal2 s 0 716 90 796 0 FreeSans 320 0 0 0 FrameData[0]
port 0 nsew signal input
flabel metal2 s 0 4076 90 4156 0 FreeSans 320 0 0 0 FrameData[10]
port 1 nsew signal input
flabel metal2 s 0 4412 90 4492 0 FreeSans 320 0 0 0 FrameData[11]
port 2 nsew signal input
flabel metal2 s 0 4748 90 4828 0 FreeSans 320 0 0 0 FrameData[12]
port 3 nsew signal input
flabel metal2 s 0 5084 90 5164 0 FreeSans 320 0 0 0 FrameData[13]
port 4 nsew signal input
flabel metal2 s 0 5420 90 5500 0 FreeSans 320 0 0 0 FrameData[14]
port 5 nsew signal input
flabel metal2 s 0 5756 90 5836 0 FreeSans 320 0 0 0 FrameData[15]
port 6 nsew signal input
flabel metal2 s 0 6092 90 6172 0 FreeSans 320 0 0 0 FrameData[16]
port 7 nsew signal input
flabel metal2 s 0 6428 90 6508 0 FreeSans 320 0 0 0 FrameData[17]
port 8 nsew signal input
flabel metal2 s 0 6764 90 6844 0 FreeSans 320 0 0 0 FrameData[18]
port 9 nsew signal input
flabel metal2 s 0 7100 90 7180 0 FreeSans 320 0 0 0 FrameData[19]
port 10 nsew signal input
flabel metal2 s 0 1052 90 1132 0 FreeSans 320 0 0 0 FrameData[1]
port 11 nsew signal input
flabel metal2 s 0 7436 90 7516 0 FreeSans 320 0 0 0 FrameData[20]
port 12 nsew signal input
flabel metal2 s 0 7772 90 7852 0 FreeSans 320 0 0 0 FrameData[21]
port 13 nsew signal input
flabel metal2 s 0 8108 90 8188 0 FreeSans 320 0 0 0 FrameData[22]
port 14 nsew signal input
flabel metal2 s 0 8444 90 8524 0 FreeSans 320 0 0 0 FrameData[23]
port 15 nsew signal input
flabel metal2 s 0 8780 90 8860 0 FreeSans 320 0 0 0 FrameData[24]
port 16 nsew signal input
flabel metal2 s 0 9116 90 9196 0 FreeSans 320 0 0 0 FrameData[25]
port 17 nsew signal input
flabel metal2 s 0 9452 90 9532 0 FreeSans 320 0 0 0 FrameData[26]
port 18 nsew signal input
flabel metal2 s 0 9788 90 9868 0 FreeSans 320 0 0 0 FrameData[27]
port 19 nsew signal input
flabel metal2 s 0 10124 90 10204 0 FreeSans 320 0 0 0 FrameData[28]
port 20 nsew signal input
flabel metal2 s 0 10460 90 10540 0 FreeSans 320 0 0 0 FrameData[29]
port 21 nsew signal input
flabel metal2 s 0 1388 90 1468 0 FreeSans 320 0 0 0 FrameData[2]
port 22 nsew signal input
flabel metal2 s 0 10796 90 10876 0 FreeSans 320 0 0 0 FrameData[30]
port 23 nsew signal input
flabel metal2 s 0 11132 90 11212 0 FreeSans 320 0 0 0 FrameData[31]
port 24 nsew signal input
flabel metal2 s 0 1724 90 1804 0 FreeSans 320 0 0 0 FrameData[3]
port 25 nsew signal input
flabel metal2 s 0 2060 90 2140 0 FreeSans 320 0 0 0 FrameData[4]
port 26 nsew signal input
flabel metal2 s 0 2396 90 2476 0 FreeSans 320 0 0 0 FrameData[5]
port 27 nsew signal input
flabel metal2 s 0 2732 90 2812 0 FreeSans 320 0 0 0 FrameData[6]
port 28 nsew signal input
flabel metal2 s 0 3068 90 3148 0 FreeSans 320 0 0 0 FrameData[7]
port 29 nsew signal input
flabel metal2 s 0 3404 90 3484 0 FreeSans 320 0 0 0 FrameData[8]
port 30 nsew signal input
flabel metal2 s 0 3740 90 3820 0 FreeSans 320 0 0 0 FrameData[9]
port 31 nsew signal input
flabel metal2 s 53190 716 53280 796 0 FreeSans 320 0 0 0 FrameData_O[0]
port 32 nsew signal output
flabel metal2 s 53190 4076 53280 4156 0 FreeSans 320 0 0 0 FrameData_O[10]
port 33 nsew signal output
flabel metal2 s 53190 4412 53280 4492 0 FreeSans 320 0 0 0 FrameData_O[11]
port 34 nsew signal output
flabel metal2 s 53190 4748 53280 4828 0 FreeSans 320 0 0 0 FrameData_O[12]
port 35 nsew signal output
flabel metal2 s 53190 5084 53280 5164 0 FreeSans 320 0 0 0 FrameData_O[13]
port 36 nsew signal output
flabel metal2 s 53190 5420 53280 5500 0 FreeSans 320 0 0 0 FrameData_O[14]
port 37 nsew signal output
flabel metal2 s 53190 5756 53280 5836 0 FreeSans 320 0 0 0 FrameData_O[15]
port 38 nsew signal output
flabel metal2 s 53190 6092 53280 6172 0 FreeSans 320 0 0 0 FrameData_O[16]
port 39 nsew signal output
flabel metal2 s 53190 6428 53280 6508 0 FreeSans 320 0 0 0 FrameData_O[17]
port 40 nsew signal output
flabel metal2 s 53190 6764 53280 6844 0 FreeSans 320 0 0 0 FrameData_O[18]
port 41 nsew signal output
flabel metal2 s 53190 7100 53280 7180 0 FreeSans 320 0 0 0 FrameData_O[19]
port 42 nsew signal output
flabel metal2 s 53190 1052 53280 1132 0 FreeSans 320 0 0 0 FrameData_O[1]
port 43 nsew signal output
flabel metal2 s 53190 7436 53280 7516 0 FreeSans 320 0 0 0 FrameData_O[20]
port 44 nsew signal output
flabel metal2 s 53190 7772 53280 7852 0 FreeSans 320 0 0 0 FrameData_O[21]
port 45 nsew signal output
flabel metal2 s 53190 8108 53280 8188 0 FreeSans 320 0 0 0 FrameData_O[22]
port 46 nsew signal output
flabel metal2 s 53190 8444 53280 8524 0 FreeSans 320 0 0 0 FrameData_O[23]
port 47 nsew signal output
flabel metal2 s 53190 8780 53280 8860 0 FreeSans 320 0 0 0 FrameData_O[24]
port 48 nsew signal output
flabel metal2 s 53190 9116 53280 9196 0 FreeSans 320 0 0 0 FrameData_O[25]
port 49 nsew signal output
flabel metal2 s 53190 9452 53280 9532 0 FreeSans 320 0 0 0 FrameData_O[26]
port 50 nsew signal output
flabel metal2 s 53190 9788 53280 9868 0 FreeSans 320 0 0 0 FrameData_O[27]
port 51 nsew signal output
flabel metal2 s 53190 10124 53280 10204 0 FreeSans 320 0 0 0 FrameData_O[28]
port 52 nsew signal output
flabel metal2 s 53190 10460 53280 10540 0 FreeSans 320 0 0 0 FrameData_O[29]
port 53 nsew signal output
flabel metal2 s 53190 1388 53280 1468 0 FreeSans 320 0 0 0 FrameData_O[2]
port 54 nsew signal output
flabel metal2 s 53190 10796 53280 10876 0 FreeSans 320 0 0 0 FrameData_O[30]
port 55 nsew signal output
flabel metal2 s 53190 11132 53280 11212 0 FreeSans 320 0 0 0 FrameData_O[31]
port 56 nsew signal output
flabel metal2 s 53190 1724 53280 1804 0 FreeSans 320 0 0 0 FrameData_O[3]
port 57 nsew signal output
flabel metal2 s 53190 2060 53280 2140 0 FreeSans 320 0 0 0 FrameData_O[4]
port 58 nsew signal output
flabel metal2 s 53190 2396 53280 2476 0 FreeSans 320 0 0 0 FrameData_O[5]
port 59 nsew signal output
flabel metal2 s 53190 2732 53280 2812 0 FreeSans 320 0 0 0 FrameData_O[6]
port 60 nsew signal output
flabel metal2 s 53190 3068 53280 3148 0 FreeSans 320 0 0 0 FrameData_O[7]
port 61 nsew signal output
flabel metal2 s 53190 3404 53280 3484 0 FreeSans 320 0 0 0 FrameData_O[8]
port 62 nsew signal output
flabel metal2 s 53190 3740 53280 3820 0 FreeSans 320 0 0 0 FrameData_O[9]
port 63 nsew signal output
flabel metal3 s 43064 0 43144 80 0 FreeSans 320 0 0 0 FrameStrobe[0]
port 64 nsew signal input
flabel metal3 s 46904 0 46984 80 0 FreeSans 320 0 0 0 FrameStrobe[10]
port 65 nsew signal input
flabel metal3 s 47288 0 47368 80 0 FreeSans 320 0 0 0 FrameStrobe[11]
port 66 nsew signal input
flabel metal3 s 47672 0 47752 80 0 FreeSans 320 0 0 0 FrameStrobe[12]
port 67 nsew signal input
flabel metal3 s 48056 0 48136 80 0 FreeSans 320 0 0 0 FrameStrobe[13]
port 68 nsew signal input
flabel metal3 s 48440 0 48520 80 0 FreeSans 320 0 0 0 FrameStrobe[14]
port 69 nsew signal input
flabel metal3 s 48824 0 48904 80 0 FreeSans 320 0 0 0 FrameStrobe[15]
port 70 nsew signal input
flabel metal3 s 49208 0 49288 80 0 FreeSans 320 0 0 0 FrameStrobe[16]
port 71 nsew signal input
flabel metal3 s 49592 0 49672 80 0 FreeSans 320 0 0 0 FrameStrobe[17]
port 72 nsew signal input
flabel metal3 s 49976 0 50056 80 0 FreeSans 320 0 0 0 FrameStrobe[18]
port 73 nsew signal input
flabel metal3 s 50360 0 50440 80 0 FreeSans 320 0 0 0 FrameStrobe[19]
port 74 nsew signal input
flabel metal3 s 43448 0 43528 80 0 FreeSans 320 0 0 0 FrameStrobe[1]
port 75 nsew signal input
flabel metal3 s 43832 0 43912 80 0 FreeSans 320 0 0 0 FrameStrobe[2]
port 76 nsew signal input
flabel metal3 s 44216 0 44296 80 0 FreeSans 320 0 0 0 FrameStrobe[3]
port 77 nsew signal input
flabel metal3 s 44600 0 44680 80 0 FreeSans 320 0 0 0 FrameStrobe[4]
port 78 nsew signal input
flabel metal3 s 44984 0 45064 80 0 FreeSans 320 0 0 0 FrameStrobe[5]
port 79 nsew signal input
flabel metal3 s 45368 0 45448 80 0 FreeSans 320 0 0 0 FrameStrobe[6]
port 80 nsew signal input
flabel metal3 s 45752 0 45832 80 0 FreeSans 320 0 0 0 FrameStrobe[7]
port 81 nsew signal input
flabel metal3 s 46136 0 46216 80 0 FreeSans 320 0 0 0 FrameStrobe[8]
port 82 nsew signal input
flabel metal3 s 46520 0 46600 80 0 FreeSans 320 0 0 0 FrameStrobe[9]
port 83 nsew signal input
flabel metal3 s 4088 12100 4168 12180 0 FreeSans 320 0 0 0 FrameStrobe_O[0]
port 84 nsew signal output
flabel metal3 s 29048 12100 29128 12180 0 FreeSans 320 0 0 0 FrameStrobe_O[10]
port 85 nsew signal output
flabel metal3 s 31544 12100 31624 12180 0 FreeSans 320 0 0 0 FrameStrobe_O[11]
port 86 nsew signal output
flabel metal3 s 34040 12100 34120 12180 0 FreeSans 320 0 0 0 FrameStrobe_O[12]
port 87 nsew signal output
flabel metal3 s 36536 12100 36616 12180 0 FreeSans 320 0 0 0 FrameStrobe_O[13]
port 88 nsew signal output
flabel metal3 s 39032 12100 39112 12180 0 FreeSans 320 0 0 0 FrameStrobe_O[14]
port 89 nsew signal output
flabel metal3 s 41528 12100 41608 12180 0 FreeSans 320 0 0 0 FrameStrobe_O[15]
port 90 nsew signal output
flabel metal3 s 44024 12100 44104 12180 0 FreeSans 320 0 0 0 FrameStrobe_O[16]
port 91 nsew signal output
flabel metal3 s 46520 12100 46600 12180 0 FreeSans 320 0 0 0 FrameStrobe_O[17]
port 92 nsew signal output
flabel metal3 s 49016 12100 49096 12180 0 FreeSans 320 0 0 0 FrameStrobe_O[18]
port 93 nsew signal output
flabel metal3 s 51512 12100 51592 12180 0 FreeSans 320 0 0 0 FrameStrobe_O[19]
port 94 nsew signal output
flabel metal3 s 6584 12100 6664 12180 0 FreeSans 320 0 0 0 FrameStrobe_O[1]
port 95 nsew signal output
flabel metal3 s 9080 12100 9160 12180 0 FreeSans 320 0 0 0 FrameStrobe_O[2]
port 96 nsew signal output
flabel metal3 s 11576 12100 11656 12180 0 FreeSans 320 0 0 0 FrameStrobe_O[3]
port 97 nsew signal output
flabel metal3 s 14072 12100 14152 12180 0 FreeSans 320 0 0 0 FrameStrobe_O[4]
port 98 nsew signal output
flabel metal3 s 16568 12100 16648 12180 0 FreeSans 320 0 0 0 FrameStrobe_O[5]
port 99 nsew signal output
flabel metal3 s 19064 12100 19144 12180 0 FreeSans 320 0 0 0 FrameStrobe_O[6]
port 100 nsew signal output
flabel metal3 s 21560 12100 21640 12180 0 FreeSans 320 0 0 0 FrameStrobe_O[7]
port 101 nsew signal output
flabel metal3 s 24056 12100 24136 12180 0 FreeSans 320 0 0 0 FrameStrobe_O[8]
port 102 nsew signal output
flabel metal3 s 26552 12100 26632 12180 0 FreeSans 320 0 0 0 FrameStrobe_O[9]
port 103 nsew signal output
flabel metal3 s 2744 0 2824 80 0 FreeSans 320 0 0 0 N1END[0]
port 104 nsew signal input
flabel metal3 s 3128 0 3208 80 0 FreeSans 320 0 0 0 N1END[1]
port 105 nsew signal input
flabel metal3 s 3512 0 3592 80 0 FreeSans 320 0 0 0 N1END[2]
port 106 nsew signal input
flabel metal3 s 3896 0 3976 80 0 FreeSans 320 0 0 0 N1END[3]
port 107 nsew signal input
flabel metal3 s 7352 0 7432 80 0 FreeSans 320 0 0 0 N2END[0]
port 108 nsew signal input
flabel metal3 s 7736 0 7816 80 0 FreeSans 320 0 0 0 N2END[1]
port 109 nsew signal input
flabel metal3 s 8120 0 8200 80 0 FreeSans 320 0 0 0 N2END[2]
port 110 nsew signal input
flabel metal3 s 8504 0 8584 80 0 FreeSans 320 0 0 0 N2END[3]
port 111 nsew signal input
flabel metal3 s 8888 0 8968 80 0 FreeSans 320 0 0 0 N2END[4]
port 112 nsew signal input
flabel metal3 s 9272 0 9352 80 0 FreeSans 320 0 0 0 N2END[5]
port 113 nsew signal input
flabel metal3 s 9656 0 9736 80 0 FreeSans 320 0 0 0 N2END[6]
port 114 nsew signal input
flabel metal3 s 10040 0 10120 80 0 FreeSans 320 0 0 0 N2END[7]
port 115 nsew signal input
flabel metal3 s 4280 0 4360 80 0 FreeSans 320 0 0 0 N2MID[0]
port 116 nsew signal input
flabel metal3 s 4664 0 4744 80 0 FreeSans 320 0 0 0 N2MID[1]
port 117 nsew signal input
flabel metal3 s 5048 0 5128 80 0 FreeSans 320 0 0 0 N2MID[2]
port 118 nsew signal input
flabel metal3 s 5432 0 5512 80 0 FreeSans 320 0 0 0 N2MID[3]
port 119 nsew signal input
flabel metal3 s 5816 0 5896 80 0 FreeSans 320 0 0 0 N2MID[4]
port 120 nsew signal input
flabel metal3 s 6200 0 6280 80 0 FreeSans 320 0 0 0 N2MID[5]
port 121 nsew signal input
flabel metal3 s 6584 0 6664 80 0 FreeSans 320 0 0 0 N2MID[6]
port 122 nsew signal input
flabel metal3 s 6968 0 7048 80 0 FreeSans 320 0 0 0 N2MID[7]
port 123 nsew signal input
flabel metal3 s 10424 0 10504 80 0 FreeSans 320 0 0 0 N4END[0]
port 124 nsew signal input
flabel metal3 s 14264 0 14344 80 0 FreeSans 320 0 0 0 N4END[10]
port 125 nsew signal input
flabel metal3 s 14648 0 14728 80 0 FreeSans 320 0 0 0 N4END[11]
port 126 nsew signal input
flabel metal3 s 15032 0 15112 80 0 FreeSans 320 0 0 0 N4END[12]
port 127 nsew signal input
flabel metal3 s 15416 0 15496 80 0 FreeSans 320 0 0 0 N4END[13]
port 128 nsew signal input
flabel metal3 s 15800 0 15880 80 0 FreeSans 320 0 0 0 N4END[14]
port 129 nsew signal input
flabel metal3 s 16184 0 16264 80 0 FreeSans 320 0 0 0 N4END[15]
port 130 nsew signal input
flabel metal3 s 10808 0 10888 80 0 FreeSans 320 0 0 0 N4END[1]
port 131 nsew signal input
flabel metal3 s 11192 0 11272 80 0 FreeSans 320 0 0 0 N4END[2]
port 132 nsew signal input
flabel metal3 s 11576 0 11656 80 0 FreeSans 320 0 0 0 N4END[3]
port 133 nsew signal input
flabel metal3 s 11960 0 12040 80 0 FreeSans 320 0 0 0 N4END[4]
port 134 nsew signal input
flabel metal3 s 12344 0 12424 80 0 FreeSans 320 0 0 0 N4END[5]
port 135 nsew signal input
flabel metal3 s 12728 0 12808 80 0 FreeSans 320 0 0 0 N4END[6]
port 136 nsew signal input
flabel metal3 s 13112 0 13192 80 0 FreeSans 320 0 0 0 N4END[7]
port 137 nsew signal input
flabel metal3 s 13496 0 13576 80 0 FreeSans 320 0 0 0 N4END[8]
port 138 nsew signal input
flabel metal3 s 13880 0 13960 80 0 FreeSans 320 0 0 0 N4END[9]
port 139 nsew signal input
flabel metal3 s 16568 0 16648 80 0 FreeSans 320 0 0 0 NN4END[0]
port 140 nsew signal input
flabel metal3 s 20408 0 20488 80 0 FreeSans 320 0 0 0 NN4END[10]
port 141 nsew signal input
flabel metal3 s 20792 0 20872 80 0 FreeSans 320 0 0 0 NN4END[11]
port 142 nsew signal input
flabel metal3 s 21176 0 21256 80 0 FreeSans 320 0 0 0 NN4END[12]
port 143 nsew signal input
flabel metal3 s 21560 0 21640 80 0 FreeSans 320 0 0 0 NN4END[13]
port 144 nsew signal input
flabel metal3 s 21944 0 22024 80 0 FreeSans 320 0 0 0 NN4END[14]
port 145 nsew signal input
flabel metal3 s 22328 0 22408 80 0 FreeSans 320 0 0 0 NN4END[15]
port 146 nsew signal input
flabel metal3 s 16952 0 17032 80 0 FreeSans 320 0 0 0 NN4END[1]
port 147 nsew signal input
flabel metal3 s 17336 0 17416 80 0 FreeSans 320 0 0 0 NN4END[2]
port 148 nsew signal input
flabel metal3 s 17720 0 17800 80 0 FreeSans 320 0 0 0 NN4END[3]
port 149 nsew signal input
flabel metal3 s 18104 0 18184 80 0 FreeSans 320 0 0 0 NN4END[4]
port 150 nsew signal input
flabel metal3 s 18488 0 18568 80 0 FreeSans 320 0 0 0 NN4END[5]
port 151 nsew signal input
flabel metal3 s 18872 0 18952 80 0 FreeSans 320 0 0 0 NN4END[6]
port 152 nsew signal input
flabel metal3 s 19256 0 19336 80 0 FreeSans 320 0 0 0 NN4END[7]
port 153 nsew signal input
flabel metal3 s 19640 0 19720 80 0 FreeSans 320 0 0 0 NN4END[8]
port 154 nsew signal input
flabel metal3 s 20024 0 20104 80 0 FreeSans 320 0 0 0 NN4END[9]
port 155 nsew signal input
flabel metal3 s 22712 0 22792 80 0 FreeSans 320 0 0 0 S1BEG[0]
port 156 nsew signal output
flabel metal3 s 23096 0 23176 80 0 FreeSans 320 0 0 0 S1BEG[1]
port 157 nsew signal output
flabel metal3 s 23480 0 23560 80 0 FreeSans 320 0 0 0 S1BEG[2]
port 158 nsew signal output
flabel metal3 s 23864 0 23944 80 0 FreeSans 320 0 0 0 S1BEG[3]
port 159 nsew signal output
flabel metal3 s 24248 0 24328 80 0 FreeSans 320 0 0 0 S2BEG[0]
port 160 nsew signal output
flabel metal3 s 24632 0 24712 80 0 FreeSans 320 0 0 0 S2BEG[1]
port 161 nsew signal output
flabel metal3 s 25016 0 25096 80 0 FreeSans 320 0 0 0 S2BEG[2]
port 162 nsew signal output
flabel metal3 s 25400 0 25480 80 0 FreeSans 320 0 0 0 S2BEG[3]
port 163 nsew signal output
flabel metal3 s 25784 0 25864 80 0 FreeSans 320 0 0 0 S2BEG[4]
port 164 nsew signal output
flabel metal3 s 26168 0 26248 80 0 FreeSans 320 0 0 0 S2BEG[5]
port 165 nsew signal output
flabel metal3 s 26552 0 26632 80 0 FreeSans 320 0 0 0 S2BEG[6]
port 166 nsew signal output
flabel metal3 s 26936 0 27016 80 0 FreeSans 320 0 0 0 S2BEG[7]
port 167 nsew signal output
flabel metal3 s 27320 0 27400 80 0 FreeSans 320 0 0 0 S2BEGb[0]
port 168 nsew signal output
flabel metal3 s 27704 0 27784 80 0 FreeSans 320 0 0 0 S2BEGb[1]
port 169 nsew signal output
flabel metal3 s 28088 0 28168 80 0 FreeSans 320 0 0 0 S2BEGb[2]
port 170 nsew signal output
flabel metal3 s 28472 0 28552 80 0 FreeSans 320 0 0 0 S2BEGb[3]
port 171 nsew signal output
flabel metal3 s 28856 0 28936 80 0 FreeSans 320 0 0 0 S2BEGb[4]
port 172 nsew signal output
flabel metal3 s 29240 0 29320 80 0 FreeSans 320 0 0 0 S2BEGb[5]
port 173 nsew signal output
flabel metal3 s 29624 0 29704 80 0 FreeSans 320 0 0 0 S2BEGb[6]
port 174 nsew signal output
flabel metal3 s 30008 0 30088 80 0 FreeSans 320 0 0 0 S2BEGb[7]
port 175 nsew signal output
flabel metal3 s 30392 0 30472 80 0 FreeSans 320 0 0 0 S4BEG[0]
port 176 nsew signal output
flabel metal3 s 34232 0 34312 80 0 FreeSans 320 0 0 0 S4BEG[10]
port 177 nsew signal output
flabel metal3 s 34616 0 34696 80 0 FreeSans 320 0 0 0 S4BEG[11]
port 178 nsew signal output
flabel metal3 s 35000 0 35080 80 0 FreeSans 320 0 0 0 S4BEG[12]
port 179 nsew signal output
flabel metal3 s 35384 0 35464 80 0 FreeSans 320 0 0 0 S4BEG[13]
port 180 nsew signal output
flabel metal3 s 35768 0 35848 80 0 FreeSans 320 0 0 0 S4BEG[14]
port 181 nsew signal output
flabel metal3 s 36152 0 36232 80 0 FreeSans 320 0 0 0 S4BEG[15]
port 182 nsew signal output
flabel metal3 s 30776 0 30856 80 0 FreeSans 320 0 0 0 S4BEG[1]
port 183 nsew signal output
flabel metal3 s 31160 0 31240 80 0 FreeSans 320 0 0 0 S4BEG[2]
port 184 nsew signal output
flabel metal3 s 31544 0 31624 80 0 FreeSans 320 0 0 0 S4BEG[3]
port 185 nsew signal output
flabel metal3 s 31928 0 32008 80 0 FreeSans 320 0 0 0 S4BEG[4]
port 186 nsew signal output
flabel metal3 s 32312 0 32392 80 0 FreeSans 320 0 0 0 S4BEG[5]
port 187 nsew signal output
flabel metal3 s 32696 0 32776 80 0 FreeSans 320 0 0 0 S4BEG[6]
port 188 nsew signal output
flabel metal3 s 33080 0 33160 80 0 FreeSans 320 0 0 0 S4BEG[7]
port 189 nsew signal output
flabel metal3 s 33464 0 33544 80 0 FreeSans 320 0 0 0 S4BEG[8]
port 190 nsew signal output
flabel metal3 s 33848 0 33928 80 0 FreeSans 320 0 0 0 S4BEG[9]
port 191 nsew signal output
flabel metal3 s 36536 0 36616 80 0 FreeSans 320 0 0 0 SS4BEG[0]
port 192 nsew signal output
flabel metal3 s 40376 0 40456 80 0 FreeSans 320 0 0 0 SS4BEG[10]
port 193 nsew signal output
flabel metal3 s 40760 0 40840 80 0 FreeSans 320 0 0 0 SS4BEG[11]
port 194 nsew signal output
flabel metal3 s 41144 0 41224 80 0 FreeSans 320 0 0 0 SS4BEG[12]
port 195 nsew signal output
flabel metal3 s 41528 0 41608 80 0 FreeSans 320 0 0 0 SS4BEG[13]
port 196 nsew signal output
flabel metal3 s 41912 0 41992 80 0 FreeSans 320 0 0 0 SS4BEG[14]
port 197 nsew signal output
flabel metal3 s 42296 0 42376 80 0 FreeSans 320 0 0 0 SS4BEG[15]
port 198 nsew signal output
flabel metal3 s 36920 0 37000 80 0 FreeSans 320 0 0 0 SS4BEG[1]
port 199 nsew signal output
flabel metal3 s 37304 0 37384 80 0 FreeSans 320 0 0 0 SS4BEG[2]
port 200 nsew signal output
flabel metal3 s 37688 0 37768 80 0 FreeSans 320 0 0 0 SS4BEG[3]
port 201 nsew signal output
flabel metal3 s 38072 0 38152 80 0 FreeSans 320 0 0 0 SS4BEG[4]
port 202 nsew signal output
flabel metal3 s 38456 0 38536 80 0 FreeSans 320 0 0 0 SS4BEG[5]
port 203 nsew signal output
flabel metal3 s 38840 0 38920 80 0 FreeSans 320 0 0 0 SS4BEG[6]
port 204 nsew signal output
flabel metal3 s 39224 0 39304 80 0 FreeSans 320 0 0 0 SS4BEG[7]
port 205 nsew signal output
flabel metal3 s 39608 0 39688 80 0 FreeSans 320 0 0 0 SS4BEG[8]
port 206 nsew signal output
flabel metal3 s 39992 0 40072 80 0 FreeSans 320 0 0 0 SS4BEG[9]
port 207 nsew signal output
flabel metal3 s 42680 0 42760 80 0 FreeSans 320 0 0 0 UserCLK
port 208 nsew signal input
flabel metal3 s 1592 12100 1672 12180 0 FreeSans 320 0 0 0 UserCLKo
port 209 nsew signal output
flabel metal5 s 4892 0 5332 12180 0 FreeSans 2560 90 0 0 VGND
port 210 nsew ground bidirectional
flabel metal5 s 4892 0 5332 40 0 FreeSans 320 0 0 0 VGND
port 210 nsew ground bidirectional
flabel metal5 s 4892 12140 5332 12180 0 FreeSans 320 0 0 0 VGND
port 210 nsew ground bidirectional
flabel metal5 s 20012 0 20452 12180 0 FreeSans 2560 90 0 0 VGND
port 210 nsew ground bidirectional
flabel metal5 s 20012 0 20452 40 0 FreeSans 320 0 0 0 VGND
port 210 nsew ground bidirectional
flabel metal5 s 20012 12140 20452 12180 0 FreeSans 320 0 0 0 VGND
port 210 nsew ground bidirectional
flabel metal5 s 35132 0 35572 12180 0 FreeSans 2560 90 0 0 VGND
port 210 nsew ground bidirectional
flabel metal5 s 35132 0 35572 40 0 FreeSans 320 0 0 0 VGND
port 210 nsew ground bidirectional
flabel metal5 s 35132 12140 35572 12180 0 FreeSans 320 0 0 0 VGND
port 210 nsew ground bidirectional
flabel metal5 s 50252 0 50692 12180 0 FreeSans 2560 90 0 0 VGND
port 210 nsew ground bidirectional
flabel metal5 s 50252 0 50692 40 0 FreeSans 320 0 0 0 VGND
port 210 nsew ground bidirectional
flabel metal5 s 50252 12140 50692 12180 0 FreeSans 320 0 0 0 VGND
port 210 nsew ground bidirectional
flabel metal5 s 3652 0 4092 12180 0 FreeSans 2560 90 0 0 VPWR
port 211 nsew power bidirectional
flabel metal5 s 3652 0 4092 40 0 FreeSans 320 0 0 0 VPWR
port 211 nsew power bidirectional
flabel metal5 s 3652 12140 4092 12180 0 FreeSans 320 0 0 0 VPWR
port 211 nsew power bidirectional
flabel metal5 s 18772 0 19212 12180 0 FreeSans 2560 90 0 0 VPWR
port 211 nsew power bidirectional
flabel metal5 s 18772 0 19212 40 0 FreeSans 320 0 0 0 VPWR
port 211 nsew power bidirectional
flabel metal5 s 18772 12140 19212 12180 0 FreeSans 320 0 0 0 VPWR
port 211 nsew power bidirectional
flabel metal5 s 33892 0 34332 12180 0 FreeSans 2560 90 0 0 VPWR
port 211 nsew power bidirectional
flabel metal5 s 33892 0 34332 40 0 FreeSans 320 0 0 0 VPWR
port 211 nsew power bidirectional
flabel metal5 s 33892 12140 34332 12180 0 FreeSans 320 0 0 0 VPWR
port 211 nsew power bidirectional
flabel metal5 s 49012 0 49452 12180 0 FreeSans 2560 90 0 0 VPWR
port 211 nsew power bidirectional
flabel metal5 s 49012 0 49452 40 0 FreeSans 320 0 0 0 VPWR
port 211 nsew power bidirectional
flabel metal5 s 49012 12140 49452 12180 0 FreeSans 320 0 0 0 VPWR
port 211 nsew power bidirectional
rlabel metal1 26640 10584 26640 10584 0 VGND
rlabel metal1 26640 9828 26640 9828 0 VPWR
rlabel metal2 416 756 416 756 0 FrameData[0]
rlabel metal2 272 4116 272 4116 0 FrameData[10]
rlabel metal2 224 4452 224 4452 0 FrameData[11]
rlabel metal2 560 4788 560 4788 0 FrameData[12]
rlabel metal2 608 5124 608 5124 0 FrameData[13]
rlabel metal3 10752 6300 10752 6300 0 FrameData[14]
rlabel metal3 22752 6132 22752 6132 0 FrameData[15]
rlabel metal3 25824 6300 25824 6300 0 FrameData[16]
rlabel metal2 752 6468 752 6468 0 FrameData[17]
rlabel metal2 1808 6804 1808 6804 0 FrameData[18]
rlabel metal2 656 7140 656 7140 0 FrameData[19]
rlabel metal2 752 1092 752 1092 0 FrameData[1]
rlabel metal3 22944 6972 22944 6972 0 FrameData[20]
rlabel metal3 21600 7476 21600 7476 0 FrameData[21]
rlabel metal2 704 8148 704 8148 0 FrameData[22]
rlabel metal2 23328 8232 23328 8232 0 FrameData[23]
rlabel metal2 656 8820 656 8820 0 FrameData[24]
rlabel metal2 128 9156 128 9156 0 FrameData[25]
rlabel metal2 3632 9492 3632 9492 0 FrameData[26]
rlabel metal2 128 9828 128 9828 0 FrameData[27]
rlabel metal2 848 10164 848 10164 0 FrameData[28]
rlabel metal3 14304 9996 14304 9996 0 FrameData[29]
rlabel metal2 752 1428 752 1428 0 FrameData[2]
rlabel metal3 23616 10164 23616 10164 0 FrameData[30]
rlabel metal2 464 11172 464 11172 0 FrameData[31]
rlabel metal2 752 1764 752 1764 0 FrameData[3]
rlabel metal2 1376 2100 1376 2100 0 FrameData[4]
rlabel metal2 752 2436 752 2436 0 FrameData[5]
rlabel metal2 752 2772 752 2772 0 FrameData[6]
rlabel metal2 33360 7728 33360 7728 0 FrameData[7]
rlabel metal2 176 3444 176 3444 0 FrameData[8]
rlabel metal2 416 3780 416 3780 0 FrameData[9]
rlabel metal2 52767 756 52767 756 0 FrameData_O[0]
rlabel metal2 52863 4116 52863 4116 0 FrameData_O[10]
rlabel metal2 52080 4368 52080 4368 0 FrameData_O[11]
rlabel metal2 52455 4788 52455 4788 0 FrameData_O[12]
rlabel metal2 52647 5124 52647 5124 0 FrameData_O[13]
rlabel metal2 52863 5460 52863 5460 0 FrameData_O[14]
rlabel metal2 52647 5796 52647 5796 0 FrameData_O[15]
rlabel metal2 52455 6132 52455 6132 0 FrameData_O[16]
rlabel metal2 52647 6468 52647 6468 0 FrameData_O[17]
rlabel metal2 53151 6804 53151 6804 0 FrameData_O[18]
rlabel metal2 52647 7140 52647 7140 0 FrameData_O[19]
rlabel metal2 52575 1092 52575 1092 0 FrameData_O[1]
rlabel via2 53199 7476 53199 7476 0 FrameData_O[20]
rlabel metal2 52455 7812 52455 7812 0 FrameData_O[21]
rlabel via2 53199 8148 53199 8148 0 FrameData_O[22]
rlabel metal2 52863 8484 52863 8484 0 FrameData_O[23]
rlabel metal2 52959 8820 52959 8820 0 FrameData_O[24]
rlabel metal2 52455 9156 52455 9156 0 FrameData_O[25]
rlabel metal2 52575 9492 52575 9492 0 FrameData_O[26]
rlabel metal2 53151 9828 53151 9828 0 FrameData_O[27]
rlabel metal2 53151 10164 53151 10164 0 FrameData_O[28]
rlabel metal2 50544 10458 50544 10458 0 FrameData_O[29]
rlabel metal2 52911 1428 52911 1428 0 FrameData_O[2]
rlabel metal2 51000 10416 51000 10416 0 FrameData_O[30]
rlabel metal2 50904 9660 50904 9660 0 FrameData_O[31]
rlabel metal2 52815 1764 52815 1764 0 FrameData_O[3]
rlabel metal2 52647 2100 52647 2100 0 FrameData_O[4]
rlabel metal2 52959 2436 52959 2436 0 FrameData_O[5]
rlabel metal2 52647 2772 52647 2772 0 FrameData_O[6]
rlabel metal2 52455 3108 52455 3108 0 FrameData_O[7]
rlabel metal2 52575 3444 52575 3444 0 FrameData_O[8]
rlabel metal2 52080 3696 52080 3696 0 FrameData_O[9]
rlabel metal2 42432 9660 42432 9660 0 FrameStrobe[0]
rlabel metal3 38016 8820 38016 8820 0 FrameStrobe[10]
rlabel metal2 46752 9156 46752 9156 0 FrameStrobe[11]
rlabel metal2 46464 9576 46464 9576 0 FrameStrobe[12]
rlabel metal3 48096 4692 48096 4692 0 FrameStrobe[13]
rlabel metal2 47904 9408 47904 9408 0 FrameStrobe[14]
rlabel metal2 46512 9072 46512 9072 0 FrameStrobe[15]
rlabel metal3 49248 1080 49248 1080 0 FrameStrobe[16]
rlabel metal2 49104 9408 49104 9408 0 FrameStrobe[17]
rlabel metal2 49344 9492 49344 9492 0 FrameStrobe[18]
rlabel via3 50400 72 50400 72 0 FrameStrobe[19]
rlabel metal2 41856 9534 41856 9534 0 FrameStrobe[1]
rlabel metal2 43584 9534 43584 9534 0 FrameStrobe[2]
rlabel via3 44256 72 44256 72 0 FrameStrobe[3]
rlabel metal2 15840 9492 15840 9492 0 FrameStrobe[4]
rlabel metal3 45024 114 45024 114 0 FrameStrobe[5]
rlabel via2 45408 72 45408 72 0 FrameStrobe[6]
rlabel metal3 45792 114 45792 114 0 FrameStrobe[7]
rlabel metal3 46176 156 46176 156 0 FrameStrobe[8]
rlabel metal2 38208 9156 38208 9156 0 FrameStrobe[9]
rlabel metal2 4152 10416 4152 10416 0 FrameStrobe_O[0]
rlabel metal2 29112 10416 29112 10416 0 FrameStrobe_O[10]
rlabel metal2 31608 10416 31608 10416 0 FrameStrobe_O[11]
rlabel metal2 34104 10416 34104 10416 0 FrameStrobe_O[12]
rlabel metal2 36600 10164 36600 10164 0 FrameStrobe_O[13]
rlabel metal2 39096 10416 39096 10416 0 FrameStrobe_O[14]
rlabel metal2 41592 10416 41592 10416 0 FrameStrobe_O[15]
rlabel metal2 44088 10416 44088 10416 0 FrameStrobe_O[16]
rlabel metal2 46584 10416 46584 10416 0 FrameStrobe_O[17]
rlabel metal2 49080 10416 49080 10416 0 FrameStrobe_O[18]
rlabel metal2 51672 10416 51672 10416 0 FrameStrobe_O[19]
rlabel metal2 6648 10416 6648 10416 0 FrameStrobe_O[1]
rlabel metal2 9144 10416 9144 10416 0 FrameStrobe_O[2]
rlabel metal2 11640 10416 11640 10416 0 FrameStrobe_O[3]
rlabel metal2 14136 10416 14136 10416 0 FrameStrobe_O[4]
rlabel metal2 16632 10416 16632 10416 0 FrameStrobe_O[5]
rlabel metal2 19128 10416 19128 10416 0 FrameStrobe_O[6]
rlabel metal2 21624 10416 21624 10416 0 FrameStrobe_O[7]
rlabel metal2 24120 10416 24120 10416 0 FrameStrobe_O[8]
rlabel metal2 26616 10416 26616 10416 0 FrameStrobe_O[9]
rlabel metal3 2784 1122 2784 1122 0 N1END[0]
rlabel metal3 3168 954 3168 954 0 N1END[1]
rlabel metal3 3552 954 3552 954 0 N1END[2]
rlabel metal3 3936 114 3936 114 0 N1END[3]
rlabel metal3 7392 1332 7392 1332 0 N2END[0]
rlabel metal3 7776 828 7776 828 0 N2END[1]
rlabel metal3 8160 1500 8160 1500 0 N2END[2]
rlabel metal3 8544 2088 8544 2088 0 N2END[3]
rlabel metal3 8928 1038 8928 1038 0 N2END[4]
rlabel metal3 9312 996 9312 996 0 N2END[5]
rlabel metal3 9696 156 9696 156 0 N2END[6]
rlabel metal3 22560 1974 22560 1974 0 N2END[7]
rlabel metal3 4320 828 4320 828 0 N2MID[0]
rlabel metal3 4704 282 4704 282 0 N2MID[1]
rlabel metal3 5088 240 5088 240 0 N2MID[2]
rlabel metal3 5472 2466 5472 2466 0 N2MID[3]
rlabel metal3 5856 2424 5856 2424 0 N2MID[4]
rlabel metal3 6240 2256 6240 2256 0 N2MID[5]
rlabel metal3 6624 2172 6624 2172 0 N2MID[6]
rlabel metal3 7008 1500 7008 1500 0 N2MID[7]
rlabel metal3 10464 1794 10464 1794 0 N4END[0]
rlabel metal2 16512 3780 16512 3780 0 N4END[10]
rlabel metal3 14688 324 14688 324 0 N4END[11]
rlabel metal2 11808 2730 11808 2730 0 N4END[12]
rlabel metal3 15456 1416 15456 1416 0 N4END[13]
rlabel metal3 15840 1332 15840 1332 0 N4END[14]
rlabel metal3 16224 1374 16224 1374 0 N4END[15]
rlabel metal3 10848 1710 10848 1710 0 N4END[1]
rlabel metal3 11232 1668 11232 1668 0 N4END[2]
rlabel metal3 11616 2130 11616 2130 0 N4END[3]
rlabel metal3 12000 156 12000 156 0 N4END[4]
rlabel metal3 12384 1290 12384 1290 0 N4END[5]
rlabel metal3 12768 1962 12768 1962 0 N4END[6]
rlabel metal3 13152 870 13152 870 0 N4END[7]
rlabel metal3 13536 114 13536 114 0 N4END[8]
rlabel metal4 15600 3528 15600 3528 0 N4END[9]
rlabel metal3 16608 1470 16608 1470 0 NN4END[0]
rlabel metal3 20448 576 20448 576 0 NN4END[10]
rlabel metal2 21696 3612 21696 3612 0 NN4END[11]
rlabel metal3 39744 1470 39744 1470 0 NN4END[12]
rlabel metal3 36288 1470 36288 1470 0 NN4END[13]
rlabel metal2 22416 3780 22416 3780 0 NN4END[14]
rlabel metal3 22368 1248 22368 1248 0 NN4END[15]
rlabel metal2 15600 3528 15600 3528 0 NN4END[1]
rlabel metal3 17376 1470 17376 1470 0 NN4END[2]
rlabel metal2 16224 4620 16224 4620 0 NN4END[3]
rlabel metal2 16704 4956 16704 4956 0 NN4END[4]
rlabel metal2 17472 4200 17472 4200 0 NN4END[5]
rlabel metal3 18912 114 18912 114 0 NN4END[6]
rlabel metal3 19296 1332 19296 1332 0 NN4END[7]
rlabel metal3 19680 1080 19680 1080 0 NN4END[8]
rlabel metal3 20064 702 20064 702 0 NN4END[9]
rlabel metal3 22752 870 22752 870 0 S1BEG[0]
rlabel metal3 23136 870 23136 870 0 S1BEG[1]
rlabel metal3 23520 870 23520 870 0 S1BEG[2]
rlabel metal3 23904 870 23904 870 0 S1BEG[3]
rlabel metal3 24288 870 24288 870 0 S2BEG[0]
rlabel metal3 24672 870 24672 870 0 S2BEG[1]
rlabel metal3 25056 870 25056 870 0 S2BEG[2]
rlabel metal3 25440 870 25440 870 0 S2BEG[3]
rlabel metal3 25824 870 25824 870 0 S2BEG[4]
rlabel metal3 26208 870 26208 870 0 S2BEG[5]
rlabel metal3 26592 870 26592 870 0 S2BEG[6]
rlabel metal3 26976 870 26976 870 0 S2BEG[7]
rlabel metal3 27360 870 27360 870 0 S2BEGb[0]
rlabel metal3 27744 870 27744 870 0 S2BEGb[1]
rlabel metal3 28128 870 28128 870 0 S2BEGb[2]
rlabel metal3 28512 870 28512 870 0 S2BEGb[3]
rlabel metal3 28896 870 28896 870 0 S2BEGb[4]
rlabel metal3 29280 870 29280 870 0 S2BEGb[5]
rlabel metal3 29664 870 29664 870 0 S2BEGb[6]
rlabel metal3 30048 870 30048 870 0 S2BEGb[7]
rlabel metal3 30432 870 30432 870 0 S4BEG[0]
rlabel metal3 34272 870 34272 870 0 S4BEG[10]
rlabel metal3 34656 870 34656 870 0 S4BEG[11]
rlabel metal3 35040 870 35040 870 0 S4BEG[12]
rlabel metal3 35424 114 35424 114 0 S4BEG[13]
rlabel metal3 35808 870 35808 870 0 S4BEG[14]
rlabel metal3 36192 870 36192 870 0 S4BEG[15]
rlabel metal3 30816 870 30816 870 0 S4BEG[1]
rlabel metal3 31200 870 31200 870 0 S4BEG[2]
rlabel metal3 31584 870 31584 870 0 S4BEG[3]
rlabel metal3 31968 870 31968 870 0 S4BEG[4]
rlabel metal3 32352 870 32352 870 0 S4BEG[5]
rlabel metal3 32736 870 32736 870 0 S4BEG[6]
rlabel metal2 33144 1680 33144 1680 0 S4BEG[7]
rlabel metal3 33504 870 33504 870 0 S4BEG[8]
rlabel metal3 33888 870 33888 870 0 S4BEG[9]
rlabel metal3 36576 870 36576 870 0 SS4BEG[0]
rlabel metal3 40416 870 40416 870 0 SS4BEG[10]
rlabel metal3 40800 870 40800 870 0 SS4BEG[11]
rlabel metal3 41184 870 41184 870 0 SS4BEG[12]
rlabel metal3 41568 870 41568 870 0 SS4BEG[13]
rlabel metal3 41952 870 41952 870 0 SS4BEG[14]
rlabel metal3 42336 870 42336 870 0 SS4BEG[15]
rlabel metal3 36960 870 36960 870 0 SS4BEG[1]
rlabel metal3 37344 870 37344 870 0 SS4BEG[2]
rlabel metal3 37728 870 37728 870 0 SS4BEG[3]
rlabel metal3 38112 870 38112 870 0 SS4BEG[4]
rlabel metal3 38496 870 38496 870 0 SS4BEG[5]
rlabel metal3 38880 870 38880 870 0 SS4BEG[6]
rlabel metal3 39264 870 39264 870 0 SS4BEG[7]
rlabel metal3 39648 870 39648 870 0 SS4BEG[8]
rlabel metal3 40032 870 40032 870 0 SS4BEG[9]
rlabel metal2 41520 9408 41520 9408 0 UserCLK
rlabel metal2 1656 10416 1656 10416 0 UserCLKo
rlabel metal3 4800 2100 4800 2100 0 net1
rlabel metal2 35136 7182 35136 7182 0 net10
rlabel metal3 37968 1512 37968 1512 0 net100
rlabel metal3 39168 2310 39168 2310 0 net101
rlabel metal3 39552 1764 39552 1764 0 net102
rlabel metal2 39552 2058 39552 2058 0 net103
rlabel metal3 40320 2310 40320 2310 0 net104
rlabel metal3 1920 9702 1920 9702 0 net105
rlabel metal2 33120 5418 33120 5418 0 net11
rlabel metal3 42432 2436 42432 2436 0 net12
rlabel metal2 25704 6552 25704 6552 0 net13
rlabel metal3 35136 7896 35136 7896 0 net14
rlabel metal3 51840 7854 51840 7854 0 net15
rlabel metal3 35040 9450 35040 9450 0 net16
rlabel metal3 51648 8820 51648 8820 0 net17
rlabel metal2 51456 9156 51456 9156 0 net18
rlabel metal3 38304 9660 38304 9660 0 net19
rlabel metal3 44256 6006 44256 6006 0 net2
rlabel metal2 28224 8778 28224 8778 0 net20
rlabel metal2 38112 9954 38112 9954 0 net21
rlabel metal2 15048 9492 15048 9492 0 net22
rlabel metal2 51072 2688 51072 2688 0 net23
rlabel metal2 36768 10374 36768 10374 0 net24
rlabel metal3 38064 9996 38064 9996 0 net25
rlabel metal2 49776 1932 49776 1932 0 net26
rlabel metal2 49056 2562 49056 2562 0 net27
rlabel metal2 50448 2520 50448 2520 0 net28
rlabel metal2 51984 2604 51984 2604 0 net29
rlabel metal3 38112 7854 38112 7854 0 net3
rlabel metal3 47232 6174 47232 6174 0 net30
rlabel metal3 47520 5208 47520 5208 0 net31
rlabel metal2 33024 4326 33024 4326 0 net32
rlabel metal3 4416 9744 4416 9744 0 net33
rlabel metal2 29544 9660 29544 9660 0 net34
rlabel metal2 33120 10122 33120 10122 0 net35
rlabel metal3 36864 10500 36864 10500 0 net36
rlabel metal3 39168 10374 39168 10374 0 net37
rlabel metal2 39360 10206 39360 10206 0 net38
rlabel metal2 43416 9660 43416 9660 0 net39
rlabel metal2 33120 6930 33120 6930 0 net4
rlabel metal2 46680 9660 46680 9660 0 net40
rlabel metal2 48216 9660 48216 9660 0 net41
rlabel metal2 48936 9660 48936 9660 0 net42
rlabel metal2 51432 9660 51432 9660 0 net43
rlabel metal3 6912 9870 6912 9870 0 net44
rlabel metal3 9408 9954 9408 9954 0 net45
rlabel metal2 13752 9660 13752 9660 0 net46
rlabel metal2 15096 9660 15096 9660 0 net47
rlabel metal2 18456 9660 18456 9660 0 net48
rlabel metal2 20856 9660 20856 9660 0 net49
rlabel metal2 33120 5040 33120 5040 0 net5
rlabel metal2 23160 9660 23160 9660 0 net50
rlabel metal2 25320 9660 25320 9660 0 net51
rlabel metal2 27864 9660 27864 9660 0 net52
rlabel metal2 19464 3192 19464 3192 0 net53
rlabel metal3 21216 2352 21216 2352 0 net54
rlabel metal3 22080 2688 22080 2688 0 net55
rlabel metal3 21888 2352 21888 2352 0 net56
rlabel metal3 22464 3066 22464 3066 0 net57
rlabel metal2 24528 1848 24528 1848 0 net58
rlabel metal2 25104 2016 25104 2016 0 net59
rlabel metal3 19968 6258 19968 6258 0 net6
rlabel metal2 25632 1932 25632 1932 0 net60
rlabel metal2 25728 4620 25728 4620 0 net61
rlabel metal3 26496 2352 26496 2352 0 net62
rlabel metal3 26880 2394 26880 2394 0 net63
rlabel metal2 27120 1932 27120 1932 0 net64
rlabel metal2 27648 1890 27648 1890 0 net65
rlabel metal3 28032 2310 28032 2310 0 net66
rlabel metal3 28416 2142 28416 2142 0 net67
rlabel metal2 28824 1932 28824 1932 0 net68
rlabel metal3 29184 2940 29184 2940 0 net69
rlabel metal3 22944 5964 22944 5964 0 net7
rlabel metal2 29136 1848 29136 1848 0 net70
rlabel metal2 29904 1932 29904 1932 0 net71
rlabel metal3 30336 2184 30336 2184 0 net72
rlabel metal2 21312 2772 21312 2772 0 net73
rlabel via1 34488 1932 34488 1932 0 net74
rlabel via1 34872 1932 34872 1932 0 net75
rlabel metal2 35184 1932 35184 1932 0 net76
rlabel metal2 35640 3192 35640 3192 0 net77
rlabel metal2 36072 3192 36072 3192 0 net78
rlabel metal2 36600 3192 36600 3192 0 net79
rlabel metal2 34632 6300 34632 6300 0 net8
rlabel metal2 14928 2394 14928 2394 0 net80
rlabel metal3 18432 2058 18432 2058 0 net81
rlabel metal2 13248 2310 13248 2310 0 net82
rlabel metal2 31848 3276 31848 3276 0 net83
rlabel metal2 32592 1932 32592 1932 0 net84
rlabel metal2 32856 3192 32856 3192 0 net85
rlabel metal2 33288 3192 33288 3192 0 net86
rlabel metal2 33744 1932 33744 1932 0 net87
rlabel metal2 34272 1932 34272 1932 0 net88
rlabel metal2 36864 1974 36864 1974 0 net89
rlabel metal2 36744 4788 36744 4788 0 net9
rlabel metal3 40032 2436 40032 2436 0 net90
rlabel metal3 41088 2142 41088 2142 0 net91
rlabel metal3 41472 2058 41472 2058 0 net92
rlabel metal3 41856 2016 41856 2016 0 net93
rlabel metal3 42240 1974 42240 1974 0 net94
rlabel metal4 17136 1512 17136 1512 0 net95
rlabel metal2 37632 1848 37632 1848 0 net96
rlabel metal3 37632 2184 37632 2184 0 net97
rlabel metal2 38016 1974 38016 1974 0 net98
rlabel metal2 22872 3612 22872 3612 0 net99
<< properties >>
string FIXED_BBOX 0 0 53280 12180
<< end >>
