VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO N_IO
  CLASS BLOCK ;
  FOREIGN N_IO ;
  ORIGIN 0.000 0.000 ;
  SIZE 231.840 BY 60.900 ;
  PIN A_I_top
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 23.320 60.500 23.720 60.900 ;
    END
  END A_I_top
  PIN A_O_top
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 17.560 60.500 17.960 60.900 ;
    END
  END A_O_top
  PIN A_T_top
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 29.080 60.500 29.480 60.900 ;
    END
  END A_T_top
  PIN A_config_C_bit0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 52.120 60.500 52.520 60.900 ;
    END
  END A_config_C_bit0
  PIN A_config_C_bit1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 57.880 60.500 58.280 60.900 ;
    END
  END A_config_C_bit1
  PIN A_config_C_bit2
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 63.640 60.500 64.040 60.900 ;
    END
  END A_config_C_bit2
  PIN A_config_C_bit3
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 69.400 60.500 69.800 60.900 ;
    END
  END A_config_C_bit3
  PIN B_I_top
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 40.600 60.500 41.000 60.900 ;
    END
  END B_I_top
  PIN B_O_top
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 34.840 60.500 35.240 60.900 ;
    END
  END B_O_top
  PIN B_T_top
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 46.360 60.500 46.760 60.900 ;
    END
  END B_T_top
  PIN B_config_C_bit0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 75.160 60.500 75.560 60.900 ;
    END
  END B_config_C_bit0
  PIN B_config_C_bit1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 80.920 60.500 81.320 60.900 ;
    END
  END B_config_C_bit1
  PIN B_config_C_bit2
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 86.680 60.500 87.080 60.900 ;
    END
  END B_config_C_bit2
  PIN B_config_C_bit3
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 92.440 60.500 92.840 60.900 ;
    END
  END B_config_C_bit3
  PIN Ci
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 104.920 0.000 105.320 0.400 ;
    END
  END Ci
  PIN FrameData[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 3.580 0.450 3.980 ;
    END
  END FrameData[0]
  PIN FrameData[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 20.380 0.450 20.780 ;
    END
  END FrameData[10]
  PIN FrameData[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 22.060 0.450 22.460 ;
    END
  END FrameData[11]
  PIN FrameData[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 23.740 0.450 24.140 ;
    END
  END FrameData[12]
  PIN FrameData[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 25.420 0.450 25.820 ;
    END
  END FrameData[13]
  PIN FrameData[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 27.100 0.450 27.500 ;
    END
  END FrameData[14]
  PIN FrameData[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 28.780 0.450 29.180 ;
    END
  END FrameData[15]
  PIN FrameData[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 30.460 0.450 30.860 ;
    END
  END FrameData[16]
  PIN FrameData[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 32.140 0.450 32.540 ;
    END
  END FrameData[17]
  PIN FrameData[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 33.820 0.450 34.220 ;
    END
  END FrameData[18]
  PIN FrameData[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 35.500 0.450 35.900 ;
    END
  END FrameData[19]
  PIN FrameData[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 5.260 0.450 5.660 ;
    END
  END FrameData[1]
  PIN FrameData[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 37.180 0.450 37.580 ;
    END
  END FrameData[20]
  PIN FrameData[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 38.860 0.450 39.260 ;
    END
  END FrameData[21]
  PIN FrameData[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 40.540 0.450 40.940 ;
    END
  END FrameData[22]
  PIN FrameData[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 42.220 0.450 42.620 ;
    END
  END FrameData[23]
  PIN FrameData[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 43.900 0.450 44.300 ;
    END
  END FrameData[24]
  PIN FrameData[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 45.580 0.450 45.980 ;
    END
  END FrameData[25]
  PIN FrameData[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 47.260 0.450 47.660 ;
    END
  END FrameData[26]
  PIN FrameData[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 48.940 0.450 49.340 ;
    END
  END FrameData[27]
  PIN FrameData[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 50.620 0.450 51.020 ;
    END
  END FrameData[28]
  PIN FrameData[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 52.300 0.450 52.700 ;
    END
  END FrameData[29]
  PIN FrameData[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 6.940 0.450 7.340 ;
    END
  END FrameData[2]
  PIN FrameData[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 53.980 0.450 54.380 ;
    END
  END FrameData[30]
  PIN FrameData[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 55.660 0.450 56.060 ;
    END
  END FrameData[31]
  PIN FrameData[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 8.620 0.450 9.020 ;
    END
  END FrameData[3]
  PIN FrameData[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 10.300 0.450 10.700 ;
    END
  END FrameData[4]
  PIN FrameData[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 11.980 0.450 12.380 ;
    END
  END FrameData[5]
  PIN FrameData[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 13.660 0.450 14.060 ;
    END
  END FrameData[6]
  PIN FrameData[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 15.340 0.450 15.740 ;
    END
  END FrameData[7]
  PIN FrameData[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 17.020 0.450 17.420 ;
    END
  END FrameData[8]
  PIN FrameData[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 18.700 0.450 19.100 ;
    END
  END FrameData[9]
  PIN FrameData_O[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 231.390 3.580 231.840 3.980 ;
    END
  END FrameData_O[0]
  PIN FrameData_O[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 231.390 20.380 231.840 20.780 ;
    END
  END FrameData_O[10]
  PIN FrameData_O[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 231.390 22.060 231.840 22.460 ;
    END
  END FrameData_O[11]
  PIN FrameData_O[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 231.390 23.740 231.840 24.140 ;
    END
  END FrameData_O[12]
  PIN FrameData_O[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 231.390 25.420 231.840 25.820 ;
    END
  END FrameData_O[13]
  PIN FrameData_O[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 231.390 27.100 231.840 27.500 ;
    END
  END FrameData_O[14]
  PIN FrameData_O[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 231.390 28.780 231.840 29.180 ;
    END
  END FrameData_O[15]
  PIN FrameData_O[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 231.390 30.460 231.840 30.860 ;
    END
  END FrameData_O[16]
  PIN FrameData_O[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 231.390 32.140 231.840 32.540 ;
    END
  END FrameData_O[17]
  PIN FrameData_O[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 231.390 33.820 231.840 34.220 ;
    END
  END FrameData_O[18]
  PIN FrameData_O[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 231.390 35.500 231.840 35.900 ;
    END
  END FrameData_O[19]
  PIN FrameData_O[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 231.390 5.260 231.840 5.660 ;
    END
  END FrameData_O[1]
  PIN FrameData_O[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 231.390 37.180 231.840 37.580 ;
    END
  END FrameData_O[20]
  PIN FrameData_O[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 231.390 38.860 231.840 39.260 ;
    END
  END FrameData_O[21]
  PIN FrameData_O[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 231.390 40.540 231.840 40.940 ;
    END
  END FrameData_O[22]
  PIN FrameData_O[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 231.390 42.220 231.840 42.620 ;
    END
  END FrameData_O[23]
  PIN FrameData_O[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 231.390 43.900 231.840 44.300 ;
    END
  END FrameData_O[24]
  PIN FrameData_O[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 231.390 45.580 231.840 45.980 ;
    END
  END FrameData_O[25]
  PIN FrameData_O[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 231.390 47.260 231.840 47.660 ;
    END
  END FrameData_O[26]
  PIN FrameData_O[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 231.390 48.940 231.840 49.340 ;
    END
  END FrameData_O[27]
  PIN FrameData_O[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 231.390 50.620 231.840 51.020 ;
    END
  END FrameData_O[28]
  PIN FrameData_O[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 231.390 52.300 231.840 52.700 ;
    END
  END FrameData_O[29]
  PIN FrameData_O[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 231.390 6.940 231.840 7.340 ;
    END
  END FrameData_O[2]
  PIN FrameData_O[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 231.390 53.980 231.840 54.380 ;
    END
  END FrameData_O[30]
  PIN FrameData_O[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 231.390 55.660 231.840 56.060 ;
    END
  END FrameData_O[31]
  PIN FrameData_O[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 231.390 8.620 231.840 9.020 ;
    END
  END FrameData_O[3]
  PIN FrameData_O[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 231.390 10.300 231.840 10.700 ;
    END
  END FrameData_O[4]
  PIN FrameData_O[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 231.390 11.980 231.840 12.380 ;
    END
  END FrameData_O[5]
  PIN FrameData_O[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 231.390 13.660 231.840 14.060 ;
    END
  END FrameData_O[6]
  PIN FrameData_O[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 231.390 15.340 231.840 15.740 ;
    END
  END FrameData_O[7]
  PIN FrameData_O[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 231.390 17.020 231.840 17.420 ;
    END
  END FrameData_O[8]
  PIN FrameData_O[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 231.390 18.700 231.840 19.100 ;
    END
  END FrameData_O[9]
  PIN FrameStrobe[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.542100 ;
    PORT
      LAYER Metal3 ;
        RECT 156.760 0.000 157.160 0.400 ;
    END
  END FrameStrobe[0]
  PIN FrameStrobe[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 166.360 0.000 166.760 0.400 ;
    END
  END FrameStrobe[10]
  PIN FrameStrobe[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 167.320 0.000 167.720 0.400 ;
    END
  END FrameStrobe[11]
  PIN FrameStrobe[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 168.280 0.000 168.680 0.400 ;
    END
  END FrameStrobe[12]
  PIN FrameStrobe[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 169.240 0.000 169.640 0.400 ;
    END
  END FrameStrobe[13]
  PIN FrameStrobe[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 170.200 0.000 170.600 0.400 ;
    END
  END FrameStrobe[14]
  PIN FrameStrobe[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 171.160 0.000 171.560 0.400 ;
    END
  END FrameStrobe[15]
  PIN FrameStrobe[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 172.120 0.000 172.520 0.400 ;
    END
  END FrameStrobe[16]
  PIN FrameStrobe[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 173.080 0.000 173.480 0.400 ;
    END
  END FrameStrobe[17]
  PIN FrameStrobe[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 174.040 0.000 174.440 0.400 ;
    END
  END FrameStrobe[18]
  PIN FrameStrobe[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 175.000 0.000 175.400 0.400 ;
    END
  END FrameStrobe[19]
  PIN FrameStrobe[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 157.720 0.000 158.120 0.400 ;
    END
  END FrameStrobe[1]
  PIN FrameStrobe[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.361400 ;
    PORT
      LAYER Metal3 ;
        RECT 158.680 0.000 159.080 0.400 ;
    END
  END FrameStrobe[2]
  PIN FrameStrobe[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 159.640 0.000 160.040 0.400 ;
    END
  END FrameStrobe[3]
  PIN FrameStrobe[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 160.600 0.000 161.000 0.400 ;
    END
  END FrameStrobe[4]
  PIN FrameStrobe[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 161.560 0.000 161.960 0.400 ;
    END
  END FrameStrobe[5]
  PIN FrameStrobe[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 162.520 0.000 162.920 0.400 ;
    END
  END FrameStrobe[6]
  PIN FrameStrobe[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 163.480 0.000 163.880 0.400 ;
    END
  END FrameStrobe[7]
  PIN FrameStrobe[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 164.440 0.000 164.840 0.400 ;
    END
  END FrameStrobe[8]
  PIN FrameStrobe[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 165.400 0.000 165.800 0.400 ;
    END
  END FrameStrobe[9]
  PIN FrameStrobe_O[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 103.960 60.500 104.360 60.900 ;
    END
  END FrameStrobe_O[0]
  PIN FrameStrobe_O[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 161.560 60.500 161.960 60.900 ;
    END
  END FrameStrobe_O[10]
  PIN FrameStrobe_O[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 167.320 60.500 167.720 60.900 ;
    END
  END FrameStrobe_O[11]
  PIN FrameStrobe_O[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 173.080 60.500 173.480 60.900 ;
    END
  END FrameStrobe_O[12]
  PIN FrameStrobe_O[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 178.840 60.500 179.240 60.900 ;
    END
  END FrameStrobe_O[13]
  PIN FrameStrobe_O[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 184.600 60.500 185.000 60.900 ;
    END
  END FrameStrobe_O[14]
  PIN FrameStrobe_O[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 190.360 60.500 190.760 60.900 ;
    END
  END FrameStrobe_O[15]
  PIN FrameStrobe_O[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 196.120 60.500 196.520 60.900 ;
    END
  END FrameStrobe_O[16]
  PIN FrameStrobe_O[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 201.880 60.500 202.280 60.900 ;
    END
  END FrameStrobe_O[17]
  PIN FrameStrobe_O[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 207.640 60.500 208.040 60.900 ;
    END
  END FrameStrobe_O[18]
  PIN FrameStrobe_O[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 213.400 60.500 213.800 60.900 ;
    END
  END FrameStrobe_O[19]
  PIN FrameStrobe_O[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 109.720 60.500 110.120 60.900 ;
    END
  END FrameStrobe_O[1]
  PIN FrameStrobe_O[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 115.480 60.500 115.880 60.900 ;
    END
  END FrameStrobe_O[2]
  PIN FrameStrobe_O[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 121.240 60.500 121.640 60.900 ;
    END
  END FrameStrobe_O[3]
  PIN FrameStrobe_O[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 127.000 60.500 127.400 60.900 ;
    END
  END FrameStrobe_O[4]
  PIN FrameStrobe_O[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 132.760 60.500 133.160 60.900 ;
    END
  END FrameStrobe_O[5]
  PIN FrameStrobe_O[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 138.520 60.500 138.920 60.900 ;
    END
  END FrameStrobe_O[6]
  PIN FrameStrobe_O[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 144.280 60.500 144.680 60.900 ;
    END
  END FrameStrobe_O[7]
  PIN FrameStrobe_O[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 150.040 60.500 150.440 60.900 ;
    END
  END FrameStrobe_O[8]
  PIN FrameStrobe_O[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 155.800 60.500 156.200 60.900 ;
    END
  END FrameStrobe_O[9]
  PIN N1END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 55.000 0.000 55.400 0.400 ;
    END
  END N1END[0]
  PIN N1END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 55.960 0.000 56.360 0.400 ;
    END
  END N1END[1]
  PIN N1END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 56.920 0.000 57.320 0.400 ;
    END
  END N1END[2]
  PIN N1END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 57.880 0.000 58.280 0.400 ;
    END
  END N1END[3]
  PIN N2END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 66.520 0.000 66.920 0.400 ;
    END
  END N2END[0]
  PIN N2END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 67.480 0.000 67.880 0.400 ;
    END
  END N2END[1]
  PIN N2END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 68.440 0.000 68.840 0.400 ;
    END
  END N2END[2]
  PIN N2END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 69.400 0.000 69.800 0.400 ;
    END
  END N2END[3]
  PIN N2END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 70.360 0.000 70.760 0.400 ;
    END
  END N2END[4]
  PIN N2END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 71.320 0.000 71.720 0.400 ;
    END
  END N2END[5]
  PIN N2END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 72.280 0.000 72.680 0.400 ;
    END
  END N2END[6]
  PIN N2END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 73.240 0.000 73.640 0.400 ;
    END
  END N2END[7]
  PIN N2MID[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 58.840 0.000 59.240 0.400 ;
    END
  END N2MID[0]
  PIN N2MID[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 59.800 0.000 60.200 0.400 ;
    END
  END N2MID[1]
  PIN N2MID[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 60.760 0.000 61.160 0.400 ;
    END
  END N2MID[2]
  PIN N2MID[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 61.720 0.000 62.120 0.400 ;
    END
  END N2MID[3]
  PIN N2MID[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 62.680 0.000 63.080 0.400 ;
    END
  END N2MID[4]
  PIN N2MID[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 63.640 0.000 64.040 0.400 ;
    END
  END N2MID[5]
  PIN N2MID[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 64.600 0.000 65.000 0.400 ;
    END
  END N2MID[6]
  PIN N2MID[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 65.560 0.000 65.960 0.400 ;
    END
  END N2MID[7]
  PIN N4END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 74.200 0.000 74.600 0.400 ;
    END
  END N4END[0]
  PIN N4END[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 83.800 0.000 84.200 0.400 ;
    END
  END N4END[10]
  PIN N4END[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 84.760 0.000 85.160 0.400 ;
    END
  END N4END[11]
  PIN N4END[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 85.720 0.000 86.120 0.400 ;
    END
  END N4END[12]
  PIN N4END[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 86.680 0.000 87.080 0.400 ;
    END
  END N4END[13]
  PIN N4END[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 87.640 0.000 88.040 0.400 ;
    END
  END N4END[14]
  PIN N4END[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 88.600 0.000 89.000 0.400 ;
    END
  END N4END[15]
  PIN N4END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 75.160 0.000 75.560 0.400 ;
    END
  END N4END[1]
  PIN N4END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 76.120 0.000 76.520 0.400 ;
    END
  END N4END[2]
  PIN N4END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 77.080 0.000 77.480 0.400 ;
    END
  END N4END[3]
  PIN N4END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 78.040 0.000 78.440 0.400 ;
    END
  END N4END[4]
  PIN N4END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 79.000 0.000 79.400 0.400 ;
    END
  END N4END[5]
  PIN N4END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 79.960 0.000 80.360 0.400 ;
    END
  END N4END[6]
  PIN N4END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 80.920 0.000 81.320 0.400 ;
    END
  END N4END[7]
  PIN N4END[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 81.880 0.000 82.280 0.400 ;
    END
  END N4END[8]
  PIN N4END[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 82.840 0.000 83.240 0.400 ;
    END
  END N4END[9]
  PIN NN4END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 89.560 0.000 89.960 0.400 ;
    END
  END NN4END[0]
  PIN NN4END[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 99.160 0.000 99.560 0.400 ;
    END
  END NN4END[10]
  PIN NN4END[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 100.120 0.000 100.520 0.400 ;
    END
  END NN4END[11]
  PIN NN4END[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 101.080 0.000 101.480 0.400 ;
    END
  END NN4END[12]
  PIN NN4END[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 102.040 0.000 102.440 0.400 ;
    END
  END NN4END[13]
  PIN NN4END[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 103.000 0.000 103.400 0.400 ;
    END
  END NN4END[14]
  PIN NN4END[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 103.960 0.000 104.360 0.400 ;
    END
  END NN4END[15]
  PIN NN4END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 90.520 0.000 90.920 0.400 ;
    END
  END NN4END[1]
  PIN NN4END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 91.480 0.000 91.880 0.400 ;
    END
  END NN4END[2]
  PIN NN4END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 92.440 0.000 92.840 0.400 ;
    END
  END NN4END[3]
  PIN NN4END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 93.400 0.000 93.800 0.400 ;
    END
  END NN4END[4]
  PIN NN4END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 94.360 0.000 94.760 0.400 ;
    END
  END NN4END[5]
  PIN NN4END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 95.320 0.000 95.720 0.400 ;
    END
  END NN4END[6]
  PIN NN4END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 96.280 0.000 96.680 0.400 ;
    END
  END NN4END[7]
  PIN NN4END[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 97.240 0.000 97.640 0.400 ;
    END
  END NN4END[8]
  PIN NN4END[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 98.200 0.000 98.600 0.400 ;
    END
  END NN4END[9]
  PIN S1BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 105.880 0.000 106.280 0.400 ;
    END
  END S1BEG[0]
  PIN S1BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 106.840 0.000 107.240 0.400 ;
    END
  END S1BEG[1]
  PIN S1BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 107.800 0.000 108.200 0.400 ;
    END
  END S1BEG[2]
  PIN S1BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 108.760 0.000 109.160 0.400 ;
    END
  END S1BEG[3]
  PIN S2BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 109.720 0.000 110.120 0.400 ;
    END
  END S2BEG[0]
  PIN S2BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 110.680 0.000 111.080 0.400 ;
    END
  END S2BEG[1]
  PIN S2BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 111.640 0.000 112.040 0.400 ;
    END
  END S2BEG[2]
  PIN S2BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 112.600 0.000 113.000 0.400 ;
    END
  END S2BEG[3]
  PIN S2BEG[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 113.560 0.000 113.960 0.400 ;
    END
  END S2BEG[4]
  PIN S2BEG[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 114.520 0.000 114.920 0.400 ;
    END
  END S2BEG[5]
  PIN S2BEG[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 115.480 0.000 115.880 0.400 ;
    END
  END S2BEG[6]
  PIN S2BEG[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 116.440 0.000 116.840 0.400 ;
    END
  END S2BEG[7]
  PIN S2BEGb[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 117.400 0.000 117.800 0.400 ;
    END
  END S2BEGb[0]
  PIN S2BEGb[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 118.360 0.000 118.760 0.400 ;
    END
  END S2BEGb[1]
  PIN S2BEGb[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 119.320 0.000 119.720 0.400 ;
    END
  END S2BEGb[2]
  PIN S2BEGb[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 120.280 0.000 120.680 0.400 ;
    END
  END S2BEGb[3]
  PIN S2BEGb[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 121.240 0.000 121.640 0.400 ;
    END
  END S2BEGb[4]
  PIN S2BEGb[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 122.200 0.000 122.600 0.400 ;
    END
  END S2BEGb[5]
  PIN S2BEGb[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 123.160 0.000 123.560 0.400 ;
    END
  END S2BEGb[6]
  PIN S2BEGb[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 124.120 0.000 124.520 0.400 ;
    END
  END S2BEGb[7]
  PIN S4BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 125.080 0.000 125.480 0.400 ;
    END
  END S4BEG[0]
  PIN S4BEG[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 134.680 0.000 135.080 0.400 ;
    END
  END S4BEG[10]
  PIN S4BEG[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 135.640 0.000 136.040 0.400 ;
    END
  END S4BEG[11]
  PIN S4BEG[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 136.600 0.000 137.000 0.400 ;
    END
  END S4BEG[12]
  PIN S4BEG[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 137.560 0.000 137.960 0.400 ;
    END
  END S4BEG[13]
  PIN S4BEG[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 138.520 0.000 138.920 0.400 ;
    END
  END S4BEG[14]
  PIN S4BEG[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 139.480 0.000 139.880 0.400 ;
    END
  END S4BEG[15]
  PIN S4BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 126.040 0.000 126.440 0.400 ;
    END
  END S4BEG[1]
  PIN S4BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 127.000 0.000 127.400 0.400 ;
    END
  END S4BEG[2]
  PIN S4BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 127.960 0.000 128.360 0.400 ;
    END
  END S4BEG[3]
  PIN S4BEG[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 128.920 0.000 129.320 0.400 ;
    END
  END S4BEG[4]
  PIN S4BEG[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 129.880 0.000 130.280 0.400 ;
    END
  END S4BEG[5]
  PIN S4BEG[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 130.840 0.000 131.240 0.400 ;
    END
  END S4BEG[6]
  PIN S4BEG[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 131.800 0.000 132.200 0.400 ;
    END
  END S4BEG[7]
  PIN S4BEG[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 132.760 0.000 133.160 0.400 ;
    END
  END S4BEG[8]
  PIN S4BEG[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 133.720 0.000 134.120 0.400 ;
    END
  END S4BEG[9]
  PIN SS4BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 140.440 0.000 140.840 0.400 ;
    END
  END SS4BEG[0]
  PIN SS4BEG[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 150.040 0.000 150.440 0.400 ;
    END
  END SS4BEG[10]
  PIN SS4BEG[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 151.000 0.000 151.400 0.400 ;
    END
  END SS4BEG[11]
  PIN SS4BEG[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 151.960 0.000 152.360 0.400 ;
    END
  END SS4BEG[12]
  PIN SS4BEG[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 152.920 0.000 153.320 0.400 ;
    END
  END SS4BEG[13]
  PIN SS4BEG[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 153.880 0.000 154.280 0.400 ;
    END
  END SS4BEG[14]
  PIN SS4BEG[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 154.840 0.000 155.240 0.400 ;
    END
  END SS4BEG[15]
  PIN SS4BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 141.400 0.000 141.800 0.400 ;
    END
  END SS4BEG[1]
  PIN SS4BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 142.360 0.000 142.760 0.400 ;
    END
  END SS4BEG[2]
  PIN SS4BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 143.320 0.000 143.720 0.400 ;
    END
  END SS4BEG[3]
  PIN SS4BEG[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 144.280 0.000 144.680 0.400 ;
    END
  END SS4BEG[4]
  PIN SS4BEG[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 145.240 0.000 145.640 0.400 ;
    END
  END SS4BEG[5]
  PIN SS4BEG[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 146.200 0.000 146.600 0.400 ;
    END
  END SS4BEG[6]
  PIN SS4BEG[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 147.160 0.000 147.560 0.400 ;
    END
  END SS4BEG[7]
  PIN SS4BEG[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 148.120 0.000 148.520 0.400 ;
    END
  END SS4BEG[8]
  PIN SS4BEG[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 149.080 0.000 149.480 0.400 ;
    END
  END SS4BEG[9]
  PIN UserCLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.633100 ;
    PORT
      LAYER Metal3 ;
        RECT 155.800 0.000 156.200 0.400 ;
    END
  END UserCLK
  PIN UserCLKo
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 98.200 60.500 98.600 60.900 ;
    END
  END UserCLKo
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal5 ;
        RECT 24.460 0.000 26.660 60.900 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 100.060 0.000 102.260 60.900 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 175.660 0.000 177.860 60.900 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal5 ;
        RECT 18.260 0.000 20.460 60.900 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 93.860 0.000 96.060 60.900 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 169.460 0.000 171.660 60.900 ;
    END
  END VPWR
  OBS
      LAYER GatPoly ;
        RECT 5.760 7.410 226.080 53.070 ;
      LAYER Metal1 ;
        RECT 5.760 7.340 226.080 53.140 ;
      LAYER Metal2 ;
        RECT 0.335 56.270 231.505 58.480 ;
        RECT 0.660 55.450 231.180 56.270 ;
        RECT 0.335 54.590 231.505 55.450 ;
        RECT 0.660 53.770 231.180 54.590 ;
        RECT 0.335 52.910 231.505 53.770 ;
        RECT 0.660 52.090 231.180 52.910 ;
        RECT 0.335 51.230 231.505 52.090 ;
        RECT 0.660 50.410 231.180 51.230 ;
        RECT 0.335 49.550 231.505 50.410 ;
        RECT 0.660 48.730 231.180 49.550 ;
        RECT 0.335 47.870 231.505 48.730 ;
        RECT 0.660 47.050 231.180 47.870 ;
        RECT 0.335 46.190 231.505 47.050 ;
        RECT 0.660 45.370 231.180 46.190 ;
        RECT 0.335 44.510 231.505 45.370 ;
        RECT 0.660 43.690 231.180 44.510 ;
        RECT 0.335 42.830 231.505 43.690 ;
        RECT 0.660 42.010 231.180 42.830 ;
        RECT 0.335 41.150 231.505 42.010 ;
        RECT 0.660 40.330 231.180 41.150 ;
        RECT 0.335 39.470 231.505 40.330 ;
        RECT 0.660 38.650 231.180 39.470 ;
        RECT 0.335 37.790 231.505 38.650 ;
        RECT 0.660 36.970 231.180 37.790 ;
        RECT 0.335 36.110 231.505 36.970 ;
        RECT 0.660 35.290 231.180 36.110 ;
        RECT 0.335 34.430 231.505 35.290 ;
        RECT 0.660 33.610 231.180 34.430 ;
        RECT 0.335 32.750 231.505 33.610 ;
        RECT 0.660 31.930 231.180 32.750 ;
        RECT 0.335 31.070 231.505 31.930 ;
        RECT 0.660 30.250 231.180 31.070 ;
        RECT 0.335 29.390 231.505 30.250 ;
        RECT 0.660 28.570 231.180 29.390 ;
        RECT 0.335 27.710 231.505 28.570 ;
        RECT 0.660 26.890 231.180 27.710 ;
        RECT 0.335 26.030 231.505 26.890 ;
        RECT 0.660 25.210 231.180 26.030 ;
        RECT 0.335 24.350 231.505 25.210 ;
        RECT 0.660 23.530 231.180 24.350 ;
        RECT 0.335 22.670 231.505 23.530 ;
        RECT 0.660 21.850 231.180 22.670 ;
        RECT 0.335 20.990 231.505 21.850 ;
        RECT 0.660 20.170 231.180 20.990 ;
        RECT 0.335 19.310 231.505 20.170 ;
        RECT 0.660 18.490 231.180 19.310 ;
        RECT 0.335 17.630 231.505 18.490 ;
        RECT 0.660 16.810 231.180 17.630 ;
        RECT 0.335 15.950 231.505 16.810 ;
        RECT 0.660 15.130 231.180 15.950 ;
        RECT 0.335 14.270 231.505 15.130 ;
        RECT 0.660 13.450 231.180 14.270 ;
        RECT 0.335 12.590 231.505 13.450 ;
        RECT 0.660 11.770 231.180 12.590 ;
        RECT 0.335 10.910 231.505 11.770 ;
        RECT 0.660 10.090 231.180 10.910 ;
        RECT 0.335 9.230 231.505 10.090 ;
        RECT 0.660 8.410 231.180 9.230 ;
        RECT 0.335 7.550 231.505 8.410 ;
        RECT 0.660 6.730 231.180 7.550 ;
        RECT 0.335 5.870 231.505 6.730 ;
        RECT 0.660 5.050 231.180 5.870 ;
        RECT 0.335 4.190 231.505 5.050 ;
        RECT 0.660 3.370 231.180 4.190 ;
        RECT 0.335 0.320 231.505 3.370 ;
      LAYER Metal3 ;
        RECT 0.380 60.290 17.350 60.500 ;
        RECT 18.170 60.290 23.110 60.500 ;
        RECT 23.930 60.290 28.870 60.500 ;
        RECT 29.690 60.290 34.630 60.500 ;
        RECT 35.450 60.290 40.390 60.500 ;
        RECT 41.210 60.290 46.150 60.500 ;
        RECT 46.970 60.290 51.910 60.500 ;
        RECT 52.730 60.290 57.670 60.500 ;
        RECT 58.490 60.290 63.430 60.500 ;
        RECT 64.250 60.290 69.190 60.500 ;
        RECT 70.010 60.290 74.950 60.500 ;
        RECT 75.770 60.290 80.710 60.500 ;
        RECT 81.530 60.290 86.470 60.500 ;
        RECT 87.290 60.290 92.230 60.500 ;
        RECT 93.050 60.290 97.990 60.500 ;
        RECT 98.810 60.290 103.750 60.500 ;
        RECT 104.570 60.290 109.510 60.500 ;
        RECT 110.330 60.290 115.270 60.500 ;
        RECT 116.090 60.290 121.030 60.500 ;
        RECT 121.850 60.290 126.790 60.500 ;
        RECT 127.610 60.290 132.550 60.500 ;
        RECT 133.370 60.290 138.310 60.500 ;
        RECT 139.130 60.290 144.070 60.500 ;
        RECT 144.890 60.290 149.830 60.500 ;
        RECT 150.650 60.290 155.590 60.500 ;
        RECT 156.410 60.290 161.350 60.500 ;
        RECT 162.170 60.290 167.110 60.500 ;
        RECT 167.930 60.290 172.870 60.500 ;
        RECT 173.690 60.290 178.630 60.500 ;
        RECT 179.450 60.290 184.390 60.500 ;
        RECT 185.210 60.290 190.150 60.500 ;
        RECT 190.970 60.290 195.910 60.500 ;
        RECT 196.730 60.290 201.670 60.500 ;
        RECT 202.490 60.290 207.430 60.500 ;
        RECT 208.250 60.290 213.190 60.500 ;
        RECT 214.010 60.290 231.460 60.500 ;
        RECT 0.380 0.610 231.460 60.290 ;
        RECT 0.380 0.180 54.790 0.610 ;
        RECT 55.610 0.180 55.750 0.610 ;
        RECT 56.570 0.180 56.710 0.610 ;
        RECT 57.530 0.180 57.670 0.610 ;
        RECT 58.490 0.180 58.630 0.610 ;
        RECT 59.450 0.180 59.590 0.610 ;
        RECT 60.410 0.180 60.550 0.610 ;
        RECT 61.370 0.180 61.510 0.610 ;
        RECT 62.330 0.180 62.470 0.610 ;
        RECT 63.290 0.180 63.430 0.610 ;
        RECT 64.250 0.180 64.390 0.610 ;
        RECT 65.210 0.180 65.350 0.610 ;
        RECT 66.170 0.180 66.310 0.610 ;
        RECT 67.130 0.180 67.270 0.610 ;
        RECT 68.090 0.180 68.230 0.610 ;
        RECT 69.050 0.180 69.190 0.610 ;
        RECT 70.010 0.180 70.150 0.610 ;
        RECT 70.970 0.180 71.110 0.610 ;
        RECT 71.930 0.180 72.070 0.610 ;
        RECT 72.890 0.180 73.030 0.610 ;
        RECT 73.850 0.180 73.990 0.610 ;
        RECT 74.810 0.180 74.950 0.610 ;
        RECT 75.770 0.180 75.910 0.610 ;
        RECT 76.730 0.180 76.870 0.610 ;
        RECT 77.690 0.180 77.830 0.610 ;
        RECT 78.650 0.180 78.790 0.610 ;
        RECT 79.610 0.180 79.750 0.610 ;
        RECT 80.570 0.180 80.710 0.610 ;
        RECT 81.530 0.180 81.670 0.610 ;
        RECT 82.490 0.180 82.630 0.610 ;
        RECT 83.450 0.180 83.590 0.610 ;
        RECT 84.410 0.180 84.550 0.610 ;
        RECT 85.370 0.180 85.510 0.610 ;
        RECT 86.330 0.180 86.470 0.610 ;
        RECT 87.290 0.180 87.430 0.610 ;
        RECT 88.250 0.180 88.390 0.610 ;
        RECT 89.210 0.180 89.350 0.610 ;
        RECT 90.170 0.180 90.310 0.610 ;
        RECT 91.130 0.180 91.270 0.610 ;
        RECT 92.090 0.180 92.230 0.610 ;
        RECT 93.050 0.180 93.190 0.610 ;
        RECT 94.010 0.180 94.150 0.610 ;
        RECT 94.970 0.180 95.110 0.610 ;
        RECT 95.930 0.180 96.070 0.610 ;
        RECT 96.890 0.180 97.030 0.610 ;
        RECT 97.850 0.180 97.990 0.610 ;
        RECT 98.810 0.180 98.950 0.610 ;
        RECT 99.770 0.180 99.910 0.610 ;
        RECT 100.730 0.180 100.870 0.610 ;
        RECT 101.690 0.180 101.830 0.610 ;
        RECT 102.650 0.180 102.790 0.610 ;
        RECT 103.610 0.180 103.750 0.610 ;
        RECT 104.570 0.180 104.710 0.610 ;
        RECT 105.530 0.180 105.670 0.610 ;
        RECT 106.490 0.180 106.630 0.610 ;
        RECT 107.450 0.180 107.590 0.610 ;
        RECT 108.410 0.180 108.550 0.610 ;
        RECT 109.370 0.180 109.510 0.610 ;
        RECT 110.330 0.180 110.470 0.610 ;
        RECT 111.290 0.180 111.430 0.610 ;
        RECT 112.250 0.180 112.390 0.610 ;
        RECT 113.210 0.180 113.350 0.610 ;
        RECT 114.170 0.180 114.310 0.610 ;
        RECT 115.130 0.180 115.270 0.610 ;
        RECT 116.090 0.180 116.230 0.610 ;
        RECT 117.050 0.180 117.190 0.610 ;
        RECT 118.010 0.180 118.150 0.610 ;
        RECT 118.970 0.180 119.110 0.610 ;
        RECT 119.930 0.180 120.070 0.610 ;
        RECT 120.890 0.180 121.030 0.610 ;
        RECT 121.850 0.180 121.990 0.610 ;
        RECT 122.810 0.180 122.950 0.610 ;
        RECT 123.770 0.180 123.910 0.610 ;
        RECT 124.730 0.180 124.870 0.610 ;
        RECT 125.690 0.180 125.830 0.610 ;
        RECT 126.650 0.180 126.790 0.610 ;
        RECT 127.610 0.180 127.750 0.610 ;
        RECT 128.570 0.180 128.710 0.610 ;
        RECT 129.530 0.180 129.670 0.610 ;
        RECT 130.490 0.180 130.630 0.610 ;
        RECT 131.450 0.180 131.590 0.610 ;
        RECT 132.410 0.180 132.550 0.610 ;
        RECT 133.370 0.180 133.510 0.610 ;
        RECT 134.330 0.180 134.470 0.610 ;
        RECT 135.290 0.180 135.430 0.610 ;
        RECT 136.250 0.180 136.390 0.610 ;
        RECT 137.210 0.180 137.350 0.610 ;
        RECT 138.170 0.180 138.310 0.610 ;
        RECT 139.130 0.180 139.270 0.610 ;
        RECT 140.090 0.180 140.230 0.610 ;
        RECT 141.050 0.180 141.190 0.610 ;
        RECT 142.010 0.180 142.150 0.610 ;
        RECT 142.970 0.180 143.110 0.610 ;
        RECT 143.930 0.180 144.070 0.610 ;
        RECT 144.890 0.180 145.030 0.610 ;
        RECT 145.850 0.180 145.990 0.610 ;
        RECT 146.810 0.180 146.950 0.610 ;
        RECT 147.770 0.180 147.910 0.610 ;
        RECT 148.730 0.180 148.870 0.610 ;
        RECT 149.690 0.180 149.830 0.610 ;
        RECT 150.650 0.180 150.790 0.610 ;
        RECT 151.610 0.180 151.750 0.610 ;
        RECT 152.570 0.180 152.710 0.610 ;
        RECT 153.530 0.180 153.670 0.610 ;
        RECT 154.490 0.180 154.630 0.610 ;
        RECT 155.450 0.180 155.590 0.610 ;
        RECT 156.410 0.180 156.550 0.610 ;
        RECT 157.370 0.180 157.510 0.610 ;
        RECT 158.330 0.180 158.470 0.610 ;
        RECT 159.290 0.180 159.430 0.610 ;
        RECT 160.250 0.180 160.390 0.610 ;
        RECT 161.210 0.180 161.350 0.610 ;
        RECT 162.170 0.180 162.310 0.610 ;
        RECT 163.130 0.180 163.270 0.610 ;
        RECT 164.090 0.180 164.230 0.610 ;
        RECT 165.050 0.180 165.190 0.610 ;
        RECT 166.010 0.180 166.150 0.610 ;
        RECT 166.970 0.180 167.110 0.610 ;
        RECT 167.930 0.180 168.070 0.610 ;
        RECT 168.890 0.180 169.030 0.610 ;
        RECT 169.850 0.180 169.990 0.610 ;
        RECT 170.810 0.180 170.950 0.610 ;
        RECT 171.770 0.180 171.910 0.610 ;
        RECT 172.730 0.180 172.870 0.610 ;
        RECT 173.690 0.180 173.830 0.610 ;
        RECT 174.650 0.180 174.790 0.610 ;
        RECT 175.610 0.180 231.460 0.610 ;
      LAYER Metal4 ;
        RECT 7.055 0.320 224.785 54.700 ;
      LAYER Metal5 ;
        RECT 72.380 6.575 93.650 47.185 ;
        RECT 96.270 6.575 99.850 47.185 ;
        RECT 102.470 6.575 169.250 47.185 ;
        RECT 171.870 6.575 173.380 47.185 ;
  END
END N_IO
END LIBRARY

