module S_term_single (Co,
    UserCLK,
    UserCLKo,
    VPWR,
    VGND,
    FrameData,
    FrameData_O,
    FrameStrobe,
    FrameStrobe_O,
    N1BEG,
    N2BEG,
    N2BEGb,
    N4BEG,
    NN4BEG,
    S1END,
    S2END,
    S2MID,
    S4END,
    SS4END);
 output Co;
 input UserCLK;
 output UserCLKo;
 inout VPWR;
 inout VGND;
 input [31:0] FrameData;
 output [31:0] FrameData_O;
 input [19:0] FrameStrobe;
 output [19:0] FrameStrobe_O;
 output [3:0] N1BEG;
 output [7:0] N2BEG;
 output [7:0] N2BEGb;
 output [15:0] N4BEG;
 output [15:0] NN4BEG;
 input [3:0] S1END;
 input [7:0] S2END;
 input [7:0] S2MID;
 input [15:0] S4END;
 input [15:0] SS4END;

 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;

 sg13g2_antennanp ANTENNA_1 (.VDD(VPWR),
    .VSS(VGND),
    .A(FrameData[16]));
 sg13g2_buf_1 _001_ (.A(FrameData[0]),
    .X(net1),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _002_ (.A(FrameData[1]),
    .X(net12),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _003_ (.A(FrameData[2]),
    .X(net23),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _004_ (.A(FrameData[3]),
    .X(net26),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _005_ (.A(FrameData[4]),
    .X(net27),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _006_ (.A(FrameData[5]),
    .X(net28),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _007_ (.A(FrameData[6]),
    .X(net29),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _008_ (.A(FrameData[7]),
    .X(net30),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _009_ (.A(FrameData[8]),
    .X(net31),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _010_ (.A(FrameData[9]),
    .X(net32),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _011_ (.A(FrameData[10]),
    .X(net2),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _012_ (.A(FrameData[11]),
    .X(net3),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _013_ (.A(FrameData[12]),
    .X(net4),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _014_ (.A(FrameData[13]),
    .X(net5),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _015_ (.A(FrameData[14]),
    .X(net6),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _016_ (.A(FrameData[15]),
    .X(net7),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _017_ (.A(FrameData[16]),
    .X(net8),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _018_ (.A(FrameData[17]),
    .X(net9),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _019_ (.A(FrameData[18]),
    .X(net10),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _020_ (.A(FrameData[19]),
    .X(net11),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _021_ (.A(FrameData[20]),
    .X(net13),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _022_ (.A(FrameData[21]),
    .X(net14),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _023_ (.A(FrameData[22]),
    .X(net15),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _024_ (.A(FrameData[23]),
    .X(net16),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _025_ (.A(FrameData[24]),
    .X(net17),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _026_ (.A(FrameData[25]),
    .X(net18),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _027_ (.A(FrameData[26]),
    .X(net19),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _028_ (.A(FrameData[27]),
    .X(net20),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _029_ (.A(FrameData[28]),
    .X(net21),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _030_ (.A(FrameData[29]),
    .X(net22),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _031_ (.A(FrameData[30]),
    .X(net24),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _032_ (.A(FrameData[31]),
    .X(net25),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _033_ (.A(FrameStrobe[0]),
    .X(net33),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _034_ (.A(FrameStrobe[1]),
    .X(net44),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _035_ (.A(FrameStrobe[2]),
    .X(net45),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _036_ (.A(FrameStrobe[3]),
    .X(net46),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _037_ (.A(FrameStrobe[4]),
    .X(net47),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _038_ (.A(FrameStrobe[5]),
    .X(net48),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _039_ (.A(FrameStrobe[6]),
    .X(net49),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _040_ (.A(FrameStrobe[7]),
    .X(net50),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _041_ (.A(FrameStrobe[8]),
    .X(net51),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _042_ (.A(FrameStrobe[9]),
    .X(net52),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _043_ (.A(FrameStrobe[10]),
    .X(net34),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _044_ (.A(FrameStrobe[11]),
    .X(net35),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _045_ (.A(FrameStrobe[12]),
    .X(net36),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _046_ (.A(FrameStrobe[13]),
    .X(net37),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _047_ (.A(FrameStrobe[14]),
    .X(net38),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _048_ (.A(FrameStrobe[15]),
    .X(net39),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _049_ (.A(FrameStrobe[16]),
    .X(net40),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _050_ (.A(FrameStrobe[17]),
    .X(net41),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _051_ (.A(FrameStrobe[18]),
    .X(net42),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _052_ (.A(FrameStrobe[19]),
    .X(net43),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _053_ (.A(S1END[3]),
    .X(net53),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _054_ (.A(S1END[2]),
    .X(net54),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _055_ (.A(S1END[1]),
    .X(net55),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _056_ (.A(S1END[0]),
    .X(net56),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _057_ (.A(S2MID[7]),
    .X(net57),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _058_ (.A(S2MID[6]),
    .X(net58),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _059_ (.A(S2MID[5]),
    .X(net59),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _060_ (.A(S2MID[4]),
    .X(net60),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _061_ (.A(S2MID[3]),
    .X(net61),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _062_ (.A(S2MID[2]),
    .X(net62),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _063_ (.A(S2MID[1]),
    .X(net63),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _064_ (.A(S2MID[0]),
    .X(net64),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _065_ (.A(S2END[7]),
    .X(net65),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _066_ (.A(S2END[6]),
    .X(net66),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _067_ (.A(S2END[5]),
    .X(net67),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _068_ (.A(S2END[4]),
    .X(net68),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _069_ (.A(S2END[3]),
    .X(net69),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _070_ (.A(S2END[2]),
    .X(net70),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _071_ (.A(S2END[1]),
    .X(net71),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _072_ (.A(S2END[0]),
    .X(net72),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _073_ (.A(S4END[15]),
    .X(net73),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _074_ (.A(S4END[14]),
    .X(net80),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _075_ (.A(S4END[13]),
    .X(net81),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _076_ (.A(S4END[12]),
    .X(net82),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _077_ (.A(S4END[11]),
    .X(net83),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _078_ (.A(S4END[10]),
    .X(net84),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _079_ (.A(S4END[9]),
    .X(net85),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _080_ (.A(S4END[8]),
    .X(net86),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _081_ (.A(S4END[7]),
    .X(net87),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _082_ (.A(S4END[6]),
    .X(net88),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _083_ (.A(S4END[5]),
    .X(net74),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _084_ (.A(S4END[4]),
    .X(net75),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _085_ (.A(S4END[3]),
    .X(net76),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _086_ (.A(S4END[2]),
    .X(net77),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _087_ (.A(S4END[1]),
    .X(net78),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _088_ (.A(S4END[0]),
    .X(net79),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _089_ (.A(SS4END[15]),
    .X(net89),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _090_ (.A(SS4END[14]),
    .X(net96),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _091_ (.A(SS4END[13]),
    .X(net97),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _092_ (.A(SS4END[12]),
    .X(net98),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _093_ (.A(SS4END[11]),
    .X(net99),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _094_ (.A(SS4END[10]),
    .X(net100),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _095_ (.A(SS4END[9]),
    .X(net101),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _096_ (.A(SS4END[8]),
    .X(net102),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _097_ (.A(SS4END[7]),
    .X(net103),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _098_ (.A(SS4END[6]),
    .X(net104),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _099_ (.A(SS4END[5]),
    .X(net90),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _100_ (.A(SS4END[4]),
    .X(net91),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _101_ (.A(SS4END[3]),
    .X(net92),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _102_ (.A(SS4END[2]),
    .X(net93),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _103_ (.A(SS4END[1]),
    .X(net94),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _104_ (.A(SS4END[0]),
    .X(net95),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _105_ (.A(UserCLK),
    .X(net105),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output1 (.A(net1),
    .X(FrameData_O[0]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output2 (.A(net2),
    .X(FrameData_O[10]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output3 (.A(net3),
    .X(FrameData_O[11]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output4 (.A(net4),
    .X(FrameData_O[12]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output5 (.A(net5),
    .X(FrameData_O[13]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output6 (.A(net6),
    .X(FrameData_O[14]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output7 (.A(net7),
    .X(FrameData_O[15]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output8 (.A(net8),
    .X(FrameData_O[16]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output9 (.A(net9),
    .X(FrameData_O[17]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output10 (.A(net10),
    .X(FrameData_O[18]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output11 (.A(net11),
    .X(FrameData_O[19]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output12 (.A(net12),
    .X(FrameData_O[1]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output13 (.A(net13),
    .X(FrameData_O[20]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output14 (.A(net14),
    .X(FrameData_O[21]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output15 (.A(net15),
    .X(FrameData_O[22]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output16 (.A(net16),
    .X(FrameData_O[23]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output17 (.A(net17),
    .X(FrameData_O[24]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output18 (.A(net18),
    .X(FrameData_O[25]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output19 (.A(net19),
    .X(FrameData_O[26]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output20 (.A(net20),
    .X(FrameData_O[27]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output21 (.A(net21),
    .X(FrameData_O[28]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output22 (.A(net22),
    .X(FrameData_O[29]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output23 (.A(net23),
    .X(FrameData_O[2]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output24 (.A(net24),
    .X(FrameData_O[30]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output25 (.A(net25),
    .X(FrameData_O[31]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output26 (.A(net26),
    .X(FrameData_O[3]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output27 (.A(net27),
    .X(FrameData_O[4]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output28 (.A(net28),
    .X(FrameData_O[5]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output29 (.A(net29),
    .X(FrameData_O[6]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output30 (.A(net30),
    .X(FrameData_O[7]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output31 (.A(net31),
    .X(FrameData_O[8]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output32 (.A(net32),
    .X(FrameData_O[9]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output33 (.A(net33),
    .X(FrameStrobe_O[0]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output34 (.A(net34),
    .X(FrameStrobe_O[10]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output35 (.A(net35),
    .X(FrameStrobe_O[11]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output36 (.A(net36),
    .X(FrameStrobe_O[12]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output37 (.A(net37),
    .X(FrameStrobe_O[13]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output38 (.A(net38),
    .X(FrameStrobe_O[14]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output39 (.A(net39),
    .X(FrameStrobe_O[15]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output40 (.A(net40),
    .X(FrameStrobe_O[16]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output41 (.A(net41),
    .X(FrameStrobe_O[17]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output42 (.A(net42),
    .X(FrameStrobe_O[18]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output43 (.A(net43),
    .X(FrameStrobe_O[19]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output44 (.A(net44),
    .X(FrameStrobe_O[1]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output45 (.A(net45),
    .X(FrameStrobe_O[2]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output46 (.A(net46),
    .X(FrameStrobe_O[3]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output47 (.A(net47),
    .X(FrameStrobe_O[4]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output48 (.A(net48),
    .X(FrameStrobe_O[5]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output49 (.A(net49),
    .X(FrameStrobe_O[6]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output50 (.A(net50),
    .X(FrameStrobe_O[7]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output51 (.A(net51),
    .X(FrameStrobe_O[8]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output52 (.A(net52),
    .X(FrameStrobe_O[9]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output53 (.A(net53),
    .X(N1BEG[0]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output54 (.A(net54),
    .X(N1BEG[1]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output55 (.A(net55),
    .X(N1BEG[2]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output56 (.A(net56),
    .X(N1BEG[3]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output57 (.A(net57),
    .X(N2BEG[0]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output58 (.A(net58),
    .X(N2BEG[1]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output59 (.A(net59),
    .X(N2BEG[2]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output60 (.A(net60),
    .X(N2BEG[3]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output61 (.A(net61),
    .X(N2BEG[4]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output62 (.A(net62),
    .X(N2BEG[5]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output63 (.A(net63),
    .X(N2BEG[6]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output64 (.A(net64),
    .X(N2BEG[7]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output65 (.A(net65),
    .X(N2BEGb[0]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output66 (.A(net66),
    .X(N2BEGb[1]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output67 (.A(net67),
    .X(N2BEGb[2]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output68 (.A(net68),
    .X(N2BEGb[3]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output69 (.A(net69),
    .X(N2BEGb[4]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output70 (.A(net70),
    .X(N2BEGb[5]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output71 (.A(net71),
    .X(N2BEGb[6]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output72 (.A(net72),
    .X(N2BEGb[7]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output73 (.A(net73),
    .X(N4BEG[0]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output74 (.A(net74),
    .X(N4BEG[10]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output75 (.A(net75),
    .X(N4BEG[11]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output76 (.A(net76),
    .X(N4BEG[12]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output77 (.A(net77),
    .X(N4BEG[13]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output78 (.A(net78),
    .X(N4BEG[14]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output79 (.A(net79),
    .X(N4BEG[15]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output80 (.A(net80),
    .X(N4BEG[1]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output81 (.A(net81),
    .X(N4BEG[2]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output82 (.A(net82),
    .X(N4BEG[3]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output83 (.A(net83),
    .X(N4BEG[4]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output84 (.A(net84),
    .X(N4BEG[5]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output85 (.A(net85),
    .X(N4BEG[6]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output86 (.A(net86),
    .X(N4BEG[7]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output87 (.A(net87),
    .X(N4BEG[8]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output88 (.A(net88),
    .X(N4BEG[9]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output89 (.A(net89),
    .X(NN4BEG[0]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output90 (.A(net90),
    .X(NN4BEG[10]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output91 (.A(net91),
    .X(NN4BEG[11]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output92 (.A(net92),
    .X(NN4BEG[12]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output93 (.A(net93),
    .X(NN4BEG[13]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output94 (.A(net94),
    .X(NN4BEG[14]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output95 (.A(net95),
    .X(NN4BEG[15]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output96 (.A(net96),
    .X(NN4BEG[1]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output97 (.A(net97),
    .X(NN4BEG[2]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output98 (.A(net98),
    .X(NN4BEG[3]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output99 (.A(net99),
    .X(NN4BEG[4]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output100 (.A(net100),
    .X(NN4BEG[5]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output101 (.A(net101),
    .X(NN4BEG[6]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output102 (.A(net102),
    .X(NN4BEG[7]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output103 (.A(net103),
    .X(NN4BEG[8]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output104 (.A(net104),
    .X(NN4BEG[9]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output105 (.A(net105),
    .X(UserCLKo),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_tielo S_term_single_106 (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(net106));
 sg13g2_antennanp ANTENNA_2 (.VDD(VPWR),
    .VSS(VGND),
    .A(FrameData[21]));
 sg13g2_antennanp ANTENNA_3 (.VDD(VPWR),
    .VSS(VGND),
    .A(FrameData[24]));
 sg13g2_antennanp ANTENNA_4 (.VDD(VPWR),
    .VSS(VGND),
    .A(FrameData[25]));
 sg13g2_antennanp ANTENNA_5 (.VDD(VPWR),
    .VSS(VGND),
    .A(FrameData[26]));
 sg13g2_antennanp ANTENNA_6 (.VDD(VPWR),
    .VSS(VGND),
    .A(FrameData[29]));
 sg13g2_antennanp ANTENNA_7 (.VDD(VPWR),
    .VSS(VGND),
    .A(FrameData[16]));
 sg13g2_antennanp ANTENNA_8 (.VDD(VPWR),
    .VSS(VGND),
    .A(FrameData[21]));
 sg13g2_antennanp ANTENNA_9 (.VDD(VPWR),
    .VSS(VGND),
    .A(FrameData[24]));
 sg13g2_antennanp ANTENNA_10 (.VDD(VPWR),
    .VSS(VGND),
    .A(FrameData[25]));
 sg13g2_antennanp ANTENNA_11 (.VDD(VPWR),
    .VSS(VGND),
    .A(FrameData[26]));
 sg13g2_antennanp ANTENNA_12 (.VDD(VPWR),
    .VSS(VGND),
    .A(FrameData[27]));
 sg13g2_antennanp ANTENNA_13 (.VDD(VPWR),
    .VSS(VGND),
    .A(FrameData[29]));
 sg13g2_antennanp ANTENNA_14 (.VDD(VPWR),
    .VSS(VGND),
    .A(FrameData[24]));
 sg13g2_antennanp ANTENNA_15 (.VDD(VPWR),
    .VSS(VGND),
    .A(FrameData[25]));
 sg13g2_antennanp ANTENNA_16 (.VDD(VPWR),
    .VSS(VGND),
    .A(FrameData[26]));
 sg13g2_antennanp ANTENNA_17 (.VDD(VPWR),
    .VSS(VGND),
    .A(FrameData[27]));
 sg13g2_antennanp ANTENNA_18 (.VDD(VPWR),
    .VSS(VGND),
    .A(FrameData[24]));
 sg13g2_antennanp ANTENNA_19 (.VDD(VPWR),
    .VSS(VGND),
    .A(FrameData[25]));
 sg13g2_antennanp ANTENNA_20 (.VDD(VPWR),
    .VSS(VGND),
    .A(FrameData[26]));
 sg13g2_antennanp ANTENNA_21 (.VDD(VPWR),
    .VSS(VGND),
    .A(FrameData[27]));
 sg13g2_antennanp ANTENNA_22 (.VDD(VPWR),
    .VSS(VGND),
    .A(FrameData[24]));
 sg13g2_antennanp ANTENNA_23 (.VDD(VPWR),
    .VSS(VGND),
    .A(FrameData[25]));
 sg13g2_antennanp ANTENNA_24 (.VDD(VPWR),
    .VSS(VGND),
    .A(FrameData[26]));
 sg13g2_antennanp ANTENNA_25 (.VDD(VPWR),
    .VSS(VGND),
    .A(FrameData[27]));
 sg13g2_antennanp ANTENNA_26 (.VDD(VPWR),
    .VSS(VGND),
    .A(FrameData[24]));
 sg13g2_antennanp ANTENNA_27 (.VDD(VPWR),
    .VSS(VGND),
    .A(FrameData[25]));
 sg13g2_antennanp ANTENNA_28 (.VDD(VPWR),
    .VSS(VGND),
    .A(FrameData[26]));
 sg13g2_antennanp ANTENNA_29 (.VDD(VPWR),
    .VSS(VGND),
    .A(FrameData[27]));
 sg13g2_antennanp ANTENNA_30 (.VDD(VPWR),
    .VSS(VGND),
    .A(FrameData[24]));
 sg13g2_antennanp ANTENNA_31 (.VDD(VPWR),
    .VSS(VGND),
    .A(FrameData[25]));
 sg13g2_antennanp ANTENNA_32 (.VDD(VPWR),
    .VSS(VGND),
    .A(FrameData[26]));
 sg13g2_antennanp ANTENNA_33 (.VDD(VPWR),
    .VSS(VGND),
    .A(FrameData[27]));
 sg13g2_antennanp ANTENNA_34 (.VDD(VPWR),
    .VSS(VGND),
    .A(FrameData[24]));
 sg13g2_antennanp ANTENNA_35 (.VDD(VPWR),
    .VSS(VGND),
    .A(FrameData[25]));
 sg13g2_antennanp ANTENNA_36 (.VDD(VPWR),
    .VSS(VGND),
    .A(FrameData[26]));
 sg13g2_antennanp ANTENNA_37 (.VDD(VPWR),
    .VSS(VGND),
    .A(FrameData[27]));
 sg13g2_antennanp ANTENNA_38 (.VDD(VPWR),
    .VSS(VGND),
    .A(FrameData[24]));
 sg13g2_antennanp ANTENNA_39 (.VDD(VPWR),
    .VSS(VGND),
    .A(FrameData[25]));
 sg13g2_antennanp ANTENNA_40 (.VDD(VPWR),
    .VSS(VGND),
    .A(FrameData[26]));
 sg13g2_antennanp ANTENNA_41 (.VDD(VPWR),
    .VSS(VGND),
    .A(FrameData[27]));
 sg13g2_antennanp ANTENNA_42 (.VDD(VPWR),
    .VSS(VGND),
    .A(FrameData[24]));
 sg13g2_antennanp ANTENNA_43 (.VDD(VPWR),
    .VSS(VGND),
    .A(FrameData[25]));
 sg13g2_antennanp ANTENNA_44 (.VDD(VPWR),
    .VSS(VGND),
    .A(FrameData[26]));
 sg13g2_antennanp ANTENNA_45 (.VDD(VPWR),
    .VSS(VGND),
    .A(FrameData[27]));
 sg13g2_decap_8 FILLER_0_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_63 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_70 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_77 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_84 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_91 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_98 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_105 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_112 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_119 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_126 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_133 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_140 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_147 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_154 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_161 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_168 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_175 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_182 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_189 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_196 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_203 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_210 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_217 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_224 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_231 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_238 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_245 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_252 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_259 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_266 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_273 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_280 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_287 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_294 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_301 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_308 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_315 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_322 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_329 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_336 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_343 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_350 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_357 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_364 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_371 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_378 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_385 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_392 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_399 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_406 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_413 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_420 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_427 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_0_434 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_0_438 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_63 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_70 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_77 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_84 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_91 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_98 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_109 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_116 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_123 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_130 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_137 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_144 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_151 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_158 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_165 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_1_172 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_1_174 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_179 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_186 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_193 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_200 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_207 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_214 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_221 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_228 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_235 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_242 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_249 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_256 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_263 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_1_274 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_1_278 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_283 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_290 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_297 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_304 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_311 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_318 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_325 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_332 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_339 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_346 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_353 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_360 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_367 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_374 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_381 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_388 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_395 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_402 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_409 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_416 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_423 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_430 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_437 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_1_444 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_1_446 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_63 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_70 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_77 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_84 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_91 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_98 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_105 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_112 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_119 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_126 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_133 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_140 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_147 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_154 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_161 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_168 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_175 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_2_182 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_2_184 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_2_189 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_197 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_2_204 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_2_218 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_2_222 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_2_235 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_2_237 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_250 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_2_261 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_2_265 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_2_270 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_2_274 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_279 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_286 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_293 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_300 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_307 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_2_314 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_2_318 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_323 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_330 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_337 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_2_344 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_352 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_359 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_366 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_373 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_380 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_387 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_394 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_401 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_408 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_415 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_422 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_429 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_436 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_443 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_2_450 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_63 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_70 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_77 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_84 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_91 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_98 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_105 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_112 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_119 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_126 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_133 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_140 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_147 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_154 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_161 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_168 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_175 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_182 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_189 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_196 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_203 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_210 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_217 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_224 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_3_231 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_239 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_246 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_3_253 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_3_255 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_260 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_267 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_274 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_281 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_288 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_295 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_302 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_309 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_316 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_323 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_330 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_337 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_3_344 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_350 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_357 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_364 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_371 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_378 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_385 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_392 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_399 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_406 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_413 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_420 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_427 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_434 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_441 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_3_448 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_3_450 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_63 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_4_70 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_4_74 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_80 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_4_87 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_4_89 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_94 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_101 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_108 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_115 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_122 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_4_129 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_137 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_144 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_151 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_158 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_165 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_172 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_179 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_4_186 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_4_188 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_4_193 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_202 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_209 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_216 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_223 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_230 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_237 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_244 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_251 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_4_258 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_263 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_270 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_277 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_284 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_291 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_298 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_305 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_4_312 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_4_316 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_325 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_332 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_339 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_346 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_353 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_360 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_367 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_374 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_381 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_388 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_395 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_402 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_409 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_416 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_423 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_430 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_437 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_444 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_63 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_70 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_5_77 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_5_81 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_114 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_5_121 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_149 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_156 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_163 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_5_170 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_214 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_221 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_228 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_235 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_242 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_249 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_256 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_263 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_5_270 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_276 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_283 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_5_290 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_310 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_5_317 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_5_329 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_5_335 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_5_339 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_5_345 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_5_347 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_352 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_359 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_366 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_373 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_380 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_387 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_394 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_401 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_408 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_415 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_422 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_429 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_436 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_443 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_5_450 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_6_63 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_6_72 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_6_74 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_87 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_94 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_101 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_108 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_115 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_122 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_6_129 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_134 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_141 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_148 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_155 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_162 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_169 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_176 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_6_183 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_6_191 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_6_193 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_202 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_209 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_216 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_223 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_230 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_237 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_244 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_251 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_258 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_265 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_272 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_279 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_286 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_293 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_300 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_307 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_314 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_321 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_328 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_6_335 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_343 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_350 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_6_357 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_365 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_372 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_379 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_386 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_393 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_400 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_407 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_414 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_421 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_428 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_435 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_442 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_6_449 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_63 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_7_70 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_78 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_85 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_92 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_99 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_106 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_113 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_120 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_127 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_134 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_141 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_148 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_155 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_162 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_169 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_176 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_183 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_190 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_197 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_204 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_211 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_218 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_225 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_232 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_239 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_246 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_7_253 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_259 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_266 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_273 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_280 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_287 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_294 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_301 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_308 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_315 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_322 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_7_329 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_7_333 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_338 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_345 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_352 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_366 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_373 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_380 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_387 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_394 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_401 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_408 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_415 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_422 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_429 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_436 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_443 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_7_450 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_63 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_70 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_77 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_84 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_91 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_98 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_105 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_112 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_119 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_126 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_133 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_140 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_147 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_154 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_161 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_168 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_175 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_182 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_189 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_196 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_203 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_210 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_217 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_224 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_231 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_238 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_8_245 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_8_249 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_8_278 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_283 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_290 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_297 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_304 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_311 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_318 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_8_325 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_8_327 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_332 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_8_339 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_8_343 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_8_365 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_392 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_403 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_410 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_417 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_424 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_8_431 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_8_435 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_441 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_8_448 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_8_450 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_63 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_70 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_77 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_84 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_91 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_9_98 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_9_102 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_199 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_206 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_213 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_220 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_227 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_234 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_241 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_248 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_9_255 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_9_261 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_9_267 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_291 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_298 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_305 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_312 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_9_339 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_9_359 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_9_374 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_410 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_417 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_424 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_431 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_9_438 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_9_442 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_63 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_70 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_77 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_84 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_91 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_10_98 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_215 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_222 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_229 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_236 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_243 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_250 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_257 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_264 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_271 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_278 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_285 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_292 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_299 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_306 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_415 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_422 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_10_429 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_10_433 (.VDD(VPWR),
    .VSS(VGND));
 assign Co = net106;
endmodule
